
module memory_WIDTH8_SIZE16_LOGSIZE4 ( clk, data_in, data_out, addr, wr_en );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, N19, N20, N21, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N16), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N20), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n293), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n292), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n291), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n290), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n289), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n288), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n287), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n286), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n285), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n284), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n283), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n282), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n281), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n280), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n279), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n278), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n277), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n276), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n275), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n274), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n273), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n272), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n271), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n270), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n269), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n268), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n267), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n266), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n265), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n264), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n263), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n262), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n261), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n260), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n259), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n258), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n257), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n256), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n255), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n254), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n253), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n252), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n251), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n250), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n249), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n248), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n247), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n246), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n245), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n244), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n243), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n242), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n241), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n240), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n239), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n238), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n237), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n236), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n235), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n234), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n233), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n232), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n231), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n230), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n229), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n228), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n227), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n226), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n225), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n224), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n223), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n222), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n221), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n220), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n219), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n218), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n217), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n216), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n215), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n214), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n213), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n212), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n211), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n210), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n209), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n208), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n207), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n206), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n205), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n204), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n203), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n202), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n201), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n200), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n199), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n198), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n197), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n196), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n195), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n194), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n193), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n192), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n191), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n190), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n189), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n188), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n187), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n186), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n185), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n184), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n183), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n182), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n181), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n180), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n179), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n178), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n177), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n176), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n175), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n174), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n173), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n172), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n171), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n170), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n169), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n168), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n167), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n166), .CK(clk), .Q(\mem[0][0] ) );
  BUF_X1 U3 ( .A(N10), .Z(n399) );
  BUF_X1 U4 ( .A(N10), .Z(n400) );
  BUF_X1 U5 ( .A(N10), .Z(n401) );
  BUF_X1 U6 ( .A(N10), .Z(n402) );
  BUF_X1 U7 ( .A(N10), .Z(n403) );
  BUF_X1 U8 ( .A(N11), .Z(n396) );
  BUF_X1 U9 ( .A(N11), .Z(n397) );
  BUF_X1 U10 ( .A(N11), .Z(n395) );
  NAND2_X1 U11 ( .A1(n42), .A2(n22), .ZN(n33) );
  NAND2_X1 U12 ( .A1(n42), .A2(n32), .ZN(n43) );
  NAND2_X1 U13 ( .A1(n21), .A2(n22), .ZN(n12) );
  NAND2_X1 U14 ( .A1(n32), .A2(n21), .ZN(n23) );
  NAND2_X1 U15 ( .A1(n100), .A2(n21), .ZN(n91) );
  NAND2_X1 U16 ( .A1(n110), .A2(n21), .ZN(n101) );
  NAND2_X1 U17 ( .A1(n100), .A2(n42), .ZN(n111) );
  NAND2_X1 U18 ( .A1(n110), .A2(n42), .ZN(n120) );
  NAND2_X1 U19 ( .A1(n61), .A2(n22), .ZN(n52) );
  NAND2_X1 U20 ( .A1(n61), .A2(n32), .ZN(n62) );
  NAND2_X1 U21 ( .A1(n80), .A2(n22), .ZN(n71) );
  NAND2_X1 U22 ( .A1(n80), .A2(n32), .ZN(n82) );
  NAND2_X1 U23 ( .A1(n100), .A2(n61), .ZN(n129) );
  NAND2_X1 U24 ( .A1(n110), .A2(n61), .ZN(n138) );
  NAND2_X1 U25 ( .A1(n100), .A2(n80), .ZN(n147) );
  NAND2_X1 U26 ( .A1(n110), .A2(n80), .ZN(n157) );
  AND2_X1 U27 ( .A1(n156), .A2(N10), .ZN(n110) );
  AND2_X1 U28 ( .A1(n156), .A2(n404), .ZN(n100) );
  AND2_X1 U29 ( .A1(N10), .A2(n81), .ZN(n32) );
  AND2_X1 U30 ( .A1(n81), .A2(n404), .ZN(n22) );
  NOR2_X1 U31 ( .A1(N11), .A2(N12), .ZN(n21) );
  NOR2_X1 U32 ( .A1(n405), .A2(N12), .ZN(n42) );
  AND2_X1 U33 ( .A1(N12), .A2(n405), .ZN(n61) );
  AND2_X1 U34 ( .A1(N12), .A2(N11), .ZN(n80) );
  OAI21_X1 U35 ( .B1(n12), .B2(n406), .A(n13), .ZN(n166) );
  NAND2_X1 U36 ( .A1(\mem[0][0] ), .A2(n12), .ZN(n13) );
  OAI21_X1 U37 ( .B1(n12), .B2(n407), .A(n14), .ZN(n167) );
  NAND2_X1 U38 ( .A1(\mem[0][1] ), .A2(n12), .ZN(n14) );
  OAI21_X1 U39 ( .B1(n12), .B2(n408), .A(n15), .ZN(n168) );
  NAND2_X1 U40 ( .A1(\mem[0][2] ), .A2(n12), .ZN(n15) );
  OAI21_X1 U41 ( .B1(n12), .B2(n409), .A(n16), .ZN(n169) );
  NAND2_X1 U42 ( .A1(\mem[0][3] ), .A2(n12), .ZN(n16) );
  OAI21_X1 U43 ( .B1(n12), .B2(n410), .A(n17), .ZN(n170) );
  NAND2_X1 U44 ( .A1(\mem[0][4] ), .A2(n12), .ZN(n17) );
  OAI21_X1 U45 ( .B1(n12), .B2(n411), .A(n18), .ZN(n171) );
  NAND2_X1 U46 ( .A1(\mem[0][5] ), .A2(n12), .ZN(n18) );
  OAI21_X1 U47 ( .B1(n12), .B2(n412), .A(n19), .ZN(n172) );
  NAND2_X1 U48 ( .A1(\mem[0][6] ), .A2(n12), .ZN(n19) );
  OAI21_X1 U49 ( .B1(n12), .B2(n413), .A(n20), .ZN(n173) );
  NAND2_X1 U50 ( .A1(\mem[0][7] ), .A2(n12), .ZN(n20) );
  OAI21_X1 U51 ( .B1(n406), .B2(n33), .A(n34), .ZN(n182) );
  NAND2_X1 U52 ( .A1(\mem[2][0] ), .A2(n33), .ZN(n34) );
  OAI21_X1 U53 ( .B1(n407), .B2(n33), .A(n35), .ZN(n183) );
  NAND2_X1 U54 ( .A1(\mem[2][1] ), .A2(n33), .ZN(n35) );
  OAI21_X1 U55 ( .B1(n408), .B2(n33), .A(n36), .ZN(n184) );
  NAND2_X1 U56 ( .A1(\mem[2][2] ), .A2(n33), .ZN(n36) );
  OAI21_X1 U57 ( .B1(n409), .B2(n33), .A(n37), .ZN(n185) );
  NAND2_X1 U58 ( .A1(\mem[2][3] ), .A2(n33), .ZN(n37) );
  OAI21_X1 U59 ( .B1(n410), .B2(n33), .A(n38), .ZN(n186) );
  NAND2_X1 U60 ( .A1(\mem[2][4] ), .A2(n33), .ZN(n38) );
  OAI21_X1 U61 ( .B1(n411), .B2(n33), .A(n39), .ZN(n187) );
  NAND2_X1 U62 ( .A1(\mem[2][5] ), .A2(n33), .ZN(n39) );
  OAI21_X1 U63 ( .B1(n412), .B2(n33), .A(n40), .ZN(n188) );
  NAND2_X1 U64 ( .A1(\mem[2][6] ), .A2(n33), .ZN(n40) );
  OAI21_X1 U65 ( .B1(n413), .B2(n33), .A(n41), .ZN(n189) );
  NAND2_X1 U66 ( .A1(\mem[2][7] ), .A2(n33), .ZN(n41) );
  OAI21_X1 U67 ( .B1(n406), .B2(n43), .A(n44), .ZN(n190) );
  NAND2_X1 U68 ( .A1(\mem[3][0] ), .A2(n43), .ZN(n44) );
  OAI21_X1 U69 ( .B1(n407), .B2(n43), .A(n45), .ZN(n191) );
  NAND2_X1 U70 ( .A1(\mem[3][1] ), .A2(n43), .ZN(n45) );
  OAI21_X1 U71 ( .B1(n408), .B2(n43), .A(n46), .ZN(n192) );
  NAND2_X1 U72 ( .A1(\mem[3][2] ), .A2(n43), .ZN(n46) );
  OAI21_X1 U73 ( .B1(n409), .B2(n43), .A(n47), .ZN(n193) );
  NAND2_X1 U74 ( .A1(\mem[3][3] ), .A2(n43), .ZN(n47) );
  OAI21_X1 U75 ( .B1(n410), .B2(n43), .A(n48), .ZN(n194) );
  NAND2_X1 U76 ( .A1(\mem[3][4] ), .A2(n43), .ZN(n48) );
  OAI21_X1 U77 ( .B1(n411), .B2(n43), .A(n49), .ZN(n195) );
  NAND2_X1 U78 ( .A1(\mem[3][5] ), .A2(n43), .ZN(n49) );
  OAI21_X1 U79 ( .B1(n412), .B2(n43), .A(n50), .ZN(n196) );
  NAND2_X1 U80 ( .A1(\mem[3][6] ), .A2(n43), .ZN(n50) );
  OAI21_X1 U81 ( .B1(n413), .B2(n43), .A(n51), .ZN(n197) );
  NAND2_X1 U82 ( .A1(\mem[3][7] ), .A2(n43), .ZN(n51) );
  NOR2_X1 U83 ( .A1(n414), .A2(N13), .ZN(n81) );
  INV_X1 U84 ( .A(wr_en), .ZN(n414) );
  OAI21_X1 U85 ( .B1(n406), .B2(n23), .A(n24), .ZN(n174) );
  NAND2_X1 U86 ( .A1(\mem[1][0] ), .A2(n23), .ZN(n24) );
  OAI21_X1 U87 ( .B1(n407), .B2(n23), .A(n25), .ZN(n175) );
  NAND2_X1 U88 ( .A1(\mem[1][1] ), .A2(n23), .ZN(n25) );
  OAI21_X1 U89 ( .B1(n408), .B2(n23), .A(n26), .ZN(n176) );
  NAND2_X1 U90 ( .A1(\mem[1][2] ), .A2(n23), .ZN(n26) );
  OAI21_X1 U91 ( .B1(n409), .B2(n23), .A(n27), .ZN(n177) );
  NAND2_X1 U92 ( .A1(\mem[1][3] ), .A2(n23), .ZN(n27) );
  OAI21_X1 U93 ( .B1(n410), .B2(n23), .A(n28), .ZN(n178) );
  NAND2_X1 U94 ( .A1(\mem[1][4] ), .A2(n23), .ZN(n28) );
  OAI21_X1 U95 ( .B1(n411), .B2(n23), .A(n29), .ZN(n179) );
  NAND2_X1 U96 ( .A1(\mem[1][5] ), .A2(n23), .ZN(n29) );
  OAI21_X1 U97 ( .B1(n412), .B2(n23), .A(n30), .ZN(n180) );
  NAND2_X1 U98 ( .A1(\mem[1][6] ), .A2(n23), .ZN(n30) );
  OAI21_X1 U99 ( .B1(n413), .B2(n23), .A(n31), .ZN(n181) );
  NAND2_X1 U100 ( .A1(\mem[1][7] ), .A2(n23), .ZN(n31) );
  OAI21_X1 U101 ( .B1(n406), .B2(n91), .A(n92), .ZN(n230) );
  NAND2_X1 U102 ( .A1(\mem[8][0] ), .A2(n91), .ZN(n92) );
  OAI21_X1 U103 ( .B1(n407), .B2(n91), .A(n93), .ZN(n231) );
  NAND2_X1 U104 ( .A1(\mem[8][1] ), .A2(n91), .ZN(n93) );
  OAI21_X1 U105 ( .B1(n408), .B2(n91), .A(n94), .ZN(n232) );
  NAND2_X1 U106 ( .A1(\mem[8][2] ), .A2(n91), .ZN(n94) );
  OAI21_X1 U107 ( .B1(n409), .B2(n91), .A(n95), .ZN(n233) );
  NAND2_X1 U108 ( .A1(\mem[8][3] ), .A2(n91), .ZN(n95) );
  OAI21_X1 U109 ( .B1(n410), .B2(n91), .A(n96), .ZN(n234) );
  NAND2_X1 U110 ( .A1(\mem[8][4] ), .A2(n91), .ZN(n96) );
  OAI21_X1 U111 ( .B1(n411), .B2(n91), .A(n97), .ZN(n235) );
  NAND2_X1 U112 ( .A1(\mem[8][5] ), .A2(n91), .ZN(n97) );
  OAI21_X1 U113 ( .B1(n412), .B2(n91), .A(n98), .ZN(n236) );
  NAND2_X1 U114 ( .A1(\mem[8][6] ), .A2(n91), .ZN(n98) );
  OAI21_X1 U115 ( .B1(n413), .B2(n91), .A(n99), .ZN(n237) );
  NAND2_X1 U116 ( .A1(\mem[8][7] ), .A2(n91), .ZN(n99) );
  OAI21_X1 U117 ( .B1(n406), .B2(n101), .A(n102), .ZN(n238) );
  NAND2_X1 U118 ( .A1(\mem[9][0] ), .A2(n101), .ZN(n102) );
  OAI21_X1 U119 ( .B1(n407), .B2(n101), .A(n103), .ZN(n239) );
  NAND2_X1 U120 ( .A1(\mem[9][1] ), .A2(n101), .ZN(n103) );
  OAI21_X1 U121 ( .B1(n408), .B2(n101), .A(n104), .ZN(n240) );
  NAND2_X1 U122 ( .A1(\mem[9][2] ), .A2(n101), .ZN(n104) );
  OAI21_X1 U123 ( .B1(n409), .B2(n101), .A(n105), .ZN(n241) );
  NAND2_X1 U124 ( .A1(\mem[9][3] ), .A2(n101), .ZN(n105) );
  OAI21_X1 U125 ( .B1(n410), .B2(n101), .A(n106), .ZN(n242) );
  NAND2_X1 U126 ( .A1(\mem[9][4] ), .A2(n101), .ZN(n106) );
  OAI21_X1 U127 ( .B1(n411), .B2(n101), .A(n107), .ZN(n243) );
  NAND2_X1 U128 ( .A1(\mem[9][5] ), .A2(n101), .ZN(n107) );
  OAI21_X1 U129 ( .B1(n412), .B2(n101), .A(n108), .ZN(n244) );
  NAND2_X1 U130 ( .A1(\mem[9][6] ), .A2(n101), .ZN(n108) );
  OAI21_X1 U131 ( .B1(n413), .B2(n101), .A(n109), .ZN(n245) );
  NAND2_X1 U132 ( .A1(\mem[9][7] ), .A2(n101), .ZN(n109) );
  OAI21_X1 U133 ( .B1(n406), .B2(n111), .A(n112), .ZN(n246) );
  NAND2_X1 U134 ( .A1(\mem[10][0] ), .A2(n111), .ZN(n112) );
  OAI21_X1 U135 ( .B1(n407), .B2(n111), .A(n113), .ZN(n247) );
  NAND2_X1 U136 ( .A1(\mem[10][1] ), .A2(n111), .ZN(n113) );
  OAI21_X1 U137 ( .B1(n408), .B2(n111), .A(n114), .ZN(n248) );
  NAND2_X1 U138 ( .A1(\mem[10][2] ), .A2(n111), .ZN(n114) );
  OAI21_X1 U139 ( .B1(n409), .B2(n111), .A(n115), .ZN(n249) );
  NAND2_X1 U140 ( .A1(\mem[10][3] ), .A2(n111), .ZN(n115) );
  OAI21_X1 U141 ( .B1(n410), .B2(n111), .A(n116), .ZN(n250) );
  NAND2_X1 U142 ( .A1(\mem[10][4] ), .A2(n111), .ZN(n116) );
  OAI21_X1 U143 ( .B1(n411), .B2(n111), .A(n117), .ZN(n251) );
  NAND2_X1 U144 ( .A1(\mem[10][5] ), .A2(n111), .ZN(n117) );
  OAI21_X1 U145 ( .B1(n412), .B2(n111), .A(n118), .ZN(n252) );
  NAND2_X1 U146 ( .A1(\mem[10][6] ), .A2(n111), .ZN(n118) );
  OAI21_X1 U147 ( .B1(n413), .B2(n111), .A(n119), .ZN(n253) );
  NAND2_X1 U148 ( .A1(\mem[10][7] ), .A2(n111), .ZN(n119) );
  OAI21_X1 U149 ( .B1(n406), .B2(n120), .A(n121), .ZN(n254) );
  NAND2_X1 U150 ( .A1(\mem[11][0] ), .A2(n120), .ZN(n121) );
  OAI21_X1 U151 ( .B1(n407), .B2(n120), .A(n122), .ZN(n255) );
  NAND2_X1 U152 ( .A1(\mem[11][1] ), .A2(n120), .ZN(n122) );
  OAI21_X1 U153 ( .B1(n408), .B2(n120), .A(n123), .ZN(n256) );
  NAND2_X1 U154 ( .A1(\mem[11][2] ), .A2(n120), .ZN(n123) );
  OAI21_X1 U155 ( .B1(n409), .B2(n120), .A(n124), .ZN(n257) );
  NAND2_X1 U156 ( .A1(\mem[11][3] ), .A2(n120), .ZN(n124) );
  OAI21_X1 U157 ( .B1(n410), .B2(n120), .A(n125), .ZN(n258) );
  NAND2_X1 U158 ( .A1(\mem[11][4] ), .A2(n120), .ZN(n125) );
  OAI21_X1 U159 ( .B1(n411), .B2(n120), .A(n126), .ZN(n259) );
  NAND2_X1 U160 ( .A1(\mem[11][5] ), .A2(n120), .ZN(n126) );
  OAI21_X1 U161 ( .B1(n412), .B2(n120), .A(n127), .ZN(n260) );
  NAND2_X1 U162 ( .A1(\mem[11][6] ), .A2(n120), .ZN(n127) );
  OAI21_X1 U163 ( .B1(n413), .B2(n120), .A(n128), .ZN(n261) );
  NAND2_X1 U164 ( .A1(\mem[11][7] ), .A2(n120), .ZN(n128) );
  OAI21_X1 U165 ( .B1(n406), .B2(n52), .A(n53), .ZN(n198) );
  NAND2_X1 U166 ( .A1(\mem[4][0] ), .A2(n52), .ZN(n53) );
  OAI21_X1 U167 ( .B1(n407), .B2(n52), .A(n54), .ZN(n199) );
  NAND2_X1 U168 ( .A1(\mem[4][1] ), .A2(n52), .ZN(n54) );
  OAI21_X1 U169 ( .B1(n408), .B2(n52), .A(n55), .ZN(n200) );
  NAND2_X1 U170 ( .A1(\mem[4][2] ), .A2(n52), .ZN(n55) );
  OAI21_X1 U171 ( .B1(n409), .B2(n52), .A(n56), .ZN(n201) );
  NAND2_X1 U172 ( .A1(\mem[4][3] ), .A2(n52), .ZN(n56) );
  OAI21_X1 U173 ( .B1(n410), .B2(n52), .A(n57), .ZN(n202) );
  NAND2_X1 U174 ( .A1(\mem[4][4] ), .A2(n52), .ZN(n57) );
  OAI21_X1 U175 ( .B1(n411), .B2(n52), .A(n58), .ZN(n203) );
  NAND2_X1 U176 ( .A1(\mem[4][5] ), .A2(n52), .ZN(n58) );
  OAI21_X1 U177 ( .B1(n412), .B2(n52), .A(n59), .ZN(n204) );
  NAND2_X1 U178 ( .A1(\mem[4][6] ), .A2(n52), .ZN(n59) );
  OAI21_X1 U179 ( .B1(n413), .B2(n52), .A(n60), .ZN(n205) );
  NAND2_X1 U180 ( .A1(\mem[4][7] ), .A2(n52), .ZN(n60) );
  OAI21_X1 U181 ( .B1(n406), .B2(n62), .A(n63), .ZN(n206) );
  NAND2_X1 U182 ( .A1(\mem[5][0] ), .A2(n62), .ZN(n63) );
  OAI21_X1 U183 ( .B1(n407), .B2(n62), .A(n64), .ZN(n207) );
  NAND2_X1 U184 ( .A1(\mem[5][1] ), .A2(n62), .ZN(n64) );
  OAI21_X1 U185 ( .B1(n408), .B2(n62), .A(n65), .ZN(n208) );
  NAND2_X1 U186 ( .A1(\mem[5][2] ), .A2(n62), .ZN(n65) );
  OAI21_X1 U187 ( .B1(n409), .B2(n62), .A(n66), .ZN(n209) );
  NAND2_X1 U188 ( .A1(\mem[5][3] ), .A2(n62), .ZN(n66) );
  OAI21_X1 U189 ( .B1(n410), .B2(n62), .A(n67), .ZN(n210) );
  NAND2_X1 U190 ( .A1(\mem[5][4] ), .A2(n62), .ZN(n67) );
  OAI21_X1 U191 ( .B1(n411), .B2(n62), .A(n68), .ZN(n211) );
  NAND2_X1 U192 ( .A1(\mem[5][5] ), .A2(n62), .ZN(n68) );
  OAI21_X1 U193 ( .B1(n412), .B2(n62), .A(n69), .ZN(n212) );
  NAND2_X1 U194 ( .A1(\mem[5][6] ), .A2(n62), .ZN(n69) );
  OAI21_X1 U195 ( .B1(n413), .B2(n62), .A(n70), .ZN(n213) );
  NAND2_X1 U196 ( .A1(\mem[5][7] ), .A2(n62), .ZN(n70) );
  OAI21_X1 U197 ( .B1(n406), .B2(n71), .A(n72), .ZN(n214) );
  NAND2_X1 U198 ( .A1(\mem[6][0] ), .A2(n71), .ZN(n72) );
  OAI21_X1 U199 ( .B1(n407), .B2(n71), .A(n73), .ZN(n215) );
  NAND2_X1 U200 ( .A1(\mem[6][1] ), .A2(n71), .ZN(n73) );
  OAI21_X1 U201 ( .B1(n408), .B2(n71), .A(n74), .ZN(n216) );
  NAND2_X1 U202 ( .A1(\mem[6][2] ), .A2(n71), .ZN(n74) );
  OAI21_X1 U203 ( .B1(n409), .B2(n71), .A(n75), .ZN(n217) );
  NAND2_X1 U204 ( .A1(\mem[6][3] ), .A2(n71), .ZN(n75) );
  OAI21_X1 U205 ( .B1(n410), .B2(n71), .A(n76), .ZN(n218) );
  NAND2_X1 U206 ( .A1(\mem[6][4] ), .A2(n71), .ZN(n76) );
  OAI21_X1 U207 ( .B1(n411), .B2(n71), .A(n77), .ZN(n219) );
  NAND2_X1 U208 ( .A1(\mem[6][5] ), .A2(n71), .ZN(n77) );
  OAI21_X1 U209 ( .B1(n412), .B2(n71), .A(n78), .ZN(n220) );
  NAND2_X1 U210 ( .A1(\mem[6][6] ), .A2(n71), .ZN(n78) );
  OAI21_X1 U211 ( .B1(n413), .B2(n71), .A(n79), .ZN(n221) );
  NAND2_X1 U212 ( .A1(\mem[6][7] ), .A2(n71), .ZN(n79) );
  OAI21_X1 U213 ( .B1(n406), .B2(n82), .A(n83), .ZN(n222) );
  NAND2_X1 U214 ( .A1(\mem[7][0] ), .A2(n82), .ZN(n83) );
  OAI21_X1 U215 ( .B1(n407), .B2(n82), .A(n84), .ZN(n223) );
  NAND2_X1 U216 ( .A1(\mem[7][1] ), .A2(n82), .ZN(n84) );
  OAI21_X1 U217 ( .B1(n408), .B2(n82), .A(n85), .ZN(n224) );
  NAND2_X1 U218 ( .A1(\mem[7][2] ), .A2(n82), .ZN(n85) );
  OAI21_X1 U219 ( .B1(n409), .B2(n82), .A(n86), .ZN(n225) );
  NAND2_X1 U220 ( .A1(\mem[7][3] ), .A2(n82), .ZN(n86) );
  OAI21_X1 U221 ( .B1(n410), .B2(n82), .A(n87), .ZN(n226) );
  NAND2_X1 U222 ( .A1(\mem[7][4] ), .A2(n82), .ZN(n87) );
  OAI21_X1 U223 ( .B1(n411), .B2(n82), .A(n88), .ZN(n227) );
  NAND2_X1 U224 ( .A1(\mem[7][5] ), .A2(n82), .ZN(n88) );
  OAI21_X1 U225 ( .B1(n412), .B2(n82), .A(n89), .ZN(n228) );
  NAND2_X1 U226 ( .A1(\mem[7][6] ), .A2(n82), .ZN(n89) );
  OAI21_X1 U227 ( .B1(n413), .B2(n82), .A(n90), .ZN(n229) );
  NAND2_X1 U228 ( .A1(\mem[7][7] ), .A2(n82), .ZN(n90) );
  OAI21_X1 U229 ( .B1(n406), .B2(n138), .A(n139), .ZN(n270) );
  NAND2_X1 U230 ( .A1(\mem[13][0] ), .A2(n138), .ZN(n139) );
  OAI21_X1 U231 ( .B1(n407), .B2(n138), .A(n140), .ZN(n271) );
  NAND2_X1 U232 ( .A1(\mem[13][1] ), .A2(n138), .ZN(n140) );
  OAI21_X1 U233 ( .B1(n408), .B2(n138), .A(n141), .ZN(n272) );
  NAND2_X1 U234 ( .A1(\mem[13][2] ), .A2(n138), .ZN(n141) );
  OAI21_X1 U235 ( .B1(n409), .B2(n138), .A(n142), .ZN(n273) );
  NAND2_X1 U236 ( .A1(\mem[13][3] ), .A2(n138), .ZN(n142) );
  OAI21_X1 U237 ( .B1(n410), .B2(n138), .A(n143), .ZN(n274) );
  NAND2_X1 U238 ( .A1(\mem[13][4] ), .A2(n138), .ZN(n143) );
  OAI21_X1 U239 ( .B1(n411), .B2(n138), .A(n144), .ZN(n275) );
  NAND2_X1 U240 ( .A1(\mem[13][5] ), .A2(n138), .ZN(n144) );
  OAI21_X1 U241 ( .B1(n412), .B2(n138), .A(n145), .ZN(n276) );
  NAND2_X1 U242 ( .A1(\mem[13][6] ), .A2(n138), .ZN(n145) );
  OAI21_X1 U243 ( .B1(n413), .B2(n138), .A(n146), .ZN(n277) );
  NAND2_X1 U244 ( .A1(\mem[13][7] ), .A2(n138), .ZN(n146) );
  OAI21_X1 U245 ( .B1(n406), .B2(n157), .A(n158), .ZN(n286) );
  NAND2_X1 U246 ( .A1(\mem[15][0] ), .A2(n157), .ZN(n158) );
  OAI21_X1 U247 ( .B1(n407), .B2(n157), .A(n159), .ZN(n287) );
  NAND2_X1 U248 ( .A1(\mem[15][1] ), .A2(n157), .ZN(n159) );
  OAI21_X1 U249 ( .B1(n408), .B2(n157), .A(n160), .ZN(n288) );
  NAND2_X1 U250 ( .A1(\mem[15][2] ), .A2(n157), .ZN(n160) );
  OAI21_X1 U251 ( .B1(n409), .B2(n157), .A(n161), .ZN(n289) );
  NAND2_X1 U252 ( .A1(\mem[15][3] ), .A2(n157), .ZN(n161) );
  OAI21_X1 U253 ( .B1(n410), .B2(n157), .A(n162), .ZN(n290) );
  NAND2_X1 U254 ( .A1(\mem[15][4] ), .A2(n157), .ZN(n162) );
  OAI21_X1 U255 ( .B1(n411), .B2(n157), .A(n163), .ZN(n291) );
  NAND2_X1 U256 ( .A1(\mem[15][5] ), .A2(n157), .ZN(n163) );
  OAI21_X1 U257 ( .B1(n412), .B2(n157), .A(n164), .ZN(n292) );
  NAND2_X1 U258 ( .A1(\mem[15][6] ), .A2(n157), .ZN(n164) );
  OAI21_X1 U259 ( .B1(n413), .B2(n157), .A(n165), .ZN(n293) );
  NAND2_X1 U260 ( .A1(\mem[15][7] ), .A2(n157), .ZN(n165) );
  OAI21_X1 U261 ( .B1(n406), .B2(n129), .A(n130), .ZN(n262) );
  NAND2_X1 U262 ( .A1(\mem[12][0] ), .A2(n129), .ZN(n130) );
  OAI21_X1 U263 ( .B1(n407), .B2(n129), .A(n131), .ZN(n263) );
  NAND2_X1 U264 ( .A1(\mem[12][1] ), .A2(n129), .ZN(n131) );
  OAI21_X1 U265 ( .B1(n408), .B2(n129), .A(n132), .ZN(n264) );
  NAND2_X1 U266 ( .A1(\mem[12][2] ), .A2(n129), .ZN(n132) );
  OAI21_X1 U267 ( .B1(n409), .B2(n129), .A(n133), .ZN(n265) );
  NAND2_X1 U268 ( .A1(\mem[12][3] ), .A2(n129), .ZN(n133) );
  OAI21_X1 U269 ( .B1(n410), .B2(n129), .A(n134), .ZN(n266) );
  NAND2_X1 U270 ( .A1(\mem[12][4] ), .A2(n129), .ZN(n134) );
  OAI21_X1 U271 ( .B1(n411), .B2(n129), .A(n135), .ZN(n267) );
  NAND2_X1 U272 ( .A1(\mem[12][5] ), .A2(n129), .ZN(n135) );
  OAI21_X1 U273 ( .B1(n412), .B2(n129), .A(n136), .ZN(n268) );
  NAND2_X1 U274 ( .A1(\mem[12][6] ), .A2(n129), .ZN(n136) );
  OAI21_X1 U275 ( .B1(n413), .B2(n129), .A(n137), .ZN(n269) );
  NAND2_X1 U276 ( .A1(\mem[12][7] ), .A2(n129), .ZN(n137) );
  OAI21_X1 U277 ( .B1(n406), .B2(n147), .A(n148), .ZN(n278) );
  NAND2_X1 U278 ( .A1(\mem[14][0] ), .A2(n147), .ZN(n148) );
  OAI21_X1 U279 ( .B1(n407), .B2(n147), .A(n149), .ZN(n279) );
  NAND2_X1 U280 ( .A1(\mem[14][1] ), .A2(n147), .ZN(n149) );
  OAI21_X1 U281 ( .B1(n408), .B2(n147), .A(n150), .ZN(n280) );
  NAND2_X1 U282 ( .A1(\mem[14][2] ), .A2(n147), .ZN(n150) );
  OAI21_X1 U283 ( .B1(n409), .B2(n147), .A(n151), .ZN(n281) );
  NAND2_X1 U284 ( .A1(\mem[14][3] ), .A2(n147), .ZN(n151) );
  OAI21_X1 U285 ( .B1(n410), .B2(n147), .A(n152), .ZN(n282) );
  NAND2_X1 U286 ( .A1(\mem[14][4] ), .A2(n147), .ZN(n152) );
  OAI21_X1 U287 ( .B1(n411), .B2(n147), .A(n153), .ZN(n283) );
  NAND2_X1 U288 ( .A1(\mem[14][5] ), .A2(n147), .ZN(n153) );
  OAI21_X1 U289 ( .B1(n412), .B2(n147), .A(n154), .ZN(n284) );
  NAND2_X1 U290 ( .A1(\mem[14][6] ), .A2(n147), .ZN(n154) );
  OAI21_X1 U291 ( .B1(n413), .B2(n147), .A(n155), .ZN(n285) );
  NAND2_X1 U292 ( .A1(\mem[14][7] ), .A2(n147), .ZN(n155) );
  AND2_X1 U293 ( .A1(N13), .A2(wr_en), .ZN(n156) );
  INV_X1 U294 ( .A(data_in[0]), .ZN(n406) );
  INV_X1 U295 ( .A(data_in[1]), .ZN(n407) );
  INV_X1 U296 ( .A(data_in[2]), .ZN(n408) );
  INV_X1 U297 ( .A(data_in[3]), .ZN(n409) );
  INV_X1 U298 ( .A(data_in[4]), .ZN(n410) );
  INV_X1 U299 ( .A(data_in[5]), .ZN(n411) );
  INV_X1 U300 ( .A(data_in[6]), .ZN(n412) );
  INV_X1 U301 ( .A(data_in[7]), .ZN(n413) );
  MUX2_X1 U302 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n398), .Z(n1) );
  MUX2_X1 U303 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n398), .Z(n2) );
  MUX2_X1 U304 ( .A(n2), .B(n1), .S(n395), .Z(n3) );
  MUX2_X1 U305 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n398), .Z(n4) );
  MUX2_X1 U306 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n398), .Z(n5) );
  MUX2_X1 U307 ( .A(n5), .B(n4), .S(n395), .Z(n6) );
  MUX2_X1 U308 ( .A(n6), .B(n3), .S(N12), .Z(n7) );
  MUX2_X1 U309 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n399), .Z(n8) );
  MUX2_X1 U310 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n399), .Z(n9) );
  MUX2_X1 U311 ( .A(n9), .B(n8), .S(n395), .Z(n10) );
  MUX2_X1 U312 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n399), .Z(n11) );
  MUX2_X1 U313 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n399), .Z(n294) );
  MUX2_X1 U314 ( .A(n294), .B(n11), .S(n395), .Z(n295) );
  MUX2_X1 U315 ( .A(n295), .B(n10), .S(N12), .Z(n296) );
  MUX2_X1 U316 ( .A(n296), .B(n7), .S(N13), .Z(N21) );
  MUX2_X1 U317 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n399), .Z(n297) );
  MUX2_X1 U318 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n399), .Z(n298) );
  MUX2_X1 U319 ( .A(n298), .B(n297), .S(n395), .Z(n299) );
  MUX2_X1 U320 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n399), .Z(n300) );
  MUX2_X1 U321 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n399), .Z(n301) );
  MUX2_X1 U322 ( .A(n301), .B(n300), .S(n395), .Z(n302) );
  MUX2_X1 U323 ( .A(n302), .B(n299), .S(N12), .Z(n303) );
  MUX2_X1 U324 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n399), .Z(n304) );
  MUX2_X1 U325 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n399), .Z(n305) );
  MUX2_X1 U326 ( .A(n305), .B(n304), .S(n395), .Z(n306) );
  MUX2_X1 U327 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n399), .Z(n307) );
  MUX2_X1 U328 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n399), .Z(n308) );
  MUX2_X1 U329 ( .A(n308), .B(n307), .S(n395), .Z(n309) );
  MUX2_X1 U330 ( .A(n309), .B(n306), .S(N12), .Z(n310) );
  MUX2_X1 U331 ( .A(n310), .B(n303), .S(N13), .Z(N20) );
  MUX2_X1 U332 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n400), .Z(n311) );
  MUX2_X1 U333 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n400), .Z(n312) );
  MUX2_X1 U334 ( .A(n312), .B(n311), .S(n396), .Z(n313) );
  MUX2_X1 U335 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n400), .Z(n314) );
  MUX2_X1 U336 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n400), .Z(n315) );
  MUX2_X1 U337 ( .A(n315), .B(n314), .S(n396), .Z(n316) );
  MUX2_X1 U338 ( .A(n316), .B(n313), .S(N12), .Z(n317) );
  MUX2_X1 U339 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n400), .Z(n318) );
  MUX2_X1 U340 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n400), .Z(n319) );
  MUX2_X1 U341 ( .A(n319), .B(n318), .S(n396), .Z(n320) );
  MUX2_X1 U342 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n400), .Z(n321) );
  MUX2_X1 U343 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n400), .Z(n322) );
  MUX2_X1 U344 ( .A(n322), .B(n321), .S(n396), .Z(n323) );
  MUX2_X1 U345 ( .A(n323), .B(n320), .S(N12), .Z(n324) );
  MUX2_X1 U346 ( .A(n324), .B(n317), .S(N13), .Z(N19) );
  MUX2_X1 U347 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n400), .Z(n325) );
  MUX2_X1 U348 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n400), .Z(n326) );
  MUX2_X1 U349 ( .A(n326), .B(n325), .S(n396), .Z(n327) );
  MUX2_X1 U350 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n400), .Z(n328) );
  MUX2_X1 U351 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n400), .Z(n329) );
  MUX2_X1 U352 ( .A(n329), .B(n328), .S(n396), .Z(n330) );
  MUX2_X1 U353 ( .A(n330), .B(n327), .S(N12), .Z(n331) );
  MUX2_X1 U354 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n401), .Z(n332) );
  MUX2_X1 U355 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n401), .Z(n333) );
  MUX2_X1 U356 ( .A(n333), .B(n332), .S(n396), .Z(n334) );
  MUX2_X1 U357 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n401), .Z(n335) );
  MUX2_X1 U358 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n401), .Z(n336) );
  MUX2_X1 U359 ( .A(n336), .B(n335), .S(n396), .Z(n337) );
  MUX2_X1 U360 ( .A(n337), .B(n334), .S(N12), .Z(n338) );
  MUX2_X1 U361 ( .A(n338), .B(n331), .S(N13), .Z(N18) );
  MUX2_X1 U362 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n401), .Z(n339) );
  MUX2_X1 U363 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n401), .Z(n340) );
  MUX2_X1 U364 ( .A(n340), .B(n339), .S(n396), .Z(n341) );
  MUX2_X1 U365 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n401), .Z(n342) );
  MUX2_X1 U366 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n401), .Z(n343) );
  MUX2_X1 U367 ( .A(n343), .B(n342), .S(n396), .Z(n344) );
  MUX2_X1 U368 ( .A(n344), .B(n341), .S(N12), .Z(n345) );
  MUX2_X1 U369 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n401), .Z(n346) );
  MUX2_X1 U370 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n401), .Z(n347) );
  MUX2_X1 U371 ( .A(n347), .B(n346), .S(n396), .Z(n348) );
  MUX2_X1 U372 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n401), .Z(n349) );
  MUX2_X1 U373 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n401), .Z(n350) );
  MUX2_X1 U374 ( .A(n350), .B(n349), .S(n396), .Z(n351) );
  MUX2_X1 U375 ( .A(n351), .B(n348), .S(N12), .Z(n352) );
  MUX2_X1 U376 ( .A(n352), .B(n345), .S(N13), .Z(N17) );
  MUX2_X1 U377 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n402), .Z(n353) );
  MUX2_X1 U378 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n402), .Z(n354) );
  MUX2_X1 U379 ( .A(n354), .B(n353), .S(n397), .Z(n355) );
  MUX2_X1 U380 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n402), .Z(n356) );
  MUX2_X1 U381 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n402), .Z(n357) );
  MUX2_X1 U382 ( .A(n357), .B(n356), .S(n397), .Z(n358) );
  MUX2_X1 U383 ( .A(n358), .B(n355), .S(N12), .Z(n359) );
  MUX2_X1 U384 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n402), .Z(n360) );
  MUX2_X1 U385 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n402), .Z(n361) );
  MUX2_X1 U386 ( .A(n361), .B(n360), .S(n397), .Z(n362) );
  MUX2_X1 U387 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n402), .Z(n363) );
  MUX2_X1 U388 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n402), .Z(n364) );
  MUX2_X1 U389 ( .A(n364), .B(n363), .S(n397), .Z(n365) );
  MUX2_X1 U390 ( .A(n365), .B(n362), .S(N12), .Z(n366) );
  MUX2_X1 U391 ( .A(n366), .B(n359), .S(N13), .Z(N16) );
  MUX2_X1 U392 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n402), .Z(n367) );
  MUX2_X1 U393 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n402), .Z(n368) );
  MUX2_X1 U394 ( .A(n368), .B(n367), .S(n397), .Z(n369) );
  MUX2_X1 U395 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n402), .Z(n370) );
  MUX2_X1 U396 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n402), .Z(n371) );
  MUX2_X1 U397 ( .A(n371), .B(n370), .S(n397), .Z(n372) );
  MUX2_X1 U398 ( .A(n372), .B(n369), .S(N12), .Z(n373) );
  MUX2_X1 U399 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n403), .Z(n374) );
  MUX2_X1 U400 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n403), .Z(n375) );
  MUX2_X1 U401 ( .A(n375), .B(n374), .S(n397), .Z(n376) );
  MUX2_X1 U402 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n403), .Z(n377) );
  MUX2_X1 U403 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n403), .Z(n378) );
  MUX2_X1 U404 ( .A(n378), .B(n377), .S(n397), .Z(n379) );
  MUX2_X1 U405 ( .A(n379), .B(n376), .S(N12), .Z(n380) );
  MUX2_X1 U406 ( .A(n380), .B(n373), .S(N13), .Z(N15) );
  MUX2_X1 U407 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n403), .Z(n381) );
  MUX2_X1 U408 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n403), .Z(n382) );
  MUX2_X1 U409 ( .A(n382), .B(n381), .S(n397), .Z(n383) );
  MUX2_X1 U410 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n403), .Z(n384) );
  MUX2_X1 U411 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n403), .Z(n385) );
  MUX2_X1 U412 ( .A(n385), .B(n384), .S(n397), .Z(n386) );
  MUX2_X1 U413 ( .A(n386), .B(n383), .S(N12), .Z(n387) );
  MUX2_X1 U414 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n403), .Z(n388) );
  MUX2_X1 U415 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n403), .Z(n389) );
  MUX2_X1 U416 ( .A(n389), .B(n388), .S(n397), .Z(n390) );
  MUX2_X1 U417 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n403), .Z(n391) );
  MUX2_X1 U418 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n403), .Z(n392) );
  MUX2_X1 U419 ( .A(n392), .B(n391), .S(n397), .Z(n393) );
  MUX2_X1 U420 ( .A(n393), .B(n390), .S(N12), .Z(n394) );
  MUX2_X1 U421 ( .A(n394), .B(n387), .S(N13), .Z(N14) );
  CLKBUF_X1 U422 ( .A(N10), .Z(n398) );
  INV_X1 U423 ( .A(N10), .ZN(n404) );
  INV_X1 U424 ( .A(N11), .ZN(n405) );
endmodule


module memory_WIDTH8_SIZE256_LOGSIZE8 ( clk, data_in, data_out, addr, wr_en );
  input [7:0] data_in;
  output [7:0] data_out;
  input [7:0] addr;
  input clk, wr_en;
  wire   N18, N19, N20, N21, N22, N23, N24, N25, \mem[255][7] , \mem[255][6] ,
         \mem[255][5] , \mem[255][4] , \mem[255][3] , \mem[255][2] ,
         \mem[255][1] , \mem[255][0] , \mem[254][7] , \mem[254][6] ,
         \mem[254][5] , \mem[254][4] , \mem[254][3] , \mem[254][2] ,
         \mem[254][1] , \mem[254][0] , \mem[253][7] , \mem[253][6] ,
         \mem[253][5] , \mem[253][4] , \mem[253][3] , \mem[253][2] ,
         \mem[253][1] , \mem[253][0] , \mem[252][7] , \mem[252][6] ,
         \mem[252][5] , \mem[252][4] , \mem[252][3] , \mem[252][2] ,
         \mem[252][1] , \mem[252][0] , \mem[251][7] , \mem[251][6] ,
         \mem[251][5] , \mem[251][4] , \mem[251][3] , \mem[251][2] ,
         \mem[251][1] , \mem[251][0] , \mem[250][7] , \mem[250][6] ,
         \mem[250][5] , \mem[250][4] , \mem[250][3] , \mem[250][2] ,
         \mem[250][1] , \mem[250][0] , \mem[249][7] , \mem[249][6] ,
         \mem[249][5] , \mem[249][4] , \mem[249][3] , \mem[249][2] ,
         \mem[249][1] , \mem[249][0] , \mem[248][7] , \mem[248][6] ,
         \mem[248][5] , \mem[248][4] , \mem[248][3] , \mem[248][2] ,
         \mem[248][1] , \mem[248][0] , \mem[247][7] , \mem[247][6] ,
         \mem[247][5] , \mem[247][4] , \mem[247][3] , \mem[247][2] ,
         \mem[247][1] , \mem[247][0] , \mem[246][7] , \mem[246][6] ,
         \mem[246][5] , \mem[246][4] , \mem[246][3] , \mem[246][2] ,
         \mem[246][1] , \mem[246][0] , \mem[245][7] , \mem[245][6] ,
         \mem[245][5] , \mem[245][4] , \mem[245][3] , \mem[245][2] ,
         \mem[245][1] , \mem[245][0] , \mem[244][7] , \mem[244][6] ,
         \mem[244][5] , \mem[244][4] , \mem[244][3] , \mem[244][2] ,
         \mem[244][1] , \mem[244][0] , \mem[243][7] , \mem[243][6] ,
         \mem[243][5] , \mem[243][4] , \mem[243][3] , \mem[243][2] ,
         \mem[243][1] , \mem[243][0] , \mem[242][7] , \mem[242][6] ,
         \mem[242][5] , \mem[242][4] , \mem[242][3] , \mem[242][2] ,
         \mem[242][1] , \mem[242][0] , \mem[241][7] , \mem[241][6] ,
         \mem[241][5] , \mem[241][4] , \mem[241][3] , \mem[241][2] ,
         \mem[241][1] , \mem[241][0] , \mem[240][7] , \mem[240][6] ,
         \mem[240][5] , \mem[240][4] , \mem[240][3] , \mem[240][2] ,
         \mem[240][1] , \mem[240][0] , \mem[239][7] , \mem[239][6] ,
         \mem[239][5] , \mem[239][4] , \mem[239][3] , \mem[239][2] ,
         \mem[239][1] , \mem[239][0] , \mem[238][7] , \mem[238][6] ,
         \mem[238][5] , \mem[238][4] , \mem[238][3] , \mem[238][2] ,
         \mem[238][1] , \mem[238][0] , \mem[237][7] , \mem[237][6] ,
         \mem[237][5] , \mem[237][4] , \mem[237][3] , \mem[237][2] ,
         \mem[237][1] , \mem[237][0] , \mem[236][7] , \mem[236][6] ,
         \mem[236][5] , \mem[236][4] , \mem[236][3] , \mem[236][2] ,
         \mem[236][1] , \mem[236][0] , \mem[235][7] , \mem[235][6] ,
         \mem[235][5] , \mem[235][4] , \mem[235][3] , \mem[235][2] ,
         \mem[235][1] , \mem[235][0] , \mem[234][7] , \mem[234][6] ,
         \mem[234][5] , \mem[234][4] , \mem[234][3] , \mem[234][2] ,
         \mem[234][1] , \mem[234][0] , \mem[233][7] , \mem[233][6] ,
         \mem[233][5] , \mem[233][4] , \mem[233][3] , \mem[233][2] ,
         \mem[233][1] , \mem[233][0] , \mem[232][7] , \mem[232][6] ,
         \mem[232][5] , \mem[232][4] , \mem[232][3] , \mem[232][2] ,
         \mem[232][1] , \mem[232][0] , \mem[231][7] , \mem[231][6] ,
         \mem[231][5] , \mem[231][4] , \mem[231][3] , \mem[231][2] ,
         \mem[231][1] , \mem[231][0] , \mem[230][7] , \mem[230][6] ,
         \mem[230][5] , \mem[230][4] , \mem[230][3] , \mem[230][2] ,
         \mem[230][1] , \mem[230][0] , \mem[229][7] , \mem[229][6] ,
         \mem[229][5] , \mem[229][4] , \mem[229][3] , \mem[229][2] ,
         \mem[229][1] , \mem[229][0] , \mem[228][7] , \mem[228][6] ,
         \mem[228][5] , \mem[228][4] , \mem[228][3] , \mem[228][2] ,
         \mem[228][1] , \mem[228][0] , \mem[227][7] , \mem[227][6] ,
         \mem[227][5] , \mem[227][4] , \mem[227][3] , \mem[227][2] ,
         \mem[227][1] , \mem[227][0] , \mem[226][7] , \mem[226][6] ,
         \mem[226][5] , \mem[226][4] , \mem[226][3] , \mem[226][2] ,
         \mem[226][1] , \mem[226][0] , \mem[225][7] , \mem[225][6] ,
         \mem[225][5] , \mem[225][4] , \mem[225][3] , \mem[225][2] ,
         \mem[225][1] , \mem[225][0] , \mem[224][7] , \mem[224][6] ,
         \mem[224][5] , \mem[224][4] , \mem[224][3] , \mem[224][2] ,
         \mem[224][1] , \mem[224][0] , \mem[223][7] , \mem[223][6] ,
         \mem[223][5] , \mem[223][4] , \mem[223][3] , \mem[223][2] ,
         \mem[223][1] , \mem[223][0] , \mem[222][7] , \mem[222][6] ,
         \mem[222][5] , \mem[222][4] , \mem[222][3] , \mem[222][2] ,
         \mem[222][1] , \mem[222][0] , \mem[221][7] , \mem[221][6] ,
         \mem[221][5] , \mem[221][4] , \mem[221][3] , \mem[221][2] ,
         \mem[221][1] , \mem[221][0] , \mem[220][7] , \mem[220][6] ,
         \mem[220][5] , \mem[220][4] , \mem[220][3] , \mem[220][2] ,
         \mem[220][1] , \mem[220][0] , \mem[219][7] , \mem[219][6] ,
         \mem[219][5] , \mem[219][4] , \mem[219][3] , \mem[219][2] ,
         \mem[219][1] , \mem[219][0] , \mem[218][7] , \mem[218][6] ,
         \mem[218][5] , \mem[218][4] , \mem[218][3] , \mem[218][2] ,
         \mem[218][1] , \mem[218][0] , \mem[217][7] , \mem[217][6] ,
         \mem[217][5] , \mem[217][4] , \mem[217][3] , \mem[217][2] ,
         \mem[217][1] , \mem[217][0] , \mem[216][7] , \mem[216][6] ,
         \mem[216][5] , \mem[216][4] , \mem[216][3] , \mem[216][2] ,
         \mem[216][1] , \mem[216][0] , \mem[215][7] , \mem[215][6] ,
         \mem[215][5] , \mem[215][4] , \mem[215][3] , \mem[215][2] ,
         \mem[215][1] , \mem[215][0] , \mem[214][7] , \mem[214][6] ,
         \mem[214][5] , \mem[214][4] , \mem[214][3] , \mem[214][2] ,
         \mem[214][1] , \mem[214][0] , \mem[213][7] , \mem[213][6] ,
         \mem[213][5] , \mem[213][4] , \mem[213][3] , \mem[213][2] ,
         \mem[213][1] , \mem[213][0] , \mem[212][7] , \mem[212][6] ,
         \mem[212][5] , \mem[212][4] , \mem[212][3] , \mem[212][2] ,
         \mem[212][1] , \mem[212][0] , \mem[211][7] , \mem[211][6] ,
         \mem[211][5] , \mem[211][4] , \mem[211][3] , \mem[211][2] ,
         \mem[211][1] , \mem[211][0] , \mem[210][7] , \mem[210][6] ,
         \mem[210][5] , \mem[210][4] , \mem[210][3] , \mem[210][2] ,
         \mem[210][1] , \mem[210][0] , \mem[209][7] , \mem[209][6] ,
         \mem[209][5] , \mem[209][4] , \mem[209][3] , \mem[209][2] ,
         \mem[209][1] , \mem[209][0] , \mem[208][7] , \mem[208][6] ,
         \mem[208][5] , \mem[208][4] , \mem[208][3] , \mem[208][2] ,
         \mem[208][1] , \mem[208][0] , \mem[207][7] , \mem[207][6] ,
         \mem[207][5] , \mem[207][4] , \mem[207][3] , \mem[207][2] ,
         \mem[207][1] , \mem[207][0] , \mem[206][7] , \mem[206][6] ,
         \mem[206][5] , \mem[206][4] , \mem[206][3] , \mem[206][2] ,
         \mem[206][1] , \mem[206][0] , \mem[205][7] , \mem[205][6] ,
         \mem[205][5] , \mem[205][4] , \mem[205][3] , \mem[205][2] ,
         \mem[205][1] , \mem[205][0] , \mem[204][7] , \mem[204][6] ,
         \mem[204][5] , \mem[204][4] , \mem[204][3] , \mem[204][2] ,
         \mem[204][1] , \mem[204][0] , \mem[203][7] , \mem[203][6] ,
         \mem[203][5] , \mem[203][4] , \mem[203][3] , \mem[203][2] ,
         \mem[203][1] , \mem[203][0] , \mem[202][7] , \mem[202][6] ,
         \mem[202][5] , \mem[202][4] , \mem[202][3] , \mem[202][2] ,
         \mem[202][1] , \mem[202][0] , \mem[201][7] , \mem[201][6] ,
         \mem[201][5] , \mem[201][4] , \mem[201][3] , \mem[201][2] ,
         \mem[201][1] , \mem[201][0] , \mem[200][7] , \mem[200][6] ,
         \mem[200][5] , \mem[200][4] , \mem[200][3] , \mem[200][2] ,
         \mem[200][1] , \mem[200][0] , \mem[199][7] , \mem[199][6] ,
         \mem[199][5] , \mem[199][4] , \mem[199][3] , \mem[199][2] ,
         \mem[199][1] , \mem[199][0] , \mem[198][7] , \mem[198][6] ,
         \mem[198][5] , \mem[198][4] , \mem[198][3] , \mem[198][2] ,
         \mem[198][1] , \mem[198][0] , \mem[197][7] , \mem[197][6] ,
         \mem[197][5] , \mem[197][4] , \mem[197][3] , \mem[197][2] ,
         \mem[197][1] , \mem[197][0] , \mem[196][7] , \mem[196][6] ,
         \mem[196][5] , \mem[196][4] , \mem[196][3] , \mem[196][2] ,
         \mem[196][1] , \mem[196][0] , \mem[195][7] , \mem[195][6] ,
         \mem[195][5] , \mem[195][4] , \mem[195][3] , \mem[195][2] ,
         \mem[195][1] , \mem[195][0] , \mem[194][7] , \mem[194][6] ,
         \mem[194][5] , \mem[194][4] , \mem[194][3] , \mem[194][2] ,
         \mem[194][1] , \mem[194][0] , \mem[193][7] , \mem[193][6] ,
         \mem[193][5] , \mem[193][4] , \mem[193][3] , \mem[193][2] ,
         \mem[193][1] , \mem[193][0] , \mem[192][7] , \mem[192][6] ,
         \mem[192][5] , \mem[192][4] , \mem[192][3] , \mem[192][2] ,
         \mem[192][1] , \mem[192][0] , \mem[191][7] , \mem[191][6] ,
         \mem[191][5] , \mem[191][4] , \mem[191][3] , \mem[191][2] ,
         \mem[191][1] , \mem[191][0] , \mem[190][7] , \mem[190][6] ,
         \mem[190][5] , \mem[190][4] , \mem[190][3] , \mem[190][2] ,
         \mem[190][1] , \mem[190][0] , \mem[189][7] , \mem[189][6] ,
         \mem[189][5] , \mem[189][4] , \mem[189][3] , \mem[189][2] ,
         \mem[189][1] , \mem[189][0] , \mem[188][7] , \mem[188][6] ,
         \mem[188][5] , \mem[188][4] , \mem[188][3] , \mem[188][2] ,
         \mem[188][1] , \mem[188][0] , \mem[187][7] , \mem[187][6] ,
         \mem[187][5] , \mem[187][4] , \mem[187][3] , \mem[187][2] ,
         \mem[187][1] , \mem[187][0] , \mem[186][7] , \mem[186][6] ,
         \mem[186][5] , \mem[186][4] , \mem[186][3] , \mem[186][2] ,
         \mem[186][1] , \mem[186][0] , \mem[185][7] , \mem[185][6] ,
         \mem[185][5] , \mem[185][4] , \mem[185][3] , \mem[185][2] ,
         \mem[185][1] , \mem[185][0] , \mem[184][7] , \mem[184][6] ,
         \mem[184][5] , \mem[184][4] , \mem[184][3] , \mem[184][2] ,
         \mem[184][1] , \mem[184][0] , \mem[183][7] , \mem[183][6] ,
         \mem[183][5] , \mem[183][4] , \mem[183][3] , \mem[183][2] ,
         \mem[183][1] , \mem[183][0] , \mem[182][7] , \mem[182][6] ,
         \mem[182][5] , \mem[182][4] , \mem[182][3] , \mem[182][2] ,
         \mem[182][1] , \mem[182][0] , \mem[181][7] , \mem[181][6] ,
         \mem[181][5] , \mem[181][4] , \mem[181][3] , \mem[181][2] ,
         \mem[181][1] , \mem[181][0] , \mem[180][7] , \mem[180][6] ,
         \mem[180][5] , \mem[180][4] , \mem[180][3] , \mem[180][2] ,
         \mem[180][1] , \mem[180][0] , \mem[179][7] , \mem[179][6] ,
         \mem[179][5] , \mem[179][4] , \mem[179][3] , \mem[179][2] ,
         \mem[179][1] , \mem[179][0] , \mem[178][7] , \mem[178][6] ,
         \mem[178][5] , \mem[178][4] , \mem[178][3] , \mem[178][2] ,
         \mem[178][1] , \mem[178][0] , \mem[177][7] , \mem[177][6] ,
         \mem[177][5] , \mem[177][4] , \mem[177][3] , \mem[177][2] ,
         \mem[177][1] , \mem[177][0] , \mem[176][7] , \mem[176][6] ,
         \mem[176][5] , \mem[176][4] , \mem[176][3] , \mem[176][2] ,
         \mem[176][1] , \mem[176][0] , \mem[175][7] , \mem[175][6] ,
         \mem[175][5] , \mem[175][4] , \mem[175][3] , \mem[175][2] ,
         \mem[175][1] , \mem[175][0] , \mem[174][7] , \mem[174][6] ,
         \mem[174][5] , \mem[174][4] , \mem[174][3] , \mem[174][2] ,
         \mem[174][1] , \mem[174][0] , \mem[173][7] , \mem[173][6] ,
         \mem[173][5] , \mem[173][4] , \mem[173][3] , \mem[173][2] ,
         \mem[173][1] , \mem[173][0] , \mem[172][7] , \mem[172][6] ,
         \mem[172][5] , \mem[172][4] , \mem[172][3] , \mem[172][2] ,
         \mem[172][1] , \mem[172][0] , \mem[171][7] , \mem[171][6] ,
         \mem[171][5] , \mem[171][4] , \mem[171][3] , \mem[171][2] ,
         \mem[171][1] , \mem[171][0] , \mem[170][7] , \mem[170][6] ,
         \mem[170][5] , \mem[170][4] , \mem[170][3] , \mem[170][2] ,
         \mem[170][1] , \mem[170][0] , \mem[169][7] , \mem[169][6] ,
         \mem[169][5] , \mem[169][4] , \mem[169][3] , \mem[169][2] ,
         \mem[169][1] , \mem[169][0] , \mem[168][7] , \mem[168][6] ,
         \mem[168][5] , \mem[168][4] , \mem[168][3] , \mem[168][2] ,
         \mem[168][1] , \mem[168][0] , \mem[167][7] , \mem[167][6] ,
         \mem[167][5] , \mem[167][4] , \mem[167][3] , \mem[167][2] ,
         \mem[167][1] , \mem[167][0] , \mem[166][7] , \mem[166][6] ,
         \mem[166][5] , \mem[166][4] , \mem[166][3] , \mem[166][2] ,
         \mem[166][1] , \mem[166][0] , \mem[165][7] , \mem[165][6] ,
         \mem[165][5] , \mem[165][4] , \mem[165][3] , \mem[165][2] ,
         \mem[165][1] , \mem[165][0] , \mem[164][7] , \mem[164][6] ,
         \mem[164][5] , \mem[164][4] , \mem[164][3] , \mem[164][2] ,
         \mem[164][1] , \mem[164][0] , \mem[163][7] , \mem[163][6] ,
         \mem[163][5] , \mem[163][4] , \mem[163][3] , \mem[163][2] ,
         \mem[163][1] , \mem[163][0] , \mem[162][7] , \mem[162][6] ,
         \mem[162][5] , \mem[162][4] , \mem[162][3] , \mem[162][2] ,
         \mem[162][1] , \mem[162][0] , \mem[161][7] , \mem[161][6] ,
         \mem[161][5] , \mem[161][4] , \mem[161][3] , \mem[161][2] ,
         \mem[161][1] , \mem[161][0] , \mem[160][7] , \mem[160][6] ,
         \mem[160][5] , \mem[160][4] , \mem[160][3] , \mem[160][2] ,
         \mem[160][1] , \mem[160][0] , \mem[159][7] , \mem[159][6] ,
         \mem[159][5] , \mem[159][4] , \mem[159][3] , \mem[159][2] ,
         \mem[159][1] , \mem[159][0] , \mem[158][7] , \mem[158][6] ,
         \mem[158][5] , \mem[158][4] , \mem[158][3] , \mem[158][2] ,
         \mem[158][1] , \mem[158][0] , \mem[157][7] , \mem[157][6] ,
         \mem[157][5] , \mem[157][4] , \mem[157][3] , \mem[157][2] ,
         \mem[157][1] , \mem[157][0] , \mem[156][7] , \mem[156][6] ,
         \mem[156][5] , \mem[156][4] , \mem[156][3] , \mem[156][2] ,
         \mem[156][1] , \mem[156][0] , \mem[155][7] , \mem[155][6] ,
         \mem[155][5] , \mem[155][4] , \mem[155][3] , \mem[155][2] ,
         \mem[155][1] , \mem[155][0] , \mem[154][7] , \mem[154][6] ,
         \mem[154][5] , \mem[154][4] , \mem[154][3] , \mem[154][2] ,
         \mem[154][1] , \mem[154][0] , \mem[153][7] , \mem[153][6] ,
         \mem[153][5] , \mem[153][4] , \mem[153][3] , \mem[153][2] ,
         \mem[153][1] , \mem[153][0] , \mem[152][7] , \mem[152][6] ,
         \mem[152][5] , \mem[152][4] , \mem[152][3] , \mem[152][2] ,
         \mem[152][1] , \mem[152][0] , \mem[151][7] , \mem[151][6] ,
         \mem[151][5] , \mem[151][4] , \mem[151][3] , \mem[151][2] ,
         \mem[151][1] , \mem[151][0] , \mem[150][7] , \mem[150][6] ,
         \mem[150][5] , \mem[150][4] , \mem[150][3] , \mem[150][2] ,
         \mem[150][1] , \mem[150][0] , \mem[149][7] , \mem[149][6] ,
         \mem[149][5] , \mem[149][4] , \mem[149][3] , \mem[149][2] ,
         \mem[149][1] , \mem[149][0] , \mem[148][7] , \mem[148][6] ,
         \mem[148][5] , \mem[148][4] , \mem[148][3] , \mem[148][2] ,
         \mem[148][1] , \mem[148][0] , \mem[147][7] , \mem[147][6] ,
         \mem[147][5] , \mem[147][4] , \mem[147][3] , \mem[147][2] ,
         \mem[147][1] , \mem[147][0] , \mem[146][7] , \mem[146][6] ,
         \mem[146][5] , \mem[146][4] , \mem[146][3] , \mem[146][2] ,
         \mem[146][1] , \mem[146][0] , \mem[145][7] , \mem[145][6] ,
         \mem[145][5] , \mem[145][4] , \mem[145][3] , \mem[145][2] ,
         \mem[145][1] , \mem[145][0] , \mem[144][7] , \mem[144][6] ,
         \mem[144][5] , \mem[144][4] , \mem[144][3] , \mem[144][2] ,
         \mem[144][1] , \mem[144][0] , \mem[143][7] , \mem[143][6] ,
         \mem[143][5] , \mem[143][4] , \mem[143][3] , \mem[143][2] ,
         \mem[143][1] , \mem[143][0] , \mem[142][7] , \mem[142][6] ,
         \mem[142][5] , \mem[142][4] , \mem[142][3] , \mem[142][2] ,
         \mem[142][1] , \mem[142][0] , \mem[141][7] , \mem[141][6] ,
         \mem[141][5] , \mem[141][4] , \mem[141][3] , \mem[141][2] ,
         \mem[141][1] , \mem[141][0] , \mem[140][7] , \mem[140][6] ,
         \mem[140][5] , \mem[140][4] , \mem[140][3] , \mem[140][2] ,
         \mem[140][1] , \mem[140][0] , \mem[139][7] , \mem[139][6] ,
         \mem[139][5] , \mem[139][4] , \mem[139][3] , \mem[139][2] ,
         \mem[139][1] , \mem[139][0] , \mem[138][7] , \mem[138][6] ,
         \mem[138][5] , \mem[138][4] , \mem[138][3] , \mem[138][2] ,
         \mem[138][1] , \mem[138][0] , \mem[137][7] , \mem[137][6] ,
         \mem[137][5] , \mem[137][4] , \mem[137][3] , \mem[137][2] ,
         \mem[137][1] , \mem[137][0] , \mem[136][7] , \mem[136][6] ,
         \mem[136][5] , \mem[136][4] , \mem[136][3] , \mem[136][2] ,
         \mem[136][1] , \mem[136][0] , \mem[135][7] , \mem[135][6] ,
         \mem[135][5] , \mem[135][4] , \mem[135][3] , \mem[135][2] ,
         \mem[135][1] , \mem[135][0] , \mem[134][7] , \mem[134][6] ,
         \mem[134][5] , \mem[134][4] , \mem[134][3] , \mem[134][2] ,
         \mem[134][1] , \mem[134][0] , \mem[133][7] , \mem[133][6] ,
         \mem[133][5] , \mem[133][4] , \mem[133][3] , \mem[133][2] ,
         \mem[133][1] , \mem[133][0] , \mem[132][7] , \mem[132][6] ,
         \mem[132][5] , \mem[132][4] , \mem[132][3] , \mem[132][2] ,
         \mem[132][1] , \mem[132][0] , \mem[131][7] , \mem[131][6] ,
         \mem[131][5] , \mem[131][4] , \mem[131][3] , \mem[131][2] ,
         \mem[131][1] , \mem[131][0] , \mem[130][7] , \mem[130][6] ,
         \mem[130][5] , \mem[130][4] , \mem[130][3] , \mem[130][2] ,
         \mem[130][1] , \mem[130][0] , \mem[129][7] , \mem[129][6] ,
         \mem[129][5] , \mem[129][4] , \mem[129][3] , \mem[129][2] ,
         \mem[129][1] , \mem[129][0] , \mem[128][7] , \mem[128][6] ,
         \mem[128][5] , \mem[128][4] , \mem[128][3] , \mem[128][2] ,
         \mem[128][1] , \mem[128][0] , \mem[127][7] , \mem[127][6] ,
         \mem[127][5] , \mem[127][4] , \mem[127][3] , \mem[127][2] ,
         \mem[127][1] , \mem[127][0] , \mem[126][7] , \mem[126][6] ,
         \mem[126][5] , \mem[126][4] , \mem[126][3] , \mem[126][2] ,
         \mem[126][1] , \mem[126][0] , \mem[125][7] , \mem[125][6] ,
         \mem[125][5] , \mem[125][4] , \mem[125][3] , \mem[125][2] ,
         \mem[125][1] , \mem[125][0] , \mem[124][7] , \mem[124][6] ,
         \mem[124][5] , \mem[124][4] , \mem[124][3] , \mem[124][2] ,
         \mem[124][1] , \mem[124][0] , \mem[123][7] , \mem[123][6] ,
         \mem[123][5] , \mem[123][4] , \mem[123][3] , \mem[123][2] ,
         \mem[123][1] , \mem[123][0] , \mem[122][7] , \mem[122][6] ,
         \mem[122][5] , \mem[122][4] , \mem[122][3] , \mem[122][2] ,
         \mem[122][1] , \mem[122][0] , \mem[121][7] , \mem[121][6] ,
         \mem[121][5] , \mem[121][4] , \mem[121][3] , \mem[121][2] ,
         \mem[121][1] , \mem[121][0] , \mem[120][7] , \mem[120][6] ,
         \mem[120][5] , \mem[120][4] , \mem[120][3] , \mem[120][2] ,
         \mem[120][1] , \mem[120][0] , \mem[119][7] , \mem[119][6] ,
         \mem[119][5] , \mem[119][4] , \mem[119][3] , \mem[119][2] ,
         \mem[119][1] , \mem[119][0] , \mem[118][7] , \mem[118][6] ,
         \mem[118][5] , \mem[118][4] , \mem[118][3] , \mem[118][2] ,
         \mem[118][1] , \mem[118][0] , \mem[117][7] , \mem[117][6] ,
         \mem[117][5] , \mem[117][4] , \mem[117][3] , \mem[117][2] ,
         \mem[117][1] , \mem[117][0] , \mem[116][7] , \mem[116][6] ,
         \mem[116][5] , \mem[116][4] , \mem[116][3] , \mem[116][2] ,
         \mem[116][1] , \mem[116][0] , \mem[115][7] , \mem[115][6] ,
         \mem[115][5] , \mem[115][4] , \mem[115][3] , \mem[115][2] ,
         \mem[115][1] , \mem[115][0] , \mem[114][7] , \mem[114][6] ,
         \mem[114][5] , \mem[114][4] , \mem[114][3] , \mem[114][2] ,
         \mem[114][1] , \mem[114][0] , \mem[113][7] , \mem[113][6] ,
         \mem[113][5] , \mem[113][4] , \mem[113][3] , \mem[113][2] ,
         \mem[113][1] , \mem[113][0] , \mem[112][7] , \mem[112][6] ,
         \mem[112][5] , \mem[112][4] , \mem[112][3] , \mem[112][2] ,
         \mem[112][1] , \mem[112][0] , \mem[111][7] , \mem[111][6] ,
         \mem[111][5] , \mem[111][4] , \mem[111][3] , \mem[111][2] ,
         \mem[111][1] , \mem[111][0] , \mem[110][7] , \mem[110][6] ,
         \mem[110][5] , \mem[110][4] , \mem[110][3] , \mem[110][2] ,
         \mem[110][1] , \mem[110][0] , \mem[109][7] , \mem[109][6] ,
         \mem[109][5] , \mem[109][4] , \mem[109][3] , \mem[109][2] ,
         \mem[109][1] , \mem[109][0] , \mem[108][7] , \mem[108][6] ,
         \mem[108][5] , \mem[108][4] , \mem[108][3] , \mem[108][2] ,
         \mem[108][1] , \mem[108][0] , \mem[107][7] , \mem[107][6] ,
         \mem[107][5] , \mem[107][4] , \mem[107][3] , \mem[107][2] ,
         \mem[107][1] , \mem[107][0] , \mem[106][7] , \mem[106][6] ,
         \mem[106][5] , \mem[106][4] , \mem[106][3] , \mem[106][2] ,
         \mem[106][1] , \mem[106][0] , \mem[105][7] , \mem[105][6] ,
         \mem[105][5] , \mem[105][4] , \mem[105][3] , \mem[105][2] ,
         \mem[105][1] , \mem[105][0] , \mem[104][7] , \mem[104][6] ,
         \mem[104][5] , \mem[104][4] , \mem[104][3] , \mem[104][2] ,
         \mem[104][1] , \mem[104][0] , \mem[103][7] , \mem[103][6] ,
         \mem[103][5] , \mem[103][4] , \mem[103][3] , \mem[103][2] ,
         \mem[103][1] , \mem[103][0] , \mem[102][7] , \mem[102][6] ,
         \mem[102][5] , \mem[102][4] , \mem[102][3] , \mem[102][2] ,
         \mem[102][1] , \mem[102][0] , \mem[101][7] , \mem[101][6] ,
         \mem[101][5] , \mem[101][4] , \mem[101][3] , \mem[101][2] ,
         \mem[101][1] , \mem[101][0] , \mem[100][7] , \mem[100][6] ,
         \mem[100][5] , \mem[100][4] , \mem[100][3] , \mem[100][2] ,
         \mem[100][1] , \mem[100][0] , \mem[99][7] , \mem[99][6] ,
         \mem[99][5] , \mem[99][4] , \mem[99][3] , \mem[99][2] , \mem[99][1] ,
         \mem[99][0] , \mem[98][7] , \mem[98][6] , \mem[98][5] , \mem[98][4] ,
         \mem[98][3] , \mem[98][2] , \mem[98][1] , \mem[98][0] , \mem[97][7] ,
         \mem[97][6] , \mem[97][5] , \mem[97][4] , \mem[97][3] , \mem[97][2] ,
         \mem[97][1] , \mem[97][0] , \mem[96][7] , \mem[96][6] , \mem[96][5] ,
         \mem[96][4] , \mem[96][3] , \mem[96][2] , \mem[96][1] , \mem[96][0] ,
         \mem[95][7] , \mem[95][6] , \mem[95][5] , \mem[95][4] , \mem[95][3] ,
         \mem[95][2] , \mem[95][1] , \mem[95][0] , \mem[94][7] , \mem[94][6] ,
         \mem[94][5] , \mem[94][4] , \mem[94][3] , \mem[94][2] , \mem[94][1] ,
         \mem[94][0] , \mem[93][7] , \mem[93][6] , \mem[93][5] , \mem[93][4] ,
         \mem[93][3] , \mem[93][2] , \mem[93][1] , \mem[93][0] , \mem[92][7] ,
         \mem[92][6] , \mem[92][5] , \mem[92][4] , \mem[92][3] , \mem[92][2] ,
         \mem[92][1] , \mem[92][0] , \mem[91][7] , \mem[91][6] , \mem[91][5] ,
         \mem[91][4] , \mem[91][3] , \mem[91][2] , \mem[91][1] , \mem[91][0] ,
         \mem[90][7] , \mem[90][6] , \mem[90][5] , \mem[90][4] , \mem[90][3] ,
         \mem[90][2] , \mem[90][1] , \mem[90][0] , \mem[89][7] , \mem[89][6] ,
         \mem[89][5] , \mem[89][4] , \mem[89][3] , \mem[89][2] , \mem[89][1] ,
         \mem[89][0] , \mem[88][7] , \mem[88][6] , \mem[88][5] , \mem[88][4] ,
         \mem[88][3] , \mem[88][2] , \mem[88][1] , \mem[88][0] , \mem[87][7] ,
         \mem[87][6] , \mem[87][5] , \mem[87][4] , \mem[87][3] , \mem[87][2] ,
         \mem[87][1] , \mem[87][0] , \mem[86][7] , \mem[86][6] , \mem[86][5] ,
         \mem[86][4] , \mem[86][3] , \mem[86][2] , \mem[86][1] , \mem[86][0] ,
         \mem[85][7] , \mem[85][6] , \mem[85][5] , \mem[85][4] , \mem[85][3] ,
         \mem[85][2] , \mem[85][1] , \mem[85][0] , \mem[84][7] , \mem[84][6] ,
         \mem[84][5] , \mem[84][4] , \mem[84][3] , \mem[84][2] , \mem[84][1] ,
         \mem[84][0] , \mem[83][7] , \mem[83][6] , \mem[83][5] , \mem[83][4] ,
         \mem[83][3] , \mem[83][2] , \mem[83][1] , \mem[83][0] , \mem[82][7] ,
         \mem[82][6] , \mem[82][5] , \mem[82][4] , \mem[82][3] , \mem[82][2] ,
         \mem[82][1] , \mem[82][0] , \mem[81][7] , \mem[81][6] , \mem[81][5] ,
         \mem[81][4] , \mem[81][3] , \mem[81][2] , \mem[81][1] , \mem[81][0] ,
         \mem[80][7] , \mem[80][6] , \mem[80][5] , \mem[80][4] , \mem[80][3] ,
         \mem[80][2] , \mem[80][1] , \mem[80][0] , \mem[79][7] , \mem[79][6] ,
         \mem[79][5] , \mem[79][4] , \mem[79][3] , \mem[79][2] , \mem[79][1] ,
         \mem[79][0] , \mem[78][7] , \mem[78][6] , \mem[78][5] , \mem[78][4] ,
         \mem[78][3] , \mem[78][2] , \mem[78][1] , \mem[78][0] , \mem[77][7] ,
         \mem[77][6] , \mem[77][5] , \mem[77][4] , \mem[77][3] , \mem[77][2] ,
         \mem[77][1] , \mem[77][0] , \mem[76][7] , \mem[76][6] , \mem[76][5] ,
         \mem[76][4] , \mem[76][3] , \mem[76][2] , \mem[76][1] , \mem[76][0] ,
         \mem[75][7] , \mem[75][6] , \mem[75][5] , \mem[75][4] , \mem[75][3] ,
         \mem[75][2] , \mem[75][1] , \mem[75][0] , \mem[74][7] , \mem[74][6] ,
         \mem[74][5] , \mem[74][4] , \mem[74][3] , \mem[74][2] , \mem[74][1] ,
         \mem[74][0] , \mem[73][7] , \mem[73][6] , \mem[73][5] , \mem[73][4] ,
         \mem[73][3] , \mem[73][2] , \mem[73][1] , \mem[73][0] , \mem[72][7] ,
         \mem[72][6] , \mem[72][5] , \mem[72][4] , \mem[72][3] , \mem[72][2] ,
         \mem[72][1] , \mem[72][0] , \mem[71][7] , \mem[71][6] , \mem[71][5] ,
         \mem[71][4] , \mem[71][3] , \mem[71][2] , \mem[71][1] , \mem[71][0] ,
         \mem[70][7] , \mem[70][6] , \mem[70][5] , \mem[70][4] , \mem[70][3] ,
         \mem[70][2] , \mem[70][1] , \mem[70][0] , \mem[69][7] , \mem[69][6] ,
         \mem[69][5] , \mem[69][4] , \mem[69][3] , \mem[69][2] , \mem[69][1] ,
         \mem[69][0] , \mem[68][7] , \mem[68][6] , \mem[68][5] , \mem[68][4] ,
         \mem[68][3] , \mem[68][2] , \mem[68][1] , \mem[68][0] , \mem[67][7] ,
         \mem[67][6] , \mem[67][5] , \mem[67][4] , \mem[67][3] , \mem[67][2] ,
         \mem[67][1] , \mem[67][0] , \mem[66][7] , \mem[66][6] , \mem[66][5] ,
         \mem[66][4] , \mem[66][3] , \mem[66][2] , \mem[66][1] , \mem[66][0] ,
         \mem[65][7] , \mem[65][6] , \mem[65][5] , \mem[65][4] , \mem[65][3] ,
         \mem[65][2] , \mem[65][1] , \mem[65][0] , \mem[64][7] , \mem[64][6] ,
         \mem[64][5] , \mem[64][4] , \mem[64][3] , \mem[64][2] , \mem[64][1] ,
         \mem[64][0] , \mem[63][7] , \mem[63][6] , \mem[63][5] , \mem[63][4] ,
         \mem[63][3] , \mem[63][2] , \mem[63][1] , \mem[63][0] , \mem[62][7] ,
         \mem[62][6] , \mem[62][5] , \mem[62][4] , \mem[62][3] , \mem[62][2] ,
         \mem[62][1] , \mem[62][0] , \mem[61][7] , \mem[61][6] , \mem[61][5] ,
         \mem[61][4] , \mem[61][3] , \mem[61][2] , \mem[61][1] , \mem[61][0] ,
         \mem[60][7] , \mem[60][6] , \mem[60][5] , \mem[60][4] , \mem[60][3] ,
         \mem[60][2] , \mem[60][1] , \mem[60][0] , \mem[59][7] , \mem[59][6] ,
         \mem[59][5] , \mem[59][4] , \mem[59][3] , \mem[59][2] , \mem[59][1] ,
         \mem[59][0] , \mem[58][7] , \mem[58][6] , \mem[58][5] , \mem[58][4] ,
         \mem[58][3] , \mem[58][2] , \mem[58][1] , \mem[58][0] , \mem[57][7] ,
         \mem[57][6] , \mem[57][5] , \mem[57][4] , \mem[57][3] , \mem[57][2] ,
         \mem[57][1] , \mem[57][0] , \mem[56][7] , \mem[56][6] , \mem[56][5] ,
         \mem[56][4] , \mem[56][3] , \mem[56][2] , \mem[56][1] , \mem[56][0] ,
         \mem[55][7] , \mem[55][6] , \mem[55][5] , \mem[55][4] , \mem[55][3] ,
         \mem[55][2] , \mem[55][1] , \mem[55][0] , \mem[54][7] , \mem[54][6] ,
         \mem[54][5] , \mem[54][4] , \mem[54][3] , \mem[54][2] , \mem[54][1] ,
         \mem[54][0] , \mem[53][7] , \mem[53][6] , \mem[53][5] , \mem[53][4] ,
         \mem[53][3] , \mem[53][2] , \mem[53][1] , \mem[53][0] , \mem[52][7] ,
         \mem[52][6] , \mem[52][5] , \mem[52][4] , \mem[52][3] , \mem[52][2] ,
         \mem[52][1] , \mem[52][0] , \mem[51][7] , \mem[51][6] , \mem[51][5] ,
         \mem[51][4] , \mem[51][3] , \mem[51][2] , \mem[51][1] , \mem[51][0] ,
         \mem[50][7] , \mem[50][6] , \mem[50][5] , \mem[50][4] , \mem[50][3] ,
         \mem[50][2] , \mem[50][1] , \mem[50][0] , \mem[49][7] , \mem[49][6] ,
         \mem[49][5] , \mem[49][4] , \mem[49][3] , \mem[49][2] , \mem[49][1] ,
         \mem[49][0] , \mem[48][7] , \mem[48][6] , \mem[48][5] , \mem[48][4] ,
         \mem[48][3] , \mem[48][2] , \mem[48][1] , \mem[48][0] , \mem[47][7] ,
         \mem[47][6] , \mem[47][5] , \mem[47][4] , \mem[47][3] , \mem[47][2] ,
         \mem[47][1] , \mem[47][0] , \mem[46][7] , \mem[46][6] , \mem[46][5] ,
         \mem[46][4] , \mem[46][3] , \mem[46][2] , \mem[46][1] , \mem[46][0] ,
         \mem[45][7] , \mem[45][6] , \mem[45][5] , \mem[45][4] , \mem[45][3] ,
         \mem[45][2] , \mem[45][1] , \mem[45][0] , \mem[44][7] , \mem[44][6] ,
         \mem[44][5] , \mem[44][4] , \mem[44][3] , \mem[44][2] , \mem[44][1] ,
         \mem[44][0] , \mem[43][7] , \mem[43][6] , \mem[43][5] , \mem[43][4] ,
         \mem[43][3] , \mem[43][2] , \mem[43][1] , \mem[43][0] , \mem[42][7] ,
         \mem[42][6] , \mem[42][5] , \mem[42][4] , \mem[42][3] , \mem[42][2] ,
         \mem[42][1] , \mem[42][0] , \mem[41][7] , \mem[41][6] , \mem[41][5] ,
         \mem[41][4] , \mem[41][3] , \mem[41][2] , \mem[41][1] , \mem[41][0] ,
         \mem[40][7] , \mem[40][6] , \mem[40][5] , \mem[40][4] , \mem[40][3] ,
         \mem[40][2] , \mem[40][1] , \mem[40][0] , \mem[39][7] , \mem[39][6] ,
         \mem[39][5] , \mem[39][4] , \mem[39][3] , \mem[39][2] , \mem[39][1] ,
         \mem[39][0] , \mem[38][7] , \mem[38][6] , \mem[38][5] , \mem[38][4] ,
         \mem[38][3] , \mem[38][2] , \mem[38][1] , \mem[38][0] , \mem[37][7] ,
         \mem[37][6] , \mem[37][5] , \mem[37][4] , \mem[37][3] , \mem[37][2] ,
         \mem[37][1] , \mem[37][0] , \mem[36][7] , \mem[36][6] , \mem[36][5] ,
         \mem[36][4] , \mem[36][3] , \mem[36][2] , \mem[36][1] , \mem[36][0] ,
         \mem[35][7] , \mem[35][6] , \mem[35][5] , \mem[35][4] , \mem[35][3] ,
         \mem[35][2] , \mem[35][1] , \mem[35][0] , \mem[34][7] , \mem[34][6] ,
         \mem[34][5] , \mem[34][4] , \mem[34][3] , \mem[34][2] , \mem[34][1] ,
         \mem[34][0] , \mem[33][7] , \mem[33][6] , \mem[33][5] , \mem[33][4] ,
         \mem[33][3] , \mem[33][2] , \mem[33][1] , \mem[33][0] , \mem[32][7] ,
         \mem[32][6] , \mem[32][5] , \mem[32][4] , \mem[32][3] , \mem[32][2] ,
         \mem[32][1] , \mem[32][0] , \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N33, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885;
  assign N18 = addr[0];
  assign N19 = addr[1];
  assign N20 = addr[2];
  assign N21 = addr[3];
  assign N22 = addr[4];
  assign N23 = addr[5];
  assign N24 = addr[6];
  assign N25 = addr[7];

  DFF_X1 \data_out_reg[0]  ( .D(N33), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[255][7]  ( .D(n2229), .CK(clk), .Q(\mem[255][7] ) );
  DFF_X1 \mem_reg[255][6]  ( .D(n2230), .CK(clk), .Q(\mem[255][6] ) );
  DFF_X1 \mem_reg[255][5]  ( .D(n2231), .CK(clk), .Q(\mem[255][5] ) );
  DFF_X1 \mem_reg[255][4]  ( .D(n2232), .CK(clk), .Q(\mem[255][4] ) );
  DFF_X1 \mem_reg[255][3]  ( .D(n2233), .CK(clk), .Q(\mem[255][3] ) );
  DFF_X1 \mem_reg[255][2]  ( .D(n2234), .CK(clk), .Q(\mem[255][2] ) );
  DFF_X1 \mem_reg[255][1]  ( .D(n2235), .CK(clk), .Q(\mem[255][1] ) );
  DFF_X1 \mem_reg[255][0]  ( .D(n2236), .CK(clk), .Q(\mem[255][0] ) );
  DFF_X1 \mem_reg[254][7]  ( .D(n2237), .CK(clk), .Q(\mem[254][7] ) );
  DFF_X1 \mem_reg[254][6]  ( .D(n2238), .CK(clk), .Q(\mem[254][6] ) );
  DFF_X1 \mem_reg[254][5]  ( .D(n2239), .CK(clk), .Q(\mem[254][5] ) );
  DFF_X1 \mem_reg[254][4]  ( .D(n2240), .CK(clk), .Q(\mem[254][4] ) );
  DFF_X1 \mem_reg[254][3]  ( .D(n2241), .CK(clk), .Q(\mem[254][3] ) );
  DFF_X1 \mem_reg[254][2]  ( .D(n2242), .CK(clk), .Q(\mem[254][2] ) );
  DFF_X1 \mem_reg[254][1]  ( .D(n2243), .CK(clk), .Q(\mem[254][1] ) );
  DFF_X1 \mem_reg[254][0]  ( .D(n2244), .CK(clk), .Q(\mem[254][0] ) );
  DFF_X1 \mem_reg[253][7]  ( .D(n2245), .CK(clk), .Q(\mem[253][7] ) );
  DFF_X1 \mem_reg[253][6]  ( .D(n2246), .CK(clk), .Q(\mem[253][6] ) );
  DFF_X1 \mem_reg[253][5]  ( .D(n2247), .CK(clk), .Q(\mem[253][5] ) );
  DFF_X1 \mem_reg[253][4]  ( .D(n2248), .CK(clk), .Q(\mem[253][4] ) );
  DFF_X1 \mem_reg[253][3]  ( .D(n2249), .CK(clk), .Q(\mem[253][3] ) );
  DFF_X1 \mem_reg[253][2]  ( .D(n2250), .CK(clk), .Q(\mem[253][2] ) );
  DFF_X1 \mem_reg[253][1]  ( .D(n2251), .CK(clk), .Q(\mem[253][1] ) );
  DFF_X1 \mem_reg[253][0]  ( .D(n2252), .CK(clk), .Q(\mem[253][0] ) );
  DFF_X1 \mem_reg[252][7]  ( .D(n2253), .CK(clk), .Q(\mem[252][7] ) );
  DFF_X1 \mem_reg[252][6]  ( .D(n2254), .CK(clk), .Q(\mem[252][6] ) );
  DFF_X1 \mem_reg[252][5]  ( .D(n2255), .CK(clk), .Q(\mem[252][5] ) );
  DFF_X1 \mem_reg[252][4]  ( .D(n2256), .CK(clk), .Q(\mem[252][4] ) );
  DFF_X1 \mem_reg[252][3]  ( .D(n2257), .CK(clk), .Q(\mem[252][3] ) );
  DFF_X1 \mem_reg[252][2]  ( .D(n2258), .CK(clk), .Q(\mem[252][2] ) );
  DFF_X1 \mem_reg[252][1]  ( .D(n2259), .CK(clk), .Q(\mem[252][1] ) );
  DFF_X1 \mem_reg[252][0]  ( .D(n2260), .CK(clk), .Q(\mem[252][0] ) );
  DFF_X1 \mem_reg[251][7]  ( .D(n2261), .CK(clk), .Q(\mem[251][7] ) );
  DFF_X1 \mem_reg[251][6]  ( .D(n2262), .CK(clk), .Q(\mem[251][6] ) );
  DFF_X1 \mem_reg[251][5]  ( .D(n2263), .CK(clk), .Q(\mem[251][5] ) );
  DFF_X1 \mem_reg[251][4]  ( .D(n2264), .CK(clk), .Q(\mem[251][4] ) );
  DFF_X1 \mem_reg[251][3]  ( .D(n2265), .CK(clk), .Q(\mem[251][3] ) );
  DFF_X1 \mem_reg[251][2]  ( .D(n2266), .CK(clk), .Q(\mem[251][2] ) );
  DFF_X1 \mem_reg[251][1]  ( .D(n2267), .CK(clk), .Q(\mem[251][1] ) );
  DFF_X1 \mem_reg[251][0]  ( .D(n2268), .CK(clk), .Q(\mem[251][0] ) );
  DFF_X1 \mem_reg[250][7]  ( .D(n2269), .CK(clk), .Q(\mem[250][7] ) );
  DFF_X1 \mem_reg[250][6]  ( .D(n2270), .CK(clk), .Q(\mem[250][6] ) );
  DFF_X1 \mem_reg[250][5]  ( .D(n2271), .CK(clk), .Q(\mem[250][5] ) );
  DFF_X1 \mem_reg[250][4]  ( .D(n2272), .CK(clk), .Q(\mem[250][4] ) );
  DFF_X1 \mem_reg[250][3]  ( .D(n2273), .CK(clk), .Q(\mem[250][3] ) );
  DFF_X1 \mem_reg[250][2]  ( .D(n2274), .CK(clk), .Q(\mem[250][2] ) );
  DFF_X1 \mem_reg[250][1]  ( .D(n2275), .CK(clk), .Q(\mem[250][1] ) );
  DFF_X1 \mem_reg[250][0]  ( .D(n2276), .CK(clk), .Q(\mem[250][0] ) );
  DFF_X1 \mem_reg[249][7]  ( .D(n2277), .CK(clk), .Q(\mem[249][7] ) );
  DFF_X1 \mem_reg[249][6]  ( .D(n2278), .CK(clk), .Q(\mem[249][6] ) );
  DFF_X1 \mem_reg[249][5]  ( .D(n2279), .CK(clk), .Q(\mem[249][5] ) );
  DFF_X1 \mem_reg[249][4]  ( .D(n2280), .CK(clk), .Q(\mem[249][4] ) );
  DFF_X1 \mem_reg[249][3]  ( .D(n2281), .CK(clk), .Q(\mem[249][3] ) );
  DFF_X1 \mem_reg[249][2]  ( .D(n2282), .CK(clk), .Q(\mem[249][2] ) );
  DFF_X1 \mem_reg[249][1]  ( .D(n2283), .CK(clk), .Q(\mem[249][1] ) );
  DFF_X1 \mem_reg[249][0]  ( .D(n2284), .CK(clk), .Q(\mem[249][0] ) );
  DFF_X1 \mem_reg[248][7]  ( .D(n2285), .CK(clk), .Q(\mem[248][7] ) );
  DFF_X1 \mem_reg[248][6]  ( .D(n2286), .CK(clk), .Q(\mem[248][6] ) );
  DFF_X1 \mem_reg[248][5]  ( .D(n2287), .CK(clk), .Q(\mem[248][5] ) );
  DFF_X1 \mem_reg[248][4]  ( .D(n2288), .CK(clk), .Q(\mem[248][4] ) );
  DFF_X1 \mem_reg[248][3]  ( .D(n2289), .CK(clk), .Q(\mem[248][3] ) );
  DFF_X1 \mem_reg[248][2]  ( .D(n2290), .CK(clk), .Q(\mem[248][2] ) );
  DFF_X1 \mem_reg[248][1]  ( .D(n2291), .CK(clk), .Q(\mem[248][1] ) );
  DFF_X1 \mem_reg[248][0]  ( .D(n2292), .CK(clk), .Q(\mem[248][0] ) );
  DFF_X1 \mem_reg[247][7]  ( .D(n2293), .CK(clk), .Q(\mem[247][7] ) );
  DFF_X1 \mem_reg[247][6]  ( .D(n2294), .CK(clk), .Q(\mem[247][6] ) );
  DFF_X1 \mem_reg[247][5]  ( .D(n2295), .CK(clk), .Q(\mem[247][5] ) );
  DFF_X1 \mem_reg[247][4]  ( .D(n2296), .CK(clk), .Q(\mem[247][4] ) );
  DFF_X1 \mem_reg[247][3]  ( .D(n2297), .CK(clk), .Q(\mem[247][3] ) );
  DFF_X1 \mem_reg[247][2]  ( .D(n2298), .CK(clk), .Q(\mem[247][2] ) );
  DFF_X1 \mem_reg[247][1]  ( .D(n2299), .CK(clk), .Q(\mem[247][1] ) );
  DFF_X1 \mem_reg[247][0]  ( .D(n2300), .CK(clk), .Q(\mem[247][0] ) );
  DFF_X1 \mem_reg[246][7]  ( .D(n2301), .CK(clk), .Q(\mem[246][7] ) );
  DFF_X1 \mem_reg[246][6]  ( .D(n2302), .CK(clk), .Q(\mem[246][6] ) );
  DFF_X1 \mem_reg[246][5]  ( .D(n2303), .CK(clk), .Q(\mem[246][5] ) );
  DFF_X1 \mem_reg[246][4]  ( .D(n2304), .CK(clk), .Q(\mem[246][4] ) );
  DFF_X1 \mem_reg[246][3]  ( .D(n2305), .CK(clk), .Q(\mem[246][3] ) );
  DFF_X1 \mem_reg[246][2]  ( .D(n2306), .CK(clk), .Q(\mem[246][2] ) );
  DFF_X1 \mem_reg[246][1]  ( .D(n2307), .CK(clk), .Q(\mem[246][1] ) );
  DFF_X1 \mem_reg[246][0]  ( .D(n2308), .CK(clk), .Q(\mem[246][0] ) );
  DFF_X1 \mem_reg[245][7]  ( .D(n2309), .CK(clk), .Q(\mem[245][7] ) );
  DFF_X1 \mem_reg[245][6]  ( .D(n2310), .CK(clk), .Q(\mem[245][6] ) );
  DFF_X1 \mem_reg[245][5]  ( .D(n2311), .CK(clk), .Q(\mem[245][5] ) );
  DFF_X1 \mem_reg[245][4]  ( .D(n2312), .CK(clk), .Q(\mem[245][4] ) );
  DFF_X1 \mem_reg[245][3]  ( .D(n4665), .CK(clk), .Q(\mem[245][3] ) );
  DFF_X1 \mem_reg[245][2]  ( .D(n4666), .CK(clk), .Q(\mem[245][2] ) );
  DFF_X1 \mem_reg[245][1]  ( .D(n4667), .CK(clk), .Q(\mem[245][1] ) );
  DFF_X1 \mem_reg[245][0]  ( .D(n4668), .CK(clk), .Q(\mem[245][0] ) );
  DFF_X1 \mem_reg[244][7]  ( .D(n4669), .CK(clk), .Q(\mem[244][7] ) );
  DFF_X1 \mem_reg[244][6]  ( .D(n4670), .CK(clk), .Q(\mem[244][6] ) );
  DFF_X1 \mem_reg[244][5]  ( .D(n4671), .CK(clk), .Q(\mem[244][5] ) );
  DFF_X1 \mem_reg[244][4]  ( .D(n4672), .CK(clk), .Q(\mem[244][4] ) );
  DFF_X1 \mem_reg[244][3]  ( .D(n4673), .CK(clk), .Q(\mem[244][3] ) );
  DFF_X1 \mem_reg[244][2]  ( .D(n4674), .CK(clk), .Q(\mem[244][2] ) );
  DFF_X1 \mem_reg[244][1]  ( .D(n4675), .CK(clk), .Q(\mem[244][1] ) );
  DFF_X1 \mem_reg[244][0]  ( .D(n4676), .CK(clk), .Q(\mem[244][0] ) );
  DFF_X1 \mem_reg[243][7]  ( .D(n4677), .CK(clk), .Q(\mem[243][7] ) );
  DFF_X1 \mem_reg[243][6]  ( .D(n4678), .CK(clk), .Q(\mem[243][6] ) );
  DFF_X1 \mem_reg[243][5]  ( .D(n4679), .CK(clk), .Q(\mem[243][5] ) );
  DFF_X1 \mem_reg[243][4]  ( .D(n4680), .CK(clk), .Q(\mem[243][4] ) );
  DFF_X1 \mem_reg[243][3]  ( .D(n4681), .CK(clk), .Q(\mem[243][3] ) );
  DFF_X1 \mem_reg[243][2]  ( .D(n4682), .CK(clk), .Q(\mem[243][2] ) );
  DFF_X1 \mem_reg[243][1]  ( .D(n4683), .CK(clk), .Q(\mem[243][1] ) );
  DFF_X1 \mem_reg[243][0]  ( .D(n4684), .CK(clk), .Q(\mem[243][0] ) );
  DFF_X1 \mem_reg[242][7]  ( .D(n4685), .CK(clk), .Q(\mem[242][7] ) );
  DFF_X1 \mem_reg[242][6]  ( .D(n4686), .CK(clk), .Q(\mem[242][6] ) );
  DFF_X1 \mem_reg[242][5]  ( .D(n4687), .CK(clk), .Q(\mem[242][5] ) );
  DFF_X1 \mem_reg[242][4]  ( .D(n4688), .CK(clk), .Q(\mem[242][4] ) );
  DFF_X1 \mem_reg[242][3]  ( .D(n4689), .CK(clk), .Q(\mem[242][3] ) );
  DFF_X1 \mem_reg[242][2]  ( .D(n4690), .CK(clk), .Q(\mem[242][2] ) );
  DFF_X1 \mem_reg[242][1]  ( .D(n4691), .CK(clk), .Q(\mem[242][1] ) );
  DFF_X1 \mem_reg[242][0]  ( .D(n4692), .CK(clk), .Q(\mem[242][0] ) );
  DFF_X1 \mem_reg[241][7]  ( .D(n4693), .CK(clk), .Q(\mem[241][7] ) );
  DFF_X1 \mem_reg[241][6]  ( .D(n4694), .CK(clk), .Q(\mem[241][6] ) );
  DFF_X1 \mem_reg[241][5]  ( .D(n4695), .CK(clk), .Q(\mem[241][5] ) );
  DFF_X1 \mem_reg[241][4]  ( .D(n4696), .CK(clk), .Q(\mem[241][4] ) );
  DFF_X1 \mem_reg[241][3]  ( .D(n4697), .CK(clk), .Q(\mem[241][3] ) );
  DFF_X1 \mem_reg[241][2]  ( .D(n4698), .CK(clk), .Q(\mem[241][2] ) );
  DFF_X1 \mem_reg[241][1]  ( .D(n4699), .CK(clk), .Q(\mem[241][1] ) );
  DFF_X1 \mem_reg[241][0]  ( .D(n4700), .CK(clk), .Q(\mem[241][0] ) );
  DFF_X1 \mem_reg[240][7]  ( .D(n4701), .CK(clk), .Q(\mem[240][7] ) );
  DFF_X1 \mem_reg[240][6]  ( .D(n4702), .CK(clk), .Q(\mem[240][6] ) );
  DFF_X1 \mem_reg[240][5]  ( .D(n4703), .CK(clk), .Q(\mem[240][5] ) );
  DFF_X1 \mem_reg[240][4]  ( .D(n4704), .CK(clk), .Q(\mem[240][4] ) );
  DFF_X1 \mem_reg[240][3]  ( .D(n4705), .CK(clk), .Q(\mem[240][3] ) );
  DFF_X1 \mem_reg[240][2]  ( .D(n4706), .CK(clk), .Q(\mem[240][2] ) );
  DFF_X1 \mem_reg[240][1]  ( .D(n4707), .CK(clk), .Q(\mem[240][1] ) );
  DFF_X1 \mem_reg[240][0]  ( .D(n4708), .CK(clk), .Q(\mem[240][0] ) );
  DFF_X1 \mem_reg[239][7]  ( .D(n4709), .CK(clk), .Q(\mem[239][7] ) );
  DFF_X1 \mem_reg[239][6]  ( .D(n4710), .CK(clk), .Q(\mem[239][6] ) );
  DFF_X1 \mem_reg[239][5]  ( .D(n4711), .CK(clk), .Q(\mem[239][5] ) );
  DFF_X1 \mem_reg[239][4]  ( .D(n4712), .CK(clk), .Q(\mem[239][4] ) );
  DFF_X1 \mem_reg[239][3]  ( .D(n4713), .CK(clk), .Q(\mem[239][3] ) );
  DFF_X1 \mem_reg[239][2]  ( .D(n4714), .CK(clk), .Q(\mem[239][2] ) );
  DFF_X1 \mem_reg[239][1]  ( .D(n4715), .CK(clk), .Q(\mem[239][1] ) );
  DFF_X1 \mem_reg[239][0]  ( .D(n4716), .CK(clk), .Q(\mem[239][0] ) );
  DFF_X1 \mem_reg[238][7]  ( .D(n4717), .CK(clk), .Q(\mem[238][7] ) );
  DFF_X1 \mem_reg[238][6]  ( .D(n4718), .CK(clk), .Q(\mem[238][6] ) );
  DFF_X1 \mem_reg[238][5]  ( .D(n4719), .CK(clk), .Q(\mem[238][5] ) );
  DFF_X1 \mem_reg[238][4]  ( .D(n4720), .CK(clk), .Q(\mem[238][4] ) );
  DFF_X1 \mem_reg[238][3]  ( .D(n4721), .CK(clk), .Q(\mem[238][3] ) );
  DFF_X1 \mem_reg[238][2]  ( .D(n4722), .CK(clk), .Q(\mem[238][2] ) );
  DFF_X1 \mem_reg[238][1]  ( .D(n4723), .CK(clk), .Q(\mem[238][1] ) );
  DFF_X1 \mem_reg[238][0]  ( .D(n4724), .CK(clk), .Q(\mem[238][0] ) );
  DFF_X1 \mem_reg[237][7]  ( .D(n4725), .CK(clk), .Q(\mem[237][7] ) );
  DFF_X1 \mem_reg[237][6]  ( .D(n4726), .CK(clk), .Q(\mem[237][6] ) );
  DFF_X1 \mem_reg[237][5]  ( .D(n4727), .CK(clk), .Q(\mem[237][5] ) );
  DFF_X1 \mem_reg[237][4]  ( .D(n4728), .CK(clk), .Q(\mem[237][4] ) );
  DFF_X1 \mem_reg[237][3]  ( .D(n4729), .CK(clk), .Q(\mem[237][3] ) );
  DFF_X1 \mem_reg[237][2]  ( .D(n4730), .CK(clk), .Q(\mem[237][2] ) );
  DFF_X1 \mem_reg[237][1]  ( .D(n4731), .CK(clk), .Q(\mem[237][1] ) );
  DFF_X1 \mem_reg[237][0]  ( .D(n4732), .CK(clk), .Q(\mem[237][0] ) );
  DFF_X1 \mem_reg[236][7]  ( .D(n4733), .CK(clk), .Q(\mem[236][7] ) );
  DFF_X1 \mem_reg[236][6]  ( .D(n4734), .CK(clk), .Q(\mem[236][6] ) );
  DFF_X1 \mem_reg[236][5]  ( .D(n4735), .CK(clk), .Q(\mem[236][5] ) );
  DFF_X1 \mem_reg[236][4]  ( .D(n4736), .CK(clk), .Q(\mem[236][4] ) );
  DFF_X1 \mem_reg[236][3]  ( .D(n4737), .CK(clk), .Q(\mem[236][3] ) );
  DFF_X1 \mem_reg[236][2]  ( .D(n4738), .CK(clk), .Q(\mem[236][2] ) );
  DFF_X1 \mem_reg[236][1]  ( .D(n4739), .CK(clk), .Q(\mem[236][1] ) );
  DFF_X1 \mem_reg[236][0]  ( .D(n4740), .CK(clk), .Q(\mem[236][0] ) );
  DFF_X1 \mem_reg[235][7]  ( .D(n4741), .CK(clk), .Q(\mem[235][7] ) );
  DFF_X1 \mem_reg[235][6]  ( .D(n4742), .CK(clk), .Q(\mem[235][6] ) );
  DFF_X1 \mem_reg[235][5]  ( .D(n4743), .CK(clk), .Q(\mem[235][5] ) );
  DFF_X1 \mem_reg[235][4]  ( .D(n4744), .CK(clk), .Q(\mem[235][4] ) );
  DFF_X1 \mem_reg[235][3]  ( .D(n4745), .CK(clk), .Q(\mem[235][3] ) );
  DFF_X1 \mem_reg[235][2]  ( .D(n4746), .CK(clk), .Q(\mem[235][2] ) );
  DFF_X1 \mem_reg[235][1]  ( .D(n4747), .CK(clk), .Q(\mem[235][1] ) );
  DFF_X1 \mem_reg[235][0]  ( .D(n4748), .CK(clk), .Q(\mem[235][0] ) );
  DFF_X1 \mem_reg[234][7]  ( .D(n4749), .CK(clk), .Q(\mem[234][7] ) );
  DFF_X1 \mem_reg[234][6]  ( .D(n4750), .CK(clk), .Q(\mem[234][6] ) );
  DFF_X1 \mem_reg[234][5]  ( .D(n4751), .CK(clk), .Q(\mem[234][5] ) );
  DFF_X1 \mem_reg[234][4]  ( .D(n4752), .CK(clk), .Q(\mem[234][4] ) );
  DFF_X1 \mem_reg[234][3]  ( .D(n4753), .CK(clk), .Q(\mem[234][3] ) );
  DFF_X1 \mem_reg[234][2]  ( .D(n4754), .CK(clk), .Q(\mem[234][2] ) );
  DFF_X1 \mem_reg[234][1]  ( .D(n4755), .CK(clk), .Q(\mem[234][1] ) );
  DFF_X1 \mem_reg[234][0]  ( .D(n4756), .CK(clk), .Q(\mem[234][0] ) );
  DFF_X1 \mem_reg[233][7]  ( .D(n4757), .CK(clk), .Q(\mem[233][7] ) );
  DFF_X1 \mem_reg[233][6]  ( .D(n4758), .CK(clk), .Q(\mem[233][6] ) );
  DFF_X1 \mem_reg[233][5]  ( .D(n4759), .CK(clk), .Q(\mem[233][5] ) );
  DFF_X1 \mem_reg[233][4]  ( .D(n4760), .CK(clk), .Q(\mem[233][4] ) );
  DFF_X1 \mem_reg[233][3]  ( .D(n4761), .CK(clk), .Q(\mem[233][3] ) );
  DFF_X1 \mem_reg[233][2]  ( .D(n4762), .CK(clk), .Q(\mem[233][2] ) );
  DFF_X1 \mem_reg[233][1]  ( .D(n4763), .CK(clk), .Q(\mem[233][1] ) );
  DFF_X1 \mem_reg[233][0]  ( .D(n4764), .CK(clk), .Q(\mem[233][0] ) );
  DFF_X1 \mem_reg[232][7]  ( .D(n4765), .CK(clk), .Q(\mem[232][7] ) );
  DFF_X1 \mem_reg[232][6]  ( .D(n4766), .CK(clk), .Q(\mem[232][6] ) );
  DFF_X1 \mem_reg[232][5]  ( .D(n4767), .CK(clk), .Q(\mem[232][5] ) );
  DFF_X1 \mem_reg[232][4]  ( .D(n4768), .CK(clk), .Q(\mem[232][4] ) );
  DFF_X1 \mem_reg[232][3]  ( .D(n4769), .CK(clk), .Q(\mem[232][3] ) );
  DFF_X1 \mem_reg[232][2]  ( .D(n4770), .CK(clk), .Q(\mem[232][2] ) );
  DFF_X1 \mem_reg[232][1]  ( .D(n4771), .CK(clk), .Q(\mem[232][1] ) );
  DFF_X1 \mem_reg[232][0]  ( .D(n4772), .CK(clk), .Q(\mem[232][0] ) );
  DFF_X1 \mem_reg[231][7]  ( .D(n4773), .CK(clk), .Q(\mem[231][7] ) );
  DFF_X1 \mem_reg[231][6]  ( .D(n4774), .CK(clk), .Q(\mem[231][6] ) );
  DFF_X1 \mem_reg[231][5]  ( .D(n4775), .CK(clk), .Q(\mem[231][5] ) );
  DFF_X1 \mem_reg[231][4]  ( .D(n4776), .CK(clk), .Q(\mem[231][4] ) );
  DFF_X1 \mem_reg[231][3]  ( .D(n4777), .CK(clk), .Q(\mem[231][3] ) );
  DFF_X1 \mem_reg[231][2]  ( .D(n4778), .CK(clk), .Q(\mem[231][2] ) );
  DFF_X1 \mem_reg[231][1]  ( .D(n4779), .CK(clk), .Q(\mem[231][1] ) );
  DFF_X1 \mem_reg[231][0]  ( .D(n4780), .CK(clk), .Q(\mem[231][0] ) );
  DFF_X1 \mem_reg[230][7]  ( .D(n4781), .CK(clk), .Q(\mem[230][7] ) );
  DFF_X1 \mem_reg[230][6]  ( .D(n4782), .CK(clk), .Q(\mem[230][6] ) );
  DFF_X1 \mem_reg[230][5]  ( .D(n4783), .CK(clk), .Q(\mem[230][5] ) );
  DFF_X1 \mem_reg[230][4]  ( .D(n4784), .CK(clk), .Q(\mem[230][4] ) );
  DFF_X1 \mem_reg[230][3]  ( .D(n4785), .CK(clk), .Q(\mem[230][3] ) );
  DFF_X1 \mem_reg[230][2]  ( .D(n4786), .CK(clk), .Q(\mem[230][2] ) );
  DFF_X1 \mem_reg[230][1]  ( .D(n4787), .CK(clk), .Q(\mem[230][1] ) );
  DFF_X1 \mem_reg[230][0]  ( .D(n4788), .CK(clk), .Q(\mem[230][0] ) );
  DFF_X1 \mem_reg[229][7]  ( .D(n4789), .CK(clk), .Q(\mem[229][7] ) );
  DFF_X1 \mem_reg[229][6]  ( .D(n4790), .CK(clk), .Q(\mem[229][6] ) );
  DFF_X1 \mem_reg[229][5]  ( .D(n4791), .CK(clk), .Q(\mem[229][5] ) );
  DFF_X1 \mem_reg[229][4]  ( .D(n4792), .CK(clk), .Q(\mem[229][4] ) );
  DFF_X1 \mem_reg[229][3]  ( .D(n4793), .CK(clk), .Q(\mem[229][3] ) );
  DFF_X1 \mem_reg[229][2]  ( .D(n4794), .CK(clk), .Q(\mem[229][2] ) );
  DFF_X1 \mem_reg[229][1]  ( .D(n4795), .CK(clk), .Q(\mem[229][1] ) );
  DFF_X1 \mem_reg[229][0]  ( .D(n4796), .CK(clk), .Q(\mem[229][0] ) );
  DFF_X1 \mem_reg[228][7]  ( .D(n4797), .CK(clk), .Q(\mem[228][7] ) );
  DFF_X1 \mem_reg[228][6]  ( .D(n4798), .CK(clk), .Q(\mem[228][6] ) );
  DFF_X1 \mem_reg[228][5]  ( .D(n4799), .CK(clk), .Q(\mem[228][5] ) );
  DFF_X1 \mem_reg[228][4]  ( .D(n4800), .CK(clk), .Q(\mem[228][4] ) );
  DFF_X1 \mem_reg[228][3]  ( .D(n4801), .CK(clk), .Q(\mem[228][3] ) );
  DFF_X1 \mem_reg[228][2]  ( .D(n4802), .CK(clk), .Q(\mem[228][2] ) );
  DFF_X1 \mem_reg[228][1]  ( .D(n4803), .CK(clk), .Q(\mem[228][1] ) );
  DFF_X1 \mem_reg[228][0]  ( .D(n4804), .CK(clk), .Q(\mem[228][0] ) );
  DFF_X1 \mem_reg[227][7]  ( .D(n4805), .CK(clk), .Q(\mem[227][7] ) );
  DFF_X1 \mem_reg[227][6]  ( .D(n4806), .CK(clk), .Q(\mem[227][6] ) );
  DFF_X1 \mem_reg[227][5]  ( .D(n4807), .CK(clk), .Q(\mem[227][5] ) );
  DFF_X1 \mem_reg[227][4]  ( .D(n4808), .CK(clk), .Q(\mem[227][4] ) );
  DFF_X1 \mem_reg[227][3]  ( .D(n4809), .CK(clk), .Q(\mem[227][3] ) );
  DFF_X1 \mem_reg[227][2]  ( .D(n4810), .CK(clk), .Q(\mem[227][2] ) );
  DFF_X1 \mem_reg[227][1]  ( .D(n4811), .CK(clk), .Q(\mem[227][1] ) );
  DFF_X1 \mem_reg[227][0]  ( .D(n4812), .CK(clk), .Q(\mem[227][0] ) );
  DFF_X1 \mem_reg[226][7]  ( .D(n4813), .CK(clk), .Q(\mem[226][7] ) );
  DFF_X1 \mem_reg[226][6]  ( .D(n4814), .CK(clk), .Q(\mem[226][6] ) );
  DFF_X1 \mem_reg[226][5]  ( .D(n4815), .CK(clk), .Q(\mem[226][5] ) );
  DFF_X1 \mem_reg[226][4]  ( .D(n4816), .CK(clk), .Q(\mem[226][4] ) );
  DFF_X1 \mem_reg[226][3]  ( .D(n4817), .CK(clk), .Q(\mem[226][3] ) );
  DFF_X1 \mem_reg[226][2]  ( .D(n4818), .CK(clk), .Q(\mem[226][2] ) );
  DFF_X1 \mem_reg[226][1]  ( .D(n4819), .CK(clk), .Q(\mem[226][1] ) );
  DFF_X1 \mem_reg[226][0]  ( .D(n4820), .CK(clk), .Q(\mem[226][0] ) );
  DFF_X1 \mem_reg[225][7]  ( .D(n4821), .CK(clk), .Q(\mem[225][7] ) );
  DFF_X1 \mem_reg[225][6]  ( .D(n4822), .CK(clk), .Q(\mem[225][6] ) );
  DFF_X1 \mem_reg[225][5]  ( .D(n4823), .CK(clk), .Q(\mem[225][5] ) );
  DFF_X1 \mem_reg[225][4]  ( .D(n4824), .CK(clk), .Q(\mem[225][4] ) );
  DFF_X1 \mem_reg[225][3]  ( .D(n4825), .CK(clk), .Q(\mem[225][3] ) );
  DFF_X1 \mem_reg[225][2]  ( .D(n4826), .CK(clk), .Q(\mem[225][2] ) );
  DFF_X1 \mem_reg[225][1]  ( .D(n4827), .CK(clk), .Q(\mem[225][1] ) );
  DFF_X1 \mem_reg[225][0]  ( .D(n4828), .CK(clk), .Q(\mem[225][0] ) );
  DFF_X1 \mem_reg[224][7]  ( .D(n4829), .CK(clk), .Q(\mem[224][7] ) );
  DFF_X1 \mem_reg[224][6]  ( .D(n4830), .CK(clk), .Q(\mem[224][6] ) );
  DFF_X1 \mem_reg[224][5]  ( .D(n4831), .CK(clk), .Q(\mem[224][5] ) );
  DFF_X1 \mem_reg[224][4]  ( .D(n4832), .CK(clk), .Q(\mem[224][4] ) );
  DFF_X1 \mem_reg[224][3]  ( .D(n4833), .CK(clk), .Q(\mem[224][3] ) );
  DFF_X1 \mem_reg[224][2]  ( .D(n4834), .CK(clk), .Q(\mem[224][2] ) );
  DFF_X1 \mem_reg[224][1]  ( .D(n4835), .CK(clk), .Q(\mem[224][1] ) );
  DFF_X1 \mem_reg[224][0]  ( .D(n4836), .CK(clk), .Q(\mem[224][0] ) );
  DFF_X1 \mem_reg[223][7]  ( .D(n4837), .CK(clk), .Q(\mem[223][7] ) );
  DFF_X1 \mem_reg[223][6]  ( .D(n4838), .CK(clk), .Q(\mem[223][6] ) );
  DFF_X1 \mem_reg[223][5]  ( .D(n4839), .CK(clk), .Q(\mem[223][5] ) );
  DFF_X1 \mem_reg[223][4]  ( .D(n4840), .CK(clk), .Q(\mem[223][4] ) );
  DFF_X1 \mem_reg[223][3]  ( .D(n4841), .CK(clk), .Q(\mem[223][3] ) );
  DFF_X1 \mem_reg[223][2]  ( .D(n4842), .CK(clk), .Q(\mem[223][2] ) );
  DFF_X1 \mem_reg[223][1]  ( .D(n4843), .CK(clk), .Q(\mem[223][1] ) );
  DFF_X1 \mem_reg[223][0]  ( .D(n4844), .CK(clk), .Q(\mem[223][0] ) );
  DFF_X1 \mem_reg[222][7]  ( .D(n4845), .CK(clk), .Q(\mem[222][7] ) );
  DFF_X1 \mem_reg[222][6]  ( .D(n4846), .CK(clk), .Q(\mem[222][6] ) );
  DFF_X1 \mem_reg[222][5]  ( .D(n4847), .CK(clk), .Q(\mem[222][5] ) );
  DFF_X1 \mem_reg[222][4]  ( .D(n4848), .CK(clk), .Q(\mem[222][4] ) );
  DFF_X1 \mem_reg[222][3]  ( .D(n4849), .CK(clk), .Q(\mem[222][3] ) );
  DFF_X1 \mem_reg[222][2]  ( .D(n4850), .CK(clk), .Q(\mem[222][2] ) );
  DFF_X1 \mem_reg[222][1]  ( .D(n4851), .CK(clk), .Q(\mem[222][1] ) );
  DFF_X1 \mem_reg[222][0]  ( .D(n4852), .CK(clk), .Q(\mem[222][0] ) );
  DFF_X1 \mem_reg[221][7]  ( .D(n4853), .CK(clk), .Q(\mem[221][7] ) );
  DFF_X1 \mem_reg[221][6]  ( .D(n4854), .CK(clk), .Q(\mem[221][6] ) );
  DFF_X1 \mem_reg[221][5]  ( .D(n4855), .CK(clk), .Q(\mem[221][5] ) );
  DFF_X1 \mem_reg[221][4]  ( .D(n4856), .CK(clk), .Q(\mem[221][4] ) );
  DFF_X1 \mem_reg[221][3]  ( .D(n4857), .CK(clk), .Q(\mem[221][3] ) );
  DFF_X1 \mem_reg[221][2]  ( .D(n4858), .CK(clk), .Q(\mem[221][2] ) );
  DFF_X1 \mem_reg[221][1]  ( .D(n4859), .CK(clk), .Q(\mem[221][1] ) );
  DFF_X1 \mem_reg[221][0]  ( .D(n4860), .CK(clk), .Q(\mem[221][0] ) );
  DFF_X1 \mem_reg[220][7]  ( .D(n4861), .CK(clk), .Q(\mem[220][7] ) );
  DFF_X1 \mem_reg[220][6]  ( .D(n4862), .CK(clk), .Q(\mem[220][6] ) );
  DFF_X1 \mem_reg[220][5]  ( .D(n4863), .CK(clk), .Q(\mem[220][5] ) );
  DFF_X1 \mem_reg[220][4]  ( .D(n4864), .CK(clk), .Q(\mem[220][4] ) );
  DFF_X1 \mem_reg[220][3]  ( .D(n4865), .CK(clk), .Q(\mem[220][3] ) );
  DFF_X1 \mem_reg[220][2]  ( .D(n4866), .CK(clk), .Q(\mem[220][2] ) );
  DFF_X1 \mem_reg[220][1]  ( .D(n4867), .CK(clk), .Q(\mem[220][1] ) );
  DFF_X1 \mem_reg[220][0]  ( .D(n4868), .CK(clk), .Q(\mem[220][0] ) );
  DFF_X1 \mem_reg[219][7]  ( .D(n4869), .CK(clk), .Q(\mem[219][7] ) );
  DFF_X1 \mem_reg[219][6]  ( .D(n4870), .CK(clk), .Q(\mem[219][6] ) );
  DFF_X1 \mem_reg[219][5]  ( .D(n4871), .CK(clk), .Q(\mem[219][5] ) );
  DFF_X1 \mem_reg[219][4]  ( .D(n4872), .CK(clk), .Q(\mem[219][4] ) );
  DFF_X1 \mem_reg[219][3]  ( .D(n4873), .CK(clk), .Q(\mem[219][3] ) );
  DFF_X1 \mem_reg[219][2]  ( .D(n4874), .CK(clk), .Q(\mem[219][2] ) );
  DFF_X1 \mem_reg[219][1]  ( .D(n4875), .CK(clk), .Q(\mem[219][1] ) );
  DFF_X1 \mem_reg[219][0]  ( .D(n4876), .CK(clk), .Q(\mem[219][0] ) );
  DFF_X1 \mem_reg[218][7]  ( .D(n4877), .CK(clk), .Q(\mem[218][7] ) );
  DFF_X1 \mem_reg[218][6]  ( .D(n4878), .CK(clk), .Q(\mem[218][6] ) );
  DFF_X1 \mem_reg[218][5]  ( .D(n4879), .CK(clk), .Q(\mem[218][5] ) );
  DFF_X1 \mem_reg[218][4]  ( .D(n4880), .CK(clk), .Q(\mem[218][4] ) );
  DFF_X1 \mem_reg[218][3]  ( .D(n4881), .CK(clk), .Q(\mem[218][3] ) );
  DFF_X1 \mem_reg[218][2]  ( .D(n4882), .CK(clk), .Q(\mem[218][2] ) );
  DFF_X1 \mem_reg[218][1]  ( .D(n4883), .CK(clk), .Q(\mem[218][1] ) );
  DFF_X1 \mem_reg[218][0]  ( .D(n4884), .CK(clk), .Q(\mem[218][0] ) );
  DFF_X1 \mem_reg[217][7]  ( .D(n4885), .CK(clk), .Q(\mem[217][7] ) );
  DFF_X1 \mem_reg[217][6]  ( .D(n4886), .CK(clk), .Q(\mem[217][6] ) );
  DFF_X1 \mem_reg[217][5]  ( .D(n4887), .CK(clk), .Q(\mem[217][5] ) );
  DFF_X1 \mem_reg[217][4]  ( .D(n4888), .CK(clk), .Q(\mem[217][4] ) );
  DFF_X1 \mem_reg[217][3]  ( .D(n4889), .CK(clk), .Q(\mem[217][3] ) );
  DFF_X1 \mem_reg[217][2]  ( .D(n4890), .CK(clk), .Q(\mem[217][2] ) );
  DFF_X1 \mem_reg[217][1]  ( .D(n4891), .CK(clk), .Q(\mem[217][1] ) );
  DFF_X1 \mem_reg[217][0]  ( .D(n4892), .CK(clk), .Q(\mem[217][0] ) );
  DFF_X1 \mem_reg[216][7]  ( .D(n4893), .CK(clk), .Q(\mem[216][7] ) );
  DFF_X1 \mem_reg[216][6]  ( .D(n4894), .CK(clk), .Q(\mem[216][6] ) );
  DFF_X1 \mem_reg[216][5]  ( .D(n4895), .CK(clk), .Q(\mem[216][5] ) );
  DFF_X1 \mem_reg[216][4]  ( .D(n4896), .CK(clk), .Q(\mem[216][4] ) );
  DFF_X1 \mem_reg[216][3]  ( .D(n4897), .CK(clk), .Q(\mem[216][3] ) );
  DFF_X1 \mem_reg[216][2]  ( .D(n4898), .CK(clk), .Q(\mem[216][2] ) );
  DFF_X1 \mem_reg[216][1]  ( .D(n4899), .CK(clk), .Q(\mem[216][1] ) );
  DFF_X1 \mem_reg[216][0]  ( .D(n4900), .CK(clk), .Q(\mem[216][0] ) );
  DFF_X1 \mem_reg[215][7]  ( .D(n4901), .CK(clk), .Q(\mem[215][7] ) );
  DFF_X1 \mem_reg[215][6]  ( .D(n4902), .CK(clk), .Q(\mem[215][6] ) );
  DFF_X1 \mem_reg[215][5]  ( .D(n4903), .CK(clk), .Q(\mem[215][5] ) );
  DFF_X1 \mem_reg[215][4]  ( .D(n4904), .CK(clk), .Q(\mem[215][4] ) );
  DFF_X1 \mem_reg[215][3]  ( .D(n4905), .CK(clk), .Q(\mem[215][3] ) );
  DFF_X1 \mem_reg[215][2]  ( .D(n4906), .CK(clk), .Q(\mem[215][2] ) );
  DFF_X1 \mem_reg[215][1]  ( .D(n4907), .CK(clk), .Q(\mem[215][1] ) );
  DFF_X1 \mem_reg[215][0]  ( .D(n4908), .CK(clk), .Q(\mem[215][0] ) );
  DFF_X1 \mem_reg[214][7]  ( .D(n4909), .CK(clk), .Q(\mem[214][7] ) );
  DFF_X1 \mem_reg[214][6]  ( .D(n4910), .CK(clk), .Q(\mem[214][6] ) );
  DFF_X1 \mem_reg[214][5]  ( .D(n4911), .CK(clk), .Q(\mem[214][5] ) );
  DFF_X1 \mem_reg[214][4]  ( .D(n4912), .CK(clk), .Q(\mem[214][4] ) );
  DFF_X1 \mem_reg[214][3]  ( .D(n4913), .CK(clk), .Q(\mem[214][3] ) );
  DFF_X1 \mem_reg[214][2]  ( .D(n4914), .CK(clk), .Q(\mem[214][2] ) );
  DFF_X1 \mem_reg[214][1]  ( .D(n4915), .CK(clk), .Q(\mem[214][1] ) );
  DFF_X1 \mem_reg[214][0]  ( .D(n4916), .CK(clk), .Q(\mem[214][0] ) );
  DFF_X1 \mem_reg[213][7]  ( .D(n4917), .CK(clk), .Q(\mem[213][7] ) );
  DFF_X1 \mem_reg[213][6]  ( .D(n4918), .CK(clk), .Q(\mem[213][6] ) );
  DFF_X1 \mem_reg[213][5]  ( .D(n4919), .CK(clk), .Q(\mem[213][5] ) );
  DFF_X1 \mem_reg[213][4]  ( .D(n4920), .CK(clk), .Q(\mem[213][4] ) );
  DFF_X1 \mem_reg[213][3]  ( .D(n4921), .CK(clk), .Q(\mem[213][3] ) );
  DFF_X1 \mem_reg[213][2]  ( .D(n4922), .CK(clk), .Q(\mem[213][2] ) );
  DFF_X1 \mem_reg[213][1]  ( .D(n4923), .CK(clk), .Q(\mem[213][1] ) );
  DFF_X1 \mem_reg[213][0]  ( .D(n4924), .CK(clk), .Q(\mem[213][0] ) );
  DFF_X1 \mem_reg[212][7]  ( .D(n4925), .CK(clk), .Q(\mem[212][7] ) );
  DFF_X1 \mem_reg[212][6]  ( .D(n4926), .CK(clk), .Q(\mem[212][6] ) );
  DFF_X1 \mem_reg[212][5]  ( .D(n4927), .CK(clk), .Q(\mem[212][5] ) );
  DFF_X1 \mem_reg[212][4]  ( .D(n4928), .CK(clk), .Q(\mem[212][4] ) );
  DFF_X1 \mem_reg[212][3]  ( .D(n4929), .CK(clk), .Q(\mem[212][3] ) );
  DFF_X1 \mem_reg[212][2]  ( .D(n4930), .CK(clk), .Q(\mem[212][2] ) );
  DFF_X1 \mem_reg[212][1]  ( .D(n4931), .CK(clk), .Q(\mem[212][1] ) );
  DFF_X1 \mem_reg[212][0]  ( .D(n4932), .CK(clk), .Q(\mem[212][0] ) );
  DFF_X1 \mem_reg[211][7]  ( .D(n4933), .CK(clk), .Q(\mem[211][7] ) );
  DFF_X1 \mem_reg[211][6]  ( .D(n4934), .CK(clk), .Q(\mem[211][6] ) );
  DFF_X1 \mem_reg[211][5]  ( .D(n4935), .CK(clk), .Q(\mem[211][5] ) );
  DFF_X1 \mem_reg[211][4]  ( .D(n4936), .CK(clk), .Q(\mem[211][4] ) );
  DFF_X1 \mem_reg[211][3]  ( .D(n4937), .CK(clk), .Q(\mem[211][3] ) );
  DFF_X1 \mem_reg[211][2]  ( .D(n4938), .CK(clk), .Q(\mem[211][2] ) );
  DFF_X1 \mem_reg[211][1]  ( .D(n4939), .CK(clk), .Q(\mem[211][1] ) );
  DFF_X1 \mem_reg[211][0]  ( .D(n4940), .CK(clk), .Q(\mem[211][0] ) );
  DFF_X1 \mem_reg[210][7]  ( .D(n4941), .CK(clk), .Q(\mem[210][7] ) );
  DFF_X1 \mem_reg[210][6]  ( .D(n4942), .CK(clk), .Q(\mem[210][6] ) );
  DFF_X1 \mem_reg[210][5]  ( .D(n4943), .CK(clk), .Q(\mem[210][5] ) );
  DFF_X1 \mem_reg[210][4]  ( .D(n4944), .CK(clk), .Q(\mem[210][4] ) );
  DFF_X1 \mem_reg[210][3]  ( .D(n4945), .CK(clk), .Q(\mem[210][3] ) );
  DFF_X1 \mem_reg[210][2]  ( .D(n4946), .CK(clk), .Q(\mem[210][2] ) );
  DFF_X1 \mem_reg[210][1]  ( .D(n4947), .CK(clk), .Q(\mem[210][1] ) );
  DFF_X1 \mem_reg[210][0]  ( .D(n4948), .CK(clk), .Q(\mem[210][0] ) );
  DFF_X1 \mem_reg[209][7]  ( .D(n4949), .CK(clk), .Q(\mem[209][7] ) );
  DFF_X1 \mem_reg[209][6]  ( .D(n4950), .CK(clk), .Q(\mem[209][6] ) );
  DFF_X1 \mem_reg[209][5]  ( .D(n4951), .CK(clk), .Q(\mem[209][5] ) );
  DFF_X1 \mem_reg[209][4]  ( .D(n4952), .CK(clk), .Q(\mem[209][4] ) );
  DFF_X1 \mem_reg[209][3]  ( .D(n4953), .CK(clk), .Q(\mem[209][3] ) );
  DFF_X1 \mem_reg[209][2]  ( .D(n4954), .CK(clk), .Q(\mem[209][2] ) );
  DFF_X1 \mem_reg[209][1]  ( .D(n4955), .CK(clk), .Q(\mem[209][1] ) );
  DFF_X1 \mem_reg[209][0]  ( .D(n4956), .CK(clk), .Q(\mem[209][0] ) );
  DFF_X1 \mem_reg[208][7]  ( .D(n4957), .CK(clk), .Q(\mem[208][7] ) );
  DFF_X1 \mem_reg[208][6]  ( .D(n4958), .CK(clk), .Q(\mem[208][6] ) );
  DFF_X1 \mem_reg[208][5]  ( .D(n4959), .CK(clk), .Q(\mem[208][5] ) );
  DFF_X1 \mem_reg[208][4]  ( .D(n4960), .CK(clk), .Q(\mem[208][4] ) );
  DFF_X1 \mem_reg[208][3]  ( .D(n4961), .CK(clk), .Q(\mem[208][3] ) );
  DFF_X1 \mem_reg[208][2]  ( .D(n4962), .CK(clk), .Q(\mem[208][2] ) );
  DFF_X1 \mem_reg[208][1]  ( .D(n4963), .CK(clk), .Q(\mem[208][1] ) );
  DFF_X1 \mem_reg[208][0]  ( .D(n4964), .CK(clk), .Q(\mem[208][0] ) );
  DFF_X1 \mem_reg[207][7]  ( .D(n4965), .CK(clk), .Q(\mem[207][7] ) );
  DFF_X1 \mem_reg[207][6]  ( .D(n4966), .CK(clk), .Q(\mem[207][6] ) );
  DFF_X1 \mem_reg[207][5]  ( .D(n4967), .CK(clk), .Q(\mem[207][5] ) );
  DFF_X1 \mem_reg[207][4]  ( .D(n4968), .CK(clk), .Q(\mem[207][4] ) );
  DFF_X1 \mem_reg[207][3]  ( .D(n4969), .CK(clk), .Q(\mem[207][3] ) );
  DFF_X1 \mem_reg[207][2]  ( .D(n4970), .CK(clk), .Q(\mem[207][2] ) );
  DFF_X1 \mem_reg[207][1]  ( .D(n4971), .CK(clk), .Q(\mem[207][1] ) );
  DFF_X1 \mem_reg[207][0]  ( .D(n4972), .CK(clk), .Q(\mem[207][0] ) );
  DFF_X1 \mem_reg[206][7]  ( .D(n4973), .CK(clk), .Q(\mem[206][7] ) );
  DFF_X1 \mem_reg[206][6]  ( .D(n4974), .CK(clk), .Q(\mem[206][6] ) );
  DFF_X1 \mem_reg[206][5]  ( .D(n4975), .CK(clk), .Q(\mem[206][5] ) );
  DFF_X1 \mem_reg[206][4]  ( .D(n4976), .CK(clk), .Q(\mem[206][4] ) );
  DFF_X1 \mem_reg[206][3]  ( .D(n4977), .CK(clk), .Q(\mem[206][3] ) );
  DFF_X1 \mem_reg[206][2]  ( .D(n4978), .CK(clk), .Q(\mem[206][2] ) );
  DFF_X1 \mem_reg[206][1]  ( .D(n4979), .CK(clk), .Q(\mem[206][1] ) );
  DFF_X1 \mem_reg[206][0]  ( .D(n4980), .CK(clk), .Q(\mem[206][0] ) );
  DFF_X1 \mem_reg[205][7]  ( .D(n4981), .CK(clk), .Q(\mem[205][7] ) );
  DFF_X1 \mem_reg[205][6]  ( .D(n4982), .CK(clk), .Q(\mem[205][6] ) );
  DFF_X1 \mem_reg[205][5]  ( .D(n4983), .CK(clk), .Q(\mem[205][5] ) );
  DFF_X1 \mem_reg[205][4]  ( .D(n4984), .CK(clk), .Q(\mem[205][4] ) );
  DFF_X1 \mem_reg[205][3]  ( .D(n4985), .CK(clk), .Q(\mem[205][3] ) );
  DFF_X1 \mem_reg[205][2]  ( .D(n4986), .CK(clk), .Q(\mem[205][2] ) );
  DFF_X1 \mem_reg[205][1]  ( .D(n4987), .CK(clk), .Q(\mem[205][1] ) );
  DFF_X1 \mem_reg[205][0]  ( .D(n4988), .CK(clk), .Q(\mem[205][0] ) );
  DFF_X1 \mem_reg[204][7]  ( .D(n4989), .CK(clk), .Q(\mem[204][7] ) );
  DFF_X1 \mem_reg[204][6]  ( .D(n4990), .CK(clk), .Q(\mem[204][6] ) );
  DFF_X1 \mem_reg[204][5]  ( .D(n4991), .CK(clk), .Q(\mem[204][5] ) );
  DFF_X1 \mem_reg[204][4]  ( .D(n4992), .CK(clk), .Q(\mem[204][4] ) );
  DFF_X1 \mem_reg[204][3]  ( .D(n4993), .CK(clk), .Q(\mem[204][3] ) );
  DFF_X1 \mem_reg[204][2]  ( .D(n4994), .CK(clk), .Q(\mem[204][2] ) );
  DFF_X1 \mem_reg[204][1]  ( .D(n4995), .CK(clk), .Q(\mem[204][1] ) );
  DFF_X1 \mem_reg[204][0]  ( .D(n4996), .CK(clk), .Q(\mem[204][0] ) );
  DFF_X1 \mem_reg[203][7]  ( .D(n4997), .CK(clk), .Q(\mem[203][7] ) );
  DFF_X1 \mem_reg[203][6]  ( .D(n4998), .CK(clk), .Q(\mem[203][6] ) );
  DFF_X1 \mem_reg[203][5]  ( .D(n4999), .CK(clk), .Q(\mem[203][5] ) );
  DFF_X1 \mem_reg[203][4]  ( .D(n5000), .CK(clk), .Q(\mem[203][4] ) );
  DFF_X1 \mem_reg[203][3]  ( .D(n5001), .CK(clk), .Q(\mem[203][3] ) );
  DFF_X1 \mem_reg[203][2]  ( .D(n5002), .CK(clk), .Q(\mem[203][2] ) );
  DFF_X1 \mem_reg[203][1]  ( .D(n5003), .CK(clk), .Q(\mem[203][1] ) );
  DFF_X1 \mem_reg[203][0]  ( .D(n5004), .CK(clk), .Q(\mem[203][0] ) );
  DFF_X1 \mem_reg[202][7]  ( .D(n5005), .CK(clk), .Q(\mem[202][7] ) );
  DFF_X1 \mem_reg[202][6]  ( .D(n5006), .CK(clk), .Q(\mem[202][6] ) );
  DFF_X1 \mem_reg[202][5]  ( .D(n5007), .CK(clk), .Q(\mem[202][5] ) );
  DFF_X1 \mem_reg[202][4]  ( .D(n5008), .CK(clk), .Q(\mem[202][4] ) );
  DFF_X1 \mem_reg[202][3]  ( .D(n5009), .CK(clk), .Q(\mem[202][3] ) );
  DFF_X1 \mem_reg[202][2]  ( .D(n5010), .CK(clk), .Q(\mem[202][2] ) );
  DFF_X1 \mem_reg[202][1]  ( .D(n5011), .CK(clk), .Q(\mem[202][1] ) );
  DFF_X1 \mem_reg[202][0]  ( .D(n5012), .CK(clk), .Q(\mem[202][0] ) );
  DFF_X1 \mem_reg[201][7]  ( .D(n5013), .CK(clk), .Q(\mem[201][7] ) );
  DFF_X1 \mem_reg[201][6]  ( .D(n5014), .CK(clk), .Q(\mem[201][6] ) );
  DFF_X1 \mem_reg[201][5]  ( .D(n5015), .CK(clk), .Q(\mem[201][5] ) );
  DFF_X1 \mem_reg[201][4]  ( .D(n5016), .CK(clk), .Q(\mem[201][4] ) );
  DFF_X1 \mem_reg[201][3]  ( .D(n5017), .CK(clk), .Q(\mem[201][3] ) );
  DFF_X1 \mem_reg[201][2]  ( .D(n5018), .CK(clk), .Q(\mem[201][2] ) );
  DFF_X1 \mem_reg[201][1]  ( .D(n5019), .CK(clk), .Q(\mem[201][1] ) );
  DFF_X1 \mem_reg[201][0]  ( .D(n5020), .CK(clk), .Q(\mem[201][0] ) );
  DFF_X1 \mem_reg[200][7]  ( .D(n5021), .CK(clk), .Q(\mem[200][7] ) );
  DFF_X1 \mem_reg[200][6]  ( .D(n5022), .CK(clk), .Q(\mem[200][6] ) );
  DFF_X1 \mem_reg[200][5]  ( .D(n5023), .CK(clk), .Q(\mem[200][5] ) );
  DFF_X1 \mem_reg[200][4]  ( .D(n5024), .CK(clk), .Q(\mem[200][4] ) );
  DFF_X1 \mem_reg[200][3]  ( .D(n5025), .CK(clk), .Q(\mem[200][3] ) );
  DFF_X1 \mem_reg[200][2]  ( .D(n5026), .CK(clk), .Q(\mem[200][2] ) );
  DFF_X1 \mem_reg[200][1]  ( .D(n5027), .CK(clk), .Q(\mem[200][1] ) );
  DFF_X1 \mem_reg[200][0]  ( .D(n5028), .CK(clk), .Q(\mem[200][0] ) );
  DFF_X1 \mem_reg[199][7]  ( .D(n5029), .CK(clk), .Q(\mem[199][7] ) );
  DFF_X1 \mem_reg[199][6]  ( .D(n5030), .CK(clk), .Q(\mem[199][6] ) );
  DFF_X1 \mem_reg[199][5]  ( .D(n5031), .CK(clk), .Q(\mem[199][5] ) );
  DFF_X1 \mem_reg[199][4]  ( .D(n5032), .CK(clk), .Q(\mem[199][4] ) );
  DFF_X1 \mem_reg[199][3]  ( .D(n5033), .CK(clk), .Q(\mem[199][3] ) );
  DFF_X1 \mem_reg[199][2]  ( .D(n5034), .CK(clk), .Q(\mem[199][2] ) );
  DFF_X1 \mem_reg[199][1]  ( .D(n5035), .CK(clk), .Q(\mem[199][1] ) );
  DFF_X1 \mem_reg[199][0]  ( .D(n5036), .CK(clk), .Q(\mem[199][0] ) );
  DFF_X1 \mem_reg[198][7]  ( .D(n5037), .CK(clk), .Q(\mem[198][7] ) );
  DFF_X1 \mem_reg[198][6]  ( .D(n5038), .CK(clk), .Q(\mem[198][6] ) );
  DFF_X1 \mem_reg[198][5]  ( .D(n5039), .CK(clk), .Q(\mem[198][5] ) );
  DFF_X1 \mem_reg[198][4]  ( .D(n5040), .CK(clk), .Q(\mem[198][4] ) );
  DFF_X1 \mem_reg[198][3]  ( .D(n5041), .CK(clk), .Q(\mem[198][3] ) );
  DFF_X1 \mem_reg[198][2]  ( .D(n5042), .CK(clk), .Q(\mem[198][2] ) );
  DFF_X1 \mem_reg[198][1]  ( .D(n5043), .CK(clk), .Q(\mem[198][1] ) );
  DFF_X1 \mem_reg[198][0]  ( .D(n5044), .CK(clk), .Q(\mem[198][0] ) );
  DFF_X1 \mem_reg[197][7]  ( .D(n5045), .CK(clk), .Q(\mem[197][7] ) );
  DFF_X1 \mem_reg[197][6]  ( .D(n5046), .CK(clk), .Q(\mem[197][6] ) );
  DFF_X1 \mem_reg[197][5]  ( .D(n5047), .CK(clk), .Q(\mem[197][5] ) );
  DFF_X1 \mem_reg[197][4]  ( .D(n5048), .CK(clk), .Q(\mem[197][4] ) );
  DFF_X1 \mem_reg[197][3]  ( .D(n5049), .CK(clk), .Q(\mem[197][3] ) );
  DFF_X1 \mem_reg[197][2]  ( .D(n5050), .CK(clk), .Q(\mem[197][2] ) );
  DFF_X1 \mem_reg[197][1]  ( .D(n5051), .CK(clk), .Q(\mem[197][1] ) );
  DFF_X1 \mem_reg[197][0]  ( .D(n5052), .CK(clk), .Q(\mem[197][0] ) );
  DFF_X1 \mem_reg[196][7]  ( .D(n5053), .CK(clk), .Q(\mem[196][7] ) );
  DFF_X1 \mem_reg[196][6]  ( .D(n5054), .CK(clk), .Q(\mem[196][6] ) );
  DFF_X1 \mem_reg[196][5]  ( .D(n5055), .CK(clk), .Q(\mem[196][5] ) );
  DFF_X1 \mem_reg[196][4]  ( .D(n5056), .CK(clk), .Q(\mem[196][4] ) );
  DFF_X1 \mem_reg[196][3]  ( .D(n5057), .CK(clk), .Q(\mem[196][3] ) );
  DFF_X1 \mem_reg[196][2]  ( .D(n5058), .CK(clk), .Q(\mem[196][2] ) );
  DFF_X1 \mem_reg[196][1]  ( .D(n5059), .CK(clk), .Q(\mem[196][1] ) );
  DFF_X1 \mem_reg[196][0]  ( .D(n5060), .CK(clk), .Q(\mem[196][0] ) );
  DFF_X1 \mem_reg[195][7]  ( .D(n5061), .CK(clk), .Q(\mem[195][7] ) );
  DFF_X1 \mem_reg[195][6]  ( .D(n5062), .CK(clk), .Q(\mem[195][6] ) );
  DFF_X1 \mem_reg[195][5]  ( .D(n5063), .CK(clk), .Q(\mem[195][5] ) );
  DFF_X1 \mem_reg[195][4]  ( .D(n5064), .CK(clk), .Q(\mem[195][4] ) );
  DFF_X1 \mem_reg[195][3]  ( .D(n5065), .CK(clk), .Q(\mem[195][3] ) );
  DFF_X1 \mem_reg[195][2]  ( .D(n5066), .CK(clk), .Q(\mem[195][2] ) );
  DFF_X1 \mem_reg[195][1]  ( .D(n5067), .CK(clk), .Q(\mem[195][1] ) );
  DFF_X1 \mem_reg[195][0]  ( .D(n5068), .CK(clk), .Q(\mem[195][0] ) );
  DFF_X1 \mem_reg[194][7]  ( .D(n5069), .CK(clk), .Q(\mem[194][7] ) );
  DFF_X1 \mem_reg[194][6]  ( .D(n5070), .CK(clk), .Q(\mem[194][6] ) );
  DFF_X1 \mem_reg[194][5]  ( .D(n5071), .CK(clk), .Q(\mem[194][5] ) );
  DFF_X1 \mem_reg[194][4]  ( .D(n5072), .CK(clk), .Q(\mem[194][4] ) );
  DFF_X1 \mem_reg[194][3]  ( .D(n5073), .CK(clk), .Q(\mem[194][3] ) );
  DFF_X1 \mem_reg[194][2]  ( .D(n5074), .CK(clk), .Q(\mem[194][2] ) );
  DFF_X1 \mem_reg[194][1]  ( .D(n5075), .CK(clk), .Q(\mem[194][1] ) );
  DFF_X1 \mem_reg[194][0]  ( .D(n5076), .CK(clk), .Q(\mem[194][0] ) );
  DFF_X1 \mem_reg[193][7]  ( .D(n5077), .CK(clk), .Q(\mem[193][7] ) );
  DFF_X1 \mem_reg[193][6]  ( .D(n5078), .CK(clk), .Q(\mem[193][6] ) );
  DFF_X1 \mem_reg[193][5]  ( .D(n5079), .CK(clk), .Q(\mem[193][5] ) );
  DFF_X1 \mem_reg[193][4]  ( .D(n5080), .CK(clk), .Q(\mem[193][4] ) );
  DFF_X1 \mem_reg[193][3]  ( .D(n5081), .CK(clk), .Q(\mem[193][3] ) );
  DFF_X1 \mem_reg[193][2]  ( .D(n5082), .CK(clk), .Q(\mem[193][2] ) );
  DFF_X1 \mem_reg[193][1]  ( .D(n5083), .CK(clk), .Q(\mem[193][1] ) );
  DFF_X1 \mem_reg[193][0]  ( .D(n5084), .CK(clk), .Q(\mem[193][0] ) );
  DFF_X1 \mem_reg[192][7]  ( .D(n5085), .CK(clk), .Q(\mem[192][7] ) );
  DFF_X1 \mem_reg[192][6]  ( .D(n5086), .CK(clk), .Q(\mem[192][6] ) );
  DFF_X1 \mem_reg[192][5]  ( .D(n5087), .CK(clk), .Q(\mem[192][5] ) );
  DFF_X1 \mem_reg[192][4]  ( .D(n5088), .CK(clk), .Q(\mem[192][4] ) );
  DFF_X1 \mem_reg[192][3]  ( .D(n5089), .CK(clk), .Q(\mem[192][3] ) );
  DFF_X1 \mem_reg[192][2]  ( .D(n5090), .CK(clk), .Q(\mem[192][2] ) );
  DFF_X1 \mem_reg[192][1]  ( .D(n5091), .CK(clk), .Q(\mem[192][1] ) );
  DFF_X1 \mem_reg[192][0]  ( .D(n5092), .CK(clk), .Q(\mem[192][0] ) );
  DFF_X1 \mem_reg[191][7]  ( .D(n5093), .CK(clk), .Q(\mem[191][7] ) );
  DFF_X1 \mem_reg[191][6]  ( .D(n5094), .CK(clk), .Q(\mem[191][6] ) );
  DFF_X1 \mem_reg[191][5]  ( .D(n5095), .CK(clk), .Q(\mem[191][5] ) );
  DFF_X1 \mem_reg[191][4]  ( .D(n5096), .CK(clk), .Q(\mem[191][4] ) );
  DFF_X1 \mem_reg[191][3]  ( .D(n5097), .CK(clk), .Q(\mem[191][3] ) );
  DFF_X1 \mem_reg[191][2]  ( .D(n5098), .CK(clk), .Q(\mem[191][2] ) );
  DFF_X1 \mem_reg[191][1]  ( .D(n5099), .CK(clk), .Q(\mem[191][1] ) );
  DFF_X1 \mem_reg[191][0]  ( .D(n5100), .CK(clk), .Q(\mem[191][0] ) );
  DFF_X1 \mem_reg[190][7]  ( .D(n5101), .CK(clk), .Q(\mem[190][7] ) );
  DFF_X1 \mem_reg[190][6]  ( .D(n5102), .CK(clk), .Q(\mem[190][6] ) );
  DFF_X1 \mem_reg[190][5]  ( .D(n5103), .CK(clk), .Q(\mem[190][5] ) );
  DFF_X1 \mem_reg[190][4]  ( .D(n5104), .CK(clk), .Q(\mem[190][4] ) );
  DFF_X1 \mem_reg[190][3]  ( .D(n5105), .CK(clk), .Q(\mem[190][3] ) );
  DFF_X1 \mem_reg[190][2]  ( .D(n5106), .CK(clk), .Q(\mem[190][2] ) );
  DFF_X1 \mem_reg[190][1]  ( .D(n5107), .CK(clk), .Q(\mem[190][1] ) );
  DFF_X1 \mem_reg[190][0]  ( .D(n5108), .CK(clk), .Q(\mem[190][0] ) );
  DFF_X1 \mem_reg[189][7]  ( .D(n5109), .CK(clk), .Q(\mem[189][7] ) );
  DFF_X1 \mem_reg[189][6]  ( .D(n5110), .CK(clk), .Q(\mem[189][6] ) );
  DFF_X1 \mem_reg[189][5]  ( .D(n5111), .CK(clk), .Q(\mem[189][5] ) );
  DFF_X1 \mem_reg[189][4]  ( .D(n5112), .CK(clk), .Q(\mem[189][4] ) );
  DFF_X1 \mem_reg[189][3]  ( .D(n5113), .CK(clk), .Q(\mem[189][3] ) );
  DFF_X1 \mem_reg[189][2]  ( .D(n5114), .CK(clk), .Q(\mem[189][2] ) );
  DFF_X1 \mem_reg[189][1]  ( .D(n5115), .CK(clk), .Q(\mem[189][1] ) );
  DFF_X1 \mem_reg[189][0]  ( .D(n5116), .CK(clk), .Q(\mem[189][0] ) );
  DFF_X1 \mem_reg[188][7]  ( .D(n5117), .CK(clk), .Q(\mem[188][7] ) );
  DFF_X1 \mem_reg[188][6]  ( .D(n5118), .CK(clk), .Q(\mem[188][6] ) );
  DFF_X1 \mem_reg[188][5]  ( .D(n5119), .CK(clk), .Q(\mem[188][5] ) );
  DFF_X1 \mem_reg[188][4]  ( .D(n5120), .CK(clk), .Q(\mem[188][4] ) );
  DFF_X1 \mem_reg[188][3]  ( .D(n5121), .CK(clk), .Q(\mem[188][3] ) );
  DFF_X1 \mem_reg[188][2]  ( .D(n5122), .CK(clk), .Q(\mem[188][2] ) );
  DFF_X1 \mem_reg[188][1]  ( .D(n5123), .CK(clk), .Q(\mem[188][1] ) );
  DFF_X1 \mem_reg[188][0]  ( .D(n5124), .CK(clk), .Q(\mem[188][0] ) );
  DFF_X1 \mem_reg[187][7]  ( .D(n5125), .CK(clk), .Q(\mem[187][7] ) );
  DFF_X1 \mem_reg[187][6]  ( .D(n5126), .CK(clk), .Q(\mem[187][6] ) );
  DFF_X1 \mem_reg[187][5]  ( .D(n5127), .CK(clk), .Q(\mem[187][5] ) );
  DFF_X1 \mem_reg[187][4]  ( .D(n5128), .CK(clk), .Q(\mem[187][4] ) );
  DFF_X1 \mem_reg[187][3]  ( .D(n5129), .CK(clk), .Q(\mem[187][3] ) );
  DFF_X1 \mem_reg[187][2]  ( .D(n5130), .CK(clk), .Q(\mem[187][2] ) );
  DFF_X1 \mem_reg[187][1]  ( .D(n5131), .CK(clk), .Q(\mem[187][1] ) );
  DFF_X1 \mem_reg[187][0]  ( .D(n5132), .CK(clk), .Q(\mem[187][0] ) );
  DFF_X1 \mem_reg[186][7]  ( .D(n5133), .CK(clk), .Q(\mem[186][7] ) );
  DFF_X1 \mem_reg[186][6]  ( .D(n5134), .CK(clk), .Q(\mem[186][6] ) );
  DFF_X1 \mem_reg[186][5]  ( .D(n5135), .CK(clk), .Q(\mem[186][5] ) );
  DFF_X1 \mem_reg[186][4]  ( .D(n5136), .CK(clk), .Q(\mem[186][4] ) );
  DFF_X1 \mem_reg[186][3]  ( .D(n5137), .CK(clk), .Q(\mem[186][3] ) );
  DFF_X1 \mem_reg[186][2]  ( .D(n5138), .CK(clk), .Q(\mem[186][2] ) );
  DFF_X1 \mem_reg[186][1]  ( .D(n5139), .CK(clk), .Q(\mem[186][1] ) );
  DFF_X1 \mem_reg[186][0]  ( .D(n5140), .CK(clk), .Q(\mem[186][0] ) );
  DFF_X1 \mem_reg[185][7]  ( .D(n5141), .CK(clk), .Q(\mem[185][7] ) );
  DFF_X1 \mem_reg[185][6]  ( .D(n5142), .CK(clk), .Q(\mem[185][6] ) );
  DFF_X1 \mem_reg[185][5]  ( .D(n5143), .CK(clk), .Q(\mem[185][5] ) );
  DFF_X1 \mem_reg[185][4]  ( .D(n5144), .CK(clk), .Q(\mem[185][4] ) );
  DFF_X1 \mem_reg[185][3]  ( .D(n5145), .CK(clk), .Q(\mem[185][3] ) );
  DFF_X1 \mem_reg[185][2]  ( .D(n5146), .CK(clk), .Q(\mem[185][2] ) );
  DFF_X1 \mem_reg[185][1]  ( .D(n5147), .CK(clk), .Q(\mem[185][1] ) );
  DFF_X1 \mem_reg[185][0]  ( .D(n5148), .CK(clk), .Q(\mem[185][0] ) );
  DFF_X1 \mem_reg[184][7]  ( .D(n5149), .CK(clk), .Q(\mem[184][7] ) );
  DFF_X1 \mem_reg[184][6]  ( .D(n5150), .CK(clk), .Q(\mem[184][6] ) );
  DFF_X1 \mem_reg[184][5]  ( .D(n5151), .CK(clk), .Q(\mem[184][5] ) );
  DFF_X1 \mem_reg[184][4]  ( .D(n5152), .CK(clk), .Q(\mem[184][4] ) );
  DFF_X1 \mem_reg[184][3]  ( .D(n5153), .CK(clk), .Q(\mem[184][3] ) );
  DFF_X1 \mem_reg[184][2]  ( .D(n5154), .CK(clk), .Q(\mem[184][2] ) );
  DFF_X1 \mem_reg[184][1]  ( .D(n5155), .CK(clk), .Q(\mem[184][1] ) );
  DFF_X1 \mem_reg[184][0]  ( .D(n5156), .CK(clk), .Q(\mem[184][0] ) );
  DFF_X1 \mem_reg[183][7]  ( .D(n5157), .CK(clk), .Q(\mem[183][7] ) );
  DFF_X1 \mem_reg[183][6]  ( .D(n5158), .CK(clk), .Q(\mem[183][6] ) );
  DFF_X1 \mem_reg[183][5]  ( .D(n5159), .CK(clk), .Q(\mem[183][5] ) );
  DFF_X1 \mem_reg[183][4]  ( .D(n5160), .CK(clk), .Q(\mem[183][4] ) );
  DFF_X1 \mem_reg[183][3]  ( .D(n5161), .CK(clk), .Q(\mem[183][3] ) );
  DFF_X1 \mem_reg[183][2]  ( .D(n5162), .CK(clk), .Q(\mem[183][2] ) );
  DFF_X1 \mem_reg[183][1]  ( .D(n5163), .CK(clk), .Q(\mem[183][1] ) );
  DFF_X1 \mem_reg[183][0]  ( .D(n5164), .CK(clk), .Q(\mem[183][0] ) );
  DFF_X1 \mem_reg[182][7]  ( .D(n5165), .CK(clk), .Q(\mem[182][7] ) );
  DFF_X1 \mem_reg[182][6]  ( .D(n5166), .CK(clk), .Q(\mem[182][6] ) );
  DFF_X1 \mem_reg[182][5]  ( .D(n5167), .CK(clk), .Q(\mem[182][5] ) );
  DFF_X1 \mem_reg[182][4]  ( .D(n5168), .CK(clk), .Q(\mem[182][4] ) );
  DFF_X1 \mem_reg[182][3]  ( .D(n5169), .CK(clk), .Q(\mem[182][3] ) );
  DFF_X1 \mem_reg[182][2]  ( .D(n5170), .CK(clk), .Q(\mem[182][2] ) );
  DFF_X1 \mem_reg[182][1]  ( .D(n5171), .CK(clk), .Q(\mem[182][1] ) );
  DFF_X1 \mem_reg[182][0]  ( .D(n5172), .CK(clk), .Q(\mem[182][0] ) );
  DFF_X1 \mem_reg[181][7]  ( .D(n5173), .CK(clk), .Q(\mem[181][7] ) );
  DFF_X1 \mem_reg[181][6]  ( .D(n5174), .CK(clk), .Q(\mem[181][6] ) );
  DFF_X1 \mem_reg[181][5]  ( .D(n5175), .CK(clk), .Q(\mem[181][5] ) );
  DFF_X1 \mem_reg[181][4]  ( .D(n5176), .CK(clk), .Q(\mem[181][4] ) );
  DFF_X1 \mem_reg[181][3]  ( .D(n5177), .CK(clk), .Q(\mem[181][3] ) );
  DFF_X1 \mem_reg[181][2]  ( .D(n5178), .CK(clk), .Q(\mem[181][2] ) );
  DFF_X1 \mem_reg[181][1]  ( .D(n5179), .CK(clk), .Q(\mem[181][1] ) );
  DFF_X1 \mem_reg[181][0]  ( .D(n5180), .CK(clk), .Q(\mem[181][0] ) );
  DFF_X1 \mem_reg[180][7]  ( .D(n5181), .CK(clk), .Q(\mem[180][7] ) );
  DFF_X1 \mem_reg[180][6]  ( .D(n5182), .CK(clk), .Q(\mem[180][6] ) );
  DFF_X1 \mem_reg[180][5]  ( .D(n5183), .CK(clk), .Q(\mem[180][5] ) );
  DFF_X1 \mem_reg[180][4]  ( .D(n5184), .CK(clk), .Q(\mem[180][4] ) );
  DFF_X1 \mem_reg[180][3]  ( .D(n5185), .CK(clk), .Q(\mem[180][3] ) );
  DFF_X1 \mem_reg[180][2]  ( .D(n5186), .CK(clk), .Q(\mem[180][2] ) );
  DFF_X1 \mem_reg[180][1]  ( .D(n5187), .CK(clk), .Q(\mem[180][1] ) );
  DFF_X1 \mem_reg[180][0]  ( .D(n5188), .CK(clk), .Q(\mem[180][0] ) );
  DFF_X1 \mem_reg[179][7]  ( .D(n5189), .CK(clk), .Q(\mem[179][7] ) );
  DFF_X1 \mem_reg[179][6]  ( .D(n5190), .CK(clk), .Q(\mem[179][6] ) );
  DFF_X1 \mem_reg[179][5]  ( .D(n5191), .CK(clk), .Q(\mem[179][5] ) );
  DFF_X1 \mem_reg[179][4]  ( .D(n5192), .CK(clk), .Q(\mem[179][4] ) );
  DFF_X1 \mem_reg[179][3]  ( .D(n5193), .CK(clk), .Q(\mem[179][3] ) );
  DFF_X1 \mem_reg[179][2]  ( .D(n5194), .CK(clk), .Q(\mem[179][2] ) );
  DFF_X1 \mem_reg[179][1]  ( .D(n5195), .CK(clk), .Q(\mem[179][1] ) );
  DFF_X1 \mem_reg[179][0]  ( .D(n5196), .CK(clk), .Q(\mem[179][0] ) );
  DFF_X1 \mem_reg[178][7]  ( .D(n5197), .CK(clk), .Q(\mem[178][7] ) );
  DFF_X1 \mem_reg[178][6]  ( .D(n5198), .CK(clk), .Q(\mem[178][6] ) );
  DFF_X1 \mem_reg[178][5]  ( .D(n5199), .CK(clk), .Q(\mem[178][5] ) );
  DFF_X1 \mem_reg[178][4]  ( .D(n5200), .CK(clk), .Q(\mem[178][4] ) );
  DFF_X1 \mem_reg[178][3]  ( .D(n5201), .CK(clk), .Q(\mem[178][3] ) );
  DFF_X1 \mem_reg[178][2]  ( .D(n5202), .CK(clk), .Q(\mem[178][2] ) );
  DFF_X1 \mem_reg[178][1]  ( .D(n5203), .CK(clk), .Q(\mem[178][1] ) );
  DFF_X1 \mem_reg[178][0]  ( .D(n5204), .CK(clk), .Q(\mem[178][0] ) );
  DFF_X1 \mem_reg[177][7]  ( .D(n5205), .CK(clk), .Q(\mem[177][7] ) );
  DFF_X1 \mem_reg[177][6]  ( .D(n5206), .CK(clk), .Q(\mem[177][6] ) );
  DFF_X1 \mem_reg[177][5]  ( .D(n5207), .CK(clk), .Q(\mem[177][5] ) );
  DFF_X1 \mem_reg[177][4]  ( .D(n5208), .CK(clk), .Q(\mem[177][4] ) );
  DFF_X1 \mem_reg[177][3]  ( .D(n5209), .CK(clk), .Q(\mem[177][3] ) );
  DFF_X1 \mem_reg[177][2]  ( .D(n5210), .CK(clk), .Q(\mem[177][2] ) );
  DFF_X1 \mem_reg[177][1]  ( .D(n5211), .CK(clk), .Q(\mem[177][1] ) );
  DFF_X1 \mem_reg[177][0]  ( .D(n5212), .CK(clk), .Q(\mem[177][0] ) );
  DFF_X1 \mem_reg[176][7]  ( .D(n5213), .CK(clk), .Q(\mem[176][7] ) );
  DFF_X1 \mem_reg[176][6]  ( .D(n5214), .CK(clk), .Q(\mem[176][6] ) );
  DFF_X1 \mem_reg[176][5]  ( .D(n5215), .CK(clk), .Q(\mem[176][5] ) );
  DFF_X1 \mem_reg[176][4]  ( .D(n5216), .CK(clk), .Q(\mem[176][4] ) );
  DFF_X1 \mem_reg[176][3]  ( .D(n5217), .CK(clk), .Q(\mem[176][3] ) );
  DFF_X1 \mem_reg[176][2]  ( .D(n5218), .CK(clk), .Q(\mem[176][2] ) );
  DFF_X1 \mem_reg[176][1]  ( .D(n5219), .CK(clk), .Q(\mem[176][1] ) );
  DFF_X1 \mem_reg[176][0]  ( .D(n5220), .CK(clk), .Q(\mem[176][0] ) );
  DFF_X1 \mem_reg[175][7]  ( .D(n5221), .CK(clk), .Q(\mem[175][7] ) );
  DFF_X1 \mem_reg[175][6]  ( .D(n5222), .CK(clk), .Q(\mem[175][6] ) );
  DFF_X1 \mem_reg[175][5]  ( .D(n5223), .CK(clk), .Q(\mem[175][5] ) );
  DFF_X1 \mem_reg[175][4]  ( .D(n5224), .CK(clk), .Q(\mem[175][4] ) );
  DFF_X1 \mem_reg[175][3]  ( .D(n5225), .CK(clk), .Q(\mem[175][3] ) );
  DFF_X1 \mem_reg[175][2]  ( .D(n5226), .CK(clk), .Q(\mem[175][2] ) );
  DFF_X1 \mem_reg[175][1]  ( .D(n5227), .CK(clk), .Q(\mem[175][1] ) );
  DFF_X1 \mem_reg[175][0]  ( .D(n5228), .CK(clk), .Q(\mem[175][0] ) );
  DFF_X1 \mem_reg[174][7]  ( .D(n5229), .CK(clk), .Q(\mem[174][7] ) );
  DFF_X1 \mem_reg[174][6]  ( .D(n5230), .CK(clk), .Q(\mem[174][6] ) );
  DFF_X1 \mem_reg[174][5]  ( .D(n5231), .CK(clk), .Q(\mem[174][5] ) );
  DFF_X1 \mem_reg[174][4]  ( .D(n5232), .CK(clk), .Q(\mem[174][4] ) );
  DFF_X1 \mem_reg[174][3]  ( .D(n5233), .CK(clk), .Q(\mem[174][3] ) );
  DFF_X1 \mem_reg[174][2]  ( .D(n5234), .CK(clk), .Q(\mem[174][2] ) );
  DFF_X1 \mem_reg[174][1]  ( .D(n5235), .CK(clk), .Q(\mem[174][1] ) );
  DFF_X1 \mem_reg[174][0]  ( .D(n5236), .CK(clk), .Q(\mem[174][0] ) );
  DFF_X1 \mem_reg[173][7]  ( .D(n5237), .CK(clk), .Q(\mem[173][7] ) );
  DFF_X1 \mem_reg[173][6]  ( .D(n5238), .CK(clk), .Q(\mem[173][6] ) );
  DFF_X1 \mem_reg[173][5]  ( .D(n5239), .CK(clk), .Q(\mem[173][5] ) );
  DFF_X1 \mem_reg[173][4]  ( .D(n5240), .CK(clk), .Q(\mem[173][4] ) );
  DFF_X1 \mem_reg[173][3]  ( .D(n5241), .CK(clk), .Q(\mem[173][3] ) );
  DFF_X1 \mem_reg[173][2]  ( .D(n5242), .CK(clk), .Q(\mem[173][2] ) );
  DFF_X1 \mem_reg[173][1]  ( .D(n5243), .CK(clk), .Q(\mem[173][1] ) );
  DFF_X1 \mem_reg[173][0]  ( .D(n5244), .CK(clk), .Q(\mem[173][0] ) );
  DFF_X1 \mem_reg[172][7]  ( .D(n5245), .CK(clk), .Q(\mem[172][7] ) );
  DFF_X1 \mem_reg[172][6]  ( .D(n5246), .CK(clk), .Q(\mem[172][6] ) );
  DFF_X1 \mem_reg[172][5]  ( .D(n5247), .CK(clk), .Q(\mem[172][5] ) );
  DFF_X1 \mem_reg[172][4]  ( .D(n5248), .CK(clk), .Q(\mem[172][4] ) );
  DFF_X1 \mem_reg[172][3]  ( .D(n5249), .CK(clk), .Q(\mem[172][3] ) );
  DFF_X1 \mem_reg[172][2]  ( .D(n5250), .CK(clk), .Q(\mem[172][2] ) );
  DFF_X1 \mem_reg[172][1]  ( .D(n5251), .CK(clk), .Q(\mem[172][1] ) );
  DFF_X1 \mem_reg[172][0]  ( .D(n5252), .CK(clk), .Q(\mem[172][0] ) );
  DFF_X1 \mem_reg[171][7]  ( .D(n5253), .CK(clk), .Q(\mem[171][7] ) );
  DFF_X1 \mem_reg[171][6]  ( .D(n5254), .CK(clk), .Q(\mem[171][6] ) );
  DFF_X1 \mem_reg[171][5]  ( .D(n5255), .CK(clk), .Q(\mem[171][5] ) );
  DFF_X1 \mem_reg[171][4]  ( .D(n5256), .CK(clk), .Q(\mem[171][4] ) );
  DFF_X1 \mem_reg[171][3]  ( .D(n5257), .CK(clk), .Q(\mem[171][3] ) );
  DFF_X1 \mem_reg[171][2]  ( .D(n5258), .CK(clk), .Q(\mem[171][2] ) );
  DFF_X1 \mem_reg[171][1]  ( .D(n5259), .CK(clk), .Q(\mem[171][1] ) );
  DFF_X1 \mem_reg[171][0]  ( .D(n5260), .CK(clk), .Q(\mem[171][0] ) );
  DFF_X1 \mem_reg[170][7]  ( .D(n5261), .CK(clk), .Q(\mem[170][7] ) );
  DFF_X1 \mem_reg[170][6]  ( .D(n5262), .CK(clk), .Q(\mem[170][6] ) );
  DFF_X1 \mem_reg[170][5]  ( .D(n5263), .CK(clk), .Q(\mem[170][5] ) );
  DFF_X1 \mem_reg[170][4]  ( .D(n5264), .CK(clk), .Q(\mem[170][4] ) );
  DFF_X1 \mem_reg[170][3]  ( .D(n5265), .CK(clk), .Q(\mem[170][3] ) );
  DFF_X1 \mem_reg[170][2]  ( .D(n5266), .CK(clk), .Q(\mem[170][2] ) );
  DFF_X1 \mem_reg[170][1]  ( .D(n5267), .CK(clk), .Q(\mem[170][1] ) );
  DFF_X1 \mem_reg[170][0]  ( .D(n5268), .CK(clk), .Q(\mem[170][0] ) );
  DFF_X1 \mem_reg[169][7]  ( .D(n5269), .CK(clk), .Q(\mem[169][7] ) );
  DFF_X1 \mem_reg[169][6]  ( .D(n5270), .CK(clk), .Q(\mem[169][6] ) );
  DFF_X1 \mem_reg[169][5]  ( .D(n5271), .CK(clk), .Q(\mem[169][5] ) );
  DFF_X1 \mem_reg[169][4]  ( .D(n5272), .CK(clk), .Q(\mem[169][4] ) );
  DFF_X1 \mem_reg[169][3]  ( .D(n5273), .CK(clk), .Q(\mem[169][3] ) );
  DFF_X1 \mem_reg[169][2]  ( .D(n5274), .CK(clk), .Q(\mem[169][2] ) );
  DFF_X1 \mem_reg[169][1]  ( .D(n5275), .CK(clk), .Q(\mem[169][1] ) );
  DFF_X1 \mem_reg[169][0]  ( .D(n5276), .CK(clk), .Q(\mem[169][0] ) );
  DFF_X1 \mem_reg[168][7]  ( .D(n5277), .CK(clk), .Q(\mem[168][7] ) );
  DFF_X1 \mem_reg[168][6]  ( .D(n5278), .CK(clk), .Q(\mem[168][6] ) );
  DFF_X1 \mem_reg[168][5]  ( .D(n5279), .CK(clk), .Q(\mem[168][5] ) );
  DFF_X1 \mem_reg[168][4]  ( .D(n5280), .CK(clk), .Q(\mem[168][4] ) );
  DFF_X1 \mem_reg[168][3]  ( .D(n5281), .CK(clk), .Q(\mem[168][3] ) );
  DFF_X1 \mem_reg[168][2]  ( .D(n5282), .CK(clk), .Q(\mem[168][2] ) );
  DFF_X1 \mem_reg[168][1]  ( .D(n5283), .CK(clk), .Q(\mem[168][1] ) );
  DFF_X1 \mem_reg[168][0]  ( .D(n5284), .CK(clk), .Q(\mem[168][0] ) );
  DFF_X1 \mem_reg[167][7]  ( .D(n5285), .CK(clk), .Q(\mem[167][7] ) );
  DFF_X1 \mem_reg[167][6]  ( .D(n5286), .CK(clk), .Q(\mem[167][6] ) );
  DFF_X1 \mem_reg[167][5]  ( .D(n5287), .CK(clk), .Q(\mem[167][5] ) );
  DFF_X1 \mem_reg[167][4]  ( .D(n5288), .CK(clk), .Q(\mem[167][4] ) );
  DFF_X1 \mem_reg[167][3]  ( .D(n5289), .CK(clk), .Q(\mem[167][3] ) );
  DFF_X1 \mem_reg[167][2]  ( .D(n5290), .CK(clk), .Q(\mem[167][2] ) );
  DFF_X1 \mem_reg[167][1]  ( .D(n5291), .CK(clk), .Q(\mem[167][1] ) );
  DFF_X1 \mem_reg[167][0]  ( .D(n5292), .CK(clk), .Q(\mem[167][0] ) );
  DFF_X1 \mem_reg[166][7]  ( .D(n5293), .CK(clk), .Q(\mem[166][7] ) );
  DFF_X1 \mem_reg[166][6]  ( .D(n5294), .CK(clk), .Q(\mem[166][6] ) );
  DFF_X1 \mem_reg[166][5]  ( .D(n5295), .CK(clk), .Q(\mem[166][5] ) );
  DFF_X1 \mem_reg[166][4]  ( .D(n5296), .CK(clk), .Q(\mem[166][4] ) );
  DFF_X1 \mem_reg[166][3]  ( .D(n5297), .CK(clk), .Q(\mem[166][3] ) );
  DFF_X1 \mem_reg[166][2]  ( .D(n5298), .CK(clk), .Q(\mem[166][2] ) );
  DFF_X1 \mem_reg[166][1]  ( .D(n5299), .CK(clk), .Q(\mem[166][1] ) );
  DFF_X1 \mem_reg[166][0]  ( .D(n5300), .CK(clk), .Q(\mem[166][0] ) );
  DFF_X1 \mem_reg[165][7]  ( .D(n5301), .CK(clk), .Q(\mem[165][7] ) );
  DFF_X1 \mem_reg[165][6]  ( .D(n5302), .CK(clk), .Q(\mem[165][6] ) );
  DFF_X1 \mem_reg[165][5]  ( .D(n5303), .CK(clk), .Q(\mem[165][5] ) );
  DFF_X1 \mem_reg[165][4]  ( .D(n5304), .CK(clk), .Q(\mem[165][4] ) );
  DFF_X1 \mem_reg[165][3]  ( .D(n5305), .CK(clk), .Q(\mem[165][3] ) );
  DFF_X1 \mem_reg[165][2]  ( .D(n5306), .CK(clk), .Q(\mem[165][2] ) );
  DFF_X1 \mem_reg[165][1]  ( .D(n5307), .CK(clk), .Q(\mem[165][1] ) );
  DFF_X1 \mem_reg[165][0]  ( .D(n5308), .CK(clk), .Q(\mem[165][0] ) );
  DFF_X1 \mem_reg[164][7]  ( .D(n5309), .CK(clk), .Q(\mem[164][7] ) );
  DFF_X1 \mem_reg[164][6]  ( .D(n5310), .CK(clk), .Q(\mem[164][6] ) );
  DFF_X1 \mem_reg[164][5]  ( .D(n5311), .CK(clk), .Q(\mem[164][5] ) );
  DFF_X1 \mem_reg[164][4]  ( .D(n5312), .CK(clk), .Q(\mem[164][4] ) );
  DFF_X1 \mem_reg[164][3]  ( .D(n5313), .CK(clk), .Q(\mem[164][3] ) );
  DFF_X1 \mem_reg[164][2]  ( .D(n5314), .CK(clk), .Q(\mem[164][2] ) );
  DFF_X1 \mem_reg[164][1]  ( .D(n5315), .CK(clk), .Q(\mem[164][1] ) );
  DFF_X1 \mem_reg[164][0]  ( .D(n5316), .CK(clk), .Q(\mem[164][0] ) );
  DFF_X1 \mem_reg[163][7]  ( .D(n5317), .CK(clk), .Q(\mem[163][7] ) );
  DFF_X1 \mem_reg[163][6]  ( .D(n5318), .CK(clk), .Q(\mem[163][6] ) );
  DFF_X1 \mem_reg[163][5]  ( .D(n5319), .CK(clk), .Q(\mem[163][5] ) );
  DFF_X1 \mem_reg[163][4]  ( .D(n5320), .CK(clk), .Q(\mem[163][4] ) );
  DFF_X1 \mem_reg[163][3]  ( .D(n5321), .CK(clk), .Q(\mem[163][3] ) );
  DFF_X1 \mem_reg[163][2]  ( .D(n5322), .CK(clk), .Q(\mem[163][2] ) );
  DFF_X1 \mem_reg[163][1]  ( .D(n5323), .CK(clk), .Q(\mem[163][1] ) );
  DFF_X1 \mem_reg[163][0]  ( .D(n5324), .CK(clk), .Q(\mem[163][0] ) );
  DFF_X1 \mem_reg[162][7]  ( .D(n5325), .CK(clk), .Q(\mem[162][7] ) );
  DFF_X1 \mem_reg[162][6]  ( .D(n5326), .CK(clk), .Q(\mem[162][6] ) );
  DFF_X1 \mem_reg[162][5]  ( .D(n5327), .CK(clk), .Q(\mem[162][5] ) );
  DFF_X1 \mem_reg[162][4]  ( .D(n5328), .CK(clk), .Q(\mem[162][4] ) );
  DFF_X1 \mem_reg[162][3]  ( .D(n5329), .CK(clk), .Q(\mem[162][3] ) );
  DFF_X1 \mem_reg[162][2]  ( .D(n5330), .CK(clk), .Q(\mem[162][2] ) );
  DFF_X1 \mem_reg[162][1]  ( .D(n5331), .CK(clk), .Q(\mem[162][1] ) );
  DFF_X1 \mem_reg[162][0]  ( .D(n5332), .CK(clk), .Q(\mem[162][0] ) );
  DFF_X1 \mem_reg[161][7]  ( .D(n5333), .CK(clk), .Q(\mem[161][7] ) );
  DFF_X1 \mem_reg[161][6]  ( .D(n5334), .CK(clk), .Q(\mem[161][6] ) );
  DFF_X1 \mem_reg[161][5]  ( .D(n5335), .CK(clk), .Q(\mem[161][5] ) );
  DFF_X1 \mem_reg[161][4]  ( .D(n5336), .CK(clk), .Q(\mem[161][4] ) );
  DFF_X1 \mem_reg[161][3]  ( .D(n5337), .CK(clk), .Q(\mem[161][3] ) );
  DFF_X1 \mem_reg[161][2]  ( .D(n5338), .CK(clk), .Q(\mem[161][2] ) );
  DFF_X1 \mem_reg[161][1]  ( .D(n5339), .CK(clk), .Q(\mem[161][1] ) );
  DFF_X1 \mem_reg[161][0]  ( .D(n5340), .CK(clk), .Q(\mem[161][0] ) );
  DFF_X1 \mem_reg[160][7]  ( .D(n5341), .CK(clk), .Q(\mem[160][7] ) );
  DFF_X1 \mem_reg[160][6]  ( .D(n5342), .CK(clk), .Q(\mem[160][6] ) );
  DFF_X1 \mem_reg[160][5]  ( .D(n5343), .CK(clk), .Q(\mem[160][5] ) );
  DFF_X1 \mem_reg[160][4]  ( .D(n5344), .CK(clk), .Q(\mem[160][4] ) );
  DFF_X1 \mem_reg[160][3]  ( .D(n5345), .CK(clk), .Q(\mem[160][3] ) );
  DFF_X1 \mem_reg[160][2]  ( .D(n5346), .CK(clk), .Q(\mem[160][2] ) );
  DFF_X1 \mem_reg[160][1]  ( .D(n5347), .CK(clk), .Q(\mem[160][1] ) );
  DFF_X1 \mem_reg[160][0]  ( .D(n5348), .CK(clk), .Q(\mem[160][0] ) );
  DFF_X1 \mem_reg[159][7]  ( .D(n5349), .CK(clk), .Q(\mem[159][7] ) );
  DFF_X1 \mem_reg[159][6]  ( .D(n5350), .CK(clk), .Q(\mem[159][6] ) );
  DFF_X1 \mem_reg[159][5]  ( .D(n5351), .CK(clk), .Q(\mem[159][5] ) );
  DFF_X1 \mem_reg[159][4]  ( .D(n5352), .CK(clk), .Q(\mem[159][4] ) );
  DFF_X1 \mem_reg[159][3]  ( .D(n5353), .CK(clk), .Q(\mem[159][3] ) );
  DFF_X1 \mem_reg[159][2]  ( .D(n5354), .CK(clk), .Q(\mem[159][2] ) );
  DFF_X1 \mem_reg[159][1]  ( .D(n5355), .CK(clk), .Q(\mem[159][1] ) );
  DFF_X1 \mem_reg[159][0]  ( .D(n5356), .CK(clk), .Q(\mem[159][0] ) );
  DFF_X1 \mem_reg[158][7]  ( .D(n5357), .CK(clk), .Q(\mem[158][7] ) );
  DFF_X1 \mem_reg[158][6]  ( .D(n5358), .CK(clk), .Q(\mem[158][6] ) );
  DFF_X1 \mem_reg[158][5]  ( .D(n5359), .CK(clk), .Q(\mem[158][5] ) );
  DFF_X1 \mem_reg[158][4]  ( .D(n5360), .CK(clk), .Q(\mem[158][4] ) );
  DFF_X1 \mem_reg[158][3]  ( .D(n5361), .CK(clk), .Q(\mem[158][3] ) );
  DFF_X1 \mem_reg[158][2]  ( .D(n5362), .CK(clk), .Q(\mem[158][2] ) );
  DFF_X1 \mem_reg[158][1]  ( .D(n5363), .CK(clk), .Q(\mem[158][1] ) );
  DFF_X1 \mem_reg[158][0]  ( .D(n5364), .CK(clk), .Q(\mem[158][0] ) );
  DFF_X1 \mem_reg[157][7]  ( .D(n5365), .CK(clk), .Q(\mem[157][7] ) );
  DFF_X1 \mem_reg[157][6]  ( .D(n5366), .CK(clk), .Q(\mem[157][6] ) );
  DFF_X1 \mem_reg[157][5]  ( .D(n5367), .CK(clk), .Q(\mem[157][5] ) );
  DFF_X1 \mem_reg[157][4]  ( .D(n5368), .CK(clk), .Q(\mem[157][4] ) );
  DFF_X1 \mem_reg[157][3]  ( .D(n5369), .CK(clk), .Q(\mem[157][3] ) );
  DFF_X1 \mem_reg[157][2]  ( .D(n5370), .CK(clk), .Q(\mem[157][2] ) );
  DFF_X1 \mem_reg[157][1]  ( .D(n5371), .CK(clk), .Q(\mem[157][1] ) );
  DFF_X1 \mem_reg[157][0]  ( .D(n5372), .CK(clk), .Q(\mem[157][0] ) );
  DFF_X1 \mem_reg[156][7]  ( .D(n5373), .CK(clk), .Q(\mem[156][7] ) );
  DFF_X1 \mem_reg[156][6]  ( .D(n5374), .CK(clk), .Q(\mem[156][6] ) );
  DFF_X1 \mem_reg[156][5]  ( .D(n5375), .CK(clk), .Q(\mem[156][5] ) );
  DFF_X1 \mem_reg[156][4]  ( .D(n5376), .CK(clk), .Q(\mem[156][4] ) );
  DFF_X1 \mem_reg[156][3]  ( .D(n5377), .CK(clk), .Q(\mem[156][3] ) );
  DFF_X1 \mem_reg[156][2]  ( .D(n5378), .CK(clk), .Q(\mem[156][2] ) );
  DFF_X1 \mem_reg[156][1]  ( .D(n5379), .CK(clk), .Q(\mem[156][1] ) );
  DFF_X1 \mem_reg[156][0]  ( .D(n5380), .CK(clk), .Q(\mem[156][0] ) );
  DFF_X1 \mem_reg[155][7]  ( .D(n5381), .CK(clk), .Q(\mem[155][7] ) );
  DFF_X1 \mem_reg[155][6]  ( .D(n5382), .CK(clk), .Q(\mem[155][6] ) );
  DFF_X1 \mem_reg[155][5]  ( .D(n5383), .CK(clk), .Q(\mem[155][5] ) );
  DFF_X1 \mem_reg[155][4]  ( .D(n5384), .CK(clk), .Q(\mem[155][4] ) );
  DFF_X1 \mem_reg[155][3]  ( .D(n5385), .CK(clk), .Q(\mem[155][3] ) );
  DFF_X1 \mem_reg[155][2]  ( .D(n5386), .CK(clk), .Q(\mem[155][2] ) );
  DFF_X1 \mem_reg[155][1]  ( .D(n5387), .CK(clk), .Q(\mem[155][1] ) );
  DFF_X1 \mem_reg[155][0]  ( .D(n5388), .CK(clk), .Q(\mem[155][0] ) );
  DFF_X1 \mem_reg[154][7]  ( .D(n5389), .CK(clk), .Q(\mem[154][7] ) );
  DFF_X1 \mem_reg[154][6]  ( .D(n5390), .CK(clk), .Q(\mem[154][6] ) );
  DFF_X1 \mem_reg[154][5]  ( .D(n5391), .CK(clk), .Q(\mem[154][5] ) );
  DFF_X1 \mem_reg[154][4]  ( .D(n5392), .CK(clk), .Q(\mem[154][4] ) );
  DFF_X1 \mem_reg[154][3]  ( .D(n5393), .CK(clk), .Q(\mem[154][3] ) );
  DFF_X1 \mem_reg[154][2]  ( .D(n5394), .CK(clk), .Q(\mem[154][2] ) );
  DFF_X1 \mem_reg[154][1]  ( .D(n5395), .CK(clk), .Q(\mem[154][1] ) );
  DFF_X1 \mem_reg[154][0]  ( .D(n5396), .CK(clk), .Q(\mem[154][0] ) );
  DFF_X1 \mem_reg[153][7]  ( .D(n5397), .CK(clk), .Q(\mem[153][7] ) );
  DFF_X1 \mem_reg[153][6]  ( .D(n5398), .CK(clk), .Q(\mem[153][6] ) );
  DFF_X1 \mem_reg[153][5]  ( .D(n5399), .CK(clk), .Q(\mem[153][5] ) );
  DFF_X1 \mem_reg[153][4]  ( .D(n5400), .CK(clk), .Q(\mem[153][4] ) );
  DFF_X1 \mem_reg[153][3]  ( .D(n5401), .CK(clk), .Q(\mem[153][3] ) );
  DFF_X1 \mem_reg[153][2]  ( .D(n5402), .CK(clk), .Q(\mem[153][2] ) );
  DFF_X1 \mem_reg[153][1]  ( .D(n5403), .CK(clk), .Q(\mem[153][1] ) );
  DFF_X1 \mem_reg[153][0]  ( .D(n5404), .CK(clk), .Q(\mem[153][0] ) );
  DFF_X1 \mem_reg[152][7]  ( .D(n5405), .CK(clk), .Q(\mem[152][7] ) );
  DFF_X1 \mem_reg[152][6]  ( .D(n5406), .CK(clk), .Q(\mem[152][6] ) );
  DFF_X1 \mem_reg[152][5]  ( .D(n5407), .CK(clk), .Q(\mem[152][5] ) );
  DFF_X1 \mem_reg[152][4]  ( .D(n5408), .CK(clk), .Q(\mem[152][4] ) );
  DFF_X1 \mem_reg[152][3]  ( .D(n5409), .CK(clk), .Q(\mem[152][3] ) );
  DFF_X1 \mem_reg[152][2]  ( .D(n5410), .CK(clk), .Q(\mem[152][2] ) );
  DFF_X1 \mem_reg[152][1]  ( .D(n5411), .CK(clk), .Q(\mem[152][1] ) );
  DFF_X1 \mem_reg[152][0]  ( .D(n5412), .CK(clk), .Q(\mem[152][0] ) );
  DFF_X1 \mem_reg[151][7]  ( .D(n5413), .CK(clk), .Q(\mem[151][7] ) );
  DFF_X1 \mem_reg[151][6]  ( .D(n5414), .CK(clk), .Q(\mem[151][6] ) );
  DFF_X1 \mem_reg[151][5]  ( .D(n5415), .CK(clk), .Q(\mem[151][5] ) );
  DFF_X1 \mem_reg[151][4]  ( .D(n5416), .CK(clk), .Q(\mem[151][4] ) );
  DFF_X1 \mem_reg[151][3]  ( .D(n5417), .CK(clk), .Q(\mem[151][3] ) );
  DFF_X1 \mem_reg[151][2]  ( .D(n5418), .CK(clk), .Q(\mem[151][2] ) );
  DFF_X1 \mem_reg[151][1]  ( .D(n5419), .CK(clk), .Q(\mem[151][1] ) );
  DFF_X1 \mem_reg[151][0]  ( .D(n5420), .CK(clk), .Q(\mem[151][0] ) );
  DFF_X1 \mem_reg[150][7]  ( .D(n5421), .CK(clk), .Q(\mem[150][7] ) );
  DFF_X1 \mem_reg[150][6]  ( .D(n5422), .CK(clk), .Q(\mem[150][6] ) );
  DFF_X1 \mem_reg[150][5]  ( .D(n5423), .CK(clk), .Q(\mem[150][5] ) );
  DFF_X1 \mem_reg[150][4]  ( .D(n5424), .CK(clk), .Q(\mem[150][4] ) );
  DFF_X1 \mem_reg[150][3]  ( .D(n5425), .CK(clk), .Q(\mem[150][3] ) );
  DFF_X1 \mem_reg[150][2]  ( .D(n5426), .CK(clk), .Q(\mem[150][2] ) );
  DFF_X1 \mem_reg[150][1]  ( .D(n5427), .CK(clk), .Q(\mem[150][1] ) );
  DFF_X1 \mem_reg[150][0]  ( .D(n5428), .CK(clk), .Q(\mem[150][0] ) );
  DFF_X1 \mem_reg[149][7]  ( .D(n5429), .CK(clk), .Q(\mem[149][7] ) );
  DFF_X1 \mem_reg[149][6]  ( .D(n5430), .CK(clk), .Q(\mem[149][6] ) );
  DFF_X1 \mem_reg[149][5]  ( .D(n5431), .CK(clk), .Q(\mem[149][5] ) );
  DFF_X1 \mem_reg[149][4]  ( .D(n5432), .CK(clk), .Q(\mem[149][4] ) );
  DFF_X1 \mem_reg[149][3]  ( .D(n5433), .CK(clk), .Q(\mem[149][3] ) );
  DFF_X1 \mem_reg[149][2]  ( .D(n5434), .CK(clk), .Q(\mem[149][2] ) );
  DFF_X1 \mem_reg[149][1]  ( .D(n5435), .CK(clk), .Q(\mem[149][1] ) );
  DFF_X1 \mem_reg[149][0]  ( .D(n5436), .CK(clk), .Q(\mem[149][0] ) );
  DFF_X1 \mem_reg[148][7]  ( .D(n5437), .CK(clk), .Q(\mem[148][7] ) );
  DFF_X1 \mem_reg[148][6]  ( .D(n5438), .CK(clk), .Q(\mem[148][6] ) );
  DFF_X1 \mem_reg[148][5]  ( .D(n5439), .CK(clk), .Q(\mem[148][5] ) );
  DFF_X1 \mem_reg[148][4]  ( .D(n5440), .CK(clk), .Q(\mem[148][4] ) );
  DFF_X1 \mem_reg[148][3]  ( .D(n5441), .CK(clk), .Q(\mem[148][3] ) );
  DFF_X1 \mem_reg[148][2]  ( .D(n5442), .CK(clk), .Q(\mem[148][2] ) );
  DFF_X1 \mem_reg[148][1]  ( .D(n5443), .CK(clk), .Q(\mem[148][1] ) );
  DFF_X1 \mem_reg[148][0]  ( .D(n5444), .CK(clk), .Q(\mem[148][0] ) );
  DFF_X1 \mem_reg[147][7]  ( .D(n5445), .CK(clk), .Q(\mem[147][7] ) );
  DFF_X1 \mem_reg[147][6]  ( .D(n5446), .CK(clk), .Q(\mem[147][6] ) );
  DFF_X1 \mem_reg[147][5]  ( .D(n5447), .CK(clk), .Q(\mem[147][5] ) );
  DFF_X1 \mem_reg[147][4]  ( .D(n5448), .CK(clk), .Q(\mem[147][4] ) );
  DFF_X1 \mem_reg[147][3]  ( .D(n5449), .CK(clk), .Q(\mem[147][3] ) );
  DFF_X1 \mem_reg[147][2]  ( .D(n5450), .CK(clk), .Q(\mem[147][2] ) );
  DFF_X1 \mem_reg[147][1]  ( .D(n5451), .CK(clk), .Q(\mem[147][1] ) );
  DFF_X1 \mem_reg[147][0]  ( .D(n5452), .CK(clk), .Q(\mem[147][0] ) );
  DFF_X1 \mem_reg[146][7]  ( .D(n5453), .CK(clk), .Q(\mem[146][7] ) );
  DFF_X1 \mem_reg[146][6]  ( .D(n5454), .CK(clk), .Q(\mem[146][6] ) );
  DFF_X1 \mem_reg[146][5]  ( .D(n5455), .CK(clk), .Q(\mem[146][5] ) );
  DFF_X1 \mem_reg[146][4]  ( .D(n5456), .CK(clk), .Q(\mem[146][4] ) );
  DFF_X1 \mem_reg[146][3]  ( .D(n5457), .CK(clk), .Q(\mem[146][3] ) );
  DFF_X1 \mem_reg[146][2]  ( .D(n5458), .CK(clk), .Q(\mem[146][2] ) );
  DFF_X1 \mem_reg[146][1]  ( .D(n5459), .CK(clk), .Q(\mem[146][1] ) );
  DFF_X1 \mem_reg[146][0]  ( .D(n5460), .CK(clk), .Q(\mem[146][0] ) );
  DFF_X1 \mem_reg[145][7]  ( .D(n5461), .CK(clk), .Q(\mem[145][7] ) );
  DFF_X1 \mem_reg[145][6]  ( .D(n5462), .CK(clk), .Q(\mem[145][6] ) );
  DFF_X1 \mem_reg[145][5]  ( .D(n5463), .CK(clk), .Q(\mem[145][5] ) );
  DFF_X1 \mem_reg[145][4]  ( .D(n5464), .CK(clk), .Q(\mem[145][4] ) );
  DFF_X1 \mem_reg[145][3]  ( .D(n5465), .CK(clk), .Q(\mem[145][3] ) );
  DFF_X1 \mem_reg[145][2]  ( .D(n5466), .CK(clk), .Q(\mem[145][2] ) );
  DFF_X1 \mem_reg[145][1]  ( .D(n5467), .CK(clk), .Q(\mem[145][1] ) );
  DFF_X1 \mem_reg[145][0]  ( .D(n5468), .CK(clk), .Q(\mem[145][0] ) );
  DFF_X1 \mem_reg[144][7]  ( .D(n5469), .CK(clk), .Q(\mem[144][7] ) );
  DFF_X1 \mem_reg[144][6]  ( .D(n5470), .CK(clk), .Q(\mem[144][6] ) );
  DFF_X1 \mem_reg[144][5]  ( .D(n5471), .CK(clk), .Q(\mem[144][5] ) );
  DFF_X1 \mem_reg[144][4]  ( .D(n5472), .CK(clk), .Q(\mem[144][4] ) );
  DFF_X1 \mem_reg[144][3]  ( .D(n5473), .CK(clk), .Q(\mem[144][3] ) );
  DFF_X1 \mem_reg[144][2]  ( .D(n5474), .CK(clk), .Q(\mem[144][2] ) );
  DFF_X1 \mem_reg[144][1]  ( .D(n5475), .CK(clk), .Q(\mem[144][1] ) );
  DFF_X1 \mem_reg[144][0]  ( .D(n5476), .CK(clk), .Q(\mem[144][0] ) );
  DFF_X1 \mem_reg[143][7]  ( .D(n5477), .CK(clk), .Q(\mem[143][7] ) );
  DFF_X1 \mem_reg[143][6]  ( .D(n5478), .CK(clk), .Q(\mem[143][6] ) );
  DFF_X1 \mem_reg[143][5]  ( .D(n5479), .CK(clk), .Q(\mem[143][5] ) );
  DFF_X1 \mem_reg[143][4]  ( .D(n5480), .CK(clk), .Q(\mem[143][4] ) );
  DFF_X1 \mem_reg[143][3]  ( .D(n5481), .CK(clk), .Q(\mem[143][3] ) );
  DFF_X1 \mem_reg[143][2]  ( .D(n5482), .CK(clk), .Q(\mem[143][2] ) );
  DFF_X1 \mem_reg[143][1]  ( .D(n5483), .CK(clk), .Q(\mem[143][1] ) );
  DFF_X1 \mem_reg[143][0]  ( .D(n5484), .CK(clk), .Q(\mem[143][0] ) );
  DFF_X1 \mem_reg[142][7]  ( .D(n5485), .CK(clk), .Q(\mem[142][7] ) );
  DFF_X1 \mem_reg[142][6]  ( .D(n5486), .CK(clk), .Q(\mem[142][6] ) );
  DFF_X1 \mem_reg[142][5]  ( .D(n5487), .CK(clk), .Q(\mem[142][5] ) );
  DFF_X1 \mem_reg[142][4]  ( .D(n5488), .CK(clk), .Q(\mem[142][4] ) );
  DFF_X1 \mem_reg[142][3]  ( .D(n5489), .CK(clk), .Q(\mem[142][3] ) );
  DFF_X1 \mem_reg[142][2]  ( .D(n5490), .CK(clk), .Q(\mem[142][2] ) );
  DFF_X1 \mem_reg[142][1]  ( .D(n5491), .CK(clk), .Q(\mem[142][1] ) );
  DFF_X1 \mem_reg[142][0]  ( .D(n5492), .CK(clk), .Q(\mem[142][0] ) );
  DFF_X1 \mem_reg[141][7]  ( .D(n5493), .CK(clk), .Q(\mem[141][7] ) );
  DFF_X1 \mem_reg[141][6]  ( .D(n5494), .CK(clk), .Q(\mem[141][6] ) );
  DFF_X1 \mem_reg[141][5]  ( .D(n5495), .CK(clk), .Q(\mem[141][5] ) );
  DFF_X1 \mem_reg[141][4]  ( .D(n5496), .CK(clk), .Q(\mem[141][4] ) );
  DFF_X1 \mem_reg[141][3]  ( .D(n5497), .CK(clk), .Q(\mem[141][3] ) );
  DFF_X1 \mem_reg[141][2]  ( .D(n5498), .CK(clk), .Q(\mem[141][2] ) );
  DFF_X1 \mem_reg[141][1]  ( .D(n5499), .CK(clk), .Q(\mem[141][1] ) );
  DFF_X1 \mem_reg[141][0]  ( .D(n5500), .CK(clk), .Q(\mem[141][0] ) );
  DFF_X1 \mem_reg[140][7]  ( .D(n5501), .CK(clk), .Q(\mem[140][7] ) );
  DFF_X1 \mem_reg[140][6]  ( .D(n5502), .CK(clk), .Q(\mem[140][6] ) );
  DFF_X1 \mem_reg[140][5]  ( .D(n5503), .CK(clk), .Q(\mem[140][5] ) );
  DFF_X1 \mem_reg[140][4]  ( .D(n5504), .CK(clk), .Q(\mem[140][4] ) );
  DFF_X1 \mem_reg[140][3]  ( .D(n5505), .CK(clk), .Q(\mem[140][3] ) );
  DFF_X1 \mem_reg[140][2]  ( .D(n5506), .CK(clk), .Q(\mem[140][2] ) );
  DFF_X1 \mem_reg[140][1]  ( .D(n5507), .CK(clk), .Q(\mem[140][1] ) );
  DFF_X1 \mem_reg[140][0]  ( .D(n5508), .CK(clk), .Q(\mem[140][0] ) );
  DFF_X1 \mem_reg[139][7]  ( .D(n5509), .CK(clk), .Q(\mem[139][7] ) );
  DFF_X1 \mem_reg[139][6]  ( .D(n5510), .CK(clk), .Q(\mem[139][6] ) );
  DFF_X1 \mem_reg[139][5]  ( .D(n5511), .CK(clk), .Q(\mem[139][5] ) );
  DFF_X1 \mem_reg[139][4]  ( .D(n5512), .CK(clk), .Q(\mem[139][4] ) );
  DFF_X1 \mem_reg[139][3]  ( .D(n5513), .CK(clk), .Q(\mem[139][3] ) );
  DFF_X1 \mem_reg[139][2]  ( .D(n5514), .CK(clk), .Q(\mem[139][2] ) );
  DFF_X1 \mem_reg[139][1]  ( .D(n5515), .CK(clk), .Q(\mem[139][1] ) );
  DFF_X1 \mem_reg[139][0]  ( .D(n5516), .CK(clk), .Q(\mem[139][0] ) );
  DFF_X1 \mem_reg[138][7]  ( .D(n5517), .CK(clk), .Q(\mem[138][7] ) );
  DFF_X1 \mem_reg[138][6]  ( .D(n5518), .CK(clk), .Q(\mem[138][6] ) );
  DFF_X1 \mem_reg[138][5]  ( .D(n5519), .CK(clk), .Q(\mem[138][5] ) );
  DFF_X1 \mem_reg[138][4]  ( .D(n5520), .CK(clk), .Q(\mem[138][4] ) );
  DFF_X1 \mem_reg[138][3]  ( .D(n5521), .CK(clk), .Q(\mem[138][3] ) );
  DFF_X1 \mem_reg[138][2]  ( .D(n5522), .CK(clk), .Q(\mem[138][2] ) );
  DFF_X1 \mem_reg[138][1]  ( .D(n5523), .CK(clk), .Q(\mem[138][1] ) );
  DFF_X1 \mem_reg[138][0]  ( .D(n5524), .CK(clk), .Q(\mem[138][0] ) );
  DFF_X1 \mem_reg[137][7]  ( .D(n5525), .CK(clk), .Q(\mem[137][7] ) );
  DFF_X1 \mem_reg[137][6]  ( .D(n5526), .CK(clk), .Q(\mem[137][6] ) );
  DFF_X1 \mem_reg[137][5]  ( .D(n5527), .CK(clk), .Q(\mem[137][5] ) );
  DFF_X1 \mem_reg[137][4]  ( .D(n5528), .CK(clk), .Q(\mem[137][4] ) );
  DFF_X1 \mem_reg[137][3]  ( .D(n5529), .CK(clk), .Q(\mem[137][3] ) );
  DFF_X1 \mem_reg[137][2]  ( .D(n5530), .CK(clk), .Q(\mem[137][2] ) );
  DFF_X1 \mem_reg[137][1]  ( .D(n5531), .CK(clk), .Q(\mem[137][1] ) );
  DFF_X1 \mem_reg[137][0]  ( .D(n5532), .CK(clk), .Q(\mem[137][0] ) );
  DFF_X1 \mem_reg[136][7]  ( .D(n5533), .CK(clk), .Q(\mem[136][7] ) );
  DFF_X1 \mem_reg[136][6]  ( .D(n5534), .CK(clk), .Q(\mem[136][6] ) );
  DFF_X1 \mem_reg[136][5]  ( .D(n5535), .CK(clk), .Q(\mem[136][5] ) );
  DFF_X1 \mem_reg[136][4]  ( .D(n5536), .CK(clk), .Q(\mem[136][4] ) );
  DFF_X1 \mem_reg[136][3]  ( .D(n5537), .CK(clk), .Q(\mem[136][3] ) );
  DFF_X1 \mem_reg[136][2]  ( .D(n5538), .CK(clk), .Q(\mem[136][2] ) );
  DFF_X1 \mem_reg[136][1]  ( .D(n5539), .CK(clk), .Q(\mem[136][1] ) );
  DFF_X1 \mem_reg[136][0]  ( .D(n5540), .CK(clk), .Q(\mem[136][0] ) );
  DFF_X1 \mem_reg[135][7]  ( .D(n5541), .CK(clk), .Q(\mem[135][7] ) );
  DFF_X1 \mem_reg[135][6]  ( .D(n5542), .CK(clk), .Q(\mem[135][6] ) );
  DFF_X1 \mem_reg[135][5]  ( .D(n5543), .CK(clk), .Q(\mem[135][5] ) );
  DFF_X1 \mem_reg[135][4]  ( .D(n5544), .CK(clk), .Q(\mem[135][4] ) );
  DFF_X1 \mem_reg[135][3]  ( .D(n5545), .CK(clk), .Q(\mem[135][3] ) );
  DFF_X1 \mem_reg[135][2]  ( .D(n5546), .CK(clk), .Q(\mem[135][2] ) );
  DFF_X1 \mem_reg[135][1]  ( .D(n5547), .CK(clk), .Q(\mem[135][1] ) );
  DFF_X1 \mem_reg[135][0]  ( .D(n5548), .CK(clk), .Q(\mem[135][0] ) );
  DFF_X1 \mem_reg[134][7]  ( .D(n5549), .CK(clk), .Q(\mem[134][7] ) );
  DFF_X1 \mem_reg[134][6]  ( .D(n5550), .CK(clk), .Q(\mem[134][6] ) );
  DFF_X1 \mem_reg[134][5]  ( .D(n5551), .CK(clk), .Q(\mem[134][5] ) );
  DFF_X1 \mem_reg[134][4]  ( .D(n5552), .CK(clk), .Q(\mem[134][4] ) );
  DFF_X1 \mem_reg[134][3]  ( .D(n5553), .CK(clk), .Q(\mem[134][3] ) );
  DFF_X1 \mem_reg[134][2]  ( .D(n5554), .CK(clk), .Q(\mem[134][2] ) );
  DFF_X1 \mem_reg[134][1]  ( .D(n5555), .CK(clk), .Q(\mem[134][1] ) );
  DFF_X1 \mem_reg[134][0]  ( .D(n5556), .CK(clk), .Q(\mem[134][0] ) );
  DFF_X1 \mem_reg[133][7]  ( .D(n5557), .CK(clk), .Q(\mem[133][7] ) );
  DFF_X1 \mem_reg[133][6]  ( .D(n5558), .CK(clk), .Q(\mem[133][6] ) );
  DFF_X1 \mem_reg[133][5]  ( .D(n5559), .CK(clk), .Q(\mem[133][5] ) );
  DFF_X1 \mem_reg[133][4]  ( .D(n5560), .CK(clk), .Q(\mem[133][4] ) );
  DFF_X1 \mem_reg[133][3]  ( .D(n5561), .CK(clk), .Q(\mem[133][3] ) );
  DFF_X1 \mem_reg[133][2]  ( .D(n5562), .CK(clk), .Q(\mem[133][2] ) );
  DFF_X1 \mem_reg[133][1]  ( .D(n5563), .CK(clk), .Q(\mem[133][1] ) );
  DFF_X1 \mem_reg[133][0]  ( .D(n5564), .CK(clk), .Q(\mem[133][0] ) );
  DFF_X1 \mem_reg[132][7]  ( .D(n5565), .CK(clk), .Q(\mem[132][7] ) );
  DFF_X1 \mem_reg[132][6]  ( .D(n5566), .CK(clk), .Q(\mem[132][6] ) );
  DFF_X1 \mem_reg[132][5]  ( .D(n5567), .CK(clk), .Q(\mem[132][5] ) );
  DFF_X1 \mem_reg[132][4]  ( .D(n5568), .CK(clk), .Q(\mem[132][4] ) );
  DFF_X1 \mem_reg[132][3]  ( .D(n5569), .CK(clk), .Q(\mem[132][3] ) );
  DFF_X1 \mem_reg[132][2]  ( .D(n5570), .CK(clk), .Q(\mem[132][2] ) );
  DFF_X1 \mem_reg[132][1]  ( .D(n5571), .CK(clk), .Q(\mem[132][1] ) );
  DFF_X1 \mem_reg[132][0]  ( .D(n5572), .CK(clk), .Q(\mem[132][0] ) );
  DFF_X1 \mem_reg[131][7]  ( .D(n5573), .CK(clk), .Q(\mem[131][7] ) );
  DFF_X1 \mem_reg[131][6]  ( .D(n5574), .CK(clk), .Q(\mem[131][6] ) );
  DFF_X1 \mem_reg[131][5]  ( .D(n5575), .CK(clk), .Q(\mem[131][5] ) );
  DFF_X1 \mem_reg[131][4]  ( .D(n5576), .CK(clk), .Q(\mem[131][4] ) );
  DFF_X1 \mem_reg[131][3]  ( .D(n5577), .CK(clk), .Q(\mem[131][3] ) );
  DFF_X1 \mem_reg[131][2]  ( .D(n5578), .CK(clk), .Q(\mem[131][2] ) );
  DFF_X1 \mem_reg[131][1]  ( .D(n5579), .CK(clk), .Q(\mem[131][1] ) );
  DFF_X1 \mem_reg[131][0]  ( .D(n5580), .CK(clk), .Q(\mem[131][0] ) );
  DFF_X1 \mem_reg[130][7]  ( .D(n5581), .CK(clk), .Q(\mem[130][7] ) );
  DFF_X1 \mem_reg[130][6]  ( .D(n5582), .CK(clk), .Q(\mem[130][6] ) );
  DFF_X1 \mem_reg[130][5]  ( .D(n5583), .CK(clk), .Q(\mem[130][5] ) );
  DFF_X1 \mem_reg[130][4]  ( .D(n5584), .CK(clk), .Q(\mem[130][4] ) );
  DFF_X1 \mem_reg[130][3]  ( .D(n5585), .CK(clk), .Q(\mem[130][3] ) );
  DFF_X1 \mem_reg[130][2]  ( .D(n5586), .CK(clk), .Q(\mem[130][2] ) );
  DFF_X1 \mem_reg[130][1]  ( .D(n5587), .CK(clk), .Q(\mem[130][1] ) );
  DFF_X1 \mem_reg[130][0]  ( .D(n5588), .CK(clk), .Q(\mem[130][0] ) );
  DFF_X1 \mem_reg[129][7]  ( .D(n5589), .CK(clk), .Q(\mem[129][7] ) );
  DFF_X1 \mem_reg[129][6]  ( .D(n5590), .CK(clk), .Q(\mem[129][6] ) );
  DFF_X1 \mem_reg[129][5]  ( .D(n5591), .CK(clk), .Q(\mem[129][5] ) );
  DFF_X1 \mem_reg[129][4]  ( .D(n5592), .CK(clk), .Q(\mem[129][4] ) );
  DFF_X1 \mem_reg[129][3]  ( .D(n5593), .CK(clk), .Q(\mem[129][3] ) );
  DFF_X1 \mem_reg[129][2]  ( .D(n5594), .CK(clk), .Q(\mem[129][2] ) );
  DFF_X1 \mem_reg[129][1]  ( .D(n5595), .CK(clk), .Q(\mem[129][1] ) );
  DFF_X1 \mem_reg[129][0]  ( .D(n5596), .CK(clk), .Q(\mem[129][0] ) );
  DFF_X1 \mem_reg[128][7]  ( .D(n5597), .CK(clk), .Q(\mem[128][7] ) );
  DFF_X1 \mem_reg[128][6]  ( .D(n5598), .CK(clk), .Q(\mem[128][6] ) );
  DFF_X1 \mem_reg[128][5]  ( .D(n5599), .CK(clk), .Q(\mem[128][5] ) );
  DFF_X1 \mem_reg[128][4]  ( .D(n5600), .CK(clk), .Q(\mem[128][4] ) );
  DFF_X1 \mem_reg[128][3]  ( .D(n5601), .CK(clk), .Q(\mem[128][3] ) );
  DFF_X1 \mem_reg[128][2]  ( .D(n5602), .CK(clk), .Q(\mem[128][2] ) );
  DFF_X1 \mem_reg[128][1]  ( .D(n5603), .CK(clk), .Q(\mem[128][1] ) );
  DFF_X1 \mem_reg[128][0]  ( .D(n5604), .CK(clk), .Q(\mem[128][0] ) );
  DFF_X1 \mem_reg[127][7]  ( .D(n5605), .CK(clk), .Q(\mem[127][7] ) );
  DFF_X1 \mem_reg[127][6]  ( .D(n5606), .CK(clk), .Q(\mem[127][6] ) );
  DFF_X1 \mem_reg[127][5]  ( .D(n5607), .CK(clk), .Q(\mem[127][5] ) );
  DFF_X1 \mem_reg[127][4]  ( .D(n5608), .CK(clk), .Q(\mem[127][4] ) );
  DFF_X1 \mem_reg[127][3]  ( .D(n5609), .CK(clk), .Q(\mem[127][3] ) );
  DFF_X1 \mem_reg[127][2]  ( .D(n5610), .CK(clk), .Q(\mem[127][2] ) );
  DFF_X1 \mem_reg[127][1]  ( .D(n5611), .CK(clk), .Q(\mem[127][1] ) );
  DFF_X1 \mem_reg[127][0]  ( .D(n5612), .CK(clk), .Q(\mem[127][0] ) );
  DFF_X1 \mem_reg[126][7]  ( .D(n5613), .CK(clk), .Q(\mem[126][7] ) );
  DFF_X1 \mem_reg[126][6]  ( .D(n5614), .CK(clk), .Q(\mem[126][6] ) );
  DFF_X1 \mem_reg[126][5]  ( .D(n5615), .CK(clk), .Q(\mem[126][5] ) );
  DFF_X1 \mem_reg[126][4]  ( .D(n5616), .CK(clk), .Q(\mem[126][4] ) );
  DFF_X1 \mem_reg[126][3]  ( .D(n5617), .CK(clk), .Q(\mem[126][3] ) );
  DFF_X1 \mem_reg[126][2]  ( .D(n5618), .CK(clk), .Q(\mem[126][2] ) );
  DFF_X1 \mem_reg[126][1]  ( .D(n5619), .CK(clk), .Q(\mem[126][1] ) );
  DFF_X1 \mem_reg[126][0]  ( .D(n5620), .CK(clk), .Q(\mem[126][0] ) );
  DFF_X1 \mem_reg[125][7]  ( .D(n5621), .CK(clk), .Q(\mem[125][7] ) );
  DFF_X1 \mem_reg[125][6]  ( .D(n5622), .CK(clk), .Q(\mem[125][6] ) );
  DFF_X1 \mem_reg[125][5]  ( .D(n5623), .CK(clk), .Q(\mem[125][5] ) );
  DFF_X1 \mem_reg[125][4]  ( .D(n5624), .CK(clk), .Q(\mem[125][4] ) );
  DFF_X1 \mem_reg[125][3]  ( .D(n5625), .CK(clk), .Q(\mem[125][3] ) );
  DFF_X1 \mem_reg[125][2]  ( .D(n5626), .CK(clk), .Q(\mem[125][2] ) );
  DFF_X1 \mem_reg[125][1]  ( .D(n5627), .CK(clk), .Q(\mem[125][1] ) );
  DFF_X1 \mem_reg[125][0]  ( .D(n5628), .CK(clk), .Q(\mem[125][0] ) );
  DFF_X1 \mem_reg[124][7]  ( .D(n5629), .CK(clk), .Q(\mem[124][7] ) );
  DFF_X1 \mem_reg[124][6]  ( .D(n5630), .CK(clk), .Q(\mem[124][6] ) );
  DFF_X1 \mem_reg[124][5]  ( .D(n5631), .CK(clk), .Q(\mem[124][5] ) );
  DFF_X1 \mem_reg[124][4]  ( .D(n5632), .CK(clk), .Q(\mem[124][4] ) );
  DFF_X1 \mem_reg[124][3]  ( .D(n5633), .CK(clk), .Q(\mem[124][3] ) );
  DFF_X1 \mem_reg[124][2]  ( .D(n5634), .CK(clk), .Q(\mem[124][2] ) );
  DFF_X1 \mem_reg[124][1]  ( .D(n5635), .CK(clk), .Q(\mem[124][1] ) );
  DFF_X1 \mem_reg[124][0]  ( .D(n5636), .CK(clk), .Q(\mem[124][0] ) );
  DFF_X1 \mem_reg[123][7]  ( .D(n5637), .CK(clk), .Q(\mem[123][7] ) );
  DFF_X1 \mem_reg[123][6]  ( .D(n5638), .CK(clk), .Q(\mem[123][6] ) );
  DFF_X1 \mem_reg[123][5]  ( .D(n5639), .CK(clk), .Q(\mem[123][5] ) );
  DFF_X1 \mem_reg[123][4]  ( .D(n5640), .CK(clk), .Q(\mem[123][4] ) );
  DFF_X1 \mem_reg[123][3]  ( .D(n5641), .CK(clk), .Q(\mem[123][3] ) );
  DFF_X1 \mem_reg[123][2]  ( .D(n5642), .CK(clk), .Q(\mem[123][2] ) );
  DFF_X1 \mem_reg[123][1]  ( .D(n5643), .CK(clk), .Q(\mem[123][1] ) );
  DFF_X1 \mem_reg[123][0]  ( .D(n5644), .CK(clk), .Q(\mem[123][0] ) );
  DFF_X1 \mem_reg[122][7]  ( .D(n5645), .CK(clk), .Q(\mem[122][7] ) );
  DFF_X1 \mem_reg[122][6]  ( .D(n5646), .CK(clk), .Q(\mem[122][6] ) );
  DFF_X1 \mem_reg[122][5]  ( .D(n5647), .CK(clk), .Q(\mem[122][5] ) );
  DFF_X1 \mem_reg[122][4]  ( .D(n5648), .CK(clk), .Q(\mem[122][4] ) );
  DFF_X1 \mem_reg[122][3]  ( .D(n5649), .CK(clk), .Q(\mem[122][3] ) );
  DFF_X1 \mem_reg[122][2]  ( .D(n5650), .CK(clk), .Q(\mem[122][2] ) );
  DFF_X1 \mem_reg[122][1]  ( .D(n5651), .CK(clk), .Q(\mem[122][1] ) );
  DFF_X1 \mem_reg[122][0]  ( .D(n5652), .CK(clk), .Q(\mem[122][0] ) );
  DFF_X1 \mem_reg[121][7]  ( .D(n5653), .CK(clk), .Q(\mem[121][7] ) );
  DFF_X1 \mem_reg[121][6]  ( .D(n5654), .CK(clk), .Q(\mem[121][6] ) );
  DFF_X1 \mem_reg[121][5]  ( .D(n5655), .CK(clk), .Q(\mem[121][5] ) );
  DFF_X1 \mem_reg[121][4]  ( .D(n5656), .CK(clk), .Q(\mem[121][4] ) );
  DFF_X1 \mem_reg[121][3]  ( .D(n5657), .CK(clk), .Q(\mem[121][3] ) );
  DFF_X1 \mem_reg[121][2]  ( .D(n5658), .CK(clk), .Q(\mem[121][2] ) );
  DFF_X1 \mem_reg[121][1]  ( .D(n5659), .CK(clk), .Q(\mem[121][1] ) );
  DFF_X1 \mem_reg[121][0]  ( .D(n5660), .CK(clk), .Q(\mem[121][0] ) );
  DFF_X1 \mem_reg[120][7]  ( .D(n5661), .CK(clk), .Q(\mem[120][7] ) );
  DFF_X1 \mem_reg[120][6]  ( .D(n5662), .CK(clk), .Q(\mem[120][6] ) );
  DFF_X1 \mem_reg[120][5]  ( .D(n5663), .CK(clk), .Q(\mem[120][5] ) );
  DFF_X1 \mem_reg[120][4]  ( .D(n5664), .CK(clk), .Q(\mem[120][4] ) );
  DFF_X1 \mem_reg[120][3]  ( .D(n5665), .CK(clk), .Q(\mem[120][3] ) );
  DFF_X1 \mem_reg[120][2]  ( .D(n5666), .CK(clk), .Q(\mem[120][2] ) );
  DFF_X1 \mem_reg[120][1]  ( .D(n5667), .CK(clk), .Q(\mem[120][1] ) );
  DFF_X1 \mem_reg[120][0]  ( .D(n5668), .CK(clk), .Q(\mem[120][0] ) );
  DFF_X1 \mem_reg[119][7]  ( .D(n5669), .CK(clk), .Q(\mem[119][7] ) );
  DFF_X1 \mem_reg[119][6]  ( .D(n5670), .CK(clk), .Q(\mem[119][6] ) );
  DFF_X1 \mem_reg[119][5]  ( .D(n5671), .CK(clk), .Q(\mem[119][5] ) );
  DFF_X1 \mem_reg[119][4]  ( .D(n5672), .CK(clk), .Q(\mem[119][4] ) );
  DFF_X1 \mem_reg[119][3]  ( .D(n5673), .CK(clk), .Q(\mem[119][3] ) );
  DFF_X1 \mem_reg[119][2]  ( .D(n5674), .CK(clk), .Q(\mem[119][2] ) );
  DFF_X1 \mem_reg[119][1]  ( .D(n5675), .CK(clk), .Q(\mem[119][1] ) );
  DFF_X1 \mem_reg[119][0]  ( .D(n5676), .CK(clk), .Q(\mem[119][0] ) );
  DFF_X1 \mem_reg[118][7]  ( .D(n5677), .CK(clk), .Q(\mem[118][7] ) );
  DFF_X1 \mem_reg[118][6]  ( .D(n5678), .CK(clk), .Q(\mem[118][6] ) );
  DFF_X1 \mem_reg[118][5]  ( .D(n5679), .CK(clk), .Q(\mem[118][5] ) );
  DFF_X1 \mem_reg[118][4]  ( .D(n5680), .CK(clk), .Q(\mem[118][4] ) );
  DFF_X1 \mem_reg[118][3]  ( .D(n5681), .CK(clk), .Q(\mem[118][3] ) );
  DFF_X1 \mem_reg[118][2]  ( .D(n5682), .CK(clk), .Q(\mem[118][2] ) );
  DFF_X1 \mem_reg[118][1]  ( .D(n5683), .CK(clk), .Q(\mem[118][1] ) );
  DFF_X1 \mem_reg[118][0]  ( .D(n5684), .CK(clk), .Q(\mem[118][0] ) );
  DFF_X1 \mem_reg[117][7]  ( .D(n5685), .CK(clk), .Q(\mem[117][7] ) );
  DFF_X1 \mem_reg[117][6]  ( .D(n5686), .CK(clk), .Q(\mem[117][6] ) );
  DFF_X1 \mem_reg[117][5]  ( .D(n5687), .CK(clk), .Q(\mem[117][5] ) );
  DFF_X1 \mem_reg[117][4]  ( .D(n5688), .CK(clk), .Q(\mem[117][4] ) );
  DFF_X1 \mem_reg[117][3]  ( .D(n5689), .CK(clk), .Q(\mem[117][3] ) );
  DFF_X1 \mem_reg[117][2]  ( .D(n5690), .CK(clk), .Q(\mem[117][2] ) );
  DFF_X1 \mem_reg[117][1]  ( .D(n5691), .CK(clk), .Q(\mem[117][1] ) );
  DFF_X1 \mem_reg[117][0]  ( .D(n5692), .CK(clk), .Q(\mem[117][0] ) );
  DFF_X1 \mem_reg[116][7]  ( .D(n5693), .CK(clk), .Q(\mem[116][7] ) );
  DFF_X1 \mem_reg[116][6]  ( .D(n5694), .CK(clk), .Q(\mem[116][6] ) );
  DFF_X1 \mem_reg[116][5]  ( .D(n5695), .CK(clk), .Q(\mem[116][5] ) );
  DFF_X1 \mem_reg[116][4]  ( .D(n5696), .CK(clk), .Q(\mem[116][4] ) );
  DFF_X1 \mem_reg[116][3]  ( .D(n5697), .CK(clk), .Q(\mem[116][3] ) );
  DFF_X1 \mem_reg[116][2]  ( .D(n5698), .CK(clk), .Q(\mem[116][2] ) );
  DFF_X1 \mem_reg[116][1]  ( .D(n5699), .CK(clk), .Q(\mem[116][1] ) );
  DFF_X1 \mem_reg[116][0]  ( .D(n5700), .CK(clk), .Q(\mem[116][0] ) );
  DFF_X1 \mem_reg[115][7]  ( .D(n5701), .CK(clk), .Q(\mem[115][7] ) );
  DFF_X1 \mem_reg[115][6]  ( .D(n5702), .CK(clk), .Q(\mem[115][6] ) );
  DFF_X1 \mem_reg[115][5]  ( .D(n5703), .CK(clk), .Q(\mem[115][5] ) );
  DFF_X1 \mem_reg[115][4]  ( .D(n5704), .CK(clk), .Q(\mem[115][4] ) );
  DFF_X1 \mem_reg[115][3]  ( .D(n5705), .CK(clk), .Q(\mem[115][3] ) );
  DFF_X1 \mem_reg[115][2]  ( .D(n5706), .CK(clk), .Q(\mem[115][2] ) );
  DFF_X1 \mem_reg[115][1]  ( .D(n5707), .CK(clk), .Q(\mem[115][1] ) );
  DFF_X1 \mem_reg[115][0]  ( .D(n5708), .CK(clk), .Q(\mem[115][0] ) );
  DFF_X1 \mem_reg[114][7]  ( .D(n5709), .CK(clk), .Q(\mem[114][7] ) );
  DFF_X1 \mem_reg[114][6]  ( .D(n5710), .CK(clk), .Q(\mem[114][6] ) );
  DFF_X1 \mem_reg[114][5]  ( .D(n5711), .CK(clk), .Q(\mem[114][5] ) );
  DFF_X1 \mem_reg[114][4]  ( .D(n5712), .CK(clk), .Q(\mem[114][4] ) );
  DFF_X1 \mem_reg[114][3]  ( .D(n5713), .CK(clk), .Q(\mem[114][3] ) );
  DFF_X1 \mem_reg[114][2]  ( .D(n5714), .CK(clk), .Q(\mem[114][2] ) );
  DFF_X1 \mem_reg[114][1]  ( .D(n5715), .CK(clk), .Q(\mem[114][1] ) );
  DFF_X1 \mem_reg[114][0]  ( .D(n5716), .CK(clk), .Q(\mem[114][0] ) );
  DFF_X1 \mem_reg[113][7]  ( .D(n5717), .CK(clk), .Q(\mem[113][7] ) );
  DFF_X1 \mem_reg[113][6]  ( .D(n5718), .CK(clk), .Q(\mem[113][6] ) );
  DFF_X1 \mem_reg[113][5]  ( .D(n5719), .CK(clk), .Q(\mem[113][5] ) );
  DFF_X1 \mem_reg[113][4]  ( .D(n5720), .CK(clk), .Q(\mem[113][4] ) );
  DFF_X1 \mem_reg[113][3]  ( .D(n5721), .CK(clk), .Q(\mem[113][3] ) );
  DFF_X1 \mem_reg[113][2]  ( .D(n5722), .CK(clk), .Q(\mem[113][2] ) );
  DFF_X1 \mem_reg[113][1]  ( .D(n5723), .CK(clk), .Q(\mem[113][1] ) );
  DFF_X1 \mem_reg[113][0]  ( .D(n5724), .CK(clk), .Q(\mem[113][0] ) );
  DFF_X1 \mem_reg[112][7]  ( .D(n5725), .CK(clk), .Q(\mem[112][7] ) );
  DFF_X1 \mem_reg[112][6]  ( .D(n5726), .CK(clk), .Q(\mem[112][6] ) );
  DFF_X1 \mem_reg[112][5]  ( .D(n5727), .CK(clk), .Q(\mem[112][5] ) );
  DFF_X1 \mem_reg[112][4]  ( .D(n5728), .CK(clk), .Q(\mem[112][4] ) );
  DFF_X1 \mem_reg[112][3]  ( .D(n5729), .CK(clk), .Q(\mem[112][3] ) );
  DFF_X1 \mem_reg[112][2]  ( .D(n5730), .CK(clk), .Q(\mem[112][2] ) );
  DFF_X1 \mem_reg[112][1]  ( .D(n5731), .CK(clk), .Q(\mem[112][1] ) );
  DFF_X1 \mem_reg[112][0]  ( .D(n5732), .CK(clk), .Q(\mem[112][0] ) );
  DFF_X1 \mem_reg[111][7]  ( .D(n5733), .CK(clk), .Q(\mem[111][7] ) );
  DFF_X1 \mem_reg[111][6]  ( .D(n5734), .CK(clk), .Q(\mem[111][6] ) );
  DFF_X1 \mem_reg[111][5]  ( .D(n5735), .CK(clk), .Q(\mem[111][5] ) );
  DFF_X1 \mem_reg[111][4]  ( .D(n5736), .CK(clk), .Q(\mem[111][4] ) );
  DFF_X1 \mem_reg[111][3]  ( .D(n5737), .CK(clk), .Q(\mem[111][3] ) );
  DFF_X1 \mem_reg[111][2]  ( .D(n5738), .CK(clk), .Q(\mem[111][2] ) );
  DFF_X1 \mem_reg[111][1]  ( .D(n5739), .CK(clk), .Q(\mem[111][1] ) );
  DFF_X1 \mem_reg[111][0]  ( .D(n5740), .CK(clk), .Q(\mem[111][0] ) );
  DFF_X1 \mem_reg[110][7]  ( .D(n5741), .CK(clk), .Q(\mem[110][7] ) );
  DFF_X1 \mem_reg[110][6]  ( .D(n5742), .CK(clk), .Q(\mem[110][6] ) );
  DFF_X1 \mem_reg[110][5]  ( .D(n5743), .CK(clk), .Q(\mem[110][5] ) );
  DFF_X1 \mem_reg[110][4]  ( .D(n5744), .CK(clk), .Q(\mem[110][4] ) );
  DFF_X1 \mem_reg[110][3]  ( .D(n5745), .CK(clk), .Q(\mem[110][3] ) );
  DFF_X1 \mem_reg[110][2]  ( .D(n5746), .CK(clk), .Q(\mem[110][2] ) );
  DFF_X1 \mem_reg[110][1]  ( .D(n5747), .CK(clk), .Q(\mem[110][1] ) );
  DFF_X1 \mem_reg[110][0]  ( .D(n5748), .CK(clk), .Q(\mem[110][0] ) );
  DFF_X1 \mem_reg[109][7]  ( .D(n5749), .CK(clk), .Q(\mem[109][7] ) );
  DFF_X1 \mem_reg[109][6]  ( .D(n5750), .CK(clk), .Q(\mem[109][6] ) );
  DFF_X1 \mem_reg[109][5]  ( .D(n5751), .CK(clk), .Q(\mem[109][5] ) );
  DFF_X1 \mem_reg[109][4]  ( .D(n5752), .CK(clk), .Q(\mem[109][4] ) );
  DFF_X1 \mem_reg[109][3]  ( .D(n5753), .CK(clk), .Q(\mem[109][3] ) );
  DFF_X1 \mem_reg[109][2]  ( .D(n5754), .CK(clk), .Q(\mem[109][2] ) );
  DFF_X1 \mem_reg[109][1]  ( .D(n5755), .CK(clk), .Q(\mem[109][1] ) );
  DFF_X1 \mem_reg[109][0]  ( .D(n5756), .CK(clk), .Q(\mem[109][0] ) );
  DFF_X1 \mem_reg[108][7]  ( .D(n5757), .CK(clk), .Q(\mem[108][7] ) );
  DFF_X1 \mem_reg[108][6]  ( .D(n5758), .CK(clk), .Q(\mem[108][6] ) );
  DFF_X1 \mem_reg[108][5]  ( .D(n5759), .CK(clk), .Q(\mem[108][5] ) );
  DFF_X1 \mem_reg[108][4]  ( .D(n5760), .CK(clk), .Q(\mem[108][4] ) );
  DFF_X1 \mem_reg[108][3]  ( .D(n5761), .CK(clk), .Q(\mem[108][3] ) );
  DFF_X1 \mem_reg[108][2]  ( .D(n5762), .CK(clk), .Q(\mem[108][2] ) );
  DFF_X1 \mem_reg[108][1]  ( .D(n5763), .CK(clk), .Q(\mem[108][1] ) );
  DFF_X1 \mem_reg[108][0]  ( .D(n5764), .CK(clk), .Q(\mem[108][0] ) );
  DFF_X1 \mem_reg[107][7]  ( .D(n5765), .CK(clk), .Q(\mem[107][7] ) );
  DFF_X1 \mem_reg[107][6]  ( .D(n5766), .CK(clk), .Q(\mem[107][6] ) );
  DFF_X1 \mem_reg[107][5]  ( .D(n5767), .CK(clk), .Q(\mem[107][5] ) );
  DFF_X1 \mem_reg[107][4]  ( .D(n5768), .CK(clk), .Q(\mem[107][4] ) );
  DFF_X1 \mem_reg[107][3]  ( .D(n5769), .CK(clk), .Q(\mem[107][3] ) );
  DFF_X1 \mem_reg[107][2]  ( .D(n5770), .CK(clk), .Q(\mem[107][2] ) );
  DFF_X1 \mem_reg[107][1]  ( .D(n5771), .CK(clk), .Q(\mem[107][1] ) );
  DFF_X1 \mem_reg[107][0]  ( .D(n5772), .CK(clk), .Q(\mem[107][0] ) );
  DFF_X1 \mem_reg[106][7]  ( .D(n5773), .CK(clk), .Q(\mem[106][7] ) );
  DFF_X1 \mem_reg[106][6]  ( .D(n5774), .CK(clk), .Q(\mem[106][6] ) );
  DFF_X1 \mem_reg[106][5]  ( .D(n5775), .CK(clk), .Q(\mem[106][5] ) );
  DFF_X1 \mem_reg[106][4]  ( .D(n5776), .CK(clk), .Q(\mem[106][4] ) );
  DFF_X1 \mem_reg[106][3]  ( .D(n5777), .CK(clk), .Q(\mem[106][3] ) );
  DFF_X1 \mem_reg[106][2]  ( .D(n5778), .CK(clk), .Q(\mem[106][2] ) );
  DFF_X1 \mem_reg[106][1]  ( .D(n5779), .CK(clk), .Q(\mem[106][1] ) );
  DFF_X1 \mem_reg[106][0]  ( .D(n5780), .CK(clk), .Q(\mem[106][0] ) );
  DFF_X1 \mem_reg[105][7]  ( .D(n5781), .CK(clk), .Q(\mem[105][7] ) );
  DFF_X1 \mem_reg[105][6]  ( .D(n5782), .CK(clk), .Q(\mem[105][6] ) );
  DFF_X1 \mem_reg[105][5]  ( .D(n5783), .CK(clk), .Q(\mem[105][5] ) );
  DFF_X1 \mem_reg[105][4]  ( .D(n5784), .CK(clk), .Q(\mem[105][4] ) );
  DFF_X1 \mem_reg[105][3]  ( .D(n5785), .CK(clk), .Q(\mem[105][3] ) );
  DFF_X1 \mem_reg[105][2]  ( .D(n5786), .CK(clk), .Q(\mem[105][2] ) );
  DFF_X1 \mem_reg[105][1]  ( .D(n5787), .CK(clk), .Q(\mem[105][1] ) );
  DFF_X1 \mem_reg[105][0]  ( .D(n5788), .CK(clk), .Q(\mem[105][0] ) );
  DFF_X1 \mem_reg[104][7]  ( .D(n5789), .CK(clk), .Q(\mem[104][7] ) );
  DFF_X1 \mem_reg[104][6]  ( .D(n5790), .CK(clk), .Q(\mem[104][6] ) );
  DFF_X1 \mem_reg[104][5]  ( .D(n5791), .CK(clk), .Q(\mem[104][5] ) );
  DFF_X1 \mem_reg[104][4]  ( .D(n5792), .CK(clk), .Q(\mem[104][4] ) );
  DFF_X1 \mem_reg[104][3]  ( .D(n5793), .CK(clk), .Q(\mem[104][3] ) );
  DFF_X1 \mem_reg[104][2]  ( .D(n5794), .CK(clk), .Q(\mem[104][2] ) );
  DFF_X1 \mem_reg[104][1]  ( .D(n5795), .CK(clk), .Q(\mem[104][1] ) );
  DFF_X1 \mem_reg[104][0]  ( .D(n5796), .CK(clk), .Q(\mem[104][0] ) );
  DFF_X1 \mem_reg[103][7]  ( .D(n5797), .CK(clk), .Q(\mem[103][7] ) );
  DFF_X1 \mem_reg[103][6]  ( .D(n5798), .CK(clk), .Q(\mem[103][6] ) );
  DFF_X1 \mem_reg[103][5]  ( .D(n5799), .CK(clk), .Q(\mem[103][5] ) );
  DFF_X1 \mem_reg[103][4]  ( .D(n5800), .CK(clk), .Q(\mem[103][4] ) );
  DFF_X1 \mem_reg[103][3]  ( .D(n5801), .CK(clk), .Q(\mem[103][3] ) );
  DFF_X1 \mem_reg[103][2]  ( .D(n5802), .CK(clk), .Q(\mem[103][2] ) );
  DFF_X1 \mem_reg[103][1]  ( .D(n5803), .CK(clk), .Q(\mem[103][1] ) );
  DFF_X1 \mem_reg[103][0]  ( .D(n5804), .CK(clk), .Q(\mem[103][0] ) );
  DFF_X1 \mem_reg[102][7]  ( .D(n5805), .CK(clk), .Q(\mem[102][7] ) );
  DFF_X1 \mem_reg[102][6]  ( .D(n5806), .CK(clk), .Q(\mem[102][6] ) );
  DFF_X1 \mem_reg[102][5]  ( .D(n5807), .CK(clk), .Q(\mem[102][5] ) );
  DFF_X1 \mem_reg[102][4]  ( .D(n5808), .CK(clk), .Q(\mem[102][4] ) );
  DFF_X1 \mem_reg[102][3]  ( .D(n5809), .CK(clk), .Q(\mem[102][3] ) );
  DFF_X1 \mem_reg[102][2]  ( .D(n5810), .CK(clk), .Q(\mem[102][2] ) );
  DFF_X1 \mem_reg[102][1]  ( .D(n5811), .CK(clk), .Q(\mem[102][1] ) );
  DFF_X1 \mem_reg[102][0]  ( .D(n5812), .CK(clk), .Q(\mem[102][0] ) );
  DFF_X1 \mem_reg[101][7]  ( .D(n5813), .CK(clk), .Q(\mem[101][7] ) );
  DFF_X1 \mem_reg[101][6]  ( .D(n5814), .CK(clk), .Q(\mem[101][6] ) );
  DFF_X1 \mem_reg[101][5]  ( .D(n5815), .CK(clk), .Q(\mem[101][5] ) );
  DFF_X1 \mem_reg[101][4]  ( .D(n5816), .CK(clk), .Q(\mem[101][4] ) );
  DFF_X1 \mem_reg[101][3]  ( .D(n5817), .CK(clk), .Q(\mem[101][3] ) );
  DFF_X1 \mem_reg[101][2]  ( .D(n5818), .CK(clk), .Q(\mem[101][2] ) );
  DFF_X1 \mem_reg[101][1]  ( .D(n5819), .CK(clk), .Q(\mem[101][1] ) );
  DFF_X1 \mem_reg[101][0]  ( .D(n5820), .CK(clk), .Q(\mem[101][0] ) );
  DFF_X1 \mem_reg[100][7]  ( .D(n5821), .CK(clk), .Q(\mem[100][7] ) );
  DFF_X1 \mem_reg[100][6]  ( .D(n5822), .CK(clk), .Q(\mem[100][6] ) );
  DFF_X1 \mem_reg[100][5]  ( .D(n5823), .CK(clk), .Q(\mem[100][5] ) );
  DFF_X1 \mem_reg[100][4]  ( .D(n5824), .CK(clk), .Q(\mem[100][4] ) );
  DFF_X1 \mem_reg[100][3]  ( .D(n5825), .CK(clk), .Q(\mem[100][3] ) );
  DFF_X1 \mem_reg[100][2]  ( .D(n5826), .CK(clk), .Q(\mem[100][2] ) );
  DFF_X1 \mem_reg[100][1]  ( .D(n5827), .CK(clk), .Q(\mem[100][1] ) );
  DFF_X1 \mem_reg[100][0]  ( .D(n5828), .CK(clk), .Q(\mem[100][0] ) );
  DFF_X1 \mem_reg[99][7]  ( .D(n5829), .CK(clk), .Q(\mem[99][7] ) );
  DFF_X1 \mem_reg[99][6]  ( .D(n5830), .CK(clk), .Q(\mem[99][6] ) );
  DFF_X1 \mem_reg[99][5]  ( .D(n5831), .CK(clk), .Q(\mem[99][5] ) );
  DFF_X1 \mem_reg[99][4]  ( .D(n5832), .CK(clk), .Q(\mem[99][4] ) );
  DFF_X1 \mem_reg[99][3]  ( .D(n5833), .CK(clk), .Q(\mem[99][3] ) );
  DFF_X1 \mem_reg[99][2]  ( .D(n5834), .CK(clk), .Q(\mem[99][2] ) );
  DFF_X1 \mem_reg[99][1]  ( .D(n5835), .CK(clk), .Q(\mem[99][1] ) );
  DFF_X1 \mem_reg[99][0]  ( .D(n5836), .CK(clk), .Q(\mem[99][0] ) );
  DFF_X1 \mem_reg[98][7]  ( .D(n5837), .CK(clk), .Q(\mem[98][7] ) );
  DFF_X1 \mem_reg[98][6]  ( .D(n5838), .CK(clk), .Q(\mem[98][6] ) );
  DFF_X1 \mem_reg[98][5]  ( .D(n5839), .CK(clk), .Q(\mem[98][5] ) );
  DFF_X1 \mem_reg[98][4]  ( .D(n5840), .CK(clk), .Q(\mem[98][4] ) );
  DFF_X1 \mem_reg[98][3]  ( .D(n5841), .CK(clk), .Q(\mem[98][3] ) );
  DFF_X1 \mem_reg[98][2]  ( .D(n5842), .CK(clk), .Q(\mem[98][2] ) );
  DFF_X1 \mem_reg[98][1]  ( .D(n5843), .CK(clk), .Q(\mem[98][1] ) );
  DFF_X1 \mem_reg[98][0]  ( .D(n5844), .CK(clk), .Q(\mem[98][0] ) );
  DFF_X1 \mem_reg[97][7]  ( .D(n5845), .CK(clk), .Q(\mem[97][7] ) );
  DFF_X1 \mem_reg[97][6]  ( .D(n5846), .CK(clk), .Q(\mem[97][6] ) );
  DFF_X1 \mem_reg[97][5]  ( .D(n5847), .CK(clk), .Q(\mem[97][5] ) );
  DFF_X1 \mem_reg[97][4]  ( .D(n5848), .CK(clk), .Q(\mem[97][4] ) );
  DFF_X1 \mem_reg[97][3]  ( .D(n5849), .CK(clk), .Q(\mem[97][3] ) );
  DFF_X1 \mem_reg[97][2]  ( .D(n5850), .CK(clk), .Q(\mem[97][2] ) );
  DFF_X1 \mem_reg[97][1]  ( .D(n5851), .CK(clk), .Q(\mem[97][1] ) );
  DFF_X1 \mem_reg[97][0]  ( .D(n5852), .CK(clk), .Q(\mem[97][0] ) );
  DFF_X1 \mem_reg[96][7]  ( .D(n5853), .CK(clk), .Q(\mem[96][7] ) );
  DFF_X1 \mem_reg[96][6]  ( .D(n5854), .CK(clk), .Q(\mem[96][6] ) );
  DFF_X1 \mem_reg[96][5]  ( .D(n5855), .CK(clk), .Q(\mem[96][5] ) );
  DFF_X1 \mem_reg[96][4]  ( .D(n5856), .CK(clk), .Q(\mem[96][4] ) );
  DFF_X1 \mem_reg[96][3]  ( .D(n5857), .CK(clk), .Q(\mem[96][3] ) );
  DFF_X1 \mem_reg[96][2]  ( .D(n5858), .CK(clk), .Q(\mem[96][2] ) );
  DFF_X1 \mem_reg[96][1]  ( .D(n5859), .CK(clk), .Q(\mem[96][1] ) );
  DFF_X1 \mem_reg[96][0]  ( .D(n5860), .CK(clk), .Q(\mem[96][0] ) );
  DFF_X1 \mem_reg[95][7]  ( .D(n5861), .CK(clk), .Q(\mem[95][7] ) );
  DFF_X1 \mem_reg[95][6]  ( .D(n5862), .CK(clk), .Q(\mem[95][6] ) );
  DFF_X1 \mem_reg[95][5]  ( .D(n5863), .CK(clk), .Q(\mem[95][5] ) );
  DFF_X1 \mem_reg[95][4]  ( .D(n5864), .CK(clk), .Q(\mem[95][4] ) );
  DFF_X1 \mem_reg[95][3]  ( .D(n5865), .CK(clk), .Q(\mem[95][3] ) );
  DFF_X1 \mem_reg[95][2]  ( .D(n5866), .CK(clk), .Q(\mem[95][2] ) );
  DFF_X1 \mem_reg[95][1]  ( .D(n5867), .CK(clk), .Q(\mem[95][1] ) );
  DFF_X1 \mem_reg[95][0]  ( .D(n5868), .CK(clk), .Q(\mem[95][0] ) );
  DFF_X1 \mem_reg[94][7]  ( .D(n5869), .CK(clk), .Q(\mem[94][7] ) );
  DFF_X1 \mem_reg[94][6]  ( .D(n5870), .CK(clk), .Q(\mem[94][6] ) );
  DFF_X1 \mem_reg[94][5]  ( .D(n5871), .CK(clk), .Q(\mem[94][5] ) );
  DFF_X1 \mem_reg[94][4]  ( .D(n5872), .CK(clk), .Q(\mem[94][4] ) );
  DFF_X1 \mem_reg[94][3]  ( .D(n5873), .CK(clk), .Q(\mem[94][3] ) );
  DFF_X1 \mem_reg[94][2]  ( .D(n5874), .CK(clk), .Q(\mem[94][2] ) );
  DFF_X1 \mem_reg[94][1]  ( .D(n5875), .CK(clk), .Q(\mem[94][1] ) );
  DFF_X1 \mem_reg[94][0]  ( .D(n5876), .CK(clk), .Q(\mem[94][0] ) );
  DFF_X1 \mem_reg[93][7]  ( .D(n5877), .CK(clk), .Q(\mem[93][7] ) );
  DFF_X1 \mem_reg[93][6]  ( .D(n5878), .CK(clk), .Q(\mem[93][6] ) );
  DFF_X1 \mem_reg[93][5]  ( .D(n5879), .CK(clk), .Q(\mem[93][5] ) );
  DFF_X1 \mem_reg[93][4]  ( .D(n5880), .CK(clk), .Q(\mem[93][4] ) );
  DFF_X1 \mem_reg[93][3]  ( .D(n5881), .CK(clk), .Q(\mem[93][3] ) );
  DFF_X1 \mem_reg[93][2]  ( .D(n5882), .CK(clk), .Q(\mem[93][2] ) );
  DFF_X1 \mem_reg[93][1]  ( .D(n5883), .CK(clk), .Q(\mem[93][1] ) );
  DFF_X1 \mem_reg[93][0]  ( .D(n5884), .CK(clk), .Q(\mem[93][0] ) );
  DFF_X1 \mem_reg[92][7]  ( .D(n5885), .CK(clk), .Q(\mem[92][7] ) );
  DFF_X1 \mem_reg[92][6]  ( .D(n5886), .CK(clk), .Q(\mem[92][6] ) );
  DFF_X1 \mem_reg[92][5]  ( .D(n5887), .CK(clk), .Q(\mem[92][5] ) );
  DFF_X1 \mem_reg[92][4]  ( .D(n5888), .CK(clk), .Q(\mem[92][4] ) );
  DFF_X1 \mem_reg[92][3]  ( .D(n5889), .CK(clk), .Q(\mem[92][3] ) );
  DFF_X1 \mem_reg[92][2]  ( .D(n5890), .CK(clk), .Q(\mem[92][2] ) );
  DFF_X1 \mem_reg[92][1]  ( .D(n5891), .CK(clk), .Q(\mem[92][1] ) );
  DFF_X1 \mem_reg[92][0]  ( .D(n5892), .CK(clk), .Q(\mem[92][0] ) );
  DFF_X1 \mem_reg[91][7]  ( .D(n5893), .CK(clk), .Q(\mem[91][7] ) );
  DFF_X1 \mem_reg[91][6]  ( .D(n5894), .CK(clk), .Q(\mem[91][6] ) );
  DFF_X1 \mem_reg[91][5]  ( .D(n5895), .CK(clk), .Q(\mem[91][5] ) );
  DFF_X1 \mem_reg[91][4]  ( .D(n5896), .CK(clk), .Q(\mem[91][4] ) );
  DFF_X1 \mem_reg[91][3]  ( .D(n5897), .CK(clk), .Q(\mem[91][3] ) );
  DFF_X1 \mem_reg[91][2]  ( .D(n5898), .CK(clk), .Q(\mem[91][2] ) );
  DFF_X1 \mem_reg[91][1]  ( .D(n5899), .CK(clk), .Q(\mem[91][1] ) );
  DFF_X1 \mem_reg[91][0]  ( .D(n5900), .CK(clk), .Q(\mem[91][0] ) );
  DFF_X1 \mem_reg[90][7]  ( .D(n5901), .CK(clk), .Q(\mem[90][7] ) );
  DFF_X1 \mem_reg[90][6]  ( .D(n5902), .CK(clk), .Q(\mem[90][6] ) );
  DFF_X1 \mem_reg[90][5]  ( .D(n5903), .CK(clk), .Q(\mem[90][5] ) );
  DFF_X1 \mem_reg[90][4]  ( .D(n5904), .CK(clk), .Q(\mem[90][4] ) );
  DFF_X1 \mem_reg[90][3]  ( .D(n5905), .CK(clk), .Q(\mem[90][3] ) );
  DFF_X1 \mem_reg[90][2]  ( .D(n5906), .CK(clk), .Q(\mem[90][2] ) );
  DFF_X1 \mem_reg[90][1]  ( .D(n5907), .CK(clk), .Q(\mem[90][1] ) );
  DFF_X1 \mem_reg[90][0]  ( .D(n5908), .CK(clk), .Q(\mem[90][0] ) );
  DFF_X1 \mem_reg[89][7]  ( .D(n5909), .CK(clk), .Q(\mem[89][7] ) );
  DFF_X1 \mem_reg[89][6]  ( .D(n5910), .CK(clk), .Q(\mem[89][6] ) );
  DFF_X1 \mem_reg[89][5]  ( .D(n5911), .CK(clk), .Q(\mem[89][5] ) );
  DFF_X1 \mem_reg[89][4]  ( .D(n5912), .CK(clk), .Q(\mem[89][4] ) );
  DFF_X1 \mem_reg[89][3]  ( .D(n5913), .CK(clk), .Q(\mem[89][3] ) );
  DFF_X1 \mem_reg[89][2]  ( .D(n5914), .CK(clk), .Q(\mem[89][2] ) );
  DFF_X1 \mem_reg[89][1]  ( .D(n5915), .CK(clk), .Q(\mem[89][1] ) );
  DFF_X1 \mem_reg[89][0]  ( .D(n5916), .CK(clk), .Q(\mem[89][0] ) );
  DFF_X1 \mem_reg[88][7]  ( .D(n5917), .CK(clk), .Q(\mem[88][7] ) );
  DFF_X1 \mem_reg[88][6]  ( .D(n5918), .CK(clk), .Q(\mem[88][6] ) );
  DFF_X1 \mem_reg[88][5]  ( .D(n5919), .CK(clk), .Q(\mem[88][5] ) );
  DFF_X1 \mem_reg[88][4]  ( .D(n5920), .CK(clk), .Q(\mem[88][4] ) );
  DFF_X1 \mem_reg[88][3]  ( .D(n5921), .CK(clk), .Q(\mem[88][3] ) );
  DFF_X1 \mem_reg[88][2]  ( .D(n5922), .CK(clk), .Q(\mem[88][2] ) );
  DFF_X1 \mem_reg[88][1]  ( .D(n5923), .CK(clk), .Q(\mem[88][1] ) );
  DFF_X1 \mem_reg[88][0]  ( .D(n5924), .CK(clk), .Q(\mem[88][0] ) );
  DFF_X1 \mem_reg[87][7]  ( .D(n5925), .CK(clk), .Q(\mem[87][7] ) );
  DFF_X1 \mem_reg[87][6]  ( .D(n5926), .CK(clk), .Q(\mem[87][6] ) );
  DFF_X1 \mem_reg[87][5]  ( .D(n5927), .CK(clk), .Q(\mem[87][5] ) );
  DFF_X1 \mem_reg[87][4]  ( .D(n5928), .CK(clk), .Q(\mem[87][4] ) );
  DFF_X1 \mem_reg[87][3]  ( .D(n5929), .CK(clk), .Q(\mem[87][3] ) );
  DFF_X1 \mem_reg[87][2]  ( .D(n5930), .CK(clk), .Q(\mem[87][2] ) );
  DFF_X1 \mem_reg[87][1]  ( .D(n5931), .CK(clk), .Q(\mem[87][1] ) );
  DFF_X1 \mem_reg[87][0]  ( .D(n5932), .CK(clk), .Q(\mem[87][0] ) );
  DFF_X1 \mem_reg[86][7]  ( .D(n5933), .CK(clk), .Q(\mem[86][7] ) );
  DFF_X1 \mem_reg[86][6]  ( .D(n5934), .CK(clk), .Q(\mem[86][6] ) );
  DFF_X1 \mem_reg[86][5]  ( .D(n5935), .CK(clk), .Q(\mem[86][5] ) );
  DFF_X1 \mem_reg[86][4]  ( .D(n5936), .CK(clk), .Q(\mem[86][4] ) );
  DFF_X1 \mem_reg[86][3]  ( .D(n5937), .CK(clk), .Q(\mem[86][3] ) );
  DFF_X1 \mem_reg[86][2]  ( .D(n5938), .CK(clk), .Q(\mem[86][2] ) );
  DFF_X1 \mem_reg[86][1]  ( .D(n5939), .CK(clk), .Q(\mem[86][1] ) );
  DFF_X1 \mem_reg[86][0]  ( .D(n5940), .CK(clk), .Q(\mem[86][0] ) );
  DFF_X1 \mem_reg[85][7]  ( .D(n5941), .CK(clk), .Q(\mem[85][7] ) );
  DFF_X1 \mem_reg[85][6]  ( .D(n5942), .CK(clk), .Q(\mem[85][6] ) );
  DFF_X1 \mem_reg[85][5]  ( .D(n5943), .CK(clk), .Q(\mem[85][5] ) );
  DFF_X1 \mem_reg[85][4]  ( .D(n5944), .CK(clk), .Q(\mem[85][4] ) );
  DFF_X1 \mem_reg[85][3]  ( .D(n5945), .CK(clk), .Q(\mem[85][3] ) );
  DFF_X1 \mem_reg[85][2]  ( .D(n5946), .CK(clk), .Q(\mem[85][2] ) );
  DFF_X1 \mem_reg[85][1]  ( .D(n5947), .CK(clk), .Q(\mem[85][1] ) );
  DFF_X1 \mem_reg[85][0]  ( .D(n5948), .CK(clk), .Q(\mem[85][0] ) );
  DFF_X1 \mem_reg[84][7]  ( .D(n5949), .CK(clk), .Q(\mem[84][7] ) );
  DFF_X1 \mem_reg[84][6]  ( .D(n5950), .CK(clk), .Q(\mem[84][6] ) );
  DFF_X1 \mem_reg[84][5]  ( .D(n5951), .CK(clk), .Q(\mem[84][5] ) );
  DFF_X1 \mem_reg[84][4]  ( .D(n5952), .CK(clk), .Q(\mem[84][4] ) );
  DFF_X1 \mem_reg[84][3]  ( .D(n5953), .CK(clk), .Q(\mem[84][3] ) );
  DFF_X1 \mem_reg[84][2]  ( .D(n5954), .CK(clk), .Q(\mem[84][2] ) );
  DFF_X1 \mem_reg[84][1]  ( .D(n5955), .CK(clk), .Q(\mem[84][1] ) );
  DFF_X1 \mem_reg[84][0]  ( .D(n5956), .CK(clk), .Q(\mem[84][0] ) );
  DFF_X1 \mem_reg[83][7]  ( .D(n5957), .CK(clk), .Q(\mem[83][7] ) );
  DFF_X1 \mem_reg[83][6]  ( .D(n5958), .CK(clk), .Q(\mem[83][6] ) );
  DFF_X1 \mem_reg[83][5]  ( .D(n5959), .CK(clk), .Q(\mem[83][5] ) );
  DFF_X1 \mem_reg[83][4]  ( .D(n5960), .CK(clk), .Q(\mem[83][4] ) );
  DFF_X1 \mem_reg[83][3]  ( .D(n5961), .CK(clk), .Q(\mem[83][3] ) );
  DFF_X1 \mem_reg[83][2]  ( .D(n5962), .CK(clk), .Q(\mem[83][2] ) );
  DFF_X1 \mem_reg[83][1]  ( .D(n5963), .CK(clk), .Q(\mem[83][1] ) );
  DFF_X1 \mem_reg[83][0]  ( .D(n5964), .CK(clk), .Q(\mem[83][0] ) );
  DFF_X1 \mem_reg[82][7]  ( .D(n5965), .CK(clk), .Q(\mem[82][7] ) );
  DFF_X1 \mem_reg[82][6]  ( .D(n5966), .CK(clk), .Q(\mem[82][6] ) );
  DFF_X1 \mem_reg[82][5]  ( .D(n5967), .CK(clk), .Q(\mem[82][5] ) );
  DFF_X1 \mem_reg[82][4]  ( .D(n5968), .CK(clk), .Q(\mem[82][4] ) );
  DFF_X1 \mem_reg[82][3]  ( .D(n5969), .CK(clk), .Q(\mem[82][3] ) );
  DFF_X1 \mem_reg[82][2]  ( .D(n5970), .CK(clk), .Q(\mem[82][2] ) );
  DFF_X1 \mem_reg[82][1]  ( .D(n5971), .CK(clk), .Q(\mem[82][1] ) );
  DFF_X1 \mem_reg[82][0]  ( .D(n5972), .CK(clk), .Q(\mem[82][0] ) );
  DFF_X1 \mem_reg[81][7]  ( .D(n5973), .CK(clk), .Q(\mem[81][7] ) );
  DFF_X1 \mem_reg[81][6]  ( .D(n5974), .CK(clk), .Q(\mem[81][6] ) );
  DFF_X1 \mem_reg[81][5]  ( .D(n5975), .CK(clk), .Q(\mem[81][5] ) );
  DFF_X1 \mem_reg[81][4]  ( .D(n5976), .CK(clk), .Q(\mem[81][4] ) );
  DFF_X1 \mem_reg[81][3]  ( .D(n5977), .CK(clk), .Q(\mem[81][3] ) );
  DFF_X1 \mem_reg[81][2]  ( .D(n5978), .CK(clk), .Q(\mem[81][2] ) );
  DFF_X1 \mem_reg[81][1]  ( .D(n5979), .CK(clk), .Q(\mem[81][1] ) );
  DFF_X1 \mem_reg[81][0]  ( .D(n5980), .CK(clk), .Q(\mem[81][0] ) );
  DFF_X1 \mem_reg[80][7]  ( .D(n5981), .CK(clk), .Q(\mem[80][7] ) );
  DFF_X1 \mem_reg[80][6]  ( .D(n5982), .CK(clk), .Q(\mem[80][6] ) );
  DFF_X1 \mem_reg[80][5]  ( .D(n5983), .CK(clk), .Q(\mem[80][5] ) );
  DFF_X1 \mem_reg[80][4]  ( .D(n5984), .CK(clk), .Q(\mem[80][4] ) );
  DFF_X1 \mem_reg[80][3]  ( .D(n5985), .CK(clk), .Q(\mem[80][3] ) );
  DFF_X1 \mem_reg[80][2]  ( .D(n5986), .CK(clk), .Q(\mem[80][2] ) );
  DFF_X1 \mem_reg[80][1]  ( .D(n5987), .CK(clk), .Q(\mem[80][1] ) );
  DFF_X1 \mem_reg[80][0]  ( .D(n5988), .CK(clk), .Q(\mem[80][0] ) );
  DFF_X1 \mem_reg[79][7]  ( .D(n5989), .CK(clk), .Q(\mem[79][7] ) );
  DFF_X1 \mem_reg[79][6]  ( .D(n5990), .CK(clk), .Q(\mem[79][6] ) );
  DFF_X1 \mem_reg[79][5]  ( .D(n5991), .CK(clk), .Q(\mem[79][5] ) );
  DFF_X1 \mem_reg[79][4]  ( .D(n5992), .CK(clk), .Q(\mem[79][4] ) );
  DFF_X1 \mem_reg[79][3]  ( .D(n5993), .CK(clk), .Q(\mem[79][3] ) );
  DFF_X1 \mem_reg[79][2]  ( .D(n5994), .CK(clk), .Q(\mem[79][2] ) );
  DFF_X1 \mem_reg[79][1]  ( .D(n5995), .CK(clk), .Q(\mem[79][1] ) );
  DFF_X1 \mem_reg[79][0]  ( .D(n5996), .CK(clk), .Q(\mem[79][0] ) );
  DFF_X1 \mem_reg[78][7]  ( .D(n5997), .CK(clk), .Q(\mem[78][7] ) );
  DFF_X1 \mem_reg[78][6]  ( .D(n5998), .CK(clk), .Q(\mem[78][6] ) );
  DFF_X1 \mem_reg[78][5]  ( .D(n5999), .CK(clk), .Q(\mem[78][5] ) );
  DFF_X1 \mem_reg[78][4]  ( .D(n6000), .CK(clk), .Q(\mem[78][4] ) );
  DFF_X1 \mem_reg[78][3]  ( .D(n6001), .CK(clk), .Q(\mem[78][3] ) );
  DFF_X1 \mem_reg[78][2]  ( .D(n6002), .CK(clk), .Q(\mem[78][2] ) );
  DFF_X1 \mem_reg[78][1]  ( .D(n6003), .CK(clk), .Q(\mem[78][1] ) );
  DFF_X1 \mem_reg[78][0]  ( .D(n6004), .CK(clk), .Q(\mem[78][0] ) );
  DFF_X1 \mem_reg[77][7]  ( .D(n6005), .CK(clk), .Q(\mem[77][7] ) );
  DFF_X1 \mem_reg[77][6]  ( .D(n6006), .CK(clk), .Q(\mem[77][6] ) );
  DFF_X1 \mem_reg[77][5]  ( .D(n6007), .CK(clk), .Q(\mem[77][5] ) );
  DFF_X1 \mem_reg[77][4]  ( .D(n6008), .CK(clk), .Q(\mem[77][4] ) );
  DFF_X1 \mem_reg[77][3]  ( .D(n6009), .CK(clk), .Q(\mem[77][3] ) );
  DFF_X1 \mem_reg[77][2]  ( .D(n6010), .CK(clk), .Q(\mem[77][2] ) );
  DFF_X1 \mem_reg[77][1]  ( .D(n6011), .CK(clk), .Q(\mem[77][1] ) );
  DFF_X1 \mem_reg[77][0]  ( .D(n6012), .CK(clk), .Q(\mem[77][0] ) );
  DFF_X1 \mem_reg[76][7]  ( .D(n6013), .CK(clk), .Q(\mem[76][7] ) );
  DFF_X1 \mem_reg[76][6]  ( .D(n6014), .CK(clk), .Q(\mem[76][6] ) );
  DFF_X1 \mem_reg[76][5]  ( .D(n6015), .CK(clk), .Q(\mem[76][5] ) );
  DFF_X1 \mem_reg[76][4]  ( .D(n6016), .CK(clk), .Q(\mem[76][4] ) );
  DFF_X1 \mem_reg[76][3]  ( .D(n6017), .CK(clk), .Q(\mem[76][3] ) );
  DFF_X1 \mem_reg[76][2]  ( .D(n6018), .CK(clk), .Q(\mem[76][2] ) );
  DFF_X1 \mem_reg[76][1]  ( .D(n6019), .CK(clk), .Q(\mem[76][1] ) );
  DFF_X1 \mem_reg[76][0]  ( .D(n6020), .CK(clk), .Q(\mem[76][0] ) );
  DFF_X1 \mem_reg[75][7]  ( .D(n6021), .CK(clk), .Q(\mem[75][7] ) );
  DFF_X1 \mem_reg[75][6]  ( .D(n6022), .CK(clk), .Q(\mem[75][6] ) );
  DFF_X1 \mem_reg[75][5]  ( .D(n6023), .CK(clk), .Q(\mem[75][5] ) );
  DFF_X1 \mem_reg[75][4]  ( .D(n6024), .CK(clk), .Q(\mem[75][4] ) );
  DFF_X1 \mem_reg[75][3]  ( .D(n6025), .CK(clk), .Q(\mem[75][3] ) );
  DFF_X1 \mem_reg[75][2]  ( .D(n6026), .CK(clk), .Q(\mem[75][2] ) );
  DFF_X1 \mem_reg[75][1]  ( .D(n6027), .CK(clk), .Q(\mem[75][1] ) );
  DFF_X1 \mem_reg[75][0]  ( .D(n6028), .CK(clk), .Q(\mem[75][0] ) );
  DFF_X1 \mem_reg[74][7]  ( .D(n6029), .CK(clk), .Q(\mem[74][7] ) );
  DFF_X1 \mem_reg[74][6]  ( .D(n6030), .CK(clk), .Q(\mem[74][6] ) );
  DFF_X1 \mem_reg[74][5]  ( .D(n6031), .CK(clk), .Q(\mem[74][5] ) );
  DFF_X1 \mem_reg[74][4]  ( .D(n6032), .CK(clk), .Q(\mem[74][4] ) );
  DFF_X1 \mem_reg[74][3]  ( .D(n6033), .CK(clk), .Q(\mem[74][3] ) );
  DFF_X1 \mem_reg[74][2]  ( .D(n6034), .CK(clk), .Q(\mem[74][2] ) );
  DFF_X1 \mem_reg[74][1]  ( .D(n6035), .CK(clk), .Q(\mem[74][1] ) );
  DFF_X1 \mem_reg[74][0]  ( .D(n6036), .CK(clk), .Q(\mem[74][0] ) );
  DFF_X1 \mem_reg[73][7]  ( .D(n6037), .CK(clk), .Q(\mem[73][7] ) );
  DFF_X1 \mem_reg[73][6]  ( .D(n6038), .CK(clk), .Q(\mem[73][6] ) );
  DFF_X1 \mem_reg[73][5]  ( .D(n6039), .CK(clk), .Q(\mem[73][5] ) );
  DFF_X1 \mem_reg[73][4]  ( .D(n6040), .CK(clk), .Q(\mem[73][4] ) );
  DFF_X1 \mem_reg[73][3]  ( .D(n6041), .CK(clk), .Q(\mem[73][3] ) );
  DFF_X1 \mem_reg[73][2]  ( .D(n6042), .CK(clk), .Q(\mem[73][2] ) );
  DFF_X1 \mem_reg[73][1]  ( .D(n6043), .CK(clk), .Q(\mem[73][1] ) );
  DFF_X1 \mem_reg[73][0]  ( .D(n6044), .CK(clk), .Q(\mem[73][0] ) );
  DFF_X1 \mem_reg[72][7]  ( .D(n6045), .CK(clk), .Q(\mem[72][7] ) );
  DFF_X1 \mem_reg[72][6]  ( .D(n6046), .CK(clk), .Q(\mem[72][6] ) );
  DFF_X1 \mem_reg[72][5]  ( .D(n6047), .CK(clk), .Q(\mem[72][5] ) );
  DFF_X1 \mem_reg[72][4]  ( .D(n6048), .CK(clk), .Q(\mem[72][4] ) );
  DFF_X1 \mem_reg[72][3]  ( .D(n6049), .CK(clk), .Q(\mem[72][3] ) );
  DFF_X1 \mem_reg[72][2]  ( .D(n6050), .CK(clk), .Q(\mem[72][2] ) );
  DFF_X1 \mem_reg[72][1]  ( .D(n6051), .CK(clk), .Q(\mem[72][1] ) );
  DFF_X1 \mem_reg[72][0]  ( .D(n6052), .CK(clk), .Q(\mem[72][0] ) );
  DFF_X1 \mem_reg[71][7]  ( .D(n6053), .CK(clk), .Q(\mem[71][7] ) );
  DFF_X1 \mem_reg[71][6]  ( .D(n6054), .CK(clk), .Q(\mem[71][6] ) );
  DFF_X1 \mem_reg[71][5]  ( .D(n6055), .CK(clk), .Q(\mem[71][5] ) );
  DFF_X1 \mem_reg[71][4]  ( .D(n6056), .CK(clk), .Q(\mem[71][4] ) );
  DFF_X1 \mem_reg[71][3]  ( .D(n6057), .CK(clk), .Q(\mem[71][3] ) );
  DFF_X1 \mem_reg[71][2]  ( .D(n6058), .CK(clk), .Q(\mem[71][2] ) );
  DFF_X1 \mem_reg[71][1]  ( .D(n6059), .CK(clk), .Q(\mem[71][1] ) );
  DFF_X1 \mem_reg[71][0]  ( .D(n6060), .CK(clk), .Q(\mem[71][0] ) );
  DFF_X1 \mem_reg[70][7]  ( .D(n6061), .CK(clk), .Q(\mem[70][7] ) );
  DFF_X1 \mem_reg[70][6]  ( .D(n6062), .CK(clk), .Q(\mem[70][6] ) );
  DFF_X1 \mem_reg[70][5]  ( .D(n6063), .CK(clk), .Q(\mem[70][5] ) );
  DFF_X1 \mem_reg[70][4]  ( .D(n6064), .CK(clk), .Q(\mem[70][4] ) );
  DFF_X1 \mem_reg[70][3]  ( .D(n6065), .CK(clk), .Q(\mem[70][3] ) );
  DFF_X1 \mem_reg[70][2]  ( .D(n6066), .CK(clk), .Q(\mem[70][2] ) );
  DFF_X1 \mem_reg[70][1]  ( .D(n6067), .CK(clk), .Q(\mem[70][1] ) );
  DFF_X1 \mem_reg[70][0]  ( .D(n6068), .CK(clk), .Q(\mem[70][0] ) );
  DFF_X1 \mem_reg[69][7]  ( .D(n6069), .CK(clk), .Q(\mem[69][7] ) );
  DFF_X1 \mem_reg[69][6]  ( .D(n6070), .CK(clk), .Q(\mem[69][6] ) );
  DFF_X1 \mem_reg[69][5]  ( .D(n6071), .CK(clk), .Q(\mem[69][5] ) );
  DFF_X1 \mem_reg[69][4]  ( .D(n6072), .CK(clk), .Q(\mem[69][4] ) );
  DFF_X1 \mem_reg[69][3]  ( .D(n6073), .CK(clk), .Q(\mem[69][3] ) );
  DFF_X1 \mem_reg[69][2]  ( .D(n6074), .CK(clk), .Q(\mem[69][2] ) );
  DFF_X1 \mem_reg[69][1]  ( .D(n6075), .CK(clk), .Q(\mem[69][1] ) );
  DFF_X1 \mem_reg[69][0]  ( .D(n6076), .CK(clk), .Q(\mem[69][0] ) );
  DFF_X1 \mem_reg[68][7]  ( .D(n6077), .CK(clk), .Q(\mem[68][7] ) );
  DFF_X1 \mem_reg[68][6]  ( .D(n6078), .CK(clk), .Q(\mem[68][6] ) );
  DFF_X1 \mem_reg[68][5]  ( .D(n6079), .CK(clk), .Q(\mem[68][5] ) );
  DFF_X1 \mem_reg[68][4]  ( .D(n6080), .CK(clk), .Q(\mem[68][4] ) );
  DFF_X1 \mem_reg[68][3]  ( .D(n6081), .CK(clk), .Q(\mem[68][3] ) );
  DFF_X1 \mem_reg[68][2]  ( .D(n6082), .CK(clk), .Q(\mem[68][2] ) );
  DFF_X1 \mem_reg[68][1]  ( .D(n6083), .CK(clk), .Q(\mem[68][1] ) );
  DFF_X1 \mem_reg[68][0]  ( .D(n6084), .CK(clk), .Q(\mem[68][0] ) );
  DFF_X1 \mem_reg[67][7]  ( .D(n6085), .CK(clk), .Q(\mem[67][7] ) );
  DFF_X1 \mem_reg[67][6]  ( .D(n6086), .CK(clk), .Q(\mem[67][6] ) );
  DFF_X1 \mem_reg[67][5]  ( .D(n6087), .CK(clk), .Q(\mem[67][5] ) );
  DFF_X1 \mem_reg[67][4]  ( .D(n6088), .CK(clk), .Q(\mem[67][4] ) );
  DFF_X1 \mem_reg[67][3]  ( .D(n6089), .CK(clk), .Q(\mem[67][3] ) );
  DFF_X1 \mem_reg[67][2]  ( .D(n6090), .CK(clk), .Q(\mem[67][2] ) );
  DFF_X1 \mem_reg[67][1]  ( .D(n6091), .CK(clk), .Q(\mem[67][1] ) );
  DFF_X1 \mem_reg[67][0]  ( .D(n6092), .CK(clk), .Q(\mem[67][0] ) );
  DFF_X1 \mem_reg[66][7]  ( .D(n6093), .CK(clk), .Q(\mem[66][7] ) );
  DFF_X1 \mem_reg[66][6]  ( .D(n6094), .CK(clk), .Q(\mem[66][6] ) );
  DFF_X1 \mem_reg[66][5]  ( .D(n6095), .CK(clk), .Q(\mem[66][5] ) );
  DFF_X1 \mem_reg[66][4]  ( .D(n6096), .CK(clk), .Q(\mem[66][4] ) );
  DFF_X1 \mem_reg[66][3]  ( .D(n6097), .CK(clk), .Q(\mem[66][3] ) );
  DFF_X1 \mem_reg[66][2]  ( .D(n6098), .CK(clk), .Q(\mem[66][2] ) );
  DFF_X1 \mem_reg[66][1]  ( .D(n6099), .CK(clk), .Q(\mem[66][1] ) );
  DFF_X1 \mem_reg[66][0]  ( .D(n6100), .CK(clk), .Q(\mem[66][0] ) );
  DFF_X1 \mem_reg[65][7]  ( .D(n6101), .CK(clk), .Q(\mem[65][7] ) );
  DFF_X1 \mem_reg[65][6]  ( .D(n6102), .CK(clk), .Q(\mem[65][6] ) );
  DFF_X1 \mem_reg[65][5]  ( .D(n6103), .CK(clk), .Q(\mem[65][5] ) );
  DFF_X1 \mem_reg[65][4]  ( .D(n6104), .CK(clk), .Q(\mem[65][4] ) );
  DFF_X1 \mem_reg[65][3]  ( .D(n6105), .CK(clk), .Q(\mem[65][3] ) );
  DFF_X1 \mem_reg[65][2]  ( .D(n6106), .CK(clk), .Q(\mem[65][2] ) );
  DFF_X1 \mem_reg[65][1]  ( .D(n6107), .CK(clk), .Q(\mem[65][1] ) );
  DFF_X1 \mem_reg[65][0]  ( .D(n6108), .CK(clk), .Q(\mem[65][0] ) );
  DFF_X1 \mem_reg[64][7]  ( .D(n6109), .CK(clk), .Q(\mem[64][7] ) );
  DFF_X1 \mem_reg[64][6]  ( .D(n6110), .CK(clk), .Q(\mem[64][6] ) );
  DFF_X1 \mem_reg[64][5]  ( .D(n6111), .CK(clk), .Q(\mem[64][5] ) );
  DFF_X1 \mem_reg[64][4]  ( .D(n6112), .CK(clk), .Q(\mem[64][4] ) );
  DFF_X1 \mem_reg[64][3]  ( .D(n6113), .CK(clk), .Q(\mem[64][3] ) );
  DFF_X1 \mem_reg[64][2]  ( .D(n6114), .CK(clk), .Q(\mem[64][2] ) );
  DFF_X1 \mem_reg[64][1]  ( .D(n6115), .CK(clk), .Q(\mem[64][1] ) );
  DFF_X1 \mem_reg[64][0]  ( .D(n6116), .CK(clk), .Q(\mem[64][0] ) );
  DFF_X1 \mem_reg[63][7]  ( .D(n6117), .CK(clk), .Q(\mem[63][7] ) );
  DFF_X1 \mem_reg[63][6]  ( .D(n6118), .CK(clk), .Q(\mem[63][6] ) );
  DFF_X1 \mem_reg[63][5]  ( .D(n6119), .CK(clk), .Q(\mem[63][5] ) );
  DFF_X1 \mem_reg[63][4]  ( .D(n6120), .CK(clk), .Q(\mem[63][4] ) );
  DFF_X1 \mem_reg[63][3]  ( .D(n6121), .CK(clk), .Q(\mem[63][3] ) );
  DFF_X1 \mem_reg[63][2]  ( .D(n6122), .CK(clk), .Q(\mem[63][2] ) );
  DFF_X1 \mem_reg[63][1]  ( .D(n6123), .CK(clk), .Q(\mem[63][1] ) );
  DFF_X1 \mem_reg[63][0]  ( .D(n6124), .CK(clk), .Q(\mem[63][0] ) );
  DFF_X1 \mem_reg[62][7]  ( .D(n6125), .CK(clk), .Q(\mem[62][7] ) );
  DFF_X1 \mem_reg[62][6]  ( .D(n6126), .CK(clk), .Q(\mem[62][6] ) );
  DFF_X1 \mem_reg[62][5]  ( .D(n6127), .CK(clk), .Q(\mem[62][5] ) );
  DFF_X1 \mem_reg[62][4]  ( .D(n6128), .CK(clk), .Q(\mem[62][4] ) );
  DFF_X1 \mem_reg[62][3]  ( .D(n6129), .CK(clk), .Q(\mem[62][3] ) );
  DFF_X1 \mem_reg[62][2]  ( .D(n6130), .CK(clk), .Q(\mem[62][2] ) );
  DFF_X1 \mem_reg[62][1]  ( .D(n6131), .CK(clk), .Q(\mem[62][1] ) );
  DFF_X1 \mem_reg[62][0]  ( .D(n6132), .CK(clk), .Q(\mem[62][0] ) );
  DFF_X1 \mem_reg[61][7]  ( .D(n6133), .CK(clk), .Q(\mem[61][7] ) );
  DFF_X1 \mem_reg[61][6]  ( .D(n6134), .CK(clk), .Q(\mem[61][6] ) );
  DFF_X1 \mem_reg[61][5]  ( .D(n6135), .CK(clk), .Q(\mem[61][5] ) );
  DFF_X1 \mem_reg[61][4]  ( .D(n6136), .CK(clk), .Q(\mem[61][4] ) );
  DFF_X1 \mem_reg[61][3]  ( .D(n6137), .CK(clk), .Q(\mem[61][3] ) );
  DFF_X1 \mem_reg[61][2]  ( .D(n6138), .CK(clk), .Q(\mem[61][2] ) );
  DFF_X1 \mem_reg[61][1]  ( .D(n6139), .CK(clk), .Q(\mem[61][1] ) );
  DFF_X1 \mem_reg[61][0]  ( .D(n6140), .CK(clk), .Q(\mem[61][0] ) );
  DFF_X1 \mem_reg[60][7]  ( .D(n6141), .CK(clk), .Q(\mem[60][7] ) );
  DFF_X1 \mem_reg[60][6]  ( .D(n6142), .CK(clk), .Q(\mem[60][6] ) );
  DFF_X1 \mem_reg[60][5]  ( .D(n6143), .CK(clk), .Q(\mem[60][5] ) );
  DFF_X1 \mem_reg[60][4]  ( .D(n6144), .CK(clk), .Q(\mem[60][4] ) );
  DFF_X1 \mem_reg[60][3]  ( .D(n6145), .CK(clk), .Q(\mem[60][3] ) );
  DFF_X1 \mem_reg[60][2]  ( .D(n6146), .CK(clk), .Q(\mem[60][2] ) );
  DFF_X1 \mem_reg[60][1]  ( .D(n6147), .CK(clk), .Q(\mem[60][1] ) );
  DFF_X1 \mem_reg[60][0]  ( .D(n6148), .CK(clk), .Q(\mem[60][0] ) );
  DFF_X1 \mem_reg[59][7]  ( .D(n6149), .CK(clk), .Q(\mem[59][7] ) );
  DFF_X1 \mem_reg[59][6]  ( .D(n6150), .CK(clk), .Q(\mem[59][6] ) );
  DFF_X1 \mem_reg[59][5]  ( .D(n6151), .CK(clk), .Q(\mem[59][5] ) );
  DFF_X1 \mem_reg[59][4]  ( .D(n6152), .CK(clk), .Q(\mem[59][4] ) );
  DFF_X1 \mem_reg[59][3]  ( .D(n6153), .CK(clk), .Q(\mem[59][3] ) );
  DFF_X1 \mem_reg[59][2]  ( .D(n6154), .CK(clk), .Q(\mem[59][2] ) );
  DFF_X1 \mem_reg[59][1]  ( .D(n6155), .CK(clk), .Q(\mem[59][1] ) );
  DFF_X1 \mem_reg[59][0]  ( .D(n6156), .CK(clk), .Q(\mem[59][0] ) );
  DFF_X1 \mem_reg[58][7]  ( .D(n6157), .CK(clk), .Q(\mem[58][7] ) );
  DFF_X1 \mem_reg[58][6]  ( .D(n6158), .CK(clk), .Q(\mem[58][6] ) );
  DFF_X1 \mem_reg[58][5]  ( .D(n6159), .CK(clk), .Q(\mem[58][5] ) );
  DFF_X1 \mem_reg[58][4]  ( .D(n6160), .CK(clk), .Q(\mem[58][4] ) );
  DFF_X1 \mem_reg[58][3]  ( .D(n6161), .CK(clk), .Q(\mem[58][3] ) );
  DFF_X1 \mem_reg[58][2]  ( .D(n6162), .CK(clk), .Q(\mem[58][2] ) );
  DFF_X1 \mem_reg[58][1]  ( .D(n6163), .CK(clk), .Q(\mem[58][1] ) );
  DFF_X1 \mem_reg[58][0]  ( .D(n6164), .CK(clk), .Q(\mem[58][0] ) );
  DFF_X1 \mem_reg[57][7]  ( .D(n6165), .CK(clk), .Q(\mem[57][7] ) );
  DFF_X1 \mem_reg[57][6]  ( .D(n6166), .CK(clk), .Q(\mem[57][6] ) );
  DFF_X1 \mem_reg[57][5]  ( .D(n6167), .CK(clk), .Q(\mem[57][5] ) );
  DFF_X1 \mem_reg[57][4]  ( .D(n6168), .CK(clk), .Q(\mem[57][4] ) );
  DFF_X1 \mem_reg[57][3]  ( .D(n6169), .CK(clk), .Q(\mem[57][3] ) );
  DFF_X1 \mem_reg[57][2]  ( .D(n6170), .CK(clk), .Q(\mem[57][2] ) );
  DFF_X1 \mem_reg[57][1]  ( .D(n6171), .CK(clk), .Q(\mem[57][1] ) );
  DFF_X1 \mem_reg[57][0]  ( .D(n6172), .CK(clk), .Q(\mem[57][0] ) );
  DFF_X1 \mem_reg[56][7]  ( .D(n6173), .CK(clk), .Q(\mem[56][7] ) );
  DFF_X1 \mem_reg[56][6]  ( .D(n6174), .CK(clk), .Q(\mem[56][6] ) );
  DFF_X1 \mem_reg[56][5]  ( .D(n6175), .CK(clk), .Q(\mem[56][5] ) );
  DFF_X1 \mem_reg[56][4]  ( .D(n6176), .CK(clk), .Q(\mem[56][4] ) );
  DFF_X1 \mem_reg[56][3]  ( .D(n6177), .CK(clk), .Q(\mem[56][3] ) );
  DFF_X1 \mem_reg[56][2]  ( .D(n6178), .CK(clk), .Q(\mem[56][2] ) );
  DFF_X1 \mem_reg[56][1]  ( .D(n6179), .CK(clk), .Q(\mem[56][1] ) );
  DFF_X1 \mem_reg[56][0]  ( .D(n6180), .CK(clk), .Q(\mem[56][0] ) );
  DFF_X1 \mem_reg[55][7]  ( .D(n6181), .CK(clk), .Q(\mem[55][7] ) );
  DFF_X1 \mem_reg[55][6]  ( .D(n6182), .CK(clk), .Q(\mem[55][6] ) );
  DFF_X1 \mem_reg[55][5]  ( .D(n6183), .CK(clk), .Q(\mem[55][5] ) );
  DFF_X1 \mem_reg[55][4]  ( .D(n6184), .CK(clk), .Q(\mem[55][4] ) );
  DFF_X1 \mem_reg[55][3]  ( .D(n6185), .CK(clk), .Q(\mem[55][3] ) );
  DFF_X1 \mem_reg[55][2]  ( .D(n6186), .CK(clk), .Q(\mem[55][2] ) );
  DFF_X1 \mem_reg[55][1]  ( .D(n6187), .CK(clk), .Q(\mem[55][1] ) );
  DFF_X1 \mem_reg[55][0]  ( .D(n6188), .CK(clk), .Q(\mem[55][0] ) );
  DFF_X1 \mem_reg[54][7]  ( .D(n6189), .CK(clk), .Q(\mem[54][7] ) );
  DFF_X1 \mem_reg[54][6]  ( .D(n6190), .CK(clk), .Q(\mem[54][6] ) );
  DFF_X1 \mem_reg[54][5]  ( .D(n6191), .CK(clk), .Q(\mem[54][5] ) );
  DFF_X1 \mem_reg[54][4]  ( .D(n6192), .CK(clk), .Q(\mem[54][4] ) );
  DFF_X1 \mem_reg[54][3]  ( .D(n6193), .CK(clk), .Q(\mem[54][3] ) );
  DFF_X1 \mem_reg[54][2]  ( .D(n6194), .CK(clk), .Q(\mem[54][2] ) );
  DFF_X1 \mem_reg[54][1]  ( .D(n6195), .CK(clk), .Q(\mem[54][1] ) );
  DFF_X1 \mem_reg[54][0]  ( .D(n6196), .CK(clk), .Q(\mem[54][0] ) );
  DFF_X1 \mem_reg[53][7]  ( .D(n6197), .CK(clk), .Q(\mem[53][7] ) );
  DFF_X1 \mem_reg[53][6]  ( .D(n6198), .CK(clk), .Q(\mem[53][6] ) );
  DFF_X1 \mem_reg[53][5]  ( .D(n6199), .CK(clk), .Q(\mem[53][5] ) );
  DFF_X1 \mem_reg[53][4]  ( .D(n6200), .CK(clk), .Q(\mem[53][4] ) );
  DFF_X1 \mem_reg[53][3]  ( .D(n6201), .CK(clk), .Q(\mem[53][3] ) );
  DFF_X1 \mem_reg[53][2]  ( .D(n6202), .CK(clk), .Q(\mem[53][2] ) );
  DFF_X1 \mem_reg[53][1]  ( .D(n6203), .CK(clk), .Q(\mem[53][1] ) );
  DFF_X1 \mem_reg[53][0]  ( .D(n6204), .CK(clk), .Q(\mem[53][0] ) );
  DFF_X1 \mem_reg[52][7]  ( .D(n6205), .CK(clk), .Q(\mem[52][7] ) );
  DFF_X1 \mem_reg[52][6]  ( .D(n6206), .CK(clk), .Q(\mem[52][6] ) );
  DFF_X1 \mem_reg[52][5]  ( .D(n6207), .CK(clk), .Q(\mem[52][5] ) );
  DFF_X1 \mem_reg[52][4]  ( .D(n6208), .CK(clk), .Q(\mem[52][4] ) );
  DFF_X1 \mem_reg[52][3]  ( .D(n6209), .CK(clk), .Q(\mem[52][3] ) );
  DFF_X1 \mem_reg[52][2]  ( .D(n6210), .CK(clk), .Q(\mem[52][2] ) );
  DFF_X1 \mem_reg[52][1]  ( .D(n6211), .CK(clk), .Q(\mem[52][1] ) );
  DFF_X1 \mem_reg[52][0]  ( .D(n6212), .CK(clk), .Q(\mem[52][0] ) );
  DFF_X1 \mem_reg[51][7]  ( .D(n6213), .CK(clk), .Q(\mem[51][7] ) );
  DFF_X1 \mem_reg[51][6]  ( .D(n6214), .CK(clk), .Q(\mem[51][6] ) );
  DFF_X1 \mem_reg[51][5]  ( .D(n6215), .CK(clk), .Q(\mem[51][5] ) );
  DFF_X1 \mem_reg[51][4]  ( .D(n6216), .CK(clk), .Q(\mem[51][4] ) );
  DFF_X1 \mem_reg[51][3]  ( .D(n6217), .CK(clk), .Q(\mem[51][3] ) );
  DFF_X1 \mem_reg[51][2]  ( .D(n6218), .CK(clk), .Q(\mem[51][2] ) );
  DFF_X1 \mem_reg[51][1]  ( .D(n6219), .CK(clk), .Q(\mem[51][1] ) );
  DFF_X1 \mem_reg[51][0]  ( .D(n6220), .CK(clk), .Q(\mem[51][0] ) );
  DFF_X1 \mem_reg[50][7]  ( .D(n6221), .CK(clk), .Q(\mem[50][7] ) );
  DFF_X1 \mem_reg[50][6]  ( .D(n6222), .CK(clk), .Q(\mem[50][6] ) );
  DFF_X1 \mem_reg[50][5]  ( .D(n6223), .CK(clk), .Q(\mem[50][5] ) );
  DFF_X1 \mem_reg[50][4]  ( .D(n6224), .CK(clk), .Q(\mem[50][4] ) );
  DFF_X1 \mem_reg[50][3]  ( .D(n6225), .CK(clk), .Q(\mem[50][3] ) );
  DFF_X1 \mem_reg[50][2]  ( .D(n6226), .CK(clk), .Q(\mem[50][2] ) );
  DFF_X1 \mem_reg[50][1]  ( .D(n6227), .CK(clk), .Q(\mem[50][1] ) );
  DFF_X1 \mem_reg[50][0]  ( .D(n6228), .CK(clk), .Q(\mem[50][0] ) );
  DFF_X1 \mem_reg[49][7]  ( .D(n6229), .CK(clk), .Q(\mem[49][7] ) );
  DFF_X1 \mem_reg[49][6]  ( .D(n6230), .CK(clk), .Q(\mem[49][6] ) );
  DFF_X1 \mem_reg[49][5]  ( .D(n6231), .CK(clk), .Q(\mem[49][5] ) );
  DFF_X1 \mem_reg[49][4]  ( .D(n6232), .CK(clk), .Q(\mem[49][4] ) );
  DFF_X1 \mem_reg[49][3]  ( .D(n6233), .CK(clk), .Q(\mem[49][3] ) );
  DFF_X1 \mem_reg[49][2]  ( .D(n6234), .CK(clk), .Q(\mem[49][2] ) );
  DFF_X1 \mem_reg[49][1]  ( .D(n6235), .CK(clk), .Q(\mem[49][1] ) );
  DFF_X1 \mem_reg[49][0]  ( .D(n6236), .CK(clk), .Q(\mem[49][0] ) );
  DFF_X1 \mem_reg[48][7]  ( .D(n6237), .CK(clk), .Q(\mem[48][7] ) );
  DFF_X1 \mem_reg[48][6]  ( .D(n6238), .CK(clk), .Q(\mem[48][6] ) );
  DFF_X1 \mem_reg[48][5]  ( .D(n6239), .CK(clk), .Q(\mem[48][5] ) );
  DFF_X1 \mem_reg[48][4]  ( .D(n6240), .CK(clk), .Q(\mem[48][4] ) );
  DFF_X1 \mem_reg[48][3]  ( .D(n6241), .CK(clk), .Q(\mem[48][3] ) );
  DFF_X1 \mem_reg[48][2]  ( .D(n6242), .CK(clk), .Q(\mem[48][2] ) );
  DFF_X1 \mem_reg[48][1]  ( .D(n6243), .CK(clk), .Q(\mem[48][1] ) );
  DFF_X1 \mem_reg[48][0]  ( .D(n6244), .CK(clk), .Q(\mem[48][0] ) );
  DFF_X1 \mem_reg[47][7]  ( .D(n6245), .CK(clk), .Q(\mem[47][7] ) );
  DFF_X1 \mem_reg[47][6]  ( .D(n6246), .CK(clk), .Q(\mem[47][6] ) );
  DFF_X1 \mem_reg[47][5]  ( .D(n6247), .CK(clk), .Q(\mem[47][5] ) );
  DFF_X1 \mem_reg[47][4]  ( .D(n6248), .CK(clk), .Q(\mem[47][4] ) );
  DFF_X1 \mem_reg[47][3]  ( .D(n6249), .CK(clk), .Q(\mem[47][3] ) );
  DFF_X1 \mem_reg[47][2]  ( .D(n6250), .CK(clk), .Q(\mem[47][2] ) );
  DFF_X1 \mem_reg[47][1]  ( .D(n6251), .CK(clk), .Q(\mem[47][1] ) );
  DFF_X1 \mem_reg[47][0]  ( .D(n6252), .CK(clk), .Q(\mem[47][0] ) );
  DFF_X1 \mem_reg[46][7]  ( .D(n6253), .CK(clk), .Q(\mem[46][7] ) );
  DFF_X1 \mem_reg[46][6]  ( .D(n6254), .CK(clk), .Q(\mem[46][6] ) );
  DFF_X1 \mem_reg[46][5]  ( .D(n6255), .CK(clk), .Q(\mem[46][5] ) );
  DFF_X1 \mem_reg[46][4]  ( .D(n6256), .CK(clk), .Q(\mem[46][4] ) );
  DFF_X1 \mem_reg[46][3]  ( .D(n6257), .CK(clk), .Q(\mem[46][3] ) );
  DFF_X1 \mem_reg[46][2]  ( .D(n6258), .CK(clk), .Q(\mem[46][2] ) );
  DFF_X1 \mem_reg[46][1]  ( .D(n6259), .CK(clk), .Q(\mem[46][1] ) );
  DFF_X1 \mem_reg[46][0]  ( .D(n6260), .CK(clk), .Q(\mem[46][0] ) );
  DFF_X1 \mem_reg[45][7]  ( .D(n6261), .CK(clk), .Q(\mem[45][7] ) );
  DFF_X1 \mem_reg[45][6]  ( .D(n6262), .CK(clk), .Q(\mem[45][6] ) );
  DFF_X1 \mem_reg[45][5]  ( .D(n6263), .CK(clk), .Q(\mem[45][5] ) );
  DFF_X1 \mem_reg[45][4]  ( .D(n6264), .CK(clk), .Q(\mem[45][4] ) );
  DFF_X1 \mem_reg[45][3]  ( .D(n6265), .CK(clk), .Q(\mem[45][3] ) );
  DFF_X1 \mem_reg[45][2]  ( .D(n6266), .CK(clk), .Q(\mem[45][2] ) );
  DFF_X1 \mem_reg[45][1]  ( .D(n6267), .CK(clk), .Q(\mem[45][1] ) );
  DFF_X1 \mem_reg[45][0]  ( .D(n6268), .CK(clk), .Q(\mem[45][0] ) );
  DFF_X1 \mem_reg[44][7]  ( .D(n6269), .CK(clk), .Q(\mem[44][7] ) );
  DFF_X1 \mem_reg[44][6]  ( .D(n6270), .CK(clk), .Q(\mem[44][6] ) );
  DFF_X1 \mem_reg[44][5]  ( .D(n6271), .CK(clk), .Q(\mem[44][5] ) );
  DFF_X1 \mem_reg[44][4]  ( .D(n6272), .CK(clk), .Q(\mem[44][4] ) );
  DFF_X1 \mem_reg[44][3]  ( .D(n6273), .CK(clk), .Q(\mem[44][3] ) );
  DFF_X1 \mem_reg[44][2]  ( .D(n6274), .CK(clk), .Q(\mem[44][2] ) );
  DFF_X1 \mem_reg[44][1]  ( .D(n6275), .CK(clk), .Q(\mem[44][1] ) );
  DFF_X1 \mem_reg[44][0]  ( .D(n6276), .CK(clk), .Q(\mem[44][0] ) );
  DFF_X1 \mem_reg[43][7]  ( .D(n6277), .CK(clk), .Q(\mem[43][7] ) );
  DFF_X1 \mem_reg[43][6]  ( .D(n6278), .CK(clk), .Q(\mem[43][6] ) );
  DFF_X1 \mem_reg[43][5]  ( .D(n6279), .CK(clk), .Q(\mem[43][5] ) );
  DFF_X1 \mem_reg[43][4]  ( .D(n6280), .CK(clk), .Q(\mem[43][4] ) );
  DFF_X1 \mem_reg[43][3]  ( .D(n6281), .CK(clk), .Q(\mem[43][3] ) );
  DFF_X1 \mem_reg[43][2]  ( .D(n6282), .CK(clk), .Q(\mem[43][2] ) );
  DFF_X1 \mem_reg[43][1]  ( .D(n6283), .CK(clk), .Q(\mem[43][1] ) );
  DFF_X1 \mem_reg[43][0]  ( .D(n6284), .CK(clk), .Q(\mem[43][0] ) );
  DFF_X1 \mem_reg[42][7]  ( .D(n6285), .CK(clk), .Q(\mem[42][7] ) );
  DFF_X1 \mem_reg[42][6]  ( .D(n6286), .CK(clk), .Q(\mem[42][6] ) );
  DFF_X1 \mem_reg[42][5]  ( .D(n6287), .CK(clk), .Q(\mem[42][5] ) );
  DFF_X1 \mem_reg[42][4]  ( .D(n6288), .CK(clk), .Q(\mem[42][4] ) );
  DFF_X1 \mem_reg[42][3]  ( .D(n6289), .CK(clk), .Q(\mem[42][3] ) );
  DFF_X1 \mem_reg[42][2]  ( .D(n6290), .CK(clk), .Q(\mem[42][2] ) );
  DFF_X1 \mem_reg[42][1]  ( .D(n6291), .CK(clk), .Q(\mem[42][1] ) );
  DFF_X1 \mem_reg[42][0]  ( .D(n6292), .CK(clk), .Q(\mem[42][0] ) );
  DFF_X1 \mem_reg[41][7]  ( .D(n6293), .CK(clk), .Q(\mem[41][7] ) );
  DFF_X1 \mem_reg[41][6]  ( .D(n6294), .CK(clk), .Q(\mem[41][6] ) );
  DFF_X1 \mem_reg[41][5]  ( .D(n6295), .CK(clk), .Q(\mem[41][5] ) );
  DFF_X1 \mem_reg[41][4]  ( .D(n6296), .CK(clk), .Q(\mem[41][4] ) );
  DFF_X1 \mem_reg[41][3]  ( .D(n6297), .CK(clk), .Q(\mem[41][3] ) );
  DFF_X1 \mem_reg[41][2]  ( .D(n6298), .CK(clk), .Q(\mem[41][2] ) );
  DFF_X1 \mem_reg[41][1]  ( .D(n6299), .CK(clk), .Q(\mem[41][1] ) );
  DFF_X1 \mem_reg[41][0]  ( .D(n6300), .CK(clk), .Q(\mem[41][0] ) );
  DFF_X1 \mem_reg[40][7]  ( .D(n6301), .CK(clk), .Q(\mem[40][7] ) );
  DFF_X1 \mem_reg[40][6]  ( .D(n6302), .CK(clk), .Q(\mem[40][6] ) );
  DFF_X1 \mem_reg[40][5]  ( .D(n6303), .CK(clk), .Q(\mem[40][5] ) );
  DFF_X1 \mem_reg[40][4]  ( .D(n6304), .CK(clk), .Q(\mem[40][4] ) );
  DFF_X1 \mem_reg[40][3]  ( .D(n6305), .CK(clk), .Q(\mem[40][3] ) );
  DFF_X1 \mem_reg[40][2]  ( .D(n6306), .CK(clk), .Q(\mem[40][2] ) );
  DFF_X1 \mem_reg[40][1]  ( .D(n6307), .CK(clk), .Q(\mem[40][1] ) );
  DFF_X1 \mem_reg[40][0]  ( .D(n6308), .CK(clk), .Q(\mem[40][0] ) );
  DFF_X1 \mem_reg[39][7]  ( .D(n6309), .CK(clk), .Q(\mem[39][7] ) );
  DFF_X1 \mem_reg[39][6]  ( .D(n6310), .CK(clk), .Q(\mem[39][6] ) );
  DFF_X1 \mem_reg[39][5]  ( .D(n6311), .CK(clk), .Q(\mem[39][5] ) );
  DFF_X1 \mem_reg[39][4]  ( .D(n6312), .CK(clk), .Q(\mem[39][4] ) );
  DFF_X1 \mem_reg[39][3]  ( .D(n6313), .CK(clk), .Q(\mem[39][3] ) );
  DFF_X1 \mem_reg[39][2]  ( .D(n6314), .CK(clk), .Q(\mem[39][2] ) );
  DFF_X1 \mem_reg[39][1]  ( .D(n6315), .CK(clk), .Q(\mem[39][1] ) );
  DFF_X1 \mem_reg[39][0]  ( .D(n6316), .CK(clk), .Q(\mem[39][0] ) );
  DFF_X1 \mem_reg[38][7]  ( .D(n6317), .CK(clk), .Q(\mem[38][7] ) );
  DFF_X1 \mem_reg[38][6]  ( .D(n6318), .CK(clk), .Q(\mem[38][6] ) );
  DFF_X1 \mem_reg[38][5]  ( .D(n6319), .CK(clk), .Q(\mem[38][5] ) );
  DFF_X1 \mem_reg[38][4]  ( .D(n6320), .CK(clk), .Q(\mem[38][4] ) );
  DFF_X1 \mem_reg[38][3]  ( .D(n6321), .CK(clk), .Q(\mem[38][3] ) );
  DFF_X1 \mem_reg[38][2]  ( .D(n6322), .CK(clk), .Q(\mem[38][2] ) );
  DFF_X1 \mem_reg[38][1]  ( .D(n6323), .CK(clk), .Q(\mem[38][1] ) );
  DFF_X1 \mem_reg[38][0]  ( .D(n6324), .CK(clk), .Q(\mem[38][0] ) );
  DFF_X1 \mem_reg[37][7]  ( .D(n6325), .CK(clk), .Q(\mem[37][7] ) );
  DFF_X1 \mem_reg[37][6]  ( .D(n6326), .CK(clk), .Q(\mem[37][6] ) );
  DFF_X1 \mem_reg[37][5]  ( .D(n6327), .CK(clk), .Q(\mem[37][5] ) );
  DFF_X1 \mem_reg[37][4]  ( .D(n6328), .CK(clk), .Q(\mem[37][4] ) );
  DFF_X1 \mem_reg[37][3]  ( .D(n6329), .CK(clk), .Q(\mem[37][3] ) );
  DFF_X1 \mem_reg[37][2]  ( .D(n6330), .CK(clk), .Q(\mem[37][2] ) );
  DFF_X1 \mem_reg[37][1]  ( .D(n6331), .CK(clk), .Q(\mem[37][1] ) );
  DFF_X1 \mem_reg[37][0]  ( .D(n6332), .CK(clk), .Q(\mem[37][0] ) );
  DFF_X1 \mem_reg[36][7]  ( .D(n6333), .CK(clk), .Q(\mem[36][7] ) );
  DFF_X1 \mem_reg[36][6]  ( .D(n6334), .CK(clk), .Q(\mem[36][6] ) );
  DFF_X1 \mem_reg[36][5]  ( .D(n6335), .CK(clk), .Q(\mem[36][5] ) );
  DFF_X1 \mem_reg[36][4]  ( .D(n6336), .CK(clk), .Q(\mem[36][4] ) );
  DFF_X1 \mem_reg[36][3]  ( .D(n6337), .CK(clk), .Q(\mem[36][3] ) );
  DFF_X1 \mem_reg[36][2]  ( .D(n6338), .CK(clk), .Q(\mem[36][2] ) );
  DFF_X1 \mem_reg[36][1]  ( .D(n6339), .CK(clk), .Q(\mem[36][1] ) );
  DFF_X1 \mem_reg[36][0]  ( .D(n6340), .CK(clk), .Q(\mem[36][0] ) );
  DFF_X1 \mem_reg[35][7]  ( .D(n6341), .CK(clk), .Q(\mem[35][7] ) );
  DFF_X1 \mem_reg[35][6]  ( .D(n6342), .CK(clk), .Q(\mem[35][6] ) );
  DFF_X1 \mem_reg[35][5]  ( .D(n6343), .CK(clk), .Q(\mem[35][5] ) );
  DFF_X1 \mem_reg[35][4]  ( .D(n6344), .CK(clk), .Q(\mem[35][4] ) );
  DFF_X1 \mem_reg[35][3]  ( .D(n6345), .CK(clk), .Q(\mem[35][3] ) );
  DFF_X1 \mem_reg[35][2]  ( .D(n6346), .CK(clk), .Q(\mem[35][2] ) );
  DFF_X1 \mem_reg[35][1]  ( .D(n6347), .CK(clk), .Q(\mem[35][1] ) );
  DFF_X1 \mem_reg[35][0]  ( .D(n6348), .CK(clk), .Q(\mem[35][0] ) );
  DFF_X1 \mem_reg[34][7]  ( .D(n6349), .CK(clk), .Q(\mem[34][7] ) );
  DFF_X1 \mem_reg[34][6]  ( .D(n6350), .CK(clk), .Q(\mem[34][6] ) );
  DFF_X1 \mem_reg[34][5]  ( .D(n6351), .CK(clk), .Q(\mem[34][5] ) );
  DFF_X1 \mem_reg[34][4]  ( .D(n6352), .CK(clk), .Q(\mem[34][4] ) );
  DFF_X1 \mem_reg[34][3]  ( .D(n6353), .CK(clk), .Q(\mem[34][3] ) );
  DFF_X1 \mem_reg[34][2]  ( .D(n6354), .CK(clk), .Q(\mem[34][2] ) );
  DFF_X1 \mem_reg[34][1]  ( .D(n6355), .CK(clk), .Q(\mem[34][1] ) );
  DFF_X1 \mem_reg[34][0]  ( .D(n6356), .CK(clk), .Q(\mem[34][0] ) );
  DFF_X1 \mem_reg[33][7]  ( .D(n6357), .CK(clk), .Q(\mem[33][7] ) );
  DFF_X1 \mem_reg[33][6]  ( .D(n6358), .CK(clk), .Q(\mem[33][6] ) );
  DFF_X1 \mem_reg[33][5]  ( .D(n6359), .CK(clk), .Q(\mem[33][5] ) );
  DFF_X1 \mem_reg[33][4]  ( .D(n6360), .CK(clk), .Q(\mem[33][4] ) );
  DFF_X1 \mem_reg[33][3]  ( .D(n6361), .CK(clk), .Q(\mem[33][3] ) );
  DFF_X1 \mem_reg[33][2]  ( .D(n6362), .CK(clk), .Q(\mem[33][2] ) );
  DFF_X1 \mem_reg[33][1]  ( .D(n6363), .CK(clk), .Q(\mem[33][1] ) );
  DFF_X1 \mem_reg[33][0]  ( .D(n6364), .CK(clk), .Q(\mem[33][0] ) );
  DFF_X1 \mem_reg[32][7]  ( .D(n6365), .CK(clk), .Q(\mem[32][7] ) );
  DFF_X1 \mem_reg[32][6]  ( .D(n6366), .CK(clk), .Q(\mem[32][6] ) );
  DFF_X1 \mem_reg[32][5]  ( .D(n6367), .CK(clk), .Q(\mem[32][5] ) );
  DFF_X1 \mem_reg[32][4]  ( .D(n6368), .CK(clk), .Q(\mem[32][4] ) );
  DFF_X1 \mem_reg[32][3]  ( .D(n6369), .CK(clk), .Q(\mem[32][3] ) );
  DFF_X1 \mem_reg[32][2]  ( .D(n6370), .CK(clk), .Q(\mem[32][2] ) );
  DFF_X1 \mem_reg[32][1]  ( .D(n6371), .CK(clk), .Q(\mem[32][1] ) );
  DFF_X1 \mem_reg[32][0]  ( .D(n6372), .CK(clk), .Q(\mem[32][0] ) );
  DFF_X1 \mem_reg[31][7]  ( .D(n6373), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n6374), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n6375), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n6376), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n6377), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n6378), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n6379), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n6380), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n6381), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n6382), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n6383), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n6384), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n6385), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n6386), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n6387), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n6388), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n6389), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n6390), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n6391), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n6392), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n6393), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n6394), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n6395), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n6396), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n6397), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n6398), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n6399), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n6400), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n6401), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n6402), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n6403), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n6404), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n6405), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n6406), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n6407), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n6408), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n6409), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n6410), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n6411), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n6412), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n6413), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n6414), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n6415), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n6416), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n6417), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n6418), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n6419), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n6420), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n6421), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n6422), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n6423), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n6424), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n6425), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n6426), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n6427), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n6428), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n6429), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n6430), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n6431), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n6432), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n6433), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n6434), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n6435), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n6436), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n6437), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n6438), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n6439), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n6440), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n6441), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n6442), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n6443), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n6444), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n6445), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n6446), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n6447), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n6448), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n6449), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n6450), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n6451), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n6452), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n6453), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n6454), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n6455), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n6456), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n6457), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n6458), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n6459), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n6460), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n6461), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n6462), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n6463), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n6464), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n6465), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n6466), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n6467), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n6468), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n6469), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n6470), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n6471), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n6472), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n6473), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n6474), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n6475), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n6476), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n6477), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n6478), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n6479), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n6480), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n6481), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n6482), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n6483), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n6484), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n6485), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n6486), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n6487), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n6488), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n6489), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n6490), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n6491), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n6492), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n6493), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n6494), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n6495), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n6496), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n6497), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n6498), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n6499), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n6500), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n6501), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n6502), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n6503), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n6504), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n6505), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n6506), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n6507), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n6508), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n6509), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n6510), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n6511), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n6512), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n6513), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n6514), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n6515), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n6516), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n6517), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n6518), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n6519), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n6520), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n6521), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n6522), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n6523), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n6524), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n6525), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n6526), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n6527), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n6528), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n6529), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n6530), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n6531), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n6532), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n6533), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n6534), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n6535), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n6536), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n6537), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n6538), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n6539), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n6540), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n6541), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n6542), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n6543), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n6544), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n6545), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n6546), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n6547), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n6548), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n6549), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n6550), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n6551), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n6552), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n6553), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n6554), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n6555), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n6556), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n6557), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n6558), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n6559), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n6560), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n6561), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n6562), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n6563), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n6564), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n6565), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n6566), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n6567), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n6568), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n6569), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n6570), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n6571), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n6572), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n6573), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n6574), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n6575), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n6576), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n6577), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n6578), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n6579), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n6580), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n6581), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n6582), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n6583), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n6584), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n6585), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n6586), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n6587), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n6588), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n6589), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n6590), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n6591), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n6592), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n6593), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n6594), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n6595), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n6596), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n6597), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n6598), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n6599), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n6600), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n6601), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n6602), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n6603), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n6604), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n6605), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n6606), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n6607), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n6608), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n6609), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n6610), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n6611), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n6612), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n6613), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n6614), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n6615), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n6616), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n6617), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n6618), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n6619), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n6620), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n6621), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n6622), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n6623), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n6624), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n6625), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n6626), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n6627), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n6628), .CK(clk), .Q(\mem[0][0] ) );
  AND3_X2 U205 ( .A1(wr_en), .A2(n2534), .A3(n2535), .ZN(n2389) );
  AND3_X2 U350 ( .A1(n2681), .A2(wr_en), .A3(n2682), .ZN(n2545) );
  AND3_X2 U495 ( .A1(n2682), .A2(wr_en), .A3(n2828), .ZN(n2692) );
  AND3_X2 U640 ( .A1(wr_en), .A2(n2974), .A3(n2682), .ZN(n2838) );
  AND3_X2 U785 ( .A1(n2535), .A2(wr_en), .A3(n2682), .ZN(n2984) );
  AND3_X2 U931 ( .A1(n2681), .A2(wr_en), .A3(n3265), .ZN(n3129) );
  AND3_X2 U1076 ( .A1(n2828), .A2(wr_en), .A3(n3265), .ZN(n3275) );
  AND3_X2 U1221 ( .A1(wr_en), .A2(n2974), .A3(n3265), .ZN(n3420) );
  AND3_X2 U1366 ( .A1(n2535), .A2(wr_en), .A3(n3265), .ZN(n3565) );
  AND3_X2 U1512 ( .A1(n2681), .A2(wr_en), .A3(n3846), .ZN(n3710) );
  AND3_X2 U1657 ( .A1(n2828), .A2(wr_en), .A3(n3846), .ZN(n3856) );
  AND3_X2 U1802 ( .A1(wr_en), .A2(n2974), .A3(n3846), .ZN(n4001) );
  AND3_X2 U1947 ( .A1(n2535), .A2(wr_en), .A3(n3846), .ZN(n4146) );
  AND3_X2 U2094 ( .A1(wr_en), .A2(n2534), .A3(n2681), .ZN(n4291) );
  AND3_X2 U2247 ( .A1(wr_en), .A2(n2534), .A3(n2828), .ZN(n4436) );
  AND3_X2 U2349 ( .A1(n2534), .A2(n2974), .A3(wr_en), .ZN(n2328) );
  SDFF_X1 \data_out_reg[1]  ( .D(n396), .SI(n523), .SE(n11), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n1412), .SI(n1539), .SE(n11), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[2]  ( .D(n650), .SI(n777), .SE(n11), .CK(clk), .Q(
        data_out[2]) );
  SDFF_X1 \data_out_reg[4]  ( .D(n1158), .SI(n1285), .SE(n11), .CK(clk), .Q(
        data_out[4]) );
  SDFF_X1 \data_out_reg[6]  ( .D(n1666), .SI(n1793), .SE(n11), .CK(clk), .Q(
        data_out[6]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n1920), .SI(n2047), .SE(n11), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n904), .SI(n1031), .SE(n11), .CK(clk), .Q(
        data_out[3]) );
  BUF_X1 U3 ( .A(n2088), .Z(n2070) );
  CLKBUF_X1 U4 ( .A(n2087), .Z(n2091) );
  BUF_X1 U5 ( .A(n2099), .Z(n2100) );
  BUF_X1 U6 ( .A(n2219), .Z(n2142) );
  BUF_X2 U7 ( .A(n2143), .Z(n2177) );
  BUF_X1 U8 ( .A(n2222), .Z(n2182) );
  BUF_X2 U9 ( .A(n2144), .Z(n2153) );
  BUF_X1 U10 ( .A(n2147), .Z(n2197) );
  BUF_X1 U11 ( .A(n2141), .Z(n2191) );
  BUF_X2 U12 ( .A(n2139), .Z(n2205) );
  BUF_X2 U13 ( .A(n2139), .Z(n1) );
  NOR2_X1 U14 ( .A1(n6885), .A2(N25), .ZN(n3265) );
  AND2_X2 U15 ( .A1(n4587), .A2(n4527), .ZN(n2409) );
  AND2_X2 U16 ( .A1(n4624), .A2(n4549), .ZN(n2429) );
  AND2_X2 U17 ( .A1(n4624), .A2(n4527), .ZN(n2449) );
  AND2_X2 U18 ( .A1(n4548), .A2(n4549), .ZN(n2348) );
  AND2_X2 U19 ( .A1(n4548), .A2(n4527), .ZN(n2368) );
  BUF_X2 U20 ( .A(n14), .Z(n2147) );
  CLKBUF_X3 U21 ( .A(n2215), .Z(n2145) );
  BUF_X1 U22 ( .A(n2216), .Z(n2218) );
  BUF_X1 U23 ( .A(n2222), .Z(n2183) );
  CLKBUF_X2 U24 ( .A(n12), .Z(n2206) );
  CLKBUF_X1 U25 ( .A(n14), .Z(n2146) );
  CLKBUF_X2 U26 ( .A(n2219), .Z(n2141) );
  BUF_X1 U27 ( .A(n2217), .Z(n2138) );
  BUF_X2 U28 ( .A(n2145), .Z(n2210) );
  CLKBUF_X1 U29 ( .A(N18), .Z(n2216) );
  CLKBUF_X3 U30 ( .A(n2144), .Z(n2174) );
  BUF_X4 U31 ( .A(n13), .Z(n2154) );
  BUF_X4 U32 ( .A(n12), .Z(n2155) );
  CLKBUF_X3 U33 ( .A(n2144), .Z(n2184) );
  INV_X1 U34 ( .A(n2191), .ZN(n2) );
  BUF_X1 U35 ( .A(n2144), .Z(n3) );
  BUF_X1 U36 ( .A(n2144), .Z(n4) );
  CLKBUF_X3 U37 ( .A(n2215), .Z(n2144) );
  CLKBUF_X3 U38 ( .A(n2142), .Z(n2190) );
  CLKBUF_X3 U39 ( .A(n2144), .Z(n2175) );
  CLKBUF_X3 U40 ( .A(n2142), .Z(n2188) );
  CLKBUF_X3 U41 ( .A(n2144), .Z(n2173) );
  CLKBUF_X3 U42 ( .A(n2142), .Z(n2189) );
  CLKBUF_X3 U43 ( .A(n2144), .Z(n2172) );
  CLKBUF_X3 U44 ( .A(n2147), .Z(n2148) );
  CLKBUF_X3 U45 ( .A(n2219), .Z(n2200) );
  CLKBUF_X3 U46 ( .A(n2139), .Z(n2199) );
  NAND2_X1 U47 ( .A1(n1727), .A2(n2227), .ZN(n5) );
  NAND2_X1 U48 ( .A1(n1712), .A2(n2056), .ZN(n6) );
  NAND2_X1 U49 ( .A1(n5), .A2(n6), .ZN(n1728) );
  CLKBUF_X3 U50 ( .A(n2137), .Z(n2214) );
  BUF_X1 U51 ( .A(n2145), .Z(n7) );
  BUF_X1 U52 ( .A(n2145), .Z(n8) );
  CLKBUF_X3 U53 ( .A(n2146), .Z(n2151) );
  CLKBUF_X3 U54 ( .A(n2146), .Z(n2150) );
  CLKBUF_X3 U55 ( .A(n2146), .Z(n2152) );
  CLKBUF_X3 U56 ( .A(n2138), .Z(n2208) );
  BUF_X2 U57 ( .A(n2138), .Z(n2212) );
  BUF_X1 U58 ( .A(n2217), .Z(n2137) );
  CLKBUF_X1 U59 ( .A(N18), .Z(n2215) );
  AND2_X1 U60 ( .A1(n4587), .A2(n4538), .ZN(n2419) );
  AND2_X1 U61 ( .A1(n4624), .A2(n4538), .ZN(n2459) );
  AND2_X1 U62 ( .A1(n4548), .A2(n4538), .ZN(n2378) );
  AND2_X1 U63 ( .A1(n4538), .A2(n4528), .ZN(n2338) );
  AND2_X1 U64 ( .A1(n4587), .A2(n4559), .ZN(n2399) );
  AND2_X1 U65 ( .A1(n4624), .A2(n4559), .ZN(n2439) );
  AND2_X1 U66 ( .A1(n4548), .A2(n4559), .ZN(n2358) );
  AND2_X1 U67 ( .A1(n4528), .A2(n4559), .ZN(n2479) );
  NAND2_X1 U68 ( .A1(n680), .A2(n2227), .ZN(n9) );
  NAND2_X1 U69 ( .A1(n665), .A2(n2053), .ZN(n10) );
  NAND2_X1 U70 ( .A1(n9), .A2(n10), .ZN(n681) );
  CLKBUF_X1 U71 ( .A(n13), .Z(n2186) );
  CLKBUF_X1 U72 ( .A(n13), .Z(n2187) );
  CLKBUF_X1 U73 ( .A(n12), .Z(n2185) );
  CLKBUF_X3 U74 ( .A(n2137), .Z(n2213) );
  MUX2_X1 U75 ( .A(n713), .B(n776), .S(n6885), .Z(n777) );
  INV_X1 U76 ( .A(N25), .ZN(n11) );
  CLKBUF_X3 U77 ( .A(n2138), .Z(n2170) );
  CLKBUF_X3 U78 ( .A(n2147), .Z(n2149) );
  INV_X1 U79 ( .A(n2223), .ZN(n2222) );
  CLKBUF_X3 U80 ( .A(n2147), .Z(n2164) );
  CLKBUF_X3 U81 ( .A(n2138), .Z(n2211) );
  CLKBUF_X3 U82 ( .A(n2138), .Z(n2209) );
  CLKBUF_X3 U83 ( .A(n2141), .Z(n2196) );
  CLKBUF_X3 U84 ( .A(n2141), .Z(n2195) );
  CLKBUF_X3 U85 ( .A(n2141), .Z(n2192) );
  CLKBUF_X3 U86 ( .A(n2141), .Z(n2193) );
  CLKBUF_X3 U87 ( .A(n2141), .Z(n2194) );
  CLKBUF_X3 U88 ( .A(n2218), .Z(n2201) );
  INV_X1 U89 ( .A(n2223), .ZN(n12) );
  CLKBUF_X1 U90 ( .A(n2217), .Z(n2139) );
  INV_X1 U91 ( .A(n2223), .ZN(n13) );
  BUF_X2 U92 ( .A(n2218), .Z(n2198) );
  INV_X1 U93 ( .A(n2223), .ZN(n14) );
  BUF_X1 U94 ( .A(N21), .Z(n2068) );
  BUF_X1 U95 ( .A(n2222), .Z(n2159) );
  BUF_X1 U96 ( .A(n2143), .Z(n2181) );
  BUF_X1 U97 ( .A(n2143), .Z(n2179) );
  BUF_X1 U98 ( .A(n2145), .Z(n2169) );
  BUF_X1 U99 ( .A(n2143), .Z(n2180) );
  BUF_X1 U100 ( .A(n2145), .Z(n2165) );
  BUF_X1 U101 ( .A(n2145), .Z(n2163) );
  BUF_X1 U102 ( .A(n13), .Z(n2207) );
  BUF_X1 U103 ( .A(n12), .Z(n2157) );
  BUF_X1 U104 ( .A(n2145), .Z(n2171) );
  BUF_X1 U105 ( .A(n2222), .Z(n2158) );
  BUF_X1 U106 ( .A(n2145), .Z(n2168) );
  BUF_X1 U107 ( .A(n2143), .Z(n2178) );
  BUF_X1 U108 ( .A(n2222), .Z(n2204) );
  BUF_X1 U109 ( .A(n13), .Z(n2203) );
  BUF_X1 U110 ( .A(n12), .Z(n2202) );
  BUF_X1 U111 ( .A(n2147), .Z(n2162) );
  BUF_X1 U112 ( .A(n2145), .Z(n2167) );
  BUF_X1 U113 ( .A(n2143), .Z(n2176) );
  BUF_X1 U114 ( .A(n2145), .Z(n2166) );
  BUF_X1 U115 ( .A(n12), .Z(n2156) );
  BUF_X1 U116 ( .A(n2144), .Z(n2161) );
  BUF_X1 U117 ( .A(n2145), .Z(n2160) );
  BUF_X1 U118 ( .A(n2091), .Z(n2084) );
  BUF_X1 U119 ( .A(n2089), .Z(n2078) );
  BUF_X1 U120 ( .A(n2094), .Z(n2128) );
  BUF_X1 U121 ( .A(n2097), .Z(n2111) );
  BUF_X1 U122 ( .A(n2091), .Z(n2086) );
  BUF_X1 U123 ( .A(n2090), .Z(n2083) );
  BUF_X1 U124 ( .A(n2091), .Z(n2085) );
  BUF_X1 U125 ( .A(n2089), .Z(n2079) );
  BUF_X1 U126 ( .A(n2095), .Z(n2122) );
  BUF_X1 U127 ( .A(n2089), .Z(n2077) );
  BUF_X1 U128 ( .A(n2095), .Z(n2120) );
  BUF_X1 U129 ( .A(n2095), .Z(n2123) );
  BUF_X1 U130 ( .A(n2096), .Z(n2115) );
  BUF_X1 U131 ( .A(n2094), .Z(n2127) );
  BUF_X1 U132 ( .A(n2096), .Z(n2116) );
  BUF_X1 U133 ( .A(n2094), .Z(n2126) );
  BUF_X1 U134 ( .A(n2095), .Z(n2121) );
  BUF_X1 U135 ( .A(n2096), .Z(n2118) );
  BUF_X1 U136 ( .A(n2098), .Z(n2108) );
  BUF_X1 U137 ( .A(n2099), .Z(n2129) );
  BUF_X1 U138 ( .A(n2094), .Z(n2125) );
  BUF_X1 U139 ( .A(n2093), .Z(n2132) );
  BUF_X1 U140 ( .A(n2098), .Z(n2107) );
  BUF_X1 U141 ( .A(n2097), .Z(n2113) );
  BUF_X1 U142 ( .A(n2096), .Z(n2117) );
  BUF_X1 U143 ( .A(n2098), .Z(n2109) );
  BUF_X1 U144 ( .A(n2097), .Z(n2112) );
  BUF_X1 U145 ( .A(n2098), .Z(n2106) );
  BUF_X1 U146 ( .A(n2093), .Z(n2131) );
  BUF_X1 U147 ( .A(n2099), .Z(n2103) );
  BUF_X1 U148 ( .A(n2099), .Z(n2102) );
  BUF_X1 U149 ( .A(n2099), .Z(n2104) );
  BUF_X1 U150 ( .A(n2089), .Z(n2076) );
  BUF_X1 U151 ( .A(n2090), .Z(n2082) );
  BUF_X1 U152 ( .A(n2090), .Z(n2081) );
  BUF_X1 U153 ( .A(n2089), .Z(n2075) );
  BUF_X1 U154 ( .A(n2098), .Z(n2105) );
  BUF_X1 U155 ( .A(n2090), .Z(n2080) );
  BUF_X1 U156 ( .A(n2095), .Z(n2119) );
  BUF_X1 U157 ( .A(n2089), .Z(n2074) );
  BUF_X1 U158 ( .A(n2097), .Z(n2110) );
  BUF_X1 U159 ( .A(n2094), .Z(n2124) );
  BUF_X1 U160 ( .A(n2096), .Z(n2114) );
  BUF_X1 U161 ( .A(n2093), .Z(n2130) );
  BUF_X1 U162 ( .A(n2092), .Z(n2133) );
  BUF_X1 U163 ( .A(n2092), .Z(n2134) );
  BUF_X1 U164 ( .A(n2099), .Z(n2101) );
  BUF_X1 U165 ( .A(n2088), .Z(n2073) );
  BUF_X1 U166 ( .A(n2088), .Z(n2071) );
  BUF_X1 U167 ( .A(n2088), .Z(n2072) );
  BUF_X1 U168 ( .A(n2218), .Z(n2140) );
  BUF_X1 U169 ( .A(n2215), .Z(n2143) );
  AND2_X1 U170 ( .A1(n4587), .A2(n4549), .ZN(n2388) );
  INV_X1 U171 ( .A(n2314), .ZN(n6629) );
  INV_X1 U172 ( .A(n2319), .ZN(n6644) );
  BUF_X1 U173 ( .A(n2069), .Z(n2066) );
  BUF_X1 U174 ( .A(n2069), .Z(n2065) );
  BUF_X1 U175 ( .A(n2069), .Z(n2067) );
  INV_X1 U176 ( .A(n2471), .ZN(n6875) );
  INV_X1 U177 ( .A(n2481), .ZN(n6874) );
  INV_X1 U178 ( .A(n2490), .ZN(n6873) );
  INV_X1 U179 ( .A(n2499), .ZN(n6872) );
  INV_X1 U180 ( .A(n2508), .ZN(n6871) );
  INV_X1 U181 ( .A(n2517), .ZN(n6870) );
  INV_X1 U182 ( .A(n2526), .ZN(n6869) );
  INV_X1 U183 ( .A(n2830), .ZN(n6836) );
  INV_X1 U184 ( .A(n2840), .ZN(n6835) );
  INV_X1 U185 ( .A(n2849), .ZN(n6834) );
  INV_X1 U186 ( .A(n2858), .ZN(n6833) );
  INV_X1 U187 ( .A(n2867), .ZN(n6832) );
  INV_X1 U188 ( .A(n2876), .ZN(n6831) );
  INV_X1 U189 ( .A(n2885), .ZN(n6830) );
  INV_X1 U190 ( .A(n2894), .ZN(n6829) );
  INV_X1 U191 ( .A(n2903), .ZN(n6828) );
  INV_X1 U192 ( .A(n2912), .ZN(n6827) );
  INV_X1 U193 ( .A(n2921), .ZN(n6826) );
  INV_X1 U194 ( .A(n2930), .ZN(n6825) );
  INV_X1 U195 ( .A(n2939), .ZN(n6824) );
  INV_X1 U196 ( .A(n2948), .ZN(n6823) );
  INV_X1 U197 ( .A(n2957), .ZN(n6822) );
  INV_X1 U198 ( .A(n2966), .ZN(n6821) );
  INV_X1 U199 ( .A(n3412), .ZN(n6772) );
  INV_X1 U200 ( .A(n3422), .ZN(n6771) );
  INV_X1 U201 ( .A(n3431), .ZN(n6770) );
  INV_X1 U202 ( .A(n3440), .ZN(n6769) );
  INV_X1 U203 ( .A(n3449), .ZN(n6768) );
  INV_X1 U204 ( .A(n3458), .ZN(n6767) );
  INV_X1 U206 ( .A(n3467), .ZN(n6766) );
  INV_X1 U207 ( .A(n3476), .ZN(n6765) );
  INV_X1 U208 ( .A(n3485), .ZN(n6764) );
  INV_X1 U209 ( .A(n3494), .ZN(n6763) );
  INV_X1 U210 ( .A(n3503), .ZN(n6762) );
  INV_X1 U211 ( .A(n3512), .ZN(n6761) );
  INV_X1 U212 ( .A(n3521), .ZN(n6760) );
  INV_X1 U213 ( .A(n3530), .ZN(n6759) );
  INV_X1 U214 ( .A(n3539), .ZN(n6758) );
  INV_X1 U215 ( .A(n3548), .ZN(n6757) );
  INV_X1 U216 ( .A(n3993), .ZN(n6708) );
  INV_X1 U217 ( .A(n4003), .ZN(n6707) );
  INV_X1 U218 ( .A(n4012), .ZN(n6706) );
  INV_X1 U219 ( .A(n4021), .ZN(n6705) );
  INV_X1 U220 ( .A(n4030), .ZN(n6704) );
  INV_X1 U221 ( .A(n4039), .ZN(n6703) );
  INV_X1 U222 ( .A(n4048), .ZN(n6702) );
  INV_X1 U223 ( .A(n4057), .ZN(n6701) );
  INV_X1 U224 ( .A(n4066), .ZN(n6700) );
  INV_X1 U225 ( .A(n4075), .ZN(n6699) );
  INV_X1 U226 ( .A(n4084), .ZN(n6698) );
  INV_X1 U227 ( .A(n4093), .ZN(n6697) );
  INV_X1 U228 ( .A(n4102), .ZN(n6696) );
  INV_X1 U229 ( .A(n4111), .ZN(n6695) );
  INV_X1 U230 ( .A(n4120), .ZN(n6694) );
  INV_X1 U231 ( .A(n4129), .ZN(n6693) );
  INV_X1 U232 ( .A(n4283), .ZN(n6676) );
  INV_X1 U233 ( .A(n4293), .ZN(n6675) );
  INV_X1 U234 ( .A(n4302), .ZN(n6674) );
  INV_X1 U235 ( .A(n4311), .ZN(n6673) );
  INV_X1 U236 ( .A(n4320), .ZN(n6672) );
  INV_X1 U237 ( .A(n4329), .ZN(n6671) );
  INV_X1 U238 ( .A(n4338), .ZN(n6670) );
  INV_X1 U239 ( .A(n4347), .ZN(n6669) );
  INV_X1 U240 ( .A(n4356), .ZN(n6668) );
  INV_X1 U241 ( .A(n4365), .ZN(n6667) );
  INV_X1 U242 ( .A(n4374), .ZN(n6666) );
  INV_X1 U243 ( .A(n4383), .ZN(n6665) );
  INV_X1 U244 ( .A(n4392), .ZN(n6664) );
  INV_X1 U245 ( .A(n4401), .ZN(n6663) );
  INV_X1 U246 ( .A(n4410), .ZN(n6662) );
  INV_X1 U247 ( .A(n4419), .ZN(n6661) );
  INV_X1 U248 ( .A(n4428), .ZN(n6660) );
  INV_X1 U249 ( .A(n4438), .ZN(n6659) );
  INV_X1 U250 ( .A(n4447), .ZN(n6658) );
  INV_X1 U251 ( .A(n4456), .ZN(n6657) );
  INV_X1 U252 ( .A(n4465), .ZN(n6656) );
  INV_X1 U253 ( .A(n4474), .ZN(n6655) );
  INV_X1 U254 ( .A(n4483), .ZN(n6654) );
  INV_X1 U255 ( .A(n4492), .ZN(n6653) );
  INV_X1 U256 ( .A(n4501), .ZN(n6652) );
  INV_X1 U257 ( .A(n4510), .ZN(n6651) );
  INV_X1 U258 ( .A(n4519), .ZN(n6650) );
  INV_X1 U259 ( .A(n4530), .ZN(n6649) );
  INV_X1 U260 ( .A(n4540), .ZN(n6648) );
  INV_X1 U261 ( .A(n4551), .ZN(n6647) );
  INV_X1 U262 ( .A(n4561), .ZN(n6646) );
  INV_X1 U263 ( .A(n4570), .ZN(n6645) );
  INV_X1 U264 ( .A(n2537), .ZN(n6868) );
  INV_X1 U265 ( .A(n2547), .ZN(n6867) );
  INV_X1 U266 ( .A(n2556), .ZN(n6866) );
  INV_X1 U267 ( .A(n2565), .ZN(n6865) );
  INV_X1 U268 ( .A(n2574), .ZN(n6864) );
  INV_X1 U269 ( .A(n2583), .ZN(n6863) );
  INV_X1 U270 ( .A(n2592), .ZN(n6862) );
  INV_X1 U271 ( .A(n2601), .ZN(n6861) );
  INV_X1 U272 ( .A(n2610), .ZN(n6860) );
  INV_X1 U273 ( .A(n2619), .ZN(n6859) );
  INV_X1 U274 ( .A(n2628), .ZN(n6858) );
  INV_X1 U275 ( .A(n2637), .ZN(n6857) );
  INV_X1 U276 ( .A(n2646), .ZN(n6856) );
  INV_X1 U277 ( .A(n2655), .ZN(n6855) );
  INV_X1 U278 ( .A(n2664), .ZN(n6854) );
  INV_X1 U279 ( .A(n2673), .ZN(n6853) );
  INV_X1 U280 ( .A(n2684), .ZN(n6852) );
  INV_X1 U281 ( .A(n2694), .ZN(n6851) );
  INV_X1 U282 ( .A(n2703), .ZN(n6850) );
  INV_X1 U283 ( .A(n2712), .ZN(n6849) );
  INV_X1 U284 ( .A(n2721), .ZN(n6848) );
  INV_X1 U285 ( .A(n2730), .ZN(n6847) );
  INV_X1 U286 ( .A(n2739), .ZN(n6846) );
  INV_X1 U287 ( .A(n2748), .ZN(n6845) );
  INV_X1 U288 ( .A(n2757), .ZN(n6844) );
  INV_X1 U289 ( .A(n2766), .ZN(n6843) );
  INV_X1 U290 ( .A(n2775), .ZN(n6842) );
  INV_X1 U291 ( .A(n2784), .ZN(n6841) );
  INV_X1 U292 ( .A(n2793), .ZN(n6840) );
  INV_X1 U293 ( .A(n2802), .ZN(n6839) );
  INV_X1 U294 ( .A(n2811), .ZN(n6838) );
  INV_X1 U295 ( .A(n2820), .ZN(n6837) );
  INV_X1 U296 ( .A(n2976), .ZN(n6820) );
  INV_X1 U297 ( .A(n2986), .ZN(n6819) );
  INV_X1 U298 ( .A(n2995), .ZN(n6818) );
  INV_X1 U299 ( .A(n3004), .ZN(n6817) );
  INV_X1 U300 ( .A(n3013), .ZN(n6816) );
  INV_X1 U301 ( .A(n3022), .ZN(n6815) );
  INV_X1 U302 ( .A(n3031), .ZN(n6814) );
  INV_X1 U303 ( .A(n3040), .ZN(n6813) );
  INV_X1 U304 ( .A(n3049), .ZN(n6812) );
  INV_X1 U305 ( .A(n3058), .ZN(n6811) );
  INV_X1 U306 ( .A(n3067), .ZN(n6810) );
  INV_X1 U307 ( .A(n3076), .ZN(n6809) );
  INV_X1 U308 ( .A(n3085), .ZN(n6808) );
  INV_X1 U309 ( .A(n3094), .ZN(n6807) );
  INV_X1 U310 ( .A(n3103), .ZN(n6806) );
  INV_X1 U311 ( .A(n3112), .ZN(n6805) );
  INV_X1 U312 ( .A(n3121), .ZN(n6804) );
  INV_X1 U313 ( .A(n3131), .ZN(n6803) );
  INV_X1 U314 ( .A(n3140), .ZN(n6802) );
  INV_X1 U315 ( .A(n3149), .ZN(n6801) );
  INV_X1 U316 ( .A(n3158), .ZN(n6800) );
  INV_X1 U317 ( .A(n3167), .ZN(n6799) );
  INV_X1 U318 ( .A(n3176), .ZN(n6798) );
  INV_X1 U319 ( .A(n3185), .ZN(n6797) );
  INV_X1 U320 ( .A(n3194), .ZN(n6796) );
  INV_X1 U321 ( .A(n3203), .ZN(n6795) );
  INV_X1 U322 ( .A(n3212), .ZN(n6794) );
  INV_X1 U323 ( .A(n3221), .ZN(n6793) );
  INV_X1 U324 ( .A(n3230), .ZN(n6792) );
  INV_X1 U325 ( .A(n3239), .ZN(n6791) );
  INV_X1 U326 ( .A(n3248), .ZN(n6790) );
  INV_X1 U327 ( .A(n3257), .ZN(n6789) );
  INV_X1 U328 ( .A(n3267), .ZN(n6788) );
  INV_X1 U329 ( .A(n3277), .ZN(n6787) );
  INV_X1 U330 ( .A(n3286), .ZN(n6786) );
  INV_X1 U331 ( .A(n3295), .ZN(n6785) );
  INV_X1 U332 ( .A(n3304), .ZN(n6784) );
  INV_X1 U333 ( .A(n3313), .ZN(n6783) );
  INV_X1 U334 ( .A(n3322), .ZN(n6782) );
  INV_X1 U335 ( .A(n3331), .ZN(n6781) );
  INV_X1 U336 ( .A(n3340), .ZN(n6780) );
  INV_X1 U337 ( .A(n3349), .ZN(n6779) );
  INV_X1 U338 ( .A(n3358), .ZN(n6778) );
  INV_X1 U339 ( .A(n3367), .ZN(n6777) );
  INV_X1 U340 ( .A(n3376), .ZN(n6776) );
  INV_X1 U341 ( .A(n3385), .ZN(n6775) );
  INV_X1 U342 ( .A(n3394), .ZN(n6774) );
  INV_X1 U343 ( .A(n3403), .ZN(n6773) );
  INV_X1 U344 ( .A(n3557), .ZN(n6756) );
  INV_X1 U345 ( .A(n3567), .ZN(n6755) );
  INV_X1 U346 ( .A(n3576), .ZN(n6754) );
  INV_X1 U347 ( .A(n3585), .ZN(n6753) );
  INV_X1 U348 ( .A(n3594), .ZN(n6752) );
  INV_X1 U349 ( .A(n3603), .ZN(n6751) );
  INV_X1 U351 ( .A(n3612), .ZN(n6750) );
  INV_X1 U352 ( .A(n3621), .ZN(n6749) );
  INV_X1 U353 ( .A(n3630), .ZN(n6748) );
  INV_X1 U354 ( .A(n3639), .ZN(n6747) );
  INV_X1 U355 ( .A(n3648), .ZN(n6746) );
  INV_X1 U356 ( .A(n3657), .ZN(n6745) );
  INV_X1 U357 ( .A(n3666), .ZN(n6744) );
  INV_X1 U358 ( .A(n3675), .ZN(n6743) );
  INV_X1 U359 ( .A(n3684), .ZN(n6742) );
  INV_X1 U360 ( .A(n3693), .ZN(n6741) );
  INV_X1 U361 ( .A(n3702), .ZN(n6740) );
  INV_X1 U362 ( .A(n3712), .ZN(n6739) );
  INV_X1 U363 ( .A(n3721), .ZN(n6738) );
  INV_X1 U364 ( .A(n3730), .ZN(n6737) );
  INV_X1 U365 ( .A(n3739), .ZN(n6736) );
  INV_X1 U366 ( .A(n3748), .ZN(n6735) );
  INV_X1 U367 ( .A(n3757), .ZN(n6734) );
  INV_X1 U368 ( .A(n3766), .ZN(n6733) );
  INV_X1 U369 ( .A(n3775), .ZN(n6732) );
  INV_X1 U370 ( .A(n3784), .ZN(n6731) );
  INV_X1 U371 ( .A(n3793), .ZN(n6730) );
  INV_X1 U372 ( .A(n3802), .ZN(n6729) );
  INV_X1 U373 ( .A(n3811), .ZN(n6728) );
  INV_X1 U374 ( .A(n3820), .ZN(n6727) );
  INV_X1 U375 ( .A(n3829), .ZN(n6726) );
  INV_X1 U376 ( .A(n3838), .ZN(n6725) );
  INV_X1 U377 ( .A(n3848), .ZN(n6724) );
  INV_X1 U378 ( .A(n3858), .ZN(n6723) );
  INV_X1 U379 ( .A(n3867), .ZN(n6722) );
  INV_X1 U380 ( .A(n3876), .ZN(n6721) );
  INV_X1 U381 ( .A(n3885), .ZN(n6720) );
  INV_X1 U382 ( .A(n3894), .ZN(n6719) );
  INV_X1 U383 ( .A(n3903), .ZN(n6718) );
  INV_X1 U384 ( .A(n3912), .ZN(n6717) );
  INV_X1 U385 ( .A(n3921), .ZN(n6716) );
  INV_X1 U386 ( .A(n3930), .ZN(n6715) );
  INV_X1 U387 ( .A(n3939), .ZN(n6714) );
  INV_X1 U388 ( .A(n3948), .ZN(n6713) );
  INV_X1 U389 ( .A(n3957), .ZN(n6712) );
  INV_X1 U390 ( .A(n3966), .ZN(n6711) );
  INV_X1 U391 ( .A(n3975), .ZN(n6710) );
  INV_X1 U392 ( .A(n3984), .ZN(n6709) );
  INV_X1 U393 ( .A(n4138), .ZN(n6692) );
  INV_X1 U394 ( .A(n4148), .ZN(n6691) );
  INV_X1 U395 ( .A(n4157), .ZN(n6690) );
  INV_X1 U396 ( .A(n4166), .ZN(n6689) );
  INV_X1 U397 ( .A(n4175), .ZN(n6688) );
  INV_X1 U398 ( .A(n4184), .ZN(n6687) );
  INV_X1 U399 ( .A(n4193), .ZN(n6686) );
  INV_X1 U400 ( .A(n4202), .ZN(n6685) );
  INV_X1 U401 ( .A(n4211), .ZN(n6684) );
  INV_X1 U402 ( .A(n4220), .ZN(n6683) );
  INV_X1 U403 ( .A(n4229), .ZN(n6682) );
  INV_X1 U404 ( .A(n4238), .ZN(n6681) );
  INV_X1 U405 ( .A(n4247), .ZN(n6680) );
  INV_X1 U406 ( .A(n4256), .ZN(n6679) );
  INV_X1 U407 ( .A(n4265), .ZN(n6678) );
  INV_X1 U408 ( .A(n4274), .ZN(n6677) );
  INV_X1 U409 ( .A(n4579), .ZN(n6638) );
  INV_X1 U410 ( .A(n4589), .ZN(n6637) );
  INV_X1 U411 ( .A(n4598), .ZN(n6636) );
  INV_X1 U412 ( .A(n4607), .ZN(n6635) );
  INV_X1 U413 ( .A(n4616), .ZN(n6634) );
  INV_X1 U414 ( .A(n4626), .ZN(n6633) );
  INV_X1 U415 ( .A(n4635), .ZN(n6632) );
  INV_X1 U416 ( .A(n4644), .ZN(n6631) );
  INV_X1 U417 ( .A(n4653), .ZN(n6630) );
  INV_X1 U418 ( .A(n2330), .ZN(n6643) );
  INV_X1 U419 ( .A(n2340), .ZN(n6642) );
  INV_X1 U420 ( .A(n2350), .ZN(n6641) );
  INV_X1 U421 ( .A(n2360), .ZN(n6640) );
  INV_X1 U422 ( .A(n2370), .ZN(n6639) );
  INV_X1 U423 ( .A(n2380), .ZN(n6884) );
  INV_X1 U424 ( .A(n2391), .ZN(n6883) );
  INV_X1 U425 ( .A(n2401), .ZN(n6882) );
  INV_X1 U426 ( .A(n2411), .ZN(n6881) );
  INV_X1 U427 ( .A(n2421), .ZN(n6880) );
  INV_X1 U428 ( .A(n2431), .ZN(n6879) );
  INV_X1 U429 ( .A(n2441), .ZN(n6878) );
  INV_X1 U430 ( .A(n2451), .ZN(n6877) );
  INV_X1 U431 ( .A(n2461), .ZN(n6876) );
  BUF_X1 U432 ( .A(n2069), .Z(n2063) );
  BUF_X1 U433 ( .A(n2069), .Z(n2062) );
  BUF_X1 U434 ( .A(n2069), .Z(n2064) );
  BUF_X1 U435 ( .A(n2068), .Z(n2060) );
  BUF_X1 U436 ( .A(n2068), .Z(n2058) );
  BUF_X1 U437 ( .A(n2068), .Z(n2061) );
  BUF_X1 U438 ( .A(n2068), .Z(n2059) );
  BUF_X1 U439 ( .A(n2135), .Z(n2095) );
  BUF_X1 U440 ( .A(n2135), .Z(n2094) );
  BUF_X1 U441 ( .A(N19), .Z(n2093) );
  BUF_X1 U442 ( .A(n2136), .Z(n2097) );
  BUF_X1 U443 ( .A(n2136), .Z(n2098) );
  BUF_X1 U444 ( .A(n2135), .Z(n2096) );
  BUF_X1 U445 ( .A(n2087), .Z(n2090) );
  BUF_X1 U446 ( .A(N20), .Z(n2089) );
  BUF_X1 U447 ( .A(n2136), .Z(n2099) );
  BUF_X1 U448 ( .A(n2136), .Z(n2092) );
  BUF_X1 U449 ( .A(N20), .Z(n2088) );
  BUF_X1 U450 ( .A(n2216), .Z(n2219) );
  BUF_X1 U451 ( .A(n2216), .Z(n2217) );
  NAND2_X1 U452 ( .A1(n2388), .A2(n2328), .ZN(n4579) );
  NAND2_X1 U453 ( .A1(n2399), .A2(n2328), .ZN(n4589) );
  NAND2_X1 U454 ( .A1(n2409), .A2(n2328), .ZN(n4598) );
  NAND2_X1 U455 ( .A1(n2419), .A2(n2328), .ZN(n4607) );
  NAND2_X1 U456 ( .A1(n2429), .A2(n2328), .ZN(n4616) );
  NAND2_X1 U457 ( .A1(n2439), .A2(n2328), .ZN(n4626) );
  NAND2_X1 U458 ( .A1(n2449), .A2(n2328), .ZN(n4635) );
  NAND2_X1 U459 ( .A1(n2459), .A2(n2328), .ZN(n4644) );
  NAND2_X1 U460 ( .A1(n2469), .A2(n2328), .ZN(n4653) );
  NAND2_X1 U461 ( .A1(n2338), .A2(n2328), .ZN(n2330) );
  NAND2_X1 U462 ( .A1(n2348), .A2(n2328), .ZN(n2340) );
  NAND2_X1 U463 ( .A1(n2358), .A2(n2328), .ZN(n2350) );
  NAND2_X1 U464 ( .A1(n2368), .A2(n2328), .ZN(n2360) );
  NAND2_X1 U465 ( .A1(n2378), .A2(n2328), .ZN(n2370) );
  NAND2_X1 U466 ( .A1(n2479), .A2(n2328), .ZN(n2314) );
  NAND2_X1 U467 ( .A1(n2327), .A2(n2328), .ZN(n2319) );
  NAND2_X1 U468 ( .A1(n2388), .A2(n2389), .ZN(n2380) );
  NAND2_X1 U469 ( .A1(n2399), .A2(n2389), .ZN(n2391) );
  NAND2_X1 U470 ( .A1(n2409), .A2(n2389), .ZN(n2401) );
  NAND2_X1 U471 ( .A1(n2419), .A2(n2389), .ZN(n2411) );
  NAND2_X1 U472 ( .A1(n2429), .A2(n2389), .ZN(n2421) );
  NAND2_X1 U473 ( .A1(n2439), .A2(n2389), .ZN(n2431) );
  NAND2_X1 U474 ( .A1(n2449), .A2(n2389), .ZN(n2441) );
  NAND2_X1 U475 ( .A1(n2459), .A2(n2389), .ZN(n2451) );
  NAND2_X1 U476 ( .A1(n2469), .A2(n2389), .ZN(n2461) );
  NAND2_X1 U477 ( .A1(n2545), .A2(n2388), .ZN(n2537) );
  NAND2_X1 U478 ( .A1(n2545), .A2(n2399), .ZN(n2547) );
  NAND2_X1 U479 ( .A1(n2545), .A2(n2409), .ZN(n2556) );
  NAND2_X1 U480 ( .A1(n2545), .A2(n2419), .ZN(n2565) );
  NAND2_X1 U481 ( .A1(n2545), .A2(n2429), .ZN(n2574) );
  NAND2_X1 U482 ( .A1(n2545), .A2(n2439), .ZN(n2583) );
  NAND2_X1 U483 ( .A1(n2545), .A2(n2449), .ZN(n2592) );
  NAND2_X1 U484 ( .A1(n2545), .A2(n2459), .ZN(n2601) );
  NAND2_X1 U485 ( .A1(n2545), .A2(n2469), .ZN(n2610) );
  NAND2_X1 U486 ( .A1(n2545), .A2(n2479), .ZN(n2619) );
  NAND2_X1 U487 ( .A1(n2545), .A2(n2327), .ZN(n2628) );
  NAND2_X1 U488 ( .A1(n2545), .A2(n2338), .ZN(n2637) );
  NAND2_X1 U489 ( .A1(n2545), .A2(n2348), .ZN(n2646) );
  NAND2_X1 U490 ( .A1(n2545), .A2(n2358), .ZN(n2655) );
  NAND2_X1 U491 ( .A1(n2545), .A2(n2368), .ZN(n2664) );
  NAND2_X1 U492 ( .A1(n2545), .A2(n2378), .ZN(n2673) );
  NAND2_X1 U493 ( .A1(n2692), .A2(n2388), .ZN(n2684) );
  NAND2_X1 U494 ( .A1(n2692), .A2(n2399), .ZN(n2694) );
  NAND2_X1 U496 ( .A1(n2692), .A2(n2409), .ZN(n2703) );
  NAND2_X1 U497 ( .A1(n2692), .A2(n2419), .ZN(n2712) );
  NAND2_X1 U498 ( .A1(n2692), .A2(n2429), .ZN(n2721) );
  NAND2_X1 U499 ( .A1(n2692), .A2(n2439), .ZN(n2730) );
  NAND2_X1 U500 ( .A1(n2692), .A2(n2449), .ZN(n2739) );
  NAND2_X1 U501 ( .A1(n2692), .A2(n2459), .ZN(n2748) );
  NAND2_X1 U502 ( .A1(n2692), .A2(n2469), .ZN(n2757) );
  NAND2_X1 U503 ( .A1(n2692), .A2(n2479), .ZN(n2766) );
  NAND2_X1 U504 ( .A1(n2692), .A2(n2327), .ZN(n2775) );
  NAND2_X1 U505 ( .A1(n2692), .A2(n2338), .ZN(n2784) );
  NAND2_X1 U506 ( .A1(n2692), .A2(n2348), .ZN(n2793) );
  NAND2_X1 U507 ( .A1(n2692), .A2(n2358), .ZN(n2802) );
  NAND2_X1 U508 ( .A1(n2692), .A2(n2368), .ZN(n2811) );
  NAND2_X1 U509 ( .A1(n2692), .A2(n2378), .ZN(n2820) );
  NAND2_X1 U510 ( .A1(n2838), .A2(n2388), .ZN(n2830) );
  NAND2_X1 U511 ( .A1(n2838), .A2(n2399), .ZN(n2840) );
  NAND2_X1 U512 ( .A1(n2838), .A2(n2409), .ZN(n2849) );
  NAND2_X1 U513 ( .A1(n2838), .A2(n2419), .ZN(n2858) );
  NAND2_X1 U514 ( .A1(n2838), .A2(n2429), .ZN(n2867) );
  NAND2_X1 U515 ( .A1(n2838), .A2(n2439), .ZN(n2876) );
  NAND2_X1 U516 ( .A1(n2838), .A2(n2449), .ZN(n2885) );
  NAND2_X1 U517 ( .A1(n2838), .A2(n2459), .ZN(n2894) );
  NAND2_X1 U518 ( .A1(n2838), .A2(n2469), .ZN(n2903) );
  NAND2_X1 U519 ( .A1(n2838), .A2(n2479), .ZN(n2912) );
  NAND2_X1 U520 ( .A1(n2838), .A2(n2327), .ZN(n2921) );
  NAND2_X1 U521 ( .A1(n2838), .A2(n2338), .ZN(n2930) );
  NAND2_X1 U522 ( .A1(n2838), .A2(n2348), .ZN(n2939) );
  NAND2_X1 U523 ( .A1(n2838), .A2(n2358), .ZN(n2948) );
  NAND2_X1 U524 ( .A1(n2838), .A2(n2368), .ZN(n2957) );
  NAND2_X1 U525 ( .A1(n2838), .A2(n2378), .ZN(n2966) );
  NAND2_X1 U526 ( .A1(n2984), .A2(n2388), .ZN(n2976) );
  NAND2_X1 U527 ( .A1(n2984), .A2(n2399), .ZN(n2986) );
  NAND2_X1 U528 ( .A1(n2984), .A2(n2409), .ZN(n2995) );
  NAND2_X1 U529 ( .A1(n2984), .A2(n2419), .ZN(n3004) );
  NAND2_X1 U530 ( .A1(n2984), .A2(n2429), .ZN(n3013) );
  NAND2_X1 U531 ( .A1(n2984), .A2(n2439), .ZN(n3022) );
  NAND2_X1 U532 ( .A1(n2984), .A2(n2449), .ZN(n3031) );
  NAND2_X1 U533 ( .A1(n2984), .A2(n2459), .ZN(n3040) );
  NAND2_X1 U534 ( .A1(n2984), .A2(n2469), .ZN(n3049) );
  NAND2_X1 U535 ( .A1(n2984), .A2(n2479), .ZN(n3058) );
  NAND2_X1 U536 ( .A1(n2984), .A2(n2327), .ZN(n3067) );
  NAND2_X1 U537 ( .A1(n2984), .A2(n2338), .ZN(n3076) );
  NAND2_X1 U538 ( .A1(n2984), .A2(n2348), .ZN(n3085) );
  NAND2_X1 U539 ( .A1(n2984), .A2(n2358), .ZN(n3094) );
  NAND2_X1 U540 ( .A1(n2984), .A2(n2368), .ZN(n3103) );
  NAND2_X1 U541 ( .A1(n2984), .A2(n2378), .ZN(n3112) );
  NAND2_X1 U542 ( .A1(n3129), .A2(n2388), .ZN(n3121) );
  NAND2_X1 U543 ( .A1(n3129), .A2(n2399), .ZN(n3131) );
  NAND2_X1 U544 ( .A1(n3129), .A2(n2409), .ZN(n3140) );
  NAND2_X1 U545 ( .A1(n3129), .A2(n2419), .ZN(n3149) );
  NAND2_X1 U546 ( .A1(n3129), .A2(n2429), .ZN(n3158) );
  NAND2_X1 U547 ( .A1(n3129), .A2(n2439), .ZN(n3167) );
  NAND2_X1 U548 ( .A1(n3129), .A2(n2449), .ZN(n3176) );
  NAND2_X1 U549 ( .A1(n3129), .A2(n2459), .ZN(n3185) );
  NAND2_X1 U550 ( .A1(n3129), .A2(n2469), .ZN(n3194) );
  NAND2_X1 U551 ( .A1(n3129), .A2(n2479), .ZN(n3203) );
  NAND2_X1 U552 ( .A1(n3129), .A2(n2327), .ZN(n3212) );
  NAND2_X1 U553 ( .A1(n3129), .A2(n2338), .ZN(n3221) );
  NAND2_X1 U554 ( .A1(n3129), .A2(n2348), .ZN(n3230) );
  NAND2_X1 U555 ( .A1(n3129), .A2(n2358), .ZN(n3239) );
  NAND2_X1 U556 ( .A1(n3129), .A2(n2368), .ZN(n3248) );
  NAND2_X1 U557 ( .A1(n3129), .A2(n2378), .ZN(n3257) );
  NAND2_X1 U558 ( .A1(n3275), .A2(n2388), .ZN(n3267) );
  NAND2_X1 U559 ( .A1(n3275), .A2(n2399), .ZN(n3277) );
  NAND2_X1 U560 ( .A1(n3275), .A2(n2409), .ZN(n3286) );
  NAND2_X1 U561 ( .A1(n3275), .A2(n2419), .ZN(n3295) );
  NAND2_X1 U562 ( .A1(n3275), .A2(n2429), .ZN(n3304) );
  NAND2_X1 U563 ( .A1(n3275), .A2(n2439), .ZN(n3313) );
  NAND2_X1 U564 ( .A1(n3275), .A2(n2449), .ZN(n3322) );
  NAND2_X1 U565 ( .A1(n3275), .A2(n2459), .ZN(n3331) );
  NAND2_X1 U566 ( .A1(n3275), .A2(n2469), .ZN(n3340) );
  NAND2_X1 U567 ( .A1(n3275), .A2(n2479), .ZN(n3349) );
  NAND2_X1 U568 ( .A1(n3275), .A2(n2327), .ZN(n3358) );
  NAND2_X1 U569 ( .A1(n3275), .A2(n2338), .ZN(n3367) );
  NAND2_X1 U570 ( .A1(n3275), .A2(n2348), .ZN(n3376) );
  NAND2_X1 U571 ( .A1(n3275), .A2(n2358), .ZN(n3385) );
  NAND2_X1 U572 ( .A1(n3275), .A2(n2368), .ZN(n3394) );
  NAND2_X1 U573 ( .A1(n3275), .A2(n2378), .ZN(n3403) );
  NAND2_X1 U574 ( .A1(n3420), .A2(n2388), .ZN(n3412) );
  NAND2_X1 U575 ( .A1(n3420), .A2(n2399), .ZN(n3422) );
  NAND2_X1 U576 ( .A1(n3420), .A2(n2409), .ZN(n3431) );
  NAND2_X1 U577 ( .A1(n3420), .A2(n2419), .ZN(n3440) );
  NAND2_X1 U578 ( .A1(n3420), .A2(n2429), .ZN(n3449) );
  NAND2_X1 U579 ( .A1(n3420), .A2(n2439), .ZN(n3458) );
  NAND2_X1 U580 ( .A1(n3420), .A2(n2449), .ZN(n3467) );
  NAND2_X1 U581 ( .A1(n3420), .A2(n2459), .ZN(n3476) );
  NAND2_X1 U582 ( .A1(n3420), .A2(n2469), .ZN(n3485) );
  NAND2_X1 U583 ( .A1(n3420), .A2(n2479), .ZN(n3494) );
  NAND2_X1 U584 ( .A1(n3420), .A2(n2327), .ZN(n3503) );
  NAND2_X1 U585 ( .A1(n3420), .A2(n2338), .ZN(n3512) );
  NAND2_X1 U586 ( .A1(n3420), .A2(n2348), .ZN(n3521) );
  NAND2_X1 U587 ( .A1(n3420), .A2(n2358), .ZN(n3530) );
  NAND2_X1 U588 ( .A1(n3420), .A2(n2368), .ZN(n3539) );
  NAND2_X1 U589 ( .A1(n3420), .A2(n2378), .ZN(n3548) );
  NAND2_X1 U590 ( .A1(n3565), .A2(n2388), .ZN(n3557) );
  NAND2_X1 U591 ( .A1(n3565), .A2(n2399), .ZN(n3567) );
  NAND2_X1 U592 ( .A1(n3565), .A2(n2409), .ZN(n3576) );
  NAND2_X1 U593 ( .A1(n3565), .A2(n2419), .ZN(n3585) );
  NAND2_X1 U594 ( .A1(n3565), .A2(n2429), .ZN(n3594) );
  NAND2_X1 U595 ( .A1(n3565), .A2(n2439), .ZN(n3603) );
  NAND2_X1 U596 ( .A1(n3565), .A2(n2449), .ZN(n3612) );
  NAND2_X1 U597 ( .A1(n3565), .A2(n2459), .ZN(n3621) );
  NAND2_X1 U598 ( .A1(n3565), .A2(n2469), .ZN(n3630) );
  NAND2_X1 U599 ( .A1(n3565), .A2(n2479), .ZN(n3639) );
  NAND2_X1 U600 ( .A1(n3565), .A2(n2327), .ZN(n3648) );
  NAND2_X1 U601 ( .A1(n3565), .A2(n2338), .ZN(n3657) );
  NAND2_X1 U602 ( .A1(n3565), .A2(n2348), .ZN(n3666) );
  NAND2_X1 U603 ( .A1(n3565), .A2(n2358), .ZN(n3675) );
  NAND2_X1 U604 ( .A1(n3565), .A2(n2368), .ZN(n3684) );
  NAND2_X1 U605 ( .A1(n3565), .A2(n2378), .ZN(n3693) );
  NAND2_X1 U606 ( .A1(n3710), .A2(n2388), .ZN(n3702) );
  NAND2_X1 U607 ( .A1(n3710), .A2(n2399), .ZN(n3712) );
  NAND2_X1 U608 ( .A1(n3710), .A2(n2409), .ZN(n3721) );
  NAND2_X1 U609 ( .A1(n3710), .A2(n2419), .ZN(n3730) );
  NAND2_X1 U610 ( .A1(n3710), .A2(n2429), .ZN(n3739) );
  NAND2_X1 U611 ( .A1(n3710), .A2(n2439), .ZN(n3748) );
  NAND2_X1 U612 ( .A1(n3710), .A2(n2449), .ZN(n3757) );
  NAND2_X1 U613 ( .A1(n3710), .A2(n2459), .ZN(n3766) );
  NAND2_X1 U614 ( .A1(n3710), .A2(n2469), .ZN(n3775) );
  NAND2_X1 U615 ( .A1(n3710), .A2(n2479), .ZN(n3784) );
  NAND2_X1 U616 ( .A1(n3710), .A2(n2327), .ZN(n3793) );
  NAND2_X1 U617 ( .A1(n3710), .A2(n2338), .ZN(n3802) );
  NAND2_X1 U618 ( .A1(n3710), .A2(n2348), .ZN(n3811) );
  NAND2_X1 U619 ( .A1(n3710), .A2(n2358), .ZN(n3820) );
  NAND2_X1 U620 ( .A1(n3710), .A2(n2368), .ZN(n3829) );
  NAND2_X1 U621 ( .A1(n3710), .A2(n2378), .ZN(n3838) );
  NAND2_X1 U622 ( .A1(n3856), .A2(n2388), .ZN(n3848) );
  NAND2_X1 U623 ( .A1(n3856), .A2(n2399), .ZN(n3858) );
  NAND2_X1 U624 ( .A1(n3856), .A2(n2409), .ZN(n3867) );
  NAND2_X1 U625 ( .A1(n3856), .A2(n2419), .ZN(n3876) );
  NAND2_X1 U626 ( .A1(n3856), .A2(n2429), .ZN(n3885) );
  NAND2_X1 U627 ( .A1(n3856), .A2(n2439), .ZN(n3894) );
  NAND2_X1 U628 ( .A1(n3856), .A2(n2449), .ZN(n3903) );
  NAND2_X1 U629 ( .A1(n3856), .A2(n2459), .ZN(n3912) );
  NAND2_X1 U630 ( .A1(n3856), .A2(n2469), .ZN(n3921) );
  NAND2_X1 U631 ( .A1(n3856), .A2(n2479), .ZN(n3930) );
  NAND2_X1 U632 ( .A1(n3856), .A2(n2327), .ZN(n3939) );
  NAND2_X1 U633 ( .A1(n3856), .A2(n2338), .ZN(n3948) );
  NAND2_X1 U634 ( .A1(n3856), .A2(n2348), .ZN(n3957) );
  NAND2_X1 U635 ( .A1(n3856), .A2(n2358), .ZN(n3966) );
  NAND2_X1 U636 ( .A1(n3856), .A2(n2368), .ZN(n3975) );
  NAND2_X1 U637 ( .A1(n3856), .A2(n2378), .ZN(n3984) );
  NAND2_X1 U638 ( .A1(n4001), .A2(n2388), .ZN(n3993) );
  NAND2_X1 U639 ( .A1(n4001), .A2(n2399), .ZN(n4003) );
  NAND2_X1 U641 ( .A1(n4001), .A2(n2409), .ZN(n4012) );
  NAND2_X1 U642 ( .A1(n4001), .A2(n2419), .ZN(n4021) );
  NAND2_X1 U643 ( .A1(n4001), .A2(n2429), .ZN(n4030) );
  NAND2_X1 U644 ( .A1(n4001), .A2(n2439), .ZN(n4039) );
  NAND2_X1 U645 ( .A1(n4001), .A2(n2449), .ZN(n4048) );
  NAND2_X1 U646 ( .A1(n4001), .A2(n2459), .ZN(n4057) );
  NAND2_X1 U647 ( .A1(n4001), .A2(n2469), .ZN(n4066) );
  NAND2_X1 U648 ( .A1(n4001), .A2(n2479), .ZN(n4075) );
  NAND2_X1 U649 ( .A1(n4001), .A2(n2327), .ZN(n4084) );
  NAND2_X1 U650 ( .A1(n4001), .A2(n2338), .ZN(n4093) );
  NAND2_X1 U651 ( .A1(n4001), .A2(n2348), .ZN(n4102) );
  NAND2_X1 U652 ( .A1(n4001), .A2(n2358), .ZN(n4111) );
  NAND2_X1 U653 ( .A1(n4001), .A2(n2368), .ZN(n4120) );
  NAND2_X1 U654 ( .A1(n4001), .A2(n2378), .ZN(n4129) );
  NAND2_X1 U655 ( .A1(n4146), .A2(n2388), .ZN(n4138) );
  NAND2_X1 U656 ( .A1(n4146), .A2(n2399), .ZN(n4148) );
  NAND2_X1 U657 ( .A1(n4146), .A2(n2409), .ZN(n4157) );
  NAND2_X1 U658 ( .A1(n4146), .A2(n2419), .ZN(n4166) );
  NAND2_X1 U659 ( .A1(n4146), .A2(n2429), .ZN(n4175) );
  NAND2_X1 U660 ( .A1(n4146), .A2(n2439), .ZN(n4184) );
  NAND2_X1 U661 ( .A1(n4146), .A2(n2449), .ZN(n4193) );
  NAND2_X1 U662 ( .A1(n4146), .A2(n2459), .ZN(n4202) );
  NAND2_X1 U663 ( .A1(n4146), .A2(n2469), .ZN(n4211) );
  NAND2_X1 U664 ( .A1(n4146), .A2(n2479), .ZN(n4220) );
  NAND2_X1 U665 ( .A1(n4146), .A2(n2327), .ZN(n4229) );
  NAND2_X1 U666 ( .A1(n4146), .A2(n2338), .ZN(n4238) );
  NAND2_X1 U667 ( .A1(n4146), .A2(n2348), .ZN(n4247) );
  NAND2_X1 U668 ( .A1(n4146), .A2(n2358), .ZN(n4256) );
  NAND2_X1 U669 ( .A1(n4146), .A2(n2368), .ZN(n4265) );
  NAND2_X1 U670 ( .A1(n4146), .A2(n2378), .ZN(n4274) );
  NAND2_X1 U671 ( .A1(n4291), .A2(n2388), .ZN(n4283) );
  NAND2_X1 U672 ( .A1(n4291), .A2(n2399), .ZN(n4293) );
  NAND2_X1 U673 ( .A1(n4291), .A2(n2409), .ZN(n4302) );
  NAND2_X1 U674 ( .A1(n4291), .A2(n2419), .ZN(n4311) );
  NAND2_X1 U675 ( .A1(n4291), .A2(n2429), .ZN(n4320) );
  NAND2_X1 U676 ( .A1(n4291), .A2(n2439), .ZN(n4329) );
  NAND2_X1 U677 ( .A1(n4291), .A2(n2449), .ZN(n4338) );
  NAND2_X1 U678 ( .A1(n4291), .A2(n2459), .ZN(n4347) );
  NAND2_X1 U679 ( .A1(n4291), .A2(n2469), .ZN(n4356) );
  NAND2_X1 U680 ( .A1(n4291), .A2(n2479), .ZN(n4365) );
  NAND2_X1 U681 ( .A1(n4291), .A2(n2327), .ZN(n4374) );
  NAND2_X1 U682 ( .A1(n4291), .A2(n2338), .ZN(n4383) );
  NAND2_X1 U683 ( .A1(n4291), .A2(n2348), .ZN(n4392) );
  NAND2_X1 U684 ( .A1(n4291), .A2(n2358), .ZN(n4401) );
  NAND2_X1 U685 ( .A1(n4291), .A2(n2368), .ZN(n4410) );
  NAND2_X1 U686 ( .A1(n4291), .A2(n2378), .ZN(n4419) );
  NAND2_X1 U687 ( .A1(n4436), .A2(n2388), .ZN(n4428) );
  NAND2_X1 U688 ( .A1(n4436), .A2(n2399), .ZN(n4438) );
  NAND2_X1 U689 ( .A1(n4436), .A2(n2409), .ZN(n4447) );
  NAND2_X1 U690 ( .A1(n4436), .A2(n2419), .ZN(n4456) );
  NAND2_X1 U691 ( .A1(n4436), .A2(n2429), .ZN(n4465) );
  NAND2_X1 U692 ( .A1(n4436), .A2(n2439), .ZN(n4474) );
  NAND2_X1 U693 ( .A1(n4436), .A2(n2449), .ZN(n4483) );
  NAND2_X1 U694 ( .A1(n4436), .A2(n2459), .ZN(n4492) );
  NAND2_X1 U695 ( .A1(n4436), .A2(n2469), .ZN(n4501) );
  NAND2_X1 U696 ( .A1(n4436), .A2(n2479), .ZN(n4510) );
  NAND2_X1 U697 ( .A1(n4436), .A2(n2327), .ZN(n4519) );
  NAND2_X1 U698 ( .A1(n4436), .A2(n2338), .ZN(n4530) );
  NAND2_X1 U699 ( .A1(n4436), .A2(n2348), .ZN(n4540) );
  NAND2_X1 U700 ( .A1(n4436), .A2(n2358), .ZN(n4551) );
  NAND2_X1 U701 ( .A1(n4436), .A2(n2368), .ZN(n4561) );
  NAND2_X1 U702 ( .A1(n4436), .A2(n2378), .ZN(n4570) );
  NAND2_X1 U703 ( .A1(n2389), .A2(n2479), .ZN(n2471) );
  NAND2_X1 U704 ( .A1(n2389), .A2(n2327), .ZN(n2481) );
  NAND2_X1 U705 ( .A1(n2389), .A2(n2338), .ZN(n2490) );
  NAND2_X1 U706 ( .A1(n2389), .A2(n2348), .ZN(n2499) );
  NAND2_X1 U707 ( .A1(n2389), .A2(n2358), .ZN(n2508) );
  NAND2_X1 U708 ( .A1(n2389), .A2(n2368), .ZN(n2517) );
  NAND2_X1 U709 ( .A1(n2389), .A2(n2378), .ZN(n2526) );
  NOR2_X1 U710 ( .A1(N20), .A2(N21), .ZN(n4587) );
  NOR2_X1 U711 ( .A1(N22), .A2(N23), .ZN(n2681) );
  BUF_X1 U712 ( .A(N22), .Z(n2052) );
  BUF_X1 U713 ( .A(N22), .Z(n2053) );
  BUF_X1 U714 ( .A(N22), .Z(n2054) );
  BUF_X1 U715 ( .A(N22), .Z(n2055) );
  BUF_X1 U716 ( .A(N22), .Z(n2056) );
  BUF_X1 U717 ( .A(N23), .Z(n2049) );
  BUF_X1 U718 ( .A(N23), .Z(n2050) );
  BUF_X1 U719 ( .A(N23), .Z(n2048) );
  BUF_X1 U720 ( .A(N21), .Z(n2069) );
  BUF_X1 U721 ( .A(N19), .Z(n2135) );
  BUF_X1 U722 ( .A(N19), .Z(n2136) );
  BUF_X1 U723 ( .A(N20), .Z(n2087) );
  NOR2_X1 U724 ( .A1(n2), .A2(N19), .ZN(n4559) );
  NOR2_X1 U725 ( .A1(n2226), .A2(N20), .ZN(n4528) );
  NOR2_X1 U726 ( .A1(n2224), .A2(n2), .ZN(n4538) );
  NOR2_X1 U727 ( .A1(n2225), .A2(N21), .ZN(n4624) );
  NOR2_X1 U728 ( .A1(n2225), .A2(n2226), .ZN(n4548) );
  NOR2_X1 U729 ( .A1(n11), .A2(n6885), .ZN(n2534) );
  NOR2_X1 U730 ( .A1(n2228), .A2(N22), .ZN(n2974) );
  NOR2_X1 U731 ( .A1(n2227), .A2(N23), .ZN(n2828) );
  NOR2_X1 U732 ( .A1(n2227), .A2(n2228), .ZN(n2535) );
  NOR2_X1 U733 ( .A1(N24), .A2(N25), .ZN(n2682) );
  NOR2_X1 U734 ( .A1(n11), .A2(N24), .ZN(n3846) );
  INV_X1 U735 ( .A(N24), .ZN(n6885) );
  INV_X1 U736 ( .A(N23), .ZN(n2228) );
  INV_X1 U737 ( .A(N21), .ZN(n2226) );
  INV_X1 U738 ( .A(N20), .ZN(n2225) );
  INV_X1 U739 ( .A(N22), .ZN(n2227) );
  INV_X1 U740 ( .A(N19), .ZN(n2224) );
  INV_X1 U741 ( .A(n2323), .ZN(n4752) );
  AOI22_X1 U742 ( .A1(\mem[234][4] ), .A2(n2319), .B1(n6644), .B2(data_in[4]), 
        .ZN(n2323) );
  INV_X1 U743 ( .A(n2324), .ZN(n4751) );
  AOI22_X1 U744 ( .A1(\mem[234][5] ), .A2(n2319), .B1(n6644), .B2(data_in[5]), 
        .ZN(n2324) );
  INV_X1 U745 ( .A(n2325), .ZN(n4750) );
  AOI22_X1 U746 ( .A1(\mem[234][6] ), .A2(n2319), .B1(n6644), .B2(data_in[6]), 
        .ZN(n2325) );
  INV_X1 U747 ( .A(n2326), .ZN(n4749) );
  AOI22_X1 U748 ( .A1(\mem[234][7] ), .A2(n2319), .B1(n6644), .B2(data_in[7]), 
        .ZN(n2326) );
  INV_X1 U749 ( .A(n2313), .ZN(n4760) );
  AOI22_X1 U750 ( .A1(\mem[233][4] ), .A2(n2314), .B1(data_in[4]), .B2(n6629), 
        .ZN(n2313) );
  INV_X1 U751 ( .A(n2315), .ZN(n4759) );
  AOI22_X1 U752 ( .A1(\mem[233][5] ), .A2(n2314), .B1(data_in[5]), .B2(n6629), 
        .ZN(n2315) );
  INV_X1 U753 ( .A(n2316), .ZN(n4758) );
  AOI22_X1 U754 ( .A1(\mem[233][6] ), .A2(n2314), .B1(data_in[6]), .B2(n6629), 
        .ZN(n2316) );
  INV_X1 U755 ( .A(n2317), .ZN(n4757) );
  AOI22_X1 U756 ( .A1(\mem[233][7] ), .A2(n2314), .B1(data_in[7]), .B2(n6629), 
        .ZN(n2317) );
  INV_X1 U757 ( .A(n4661), .ZN(n4764) );
  AOI22_X1 U758 ( .A1(\mem[233][0] ), .A2(n2314), .B1(data_in[0]), .B2(n6629), 
        .ZN(n4661) );
  INV_X1 U759 ( .A(n4662), .ZN(n4763) );
  AOI22_X1 U760 ( .A1(\mem[233][1] ), .A2(n2314), .B1(data_in[1]), .B2(n6629), 
        .ZN(n4662) );
  INV_X1 U761 ( .A(n4663), .ZN(n4762) );
  AOI22_X1 U762 ( .A1(\mem[233][2] ), .A2(n2314), .B1(data_in[2]), .B2(n6629), 
        .ZN(n4663) );
  INV_X1 U763 ( .A(n4664), .ZN(n4761) );
  AOI22_X1 U764 ( .A1(\mem[233][3] ), .A2(n2314), .B1(data_in[3]), .B2(n6629), 
        .ZN(n4664) );
  INV_X1 U765 ( .A(n2318), .ZN(n4756) );
  AOI22_X1 U766 ( .A1(\mem[234][0] ), .A2(n2319), .B1(data_in[0]), .B2(n6644), 
        .ZN(n2318) );
  INV_X1 U767 ( .A(n2320), .ZN(n4755) );
  AOI22_X1 U768 ( .A1(\mem[234][1] ), .A2(n2319), .B1(data_in[1]), .B2(n6644), 
        .ZN(n2320) );
  INV_X1 U769 ( .A(n2321), .ZN(n4754) );
  AOI22_X1 U770 ( .A1(\mem[234][2] ), .A2(n2319), .B1(data_in[2]), .B2(n6644), 
        .ZN(n2321) );
  INV_X1 U771 ( .A(n2322), .ZN(n4753) );
  AOI22_X1 U772 ( .A1(\mem[234][3] ), .A2(n2319), .B1(data_in[3]), .B2(n6644), 
        .ZN(n2322) );
  INV_X1 U773 ( .A(n2470), .ZN(n2284) );
  AOI22_X1 U774 ( .A1(\mem[249][0] ), .A2(n2471), .B1(n6875), .B2(data_in[0]), 
        .ZN(n2470) );
  INV_X1 U775 ( .A(n2472), .ZN(n2283) );
  AOI22_X1 U776 ( .A1(\mem[249][1] ), .A2(n2471), .B1(n6875), .B2(data_in[1]), 
        .ZN(n2472) );
  INV_X1 U777 ( .A(n2473), .ZN(n2282) );
  AOI22_X1 U778 ( .A1(\mem[249][2] ), .A2(n2471), .B1(n6875), .B2(data_in[2]), 
        .ZN(n2473) );
  INV_X1 U779 ( .A(n2474), .ZN(n2281) );
  AOI22_X1 U780 ( .A1(\mem[249][3] ), .A2(n2471), .B1(n6875), .B2(data_in[3]), 
        .ZN(n2474) );
  INV_X1 U781 ( .A(n2475), .ZN(n2280) );
  AOI22_X1 U782 ( .A1(\mem[249][4] ), .A2(n2471), .B1(n6875), .B2(data_in[4]), 
        .ZN(n2475) );
  INV_X1 U783 ( .A(n2476), .ZN(n2279) );
  AOI22_X1 U784 ( .A1(\mem[249][5] ), .A2(n2471), .B1(n6875), .B2(data_in[5]), 
        .ZN(n2476) );
  INV_X1 U786 ( .A(n2477), .ZN(n2278) );
  AOI22_X1 U787 ( .A1(\mem[249][6] ), .A2(n2471), .B1(n6875), .B2(data_in[6]), 
        .ZN(n2477) );
  INV_X1 U788 ( .A(n2478), .ZN(n2277) );
  AOI22_X1 U789 ( .A1(\mem[249][7] ), .A2(n2471), .B1(n6875), .B2(data_in[7]), 
        .ZN(n2478) );
  INV_X1 U790 ( .A(n2480), .ZN(n2276) );
  AOI22_X1 U791 ( .A1(\mem[250][0] ), .A2(n2481), .B1(n6874), .B2(data_in[0]), 
        .ZN(n2480) );
  INV_X1 U792 ( .A(n2482), .ZN(n2275) );
  AOI22_X1 U793 ( .A1(\mem[250][1] ), .A2(n2481), .B1(n6874), .B2(data_in[1]), 
        .ZN(n2482) );
  INV_X1 U794 ( .A(n2483), .ZN(n2274) );
  AOI22_X1 U795 ( .A1(\mem[250][2] ), .A2(n2481), .B1(n6874), .B2(data_in[2]), 
        .ZN(n2483) );
  INV_X1 U796 ( .A(n2484), .ZN(n2273) );
  AOI22_X1 U797 ( .A1(\mem[250][3] ), .A2(n2481), .B1(n6874), .B2(data_in[3]), 
        .ZN(n2484) );
  INV_X1 U798 ( .A(n2485), .ZN(n2272) );
  AOI22_X1 U799 ( .A1(\mem[250][4] ), .A2(n2481), .B1(n6874), .B2(data_in[4]), 
        .ZN(n2485) );
  INV_X1 U800 ( .A(n2486), .ZN(n2271) );
  AOI22_X1 U801 ( .A1(\mem[250][5] ), .A2(n2481), .B1(n6874), .B2(data_in[5]), 
        .ZN(n2486) );
  INV_X1 U802 ( .A(n2487), .ZN(n2270) );
  AOI22_X1 U803 ( .A1(\mem[250][6] ), .A2(n2481), .B1(n6874), .B2(data_in[6]), 
        .ZN(n2487) );
  INV_X1 U804 ( .A(n2488), .ZN(n2269) );
  AOI22_X1 U805 ( .A1(\mem[250][7] ), .A2(n2481), .B1(n6874), .B2(data_in[7]), 
        .ZN(n2488) );
  INV_X1 U806 ( .A(n2489), .ZN(n2268) );
  AOI22_X1 U807 ( .A1(\mem[251][0] ), .A2(n2490), .B1(n6873), .B2(data_in[0]), 
        .ZN(n2489) );
  INV_X1 U808 ( .A(n2491), .ZN(n2267) );
  AOI22_X1 U809 ( .A1(\mem[251][1] ), .A2(n2490), .B1(n6873), .B2(data_in[1]), 
        .ZN(n2491) );
  INV_X1 U810 ( .A(n2492), .ZN(n2266) );
  AOI22_X1 U811 ( .A1(\mem[251][2] ), .A2(n2490), .B1(n6873), .B2(data_in[2]), 
        .ZN(n2492) );
  INV_X1 U812 ( .A(n2493), .ZN(n2265) );
  AOI22_X1 U813 ( .A1(\mem[251][3] ), .A2(n2490), .B1(n6873), .B2(data_in[3]), 
        .ZN(n2493) );
  INV_X1 U814 ( .A(n2494), .ZN(n2264) );
  AOI22_X1 U815 ( .A1(\mem[251][4] ), .A2(n2490), .B1(n6873), .B2(data_in[4]), 
        .ZN(n2494) );
  INV_X1 U816 ( .A(n2495), .ZN(n2263) );
  AOI22_X1 U817 ( .A1(\mem[251][5] ), .A2(n2490), .B1(n6873), .B2(data_in[5]), 
        .ZN(n2495) );
  INV_X1 U818 ( .A(n2496), .ZN(n2262) );
  AOI22_X1 U819 ( .A1(\mem[251][6] ), .A2(n2490), .B1(n6873), .B2(data_in[6]), 
        .ZN(n2496) );
  INV_X1 U820 ( .A(n2497), .ZN(n2261) );
  AOI22_X1 U821 ( .A1(\mem[251][7] ), .A2(n2490), .B1(n6873), .B2(data_in[7]), 
        .ZN(n2497) );
  INV_X1 U822 ( .A(n2498), .ZN(n2260) );
  AOI22_X1 U823 ( .A1(\mem[252][0] ), .A2(n2499), .B1(n6872), .B2(data_in[0]), 
        .ZN(n2498) );
  INV_X1 U824 ( .A(n2500), .ZN(n2259) );
  AOI22_X1 U825 ( .A1(\mem[252][1] ), .A2(n2499), .B1(n6872), .B2(data_in[1]), 
        .ZN(n2500) );
  INV_X1 U826 ( .A(n2501), .ZN(n2258) );
  AOI22_X1 U827 ( .A1(\mem[252][2] ), .A2(n2499), .B1(n6872), .B2(data_in[2]), 
        .ZN(n2501) );
  INV_X1 U828 ( .A(n2502), .ZN(n2257) );
  AOI22_X1 U829 ( .A1(\mem[252][3] ), .A2(n2499), .B1(n6872), .B2(data_in[3]), 
        .ZN(n2502) );
  INV_X1 U830 ( .A(n2503), .ZN(n2256) );
  AOI22_X1 U831 ( .A1(\mem[252][4] ), .A2(n2499), .B1(n6872), .B2(data_in[4]), 
        .ZN(n2503) );
  INV_X1 U832 ( .A(n2504), .ZN(n2255) );
  AOI22_X1 U833 ( .A1(\mem[252][5] ), .A2(n2499), .B1(n6872), .B2(data_in[5]), 
        .ZN(n2504) );
  INV_X1 U834 ( .A(n2505), .ZN(n2254) );
  AOI22_X1 U835 ( .A1(\mem[252][6] ), .A2(n2499), .B1(n6872), .B2(data_in[6]), 
        .ZN(n2505) );
  INV_X1 U836 ( .A(n2506), .ZN(n2253) );
  AOI22_X1 U837 ( .A1(\mem[252][7] ), .A2(n2499), .B1(n6872), .B2(data_in[7]), 
        .ZN(n2506) );
  INV_X1 U838 ( .A(n2507), .ZN(n2252) );
  AOI22_X1 U839 ( .A1(\mem[253][0] ), .A2(n2508), .B1(n6871), .B2(data_in[0]), 
        .ZN(n2507) );
  INV_X1 U840 ( .A(n2509), .ZN(n2251) );
  AOI22_X1 U841 ( .A1(\mem[253][1] ), .A2(n2508), .B1(n6871), .B2(data_in[1]), 
        .ZN(n2509) );
  INV_X1 U842 ( .A(n2510), .ZN(n2250) );
  AOI22_X1 U843 ( .A1(\mem[253][2] ), .A2(n2508), .B1(n6871), .B2(data_in[2]), 
        .ZN(n2510) );
  INV_X1 U844 ( .A(n2511), .ZN(n2249) );
  AOI22_X1 U845 ( .A1(\mem[253][3] ), .A2(n2508), .B1(n6871), .B2(data_in[3]), 
        .ZN(n2511) );
  INV_X1 U846 ( .A(n2512), .ZN(n2248) );
  AOI22_X1 U847 ( .A1(\mem[253][4] ), .A2(n2508), .B1(n6871), .B2(data_in[4]), 
        .ZN(n2512) );
  INV_X1 U848 ( .A(n2513), .ZN(n2247) );
  AOI22_X1 U849 ( .A1(\mem[253][5] ), .A2(n2508), .B1(n6871), .B2(data_in[5]), 
        .ZN(n2513) );
  INV_X1 U850 ( .A(n2514), .ZN(n2246) );
  AOI22_X1 U851 ( .A1(\mem[253][6] ), .A2(n2508), .B1(n6871), .B2(data_in[6]), 
        .ZN(n2514) );
  INV_X1 U852 ( .A(n2515), .ZN(n2245) );
  AOI22_X1 U853 ( .A1(\mem[253][7] ), .A2(n2508), .B1(n6871), .B2(data_in[7]), 
        .ZN(n2515) );
  INV_X1 U854 ( .A(n2516), .ZN(n2244) );
  AOI22_X1 U855 ( .A1(\mem[254][0] ), .A2(n2517), .B1(n6870), .B2(data_in[0]), 
        .ZN(n2516) );
  INV_X1 U856 ( .A(n2518), .ZN(n2243) );
  AOI22_X1 U857 ( .A1(\mem[254][1] ), .A2(n2517), .B1(n6870), .B2(data_in[1]), 
        .ZN(n2518) );
  INV_X1 U858 ( .A(n2519), .ZN(n2242) );
  AOI22_X1 U859 ( .A1(\mem[254][2] ), .A2(n2517), .B1(n6870), .B2(data_in[2]), 
        .ZN(n2519) );
  INV_X1 U860 ( .A(n2520), .ZN(n2241) );
  AOI22_X1 U861 ( .A1(\mem[254][3] ), .A2(n2517), .B1(n6870), .B2(data_in[3]), 
        .ZN(n2520) );
  INV_X1 U862 ( .A(n2521), .ZN(n2240) );
  AOI22_X1 U863 ( .A1(\mem[254][4] ), .A2(n2517), .B1(n6870), .B2(data_in[4]), 
        .ZN(n2521) );
  INV_X1 U864 ( .A(n2522), .ZN(n2239) );
  AOI22_X1 U865 ( .A1(\mem[254][5] ), .A2(n2517), .B1(n6870), .B2(data_in[5]), 
        .ZN(n2522) );
  INV_X1 U866 ( .A(n2523), .ZN(n2238) );
  AOI22_X1 U867 ( .A1(\mem[254][6] ), .A2(n2517), .B1(n6870), .B2(data_in[6]), 
        .ZN(n2523) );
  INV_X1 U868 ( .A(n2524), .ZN(n2237) );
  AOI22_X1 U869 ( .A1(\mem[254][7] ), .A2(n2517), .B1(n6870), .B2(data_in[7]), 
        .ZN(n2524) );
  INV_X1 U870 ( .A(n2525), .ZN(n2236) );
  AOI22_X1 U871 ( .A1(\mem[255][0] ), .A2(n2526), .B1(n6869), .B2(data_in[0]), 
        .ZN(n2525) );
  INV_X1 U872 ( .A(n2527), .ZN(n2235) );
  AOI22_X1 U873 ( .A1(\mem[255][1] ), .A2(n2526), .B1(n6869), .B2(data_in[1]), 
        .ZN(n2527) );
  INV_X1 U874 ( .A(n2528), .ZN(n2234) );
  AOI22_X1 U875 ( .A1(\mem[255][2] ), .A2(n2526), .B1(n6869), .B2(data_in[2]), 
        .ZN(n2528) );
  INV_X1 U876 ( .A(n2529), .ZN(n2233) );
  AOI22_X1 U877 ( .A1(\mem[255][3] ), .A2(n2526), .B1(n6869), .B2(data_in[3]), 
        .ZN(n2529) );
  INV_X1 U878 ( .A(n2530), .ZN(n2232) );
  AOI22_X1 U879 ( .A1(\mem[255][4] ), .A2(n2526), .B1(n6869), .B2(data_in[4]), 
        .ZN(n2530) );
  INV_X1 U880 ( .A(n2531), .ZN(n2231) );
  AOI22_X1 U881 ( .A1(\mem[255][5] ), .A2(n2526), .B1(n6869), .B2(data_in[5]), 
        .ZN(n2531) );
  INV_X1 U882 ( .A(n2532), .ZN(n2230) );
  AOI22_X1 U883 ( .A1(\mem[255][6] ), .A2(n2526), .B1(n6869), .B2(data_in[6]), 
        .ZN(n2532) );
  INV_X1 U884 ( .A(n2533), .ZN(n2229) );
  AOI22_X1 U885 ( .A1(\mem[255][7] ), .A2(n2526), .B1(n6869), .B2(data_in[7]), 
        .ZN(n2533) );
  INV_X1 U886 ( .A(n2536), .ZN(n6628) );
  AOI22_X1 U887 ( .A1(\mem[0][0] ), .A2(n2537), .B1(n6868), .B2(data_in[0]), 
        .ZN(n2536) );
  INV_X1 U888 ( .A(n2538), .ZN(n6627) );
  AOI22_X1 U889 ( .A1(\mem[0][1] ), .A2(n2537), .B1(n6868), .B2(data_in[1]), 
        .ZN(n2538) );
  INV_X1 U890 ( .A(n2539), .ZN(n6626) );
  AOI22_X1 U891 ( .A1(\mem[0][2] ), .A2(n2537), .B1(n6868), .B2(data_in[2]), 
        .ZN(n2539) );
  INV_X1 U892 ( .A(n2540), .ZN(n6625) );
  AOI22_X1 U893 ( .A1(\mem[0][3] ), .A2(n2537), .B1(n6868), .B2(data_in[3]), 
        .ZN(n2540) );
  INV_X1 U894 ( .A(n2541), .ZN(n6624) );
  AOI22_X1 U895 ( .A1(\mem[0][4] ), .A2(n2537), .B1(n6868), .B2(data_in[4]), 
        .ZN(n2541) );
  INV_X1 U896 ( .A(n2542), .ZN(n6623) );
  AOI22_X1 U897 ( .A1(\mem[0][5] ), .A2(n2537), .B1(n6868), .B2(data_in[5]), 
        .ZN(n2542) );
  INV_X1 U898 ( .A(n2543), .ZN(n6622) );
  AOI22_X1 U899 ( .A1(\mem[0][6] ), .A2(n2537), .B1(n6868), .B2(data_in[6]), 
        .ZN(n2543) );
  INV_X1 U900 ( .A(n2544), .ZN(n6621) );
  AOI22_X1 U901 ( .A1(\mem[0][7] ), .A2(n2537), .B1(n6868), .B2(data_in[7]), 
        .ZN(n2544) );
  INV_X1 U902 ( .A(n2546), .ZN(n6620) );
  AOI22_X1 U903 ( .A1(\mem[1][0] ), .A2(n2547), .B1(n6867), .B2(data_in[0]), 
        .ZN(n2546) );
  INV_X1 U904 ( .A(n2548), .ZN(n6619) );
  AOI22_X1 U905 ( .A1(\mem[1][1] ), .A2(n2547), .B1(n6867), .B2(data_in[1]), 
        .ZN(n2548) );
  INV_X1 U906 ( .A(n2549), .ZN(n6618) );
  AOI22_X1 U907 ( .A1(\mem[1][2] ), .A2(n2547), .B1(n6867), .B2(data_in[2]), 
        .ZN(n2549) );
  INV_X1 U908 ( .A(n2550), .ZN(n6617) );
  AOI22_X1 U909 ( .A1(\mem[1][3] ), .A2(n2547), .B1(n6867), .B2(data_in[3]), 
        .ZN(n2550) );
  INV_X1 U910 ( .A(n2551), .ZN(n6616) );
  AOI22_X1 U911 ( .A1(\mem[1][4] ), .A2(n2547), .B1(n6867), .B2(data_in[4]), 
        .ZN(n2551) );
  INV_X1 U912 ( .A(n2552), .ZN(n6615) );
  AOI22_X1 U913 ( .A1(\mem[1][5] ), .A2(n2547), .B1(n6867), .B2(data_in[5]), 
        .ZN(n2552) );
  INV_X1 U914 ( .A(n2553), .ZN(n6614) );
  AOI22_X1 U915 ( .A1(\mem[1][6] ), .A2(n2547), .B1(n6867), .B2(data_in[6]), 
        .ZN(n2553) );
  INV_X1 U916 ( .A(n2554), .ZN(n6613) );
  AOI22_X1 U917 ( .A1(\mem[1][7] ), .A2(n2547), .B1(n6867), .B2(data_in[7]), 
        .ZN(n2554) );
  INV_X1 U918 ( .A(n2555), .ZN(n6612) );
  AOI22_X1 U919 ( .A1(\mem[2][0] ), .A2(n2556), .B1(n6866), .B2(data_in[0]), 
        .ZN(n2555) );
  INV_X1 U920 ( .A(n2557), .ZN(n6611) );
  AOI22_X1 U921 ( .A1(\mem[2][1] ), .A2(n2556), .B1(n6866), .B2(data_in[1]), 
        .ZN(n2557) );
  INV_X1 U922 ( .A(n2558), .ZN(n6610) );
  AOI22_X1 U923 ( .A1(\mem[2][2] ), .A2(n2556), .B1(n6866), .B2(data_in[2]), 
        .ZN(n2558) );
  INV_X1 U924 ( .A(n2559), .ZN(n6609) );
  AOI22_X1 U925 ( .A1(\mem[2][3] ), .A2(n2556), .B1(n6866), .B2(data_in[3]), 
        .ZN(n2559) );
  INV_X1 U926 ( .A(n2560), .ZN(n6608) );
  AOI22_X1 U927 ( .A1(\mem[2][4] ), .A2(n2556), .B1(n6866), .B2(data_in[4]), 
        .ZN(n2560) );
  INV_X1 U928 ( .A(n2561), .ZN(n6607) );
  AOI22_X1 U929 ( .A1(\mem[2][5] ), .A2(n2556), .B1(n6866), .B2(data_in[5]), 
        .ZN(n2561) );
  INV_X1 U930 ( .A(n2562), .ZN(n6606) );
  AOI22_X1 U932 ( .A1(\mem[2][6] ), .A2(n2556), .B1(n6866), .B2(data_in[6]), 
        .ZN(n2562) );
  INV_X1 U933 ( .A(n2563), .ZN(n6605) );
  AOI22_X1 U934 ( .A1(\mem[2][7] ), .A2(n2556), .B1(n6866), .B2(data_in[7]), 
        .ZN(n2563) );
  INV_X1 U935 ( .A(n2564), .ZN(n6604) );
  AOI22_X1 U936 ( .A1(\mem[3][0] ), .A2(n2565), .B1(n6865), .B2(data_in[0]), 
        .ZN(n2564) );
  INV_X1 U937 ( .A(n2566), .ZN(n6603) );
  AOI22_X1 U938 ( .A1(\mem[3][1] ), .A2(n2565), .B1(n6865), .B2(data_in[1]), 
        .ZN(n2566) );
  INV_X1 U939 ( .A(n2567), .ZN(n6602) );
  AOI22_X1 U940 ( .A1(\mem[3][2] ), .A2(n2565), .B1(n6865), .B2(data_in[2]), 
        .ZN(n2567) );
  INV_X1 U941 ( .A(n2568), .ZN(n6601) );
  AOI22_X1 U942 ( .A1(\mem[3][3] ), .A2(n2565), .B1(n6865), .B2(data_in[3]), 
        .ZN(n2568) );
  INV_X1 U943 ( .A(n2569), .ZN(n6600) );
  AOI22_X1 U944 ( .A1(\mem[3][4] ), .A2(n2565), .B1(n6865), .B2(data_in[4]), 
        .ZN(n2569) );
  INV_X1 U945 ( .A(n2570), .ZN(n6599) );
  AOI22_X1 U946 ( .A1(\mem[3][5] ), .A2(n2565), .B1(n6865), .B2(data_in[5]), 
        .ZN(n2570) );
  INV_X1 U947 ( .A(n2571), .ZN(n6598) );
  AOI22_X1 U948 ( .A1(\mem[3][6] ), .A2(n2565), .B1(n6865), .B2(data_in[6]), 
        .ZN(n2571) );
  INV_X1 U949 ( .A(n2572), .ZN(n6597) );
  AOI22_X1 U950 ( .A1(\mem[3][7] ), .A2(n2565), .B1(n6865), .B2(data_in[7]), 
        .ZN(n2572) );
  INV_X1 U951 ( .A(n2573), .ZN(n6596) );
  AOI22_X1 U952 ( .A1(\mem[4][0] ), .A2(n2574), .B1(n6864), .B2(data_in[0]), 
        .ZN(n2573) );
  INV_X1 U953 ( .A(n2575), .ZN(n6595) );
  AOI22_X1 U954 ( .A1(\mem[4][1] ), .A2(n2574), .B1(n6864), .B2(data_in[1]), 
        .ZN(n2575) );
  INV_X1 U955 ( .A(n2576), .ZN(n6594) );
  AOI22_X1 U956 ( .A1(\mem[4][2] ), .A2(n2574), .B1(n6864), .B2(data_in[2]), 
        .ZN(n2576) );
  INV_X1 U957 ( .A(n2577), .ZN(n6593) );
  AOI22_X1 U958 ( .A1(\mem[4][3] ), .A2(n2574), .B1(n6864), .B2(data_in[3]), 
        .ZN(n2577) );
  INV_X1 U959 ( .A(n2578), .ZN(n6592) );
  AOI22_X1 U960 ( .A1(\mem[4][4] ), .A2(n2574), .B1(n6864), .B2(data_in[4]), 
        .ZN(n2578) );
  INV_X1 U961 ( .A(n2579), .ZN(n6591) );
  AOI22_X1 U962 ( .A1(\mem[4][5] ), .A2(n2574), .B1(n6864), .B2(data_in[5]), 
        .ZN(n2579) );
  INV_X1 U963 ( .A(n2580), .ZN(n6590) );
  AOI22_X1 U964 ( .A1(\mem[4][6] ), .A2(n2574), .B1(n6864), .B2(data_in[6]), 
        .ZN(n2580) );
  INV_X1 U965 ( .A(n2581), .ZN(n6589) );
  AOI22_X1 U966 ( .A1(\mem[4][7] ), .A2(n2574), .B1(n6864), .B2(data_in[7]), 
        .ZN(n2581) );
  INV_X1 U967 ( .A(n2582), .ZN(n6588) );
  AOI22_X1 U968 ( .A1(\mem[5][0] ), .A2(n2583), .B1(n6863), .B2(data_in[0]), 
        .ZN(n2582) );
  INV_X1 U969 ( .A(n2584), .ZN(n6587) );
  AOI22_X1 U970 ( .A1(\mem[5][1] ), .A2(n2583), .B1(n6863), .B2(data_in[1]), 
        .ZN(n2584) );
  INV_X1 U971 ( .A(n2585), .ZN(n6586) );
  AOI22_X1 U972 ( .A1(\mem[5][2] ), .A2(n2583), .B1(n6863), .B2(data_in[2]), 
        .ZN(n2585) );
  INV_X1 U973 ( .A(n2586), .ZN(n6585) );
  AOI22_X1 U974 ( .A1(\mem[5][3] ), .A2(n2583), .B1(n6863), .B2(data_in[3]), 
        .ZN(n2586) );
  INV_X1 U975 ( .A(n2587), .ZN(n6584) );
  AOI22_X1 U976 ( .A1(\mem[5][4] ), .A2(n2583), .B1(n6863), .B2(data_in[4]), 
        .ZN(n2587) );
  INV_X1 U977 ( .A(n2588), .ZN(n6583) );
  AOI22_X1 U978 ( .A1(\mem[5][5] ), .A2(n2583), .B1(n6863), .B2(data_in[5]), 
        .ZN(n2588) );
  INV_X1 U979 ( .A(n2589), .ZN(n6582) );
  AOI22_X1 U980 ( .A1(\mem[5][6] ), .A2(n2583), .B1(n6863), .B2(data_in[6]), 
        .ZN(n2589) );
  INV_X1 U981 ( .A(n2590), .ZN(n6581) );
  AOI22_X1 U982 ( .A1(\mem[5][7] ), .A2(n2583), .B1(n6863), .B2(data_in[7]), 
        .ZN(n2590) );
  INV_X1 U983 ( .A(n2591), .ZN(n6580) );
  AOI22_X1 U984 ( .A1(\mem[6][0] ), .A2(n2592), .B1(n6862), .B2(data_in[0]), 
        .ZN(n2591) );
  INV_X1 U985 ( .A(n2593), .ZN(n6579) );
  AOI22_X1 U986 ( .A1(\mem[6][1] ), .A2(n2592), .B1(n6862), .B2(data_in[1]), 
        .ZN(n2593) );
  INV_X1 U987 ( .A(n2594), .ZN(n6578) );
  AOI22_X1 U988 ( .A1(\mem[6][2] ), .A2(n2592), .B1(n6862), .B2(data_in[2]), 
        .ZN(n2594) );
  INV_X1 U989 ( .A(n2595), .ZN(n6577) );
  AOI22_X1 U990 ( .A1(\mem[6][3] ), .A2(n2592), .B1(n6862), .B2(data_in[3]), 
        .ZN(n2595) );
  INV_X1 U991 ( .A(n2596), .ZN(n6576) );
  AOI22_X1 U992 ( .A1(\mem[6][4] ), .A2(n2592), .B1(n6862), .B2(data_in[4]), 
        .ZN(n2596) );
  INV_X1 U993 ( .A(n2597), .ZN(n6575) );
  AOI22_X1 U994 ( .A1(\mem[6][5] ), .A2(n2592), .B1(n6862), .B2(data_in[5]), 
        .ZN(n2597) );
  INV_X1 U995 ( .A(n2598), .ZN(n6574) );
  AOI22_X1 U996 ( .A1(\mem[6][6] ), .A2(n2592), .B1(n6862), .B2(data_in[6]), 
        .ZN(n2598) );
  INV_X1 U997 ( .A(n2599), .ZN(n6573) );
  AOI22_X1 U998 ( .A1(\mem[6][7] ), .A2(n2592), .B1(n6862), .B2(data_in[7]), 
        .ZN(n2599) );
  INV_X1 U999 ( .A(n2600), .ZN(n6572) );
  AOI22_X1 U1000 ( .A1(\mem[7][0] ), .A2(n2601), .B1(n6861), .B2(data_in[0]), 
        .ZN(n2600) );
  INV_X1 U1001 ( .A(n2602), .ZN(n6571) );
  AOI22_X1 U1002 ( .A1(\mem[7][1] ), .A2(n2601), .B1(n6861), .B2(data_in[1]), 
        .ZN(n2602) );
  INV_X1 U1003 ( .A(n2603), .ZN(n6570) );
  AOI22_X1 U1004 ( .A1(\mem[7][2] ), .A2(n2601), .B1(n6861), .B2(data_in[2]), 
        .ZN(n2603) );
  INV_X1 U1005 ( .A(n2604), .ZN(n6569) );
  AOI22_X1 U1006 ( .A1(\mem[7][3] ), .A2(n2601), .B1(n6861), .B2(data_in[3]), 
        .ZN(n2604) );
  INV_X1 U1007 ( .A(n2605), .ZN(n6568) );
  AOI22_X1 U1008 ( .A1(\mem[7][4] ), .A2(n2601), .B1(n6861), .B2(data_in[4]), 
        .ZN(n2605) );
  INV_X1 U1009 ( .A(n2606), .ZN(n6567) );
  AOI22_X1 U1010 ( .A1(\mem[7][5] ), .A2(n2601), .B1(n6861), .B2(data_in[5]), 
        .ZN(n2606) );
  INV_X1 U1011 ( .A(n2607), .ZN(n6566) );
  AOI22_X1 U1012 ( .A1(\mem[7][6] ), .A2(n2601), .B1(n6861), .B2(data_in[6]), 
        .ZN(n2607) );
  INV_X1 U1013 ( .A(n2608), .ZN(n6565) );
  AOI22_X1 U1014 ( .A1(\mem[7][7] ), .A2(n2601), .B1(n6861), .B2(data_in[7]), 
        .ZN(n2608) );
  INV_X1 U1015 ( .A(n2609), .ZN(n6564) );
  AOI22_X1 U1016 ( .A1(\mem[8][0] ), .A2(n2610), .B1(n6860), .B2(data_in[0]), 
        .ZN(n2609) );
  INV_X1 U1017 ( .A(n2611), .ZN(n6563) );
  AOI22_X1 U1018 ( .A1(\mem[8][1] ), .A2(n2610), .B1(n6860), .B2(data_in[1]), 
        .ZN(n2611) );
  INV_X1 U1019 ( .A(n2612), .ZN(n6562) );
  AOI22_X1 U1020 ( .A1(\mem[8][2] ), .A2(n2610), .B1(n6860), .B2(data_in[2]), 
        .ZN(n2612) );
  INV_X1 U1021 ( .A(n2613), .ZN(n6561) );
  AOI22_X1 U1022 ( .A1(\mem[8][3] ), .A2(n2610), .B1(n6860), .B2(data_in[3]), 
        .ZN(n2613) );
  INV_X1 U1023 ( .A(n2614), .ZN(n6560) );
  AOI22_X1 U1024 ( .A1(\mem[8][4] ), .A2(n2610), .B1(n6860), .B2(data_in[4]), 
        .ZN(n2614) );
  INV_X1 U1025 ( .A(n2615), .ZN(n6559) );
  AOI22_X1 U1026 ( .A1(\mem[8][5] ), .A2(n2610), .B1(n6860), .B2(data_in[5]), 
        .ZN(n2615) );
  INV_X1 U1027 ( .A(n2616), .ZN(n6558) );
  AOI22_X1 U1028 ( .A1(\mem[8][6] ), .A2(n2610), .B1(n6860), .B2(data_in[6]), 
        .ZN(n2616) );
  INV_X1 U1029 ( .A(n2617), .ZN(n6557) );
  AOI22_X1 U1030 ( .A1(\mem[8][7] ), .A2(n2610), .B1(n6860), .B2(data_in[7]), 
        .ZN(n2617) );
  INV_X1 U1031 ( .A(n2618), .ZN(n6556) );
  AOI22_X1 U1032 ( .A1(\mem[9][0] ), .A2(n2619), .B1(n6859), .B2(data_in[0]), 
        .ZN(n2618) );
  INV_X1 U1033 ( .A(n2620), .ZN(n6555) );
  AOI22_X1 U1034 ( .A1(\mem[9][1] ), .A2(n2619), .B1(n6859), .B2(data_in[1]), 
        .ZN(n2620) );
  INV_X1 U1035 ( .A(n2621), .ZN(n6554) );
  AOI22_X1 U1036 ( .A1(\mem[9][2] ), .A2(n2619), .B1(n6859), .B2(data_in[2]), 
        .ZN(n2621) );
  INV_X1 U1037 ( .A(n2622), .ZN(n6553) );
  AOI22_X1 U1038 ( .A1(\mem[9][3] ), .A2(n2619), .B1(n6859), .B2(data_in[3]), 
        .ZN(n2622) );
  INV_X1 U1039 ( .A(n2623), .ZN(n6552) );
  AOI22_X1 U1040 ( .A1(\mem[9][4] ), .A2(n2619), .B1(n6859), .B2(data_in[4]), 
        .ZN(n2623) );
  INV_X1 U1041 ( .A(n2624), .ZN(n6551) );
  AOI22_X1 U1042 ( .A1(\mem[9][5] ), .A2(n2619), .B1(n6859), .B2(data_in[5]), 
        .ZN(n2624) );
  INV_X1 U1043 ( .A(n2625), .ZN(n6550) );
  AOI22_X1 U1044 ( .A1(\mem[9][6] ), .A2(n2619), .B1(n6859), .B2(data_in[6]), 
        .ZN(n2625) );
  INV_X1 U1045 ( .A(n2626), .ZN(n6549) );
  AOI22_X1 U1046 ( .A1(\mem[9][7] ), .A2(n2619), .B1(n6859), .B2(data_in[7]), 
        .ZN(n2626) );
  INV_X1 U1047 ( .A(n2627), .ZN(n6548) );
  AOI22_X1 U1048 ( .A1(\mem[10][0] ), .A2(n2628), .B1(n6858), .B2(data_in[0]), 
        .ZN(n2627) );
  INV_X1 U1049 ( .A(n2629), .ZN(n6547) );
  AOI22_X1 U1050 ( .A1(\mem[10][1] ), .A2(n2628), .B1(n6858), .B2(data_in[1]), 
        .ZN(n2629) );
  INV_X1 U1051 ( .A(n2630), .ZN(n6546) );
  AOI22_X1 U1052 ( .A1(\mem[10][2] ), .A2(n2628), .B1(n6858), .B2(data_in[2]), 
        .ZN(n2630) );
  INV_X1 U1053 ( .A(n2631), .ZN(n6545) );
  AOI22_X1 U1054 ( .A1(\mem[10][3] ), .A2(n2628), .B1(n6858), .B2(data_in[3]), 
        .ZN(n2631) );
  INV_X1 U1055 ( .A(n2632), .ZN(n6544) );
  AOI22_X1 U1056 ( .A1(\mem[10][4] ), .A2(n2628), .B1(n6858), .B2(data_in[4]), 
        .ZN(n2632) );
  INV_X1 U1057 ( .A(n2633), .ZN(n6543) );
  AOI22_X1 U1058 ( .A1(\mem[10][5] ), .A2(n2628), .B1(n6858), .B2(data_in[5]), 
        .ZN(n2633) );
  INV_X1 U1059 ( .A(n2634), .ZN(n6542) );
  AOI22_X1 U1060 ( .A1(\mem[10][6] ), .A2(n2628), .B1(n6858), .B2(data_in[6]), 
        .ZN(n2634) );
  INV_X1 U1061 ( .A(n2635), .ZN(n6541) );
  AOI22_X1 U1062 ( .A1(\mem[10][7] ), .A2(n2628), .B1(n6858), .B2(data_in[7]), 
        .ZN(n2635) );
  INV_X1 U1063 ( .A(n2636), .ZN(n6540) );
  AOI22_X1 U1064 ( .A1(\mem[11][0] ), .A2(n2637), .B1(n6857), .B2(data_in[0]), 
        .ZN(n2636) );
  INV_X1 U1065 ( .A(n2638), .ZN(n6539) );
  AOI22_X1 U1066 ( .A1(\mem[11][1] ), .A2(n2637), .B1(n6857), .B2(data_in[1]), 
        .ZN(n2638) );
  INV_X1 U1067 ( .A(n2639), .ZN(n6538) );
  AOI22_X1 U1068 ( .A1(\mem[11][2] ), .A2(n2637), .B1(n6857), .B2(data_in[2]), 
        .ZN(n2639) );
  INV_X1 U1069 ( .A(n2640), .ZN(n6537) );
  AOI22_X1 U1070 ( .A1(\mem[11][3] ), .A2(n2637), .B1(n6857), .B2(data_in[3]), 
        .ZN(n2640) );
  INV_X1 U1071 ( .A(n2641), .ZN(n6536) );
  AOI22_X1 U1072 ( .A1(\mem[11][4] ), .A2(n2637), .B1(n6857), .B2(data_in[4]), 
        .ZN(n2641) );
  INV_X1 U1073 ( .A(n2642), .ZN(n6535) );
  AOI22_X1 U1074 ( .A1(\mem[11][5] ), .A2(n2637), .B1(n6857), .B2(data_in[5]), 
        .ZN(n2642) );
  INV_X1 U1075 ( .A(n2643), .ZN(n6534) );
  AOI22_X1 U1077 ( .A1(\mem[11][6] ), .A2(n2637), .B1(n6857), .B2(data_in[6]), 
        .ZN(n2643) );
  INV_X1 U1078 ( .A(n2644), .ZN(n6533) );
  AOI22_X1 U1079 ( .A1(\mem[11][7] ), .A2(n2637), .B1(n6857), .B2(data_in[7]), 
        .ZN(n2644) );
  INV_X1 U1080 ( .A(n2645), .ZN(n6532) );
  AOI22_X1 U1081 ( .A1(\mem[12][0] ), .A2(n2646), .B1(n6856), .B2(data_in[0]), 
        .ZN(n2645) );
  INV_X1 U1082 ( .A(n2647), .ZN(n6531) );
  AOI22_X1 U1083 ( .A1(\mem[12][1] ), .A2(n2646), .B1(n6856), .B2(data_in[1]), 
        .ZN(n2647) );
  INV_X1 U1084 ( .A(n2648), .ZN(n6530) );
  AOI22_X1 U1085 ( .A1(\mem[12][2] ), .A2(n2646), .B1(n6856), .B2(data_in[2]), 
        .ZN(n2648) );
  INV_X1 U1086 ( .A(n2649), .ZN(n6529) );
  AOI22_X1 U1087 ( .A1(\mem[12][3] ), .A2(n2646), .B1(n6856), .B2(data_in[3]), 
        .ZN(n2649) );
  INV_X1 U1088 ( .A(n2650), .ZN(n6528) );
  AOI22_X1 U1089 ( .A1(\mem[12][4] ), .A2(n2646), .B1(n6856), .B2(data_in[4]), 
        .ZN(n2650) );
  INV_X1 U1090 ( .A(n2651), .ZN(n6527) );
  AOI22_X1 U1091 ( .A1(\mem[12][5] ), .A2(n2646), .B1(n6856), .B2(data_in[5]), 
        .ZN(n2651) );
  INV_X1 U1092 ( .A(n2652), .ZN(n6526) );
  AOI22_X1 U1093 ( .A1(\mem[12][6] ), .A2(n2646), .B1(n6856), .B2(data_in[6]), 
        .ZN(n2652) );
  INV_X1 U1094 ( .A(n2653), .ZN(n6525) );
  AOI22_X1 U1095 ( .A1(\mem[12][7] ), .A2(n2646), .B1(n6856), .B2(data_in[7]), 
        .ZN(n2653) );
  INV_X1 U1096 ( .A(n2654), .ZN(n6524) );
  AOI22_X1 U1097 ( .A1(\mem[13][0] ), .A2(n2655), .B1(n6855), .B2(data_in[0]), 
        .ZN(n2654) );
  INV_X1 U1098 ( .A(n2656), .ZN(n6523) );
  AOI22_X1 U1099 ( .A1(\mem[13][1] ), .A2(n2655), .B1(n6855), .B2(data_in[1]), 
        .ZN(n2656) );
  INV_X1 U1100 ( .A(n2657), .ZN(n6522) );
  AOI22_X1 U1101 ( .A1(\mem[13][2] ), .A2(n2655), .B1(n6855), .B2(data_in[2]), 
        .ZN(n2657) );
  INV_X1 U1102 ( .A(n2658), .ZN(n6521) );
  AOI22_X1 U1103 ( .A1(\mem[13][3] ), .A2(n2655), .B1(n6855), .B2(data_in[3]), 
        .ZN(n2658) );
  INV_X1 U1104 ( .A(n2659), .ZN(n6520) );
  AOI22_X1 U1105 ( .A1(\mem[13][4] ), .A2(n2655), .B1(n6855), .B2(data_in[4]), 
        .ZN(n2659) );
  INV_X1 U1106 ( .A(n2660), .ZN(n6519) );
  AOI22_X1 U1107 ( .A1(\mem[13][5] ), .A2(n2655), .B1(n6855), .B2(data_in[5]), 
        .ZN(n2660) );
  INV_X1 U1108 ( .A(n2661), .ZN(n6518) );
  AOI22_X1 U1109 ( .A1(\mem[13][6] ), .A2(n2655), .B1(n6855), .B2(data_in[6]), 
        .ZN(n2661) );
  INV_X1 U1110 ( .A(n2662), .ZN(n6517) );
  AOI22_X1 U1111 ( .A1(\mem[13][7] ), .A2(n2655), .B1(n6855), .B2(data_in[7]), 
        .ZN(n2662) );
  INV_X1 U1112 ( .A(n2663), .ZN(n6516) );
  AOI22_X1 U1113 ( .A1(\mem[14][0] ), .A2(n2664), .B1(n6854), .B2(data_in[0]), 
        .ZN(n2663) );
  INV_X1 U1114 ( .A(n2665), .ZN(n6515) );
  AOI22_X1 U1115 ( .A1(\mem[14][1] ), .A2(n2664), .B1(n6854), .B2(data_in[1]), 
        .ZN(n2665) );
  INV_X1 U1116 ( .A(n2666), .ZN(n6514) );
  AOI22_X1 U1117 ( .A1(\mem[14][2] ), .A2(n2664), .B1(n6854), .B2(data_in[2]), 
        .ZN(n2666) );
  INV_X1 U1118 ( .A(n2667), .ZN(n6513) );
  AOI22_X1 U1119 ( .A1(\mem[14][3] ), .A2(n2664), .B1(n6854), .B2(data_in[3]), 
        .ZN(n2667) );
  INV_X1 U1120 ( .A(n2668), .ZN(n6512) );
  AOI22_X1 U1121 ( .A1(\mem[14][4] ), .A2(n2664), .B1(n6854), .B2(data_in[4]), 
        .ZN(n2668) );
  INV_X1 U1122 ( .A(n2669), .ZN(n6511) );
  AOI22_X1 U1123 ( .A1(\mem[14][5] ), .A2(n2664), .B1(n6854), .B2(data_in[5]), 
        .ZN(n2669) );
  INV_X1 U1124 ( .A(n2670), .ZN(n6510) );
  AOI22_X1 U1125 ( .A1(\mem[14][6] ), .A2(n2664), .B1(n6854), .B2(data_in[6]), 
        .ZN(n2670) );
  INV_X1 U1126 ( .A(n2671), .ZN(n6509) );
  AOI22_X1 U1127 ( .A1(\mem[14][7] ), .A2(n2664), .B1(n6854), .B2(data_in[7]), 
        .ZN(n2671) );
  INV_X1 U1128 ( .A(n2672), .ZN(n6508) );
  AOI22_X1 U1129 ( .A1(\mem[15][0] ), .A2(n2673), .B1(n6853), .B2(data_in[0]), 
        .ZN(n2672) );
  INV_X1 U1130 ( .A(n2674), .ZN(n6507) );
  AOI22_X1 U1131 ( .A1(\mem[15][1] ), .A2(n2673), .B1(n6853), .B2(data_in[1]), 
        .ZN(n2674) );
  INV_X1 U1132 ( .A(n2675), .ZN(n6506) );
  AOI22_X1 U1133 ( .A1(\mem[15][2] ), .A2(n2673), .B1(n6853), .B2(data_in[2]), 
        .ZN(n2675) );
  INV_X1 U1134 ( .A(n2676), .ZN(n6505) );
  AOI22_X1 U1135 ( .A1(\mem[15][3] ), .A2(n2673), .B1(n6853), .B2(data_in[3]), 
        .ZN(n2676) );
  INV_X1 U1136 ( .A(n2677), .ZN(n6504) );
  AOI22_X1 U1137 ( .A1(\mem[15][4] ), .A2(n2673), .B1(n6853), .B2(data_in[4]), 
        .ZN(n2677) );
  INV_X1 U1138 ( .A(n2678), .ZN(n6503) );
  AOI22_X1 U1139 ( .A1(\mem[15][5] ), .A2(n2673), .B1(n6853), .B2(data_in[5]), 
        .ZN(n2678) );
  INV_X1 U1140 ( .A(n2679), .ZN(n6502) );
  AOI22_X1 U1141 ( .A1(\mem[15][6] ), .A2(n2673), .B1(n6853), .B2(data_in[6]), 
        .ZN(n2679) );
  INV_X1 U1142 ( .A(n2680), .ZN(n6501) );
  AOI22_X1 U1143 ( .A1(\mem[15][7] ), .A2(n2673), .B1(n6853), .B2(data_in[7]), 
        .ZN(n2680) );
  INV_X1 U1144 ( .A(n2683), .ZN(n6500) );
  AOI22_X1 U1145 ( .A1(\mem[16][0] ), .A2(n2684), .B1(n6852), .B2(data_in[0]), 
        .ZN(n2683) );
  INV_X1 U1146 ( .A(n2685), .ZN(n6499) );
  AOI22_X1 U1147 ( .A1(\mem[16][1] ), .A2(n2684), .B1(n6852), .B2(data_in[1]), 
        .ZN(n2685) );
  INV_X1 U1148 ( .A(n2686), .ZN(n6498) );
  AOI22_X1 U1149 ( .A1(\mem[16][2] ), .A2(n2684), .B1(n6852), .B2(data_in[2]), 
        .ZN(n2686) );
  INV_X1 U1150 ( .A(n2687), .ZN(n6497) );
  AOI22_X1 U1151 ( .A1(\mem[16][3] ), .A2(n2684), .B1(n6852), .B2(data_in[3]), 
        .ZN(n2687) );
  INV_X1 U1152 ( .A(n2688), .ZN(n6496) );
  AOI22_X1 U1153 ( .A1(\mem[16][4] ), .A2(n2684), .B1(n6852), .B2(data_in[4]), 
        .ZN(n2688) );
  INV_X1 U1154 ( .A(n2689), .ZN(n6495) );
  AOI22_X1 U1155 ( .A1(\mem[16][5] ), .A2(n2684), .B1(n6852), .B2(data_in[5]), 
        .ZN(n2689) );
  INV_X1 U1156 ( .A(n2690), .ZN(n6494) );
  AOI22_X1 U1157 ( .A1(\mem[16][6] ), .A2(n2684), .B1(n6852), .B2(data_in[6]), 
        .ZN(n2690) );
  INV_X1 U1158 ( .A(n2691), .ZN(n6493) );
  AOI22_X1 U1159 ( .A1(\mem[16][7] ), .A2(n2684), .B1(n6852), .B2(data_in[7]), 
        .ZN(n2691) );
  INV_X1 U1160 ( .A(n2693), .ZN(n6492) );
  AOI22_X1 U1161 ( .A1(\mem[17][0] ), .A2(n2694), .B1(n6851), .B2(data_in[0]), 
        .ZN(n2693) );
  INV_X1 U1162 ( .A(n2695), .ZN(n6491) );
  AOI22_X1 U1163 ( .A1(\mem[17][1] ), .A2(n2694), .B1(n6851), .B2(data_in[1]), 
        .ZN(n2695) );
  INV_X1 U1164 ( .A(n2696), .ZN(n6490) );
  AOI22_X1 U1165 ( .A1(\mem[17][2] ), .A2(n2694), .B1(n6851), .B2(data_in[2]), 
        .ZN(n2696) );
  INV_X1 U1166 ( .A(n2697), .ZN(n6489) );
  AOI22_X1 U1167 ( .A1(\mem[17][3] ), .A2(n2694), .B1(n6851), .B2(data_in[3]), 
        .ZN(n2697) );
  INV_X1 U1168 ( .A(n2698), .ZN(n6488) );
  AOI22_X1 U1169 ( .A1(\mem[17][4] ), .A2(n2694), .B1(n6851), .B2(data_in[4]), 
        .ZN(n2698) );
  INV_X1 U1170 ( .A(n2699), .ZN(n6487) );
  AOI22_X1 U1171 ( .A1(\mem[17][5] ), .A2(n2694), .B1(n6851), .B2(data_in[5]), 
        .ZN(n2699) );
  INV_X1 U1172 ( .A(n2700), .ZN(n6486) );
  AOI22_X1 U1173 ( .A1(\mem[17][6] ), .A2(n2694), .B1(n6851), .B2(data_in[6]), 
        .ZN(n2700) );
  INV_X1 U1174 ( .A(n2701), .ZN(n6485) );
  AOI22_X1 U1175 ( .A1(\mem[17][7] ), .A2(n2694), .B1(n6851), .B2(data_in[7]), 
        .ZN(n2701) );
  INV_X1 U1176 ( .A(n2702), .ZN(n6484) );
  AOI22_X1 U1177 ( .A1(\mem[18][0] ), .A2(n2703), .B1(n6850), .B2(data_in[0]), 
        .ZN(n2702) );
  INV_X1 U1178 ( .A(n2704), .ZN(n6483) );
  AOI22_X1 U1179 ( .A1(\mem[18][1] ), .A2(n2703), .B1(n6850), .B2(data_in[1]), 
        .ZN(n2704) );
  INV_X1 U1180 ( .A(n2705), .ZN(n6482) );
  AOI22_X1 U1181 ( .A1(\mem[18][2] ), .A2(n2703), .B1(n6850), .B2(data_in[2]), 
        .ZN(n2705) );
  INV_X1 U1182 ( .A(n2706), .ZN(n6481) );
  AOI22_X1 U1183 ( .A1(\mem[18][3] ), .A2(n2703), .B1(n6850), .B2(data_in[3]), 
        .ZN(n2706) );
  INV_X1 U1184 ( .A(n2707), .ZN(n6480) );
  AOI22_X1 U1185 ( .A1(\mem[18][4] ), .A2(n2703), .B1(n6850), .B2(data_in[4]), 
        .ZN(n2707) );
  INV_X1 U1186 ( .A(n2708), .ZN(n6479) );
  AOI22_X1 U1187 ( .A1(\mem[18][5] ), .A2(n2703), .B1(n6850), .B2(data_in[5]), 
        .ZN(n2708) );
  INV_X1 U1188 ( .A(n2709), .ZN(n6478) );
  AOI22_X1 U1189 ( .A1(\mem[18][6] ), .A2(n2703), .B1(n6850), .B2(data_in[6]), 
        .ZN(n2709) );
  INV_X1 U1190 ( .A(n2710), .ZN(n6477) );
  AOI22_X1 U1191 ( .A1(\mem[18][7] ), .A2(n2703), .B1(n6850), .B2(data_in[7]), 
        .ZN(n2710) );
  INV_X1 U1192 ( .A(n2711), .ZN(n6476) );
  AOI22_X1 U1193 ( .A1(\mem[19][0] ), .A2(n2712), .B1(n6849), .B2(data_in[0]), 
        .ZN(n2711) );
  INV_X1 U1194 ( .A(n2713), .ZN(n6475) );
  AOI22_X1 U1195 ( .A1(\mem[19][1] ), .A2(n2712), .B1(n6849), .B2(data_in[1]), 
        .ZN(n2713) );
  INV_X1 U1196 ( .A(n2714), .ZN(n6474) );
  AOI22_X1 U1197 ( .A1(\mem[19][2] ), .A2(n2712), .B1(n6849), .B2(data_in[2]), 
        .ZN(n2714) );
  INV_X1 U1198 ( .A(n2715), .ZN(n6473) );
  AOI22_X1 U1199 ( .A1(\mem[19][3] ), .A2(n2712), .B1(n6849), .B2(data_in[3]), 
        .ZN(n2715) );
  INV_X1 U1200 ( .A(n2716), .ZN(n6472) );
  AOI22_X1 U1201 ( .A1(\mem[19][4] ), .A2(n2712), .B1(n6849), .B2(data_in[4]), 
        .ZN(n2716) );
  INV_X1 U1202 ( .A(n2717), .ZN(n6471) );
  AOI22_X1 U1203 ( .A1(\mem[19][5] ), .A2(n2712), .B1(n6849), .B2(data_in[5]), 
        .ZN(n2717) );
  INV_X1 U1204 ( .A(n2718), .ZN(n6470) );
  AOI22_X1 U1205 ( .A1(\mem[19][6] ), .A2(n2712), .B1(n6849), .B2(data_in[6]), 
        .ZN(n2718) );
  INV_X1 U1206 ( .A(n2719), .ZN(n6469) );
  AOI22_X1 U1207 ( .A1(\mem[19][7] ), .A2(n2712), .B1(n6849), .B2(data_in[7]), 
        .ZN(n2719) );
  INV_X1 U1208 ( .A(n2720), .ZN(n6468) );
  AOI22_X1 U1209 ( .A1(\mem[20][0] ), .A2(n2721), .B1(n6848), .B2(data_in[0]), 
        .ZN(n2720) );
  INV_X1 U1210 ( .A(n2722), .ZN(n6467) );
  AOI22_X1 U1211 ( .A1(\mem[20][1] ), .A2(n2721), .B1(n6848), .B2(data_in[1]), 
        .ZN(n2722) );
  INV_X1 U1212 ( .A(n2723), .ZN(n6466) );
  AOI22_X1 U1213 ( .A1(\mem[20][2] ), .A2(n2721), .B1(n6848), .B2(data_in[2]), 
        .ZN(n2723) );
  INV_X1 U1214 ( .A(n2724), .ZN(n6465) );
  AOI22_X1 U1215 ( .A1(\mem[20][3] ), .A2(n2721), .B1(n6848), .B2(data_in[3]), 
        .ZN(n2724) );
  INV_X1 U1216 ( .A(n2725), .ZN(n6464) );
  AOI22_X1 U1217 ( .A1(\mem[20][4] ), .A2(n2721), .B1(n6848), .B2(data_in[4]), 
        .ZN(n2725) );
  INV_X1 U1218 ( .A(n2726), .ZN(n6463) );
  AOI22_X1 U1219 ( .A1(\mem[20][5] ), .A2(n2721), .B1(n6848), .B2(data_in[5]), 
        .ZN(n2726) );
  INV_X1 U1220 ( .A(n2727), .ZN(n6462) );
  AOI22_X1 U1222 ( .A1(\mem[20][6] ), .A2(n2721), .B1(n6848), .B2(data_in[6]), 
        .ZN(n2727) );
  INV_X1 U1223 ( .A(n2728), .ZN(n6461) );
  AOI22_X1 U1224 ( .A1(\mem[20][7] ), .A2(n2721), .B1(n6848), .B2(data_in[7]), 
        .ZN(n2728) );
  INV_X1 U1225 ( .A(n2729), .ZN(n6460) );
  AOI22_X1 U1226 ( .A1(\mem[21][0] ), .A2(n2730), .B1(n6847), .B2(data_in[0]), 
        .ZN(n2729) );
  INV_X1 U1227 ( .A(n2731), .ZN(n6459) );
  AOI22_X1 U1228 ( .A1(\mem[21][1] ), .A2(n2730), .B1(n6847), .B2(data_in[1]), 
        .ZN(n2731) );
  INV_X1 U1229 ( .A(n2732), .ZN(n6458) );
  AOI22_X1 U1230 ( .A1(\mem[21][2] ), .A2(n2730), .B1(n6847), .B2(data_in[2]), 
        .ZN(n2732) );
  INV_X1 U1231 ( .A(n2733), .ZN(n6457) );
  AOI22_X1 U1232 ( .A1(\mem[21][3] ), .A2(n2730), .B1(n6847), .B2(data_in[3]), 
        .ZN(n2733) );
  INV_X1 U1233 ( .A(n2734), .ZN(n6456) );
  AOI22_X1 U1234 ( .A1(\mem[21][4] ), .A2(n2730), .B1(n6847), .B2(data_in[4]), 
        .ZN(n2734) );
  INV_X1 U1235 ( .A(n2735), .ZN(n6455) );
  AOI22_X1 U1236 ( .A1(\mem[21][5] ), .A2(n2730), .B1(n6847), .B2(data_in[5]), 
        .ZN(n2735) );
  INV_X1 U1237 ( .A(n2736), .ZN(n6454) );
  AOI22_X1 U1238 ( .A1(\mem[21][6] ), .A2(n2730), .B1(n6847), .B2(data_in[6]), 
        .ZN(n2736) );
  INV_X1 U1239 ( .A(n2737), .ZN(n6453) );
  AOI22_X1 U1240 ( .A1(\mem[21][7] ), .A2(n2730), .B1(n6847), .B2(data_in[7]), 
        .ZN(n2737) );
  INV_X1 U1241 ( .A(n2738), .ZN(n6452) );
  AOI22_X1 U1242 ( .A1(\mem[22][0] ), .A2(n2739), .B1(n6846), .B2(data_in[0]), 
        .ZN(n2738) );
  INV_X1 U1243 ( .A(n2740), .ZN(n6451) );
  AOI22_X1 U1244 ( .A1(\mem[22][1] ), .A2(n2739), .B1(n6846), .B2(data_in[1]), 
        .ZN(n2740) );
  INV_X1 U1245 ( .A(n2741), .ZN(n6450) );
  AOI22_X1 U1246 ( .A1(\mem[22][2] ), .A2(n2739), .B1(n6846), .B2(data_in[2]), 
        .ZN(n2741) );
  INV_X1 U1247 ( .A(n2742), .ZN(n6449) );
  AOI22_X1 U1248 ( .A1(\mem[22][3] ), .A2(n2739), .B1(n6846), .B2(data_in[3]), 
        .ZN(n2742) );
  INV_X1 U1249 ( .A(n2743), .ZN(n6448) );
  AOI22_X1 U1250 ( .A1(\mem[22][4] ), .A2(n2739), .B1(n6846), .B2(data_in[4]), 
        .ZN(n2743) );
  INV_X1 U1251 ( .A(n2744), .ZN(n6447) );
  AOI22_X1 U1252 ( .A1(\mem[22][5] ), .A2(n2739), .B1(n6846), .B2(data_in[5]), 
        .ZN(n2744) );
  INV_X1 U1253 ( .A(n2745), .ZN(n6446) );
  AOI22_X1 U1254 ( .A1(\mem[22][6] ), .A2(n2739), .B1(n6846), .B2(data_in[6]), 
        .ZN(n2745) );
  INV_X1 U1255 ( .A(n2746), .ZN(n6445) );
  AOI22_X1 U1256 ( .A1(\mem[22][7] ), .A2(n2739), .B1(n6846), .B2(data_in[7]), 
        .ZN(n2746) );
  INV_X1 U1257 ( .A(n2747), .ZN(n6444) );
  AOI22_X1 U1258 ( .A1(\mem[23][0] ), .A2(n2748), .B1(n6845), .B2(data_in[0]), 
        .ZN(n2747) );
  INV_X1 U1259 ( .A(n2749), .ZN(n6443) );
  AOI22_X1 U1260 ( .A1(\mem[23][1] ), .A2(n2748), .B1(n6845), .B2(data_in[1]), 
        .ZN(n2749) );
  INV_X1 U1261 ( .A(n2750), .ZN(n6442) );
  AOI22_X1 U1262 ( .A1(\mem[23][2] ), .A2(n2748), .B1(n6845), .B2(data_in[2]), 
        .ZN(n2750) );
  INV_X1 U1263 ( .A(n2751), .ZN(n6441) );
  AOI22_X1 U1264 ( .A1(\mem[23][3] ), .A2(n2748), .B1(n6845), .B2(data_in[3]), 
        .ZN(n2751) );
  INV_X1 U1265 ( .A(n2752), .ZN(n6440) );
  AOI22_X1 U1266 ( .A1(\mem[23][4] ), .A2(n2748), .B1(n6845), .B2(data_in[4]), 
        .ZN(n2752) );
  INV_X1 U1267 ( .A(n2753), .ZN(n6439) );
  AOI22_X1 U1268 ( .A1(\mem[23][5] ), .A2(n2748), .B1(n6845), .B2(data_in[5]), 
        .ZN(n2753) );
  INV_X1 U1269 ( .A(n2754), .ZN(n6438) );
  AOI22_X1 U1270 ( .A1(\mem[23][6] ), .A2(n2748), .B1(n6845), .B2(data_in[6]), 
        .ZN(n2754) );
  INV_X1 U1271 ( .A(n2755), .ZN(n6437) );
  AOI22_X1 U1272 ( .A1(\mem[23][7] ), .A2(n2748), .B1(n6845), .B2(data_in[7]), 
        .ZN(n2755) );
  INV_X1 U1273 ( .A(n2756), .ZN(n6436) );
  AOI22_X1 U1274 ( .A1(\mem[24][0] ), .A2(n2757), .B1(n6844), .B2(data_in[0]), 
        .ZN(n2756) );
  INV_X1 U1275 ( .A(n2758), .ZN(n6435) );
  AOI22_X1 U1276 ( .A1(\mem[24][1] ), .A2(n2757), .B1(n6844), .B2(data_in[1]), 
        .ZN(n2758) );
  INV_X1 U1277 ( .A(n2759), .ZN(n6434) );
  AOI22_X1 U1278 ( .A1(\mem[24][2] ), .A2(n2757), .B1(n6844), .B2(data_in[2]), 
        .ZN(n2759) );
  INV_X1 U1279 ( .A(n2760), .ZN(n6433) );
  AOI22_X1 U1280 ( .A1(\mem[24][3] ), .A2(n2757), .B1(n6844), .B2(data_in[3]), 
        .ZN(n2760) );
  INV_X1 U1281 ( .A(n2761), .ZN(n6432) );
  AOI22_X1 U1282 ( .A1(\mem[24][4] ), .A2(n2757), .B1(n6844), .B2(data_in[4]), 
        .ZN(n2761) );
  INV_X1 U1283 ( .A(n2762), .ZN(n6431) );
  AOI22_X1 U1284 ( .A1(\mem[24][5] ), .A2(n2757), .B1(n6844), .B2(data_in[5]), 
        .ZN(n2762) );
  INV_X1 U1285 ( .A(n2763), .ZN(n6430) );
  AOI22_X1 U1286 ( .A1(\mem[24][6] ), .A2(n2757), .B1(n6844), .B2(data_in[6]), 
        .ZN(n2763) );
  INV_X1 U1287 ( .A(n2764), .ZN(n6429) );
  AOI22_X1 U1288 ( .A1(\mem[24][7] ), .A2(n2757), .B1(n6844), .B2(data_in[7]), 
        .ZN(n2764) );
  INV_X1 U1289 ( .A(n2765), .ZN(n6428) );
  AOI22_X1 U1290 ( .A1(\mem[25][0] ), .A2(n2766), .B1(n6843), .B2(data_in[0]), 
        .ZN(n2765) );
  INV_X1 U1291 ( .A(n2767), .ZN(n6427) );
  AOI22_X1 U1292 ( .A1(\mem[25][1] ), .A2(n2766), .B1(n6843), .B2(data_in[1]), 
        .ZN(n2767) );
  INV_X1 U1293 ( .A(n2768), .ZN(n6426) );
  AOI22_X1 U1294 ( .A1(\mem[25][2] ), .A2(n2766), .B1(n6843), .B2(data_in[2]), 
        .ZN(n2768) );
  INV_X1 U1295 ( .A(n2769), .ZN(n6425) );
  AOI22_X1 U1296 ( .A1(\mem[25][3] ), .A2(n2766), .B1(n6843), .B2(data_in[3]), 
        .ZN(n2769) );
  INV_X1 U1297 ( .A(n2770), .ZN(n6424) );
  AOI22_X1 U1298 ( .A1(\mem[25][4] ), .A2(n2766), .B1(n6843), .B2(data_in[4]), 
        .ZN(n2770) );
  INV_X1 U1299 ( .A(n2771), .ZN(n6423) );
  AOI22_X1 U1300 ( .A1(\mem[25][5] ), .A2(n2766), .B1(n6843), .B2(data_in[5]), 
        .ZN(n2771) );
  INV_X1 U1301 ( .A(n2772), .ZN(n6422) );
  AOI22_X1 U1302 ( .A1(\mem[25][6] ), .A2(n2766), .B1(n6843), .B2(data_in[6]), 
        .ZN(n2772) );
  INV_X1 U1303 ( .A(n2773), .ZN(n6421) );
  AOI22_X1 U1304 ( .A1(\mem[25][7] ), .A2(n2766), .B1(n6843), .B2(data_in[7]), 
        .ZN(n2773) );
  INV_X1 U1305 ( .A(n2774), .ZN(n6420) );
  AOI22_X1 U1306 ( .A1(\mem[26][0] ), .A2(n2775), .B1(n6842), .B2(data_in[0]), 
        .ZN(n2774) );
  INV_X1 U1307 ( .A(n2776), .ZN(n6419) );
  AOI22_X1 U1308 ( .A1(\mem[26][1] ), .A2(n2775), .B1(n6842), .B2(data_in[1]), 
        .ZN(n2776) );
  INV_X1 U1309 ( .A(n2777), .ZN(n6418) );
  AOI22_X1 U1310 ( .A1(\mem[26][2] ), .A2(n2775), .B1(n6842), .B2(data_in[2]), 
        .ZN(n2777) );
  INV_X1 U1311 ( .A(n2778), .ZN(n6417) );
  AOI22_X1 U1312 ( .A1(\mem[26][3] ), .A2(n2775), .B1(n6842), .B2(data_in[3]), 
        .ZN(n2778) );
  INV_X1 U1313 ( .A(n2779), .ZN(n6416) );
  AOI22_X1 U1314 ( .A1(\mem[26][4] ), .A2(n2775), .B1(n6842), .B2(data_in[4]), 
        .ZN(n2779) );
  INV_X1 U1315 ( .A(n2780), .ZN(n6415) );
  AOI22_X1 U1316 ( .A1(\mem[26][5] ), .A2(n2775), .B1(n6842), .B2(data_in[5]), 
        .ZN(n2780) );
  INV_X1 U1317 ( .A(n2781), .ZN(n6414) );
  AOI22_X1 U1318 ( .A1(\mem[26][6] ), .A2(n2775), .B1(n6842), .B2(data_in[6]), 
        .ZN(n2781) );
  INV_X1 U1319 ( .A(n2782), .ZN(n6413) );
  AOI22_X1 U1320 ( .A1(\mem[26][7] ), .A2(n2775), .B1(n6842), .B2(data_in[7]), 
        .ZN(n2782) );
  INV_X1 U1321 ( .A(n2783), .ZN(n6412) );
  AOI22_X1 U1322 ( .A1(\mem[27][0] ), .A2(n2784), .B1(n6841), .B2(data_in[0]), 
        .ZN(n2783) );
  INV_X1 U1323 ( .A(n2785), .ZN(n6411) );
  AOI22_X1 U1324 ( .A1(\mem[27][1] ), .A2(n2784), .B1(n6841), .B2(data_in[1]), 
        .ZN(n2785) );
  INV_X1 U1325 ( .A(n2786), .ZN(n6410) );
  AOI22_X1 U1326 ( .A1(\mem[27][2] ), .A2(n2784), .B1(n6841), .B2(data_in[2]), 
        .ZN(n2786) );
  INV_X1 U1327 ( .A(n2787), .ZN(n6409) );
  AOI22_X1 U1328 ( .A1(\mem[27][3] ), .A2(n2784), .B1(n6841), .B2(data_in[3]), 
        .ZN(n2787) );
  INV_X1 U1329 ( .A(n2788), .ZN(n6408) );
  AOI22_X1 U1330 ( .A1(\mem[27][4] ), .A2(n2784), .B1(n6841), .B2(data_in[4]), 
        .ZN(n2788) );
  INV_X1 U1331 ( .A(n2789), .ZN(n6407) );
  AOI22_X1 U1332 ( .A1(\mem[27][5] ), .A2(n2784), .B1(n6841), .B2(data_in[5]), 
        .ZN(n2789) );
  INV_X1 U1333 ( .A(n2790), .ZN(n6406) );
  AOI22_X1 U1334 ( .A1(\mem[27][6] ), .A2(n2784), .B1(n6841), .B2(data_in[6]), 
        .ZN(n2790) );
  INV_X1 U1335 ( .A(n2791), .ZN(n6405) );
  AOI22_X1 U1336 ( .A1(\mem[27][7] ), .A2(n2784), .B1(n6841), .B2(data_in[7]), 
        .ZN(n2791) );
  INV_X1 U1337 ( .A(n2792), .ZN(n6404) );
  AOI22_X1 U1338 ( .A1(\mem[28][0] ), .A2(n2793), .B1(n6840), .B2(data_in[0]), 
        .ZN(n2792) );
  INV_X1 U1339 ( .A(n2794), .ZN(n6403) );
  AOI22_X1 U1340 ( .A1(\mem[28][1] ), .A2(n2793), .B1(n6840), .B2(data_in[1]), 
        .ZN(n2794) );
  INV_X1 U1341 ( .A(n2795), .ZN(n6402) );
  AOI22_X1 U1342 ( .A1(\mem[28][2] ), .A2(n2793), .B1(n6840), .B2(data_in[2]), 
        .ZN(n2795) );
  INV_X1 U1343 ( .A(n2796), .ZN(n6401) );
  AOI22_X1 U1344 ( .A1(\mem[28][3] ), .A2(n2793), .B1(n6840), .B2(data_in[3]), 
        .ZN(n2796) );
  INV_X1 U1345 ( .A(n2797), .ZN(n6400) );
  AOI22_X1 U1346 ( .A1(\mem[28][4] ), .A2(n2793), .B1(n6840), .B2(data_in[4]), 
        .ZN(n2797) );
  INV_X1 U1347 ( .A(n2798), .ZN(n6399) );
  AOI22_X1 U1348 ( .A1(\mem[28][5] ), .A2(n2793), .B1(n6840), .B2(data_in[5]), 
        .ZN(n2798) );
  INV_X1 U1349 ( .A(n2799), .ZN(n6398) );
  AOI22_X1 U1350 ( .A1(\mem[28][6] ), .A2(n2793), .B1(n6840), .B2(data_in[6]), 
        .ZN(n2799) );
  INV_X1 U1351 ( .A(n2800), .ZN(n6397) );
  AOI22_X1 U1352 ( .A1(\mem[28][7] ), .A2(n2793), .B1(n6840), .B2(data_in[7]), 
        .ZN(n2800) );
  INV_X1 U1353 ( .A(n2801), .ZN(n6396) );
  AOI22_X1 U1354 ( .A1(\mem[29][0] ), .A2(n2802), .B1(n6839), .B2(data_in[0]), 
        .ZN(n2801) );
  INV_X1 U1355 ( .A(n2803), .ZN(n6395) );
  AOI22_X1 U1356 ( .A1(\mem[29][1] ), .A2(n2802), .B1(n6839), .B2(data_in[1]), 
        .ZN(n2803) );
  INV_X1 U1357 ( .A(n2804), .ZN(n6394) );
  AOI22_X1 U1358 ( .A1(\mem[29][2] ), .A2(n2802), .B1(n6839), .B2(data_in[2]), 
        .ZN(n2804) );
  INV_X1 U1359 ( .A(n2805), .ZN(n6393) );
  AOI22_X1 U1360 ( .A1(\mem[29][3] ), .A2(n2802), .B1(n6839), .B2(data_in[3]), 
        .ZN(n2805) );
  INV_X1 U1361 ( .A(n2806), .ZN(n6392) );
  AOI22_X1 U1362 ( .A1(\mem[29][4] ), .A2(n2802), .B1(n6839), .B2(data_in[4]), 
        .ZN(n2806) );
  INV_X1 U1363 ( .A(n2807), .ZN(n6391) );
  AOI22_X1 U1364 ( .A1(\mem[29][5] ), .A2(n2802), .B1(n6839), .B2(data_in[5]), 
        .ZN(n2807) );
  INV_X1 U1365 ( .A(n2808), .ZN(n6390) );
  AOI22_X1 U1367 ( .A1(\mem[29][6] ), .A2(n2802), .B1(n6839), .B2(data_in[6]), 
        .ZN(n2808) );
  INV_X1 U1368 ( .A(n2809), .ZN(n6389) );
  AOI22_X1 U1369 ( .A1(\mem[29][7] ), .A2(n2802), .B1(n6839), .B2(data_in[7]), 
        .ZN(n2809) );
  INV_X1 U1370 ( .A(n2810), .ZN(n6388) );
  AOI22_X1 U1371 ( .A1(\mem[30][0] ), .A2(n2811), .B1(n6838), .B2(data_in[0]), 
        .ZN(n2810) );
  INV_X1 U1372 ( .A(n2812), .ZN(n6387) );
  AOI22_X1 U1373 ( .A1(\mem[30][1] ), .A2(n2811), .B1(n6838), .B2(data_in[1]), 
        .ZN(n2812) );
  INV_X1 U1374 ( .A(n2813), .ZN(n6386) );
  AOI22_X1 U1375 ( .A1(\mem[30][2] ), .A2(n2811), .B1(n6838), .B2(data_in[2]), 
        .ZN(n2813) );
  INV_X1 U1376 ( .A(n2814), .ZN(n6385) );
  AOI22_X1 U1377 ( .A1(\mem[30][3] ), .A2(n2811), .B1(n6838), .B2(data_in[3]), 
        .ZN(n2814) );
  INV_X1 U1378 ( .A(n2815), .ZN(n6384) );
  AOI22_X1 U1379 ( .A1(\mem[30][4] ), .A2(n2811), .B1(n6838), .B2(data_in[4]), 
        .ZN(n2815) );
  INV_X1 U1380 ( .A(n2816), .ZN(n6383) );
  AOI22_X1 U1381 ( .A1(\mem[30][5] ), .A2(n2811), .B1(n6838), .B2(data_in[5]), 
        .ZN(n2816) );
  INV_X1 U1382 ( .A(n2817), .ZN(n6382) );
  AOI22_X1 U1383 ( .A1(\mem[30][6] ), .A2(n2811), .B1(n6838), .B2(data_in[6]), 
        .ZN(n2817) );
  INV_X1 U1384 ( .A(n2818), .ZN(n6381) );
  AOI22_X1 U1385 ( .A1(\mem[30][7] ), .A2(n2811), .B1(n6838), .B2(data_in[7]), 
        .ZN(n2818) );
  INV_X1 U1386 ( .A(n2819), .ZN(n6380) );
  AOI22_X1 U1387 ( .A1(\mem[31][0] ), .A2(n2820), .B1(n6837), .B2(data_in[0]), 
        .ZN(n2819) );
  INV_X1 U1388 ( .A(n2821), .ZN(n6379) );
  AOI22_X1 U1389 ( .A1(\mem[31][1] ), .A2(n2820), .B1(n6837), .B2(data_in[1]), 
        .ZN(n2821) );
  INV_X1 U1390 ( .A(n2822), .ZN(n6378) );
  AOI22_X1 U1391 ( .A1(\mem[31][2] ), .A2(n2820), .B1(n6837), .B2(data_in[2]), 
        .ZN(n2822) );
  INV_X1 U1392 ( .A(n2823), .ZN(n6377) );
  AOI22_X1 U1393 ( .A1(\mem[31][3] ), .A2(n2820), .B1(n6837), .B2(data_in[3]), 
        .ZN(n2823) );
  INV_X1 U1394 ( .A(n2824), .ZN(n6376) );
  AOI22_X1 U1395 ( .A1(\mem[31][4] ), .A2(n2820), .B1(n6837), .B2(data_in[4]), 
        .ZN(n2824) );
  INV_X1 U1396 ( .A(n2825), .ZN(n6375) );
  AOI22_X1 U1397 ( .A1(\mem[31][5] ), .A2(n2820), .B1(n6837), .B2(data_in[5]), 
        .ZN(n2825) );
  INV_X1 U1398 ( .A(n2826), .ZN(n6374) );
  AOI22_X1 U1399 ( .A1(\mem[31][6] ), .A2(n2820), .B1(n6837), .B2(data_in[6]), 
        .ZN(n2826) );
  INV_X1 U1400 ( .A(n2827), .ZN(n6373) );
  AOI22_X1 U1401 ( .A1(\mem[31][7] ), .A2(n2820), .B1(n6837), .B2(data_in[7]), 
        .ZN(n2827) );
  INV_X1 U1402 ( .A(n2829), .ZN(n6372) );
  AOI22_X1 U1403 ( .A1(\mem[32][0] ), .A2(n2830), .B1(n6836), .B2(data_in[0]), 
        .ZN(n2829) );
  INV_X1 U1404 ( .A(n2831), .ZN(n6371) );
  AOI22_X1 U1405 ( .A1(\mem[32][1] ), .A2(n2830), .B1(n6836), .B2(data_in[1]), 
        .ZN(n2831) );
  INV_X1 U1406 ( .A(n2832), .ZN(n6370) );
  AOI22_X1 U1407 ( .A1(\mem[32][2] ), .A2(n2830), .B1(n6836), .B2(data_in[2]), 
        .ZN(n2832) );
  INV_X1 U1408 ( .A(n2833), .ZN(n6369) );
  AOI22_X1 U1409 ( .A1(\mem[32][3] ), .A2(n2830), .B1(n6836), .B2(data_in[3]), 
        .ZN(n2833) );
  INV_X1 U1410 ( .A(n2834), .ZN(n6368) );
  AOI22_X1 U1411 ( .A1(\mem[32][4] ), .A2(n2830), .B1(n6836), .B2(data_in[4]), 
        .ZN(n2834) );
  INV_X1 U1412 ( .A(n2835), .ZN(n6367) );
  AOI22_X1 U1413 ( .A1(\mem[32][5] ), .A2(n2830), .B1(n6836), .B2(data_in[5]), 
        .ZN(n2835) );
  INV_X1 U1414 ( .A(n2836), .ZN(n6366) );
  AOI22_X1 U1415 ( .A1(\mem[32][6] ), .A2(n2830), .B1(n6836), .B2(data_in[6]), 
        .ZN(n2836) );
  INV_X1 U1416 ( .A(n2837), .ZN(n6365) );
  AOI22_X1 U1417 ( .A1(\mem[32][7] ), .A2(n2830), .B1(n6836), .B2(data_in[7]), 
        .ZN(n2837) );
  INV_X1 U1418 ( .A(n2839), .ZN(n6364) );
  AOI22_X1 U1419 ( .A1(\mem[33][0] ), .A2(n2840), .B1(n6835), .B2(data_in[0]), 
        .ZN(n2839) );
  INV_X1 U1420 ( .A(n2841), .ZN(n6363) );
  AOI22_X1 U1421 ( .A1(\mem[33][1] ), .A2(n2840), .B1(n6835), .B2(data_in[1]), 
        .ZN(n2841) );
  INV_X1 U1422 ( .A(n2842), .ZN(n6362) );
  AOI22_X1 U1423 ( .A1(\mem[33][2] ), .A2(n2840), .B1(n6835), .B2(data_in[2]), 
        .ZN(n2842) );
  INV_X1 U1424 ( .A(n2843), .ZN(n6361) );
  AOI22_X1 U1425 ( .A1(\mem[33][3] ), .A2(n2840), .B1(n6835), .B2(data_in[3]), 
        .ZN(n2843) );
  INV_X1 U1426 ( .A(n2844), .ZN(n6360) );
  AOI22_X1 U1427 ( .A1(\mem[33][4] ), .A2(n2840), .B1(n6835), .B2(data_in[4]), 
        .ZN(n2844) );
  INV_X1 U1428 ( .A(n2845), .ZN(n6359) );
  AOI22_X1 U1429 ( .A1(\mem[33][5] ), .A2(n2840), .B1(n6835), .B2(data_in[5]), 
        .ZN(n2845) );
  INV_X1 U1430 ( .A(n2846), .ZN(n6358) );
  AOI22_X1 U1431 ( .A1(\mem[33][6] ), .A2(n2840), .B1(n6835), .B2(data_in[6]), 
        .ZN(n2846) );
  INV_X1 U1432 ( .A(n2847), .ZN(n6357) );
  AOI22_X1 U1433 ( .A1(\mem[33][7] ), .A2(n2840), .B1(n6835), .B2(data_in[7]), 
        .ZN(n2847) );
  INV_X1 U1434 ( .A(n2848), .ZN(n6356) );
  AOI22_X1 U1435 ( .A1(\mem[34][0] ), .A2(n2849), .B1(n6834), .B2(data_in[0]), 
        .ZN(n2848) );
  INV_X1 U1436 ( .A(n2850), .ZN(n6355) );
  AOI22_X1 U1437 ( .A1(\mem[34][1] ), .A2(n2849), .B1(n6834), .B2(data_in[1]), 
        .ZN(n2850) );
  INV_X1 U1438 ( .A(n2851), .ZN(n6354) );
  AOI22_X1 U1439 ( .A1(\mem[34][2] ), .A2(n2849), .B1(n6834), .B2(data_in[2]), 
        .ZN(n2851) );
  INV_X1 U1440 ( .A(n2852), .ZN(n6353) );
  AOI22_X1 U1441 ( .A1(\mem[34][3] ), .A2(n2849), .B1(n6834), .B2(data_in[3]), 
        .ZN(n2852) );
  INV_X1 U1442 ( .A(n2853), .ZN(n6352) );
  AOI22_X1 U1443 ( .A1(\mem[34][4] ), .A2(n2849), .B1(n6834), .B2(data_in[4]), 
        .ZN(n2853) );
  INV_X1 U1444 ( .A(n2854), .ZN(n6351) );
  AOI22_X1 U1445 ( .A1(\mem[34][5] ), .A2(n2849), .B1(n6834), .B2(data_in[5]), 
        .ZN(n2854) );
  INV_X1 U1446 ( .A(n2855), .ZN(n6350) );
  AOI22_X1 U1447 ( .A1(\mem[34][6] ), .A2(n2849), .B1(n6834), .B2(data_in[6]), 
        .ZN(n2855) );
  INV_X1 U1448 ( .A(n2856), .ZN(n6349) );
  AOI22_X1 U1449 ( .A1(\mem[34][7] ), .A2(n2849), .B1(n6834), .B2(data_in[7]), 
        .ZN(n2856) );
  INV_X1 U1450 ( .A(n2857), .ZN(n6348) );
  AOI22_X1 U1451 ( .A1(\mem[35][0] ), .A2(n2858), .B1(n6833), .B2(data_in[0]), 
        .ZN(n2857) );
  INV_X1 U1452 ( .A(n2859), .ZN(n6347) );
  AOI22_X1 U1453 ( .A1(\mem[35][1] ), .A2(n2858), .B1(n6833), .B2(data_in[1]), 
        .ZN(n2859) );
  INV_X1 U1454 ( .A(n2860), .ZN(n6346) );
  AOI22_X1 U1455 ( .A1(\mem[35][2] ), .A2(n2858), .B1(n6833), .B2(data_in[2]), 
        .ZN(n2860) );
  INV_X1 U1456 ( .A(n2861), .ZN(n6345) );
  AOI22_X1 U1457 ( .A1(\mem[35][3] ), .A2(n2858), .B1(n6833), .B2(data_in[3]), 
        .ZN(n2861) );
  INV_X1 U1458 ( .A(n2862), .ZN(n6344) );
  AOI22_X1 U1459 ( .A1(\mem[35][4] ), .A2(n2858), .B1(n6833), .B2(data_in[4]), 
        .ZN(n2862) );
  INV_X1 U1460 ( .A(n2863), .ZN(n6343) );
  AOI22_X1 U1461 ( .A1(\mem[35][5] ), .A2(n2858), .B1(n6833), .B2(data_in[5]), 
        .ZN(n2863) );
  INV_X1 U1462 ( .A(n2864), .ZN(n6342) );
  AOI22_X1 U1463 ( .A1(\mem[35][6] ), .A2(n2858), .B1(n6833), .B2(data_in[6]), 
        .ZN(n2864) );
  INV_X1 U1464 ( .A(n2865), .ZN(n6341) );
  AOI22_X1 U1465 ( .A1(\mem[35][7] ), .A2(n2858), .B1(n6833), .B2(data_in[7]), 
        .ZN(n2865) );
  INV_X1 U1466 ( .A(n2866), .ZN(n6340) );
  AOI22_X1 U1467 ( .A1(\mem[36][0] ), .A2(n2867), .B1(n6832), .B2(data_in[0]), 
        .ZN(n2866) );
  INV_X1 U1468 ( .A(n2868), .ZN(n6339) );
  AOI22_X1 U1469 ( .A1(\mem[36][1] ), .A2(n2867), .B1(n6832), .B2(data_in[1]), 
        .ZN(n2868) );
  INV_X1 U1470 ( .A(n2869), .ZN(n6338) );
  AOI22_X1 U1471 ( .A1(\mem[36][2] ), .A2(n2867), .B1(n6832), .B2(data_in[2]), 
        .ZN(n2869) );
  INV_X1 U1472 ( .A(n2870), .ZN(n6337) );
  AOI22_X1 U1473 ( .A1(\mem[36][3] ), .A2(n2867), .B1(n6832), .B2(data_in[3]), 
        .ZN(n2870) );
  INV_X1 U1474 ( .A(n2871), .ZN(n6336) );
  AOI22_X1 U1475 ( .A1(\mem[36][4] ), .A2(n2867), .B1(n6832), .B2(data_in[4]), 
        .ZN(n2871) );
  INV_X1 U1476 ( .A(n2872), .ZN(n6335) );
  AOI22_X1 U1477 ( .A1(\mem[36][5] ), .A2(n2867), .B1(n6832), .B2(data_in[5]), 
        .ZN(n2872) );
  INV_X1 U1478 ( .A(n2873), .ZN(n6334) );
  AOI22_X1 U1479 ( .A1(\mem[36][6] ), .A2(n2867), .B1(n6832), .B2(data_in[6]), 
        .ZN(n2873) );
  INV_X1 U1480 ( .A(n2874), .ZN(n6333) );
  AOI22_X1 U1481 ( .A1(\mem[36][7] ), .A2(n2867), .B1(n6832), .B2(data_in[7]), 
        .ZN(n2874) );
  INV_X1 U1482 ( .A(n2875), .ZN(n6332) );
  AOI22_X1 U1483 ( .A1(\mem[37][0] ), .A2(n2876), .B1(n6831), .B2(data_in[0]), 
        .ZN(n2875) );
  INV_X1 U1484 ( .A(n2877), .ZN(n6331) );
  AOI22_X1 U1485 ( .A1(\mem[37][1] ), .A2(n2876), .B1(n6831), .B2(data_in[1]), 
        .ZN(n2877) );
  INV_X1 U1486 ( .A(n2878), .ZN(n6330) );
  AOI22_X1 U1487 ( .A1(\mem[37][2] ), .A2(n2876), .B1(n6831), .B2(data_in[2]), 
        .ZN(n2878) );
  INV_X1 U1488 ( .A(n2879), .ZN(n6329) );
  AOI22_X1 U1489 ( .A1(\mem[37][3] ), .A2(n2876), .B1(n6831), .B2(data_in[3]), 
        .ZN(n2879) );
  INV_X1 U1490 ( .A(n2880), .ZN(n6328) );
  AOI22_X1 U1491 ( .A1(\mem[37][4] ), .A2(n2876), .B1(n6831), .B2(data_in[4]), 
        .ZN(n2880) );
  INV_X1 U1492 ( .A(n2881), .ZN(n6327) );
  AOI22_X1 U1493 ( .A1(\mem[37][5] ), .A2(n2876), .B1(n6831), .B2(data_in[5]), 
        .ZN(n2881) );
  INV_X1 U1494 ( .A(n2882), .ZN(n6326) );
  AOI22_X1 U1495 ( .A1(\mem[37][6] ), .A2(n2876), .B1(n6831), .B2(data_in[6]), 
        .ZN(n2882) );
  INV_X1 U1496 ( .A(n2883), .ZN(n6325) );
  AOI22_X1 U1497 ( .A1(\mem[37][7] ), .A2(n2876), .B1(n6831), .B2(data_in[7]), 
        .ZN(n2883) );
  INV_X1 U1498 ( .A(n2884), .ZN(n6324) );
  AOI22_X1 U1499 ( .A1(\mem[38][0] ), .A2(n2885), .B1(n6830), .B2(data_in[0]), 
        .ZN(n2884) );
  INV_X1 U1500 ( .A(n2886), .ZN(n6323) );
  AOI22_X1 U1501 ( .A1(\mem[38][1] ), .A2(n2885), .B1(n6830), .B2(data_in[1]), 
        .ZN(n2886) );
  INV_X1 U1502 ( .A(n2887), .ZN(n6322) );
  AOI22_X1 U1503 ( .A1(\mem[38][2] ), .A2(n2885), .B1(n6830), .B2(data_in[2]), 
        .ZN(n2887) );
  INV_X1 U1504 ( .A(n2888), .ZN(n6321) );
  AOI22_X1 U1505 ( .A1(\mem[38][3] ), .A2(n2885), .B1(n6830), .B2(data_in[3]), 
        .ZN(n2888) );
  INV_X1 U1506 ( .A(n2889), .ZN(n6320) );
  AOI22_X1 U1507 ( .A1(\mem[38][4] ), .A2(n2885), .B1(n6830), .B2(data_in[4]), 
        .ZN(n2889) );
  INV_X1 U1508 ( .A(n2890), .ZN(n6319) );
  AOI22_X1 U1509 ( .A1(\mem[38][5] ), .A2(n2885), .B1(n6830), .B2(data_in[5]), 
        .ZN(n2890) );
  INV_X1 U1510 ( .A(n2891), .ZN(n6318) );
  AOI22_X1 U1511 ( .A1(\mem[38][6] ), .A2(n2885), .B1(n6830), .B2(data_in[6]), 
        .ZN(n2891) );
  INV_X1 U1513 ( .A(n2892), .ZN(n6317) );
  AOI22_X1 U1514 ( .A1(\mem[38][7] ), .A2(n2885), .B1(n6830), .B2(data_in[7]), 
        .ZN(n2892) );
  INV_X1 U1515 ( .A(n2893), .ZN(n6316) );
  AOI22_X1 U1516 ( .A1(\mem[39][0] ), .A2(n2894), .B1(n6829), .B2(data_in[0]), 
        .ZN(n2893) );
  INV_X1 U1517 ( .A(n2895), .ZN(n6315) );
  AOI22_X1 U1518 ( .A1(\mem[39][1] ), .A2(n2894), .B1(n6829), .B2(data_in[1]), 
        .ZN(n2895) );
  INV_X1 U1519 ( .A(n2896), .ZN(n6314) );
  AOI22_X1 U1520 ( .A1(\mem[39][2] ), .A2(n2894), .B1(n6829), .B2(data_in[2]), 
        .ZN(n2896) );
  INV_X1 U1521 ( .A(n2897), .ZN(n6313) );
  AOI22_X1 U1522 ( .A1(\mem[39][3] ), .A2(n2894), .B1(n6829), .B2(data_in[3]), 
        .ZN(n2897) );
  INV_X1 U1523 ( .A(n2898), .ZN(n6312) );
  AOI22_X1 U1524 ( .A1(\mem[39][4] ), .A2(n2894), .B1(n6829), .B2(data_in[4]), 
        .ZN(n2898) );
  INV_X1 U1525 ( .A(n2899), .ZN(n6311) );
  AOI22_X1 U1526 ( .A1(\mem[39][5] ), .A2(n2894), .B1(n6829), .B2(data_in[5]), 
        .ZN(n2899) );
  INV_X1 U1527 ( .A(n2900), .ZN(n6310) );
  AOI22_X1 U1528 ( .A1(\mem[39][6] ), .A2(n2894), .B1(n6829), .B2(data_in[6]), 
        .ZN(n2900) );
  INV_X1 U1529 ( .A(n2901), .ZN(n6309) );
  AOI22_X1 U1530 ( .A1(\mem[39][7] ), .A2(n2894), .B1(n6829), .B2(data_in[7]), 
        .ZN(n2901) );
  INV_X1 U1531 ( .A(n2902), .ZN(n6308) );
  AOI22_X1 U1532 ( .A1(\mem[40][0] ), .A2(n2903), .B1(n6828), .B2(data_in[0]), 
        .ZN(n2902) );
  INV_X1 U1533 ( .A(n2904), .ZN(n6307) );
  AOI22_X1 U1534 ( .A1(\mem[40][1] ), .A2(n2903), .B1(n6828), .B2(data_in[1]), 
        .ZN(n2904) );
  INV_X1 U1535 ( .A(n2905), .ZN(n6306) );
  AOI22_X1 U1536 ( .A1(\mem[40][2] ), .A2(n2903), .B1(n6828), .B2(data_in[2]), 
        .ZN(n2905) );
  INV_X1 U1537 ( .A(n2906), .ZN(n6305) );
  AOI22_X1 U1538 ( .A1(\mem[40][3] ), .A2(n2903), .B1(n6828), .B2(data_in[3]), 
        .ZN(n2906) );
  INV_X1 U1539 ( .A(n2907), .ZN(n6304) );
  AOI22_X1 U1540 ( .A1(\mem[40][4] ), .A2(n2903), .B1(n6828), .B2(data_in[4]), 
        .ZN(n2907) );
  INV_X1 U1541 ( .A(n2908), .ZN(n6303) );
  AOI22_X1 U1542 ( .A1(\mem[40][5] ), .A2(n2903), .B1(n6828), .B2(data_in[5]), 
        .ZN(n2908) );
  INV_X1 U1543 ( .A(n2909), .ZN(n6302) );
  AOI22_X1 U1544 ( .A1(\mem[40][6] ), .A2(n2903), .B1(n6828), .B2(data_in[6]), 
        .ZN(n2909) );
  INV_X1 U1545 ( .A(n2910), .ZN(n6301) );
  AOI22_X1 U1546 ( .A1(\mem[40][7] ), .A2(n2903), .B1(n6828), .B2(data_in[7]), 
        .ZN(n2910) );
  INV_X1 U1547 ( .A(n2911), .ZN(n6300) );
  AOI22_X1 U1548 ( .A1(\mem[41][0] ), .A2(n2912), .B1(n6827), .B2(data_in[0]), 
        .ZN(n2911) );
  INV_X1 U1549 ( .A(n2913), .ZN(n6299) );
  AOI22_X1 U1550 ( .A1(\mem[41][1] ), .A2(n2912), .B1(n6827), .B2(data_in[1]), 
        .ZN(n2913) );
  INV_X1 U1551 ( .A(n2914), .ZN(n6298) );
  AOI22_X1 U1552 ( .A1(\mem[41][2] ), .A2(n2912), .B1(n6827), .B2(data_in[2]), 
        .ZN(n2914) );
  INV_X1 U1553 ( .A(n2915), .ZN(n6297) );
  AOI22_X1 U1554 ( .A1(\mem[41][3] ), .A2(n2912), .B1(n6827), .B2(data_in[3]), 
        .ZN(n2915) );
  INV_X1 U1555 ( .A(n2916), .ZN(n6296) );
  AOI22_X1 U1556 ( .A1(\mem[41][4] ), .A2(n2912), .B1(n6827), .B2(data_in[4]), 
        .ZN(n2916) );
  INV_X1 U1557 ( .A(n2917), .ZN(n6295) );
  AOI22_X1 U1558 ( .A1(\mem[41][5] ), .A2(n2912), .B1(n6827), .B2(data_in[5]), 
        .ZN(n2917) );
  INV_X1 U1559 ( .A(n2918), .ZN(n6294) );
  AOI22_X1 U1560 ( .A1(\mem[41][6] ), .A2(n2912), .B1(n6827), .B2(data_in[6]), 
        .ZN(n2918) );
  INV_X1 U1561 ( .A(n2919), .ZN(n6293) );
  AOI22_X1 U1562 ( .A1(\mem[41][7] ), .A2(n2912), .B1(n6827), .B2(data_in[7]), 
        .ZN(n2919) );
  INV_X1 U1563 ( .A(n2920), .ZN(n6292) );
  AOI22_X1 U1564 ( .A1(\mem[42][0] ), .A2(n2921), .B1(n6826), .B2(data_in[0]), 
        .ZN(n2920) );
  INV_X1 U1565 ( .A(n2922), .ZN(n6291) );
  AOI22_X1 U1566 ( .A1(\mem[42][1] ), .A2(n2921), .B1(n6826), .B2(data_in[1]), 
        .ZN(n2922) );
  INV_X1 U1567 ( .A(n2923), .ZN(n6290) );
  AOI22_X1 U1568 ( .A1(\mem[42][2] ), .A2(n2921), .B1(n6826), .B2(data_in[2]), 
        .ZN(n2923) );
  INV_X1 U1569 ( .A(n2924), .ZN(n6289) );
  AOI22_X1 U1570 ( .A1(\mem[42][3] ), .A2(n2921), .B1(n6826), .B2(data_in[3]), 
        .ZN(n2924) );
  INV_X1 U1571 ( .A(n2925), .ZN(n6288) );
  AOI22_X1 U1572 ( .A1(\mem[42][4] ), .A2(n2921), .B1(n6826), .B2(data_in[4]), 
        .ZN(n2925) );
  INV_X1 U1573 ( .A(n2926), .ZN(n6287) );
  AOI22_X1 U1574 ( .A1(\mem[42][5] ), .A2(n2921), .B1(n6826), .B2(data_in[5]), 
        .ZN(n2926) );
  INV_X1 U1575 ( .A(n2927), .ZN(n6286) );
  AOI22_X1 U1576 ( .A1(\mem[42][6] ), .A2(n2921), .B1(n6826), .B2(data_in[6]), 
        .ZN(n2927) );
  INV_X1 U1577 ( .A(n2928), .ZN(n6285) );
  AOI22_X1 U1578 ( .A1(\mem[42][7] ), .A2(n2921), .B1(n6826), .B2(data_in[7]), 
        .ZN(n2928) );
  INV_X1 U1579 ( .A(n2929), .ZN(n6284) );
  AOI22_X1 U1580 ( .A1(\mem[43][0] ), .A2(n2930), .B1(n6825), .B2(data_in[0]), 
        .ZN(n2929) );
  INV_X1 U1581 ( .A(n2931), .ZN(n6283) );
  AOI22_X1 U1582 ( .A1(\mem[43][1] ), .A2(n2930), .B1(n6825), .B2(data_in[1]), 
        .ZN(n2931) );
  INV_X1 U1583 ( .A(n2932), .ZN(n6282) );
  AOI22_X1 U1584 ( .A1(\mem[43][2] ), .A2(n2930), .B1(n6825), .B2(data_in[2]), 
        .ZN(n2932) );
  INV_X1 U1585 ( .A(n2933), .ZN(n6281) );
  AOI22_X1 U1586 ( .A1(\mem[43][3] ), .A2(n2930), .B1(n6825), .B2(data_in[3]), 
        .ZN(n2933) );
  INV_X1 U1587 ( .A(n2934), .ZN(n6280) );
  AOI22_X1 U1588 ( .A1(\mem[43][4] ), .A2(n2930), .B1(n6825), .B2(data_in[4]), 
        .ZN(n2934) );
  INV_X1 U1589 ( .A(n2935), .ZN(n6279) );
  AOI22_X1 U1590 ( .A1(\mem[43][5] ), .A2(n2930), .B1(n6825), .B2(data_in[5]), 
        .ZN(n2935) );
  INV_X1 U1591 ( .A(n2936), .ZN(n6278) );
  AOI22_X1 U1592 ( .A1(\mem[43][6] ), .A2(n2930), .B1(n6825), .B2(data_in[6]), 
        .ZN(n2936) );
  INV_X1 U1593 ( .A(n2937), .ZN(n6277) );
  AOI22_X1 U1594 ( .A1(\mem[43][7] ), .A2(n2930), .B1(n6825), .B2(data_in[7]), 
        .ZN(n2937) );
  INV_X1 U1595 ( .A(n2938), .ZN(n6276) );
  AOI22_X1 U1596 ( .A1(\mem[44][0] ), .A2(n2939), .B1(n6824), .B2(data_in[0]), 
        .ZN(n2938) );
  INV_X1 U1597 ( .A(n2940), .ZN(n6275) );
  AOI22_X1 U1598 ( .A1(\mem[44][1] ), .A2(n2939), .B1(n6824), .B2(data_in[1]), 
        .ZN(n2940) );
  INV_X1 U1599 ( .A(n2941), .ZN(n6274) );
  AOI22_X1 U1600 ( .A1(\mem[44][2] ), .A2(n2939), .B1(n6824), .B2(data_in[2]), 
        .ZN(n2941) );
  INV_X1 U1601 ( .A(n2942), .ZN(n6273) );
  AOI22_X1 U1602 ( .A1(\mem[44][3] ), .A2(n2939), .B1(n6824), .B2(data_in[3]), 
        .ZN(n2942) );
  INV_X1 U1603 ( .A(n2943), .ZN(n6272) );
  AOI22_X1 U1604 ( .A1(\mem[44][4] ), .A2(n2939), .B1(n6824), .B2(data_in[4]), 
        .ZN(n2943) );
  INV_X1 U1605 ( .A(n2944), .ZN(n6271) );
  AOI22_X1 U1606 ( .A1(\mem[44][5] ), .A2(n2939), .B1(n6824), .B2(data_in[5]), 
        .ZN(n2944) );
  INV_X1 U1607 ( .A(n2945), .ZN(n6270) );
  AOI22_X1 U1608 ( .A1(\mem[44][6] ), .A2(n2939), .B1(n6824), .B2(data_in[6]), 
        .ZN(n2945) );
  INV_X1 U1609 ( .A(n2946), .ZN(n6269) );
  AOI22_X1 U1610 ( .A1(\mem[44][7] ), .A2(n2939), .B1(n6824), .B2(data_in[7]), 
        .ZN(n2946) );
  INV_X1 U1611 ( .A(n2947), .ZN(n6268) );
  AOI22_X1 U1612 ( .A1(\mem[45][0] ), .A2(n2948), .B1(n6823), .B2(data_in[0]), 
        .ZN(n2947) );
  INV_X1 U1613 ( .A(n2949), .ZN(n6267) );
  AOI22_X1 U1614 ( .A1(\mem[45][1] ), .A2(n2948), .B1(n6823), .B2(data_in[1]), 
        .ZN(n2949) );
  INV_X1 U1615 ( .A(n2950), .ZN(n6266) );
  AOI22_X1 U1616 ( .A1(\mem[45][2] ), .A2(n2948), .B1(n6823), .B2(data_in[2]), 
        .ZN(n2950) );
  INV_X1 U1617 ( .A(n2951), .ZN(n6265) );
  AOI22_X1 U1618 ( .A1(\mem[45][3] ), .A2(n2948), .B1(n6823), .B2(data_in[3]), 
        .ZN(n2951) );
  INV_X1 U1619 ( .A(n2952), .ZN(n6264) );
  AOI22_X1 U1620 ( .A1(\mem[45][4] ), .A2(n2948), .B1(n6823), .B2(data_in[4]), 
        .ZN(n2952) );
  INV_X1 U1621 ( .A(n2953), .ZN(n6263) );
  AOI22_X1 U1622 ( .A1(\mem[45][5] ), .A2(n2948), .B1(n6823), .B2(data_in[5]), 
        .ZN(n2953) );
  INV_X1 U1623 ( .A(n2954), .ZN(n6262) );
  AOI22_X1 U1624 ( .A1(\mem[45][6] ), .A2(n2948), .B1(n6823), .B2(data_in[6]), 
        .ZN(n2954) );
  INV_X1 U1625 ( .A(n2955), .ZN(n6261) );
  AOI22_X1 U1626 ( .A1(\mem[45][7] ), .A2(n2948), .B1(n6823), .B2(data_in[7]), 
        .ZN(n2955) );
  INV_X1 U1627 ( .A(n2956), .ZN(n6260) );
  AOI22_X1 U1628 ( .A1(\mem[46][0] ), .A2(n2957), .B1(n6822), .B2(data_in[0]), 
        .ZN(n2956) );
  INV_X1 U1629 ( .A(n2958), .ZN(n6259) );
  AOI22_X1 U1630 ( .A1(\mem[46][1] ), .A2(n2957), .B1(n6822), .B2(data_in[1]), 
        .ZN(n2958) );
  INV_X1 U1631 ( .A(n2959), .ZN(n6258) );
  AOI22_X1 U1632 ( .A1(\mem[46][2] ), .A2(n2957), .B1(n6822), .B2(data_in[2]), 
        .ZN(n2959) );
  INV_X1 U1633 ( .A(n2960), .ZN(n6257) );
  AOI22_X1 U1634 ( .A1(\mem[46][3] ), .A2(n2957), .B1(n6822), .B2(data_in[3]), 
        .ZN(n2960) );
  INV_X1 U1635 ( .A(n2961), .ZN(n6256) );
  AOI22_X1 U1636 ( .A1(\mem[46][4] ), .A2(n2957), .B1(n6822), .B2(data_in[4]), 
        .ZN(n2961) );
  INV_X1 U1637 ( .A(n2962), .ZN(n6255) );
  AOI22_X1 U1638 ( .A1(\mem[46][5] ), .A2(n2957), .B1(n6822), .B2(data_in[5]), 
        .ZN(n2962) );
  INV_X1 U1639 ( .A(n2963), .ZN(n6254) );
  AOI22_X1 U1640 ( .A1(\mem[46][6] ), .A2(n2957), .B1(n6822), .B2(data_in[6]), 
        .ZN(n2963) );
  INV_X1 U1641 ( .A(n2964), .ZN(n6253) );
  AOI22_X1 U1642 ( .A1(\mem[46][7] ), .A2(n2957), .B1(n6822), .B2(data_in[7]), 
        .ZN(n2964) );
  INV_X1 U1643 ( .A(n2965), .ZN(n6252) );
  AOI22_X1 U1644 ( .A1(\mem[47][0] ), .A2(n2966), .B1(n6821), .B2(data_in[0]), 
        .ZN(n2965) );
  INV_X1 U1645 ( .A(n2967), .ZN(n6251) );
  AOI22_X1 U1646 ( .A1(\mem[47][1] ), .A2(n2966), .B1(n6821), .B2(data_in[1]), 
        .ZN(n2967) );
  INV_X1 U1647 ( .A(n2968), .ZN(n6250) );
  AOI22_X1 U1648 ( .A1(\mem[47][2] ), .A2(n2966), .B1(n6821), .B2(data_in[2]), 
        .ZN(n2968) );
  INV_X1 U1649 ( .A(n2969), .ZN(n6249) );
  AOI22_X1 U1650 ( .A1(\mem[47][3] ), .A2(n2966), .B1(n6821), .B2(data_in[3]), 
        .ZN(n2969) );
  INV_X1 U1651 ( .A(n2970), .ZN(n6248) );
  AOI22_X1 U1652 ( .A1(\mem[47][4] ), .A2(n2966), .B1(n6821), .B2(data_in[4]), 
        .ZN(n2970) );
  INV_X1 U1653 ( .A(n2971), .ZN(n6247) );
  AOI22_X1 U1654 ( .A1(\mem[47][5] ), .A2(n2966), .B1(n6821), .B2(data_in[5]), 
        .ZN(n2971) );
  INV_X1 U1655 ( .A(n2972), .ZN(n6246) );
  AOI22_X1 U1656 ( .A1(\mem[47][6] ), .A2(n2966), .B1(n6821), .B2(data_in[6]), 
        .ZN(n2972) );
  INV_X1 U1658 ( .A(n2973), .ZN(n6245) );
  AOI22_X1 U1659 ( .A1(\mem[47][7] ), .A2(n2966), .B1(n6821), .B2(data_in[7]), 
        .ZN(n2973) );
  INV_X1 U1660 ( .A(n2975), .ZN(n6244) );
  AOI22_X1 U1661 ( .A1(\mem[48][0] ), .A2(n2976), .B1(n6820), .B2(data_in[0]), 
        .ZN(n2975) );
  INV_X1 U1662 ( .A(n2977), .ZN(n6243) );
  AOI22_X1 U1663 ( .A1(\mem[48][1] ), .A2(n2976), .B1(n6820), .B2(data_in[1]), 
        .ZN(n2977) );
  INV_X1 U1664 ( .A(n2978), .ZN(n6242) );
  AOI22_X1 U1665 ( .A1(\mem[48][2] ), .A2(n2976), .B1(n6820), .B2(data_in[2]), 
        .ZN(n2978) );
  INV_X1 U1666 ( .A(n2979), .ZN(n6241) );
  AOI22_X1 U1667 ( .A1(\mem[48][3] ), .A2(n2976), .B1(n6820), .B2(data_in[3]), 
        .ZN(n2979) );
  INV_X1 U1668 ( .A(n2980), .ZN(n6240) );
  AOI22_X1 U1669 ( .A1(\mem[48][4] ), .A2(n2976), .B1(n6820), .B2(data_in[4]), 
        .ZN(n2980) );
  INV_X1 U1670 ( .A(n2981), .ZN(n6239) );
  AOI22_X1 U1671 ( .A1(\mem[48][5] ), .A2(n2976), .B1(n6820), .B2(data_in[5]), 
        .ZN(n2981) );
  INV_X1 U1672 ( .A(n2982), .ZN(n6238) );
  AOI22_X1 U1673 ( .A1(\mem[48][6] ), .A2(n2976), .B1(n6820), .B2(data_in[6]), 
        .ZN(n2982) );
  INV_X1 U1674 ( .A(n2983), .ZN(n6237) );
  AOI22_X1 U1675 ( .A1(\mem[48][7] ), .A2(n2976), .B1(n6820), .B2(data_in[7]), 
        .ZN(n2983) );
  INV_X1 U1676 ( .A(n2985), .ZN(n6236) );
  AOI22_X1 U1677 ( .A1(\mem[49][0] ), .A2(n2986), .B1(n6819), .B2(data_in[0]), 
        .ZN(n2985) );
  INV_X1 U1678 ( .A(n2987), .ZN(n6235) );
  AOI22_X1 U1679 ( .A1(\mem[49][1] ), .A2(n2986), .B1(n6819), .B2(data_in[1]), 
        .ZN(n2987) );
  INV_X1 U1680 ( .A(n2988), .ZN(n6234) );
  AOI22_X1 U1681 ( .A1(\mem[49][2] ), .A2(n2986), .B1(n6819), .B2(data_in[2]), 
        .ZN(n2988) );
  INV_X1 U1682 ( .A(n2989), .ZN(n6233) );
  AOI22_X1 U1683 ( .A1(\mem[49][3] ), .A2(n2986), .B1(n6819), .B2(data_in[3]), 
        .ZN(n2989) );
  INV_X1 U1684 ( .A(n2990), .ZN(n6232) );
  AOI22_X1 U1685 ( .A1(\mem[49][4] ), .A2(n2986), .B1(n6819), .B2(data_in[4]), 
        .ZN(n2990) );
  INV_X1 U1686 ( .A(n2991), .ZN(n6231) );
  AOI22_X1 U1687 ( .A1(\mem[49][5] ), .A2(n2986), .B1(n6819), .B2(data_in[5]), 
        .ZN(n2991) );
  INV_X1 U1688 ( .A(n2992), .ZN(n6230) );
  AOI22_X1 U1689 ( .A1(\mem[49][6] ), .A2(n2986), .B1(n6819), .B2(data_in[6]), 
        .ZN(n2992) );
  INV_X1 U1690 ( .A(n2993), .ZN(n6229) );
  AOI22_X1 U1691 ( .A1(\mem[49][7] ), .A2(n2986), .B1(n6819), .B2(data_in[7]), 
        .ZN(n2993) );
  INV_X1 U1692 ( .A(n2994), .ZN(n6228) );
  AOI22_X1 U1693 ( .A1(\mem[50][0] ), .A2(n2995), .B1(n6818), .B2(data_in[0]), 
        .ZN(n2994) );
  INV_X1 U1694 ( .A(n2996), .ZN(n6227) );
  AOI22_X1 U1695 ( .A1(\mem[50][1] ), .A2(n2995), .B1(n6818), .B2(data_in[1]), 
        .ZN(n2996) );
  INV_X1 U1696 ( .A(n2997), .ZN(n6226) );
  AOI22_X1 U1697 ( .A1(\mem[50][2] ), .A2(n2995), .B1(n6818), .B2(data_in[2]), 
        .ZN(n2997) );
  INV_X1 U1698 ( .A(n2998), .ZN(n6225) );
  AOI22_X1 U1699 ( .A1(\mem[50][3] ), .A2(n2995), .B1(n6818), .B2(data_in[3]), 
        .ZN(n2998) );
  INV_X1 U1700 ( .A(n2999), .ZN(n6224) );
  AOI22_X1 U1701 ( .A1(\mem[50][4] ), .A2(n2995), .B1(n6818), .B2(data_in[4]), 
        .ZN(n2999) );
  INV_X1 U1702 ( .A(n3000), .ZN(n6223) );
  AOI22_X1 U1703 ( .A1(\mem[50][5] ), .A2(n2995), .B1(n6818), .B2(data_in[5]), 
        .ZN(n3000) );
  INV_X1 U1704 ( .A(n3001), .ZN(n6222) );
  AOI22_X1 U1705 ( .A1(\mem[50][6] ), .A2(n2995), .B1(n6818), .B2(data_in[6]), 
        .ZN(n3001) );
  INV_X1 U1706 ( .A(n3002), .ZN(n6221) );
  AOI22_X1 U1707 ( .A1(\mem[50][7] ), .A2(n2995), .B1(n6818), .B2(data_in[7]), 
        .ZN(n3002) );
  INV_X1 U1708 ( .A(n3003), .ZN(n6220) );
  AOI22_X1 U1709 ( .A1(\mem[51][0] ), .A2(n3004), .B1(n6817), .B2(data_in[0]), 
        .ZN(n3003) );
  INV_X1 U1710 ( .A(n3005), .ZN(n6219) );
  AOI22_X1 U1711 ( .A1(\mem[51][1] ), .A2(n3004), .B1(n6817), .B2(data_in[1]), 
        .ZN(n3005) );
  INV_X1 U1712 ( .A(n3006), .ZN(n6218) );
  AOI22_X1 U1713 ( .A1(\mem[51][2] ), .A2(n3004), .B1(n6817), .B2(data_in[2]), 
        .ZN(n3006) );
  INV_X1 U1714 ( .A(n3007), .ZN(n6217) );
  AOI22_X1 U1715 ( .A1(\mem[51][3] ), .A2(n3004), .B1(n6817), .B2(data_in[3]), 
        .ZN(n3007) );
  INV_X1 U1716 ( .A(n3008), .ZN(n6216) );
  AOI22_X1 U1717 ( .A1(\mem[51][4] ), .A2(n3004), .B1(n6817), .B2(data_in[4]), 
        .ZN(n3008) );
  INV_X1 U1718 ( .A(n3009), .ZN(n6215) );
  AOI22_X1 U1719 ( .A1(\mem[51][5] ), .A2(n3004), .B1(n6817), .B2(data_in[5]), 
        .ZN(n3009) );
  INV_X1 U1720 ( .A(n3010), .ZN(n6214) );
  AOI22_X1 U1721 ( .A1(\mem[51][6] ), .A2(n3004), .B1(n6817), .B2(data_in[6]), 
        .ZN(n3010) );
  INV_X1 U1722 ( .A(n3011), .ZN(n6213) );
  AOI22_X1 U1723 ( .A1(\mem[51][7] ), .A2(n3004), .B1(n6817), .B2(data_in[7]), 
        .ZN(n3011) );
  INV_X1 U1724 ( .A(n3012), .ZN(n6212) );
  AOI22_X1 U1725 ( .A1(\mem[52][0] ), .A2(n3013), .B1(n6816), .B2(data_in[0]), 
        .ZN(n3012) );
  INV_X1 U1726 ( .A(n3014), .ZN(n6211) );
  AOI22_X1 U1727 ( .A1(\mem[52][1] ), .A2(n3013), .B1(n6816), .B2(data_in[1]), 
        .ZN(n3014) );
  INV_X1 U1728 ( .A(n3015), .ZN(n6210) );
  AOI22_X1 U1729 ( .A1(\mem[52][2] ), .A2(n3013), .B1(n6816), .B2(data_in[2]), 
        .ZN(n3015) );
  INV_X1 U1730 ( .A(n3016), .ZN(n6209) );
  AOI22_X1 U1731 ( .A1(\mem[52][3] ), .A2(n3013), .B1(n6816), .B2(data_in[3]), 
        .ZN(n3016) );
  INV_X1 U1732 ( .A(n3017), .ZN(n6208) );
  AOI22_X1 U1733 ( .A1(\mem[52][4] ), .A2(n3013), .B1(n6816), .B2(data_in[4]), 
        .ZN(n3017) );
  INV_X1 U1734 ( .A(n3018), .ZN(n6207) );
  AOI22_X1 U1735 ( .A1(\mem[52][5] ), .A2(n3013), .B1(n6816), .B2(data_in[5]), 
        .ZN(n3018) );
  INV_X1 U1736 ( .A(n3019), .ZN(n6206) );
  AOI22_X1 U1737 ( .A1(\mem[52][6] ), .A2(n3013), .B1(n6816), .B2(data_in[6]), 
        .ZN(n3019) );
  INV_X1 U1738 ( .A(n3020), .ZN(n6205) );
  AOI22_X1 U1739 ( .A1(\mem[52][7] ), .A2(n3013), .B1(n6816), .B2(data_in[7]), 
        .ZN(n3020) );
  INV_X1 U1740 ( .A(n3021), .ZN(n6204) );
  AOI22_X1 U1741 ( .A1(\mem[53][0] ), .A2(n3022), .B1(n6815), .B2(data_in[0]), 
        .ZN(n3021) );
  INV_X1 U1742 ( .A(n3023), .ZN(n6203) );
  AOI22_X1 U1743 ( .A1(\mem[53][1] ), .A2(n3022), .B1(n6815), .B2(data_in[1]), 
        .ZN(n3023) );
  INV_X1 U1744 ( .A(n3024), .ZN(n6202) );
  AOI22_X1 U1745 ( .A1(\mem[53][2] ), .A2(n3022), .B1(n6815), .B2(data_in[2]), 
        .ZN(n3024) );
  INV_X1 U1746 ( .A(n3025), .ZN(n6201) );
  AOI22_X1 U1747 ( .A1(\mem[53][3] ), .A2(n3022), .B1(n6815), .B2(data_in[3]), 
        .ZN(n3025) );
  INV_X1 U1748 ( .A(n3026), .ZN(n6200) );
  AOI22_X1 U1749 ( .A1(\mem[53][4] ), .A2(n3022), .B1(n6815), .B2(data_in[4]), 
        .ZN(n3026) );
  INV_X1 U1750 ( .A(n3027), .ZN(n6199) );
  AOI22_X1 U1751 ( .A1(\mem[53][5] ), .A2(n3022), .B1(n6815), .B2(data_in[5]), 
        .ZN(n3027) );
  INV_X1 U1752 ( .A(n3028), .ZN(n6198) );
  AOI22_X1 U1753 ( .A1(\mem[53][6] ), .A2(n3022), .B1(n6815), .B2(data_in[6]), 
        .ZN(n3028) );
  INV_X1 U1754 ( .A(n3029), .ZN(n6197) );
  AOI22_X1 U1755 ( .A1(\mem[53][7] ), .A2(n3022), .B1(n6815), .B2(data_in[7]), 
        .ZN(n3029) );
  INV_X1 U1756 ( .A(n3030), .ZN(n6196) );
  AOI22_X1 U1757 ( .A1(\mem[54][0] ), .A2(n3031), .B1(n6814), .B2(data_in[0]), 
        .ZN(n3030) );
  INV_X1 U1758 ( .A(n3032), .ZN(n6195) );
  AOI22_X1 U1759 ( .A1(\mem[54][1] ), .A2(n3031), .B1(n6814), .B2(data_in[1]), 
        .ZN(n3032) );
  INV_X1 U1760 ( .A(n3033), .ZN(n6194) );
  AOI22_X1 U1761 ( .A1(\mem[54][2] ), .A2(n3031), .B1(n6814), .B2(data_in[2]), 
        .ZN(n3033) );
  INV_X1 U1762 ( .A(n3034), .ZN(n6193) );
  AOI22_X1 U1763 ( .A1(\mem[54][3] ), .A2(n3031), .B1(n6814), .B2(data_in[3]), 
        .ZN(n3034) );
  INV_X1 U1764 ( .A(n3035), .ZN(n6192) );
  AOI22_X1 U1765 ( .A1(\mem[54][4] ), .A2(n3031), .B1(n6814), .B2(data_in[4]), 
        .ZN(n3035) );
  INV_X1 U1766 ( .A(n3036), .ZN(n6191) );
  AOI22_X1 U1767 ( .A1(\mem[54][5] ), .A2(n3031), .B1(n6814), .B2(data_in[5]), 
        .ZN(n3036) );
  INV_X1 U1768 ( .A(n3037), .ZN(n6190) );
  AOI22_X1 U1769 ( .A1(\mem[54][6] ), .A2(n3031), .B1(n6814), .B2(data_in[6]), 
        .ZN(n3037) );
  INV_X1 U1770 ( .A(n3038), .ZN(n6189) );
  AOI22_X1 U1771 ( .A1(\mem[54][7] ), .A2(n3031), .B1(n6814), .B2(data_in[7]), 
        .ZN(n3038) );
  INV_X1 U1772 ( .A(n3039), .ZN(n6188) );
  AOI22_X1 U1773 ( .A1(\mem[55][0] ), .A2(n3040), .B1(n6813), .B2(data_in[0]), 
        .ZN(n3039) );
  INV_X1 U1774 ( .A(n3041), .ZN(n6187) );
  AOI22_X1 U1775 ( .A1(\mem[55][1] ), .A2(n3040), .B1(n6813), .B2(data_in[1]), 
        .ZN(n3041) );
  INV_X1 U1776 ( .A(n3042), .ZN(n6186) );
  AOI22_X1 U1777 ( .A1(\mem[55][2] ), .A2(n3040), .B1(n6813), .B2(data_in[2]), 
        .ZN(n3042) );
  INV_X1 U1778 ( .A(n3043), .ZN(n6185) );
  AOI22_X1 U1779 ( .A1(\mem[55][3] ), .A2(n3040), .B1(n6813), .B2(data_in[3]), 
        .ZN(n3043) );
  INV_X1 U1780 ( .A(n3044), .ZN(n6184) );
  AOI22_X1 U1781 ( .A1(\mem[55][4] ), .A2(n3040), .B1(n6813), .B2(data_in[4]), 
        .ZN(n3044) );
  INV_X1 U1782 ( .A(n3045), .ZN(n6183) );
  AOI22_X1 U1783 ( .A1(\mem[55][5] ), .A2(n3040), .B1(n6813), .B2(data_in[5]), 
        .ZN(n3045) );
  INV_X1 U1784 ( .A(n3046), .ZN(n6182) );
  AOI22_X1 U1785 ( .A1(\mem[55][6] ), .A2(n3040), .B1(n6813), .B2(data_in[6]), 
        .ZN(n3046) );
  INV_X1 U1786 ( .A(n3047), .ZN(n6181) );
  AOI22_X1 U1787 ( .A1(\mem[55][7] ), .A2(n3040), .B1(n6813), .B2(data_in[7]), 
        .ZN(n3047) );
  INV_X1 U1788 ( .A(n3048), .ZN(n6180) );
  AOI22_X1 U1789 ( .A1(\mem[56][0] ), .A2(n3049), .B1(n6812), .B2(data_in[0]), 
        .ZN(n3048) );
  INV_X1 U1790 ( .A(n3050), .ZN(n6179) );
  AOI22_X1 U1791 ( .A1(\mem[56][1] ), .A2(n3049), .B1(n6812), .B2(data_in[1]), 
        .ZN(n3050) );
  INV_X1 U1792 ( .A(n3051), .ZN(n6178) );
  AOI22_X1 U1793 ( .A1(\mem[56][2] ), .A2(n3049), .B1(n6812), .B2(data_in[2]), 
        .ZN(n3051) );
  INV_X1 U1794 ( .A(n3052), .ZN(n6177) );
  AOI22_X1 U1795 ( .A1(\mem[56][3] ), .A2(n3049), .B1(n6812), .B2(data_in[3]), 
        .ZN(n3052) );
  INV_X1 U1796 ( .A(n3053), .ZN(n6176) );
  AOI22_X1 U1797 ( .A1(\mem[56][4] ), .A2(n3049), .B1(n6812), .B2(data_in[4]), 
        .ZN(n3053) );
  INV_X1 U1798 ( .A(n3054), .ZN(n6175) );
  AOI22_X1 U1799 ( .A1(\mem[56][5] ), .A2(n3049), .B1(n6812), .B2(data_in[5]), 
        .ZN(n3054) );
  INV_X1 U1800 ( .A(n3055), .ZN(n6174) );
  AOI22_X1 U1801 ( .A1(\mem[56][6] ), .A2(n3049), .B1(n6812), .B2(data_in[6]), 
        .ZN(n3055) );
  INV_X1 U1803 ( .A(n3056), .ZN(n6173) );
  AOI22_X1 U1804 ( .A1(\mem[56][7] ), .A2(n3049), .B1(n6812), .B2(data_in[7]), 
        .ZN(n3056) );
  INV_X1 U1805 ( .A(n3057), .ZN(n6172) );
  AOI22_X1 U1806 ( .A1(\mem[57][0] ), .A2(n3058), .B1(n6811), .B2(data_in[0]), 
        .ZN(n3057) );
  INV_X1 U1807 ( .A(n3059), .ZN(n6171) );
  AOI22_X1 U1808 ( .A1(\mem[57][1] ), .A2(n3058), .B1(n6811), .B2(data_in[1]), 
        .ZN(n3059) );
  INV_X1 U1809 ( .A(n3060), .ZN(n6170) );
  AOI22_X1 U1810 ( .A1(\mem[57][2] ), .A2(n3058), .B1(n6811), .B2(data_in[2]), 
        .ZN(n3060) );
  INV_X1 U1811 ( .A(n3061), .ZN(n6169) );
  AOI22_X1 U1812 ( .A1(\mem[57][3] ), .A2(n3058), .B1(n6811), .B2(data_in[3]), 
        .ZN(n3061) );
  INV_X1 U1813 ( .A(n3062), .ZN(n6168) );
  AOI22_X1 U1814 ( .A1(\mem[57][4] ), .A2(n3058), .B1(n6811), .B2(data_in[4]), 
        .ZN(n3062) );
  INV_X1 U1815 ( .A(n3063), .ZN(n6167) );
  AOI22_X1 U1816 ( .A1(\mem[57][5] ), .A2(n3058), .B1(n6811), .B2(data_in[5]), 
        .ZN(n3063) );
  INV_X1 U1817 ( .A(n3064), .ZN(n6166) );
  AOI22_X1 U1818 ( .A1(\mem[57][6] ), .A2(n3058), .B1(n6811), .B2(data_in[6]), 
        .ZN(n3064) );
  INV_X1 U1819 ( .A(n3065), .ZN(n6165) );
  AOI22_X1 U1820 ( .A1(\mem[57][7] ), .A2(n3058), .B1(n6811), .B2(data_in[7]), 
        .ZN(n3065) );
  INV_X1 U1821 ( .A(n3066), .ZN(n6164) );
  AOI22_X1 U1822 ( .A1(\mem[58][0] ), .A2(n3067), .B1(n6810), .B2(data_in[0]), 
        .ZN(n3066) );
  INV_X1 U1823 ( .A(n3068), .ZN(n6163) );
  AOI22_X1 U1824 ( .A1(\mem[58][1] ), .A2(n3067), .B1(n6810), .B2(data_in[1]), 
        .ZN(n3068) );
  INV_X1 U1825 ( .A(n3069), .ZN(n6162) );
  AOI22_X1 U1826 ( .A1(\mem[58][2] ), .A2(n3067), .B1(n6810), .B2(data_in[2]), 
        .ZN(n3069) );
  INV_X1 U1827 ( .A(n3070), .ZN(n6161) );
  AOI22_X1 U1828 ( .A1(\mem[58][3] ), .A2(n3067), .B1(n6810), .B2(data_in[3]), 
        .ZN(n3070) );
  INV_X1 U1829 ( .A(n3071), .ZN(n6160) );
  AOI22_X1 U1830 ( .A1(\mem[58][4] ), .A2(n3067), .B1(n6810), .B2(data_in[4]), 
        .ZN(n3071) );
  INV_X1 U1831 ( .A(n3072), .ZN(n6159) );
  AOI22_X1 U1832 ( .A1(\mem[58][5] ), .A2(n3067), .B1(n6810), .B2(data_in[5]), 
        .ZN(n3072) );
  INV_X1 U1833 ( .A(n3073), .ZN(n6158) );
  AOI22_X1 U1834 ( .A1(\mem[58][6] ), .A2(n3067), .B1(n6810), .B2(data_in[6]), 
        .ZN(n3073) );
  INV_X1 U1835 ( .A(n3074), .ZN(n6157) );
  AOI22_X1 U1836 ( .A1(\mem[58][7] ), .A2(n3067), .B1(n6810), .B2(data_in[7]), 
        .ZN(n3074) );
  INV_X1 U1837 ( .A(n3075), .ZN(n6156) );
  AOI22_X1 U1838 ( .A1(\mem[59][0] ), .A2(n3076), .B1(n6809), .B2(data_in[0]), 
        .ZN(n3075) );
  INV_X1 U1839 ( .A(n3077), .ZN(n6155) );
  AOI22_X1 U1840 ( .A1(\mem[59][1] ), .A2(n3076), .B1(n6809), .B2(data_in[1]), 
        .ZN(n3077) );
  INV_X1 U1841 ( .A(n3078), .ZN(n6154) );
  AOI22_X1 U1842 ( .A1(\mem[59][2] ), .A2(n3076), .B1(n6809), .B2(data_in[2]), 
        .ZN(n3078) );
  INV_X1 U1843 ( .A(n3079), .ZN(n6153) );
  AOI22_X1 U1844 ( .A1(\mem[59][3] ), .A2(n3076), .B1(n6809), .B2(data_in[3]), 
        .ZN(n3079) );
  INV_X1 U1845 ( .A(n3080), .ZN(n6152) );
  AOI22_X1 U1846 ( .A1(\mem[59][4] ), .A2(n3076), .B1(n6809), .B2(data_in[4]), 
        .ZN(n3080) );
  INV_X1 U1847 ( .A(n3081), .ZN(n6151) );
  AOI22_X1 U1848 ( .A1(\mem[59][5] ), .A2(n3076), .B1(n6809), .B2(data_in[5]), 
        .ZN(n3081) );
  INV_X1 U1849 ( .A(n3082), .ZN(n6150) );
  AOI22_X1 U1850 ( .A1(\mem[59][6] ), .A2(n3076), .B1(n6809), .B2(data_in[6]), 
        .ZN(n3082) );
  INV_X1 U1851 ( .A(n3083), .ZN(n6149) );
  AOI22_X1 U1852 ( .A1(\mem[59][7] ), .A2(n3076), .B1(n6809), .B2(data_in[7]), 
        .ZN(n3083) );
  INV_X1 U1853 ( .A(n3084), .ZN(n6148) );
  AOI22_X1 U1854 ( .A1(\mem[60][0] ), .A2(n3085), .B1(n6808), .B2(data_in[0]), 
        .ZN(n3084) );
  INV_X1 U1855 ( .A(n3086), .ZN(n6147) );
  AOI22_X1 U1856 ( .A1(\mem[60][1] ), .A2(n3085), .B1(n6808), .B2(data_in[1]), 
        .ZN(n3086) );
  INV_X1 U1857 ( .A(n3087), .ZN(n6146) );
  AOI22_X1 U1858 ( .A1(\mem[60][2] ), .A2(n3085), .B1(n6808), .B2(data_in[2]), 
        .ZN(n3087) );
  INV_X1 U1859 ( .A(n3088), .ZN(n6145) );
  AOI22_X1 U1860 ( .A1(\mem[60][3] ), .A2(n3085), .B1(n6808), .B2(data_in[3]), 
        .ZN(n3088) );
  INV_X1 U1861 ( .A(n3089), .ZN(n6144) );
  AOI22_X1 U1862 ( .A1(\mem[60][4] ), .A2(n3085), .B1(n6808), .B2(data_in[4]), 
        .ZN(n3089) );
  INV_X1 U1863 ( .A(n3090), .ZN(n6143) );
  AOI22_X1 U1864 ( .A1(\mem[60][5] ), .A2(n3085), .B1(n6808), .B2(data_in[5]), 
        .ZN(n3090) );
  INV_X1 U1865 ( .A(n3091), .ZN(n6142) );
  AOI22_X1 U1866 ( .A1(\mem[60][6] ), .A2(n3085), .B1(n6808), .B2(data_in[6]), 
        .ZN(n3091) );
  INV_X1 U1867 ( .A(n3092), .ZN(n6141) );
  AOI22_X1 U1868 ( .A1(\mem[60][7] ), .A2(n3085), .B1(n6808), .B2(data_in[7]), 
        .ZN(n3092) );
  INV_X1 U1869 ( .A(n3093), .ZN(n6140) );
  AOI22_X1 U1870 ( .A1(\mem[61][0] ), .A2(n3094), .B1(n6807), .B2(data_in[0]), 
        .ZN(n3093) );
  INV_X1 U1871 ( .A(n3095), .ZN(n6139) );
  AOI22_X1 U1872 ( .A1(\mem[61][1] ), .A2(n3094), .B1(n6807), .B2(data_in[1]), 
        .ZN(n3095) );
  INV_X1 U1873 ( .A(n3096), .ZN(n6138) );
  AOI22_X1 U1874 ( .A1(\mem[61][2] ), .A2(n3094), .B1(n6807), .B2(data_in[2]), 
        .ZN(n3096) );
  INV_X1 U1875 ( .A(n3097), .ZN(n6137) );
  AOI22_X1 U1876 ( .A1(\mem[61][3] ), .A2(n3094), .B1(n6807), .B2(data_in[3]), 
        .ZN(n3097) );
  INV_X1 U1877 ( .A(n3098), .ZN(n6136) );
  AOI22_X1 U1878 ( .A1(\mem[61][4] ), .A2(n3094), .B1(n6807), .B2(data_in[4]), 
        .ZN(n3098) );
  INV_X1 U1879 ( .A(n3099), .ZN(n6135) );
  AOI22_X1 U1880 ( .A1(\mem[61][5] ), .A2(n3094), .B1(n6807), .B2(data_in[5]), 
        .ZN(n3099) );
  INV_X1 U1881 ( .A(n3100), .ZN(n6134) );
  AOI22_X1 U1882 ( .A1(\mem[61][6] ), .A2(n3094), .B1(n6807), .B2(data_in[6]), 
        .ZN(n3100) );
  INV_X1 U1883 ( .A(n3101), .ZN(n6133) );
  AOI22_X1 U1884 ( .A1(\mem[61][7] ), .A2(n3094), .B1(n6807), .B2(data_in[7]), 
        .ZN(n3101) );
  INV_X1 U1885 ( .A(n3102), .ZN(n6132) );
  AOI22_X1 U1886 ( .A1(\mem[62][0] ), .A2(n3103), .B1(n6806), .B2(data_in[0]), 
        .ZN(n3102) );
  INV_X1 U1887 ( .A(n3104), .ZN(n6131) );
  AOI22_X1 U1888 ( .A1(\mem[62][1] ), .A2(n3103), .B1(n6806), .B2(data_in[1]), 
        .ZN(n3104) );
  INV_X1 U1889 ( .A(n3105), .ZN(n6130) );
  AOI22_X1 U1890 ( .A1(\mem[62][2] ), .A2(n3103), .B1(n6806), .B2(data_in[2]), 
        .ZN(n3105) );
  INV_X1 U1891 ( .A(n3106), .ZN(n6129) );
  AOI22_X1 U1892 ( .A1(\mem[62][3] ), .A2(n3103), .B1(n6806), .B2(data_in[3]), 
        .ZN(n3106) );
  INV_X1 U1893 ( .A(n3107), .ZN(n6128) );
  AOI22_X1 U1894 ( .A1(\mem[62][4] ), .A2(n3103), .B1(n6806), .B2(data_in[4]), 
        .ZN(n3107) );
  INV_X1 U1895 ( .A(n3108), .ZN(n6127) );
  AOI22_X1 U1896 ( .A1(\mem[62][5] ), .A2(n3103), .B1(n6806), .B2(data_in[5]), 
        .ZN(n3108) );
  INV_X1 U1897 ( .A(n3109), .ZN(n6126) );
  AOI22_X1 U1898 ( .A1(\mem[62][6] ), .A2(n3103), .B1(n6806), .B2(data_in[6]), 
        .ZN(n3109) );
  INV_X1 U1899 ( .A(n3110), .ZN(n6125) );
  AOI22_X1 U1900 ( .A1(\mem[62][7] ), .A2(n3103), .B1(n6806), .B2(data_in[7]), 
        .ZN(n3110) );
  INV_X1 U1901 ( .A(n3111), .ZN(n6124) );
  AOI22_X1 U1902 ( .A1(\mem[63][0] ), .A2(n3112), .B1(n6805), .B2(data_in[0]), 
        .ZN(n3111) );
  INV_X1 U1903 ( .A(n3113), .ZN(n6123) );
  AOI22_X1 U1904 ( .A1(\mem[63][1] ), .A2(n3112), .B1(n6805), .B2(data_in[1]), 
        .ZN(n3113) );
  INV_X1 U1905 ( .A(n3114), .ZN(n6122) );
  AOI22_X1 U1906 ( .A1(\mem[63][2] ), .A2(n3112), .B1(n6805), .B2(data_in[2]), 
        .ZN(n3114) );
  INV_X1 U1907 ( .A(n3115), .ZN(n6121) );
  AOI22_X1 U1908 ( .A1(\mem[63][3] ), .A2(n3112), .B1(n6805), .B2(data_in[3]), 
        .ZN(n3115) );
  INV_X1 U1909 ( .A(n3116), .ZN(n6120) );
  AOI22_X1 U1910 ( .A1(\mem[63][4] ), .A2(n3112), .B1(n6805), .B2(data_in[4]), 
        .ZN(n3116) );
  INV_X1 U1911 ( .A(n3117), .ZN(n6119) );
  AOI22_X1 U1912 ( .A1(\mem[63][5] ), .A2(n3112), .B1(n6805), .B2(data_in[5]), 
        .ZN(n3117) );
  INV_X1 U1913 ( .A(n3118), .ZN(n6118) );
  AOI22_X1 U1914 ( .A1(\mem[63][6] ), .A2(n3112), .B1(n6805), .B2(data_in[6]), 
        .ZN(n3118) );
  INV_X1 U1915 ( .A(n3119), .ZN(n6117) );
  AOI22_X1 U1916 ( .A1(\mem[63][7] ), .A2(n3112), .B1(n6805), .B2(data_in[7]), 
        .ZN(n3119) );
  INV_X1 U1917 ( .A(n3120), .ZN(n6116) );
  AOI22_X1 U1918 ( .A1(\mem[64][0] ), .A2(n3121), .B1(n6804), .B2(data_in[0]), 
        .ZN(n3120) );
  INV_X1 U1919 ( .A(n3122), .ZN(n6115) );
  AOI22_X1 U1920 ( .A1(\mem[64][1] ), .A2(n3121), .B1(n6804), .B2(data_in[1]), 
        .ZN(n3122) );
  INV_X1 U1921 ( .A(n3123), .ZN(n6114) );
  AOI22_X1 U1922 ( .A1(\mem[64][2] ), .A2(n3121), .B1(n6804), .B2(data_in[2]), 
        .ZN(n3123) );
  INV_X1 U1923 ( .A(n3124), .ZN(n6113) );
  AOI22_X1 U1924 ( .A1(\mem[64][3] ), .A2(n3121), .B1(n6804), .B2(data_in[3]), 
        .ZN(n3124) );
  INV_X1 U1925 ( .A(n3125), .ZN(n6112) );
  AOI22_X1 U1926 ( .A1(\mem[64][4] ), .A2(n3121), .B1(n6804), .B2(data_in[4]), 
        .ZN(n3125) );
  INV_X1 U1927 ( .A(n3126), .ZN(n6111) );
  AOI22_X1 U1928 ( .A1(\mem[64][5] ), .A2(n3121), .B1(n6804), .B2(data_in[5]), 
        .ZN(n3126) );
  INV_X1 U1929 ( .A(n3127), .ZN(n6110) );
  AOI22_X1 U1930 ( .A1(\mem[64][6] ), .A2(n3121), .B1(n6804), .B2(data_in[6]), 
        .ZN(n3127) );
  INV_X1 U1931 ( .A(n3128), .ZN(n6109) );
  AOI22_X1 U1932 ( .A1(\mem[64][7] ), .A2(n3121), .B1(n6804), .B2(data_in[7]), 
        .ZN(n3128) );
  INV_X1 U1933 ( .A(n3130), .ZN(n6108) );
  AOI22_X1 U1934 ( .A1(\mem[65][0] ), .A2(n3131), .B1(n6803), .B2(data_in[0]), 
        .ZN(n3130) );
  INV_X1 U1935 ( .A(n3132), .ZN(n6107) );
  AOI22_X1 U1936 ( .A1(\mem[65][1] ), .A2(n3131), .B1(n6803), .B2(data_in[1]), 
        .ZN(n3132) );
  INV_X1 U1937 ( .A(n3133), .ZN(n6106) );
  AOI22_X1 U1938 ( .A1(\mem[65][2] ), .A2(n3131), .B1(n6803), .B2(data_in[2]), 
        .ZN(n3133) );
  INV_X1 U1939 ( .A(n3134), .ZN(n6105) );
  AOI22_X1 U1940 ( .A1(\mem[65][3] ), .A2(n3131), .B1(n6803), .B2(data_in[3]), 
        .ZN(n3134) );
  INV_X1 U1941 ( .A(n3135), .ZN(n6104) );
  AOI22_X1 U1942 ( .A1(\mem[65][4] ), .A2(n3131), .B1(n6803), .B2(data_in[4]), 
        .ZN(n3135) );
  INV_X1 U1943 ( .A(n3136), .ZN(n6103) );
  AOI22_X1 U1944 ( .A1(\mem[65][5] ), .A2(n3131), .B1(n6803), .B2(data_in[5]), 
        .ZN(n3136) );
  INV_X1 U1945 ( .A(n3137), .ZN(n6102) );
  AOI22_X1 U1946 ( .A1(\mem[65][6] ), .A2(n3131), .B1(n6803), .B2(data_in[6]), 
        .ZN(n3137) );
  INV_X1 U1948 ( .A(n3138), .ZN(n6101) );
  AOI22_X1 U1949 ( .A1(\mem[65][7] ), .A2(n3131), .B1(n6803), .B2(data_in[7]), 
        .ZN(n3138) );
  INV_X1 U1950 ( .A(n3139), .ZN(n6100) );
  AOI22_X1 U1951 ( .A1(\mem[66][0] ), .A2(n3140), .B1(n6802), .B2(data_in[0]), 
        .ZN(n3139) );
  INV_X1 U1952 ( .A(n3141), .ZN(n6099) );
  AOI22_X1 U1953 ( .A1(\mem[66][1] ), .A2(n3140), .B1(n6802), .B2(data_in[1]), 
        .ZN(n3141) );
  INV_X1 U1954 ( .A(n3142), .ZN(n6098) );
  AOI22_X1 U1955 ( .A1(\mem[66][2] ), .A2(n3140), .B1(n6802), .B2(data_in[2]), 
        .ZN(n3142) );
  INV_X1 U1956 ( .A(n3143), .ZN(n6097) );
  AOI22_X1 U1957 ( .A1(\mem[66][3] ), .A2(n3140), .B1(n6802), .B2(data_in[3]), 
        .ZN(n3143) );
  INV_X1 U1958 ( .A(n3144), .ZN(n6096) );
  AOI22_X1 U1959 ( .A1(\mem[66][4] ), .A2(n3140), .B1(n6802), .B2(data_in[4]), 
        .ZN(n3144) );
  INV_X1 U1960 ( .A(n3145), .ZN(n6095) );
  AOI22_X1 U1961 ( .A1(\mem[66][5] ), .A2(n3140), .B1(n6802), .B2(data_in[5]), 
        .ZN(n3145) );
  INV_X1 U1962 ( .A(n3146), .ZN(n6094) );
  AOI22_X1 U1963 ( .A1(\mem[66][6] ), .A2(n3140), .B1(n6802), .B2(data_in[6]), 
        .ZN(n3146) );
  INV_X1 U1964 ( .A(n3147), .ZN(n6093) );
  AOI22_X1 U1965 ( .A1(\mem[66][7] ), .A2(n3140), .B1(n6802), .B2(data_in[7]), 
        .ZN(n3147) );
  INV_X1 U1966 ( .A(n3148), .ZN(n6092) );
  AOI22_X1 U1967 ( .A1(\mem[67][0] ), .A2(n3149), .B1(n6801), .B2(data_in[0]), 
        .ZN(n3148) );
  INV_X1 U1968 ( .A(n3150), .ZN(n6091) );
  AOI22_X1 U1969 ( .A1(\mem[67][1] ), .A2(n3149), .B1(n6801), .B2(data_in[1]), 
        .ZN(n3150) );
  INV_X1 U1970 ( .A(n3151), .ZN(n6090) );
  AOI22_X1 U1971 ( .A1(\mem[67][2] ), .A2(n3149), .B1(n6801), .B2(data_in[2]), 
        .ZN(n3151) );
  INV_X1 U1972 ( .A(n3152), .ZN(n6089) );
  AOI22_X1 U1973 ( .A1(\mem[67][3] ), .A2(n3149), .B1(n6801), .B2(data_in[3]), 
        .ZN(n3152) );
  INV_X1 U1974 ( .A(n3153), .ZN(n6088) );
  AOI22_X1 U1975 ( .A1(\mem[67][4] ), .A2(n3149), .B1(n6801), .B2(data_in[4]), 
        .ZN(n3153) );
  INV_X1 U1976 ( .A(n3154), .ZN(n6087) );
  AOI22_X1 U1977 ( .A1(\mem[67][5] ), .A2(n3149), .B1(n6801), .B2(data_in[5]), 
        .ZN(n3154) );
  INV_X1 U1978 ( .A(n3155), .ZN(n6086) );
  AOI22_X1 U1979 ( .A1(\mem[67][6] ), .A2(n3149), .B1(n6801), .B2(data_in[6]), 
        .ZN(n3155) );
  INV_X1 U1980 ( .A(n3156), .ZN(n6085) );
  AOI22_X1 U1981 ( .A1(\mem[67][7] ), .A2(n3149), .B1(n6801), .B2(data_in[7]), 
        .ZN(n3156) );
  INV_X1 U1982 ( .A(n3157), .ZN(n6084) );
  AOI22_X1 U1983 ( .A1(\mem[68][0] ), .A2(n3158), .B1(n6800), .B2(data_in[0]), 
        .ZN(n3157) );
  INV_X1 U1984 ( .A(n3159), .ZN(n6083) );
  AOI22_X1 U1985 ( .A1(\mem[68][1] ), .A2(n3158), .B1(n6800), .B2(data_in[1]), 
        .ZN(n3159) );
  INV_X1 U1986 ( .A(n3160), .ZN(n6082) );
  AOI22_X1 U1987 ( .A1(\mem[68][2] ), .A2(n3158), .B1(n6800), .B2(data_in[2]), 
        .ZN(n3160) );
  INV_X1 U1988 ( .A(n3161), .ZN(n6081) );
  AOI22_X1 U1989 ( .A1(\mem[68][3] ), .A2(n3158), .B1(n6800), .B2(data_in[3]), 
        .ZN(n3161) );
  INV_X1 U1990 ( .A(n3162), .ZN(n6080) );
  AOI22_X1 U1991 ( .A1(\mem[68][4] ), .A2(n3158), .B1(n6800), .B2(data_in[4]), 
        .ZN(n3162) );
  INV_X1 U1992 ( .A(n3163), .ZN(n6079) );
  AOI22_X1 U1993 ( .A1(\mem[68][5] ), .A2(n3158), .B1(n6800), .B2(data_in[5]), 
        .ZN(n3163) );
  INV_X1 U1994 ( .A(n3164), .ZN(n6078) );
  AOI22_X1 U1995 ( .A1(\mem[68][6] ), .A2(n3158), .B1(n6800), .B2(data_in[6]), 
        .ZN(n3164) );
  INV_X1 U1996 ( .A(n3165), .ZN(n6077) );
  AOI22_X1 U1997 ( .A1(\mem[68][7] ), .A2(n3158), .B1(n6800), .B2(data_in[7]), 
        .ZN(n3165) );
  INV_X1 U1998 ( .A(n3166), .ZN(n6076) );
  AOI22_X1 U1999 ( .A1(\mem[69][0] ), .A2(n3167), .B1(n6799), .B2(data_in[0]), 
        .ZN(n3166) );
  INV_X1 U2000 ( .A(n3168), .ZN(n6075) );
  AOI22_X1 U2001 ( .A1(\mem[69][1] ), .A2(n3167), .B1(n6799), .B2(data_in[1]), 
        .ZN(n3168) );
  INV_X1 U2002 ( .A(n3169), .ZN(n6074) );
  AOI22_X1 U2003 ( .A1(\mem[69][2] ), .A2(n3167), .B1(n6799), .B2(data_in[2]), 
        .ZN(n3169) );
  INV_X1 U2004 ( .A(n3170), .ZN(n6073) );
  AOI22_X1 U2005 ( .A1(\mem[69][3] ), .A2(n3167), .B1(n6799), .B2(data_in[3]), 
        .ZN(n3170) );
  INV_X1 U2006 ( .A(n3171), .ZN(n6072) );
  AOI22_X1 U2007 ( .A1(\mem[69][4] ), .A2(n3167), .B1(n6799), .B2(data_in[4]), 
        .ZN(n3171) );
  INV_X1 U2008 ( .A(n3172), .ZN(n6071) );
  AOI22_X1 U2009 ( .A1(\mem[69][5] ), .A2(n3167), .B1(n6799), .B2(data_in[5]), 
        .ZN(n3172) );
  INV_X1 U2010 ( .A(n3173), .ZN(n6070) );
  AOI22_X1 U2011 ( .A1(\mem[69][6] ), .A2(n3167), .B1(n6799), .B2(data_in[6]), 
        .ZN(n3173) );
  INV_X1 U2012 ( .A(n3174), .ZN(n6069) );
  AOI22_X1 U2013 ( .A1(\mem[69][7] ), .A2(n3167), .B1(n6799), .B2(data_in[7]), 
        .ZN(n3174) );
  INV_X1 U2014 ( .A(n3175), .ZN(n6068) );
  AOI22_X1 U2015 ( .A1(\mem[70][0] ), .A2(n3176), .B1(n6798), .B2(data_in[0]), 
        .ZN(n3175) );
  INV_X1 U2016 ( .A(n3177), .ZN(n6067) );
  AOI22_X1 U2017 ( .A1(\mem[70][1] ), .A2(n3176), .B1(n6798), .B2(data_in[1]), 
        .ZN(n3177) );
  INV_X1 U2018 ( .A(n3178), .ZN(n6066) );
  AOI22_X1 U2019 ( .A1(\mem[70][2] ), .A2(n3176), .B1(n6798), .B2(data_in[2]), 
        .ZN(n3178) );
  INV_X1 U2020 ( .A(n3179), .ZN(n6065) );
  AOI22_X1 U2021 ( .A1(\mem[70][3] ), .A2(n3176), .B1(n6798), .B2(data_in[3]), 
        .ZN(n3179) );
  INV_X1 U2022 ( .A(n3180), .ZN(n6064) );
  AOI22_X1 U2023 ( .A1(\mem[70][4] ), .A2(n3176), .B1(n6798), .B2(data_in[4]), 
        .ZN(n3180) );
  INV_X1 U2024 ( .A(n3181), .ZN(n6063) );
  AOI22_X1 U2025 ( .A1(\mem[70][5] ), .A2(n3176), .B1(n6798), .B2(data_in[5]), 
        .ZN(n3181) );
  INV_X1 U2026 ( .A(n3182), .ZN(n6062) );
  AOI22_X1 U2027 ( .A1(\mem[70][6] ), .A2(n3176), .B1(n6798), .B2(data_in[6]), 
        .ZN(n3182) );
  INV_X1 U2028 ( .A(n3183), .ZN(n6061) );
  AOI22_X1 U2029 ( .A1(\mem[70][7] ), .A2(n3176), .B1(n6798), .B2(data_in[7]), 
        .ZN(n3183) );
  INV_X1 U2030 ( .A(n3184), .ZN(n6060) );
  AOI22_X1 U2031 ( .A1(\mem[71][0] ), .A2(n3185), .B1(n6797), .B2(data_in[0]), 
        .ZN(n3184) );
  INV_X1 U2032 ( .A(n3186), .ZN(n6059) );
  AOI22_X1 U2033 ( .A1(\mem[71][1] ), .A2(n3185), .B1(n6797), .B2(data_in[1]), 
        .ZN(n3186) );
  INV_X1 U2034 ( .A(n3187), .ZN(n6058) );
  AOI22_X1 U2035 ( .A1(\mem[71][2] ), .A2(n3185), .B1(n6797), .B2(data_in[2]), 
        .ZN(n3187) );
  INV_X1 U2036 ( .A(n3188), .ZN(n6057) );
  AOI22_X1 U2037 ( .A1(\mem[71][3] ), .A2(n3185), .B1(n6797), .B2(data_in[3]), 
        .ZN(n3188) );
  INV_X1 U2038 ( .A(n3189), .ZN(n6056) );
  AOI22_X1 U2039 ( .A1(\mem[71][4] ), .A2(n3185), .B1(n6797), .B2(data_in[4]), 
        .ZN(n3189) );
  INV_X1 U2040 ( .A(n3190), .ZN(n6055) );
  AOI22_X1 U2041 ( .A1(\mem[71][5] ), .A2(n3185), .B1(n6797), .B2(data_in[5]), 
        .ZN(n3190) );
  INV_X1 U2042 ( .A(n3191), .ZN(n6054) );
  AOI22_X1 U2043 ( .A1(\mem[71][6] ), .A2(n3185), .B1(n6797), .B2(data_in[6]), 
        .ZN(n3191) );
  INV_X1 U2044 ( .A(n3192), .ZN(n6053) );
  AOI22_X1 U2045 ( .A1(\mem[71][7] ), .A2(n3185), .B1(n6797), .B2(data_in[7]), 
        .ZN(n3192) );
  INV_X1 U2046 ( .A(n3193), .ZN(n6052) );
  AOI22_X1 U2047 ( .A1(\mem[72][0] ), .A2(n3194), .B1(n6796), .B2(data_in[0]), 
        .ZN(n3193) );
  INV_X1 U2048 ( .A(n3195), .ZN(n6051) );
  AOI22_X1 U2049 ( .A1(\mem[72][1] ), .A2(n3194), .B1(n6796), .B2(data_in[1]), 
        .ZN(n3195) );
  INV_X1 U2050 ( .A(n3196), .ZN(n6050) );
  AOI22_X1 U2051 ( .A1(\mem[72][2] ), .A2(n3194), .B1(n6796), .B2(data_in[2]), 
        .ZN(n3196) );
  INV_X1 U2052 ( .A(n3197), .ZN(n6049) );
  AOI22_X1 U2053 ( .A1(\mem[72][3] ), .A2(n3194), .B1(n6796), .B2(data_in[3]), 
        .ZN(n3197) );
  INV_X1 U2054 ( .A(n3198), .ZN(n6048) );
  AOI22_X1 U2055 ( .A1(\mem[72][4] ), .A2(n3194), .B1(n6796), .B2(data_in[4]), 
        .ZN(n3198) );
  INV_X1 U2056 ( .A(n3199), .ZN(n6047) );
  AOI22_X1 U2057 ( .A1(\mem[72][5] ), .A2(n3194), .B1(n6796), .B2(data_in[5]), 
        .ZN(n3199) );
  INV_X1 U2058 ( .A(n3200), .ZN(n6046) );
  AOI22_X1 U2059 ( .A1(\mem[72][6] ), .A2(n3194), .B1(n6796), .B2(data_in[6]), 
        .ZN(n3200) );
  INV_X1 U2060 ( .A(n3201), .ZN(n6045) );
  AOI22_X1 U2061 ( .A1(\mem[72][7] ), .A2(n3194), .B1(n6796), .B2(data_in[7]), 
        .ZN(n3201) );
  INV_X1 U2062 ( .A(n3202), .ZN(n6044) );
  AOI22_X1 U2063 ( .A1(\mem[73][0] ), .A2(n3203), .B1(n6795), .B2(data_in[0]), 
        .ZN(n3202) );
  INV_X1 U2064 ( .A(n3204), .ZN(n6043) );
  AOI22_X1 U2065 ( .A1(\mem[73][1] ), .A2(n3203), .B1(n6795), .B2(data_in[1]), 
        .ZN(n3204) );
  INV_X1 U2066 ( .A(n3205), .ZN(n6042) );
  AOI22_X1 U2067 ( .A1(\mem[73][2] ), .A2(n3203), .B1(n6795), .B2(data_in[2]), 
        .ZN(n3205) );
  INV_X1 U2068 ( .A(n3206), .ZN(n6041) );
  AOI22_X1 U2069 ( .A1(\mem[73][3] ), .A2(n3203), .B1(n6795), .B2(data_in[3]), 
        .ZN(n3206) );
  INV_X1 U2070 ( .A(n3207), .ZN(n6040) );
  AOI22_X1 U2071 ( .A1(\mem[73][4] ), .A2(n3203), .B1(n6795), .B2(data_in[4]), 
        .ZN(n3207) );
  INV_X1 U2072 ( .A(n3208), .ZN(n6039) );
  AOI22_X1 U2073 ( .A1(\mem[73][5] ), .A2(n3203), .B1(n6795), .B2(data_in[5]), 
        .ZN(n3208) );
  INV_X1 U2074 ( .A(n3209), .ZN(n6038) );
  AOI22_X1 U2075 ( .A1(\mem[73][6] ), .A2(n3203), .B1(n6795), .B2(data_in[6]), 
        .ZN(n3209) );
  INV_X1 U2076 ( .A(n3210), .ZN(n6037) );
  AOI22_X1 U2077 ( .A1(\mem[73][7] ), .A2(n3203), .B1(n6795), .B2(data_in[7]), 
        .ZN(n3210) );
  INV_X1 U2078 ( .A(n3211), .ZN(n6036) );
  AOI22_X1 U2079 ( .A1(\mem[74][0] ), .A2(n3212), .B1(n6794), .B2(data_in[0]), 
        .ZN(n3211) );
  INV_X1 U2080 ( .A(n3213), .ZN(n6035) );
  AOI22_X1 U2081 ( .A1(\mem[74][1] ), .A2(n3212), .B1(n6794), .B2(data_in[1]), 
        .ZN(n3213) );
  INV_X1 U2082 ( .A(n3214), .ZN(n6034) );
  AOI22_X1 U2083 ( .A1(\mem[74][2] ), .A2(n3212), .B1(n6794), .B2(data_in[2]), 
        .ZN(n3214) );
  INV_X1 U2084 ( .A(n3215), .ZN(n6033) );
  AOI22_X1 U2085 ( .A1(\mem[74][3] ), .A2(n3212), .B1(n6794), .B2(data_in[3]), 
        .ZN(n3215) );
  INV_X1 U2086 ( .A(n3216), .ZN(n6032) );
  AOI22_X1 U2087 ( .A1(\mem[74][4] ), .A2(n3212), .B1(n6794), .B2(data_in[4]), 
        .ZN(n3216) );
  INV_X1 U2088 ( .A(n3217), .ZN(n6031) );
  AOI22_X1 U2089 ( .A1(\mem[74][5] ), .A2(n3212), .B1(n6794), .B2(data_in[5]), 
        .ZN(n3217) );
  INV_X1 U2090 ( .A(n3218), .ZN(n6030) );
  AOI22_X1 U2091 ( .A1(\mem[74][6] ), .A2(n3212), .B1(n6794), .B2(data_in[6]), 
        .ZN(n3218) );
  INV_X1 U2092 ( .A(n3219), .ZN(n6029) );
  AOI22_X1 U2093 ( .A1(\mem[74][7] ), .A2(n3212), .B1(n6794), .B2(data_in[7]), 
        .ZN(n3219) );
  INV_X1 U2095 ( .A(n3220), .ZN(n6028) );
  AOI22_X1 U2096 ( .A1(\mem[75][0] ), .A2(n3221), .B1(n6793), .B2(data_in[0]), 
        .ZN(n3220) );
  INV_X1 U2097 ( .A(n3222), .ZN(n6027) );
  AOI22_X1 U2098 ( .A1(\mem[75][1] ), .A2(n3221), .B1(n6793), .B2(data_in[1]), 
        .ZN(n3222) );
  INV_X1 U2099 ( .A(n3223), .ZN(n6026) );
  AOI22_X1 U2100 ( .A1(\mem[75][2] ), .A2(n3221), .B1(n6793), .B2(data_in[2]), 
        .ZN(n3223) );
  INV_X1 U2101 ( .A(n3224), .ZN(n6025) );
  AOI22_X1 U2102 ( .A1(\mem[75][3] ), .A2(n3221), .B1(n6793), .B2(data_in[3]), 
        .ZN(n3224) );
  INV_X1 U2103 ( .A(n3225), .ZN(n6024) );
  AOI22_X1 U2104 ( .A1(\mem[75][4] ), .A2(n3221), .B1(n6793), .B2(data_in[4]), 
        .ZN(n3225) );
  INV_X1 U2105 ( .A(n3226), .ZN(n6023) );
  AOI22_X1 U2106 ( .A1(\mem[75][5] ), .A2(n3221), .B1(n6793), .B2(data_in[5]), 
        .ZN(n3226) );
  INV_X1 U2107 ( .A(n3227), .ZN(n6022) );
  AOI22_X1 U2108 ( .A1(\mem[75][6] ), .A2(n3221), .B1(n6793), .B2(data_in[6]), 
        .ZN(n3227) );
  INV_X1 U2109 ( .A(n3228), .ZN(n6021) );
  AOI22_X1 U2110 ( .A1(\mem[75][7] ), .A2(n3221), .B1(n6793), .B2(data_in[7]), 
        .ZN(n3228) );
  INV_X1 U2111 ( .A(n3229), .ZN(n6020) );
  AOI22_X1 U2112 ( .A1(\mem[76][0] ), .A2(n3230), .B1(n6792), .B2(data_in[0]), 
        .ZN(n3229) );
  INV_X1 U2113 ( .A(n3231), .ZN(n6019) );
  AOI22_X1 U2114 ( .A1(\mem[76][1] ), .A2(n3230), .B1(n6792), .B2(data_in[1]), 
        .ZN(n3231) );
  INV_X1 U2115 ( .A(n3232), .ZN(n6018) );
  AOI22_X1 U2116 ( .A1(\mem[76][2] ), .A2(n3230), .B1(n6792), .B2(data_in[2]), 
        .ZN(n3232) );
  INV_X1 U2117 ( .A(n3233), .ZN(n6017) );
  AOI22_X1 U2118 ( .A1(\mem[76][3] ), .A2(n3230), .B1(n6792), .B2(data_in[3]), 
        .ZN(n3233) );
  INV_X1 U2119 ( .A(n3234), .ZN(n6016) );
  AOI22_X1 U2120 ( .A1(\mem[76][4] ), .A2(n3230), .B1(n6792), .B2(data_in[4]), 
        .ZN(n3234) );
  INV_X1 U2121 ( .A(n3235), .ZN(n6015) );
  AOI22_X1 U2122 ( .A1(\mem[76][5] ), .A2(n3230), .B1(n6792), .B2(data_in[5]), 
        .ZN(n3235) );
  INV_X1 U2123 ( .A(n3236), .ZN(n6014) );
  AOI22_X1 U2124 ( .A1(\mem[76][6] ), .A2(n3230), .B1(n6792), .B2(data_in[6]), 
        .ZN(n3236) );
  INV_X1 U2125 ( .A(n3237), .ZN(n6013) );
  AOI22_X1 U2126 ( .A1(\mem[76][7] ), .A2(n3230), .B1(n6792), .B2(data_in[7]), 
        .ZN(n3237) );
  INV_X1 U2127 ( .A(n3238), .ZN(n6012) );
  AOI22_X1 U2128 ( .A1(\mem[77][0] ), .A2(n3239), .B1(n6791), .B2(data_in[0]), 
        .ZN(n3238) );
  INV_X1 U2129 ( .A(n3240), .ZN(n6011) );
  AOI22_X1 U2130 ( .A1(\mem[77][1] ), .A2(n3239), .B1(n6791), .B2(data_in[1]), 
        .ZN(n3240) );
  INV_X1 U2131 ( .A(n3241), .ZN(n6010) );
  AOI22_X1 U2132 ( .A1(\mem[77][2] ), .A2(n3239), .B1(n6791), .B2(data_in[2]), 
        .ZN(n3241) );
  INV_X1 U2133 ( .A(n3242), .ZN(n6009) );
  AOI22_X1 U2134 ( .A1(\mem[77][3] ), .A2(n3239), .B1(n6791), .B2(data_in[3]), 
        .ZN(n3242) );
  INV_X1 U2135 ( .A(n3243), .ZN(n6008) );
  AOI22_X1 U2136 ( .A1(\mem[77][4] ), .A2(n3239), .B1(n6791), .B2(data_in[4]), 
        .ZN(n3243) );
  INV_X1 U2137 ( .A(n3244), .ZN(n6007) );
  AOI22_X1 U2138 ( .A1(\mem[77][5] ), .A2(n3239), .B1(n6791), .B2(data_in[5]), 
        .ZN(n3244) );
  INV_X1 U2139 ( .A(n3245), .ZN(n6006) );
  AOI22_X1 U2140 ( .A1(\mem[77][6] ), .A2(n3239), .B1(n6791), .B2(data_in[6]), 
        .ZN(n3245) );
  INV_X1 U2141 ( .A(n3246), .ZN(n6005) );
  AOI22_X1 U2142 ( .A1(\mem[77][7] ), .A2(n3239), .B1(n6791), .B2(data_in[7]), 
        .ZN(n3246) );
  INV_X1 U2143 ( .A(n3247), .ZN(n6004) );
  AOI22_X1 U2144 ( .A1(\mem[78][0] ), .A2(n3248), .B1(n6790), .B2(data_in[0]), 
        .ZN(n3247) );
  INV_X1 U2145 ( .A(n3249), .ZN(n6003) );
  AOI22_X1 U2146 ( .A1(\mem[78][1] ), .A2(n3248), .B1(n6790), .B2(data_in[1]), 
        .ZN(n3249) );
  INV_X1 U2147 ( .A(n3250), .ZN(n6002) );
  AOI22_X1 U2148 ( .A1(\mem[78][2] ), .A2(n3248), .B1(n6790), .B2(data_in[2]), 
        .ZN(n3250) );
  INV_X1 U2149 ( .A(n3251), .ZN(n6001) );
  AOI22_X1 U2150 ( .A1(\mem[78][3] ), .A2(n3248), .B1(n6790), .B2(data_in[3]), 
        .ZN(n3251) );
  INV_X1 U2151 ( .A(n3252), .ZN(n6000) );
  AOI22_X1 U2152 ( .A1(\mem[78][4] ), .A2(n3248), .B1(n6790), .B2(data_in[4]), 
        .ZN(n3252) );
  INV_X1 U2153 ( .A(n3253), .ZN(n5999) );
  AOI22_X1 U2154 ( .A1(\mem[78][5] ), .A2(n3248), .B1(n6790), .B2(data_in[5]), 
        .ZN(n3253) );
  INV_X1 U2155 ( .A(n3254), .ZN(n5998) );
  AOI22_X1 U2156 ( .A1(\mem[78][6] ), .A2(n3248), .B1(n6790), .B2(data_in[6]), 
        .ZN(n3254) );
  INV_X1 U2157 ( .A(n3255), .ZN(n5997) );
  AOI22_X1 U2158 ( .A1(\mem[78][7] ), .A2(n3248), .B1(n6790), .B2(data_in[7]), 
        .ZN(n3255) );
  INV_X1 U2159 ( .A(n3256), .ZN(n5996) );
  AOI22_X1 U2160 ( .A1(\mem[79][0] ), .A2(n3257), .B1(n6789), .B2(data_in[0]), 
        .ZN(n3256) );
  INV_X1 U2161 ( .A(n3258), .ZN(n5995) );
  AOI22_X1 U2162 ( .A1(\mem[79][1] ), .A2(n3257), .B1(n6789), .B2(data_in[1]), 
        .ZN(n3258) );
  INV_X1 U2163 ( .A(n3259), .ZN(n5994) );
  AOI22_X1 U2164 ( .A1(\mem[79][2] ), .A2(n3257), .B1(n6789), .B2(data_in[2]), 
        .ZN(n3259) );
  INV_X1 U2165 ( .A(n3260), .ZN(n5993) );
  AOI22_X1 U2166 ( .A1(\mem[79][3] ), .A2(n3257), .B1(n6789), .B2(data_in[3]), 
        .ZN(n3260) );
  INV_X1 U2167 ( .A(n3261), .ZN(n5992) );
  AOI22_X1 U2168 ( .A1(\mem[79][4] ), .A2(n3257), .B1(n6789), .B2(data_in[4]), 
        .ZN(n3261) );
  INV_X1 U2169 ( .A(n3262), .ZN(n5991) );
  AOI22_X1 U2170 ( .A1(\mem[79][5] ), .A2(n3257), .B1(n6789), .B2(data_in[5]), 
        .ZN(n3262) );
  INV_X1 U2171 ( .A(n3263), .ZN(n5990) );
  AOI22_X1 U2172 ( .A1(\mem[79][6] ), .A2(n3257), .B1(n6789), .B2(data_in[6]), 
        .ZN(n3263) );
  INV_X1 U2173 ( .A(n3264), .ZN(n5989) );
  AOI22_X1 U2174 ( .A1(\mem[79][7] ), .A2(n3257), .B1(n6789), .B2(data_in[7]), 
        .ZN(n3264) );
  INV_X1 U2175 ( .A(n3266), .ZN(n5988) );
  AOI22_X1 U2176 ( .A1(\mem[80][0] ), .A2(n3267), .B1(n6788), .B2(data_in[0]), 
        .ZN(n3266) );
  INV_X1 U2177 ( .A(n3268), .ZN(n5987) );
  AOI22_X1 U2178 ( .A1(\mem[80][1] ), .A2(n3267), .B1(n6788), .B2(data_in[1]), 
        .ZN(n3268) );
  INV_X1 U2179 ( .A(n3269), .ZN(n5986) );
  AOI22_X1 U2180 ( .A1(\mem[80][2] ), .A2(n3267), .B1(n6788), .B2(data_in[2]), 
        .ZN(n3269) );
  INV_X1 U2181 ( .A(n3270), .ZN(n5985) );
  AOI22_X1 U2182 ( .A1(\mem[80][3] ), .A2(n3267), .B1(n6788), .B2(data_in[3]), 
        .ZN(n3270) );
  INV_X1 U2183 ( .A(n3271), .ZN(n5984) );
  AOI22_X1 U2184 ( .A1(\mem[80][4] ), .A2(n3267), .B1(n6788), .B2(data_in[4]), 
        .ZN(n3271) );
  INV_X1 U2185 ( .A(n3272), .ZN(n5983) );
  AOI22_X1 U2186 ( .A1(\mem[80][5] ), .A2(n3267), .B1(n6788), .B2(data_in[5]), 
        .ZN(n3272) );
  INV_X1 U2187 ( .A(n3273), .ZN(n5982) );
  AOI22_X1 U2188 ( .A1(\mem[80][6] ), .A2(n3267), .B1(n6788), .B2(data_in[6]), 
        .ZN(n3273) );
  INV_X1 U2189 ( .A(n3274), .ZN(n5981) );
  AOI22_X1 U2190 ( .A1(\mem[80][7] ), .A2(n3267), .B1(n6788), .B2(data_in[7]), 
        .ZN(n3274) );
  INV_X1 U2191 ( .A(n3276), .ZN(n5980) );
  AOI22_X1 U2192 ( .A1(\mem[81][0] ), .A2(n3277), .B1(n6787), .B2(data_in[0]), 
        .ZN(n3276) );
  INV_X1 U2193 ( .A(n3278), .ZN(n5979) );
  AOI22_X1 U2194 ( .A1(\mem[81][1] ), .A2(n3277), .B1(n6787), .B2(data_in[1]), 
        .ZN(n3278) );
  INV_X1 U2195 ( .A(n3279), .ZN(n5978) );
  AOI22_X1 U2196 ( .A1(\mem[81][2] ), .A2(n3277), .B1(n6787), .B2(data_in[2]), 
        .ZN(n3279) );
  INV_X1 U2197 ( .A(n3280), .ZN(n5977) );
  AOI22_X1 U2198 ( .A1(\mem[81][3] ), .A2(n3277), .B1(n6787), .B2(data_in[3]), 
        .ZN(n3280) );
  INV_X1 U2199 ( .A(n3281), .ZN(n5976) );
  AOI22_X1 U2200 ( .A1(\mem[81][4] ), .A2(n3277), .B1(n6787), .B2(data_in[4]), 
        .ZN(n3281) );
  INV_X1 U2201 ( .A(n3282), .ZN(n5975) );
  AOI22_X1 U2202 ( .A1(\mem[81][5] ), .A2(n3277), .B1(n6787), .B2(data_in[5]), 
        .ZN(n3282) );
  INV_X1 U2203 ( .A(n3283), .ZN(n5974) );
  AOI22_X1 U2204 ( .A1(\mem[81][6] ), .A2(n3277), .B1(n6787), .B2(data_in[6]), 
        .ZN(n3283) );
  INV_X1 U2205 ( .A(n3284), .ZN(n5973) );
  AOI22_X1 U2206 ( .A1(\mem[81][7] ), .A2(n3277), .B1(n6787), .B2(data_in[7]), 
        .ZN(n3284) );
  INV_X1 U2207 ( .A(n3285), .ZN(n5972) );
  AOI22_X1 U2208 ( .A1(\mem[82][0] ), .A2(n3286), .B1(n6786), .B2(data_in[0]), 
        .ZN(n3285) );
  INV_X1 U2209 ( .A(n3287), .ZN(n5971) );
  AOI22_X1 U2210 ( .A1(\mem[82][1] ), .A2(n3286), .B1(n6786), .B2(data_in[1]), 
        .ZN(n3287) );
  INV_X1 U2211 ( .A(n3288), .ZN(n5970) );
  AOI22_X1 U2212 ( .A1(\mem[82][2] ), .A2(n3286), .B1(n6786), .B2(data_in[2]), 
        .ZN(n3288) );
  INV_X1 U2213 ( .A(n3289), .ZN(n5969) );
  AOI22_X1 U2214 ( .A1(\mem[82][3] ), .A2(n3286), .B1(n6786), .B2(data_in[3]), 
        .ZN(n3289) );
  INV_X1 U2215 ( .A(n3290), .ZN(n5968) );
  AOI22_X1 U2216 ( .A1(\mem[82][4] ), .A2(n3286), .B1(n6786), .B2(data_in[4]), 
        .ZN(n3290) );
  INV_X1 U2217 ( .A(n3291), .ZN(n5967) );
  AOI22_X1 U2218 ( .A1(\mem[82][5] ), .A2(n3286), .B1(n6786), .B2(data_in[5]), 
        .ZN(n3291) );
  INV_X1 U2219 ( .A(n3292), .ZN(n5966) );
  AOI22_X1 U2220 ( .A1(\mem[82][6] ), .A2(n3286), .B1(n6786), .B2(data_in[6]), 
        .ZN(n3292) );
  INV_X1 U2221 ( .A(n3293), .ZN(n5965) );
  AOI22_X1 U2222 ( .A1(\mem[82][7] ), .A2(n3286), .B1(n6786), .B2(data_in[7]), 
        .ZN(n3293) );
  INV_X1 U2223 ( .A(n3294), .ZN(n5964) );
  AOI22_X1 U2224 ( .A1(\mem[83][0] ), .A2(n3295), .B1(n6785), .B2(data_in[0]), 
        .ZN(n3294) );
  INV_X1 U2225 ( .A(n3296), .ZN(n5963) );
  AOI22_X1 U2226 ( .A1(\mem[83][1] ), .A2(n3295), .B1(n6785), .B2(data_in[1]), 
        .ZN(n3296) );
  INV_X1 U2227 ( .A(n3297), .ZN(n5962) );
  AOI22_X1 U2228 ( .A1(\mem[83][2] ), .A2(n3295), .B1(n6785), .B2(data_in[2]), 
        .ZN(n3297) );
  INV_X1 U2229 ( .A(n3298), .ZN(n5961) );
  AOI22_X1 U2230 ( .A1(\mem[83][3] ), .A2(n3295), .B1(n6785), .B2(data_in[3]), 
        .ZN(n3298) );
  INV_X1 U2231 ( .A(n3299), .ZN(n5960) );
  AOI22_X1 U2232 ( .A1(\mem[83][4] ), .A2(n3295), .B1(n6785), .B2(data_in[4]), 
        .ZN(n3299) );
  INV_X1 U2233 ( .A(n3300), .ZN(n5959) );
  AOI22_X1 U2234 ( .A1(\mem[83][5] ), .A2(n3295), .B1(n6785), .B2(data_in[5]), 
        .ZN(n3300) );
  INV_X1 U2235 ( .A(n3301), .ZN(n5958) );
  AOI22_X1 U2236 ( .A1(\mem[83][6] ), .A2(n3295), .B1(n6785), .B2(data_in[6]), 
        .ZN(n3301) );
  INV_X1 U2237 ( .A(n3302), .ZN(n5957) );
  AOI22_X1 U2238 ( .A1(\mem[83][7] ), .A2(n3295), .B1(n6785), .B2(data_in[7]), 
        .ZN(n3302) );
  INV_X1 U2239 ( .A(n3303), .ZN(n5956) );
  AOI22_X1 U2240 ( .A1(\mem[84][0] ), .A2(n3304), .B1(n6784), .B2(data_in[0]), 
        .ZN(n3303) );
  INV_X1 U2241 ( .A(n3305), .ZN(n5955) );
  AOI22_X1 U2242 ( .A1(\mem[84][1] ), .A2(n3304), .B1(n6784), .B2(data_in[1]), 
        .ZN(n3305) );
  INV_X1 U2243 ( .A(n3306), .ZN(n5954) );
  AOI22_X1 U2244 ( .A1(\mem[84][2] ), .A2(n3304), .B1(n6784), .B2(data_in[2]), 
        .ZN(n3306) );
  INV_X1 U2245 ( .A(n3307), .ZN(n5953) );
  AOI22_X1 U2246 ( .A1(\mem[84][3] ), .A2(n3304), .B1(n6784), .B2(data_in[3]), 
        .ZN(n3307) );
  INV_X1 U2248 ( .A(n3308), .ZN(n5952) );
  AOI22_X1 U2249 ( .A1(\mem[84][4] ), .A2(n3304), .B1(n6784), .B2(data_in[4]), 
        .ZN(n3308) );
  INV_X1 U2250 ( .A(n3309), .ZN(n5951) );
  AOI22_X1 U2251 ( .A1(\mem[84][5] ), .A2(n3304), .B1(n6784), .B2(data_in[5]), 
        .ZN(n3309) );
  INV_X1 U2252 ( .A(n3310), .ZN(n5950) );
  AOI22_X1 U2253 ( .A1(\mem[84][6] ), .A2(n3304), .B1(n6784), .B2(data_in[6]), 
        .ZN(n3310) );
  INV_X1 U2254 ( .A(n3311), .ZN(n5949) );
  AOI22_X1 U2255 ( .A1(\mem[84][7] ), .A2(n3304), .B1(n6784), .B2(data_in[7]), 
        .ZN(n3311) );
  INV_X1 U2256 ( .A(n3312), .ZN(n5948) );
  AOI22_X1 U2257 ( .A1(\mem[85][0] ), .A2(n3313), .B1(n6783), .B2(data_in[0]), 
        .ZN(n3312) );
  INV_X1 U2258 ( .A(n3314), .ZN(n5947) );
  AOI22_X1 U2259 ( .A1(\mem[85][1] ), .A2(n3313), .B1(n6783), .B2(data_in[1]), 
        .ZN(n3314) );
  INV_X1 U2260 ( .A(n3315), .ZN(n5946) );
  AOI22_X1 U2261 ( .A1(\mem[85][2] ), .A2(n3313), .B1(n6783), .B2(data_in[2]), 
        .ZN(n3315) );
  INV_X1 U2262 ( .A(n3316), .ZN(n5945) );
  AOI22_X1 U2263 ( .A1(\mem[85][3] ), .A2(n3313), .B1(n6783), .B2(data_in[3]), 
        .ZN(n3316) );
  INV_X1 U2264 ( .A(n3317), .ZN(n5944) );
  AOI22_X1 U2265 ( .A1(\mem[85][4] ), .A2(n3313), .B1(n6783), .B2(data_in[4]), 
        .ZN(n3317) );
  INV_X1 U2266 ( .A(n3318), .ZN(n5943) );
  AOI22_X1 U2267 ( .A1(\mem[85][5] ), .A2(n3313), .B1(n6783), .B2(data_in[5]), 
        .ZN(n3318) );
  INV_X1 U2268 ( .A(n3319), .ZN(n5942) );
  AOI22_X1 U2269 ( .A1(\mem[85][6] ), .A2(n3313), .B1(n6783), .B2(data_in[6]), 
        .ZN(n3319) );
  INV_X1 U2270 ( .A(n3320), .ZN(n5941) );
  AOI22_X1 U2271 ( .A1(\mem[85][7] ), .A2(n3313), .B1(n6783), .B2(data_in[7]), 
        .ZN(n3320) );
  INV_X1 U2272 ( .A(n3321), .ZN(n5940) );
  AOI22_X1 U2273 ( .A1(\mem[86][0] ), .A2(n3322), .B1(n6782), .B2(data_in[0]), 
        .ZN(n3321) );
  INV_X1 U2274 ( .A(n3323), .ZN(n5939) );
  AOI22_X1 U2275 ( .A1(\mem[86][1] ), .A2(n3322), .B1(n6782), .B2(data_in[1]), 
        .ZN(n3323) );
  INV_X1 U2276 ( .A(n3324), .ZN(n5938) );
  AOI22_X1 U2277 ( .A1(\mem[86][2] ), .A2(n3322), .B1(n6782), .B2(data_in[2]), 
        .ZN(n3324) );
  INV_X1 U2278 ( .A(n3325), .ZN(n5937) );
  AOI22_X1 U2279 ( .A1(\mem[86][3] ), .A2(n3322), .B1(n6782), .B2(data_in[3]), 
        .ZN(n3325) );
  INV_X1 U2280 ( .A(n3326), .ZN(n5936) );
  AOI22_X1 U2281 ( .A1(\mem[86][4] ), .A2(n3322), .B1(n6782), .B2(data_in[4]), 
        .ZN(n3326) );
  INV_X1 U2282 ( .A(n3327), .ZN(n5935) );
  AOI22_X1 U2283 ( .A1(\mem[86][5] ), .A2(n3322), .B1(n6782), .B2(data_in[5]), 
        .ZN(n3327) );
  INV_X1 U2284 ( .A(n3328), .ZN(n5934) );
  AOI22_X1 U2285 ( .A1(\mem[86][6] ), .A2(n3322), .B1(n6782), .B2(data_in[6]), 
        .ZN(n3328) );
  INV_X1 U2286 ( .A(n3329), .ZN(n5933) );
  AOI22_X1 U2287 ( .A1(\mem[86][7] ), .A2(n3322), .B1(n6782), .B2(data_in[7]), 
        .ZN(n3329) );
  INV_X1 U2288 ( .A(n3330), .ZN(n5932) );
  AOI22_X1 U2289 ( .A1(\mem[87][0] ), .A2(n3331), .B1(n6781), .B2(data_in[0]), 
        .ZN(n3330) );
  INV_X1 U2290 ( .A(n3332), .ZN(n5931) );
  AOI22_X1 U2291 ( .A1(\mem[87][1] ), .A2(n3331), .B1(n6781), .B2(data_in[1]), 
        .ZN(n3332) );
  INV_X1 U2292 ( .A(n3333), .ZN(n5930) );
  AOI22_X1 U2293 ( .A1(\mem[87][2] ), .A2(n3331), .B1(n6781), .B2(data_in[2]), 
        .ZN(n3333) );
  INV_X1 U2294 ( .A(n3334), .ZN(n5929) );
  AOI22_X1 U2295 ( .A1(\mem[87][3] ), .A2(n3331), .B1(n6781), .B2(data_in[3]), 
        .ZN(n3334) );
  INV_X1 U2296 ( .A(n3335), .ZN(n5928) );
  AOI22_X1 U2297 ( .A1(\mem[87][4] ), .A2(n3331), .B1(n6781), .B2(data_in[4]), 
        .ZN(n3335) );
  INV_X1 U2298 ( .A(n3336), .ZN(n5927) );
  AOI22_X1 U2299 ( .A1(\mem[87][5] ), .A2(n3331), .B1(n6781), .B2(data_in[5]), 
        .ZN(n3336) );
  INV_X1 U2300 ( .A(n3337), .ZN(n5926) );
  AOI22_X1 U2301 ( .A1(\mem[87][6] ), .A2(n3331), .B1(n6781), .B2(data_in[6]), 
        .ZN(n3337) );
  INV_X1 U2302 ( .A(n3338), .ZN(n5925) );
  AOI22_X1 U2303 ( .A1(\mem[87][7] ), .A2(n3331), .B1(n6781), .B2(data_in[7]), 
        .ZN(n3338) );
  INV_X1 U2304 ( .A(n3339), .ZN(n5924) );
  AOI22_X1 U2305 ( .A1(\mem[88][0] ), .A2(n3340), .B1(n6780), .B2(data_in[0]), 
        .ZN(n3339) );
  INV_X1 U2306 ( .A(n3341), .ZN(n5923) );
  AOI22_X1 U2307 ( .A1(\mem[88][1] ), .A2(n3340), .B1(n6780), .B2(data_in[1]), 
        .ZN(n3341) );
  INV_X1 U2308 ( .A(n3342), .ZN(n5922) );
  AOI22_X1 U2309 ( .A1(\mem[88][2] ), .A2(n3340), .B1(n6780), .B2(data_in[2]), 
        .ZN(n3342) );
  INV_X1 U2310 ( .A(n3343), .ZN(n5921) );
  AOI22_X1 U2311 ( .A1(\mem[88][3] ), .A2(n3340), .B1(n6780), .B2(data_in[3]), 
        .ZN(n3343) );
  INV_X1 U2312 ( .A(n3344), .ZN(n5920) );
  AOI22_X1 U2313 ( .A1(\mem[88][4] ), .A2(n3340), .B1(n6780), .B2(data_in[4]), 
        .ZN(n3344) );
  INV_X1 U2314 ( .A(n3345), .ZN(n5919) );
  AOI22_X1 U2315 ( .A1(\mem[88][5] ), .A2(n3340), .B1(n6780), .B2(data_in[5]), 
        .ZN(n3345) );
  INV_X1 U2316 ( .A(n3346), .ZN(n5918) );
  AOI22_X1 U2317 ( .A1(\mem[88][6] ), .A2(n3340), .B1(n6780), .B2(data_in[6]), 
        .ZN(n3346) );
  INV_X1 U2318 ( .A(n3347), .ZN(n5917) );
  AOI22_X1 U2319 ( .A1(\mem[88][7] ), .A2(n3340), .B1(n6780), .B2(data_in[7]), 
        .ZN(n3347) );
  INV_X1 U2320 ( .A(n3348), .ZN(n5916) );
  AOI22_X1 U2321 ( .A1(\mem[89][0] ), .A2(n3349), .B1(n6779), .B2(data_in[0]), 
        .ZN(n3348) );
  INV_X1 U2322 ( .A(n3350), .ZN(n5915) );
  AOI22_X1 U2323 ( .A1(\mem[89][1] ), .A2(n3349), .B1(n6779), .B2(data_in[1]), 
        .ZN(n3350) );
  INV_X1 U2324 ( .A(n3351), .ZN(n5914) );
  AOI22_X1 U2325 ( .A1(\mem[89][2] ), .A2(n3349), .B1(n6779), .B2(data_in[2]), 
        .ZN(n3351) );
  INV_X1 U2326 ( .A(n3352), .ZN(n5913) );
  AOI22_X1 U2327 ( .A1(\mem[89][3] ), .A2(n3349), .B1(n6779), .B2(data_in[3]), 
        .ZN(n3352) );
  INV_X1 U2328 ( .A(n3353), .ZN(n5912) );
  AOI22_X1 U2329 ( .A1(\mem[89][4] ), .A2(n3349), .B1(n6779), .B2(data_in[4]), 
        .ZN(n3353) );
  INV_X1 U2330 ( .A(n3354), .ZN(n5911) );
  AOI22_X1 U2331 ( .A1(\mem[89][5] ), .A2(n3349), .B1(n6779), .B2(data_in[5]), 
        .ZN(n3354) );
  INV_X1 U2332 ( .A(n3355), .ZN(n5910) );
  AOI22_X1 U2333 ( .A1(\mem[89][6] ), .A2(n3349), .B1(n6779), .B2(data_in[6]), 
        .ZN(n3355) );
  INV_X1 U2334 ( .A(n3356), .ZN(n5909) );
  AOI22_X1 U2335 ( .A1(\mem[89][7] ), .A2(n3349), .B1(n6779), .B2(data_in[7]), 
        .ZN(n3356) );
  INV_X1 U2336 ( .A(n3357), .ZN(n5908) );
  AOI22_X1 U2337 ( .A1(\mem[90][0] ), .A2(n3358), .B1(n6778), .B2(data_in[0]), 
        .ZN(n3357) );
  INV_X1 U2338 ( .A(n3359), .ZN(n5907) );
  AOI22_X1 U2339 ( .A1(\mem[90][1] ), .A2(n3358), .B1(n6778), .B2(data_in[1]), 
        .ZN(n3359) );
  INV_X1 U2340 ( .A(n3360), .ZN(n5906) );
  AOI22_X1 U2341 ( .A1(\mem[90][2] ), .A2(n3358), .B1(n6778), .B2(data_in[2]), 
        .ZN(n3360) );
  INV_X1 U2342 ( .A(n3361), .ZN(n5905) );
  AOI22_X1 U2343 ( .A1(\mem[90][3] ), .A2(n3358), .B1(n6778), .B2(data_in[3]), 
        .ZN(n3361) );
  INV_X1 U2344 ( .A(n3362), .ZN(n5904) );
  AOI22_X1 U2345 ( .A1(\mem[90][4] ), .A2(n3358), .B1(n6778), .B2(data_in[4]), 
        .ZN(n3362) );
  INV_X1 U2346 ( .A(n3363), .ZN(n5903) );
  AOI22_X1 U2347 ( .A1(\mem[90][5] ), .A2(n3358), .B1(n6778), .B2(data_in[5]), 
        .ZN(n3363) );
  INV_X1 U2348 ( .A(n3364), .ZN(n5902) );
  AOI22_X1 U2350 ( .A1(\mem[90][6] ), .A2(n3358), .B1(n6778), .B2(data_in[6]), 
        .ZN(n3364) );
  INV_X1 U2351 ( .A(n3365), .ZN(n5901) );
  AOI22_X1 U2352 ( .A1(\mem[90][7] ), .A2(n3358), .B1(n6778), .B2(data_in[7]), 
        .ZN(n3365) );
  INV_X1 U2353 ( .A(n3366), .ZN(n5900) );
  AOI22_X1 U2354 ( .A1(\mem[91][0] ), .A2(n3367), .B1(n6777), .B2(data_in[0]), 
        .ZN(n3366) );
  INV_X1 U2355 ( .A(n3368), .ZN(n5899) );
  AOI22_X1 U2356 ( .A1(\mem[91][1] ), .A2(n3367), .B1(n6777), .B2(data_in[1]), 
        .ZN(n3368) );
  INV_X1 U2357 ( .A(n3369), .ZN(n5898) );
  AOI22_X1 U2358 ( .A1(\mem[91][2] ), .A2(n3367), .B1(n6777), .B2(data_in[2]), 
        .ZN(n3369) );
  INV_X1 U2359 ( .A(n3370), .ZN(n5897) );
  AOI22_X1 U2360 ( .A1(\mem[91][3] ), .A2(n3367), .B1(n6777), .B2(data_in[3]), 
        .ZN(n3370) );
  INV_X1 U2361 ( .A(n3371), .ZN(n5896) );
  AOI22_X1 U2362 ( .A1(\mem[91][4] ), .A2(n3367), .B1(n6777), .B2(data_in[4]), 
        .ZN(n3371) );
  INV_X1 U2363 ( .A(n3372), .ZN(n5895) );
  AOI22_X1 U2364 ( .A1(\mem[91][5] ), .A2(n3367), .B1(n6777), .B2(data_in[5]), 
        .ZN(n3372) );
  INV_X1 U2365 ( .A(n3373), .ZN(n5894) );
  AOI22_X1 U2366 ( .A1(\mem[91][6] ), .A2(n3367), .B1(n6777), .B2(data_in[6]), 
        .ZN(n3373) );
  INV_X1 U2367 ( .A(n3374), .ZN(n5893) );
  AOI22_X1 U2368 ( .A1(\mem[91][7] ), .A2(n3367), .B1(n6777), .B2(data_in[7]), 
        .ZN(n3374) );
  INV_X1 U2369 ( .A(n3375), .ZN(n5892) );
  AOI22_X1 U2370 ( .A1(\mem[92][0] ), .A2(n3376), .B1(n6776), .B2(data_in[0]), 
        .ZN(n3375) );
  INV_X1 U2371 ( .A(n3377), .ZN(n5891) );
  AOI22_X1 U2372 ( .A1(\mem[92][1] ), .A2(n3376), .B1(n6776), .B2(data_in[1]), 
        .ZN(n3377) );
  INV_X1 U2373 ( .A(n3378), .ZN(n5890) );
  AOI22_X1 U2374 ( .A1(\mem[92][2] ), .A2(n3376), .B1(n6776), .B2(data_in[2]), 
        .ZN(n3378) );
  INV_X1 U2375 ( .A(n3379), .ZN(n5889) );
  AOI22_X1 U2376 ( .A1(\mem[92][3] ), .A2(n3376), .B1(n6776), .B2(data_in[3]), 
        .ZN(n3379) );
  INV_X1 U2377 ( .A(n3380), .ZN(n5888) );
  AOI22_X1 U2378 ( .A1(\mem[92][4] ), .A2(n3376), .B1(n6776), .B2(data_in[4]), 
        .ZN(n3380) );
  INV_X1 U2379 ( .A(n3381), .ZN(n5887) );
  AOI22_X1 U2380 ( .A1(\mem[92][5] ), .A2(n3376), .B1(n6776), .B2(data_in[5]), 
        .ZN(n3381) );
  INV_X1 U2381 ( .A(n3382), .ZN(n5886) );
  AOI22_X1 U2382 ( .A1(\mem[92][6] ), .A2(n3376), .B1(n6776), .B2(data_in[6]), 
        .ZN(n3382) );
  INV_X1 U2383 ( .A(n3383), .ZN(n5885) );
  AOI22_X1 U2384 ( .A1(\mem[92][7] ), .A2(n3376), .B1(n6776), .B2(data_in[7]), 
        .ZN(n3383) );
  INV_X1 U2385 ( .A(n3384), .ZN(n5884) );
  AOI22_X1 U2386 ( .A1(\mem[93][0] ), .A2(n3385), .B1(n6775), .B2(data_in[0]), 
        .ZN(n3384) );
  INV_X1 U2387 ( .A(n3386), .ZN(n5883) );
  AOI22_X1 U2388 ( .A1(\mem[93][1] ), .A2(n3385), .B1(n6775), .B2(data_in[1]), 
        .ZN(n3386) );
  INV_X1 U2389 ( .A(n3387), .ZN(n5882) );
  AOI22_X1 U2390 ( .A1(\mem[93][2] ), .A2(n3385), .B1(n6775), .B2(data_in[2]), 
        .ZN(n3387) );
  INV_X1 U2391 ( .A(n3388), .ZN(n5881) );
  AOI22_X1 U2392 ( .A1(\mem[93][3] ), .A2(n3385), .B1(n6775), .B2(data_in[3]), 
        .ZN(n3388) );
  INV_X1 U2393 ( .A(n3389), .ZN(n5880) );
  AOI22_X1 U2394 ( .A1(\mem[93][4] ), .A2(n3385), .B1(n6775), .B2(data_in[4]), 
        .ZN(n3389) );
  INV_X1 U2395 ( .A(n3390), .ZN(n5879) );
  AOI22_X1 U2396 ( .A1(\mem[93][5] ), .A2(n3385), .B1(n6775), .B2(data_in[5]), 
        .ZN(n3390) );
  INV_X1 U2397 ( .A(n3391), .ZN(n5878) );
  AOI22_X1 U2398 ( .A1(\mem[93][6] ), .A2(n3385), .B1(n6775), .B2(data_in[6]), 
        .ZN(n3391) );
  INV_X1 U2399 ( .A(n3392), .ZN(n5877) );
  AOI22_X1 U2400 ( .A1(\mem[93][7] ), .A2(n3385), .B1(n6775), .B2(data_in[7]), 
        .ZN(n3392) );
  INV_X1 U2401 ( .A(n3393), .ZN(n5876) );
  AOI22_X1 U2402 ( .A1(\mem[94][0] ), .A2(n3394), .B1(n6774), .B2(data_in[0]), 
        .ZN(n3393) );
  INV_X1 U2403 ( .A(n3395), .ZN(n5875) );
  AOI22_X1 U2404 ( .A1(\mem[94][1] ), .A2(n3394), .B1(n6774), .B2(data_in[1]), 
        .ZN(n3395) );
  INV_X1 U2405 ( .A(n3396), .ZN(n5874) );
  AOI22_X1 U2406 ( .A1(\mem[94][2] ), .A2(n3394), .B1(n6774), .B2(data_in[2]), 
        .ZN(n3396) );
  INV_X1 U2407 ( .A(n3397), .ZN(n5873) );
  AOI22_X1 U2408 ( .A1(\mem[94][3] ), .A2(n3394), .B1(n6774), .B2(data_in[3]), 
        .ZN(n3397) );
  INV_X1 U2409 ( .A(n3398), .ZN(n5872) );
  AOI22_X1 U2410 ( .A1(\mem[94][4] ), .A2(n3394), .B1(n6774), .B2(data_in[4]), 
        .ZN(n3398) );
  INV_X1 U2411 ( .A(n3399), .ZN(n5871) );
  AOI22_X1 U2412 ( .A1(\mem[94][5] ), .A2(n3394), .B1(n6774), .B2(data_in[5]), 
        .ZN(n3399) );
  INV_X1 U2413 ( .A(n3400), .ZN(n5870) );
  AOI22_X1 U2414 ( .A1(\mem[94][6] ), .A2(n3394), .B1(n6774), .B2(data_in[6]), 
        .ZN(n3400) );
  INV_X1 U2415 ( .A(n3401), .ZN(n5869) );
  AOI22_X1 U2416 ( .A1(\mem[94][7] ), .A2(n3394), .B1(n6774), .B2(data_in[7]), 
        .ZN(n3401) );
  INV_X1 U2417 ( .A(n3402), .ZN(n5868) );
  AOI22_X1 U2418 ( .A1(\mem[95][0] ), .A2(n3403), .B1(n6773), .B2(data_in[0]), 
        .ZN(n3402) );
  INV_X1 U2419 ( .A(n3404), .ZN(n5867) );
  AOI22_X1 U2420 ( .A1(\mem[95][1] ), .A2(n3403), .B1(n6773), .B2(data_in[1]), 
        .ZN(n3404) );
  INV_X1 U2421 ( .A(n3405), .ZN(n5866) );
  AOI22_X1 U2422 ( .A1(\mem[95][2] ), .A2(n3403), .B1(n6773), .B2(data_in[2]), 
        .ZN(n3405) );
  INV_X1 U2423 ( .A(n3406), .ZN(n5865) );
  AOI22_X1 U2424 ( .A1(\mem[95][3] ), .A2(n3403), .B1(n6773), .B2(data_in[3]), 
        .ZN(n3406) );
  INV_X1 U2425 ( .A(n3407), .ZN(n5864) );
  AOI22_X1 U2426 ( .A1(\mem[95][4] ), .A2(n3403), .B1(n6773), .B2(data_in[4]), 
        .ZN(n3407) );
  INV_X1 U2427 ( .A(n3408), .ZN(n5863) );
  AOI22_X1 U2428 ( .A1(\mem[95][5] ), .A2(n3403), .B1(n6773), .B2(data_in[5]), 
        .ZN(n3408) );
  INV_X1 U2429 ( .A(n3409), .ZN(n5862) );
  AOI22_X1 U2430 ( .A1(\mem[95][6] ), .A2(n3403), .B1(n6773), .B2(data_in[6]), 
        .ZN(n3409) );
  INV_X1 U2431 ( .A(n3410), .ZN(n5861) );
  AOI22_X1 U2432 ( .A1(\mem[95][7] ), .A2(n3403), .B1(n6773), .B2(data_in[7]), 
        .ZN(n3410) );
  INV_X1 U2433 ( .A(n3411), .ZN(n5860) );
  AOI22_X1 U2434 ( .A1(\mem[96][0] ), .A2(n3412), .B1(n6772), .B2(data_in[0]), 
        .ZN(n3411) );
  INV_X1 U2435 ( .A(n3413), .ZN(n5859) );
  AOI22_X1 U2436 ( .A1(\mem[96][1] ), .A2(n3412), .B1(n6772), .B2(data_in[1]), 
        .ZN(n3413) );
  INV_X1 U2437 ( .A(n3414), .ZN(n5858) );
  AOI22_X1 U2438 ( .A1(\mem[96][2] ), .A2(n3412), .B1(n6772), .B2(data_in[2]), 
        .ZN(n3414) );
  INV_X1 U2439 ( .A(n3415), .ZN(n5857) );
  AOI22_X1 U2440 ( .A1(\mem[96][3] ), .A2(n3412), .B1(n6772), .B2(data_in[3]), 
        .ZN(n3415) );
  INV_X1 U2441 ( .A(n3416), .ZN(n5856) );
  AOI22_X1 U2442 ( .A1(\mem[96][4] ), .A2(n3412), .B1(n6772), .B2(data_in[4]), 
        .ZN(n3416) );
  INV_X1 U2443 ( .A(n3417), .ZN(n5855) );
  AOI22_X1 U2444 ( .A1(\mem[96][5] ), .A2(n3412), .B1(n6772), .B2(data_in[5]), 
        .ZN(n3417) );
  INV_X1 U2445 ( .A(n3418), .ZN(n5854) );
  AOI22_X1 U2446 ( .A1(\mem[96][6] ), .A2(n3412), .B1(n6772), .B2(data_in[6]), 
        .ZN(n3418) );
  INV_X1 U2447 ( .A(n3419), .ZN(n5853) );
  AOI22_X1 U2448 ( .A1(\mem[96][7] ), .A2(n3412), .B1(n6772), .B2(data_in[7]), 
        .ZN(n3419) );
  INV_X1 U2449 ( .A(n3421), .ZN(n5852) );
  AOI22_X1 U2450 ( .A1(\mem[97][0] ), .A2(n3422), .B1(n6771), .B2(data_in[0]), 
        .ZN(n3421) );
  INV_X1 U2451 ( .A(n3423), .ZN(n5851) );
  AOI22_X1 U2452 ( .A1(\mem[97][1] ), .A2(n3422), .B1(n6771), .B2(data_in[1]), 
        .ZN(n3423) );
  INV_X1 U2453 ( .A(n3424), .ZN(n5850) );
  AOI22_X1 U2454 ( .A1(\mem[97][2] ), .A2(n3422), .B1(n6771), .B2(data_in[2]), 
        .ZN(n3424) );
  INV_X1 U2455 ( .A(n3425), .ZN(n5849) );
  AOI22_X1 U2456 ( .A1(\mem[97][3] ), .A2(n3422), .B1(n6771), .B2(data_in[3]), 
        .ZN(n3425) );
  INV_X1 U2457 ( .A(n3426), .ZN(n5848) );
  AOI22_X1 U2458 ( .A1(\mem[97][4] ), .A2(n3422), .B1(n6771), .B2(data_in[4]), 
        .ZN(n3426) );
  INV_X1 U2459 ( .A(n3427), .ZN(n5847) );
  AOI22_X1 U2460 ( .A1(\mem[97][5] ), .A2(n3422), .B1(n6771), .B2(data_in[5]), 
        .ZN(n3427) );
  INV_X1 U2461 ( .A(n3428), .ZN(n5846) );
  AOI22_X1 U2462 ( .A1(\mem[97][6] ), .A2(n3422), .B1(n6771), .B2(data_in[6]), 
        .ZN(n3428) );
  INV_X1 U2463 ( .A(n3429), .ZN(n5845) );
  AOI22_X1 U2464 ( .A1(\mem[97][7] ), .A2(n3422), .B1(n6771), .B2(data_in[7]), 
        .ZN(n3429) );
  INV_X1 U2465 ( .A(n3430), .ZN(n5844) );
  AOI22_X1 U2466 ( .A1(\mem[98][0] ), .A2(n3431), .B1(n6770), .B2(data_in[0]), 
        .ZN(n3430) );
  INV_X1 U2467 ( .A(n3432), .ZN(n5843) );
  AOI22_X1 U2468 ( .A1(\mem[98][1] ), .A2(n3431), .B1(n6770), .B2(data_in[1]), 
        .ZN(n3432) );
  INV_X1 U2469 ( .A(n3433), .ZN(n5842) );
  AOI22_X1 U2470 ( .A1(\mem[98][2] ), .A2(n3431), .B1(n6770), .B2(data_in[2]), 
        .ZN(n3433) );
  INV_X1 U2471 ( .A(n3434), .ZN(n5841) );
  AOI22_X1 U2472 ( .A1(\mem[98][3] ), .A2(n3431), .B1(n6770), .B2(data_in[3]), 
        .ZN(n3434) );
  INV_X1 U2473 ( .A(n3435), .ZN(n5840) );
  AOI22_X1 U2474 ( .A1(\mem[98][4] ), .A2(n3431), .B1(n6770), .B2(data_in[4]), 
        .ZN(n3435) );
  INV_X1 U2475 ( .A(n3436), .ZN(n5839) );
  AOI22_X1 U2476 ( .A1(\mem[98][5] ), .A2(n3431), .B1(n6770), .B2(data_in[5]), 
        .ZN(n3436) );
  INV_X1 U2477 ( .A(n3437), .ZN(n5838) );
  AOI22_X1 U2478 ( .A1(\mem[98][6] ), .A2(n3431), .B1(n6770), .B2(data_in[6]), 
        .ZN(n3437) );
  INV_X1 U2479 ( .A(n3438), .ZN(n5837) );
  AOI22_X1 U2480 ( .A1(\mem[98][7] ), .A2(n3431), .B1(n6770), .B2(data_in[7]), 
        .ZN(n3438) );
  INV_X1 U2481 ( .A(n3439), .ZN(n5836) );
  AOI22_X1 U2482 ( .A1(\mem[99][0] ), .A2(n3440), .B1(n6769), .B2(data_in[0]), 
        .ZN(n3439) );
  INV_X1 U2483 ( .A(n3441), .ZN(n5835) );
  AOI22_X1 U2484 ( .A1(\mem[99][1] ), .A2(n3440), .B1(n6769), .B2(data_in[1]), 
        .ZN(n3441) );
  INV_X1 U2485 ( .A(n3442), .ZN(n5834) );
  AOI22_X1 U2486 ( .A1(\mem[99][2] ), .A2(n3440), .B1(n6769), .B2(data_in[2]), 
        .ZN(n3442) );
  INV_X1 U2487 ( .A(n3443), .ZN(n5833) );
  AOI22_X1 U2488 ( .A1(\mem[99][3] ), .A2(n3440), .B1(n6769), .B2(data_in[3]), 
        .ZN(n3443) );
  INV_X1 U2489 ( .A(n3444), .ZN(n5832) );
  AOI22_X1 U2490 ( .A1(\mem[99][4] ), .A2(n3440), .B1(n6769), .B2(data_in[4]), 
        .ZN(n3444) );
  INV_X1 U2491 ( .A(n3445), .ZN(n5831) );
  AOI22_X1 U2492 ( .A1(\mem[99][5] ), .A2(n3440), .B1(n6769), .B2(data_in[5]), 
        .ZN(n3445) );
  INV_X1 U2493 ( .A(n3446), .ZN(n5830) );
  AOI22_X1 U2494 ( .A1(\mem[99][6] ), .A2(n3440), .B1(n6769), .B2(data_in[6]), 
        .ZN(n3446) );
  INV_X1 U2495 ( .A(n3447), .ZN(n5829) );
  AOI22_X1 U2496 ( .A1(\mem[99][7] ), .A2(n3440), .B1(n6769), .B2(data_in[7]), 
        .ZN(n3447) );
  INV_X1 U2497 ( .A(n3448), .ZN(n5828) );
  AOI22_X1 U2498 ( .A1(\mem[100][0] ), .A2(n3449), .B1(n6768), .B2(data_in[0]), 
        .ZN(n3448) );
  INV_X1 U2499 ( .A(n3450), .ZN(n5827) );
  AOI22_X1 U2500 ( .A1(\mem[100][1] ), .A2(n3449), .B1(n6768), .B2(data_in[1]), 
        .ZN(n3450) );
  INV_X1 U2501 ( .A(n3451), .ZN(n5826) );
  AOI22_X1 U2502 ( .A1(\mem[100][2] ), .A2(n3449), .B1(n6768), .B2(data_in[2]), 
        .ZN(n3451) );
  INV_X1 U2503 ( .A(n3452), .ZN(n5825) );
  AOI22_X1 U2504 ( .A1(\mem[100][3] ), .A2(n3449), .B1(n6768), .B2(data_in[3]), 
        .ZN(n3452) );
  INV_X1 U2505 ( .A(n3453), .ZN(n5824) );
  AOI22_X1 U2506 ( .A1(\mem[100][4] ), .A2(n3449), .B1(n6768), .B2(data_in[4]), 
        .ZN(n3453) );
  INV_X1 U2507 ( .A(n3454), .ZN(n5823) );
  AOI22_X1 U2508 ( .A1(\mem[100][5] ), .A2(n3449), .B1(n6768), .B2(data_in[5]), 
        .ZN(n3454) );
  INV_X1 U2509 ( .A(n3455), .ZN(n5822) );
  AOI22_X1 U2510 ( .A1(\mem[100][6] ), .A2(n3449), .B1(n6768), .B2(data_in[6]), 
        .ZN(n3455) );
  INV_X1 U2511 ( .A(n3456), .ZN(n5821) );
  AOI22_X1 U2512 ( .A1(\mem[100][7] ), .A2(n3449), .B1(n6768), .B2(data_in[7]), 
        .ZN(n3456) );
  INV_X1 U2513 ( .A(n3457), .ZN(n5820) );
  AOI22_X1 U2514 ( .A1(\mem[101][0] ), .A2(n3458), .B1(n6767), .B2(data_in[0]), 
        .ZN(n3457) );
  INV_X1 U2515 ( .A(n3459), .ZN(n5819) );
  AOI22_X1 U2516 ( .A1(\mem[101][1] ), .A2(n3458), .B1(n6767), .B2(data_in[1]), 
        .ZN(n3459) );
  INV_X1 U2517 ( .A(n3460), .ZN(n5818) );
  AOI22_X1 U2518 ( .A1(\mem[101][2] ), .A2(n3458), .B1(n6767), .B2(data_in[2]), 
        .ZN(n3460) );
  INV_X1 U2519 ( .A(n3461), .ZN(n5817) );
  AOI22_X1 U2520 ( .A1(\mem[101][3] ), .A2(n3458), .B1(n6767), .B2(data_in[3]), 
        .ZN(n3461) );
  INV_X1 U2521 ( .A(n3462), .ZN(n5816) );
  AOI22_X1 U2522 ( .A1(\mem[101][4] ), .A2(n3458), .B1(n6767), .B2(data_in[4]), 
        .ZN(n3462) );
  INV_X1 U2523 ( .A(n3463), .ZN(n5815) );
  AOI22_X1 U2524 ( .A1(\mem[101][5] ), .A2(n3458), .B1(n6767), .B2(data_in[5]), 
        .ZN(n3463) );
  INV_X1 U2525 ( .A(n3464), .ZN(n5814) );
  AOI22_X1 U2526 ( .A1(\mem[101][6] ), .A2(n3458), .B1(n6767), .B2(data_in[6]), 
        .ZN(n3464) );
  INV_X1 U2527 ( .A(n3465), .ZN(n5813) );
  AOI22_X1 U2528 ( .A1(\mem[101][7] ), .A2(n3458), .B1(n6767), .B2(data_in[7]), 
        .ZN(n3465) );
  INV_X1 U2529 ( .A(n3466), .ZN(n5812) );
  AOI22_X1 U2530 ( .A1(\mem[102][0] ), .A2(n3467), .B1(n6766), .B2(data_in[0]), 
        .ZN(n3466) );
  INV_X1 U2531 ( .A(n3468), .ZN(n5811) );
  AOI22_X1 U2532 ( .A1(\mem[102][1] ), .A2(n3467), .B1(n6766), .B2(data_in[1]), 
        .ZN(n3468) );
  INV_X1 U2533 ( .A(n3469), .ZN(n5810) );
  AOI22_X1 U2534 ( .A1(\mem[102][2] ), .A2(n3467), .B1(n6766), .B2(data_in[2]), 
        .ZN(n3469) );
  INV_X1 U2535 ( .A(n3470), .ZN(n5809) );
  AOI22_X1 U2536 ( .A1(\mem[102][3] ), .A2(n3467), .B1(n6766), .B2(data_in[3]), 
        .ZN(n3470) );
  INV_X1 U2537 ( .A(n3471), .ZN(n5808) );
  AOI22_X1 U2538 ( .A1(\mem[102][4] ), .A2(n3467), .B1(n6766), .B2(data_in[4]), 
        .ZN(n3471) );
  INV_X1 U2539 ( .A(n3472), .ZN(n5807) );
  AOI22_X1 U2540 ( .A1(\mem[102][5] ), .A2(n3467), .B1(n6766), .B2(data_in[5]), 
        .ZN(n3472) );
  INV_X1 U2541 ( .A(n3473), .ZN(n5806) );
  AOI22_X1 U2542 ( .A1(\mem[102][6] ), .A2(n3467), .B1(n6766), .B2(data_in[6]), 
        .ZN(n3473) );
  INV_X1 U2543 ( .A(n3474), .ZN(n5805) );
  AOI22_X1 U2544 ( .A1(\mem[102][7] ), .A2(n3467), .B1(n6766), .B2(data_in[7]), 
        .ZN(n3474) );
  INV_X1 U2545 ( .A(n3475), .ZN(n5804) );
  AOI22_X1 U2546 ( .A1(\mem[103][0] ), .A2(n3476), .B1(n6765), .B2(data_in[0]), 
        .ZN(n3475) );
  INV_X1 U2547 ( .A(n3477), .ZN(n5803) );
  AOI22_X1 U2548 ( .A1(\mem[103][1] ), .A2(n3476), .B1(n6765), .B2(data_in[1]), 
        .ZN(n3477) );
  INV_X1 U2549 ( .A(n3478), .ZN(n5802) );
  AOI22_X1 U2550 ( .A1(\mem[103][2] ), .A2(n3476), .B1(n6765), .B2(data_in[2]), 
        .ZN(n3478) );
  INV_X1 U2551 ( .A(n3479), .ZN(n5801) );
  AOI22_X1 U2552 ( .A1(\mem[103][3] ), .A2(n3476), .B1(n6765), .B2(data_in[3]), 
        .ZN(n3479) );
  INV_X1 U2553 ( .A(n3480), .ZN(n5800) );
  AOI22_X1 U2554 ( .A1(\mem[103][4] ), .A2(n3476), .B1(n6765), .B2(data_in[4]), 
        .ZN(n3480) );
  INV_X1 U2555 ( .A(n3481), .ZN(n5799) );
  AOI22_X1 U2556 ( .A1(\mem[103][5] ), .A2(n3476), .B1(n6765), .B2(data_in[5]), 
        .ZN(n3481) );
  INV_X1 U2557 ( .A(n3482), .ZN(n5798) );
  AOI22_X1 U2558 ( .A1(\mem[103][6] ), .A2(n3476), .B1(n6765), .B2(data_in[6]), 
        .ZN(n3482) );
  INV_X1 U2559 ( .A(n3483), .ZN(n5797) );
  AOI22_X1 U2560 ( .A1(\mem[103][7] ), .A2(n3476), .B1(n6765), .B2(data_in[7]), 
        .ZN(n3483) );
  INV_X1 U2561 ( .A(n3484), .ZN(n5796) );
  AOI22_X1 U2562 ( .A1(\mem[104][0] ), .A2(n3485), .B1(n6764), .B2(data_in[0]), 
        .ZN(n3484) );
  INV_X1 U2563 ( .A(n3486), .ZN(n5795) );
  AOI22_X1 U2564 ( .A1(\mem[104][1] ), .A2(n3485), .B1(n6764), .B2(data_in[1]), 
        .ZN(n3486) );
  INV_X1 U2565 ( .A(n3487), .ZN(n5794) );
  AOI22_X1 U2566 ( .A1(\mem[104][2] ), .A2(n3485), .B1(n6764), .B2(data_in[2]), 
        .ZN(n3487) );
  INV_X1 U2567 ( .A(n3488), .ZN(n5793) );
  AOI22_X1 U2568 ( .A1(\mem[104][3] ), .A2(n3485), .B1(n6764), .B2(data_in[3]), 
        .ZN(n3488) );
  INV_X1 U2569 ( .A(n3489), .ZN(n5792) );
  AOI22_X1 U2570 ( .A1(\mem[104][4] ), .A2(n3485), .B1(n6764), .B2(data_in[4]), 
        .ZN(n3489) );
  INV_X1 U2571 ( .A(n3490), .ZN(n5791) );
  AOI22_X1 U2572 ( .A1(\mem[104][5] ), .A2(n3485), .B1(n6764), .B2(data_in[5]), 
        .ZN(n3490) );
  INV_X1 U2573 ( .A(n3491), .ZN(n5790) );
  AOI22_X1 U2574 ( .A1(\mem[104][6] ), .A2(n3485), .B1(n6764), .B2(data_in[6]), 
        .ZN(n3491) );
  INV_X1 U2575 ( .A(n3492), .ZN(n5789) );
  AOI22_X1 U2576 ( .A1(\mem[104][7] ), .A2(n3485), .B1(n6764), .B2(data_in[7]), 
        .ZN(n3492) );
  INV_X1 U2577 ( .A(n3493), .ZN(n5788) );
  AOI22_X1 U2578 ( .A1(\mem[105][0] ), .A2(n3494), .B1(n6763), .B2(data_in[0]), 
        .ZN(n3493) );
  INV_X1 U2579 ( .A(n3495), .ZN(n5787) );
  AOI22_X1 U2580 ( .A1(\mem[105][1] ), .A2(n3494), .B1(n6763), .B2(data_in[1]), 
        .ZN(n3495) );
  INV_X1 U2581 ( .A(n3496), .ZN(n5786) );
  AOI22_X1 U2582 ( .A1(\mem[105][2] ), .A2(n3494), .B1(n6763), .B2(data_in[2]), 
        .ZN(n3496) );
  INV_X1 U2583 ( .A(n3497), .ZN(n5785) );
  AOI22_X1 U2584 ( .A1(\mem[105][3] ), .A2(n3494), .B1(n6763), .B2(data_in[3]), 
        .ZN(n3497) );
  INV_X1 U2585 ( .A(n3498), .ZN(n5784) );
  AOI22_X1 U2586 ( .A1(\mem[105][4] ), .A2(n3494), .B1(n6763), .B2(data_in[4]), 
        .ZN(n3498) );
  INV_X1 U2587 ( .A(n3499), .ZN(n5783) );
  AOI22_X1 U2588 ( .A1(\mem[105][5] ), .A2(n3494), .B1(n6763), .B2(data_in[5]), 
        .ZN(n3499) );
  INV_X1 U2589 ( .A(n3500), .ZN(n5782) );
  AOI22_X1 U2590 ( .A1(\mem[105][6] ), .A2(n3494), .B1(n6763), .B2(data_in[6]), 
        .ZN(n3500) );
  INV_X1 U2591 ( .A(n3501), .ZN(n5781) );
  AOI22_X1 U2592 ( .A1(\mem[105][7] ), .A2(n3494), .B1(n6763), .B2(data_in[7]), 
        .ZN(n3501) );
  INV_X1 U2593 ( .A(n3502), .ZN(n5780) );
  AOI22_X1 U2594 ( .A1(\mem[106][0] ), .A2(n3503), .B1(n6762), .B2(data_in[0]), 
        .ZN(n3502) );
  INV_X1 U2595 ( .A(n3504), .ZN(n5779) );
  AOI22_X1 U2596 ( .A1(\mem[106][1] ), .A2(n3503), .B1(n6762), .B2(data_in[1]), 
        .ZN(n3504) );
  INV_X1 U2597 ( .A(n3505), .ZN(n5778) );
  AOI22_X1 U2598 ( .A1(\mem[106][2] ), .A2(n3503), .B1(n6762), .B2(data_in[2]), 
        .ZN(n3505) );
  INV_X1 U2599 ( .A(n3506), .ZN(n5777) );
  AOI22_X1 U2600 ( .A1(\mem[106][3] ), .A2(n3503), .B1(n6762), .B2(data_in[3]), 
        .ZN(n3506) );
  INV_X1 U2601 ( .A(n3507), .ZN(n5776) );
  AOI22_X1 U2602 ( .A1(\mem[106][4] ), .A2(n3503), .B1(n6762), .B2(data_in[4]), 
        .ZN(n3507) );
  INV_X1 U2603 ( .A(n3508), .ZN(n5775) );
  AOI22_X1 U2604 ( .A1(\mem[106][5] ), .A2(n3503), .B1(n6762), .B2(data_in[5]), 
        .ZN(n3508) );
  INV_X1 U2605 ( .A(n3509), .ZN(n5774) );
  AOI22_X1 U2606 ( .A1(\mem[106][6] ), .A2(n3503), .B1(n6762), .B2(data_in[6]), 
        .ZN(n3509) );
  INV_X1 U2607 ( .A(n3510), .ZN(n5773) );
  AOI22_X1 U2608 ( .A1(\mem[106][7] ), .A2(n3503), .B1(n6762), .B2(data_in[7]), 
        .ZN(n3510) );
  INV_X1 U2609 ( .A(n3511), .ZN(n5772) );
  AOI22_X1 U2610 ( .A1(\mem[107][0] ), .A2(n3512), .B1(n6761), .B2(data_in[0]), 
        .ZN(n3511) );
  INV_X1 U2611 ( .A(n3513), .ZN(n5771) );
  AOI22_X1 U2612 ( .A1(\mem[107][1] ), .A2(n3512), .B1(n6761), .B2(data_in[1]), 
        .ZN(n3513) );
  INV_X1 U2613 ( .A(n3514), .ZN(n5770) );
  AOI22_X1 U2614 ( .A1(\mem[107][2] ), .A2(n3512), .B1(n6761), .B2(data_in[2]), 
        .ZN(n3514) );
  INV_X1 U2615 ( .A(n3515), .ZN(n5769) );
  AOI22_X1 U2616 ( .A1(\mem[107][3] ), .A2(n3512), .B1(n6761), .B2(data_in[3]), 
        .ZN(n3515) );
  INV_X1 U2617 ( .A(n3516), .ZN(n5768) );
  AOI22_X1 U2618 ( .A1(\mem[107][4] ), .A2(n3512), .B1(n6761), .B2(data_in[4]), 
        .ZN(n3516) );
  INV_X1 U2619 ( .A(n3517), .ZN(n5767) );
  AOI22_X1 U2620 ( .A1(\mem[107][5] ), .A2(n3512), .B1(n6761), .B2(data_in[5]), 
        .ZN(n3517) );
  INV_X1 U2621 ( .A(n3518), .ZN(n5766) );
  AOI22_X1 U2622 ( .A1(\mem[107][6] ), .A2(n3512), .B1(n6761), .B2(data_in[6]), 
        .ZN(n3518) );
  INV_X1 U2623 ( .A(n3519), .ZN(n5765) );
  AOI22_X1 U2624 ( .A1(\mem[107][7] ), .A2(n3512), .B1(n6761), .B2(data_in[7]), 
        .ZN(n3519) );
  INV_X1 U2625 ( .A(n3520), .ZN(n5764) );
  AOI22_X1 U2626 ( .A1(\mem[108][0] ), .A2(n3521), .B1(n6760), .B2(data_in[0]), 
        .ZN(n3520) );
  INV_X1 U2627 ( .A(n3522), .ZN(n5763) );
  AOI22_X1 U2628 ( .A1(\mem[108][1] ), .A2(n3521), .B1(n6760), .B2(data_in[1]), 
        .ZN(n3522) );
  INV_X1 U2629 ( .A(n3523), .ZN(n5762) );
  AOI22_X1 U2630 ( .A1(\mem[108][2] ), .A2(n3521), .B1(n6760), .B2(data_in[2]), 
        .ZN(n3523) );
  INV_X1 U2631 ( .A(n3524), .ZN(n5761) );
  AOI22_X1 U2632 ( .A1(\mem[108][3] ), .A2(n3521), .B1(n6760), .B2(data_in[3]), 
        .ZN(n3524) );
  INV_X1 U2633 ( .A(n3525), .ZN(n5760) );
  AOI22_X1 U2634 ( .A1(\mem[108][4] ), .A2(n3521), .B1(n6760), .B2(data_in[4]), 
        .ZN(n3525) );
  INV_X1 U2635 ( .A(n3526), .ZN(n5759) );
  AOI22_X1 U2636 ( .A1(\mem[108][5] ), .A2(n3521), .B1(n6760), .B2(data_in[5]), 
        .ZN(n3526) );
  INV_X1 U2637 ( .A(n3527), .ZN(n5758) );
  AOI22_X1 U2638 ( .A1(\mem[108][6] ), .A2(n3521), .B1(n6760), .B2(data_in[6]), 
        .ZN(n3527) );
  INV_X1 U2639 ( .A(n3528), .ZN(n5757) );
  AOI22_X1 U2640 ( .A1(\mem[108][7] ), .A2(n3521), .B1(n6760), .B2(data_in[7]), 
        .ZN(n3528) );
  INV_X1 U2641 ( .A(n3529), .ZN(n5756) );
  AOI22_X1 U2642 ( .A1(\mem[109][0] ), .A2(n3530), .B1(n6759), .B2(data_in[0]), 
        .ZN(n3529) );
  INV_X1 U2643 ( .A(n3531), .ZN(n5755) );
  AOI22_X1 U2644 ( .A1(\mem[109][1] ), .A2(n3530), .B1(n6759), .B2(data_in[1]), 
        .ZN(n3531) );
  INV_X1 U2645 ( .A(n3532), .ZN(n5754) );
  AOI22_X1 U2646 ( .A1(\mem[109][2] ), .A2(n3530), .B1(n6759), .B2(data_in[2]), 
        .ZN(n3532) );
  INV_X1 U2647 ( .A(n3533), .ZN(n5753) );
  AOI22_X1 U2648 ( .A1(\mem[109][3] ), .A2(n3530), .B1(n6759), .B2(data_in[3]), 
        .ZN(n3533) );
  INV_X1 U2649 ( .A(n3534), .ZN(n5752) );
  AOI22_X1 U2650 ( .A1(\mem[109][4] ), .A2(n3530), .B1(n6759), .B2(data_in[4]), 
        .ZN(n3534) );
  INV_X1 U2651 ( .A(n3535), .ZN(n5751) );
  AOI22_X1 U2652 ( .A1(\mem[109][5] ), .A2(n3530), .B1(n6759), .B2(data_in[5]), 
        .ZN(n3535) );
  INV_X1 U2653 ( .A(n3536), .ZN(n5750) );
  AOI22_X1 U2654 ( .A1(\mem[109][6] ), .A2(n3530), .B1(n6759), .B2(data_in[6]), 
        .ZN(n3536) );
  INV_X1 U2655 ( .A(n3537), .ZN(n5749) );
  AOI22_X1 U2656 ( .A1(\mem[109][7] ), .A2(n3530), .B1(n6759), .B2(data_in[7]), 
        .ZN(n3537) );
  INV_X1 U2657 ( .A(n3538), .ZN(n5748) );
  AOI22_X1 U2658 ( .A1(\mem[110][0] ), .A2(n3539), .B1(n6758), .B2(data_in[0]), 
        .ZN(n3538) );
  INV_X1 U2659 ( .A(n3540), .ZN(n5747) );
  AOI22_X1 U2660 ( .A1(\mem[110][1] ), .A2(n3539), .B1(n6758), .B2(data_in[1]), 
        .ZN(n3540) );
  INV_X1 U2661 ( .A(n3541), .ZN(n5746) );
  AOI22_X1 U2662 ( .A1(\mem[110][2] ), .A2(n3539), .B1(n6758), .B2(data_in[2]), 
        .ZN(n3541) );
  INV_X1 U2663 ( .A(n3542), .ZN(n5745) );
  AOI22_X1 U2664 ( .A1(\mem[110][3] ), .A2(n3539), .B1(n6758), .B2(data_in[3]), 
        .ZN(n3542) );
  INV_X1 U2665 ( .A(n3543), .ZN(n5744) );
  AOI22_X1 U2666 ( .A1(\mem[110][4] ), .A2(n3539), .B1(n6758), .B2(data_in[4]), 
        .ZN(n3543) );
  INV_X1 U2667 ( .A(n3544), .ZN(n5743) );
  AOI22_X1 U2668 ( .A1(\mem[110][5] ), .A2(n3539), .B1(n6758), .B2(data_in[5]), 
        .ZN(n3544) );
  INV_X1 U2669 ( .A(n3545), .ZN(n5742) );
  AOI22_X1 U2670 ( .A1(\mem[110][6] ), .A2(n3539), .B1(n6758), .B2(data_in[6]), 
        .ZN(n3545) );
  INV_X1 U2671 ( .A(n3546), .ZN(n5741) );
  AOI22_X1 U2672 ( .A1(\mem[110][7] ), .A2(n3539), .B1(n6758), .B2(data_in[7]), 
        .ZN(n3546) );
  INV_X1 U2673 ( .A(n3547), .ZN(n5740) );
  AOI22_X1 U2674 ( .A1(\mem[111][0] ), .A2(n3548), .B1(n6757), .B2(data_in[0]), 
        .ZN(n3547) );
  INV_X1 U2675 ( .A(n3549), .ZN(n5739) );
  AOI22_X1 U2676 ( .A1(\mem[111][1] ), .A2(n3548), .B1(n6757), .B2(data_in[1]), 
        .ZN(n3549) );
  INV_X1 U2677 ( .A(n3550), .ZN(n5738) );
  AOI22_X1 U2678 ( .A1(\mem[111][2] ), .A2(n3548), .B1(n6757), .B2(data_in[2]), 
        .ZN(n3550) );
  INV_X1 U2679 ( .A(n3551), .ZN(n5737) );
  AOI22_X1 U2680 ( .A1(\mem[111][3] ), .A2(n3548), .B1(n6757), .B2(data_in[3]), 
        .ZN(n3551) );
  INV_X1 U2681 ( .A(n3552), .ZN(n5736) );
  AOI22_X1 U2682 ( .A1(\mem[111][4] ), .A2(n3548), .B1(n6757), .B2(data_in[4]), 
        .ZN(n3552) );
  INV_X1 U2683 ( .A(n3553), .ZN(n5735) );
  AOI22_X1 U2684 ( .A1(\mem[111][5] ), .A2(n3548), .B1(n6757), .B2(data_in[5]), 
        .ZN(n3553) );
  INV_X1 U2685 ( .A(n3554), .ZN(n5734) );
  AOI22_X1 U2686 ( .A1(\mem[111][6] ), .A2(n3548), .B1(n6757), .B2(data_in[6]), 
        .ZN(n3554) );
  INV_X1 U2687 ( .A(n3555), .ZN(n5733) );
  AOI22_X1 U2688 ( .A1(\mem[111][7] ), .A2(n3548), .B1(n6757), .B2(data_in[7]), 
        .ZN(n3555) );
  INV_X1 U2689 ( .A(n3556), .ZN(n5732) );
  AOI22_X1 U2690 ( .A1(\mem[112][0] ), .A2(n3557), .B1(n6756), .B2(data_in[0]), 
        .ZN(n3556) );
  INV_X1 U2691 ( .A(n3558), .ZN(n5731) );
  AOI22_X1 U2692 ( .A1(\mem[112][1] ), .A2(n3557), .B1(n6756), .B2(data_in[1]), 
        .ZN(n3558) );
  INV_X1 U2693 ( .A(n3559), .ZN(n5730) );
  AOI22_X1 U2694 ( .A1(\mem[112][2] ), .A2(n3557), .B1(n6756), .B2(data_in[2]), 
        .ZN(n3559) );
  INV_X1 U2695 ( .A(n3560), .ZN(n5729) );
  AOI22_X1 U2696 ( .A1(\mem[112][3] ), .A2(n3557), .B1(n6756), .B2(data_in[3]), 
        .ZN(n3560) );
  INV_X1 U2697 ( .A(n3561), .ZN(n5728) );
  AOI22_X1 U2698 ( .A1(\mem[112][4] ), .A2(n3557), .B1(n6756), .B2(data_in[4]), 
        .ZN(n3561) );
  INV_X1 U2699 ( .A(n3562), .ZN(n5727) );
  AOI22_X1 U2700 ( .A1(\mem[112][5] ), .A2(n3557), .B1(n6756), .B2(data_in[5]), 
        .ZN(n3562) );
  INV_X1 U2701 ( .A(n3563), .ZN(n5726) );
  AOI22_X1 U2702 ( .A1(\mem[112][6] ), .A2(n3557), .B1(n6756), .B2(data_in[6]), 
        .ZN(n3563) );
  INV_X1 U2703 ( .A(n3564), .ZN(n5725) );
  AOI22_X1 U2704 ( .A1(\mem[112][7] ), .A2(n3557), .B1(n6756), .B2(data_in[7]), 
        .ZN(n3564) );
  INV_X1 U2705 ( .A(n3566), .ZN(n5724) );
  AOI22_X1 U2706 ( .A1(\mem[113][0] ), .A2(n3567), .B1(n6755), .B2(data_in[0]), 
        .ZN(n3566) );
  INV_X1 U2707 ( .A(n3568), .ZN(n5723) );
  AOI22_X1 U2708 ( .A1(\mem[113][1] ), .A2(n3567), .B1(n6755), .B2(data_in[1]), 
        .ZN(n3568) );
  INV_X1 U2709 ( .A(n3569), .ZN(n5722) );
  AOI22_X1 U2710 ( .A1(\mem[113][2] ), .A2(n3567), .B1(n6755), .B2(data_in[2]), 
        .ZN(n3569) );
  INV_X1 U2711 ( .A(n3570), .ZN(n5721) );
  AOI22_X1 U2712 ( .A1(\mem[113][3] ), .A2(n3567), .B1(n6755), .B2(data_in[3]), 
        .ZN(n3570) );
  INV_X1 U2713 ( .A(n3571), .ZN(n5720) );
  AOI22_X1 U2714 ( .A1(\mem[113][4] ), .A2(n3567), .B1(n6755), .B2(data_in[4]), 
        .ZN(n3571) );
  INV_X1 U2715 ( .A(n3572), .ZN(n5719) );
  AOI22_X1 U2716 ( .A1(\mem[113][5] ), .A2(n3567), .B1(n6755), .B2(data_in[5]), 
        .ZN(n3572) );
  INV_X1 U2717 ( .A(n3573), .ZN(n5718) );
  AOI22_X1 U2718 ( .A1(\mem[113][6] ), .A2(n3567), .B1(n6755), .B2(data_in[6]), 
        .ZN(n3573) );
  INV_X1 U2719 ( .A(n3574), .ZN(n5717) );
  AOI22_X1 U2720 ( .A1(\mem[113][7] ), .A2(n3567), .B1(n6755), .B2(data_in[7]), 
        .ZN(n3574) );
  INV_X1 U2721 ( .A(n3575), .ZN(n5716) );
  AOI22_X1 U2722 ( .A1(\mem[114][0] ), .A2(n3576), .B1(n6754), .B2(data_in[0]), 
        .ZN(n3575) );
  INV_X1 U2723 ( .A(n3577), .ZN(n5715) );
  AOI22_X1 U2724 ( .A1(\mem[114][1] ), .A2(n3576), .B1(n6754), .B2(data_in[1]), 
        .ZN(n3577) );
  INV_X1 U2725 ( .A(n3578), .ZN(n5714) );
  AOI22_X1 U2726 ( .A1(\mem[114][2] ), .A2(n3576), .B1(n6754), .B2(data_in[2]), 
        .ZN(n3578) );
  INV_X1 U2727 ( .A(n3579), .ZN(n5713) );
  AOI22_X1 U2728 ( .A1(\mem[114][3] ), .A2(n3576), .B1(n6754), .B2(data_in[3]), 
        .ZN(n3579) );
  INV_X1 U2729 ( .A(n3580), .ZN(n5712) );
  AOI22_X1 U2730 ( .A1(\mem[114][4] ), .A2(n3576), .B1(n6754), .B2(data_in[4]), 
        .ZN(n3580) );
  INV_X1 U2731 ( .A(n3581), .ZN(n5711) );
  AOI22_X1 U2732 ( .A1(\mem[114][5] ), .A2(n3576), .B1(n6754), .B2(data_in[5]), 
        .ZN(n3581) );
  INV_X1 U2733 ( .A(n3582), .ZN(n5710) );
  AOI22_X1 U2734 ( .A1(\mem[114][6] ), .A2(n3576), .B1(n6754), .B2(data_in[6]), 
        .ZN(n3582) );
  INV_X1 U2735 ( .A(n3583), .ZN(n5709) );
  AOI22_X1 U2736 ( .A1(\mem[114][7] ), .A2(n3576), .B1(n6754), .B2(data_in[7]), 
        .ZN(n3583) );
  INV_X1 U2737 ( .A(n3584), .ZN(n5708) );
  AOI22_X1 U2738 ( .A1(\mem[115][0] ), .A2(n3585), .B1(n6753), .B2(data_in[0]), 
        .ZN(n3584) );
  INV_X1 U2739 ( .A(n3586), .ZN(n5707) );
  AOI22_X1 U2740 ( .A1(\mem[115][1] ), .A2(n3585), .B1(n6753), .B2(data_in[1]), 
        .ZN(n3586) );
  INV_X1 U2741 ( .A(n3587), .ZN(n5706) );
  AOI22_X1 U2742 ( .A1(\mem[115][2] ), .A2(n3585), .B1(n6753), .B2(data_in[2]), 
        .ZN(n3587) );
  INV_X1 U2743 ( .A(n3588), .ZN(n5705) );
  AOI22_X1 U2744 ( .A1(\mem[115][3] ), .A2(n3585), .B1(n6753), .B2(data_in[3]), 
        .ZN(n3588) );
  INV_X1 U2745 ( .A(n3589), .ZN(n5704) );
  AOI22_X1 U2746 ( .A1(\mem[115][4] ), .A2(n3585), .B1(n6753), .B2(data_in[4]), 
        .ZN(n3589) );
  INV_X1 U2747 ( .A(n3590), .ZN(n5703) );
  AOI22_X1 U2748 ( .A1(\mem[115][5] ), .A2(n3585), .B1(n6753), .B2(data_in[5]), 
        .ZN(n3590) );
  INV_X1 U2749 ( .A(n3591), .ZN(n5702) );
  AOI22_X1 U2750 ( .A1(\mem[115][6] ), .A2(n3585), .B1(n6753), .B2(data_in[6]), 
        .ZN(n3591) );
  INV_X1 U2751 ( .A(n3592), .ZN(n5701) );
  AOI22_X1 U2752 ( .A1(\mem[115][7] ), .A2(n3585), .B1(n6753), .B2(data_in[7]), 
        .ZN(n3592) );
  INV_X1 U2753 ( .A(n3593), .ZN(n5700) );
  AOI22_X1 U2754 ( .A1(\mem[116][0] ), .A2(n3594), .B1(n6752), .B2(data_in[0]), 
        .ZN(n3593) );
  INV_X1 U2755 ( .A(n3595), .ZN(n5699) );
  AOI22_X1 U2756 ( .A1(\mem[116][1] ), .A2(n3594), .B1(n6752), .B2(data_in[1]), 
        .ZN(n3595) );
  INV_X1 U2757 ( .A(n3596), .ZN(n5698) );
  AOI22_X1 U2758 ( .A1(\mem[116][2] ), .A2(n3594), .B1(n6752), .B2(data_in[2]), 
        .ZN(n3596) );
  INV_X1 U2759 ( .A(n3597), .ZN(n5697) );
  AOI22_X1 U2760 ( .A1(\mem[116][3] ), .A2(n3594), .B1(n6752), .B2(data_in[3]), 
        .ZN(n3597) );
  INV_X1 U2761 ( .A(n3598), .ZN(n5696) );
  AOI22_X1 U2762 ( .A1(\mem[116][4] ), .A2(n3594), .B1(n6752), .B2(data_in[4]), 
        .ZN(n3598) );
  INV_X1 U2763 ( .A(n3599), .ZN(n5695) );
  AOI22_X1 U2764 ( .A1(\mem[116][5] ), .A2(n3594), .B1(n6752), .B2(data_in[5]), 
        .ZN(n3599) );
  INV_X1 U2765 ( .A(n3600), .ZN(n5694) );
  AOI22_X1 U2766 ( .A1(\mem[116][6] ), .A2(n3594), .B1(n6752), .B2(data_in[6]), 
        .ZN(n3600) );
  INV_X1 U2767 ( .A(n3601), .ZN(n5693) );
  AOI22_X1 U2768 ( .A1(\mem[116][7] ), .A2(n3594), .B1(n6752), .B2(data_in[7]), 
        .ZN(n3601) );
  INV_X1 U2769 ( .A(n3602), .ZN(n5692) );
  AOI22_X1 U2770 ( .A1(\mem[117][0] ), .A2(n3603), .B1(n6751), .B2(data_in[0]), 
        .ZN(n3602) );
  INV_X1 U2771 ( .A(n3604), .ZN(n5691) );
  AOI22_X1 U2772 ( .A1(\mem[117][1] ), .A2(n3603), .B1(n6751), .B2(data_in[1]), 
        .ZN(n3604) );
  INV_X1 U2773 ( .A(n3605), .ZN(n5690) );
  AOI22_X1 U2774 ( .A1(\mem[117][2] ), .A2(n3603), .B1(n6751), .B2(data_in[2]), 
        .ZN(n3605) );
  INV_X1 U2775 ( .A(n3606), .ZN(n5689) );
  AOI22_X1 U2776 ( .A1(\mem[117][3] ), .A2(n3603), .B1(n6751), .B2(data_in[3]), 
        .ZN(n3606) );
  INV_X1 U2777 ( .A(n3607), .ZN(n5688) );
  AOI22_X1 U2778 ( .A1(\mem[117][4] ), .A2(n3603), .B1(n6751), .B2(data_in[4]), 
        .ZN(n3607) );
  INV_X1 U2779 ( .A(n3608), .ZN(n5687) );
  AOI22_X1 U2780 ( .A1(\mem[117][5] ), .A2(n3603), .B1(n6751), .B2(data_in[5]), 
        .ZN(n3608) );
  INV_X1 U2781 ( .A(n3609), .ZN(n5686) );
  AOI22_X1 U2782 ( .A1(\mem[117][6] ), .A2(n3603), .B1(n6751), .B2(data_in[6]), 
        .ZN(n3609) );
  INV_X1 U2783 ( .A(n3610), .ZN(n5685) );
  AOI22_X1 U2784 ( .A1(\mem[117][7] ), .A2(n3603), .B1(n6751), .B2(data_in[7]), 
        .ZN(n3610) );
  INV_X1 U2785 ( .A(n3611), .ZN(n5684) );
  AOI22_X1 U2786 ( .A1(\mem[118][0] ), .A2(n3612), .B1(n6750), .B2(data_in[0]), 
        .ZN(n3611) );
  INV_X1 U2787 ( .A(n3613), .ZN(n5683) );
  AOI22_X1 U2788 ( .A1(\mem[118][1] ), .A2(n3612), .B1(n6750), .B2(data_in[1]), 
        .ZN(n3613) );
  INV_X1 U2789 ( .A(n3614), .ZN(n5682) );
  AOI22_X1 U2790 ( .A1(\mem[118][2] ), .A2(n3612), .B1(n6750), .B2(data_in[2]), 
        .ZN(n3614) );
  INV_X1 U2791 ( .A(n3615), .ZN(n5681) );
  AOI22_X1 U2792 ( .A1(\mem[118][3] ), .A2(n3612), .B1(n6750), .B2(data_in[3]), 
        .ZN(n3615) );
  INV_X1 U2793 ( .A(n3616), .ZN(n5680) );
  AOI22_X1 U2794 ( .A1(\mem[118][4] ), .A2(n3612), .B1(n6750), .B2(data_in[4]), 
        .ZN(n3616) );
  INV_X1 U2795 ( .A(n3617), .ZN(n5679) );
  AOI22_X1 U2796 ( .A1(\mem[118][5] ), .A2(n3612), .B1(n6750), .B2(data_in[5]), 
        .ZN(n3617) );
  INV_X1 U2797 ( .A(n3618), .ZN(n5678) );
  AOI22_X1 U2798 ( .A1(\mem[118][6] ), .A2(n3612), .B1(n6750), .B2(data_in[6]), 
        .ZN(n3618) );
  INV_X1 U2799 ( .A(n3619), .ZN(n5677) );
  AOI22_X1 U2800 ( .A1(\mem[118][7] ), .A2(n3612), .B1(n6750), .B2(data_in[7]), 
        .ZN(n3619) );
  INV_X1 U2801 ( .A(n3620), .ZN(n5676) );
  AOI22_X1 U2802 ( .A1(\mem[119][0] ), .A2(n3621), .B1(n6749), .B2(data_in[0]), 
        .ZN(n3620) );
  INV_X1 U2803 ( .A(n3622), .ZN(n5675) );
  AOI22_X1 U2804 ( .A1(\mem[119][1] ), .A2(n3621), .B1(n6749), .B2(data_in[1]), 
        .ZN(n3622) );
  INV_X1 U2805 ( .A(n3623), .ZN(n5674) );
  AOI22_X1 U2806 ( .A1(\mem[119][2] ), .A2(n3621), .B1(n6749), .B2(data_in[2]), 
        .ZN(n3623) );
  INV_X1 U2807 ( .A(n3624), .ZN(n5673) );
  AOI22_X1 U2808 ( .A1(\mem[119][3] ), .A2(n3621), .B1(n6749), .B2(data_in[3]), 
        .ZN(n3624) );
  INV_X1 U2809 ( .A(n3625), .ZN(n5672) );
  AOI22_X1 U2810 ( .A1(\mem[119][4] ), .A2(n3621), .B1(n6749), .B2(data_in[4]), 
        .ZN(n3625) );
  INV_X1 U2811 ( .A(n3626), .ZN(n5671) );
  AOI22_X1 U2812 ( .A1(\mem[119][5] ), .A2(n3621), .B1(n6749), .B2(data_in[5]), 
        .ZN(n3626) );
  INV_X1 U2813 ( .A(n3627), .ZN(n5670) );
  AOI22_X1 U2814 ( .A1(\mem[119][6] ), .A2(n3621), .B1(n6749), .B2(data_in[6]), 
        .ZN(n3627) );
  INV_X1 U2815 ( .A(n3628), .ZN(n5669) );
  AOI22_X1 U2816 ( .A1(\mem[119][7] ), .A2(n3621), .B1(n6749), .B2(data_in[7]), 
        .ZN(n3628) );
  INV_X1 U2817 ( .A(n3629), .ZN(n5668) );
  AOI22_X1 U2818 ( .A1(\mem[120][0] ), .A2(n3630), .B1(n6748), .B2(data_in[0]), 
        .ZN(n3629) );
  INV_X1 U2819 ( .A(n3631), .ZN(n5667) );
  AOI22_X1 U2820 ( .A1(\mem[120][1] ), .A2(n3630), .B1(n6748), .B2(data_in[1]), 
        .ZN(n3631) );
  INV_X1 U2821 ( .A(n3632), .ZN(n5666) );
  AOI22_X1 U2822 ( .A1(\mem[120][2] ), .A2(n3630), .B1(n6748), .B2(data_in[2]), 
        .ZN(n3632) );
  INV_X1 U2823 ( .A(n3633), .ZN(n5665) );
  AOI22_X1 U2824 ( .A1(\mem[120][3] ), .A2(n3630), .B1(n6748), .B2(data_in[3]), 
        .ZN(n3633) );
  INV_X1 U2825 ( .A(n3634), .ZN(n5664) );
  AOI22_X1 U2826 ( .A1(\mem[120][4] ), .A2(n3630), .B1(n6748), .B2(data_in[4]), 
        .ZN(n3634) );
  INV_X1 U2827 ( .A(n3635), .ZN(n5663) );
  AOI22_X1 U2828 ( .A1(\mem[120][5] ), .A2(n3630), .B1(n6748), .B2(data_in[5]), 
        .ZN(n3635) );
  INV_X1 U2829 ( .A(n3636), .ZN(n5662) );
  AOI22_X1 U2830 ( .A1(\mem[120][6] ), .A2(n3630), .B1(n6748), .B2(data_in[6]), 
        .ZN(n3636) );
  INV_X1 U2831 ( .A(n3637), .ZN(n5661) );
  AOI22_X1 U2832 ( .A1(\mem[120][7] ), .A2(n3630), .B1(n6748), .B2(data_in[7]), 
        .ZN(n3637) );
  INV_X1 U2833 ( .A(n3638), .ZN(n5660) );
  AOI22_X1 U2834 ( .A1(\mem[121][0] ), .A2(n3639), .B1(n6747), .B2(data_in[0]), 
        .ZN(n3638) );
  INV_X1 U2835 ( .A(n3640), .ZN(n5659) );
  AOI22_X1 U2836 ( .A1(\mem[121][1] ), .A2(n3639), .B1(n6747), .B2(data_in[1]), 
        .ZN(n3640) );
  INV_X1 U2837 ( .A(n3641), .ZN(n5658) );
  AOI22_X1 U2838 ( .A1(\mem[121][2] ), .A2(n3639), .B1(n6747), .B2(data_in[2]), 
        .ZN(n3641) );
  INV_X1 U2839 ( .A(n3642), .ZN(n5657) );
  AOI22_X1 U2840 ( .A1(\mem[121][3] ), .A2(n3639), .B1(n6747), .B2(data_in[3]), 
        .ZN(n3642) );
  INV_X1 U2841 ( .A(n3643), .ZN(n5656) );
  AOI22_X1 U2842 ( .A1(\mem[121][4] ), .A2(n3639), .B1(n6747), .B2(data_in[4]), 
        .ZN(n3643) );
  INV_X1 U2843 ( .A(n3644), .ZN(n5655) );
  AOI22_X1 U2844 ( .A1(\mem[121][5] ), .A2(n3639), .B1(n6747), .B2(data_in[5]), 
        .ZN(n3644) );
  INV_X1 U2845 ( .A(n3645), .ZN(n5654) );
  AOI22_X1 U2846 ( .A1(\mem[121][6] ), .A2(n3639), .B1(n6747), .B2(data_in[6]), 
        .ZN(n3645) );
  INV_X1 U2847 ( .A(n3646), .ZN(n5653) );
  AOI22_X1 U2848 ( .A1(\mem[121][7] ), .A2(n3639), .B1(n6747), .B2(data_in[7]), 
        .ZN(n3646) );
  INV_X1 U2849 ( .A(n3647), .ZN(n5652) );
  AOI22_X1 U2850 ( .A1(\mem[122][0] ), .A2(n3648), .B1(n6746), .B2(data_in[0]), 
        .ZN(n3647) );
  INV_X1 U2851 ( .A(n3649), .ZN(n5651) );
  AOI22_X1 U2852 ( .A1(\mem[122][1] ), .A2(n3648), .B1(n6746), .B2(data_in[1]), 
        .ZN(n3649) );
  INV_X1 U2853 ( .A(n3650), .ZN(n5650) );
  AOI22_X1 U2854 ( .A1(\mem[122][2] ), .A2(n3648), .B1(n6746), .B2(data_in[2]), 
        .ZN(n3650) );
  INV_X1 U2855 ( .A(n3651), .ZN(n5649) );
  AOI22_X1 U2856 ( .A1(\mem[122][3] ), .A2(n3648), .B1(n6746), .B2(data_in[3]), 
        .ZN(n3651) );
  INV_X1 U2857 ( .A(n3652), .ZN(n5648) );
  AOI22_X1 U2858 ( .A1(\mem[122][4] ), .A2(n3648), .B1(n6746), .B2(data_in[4]), 
        .ZN(n3652) );
  INV_X1 U2859 ( .A(n3653), .ZN(n5647) );
  AOI22_X1 U2860 ( .A1(\mem[122][5] ), .A2(n3648), .B1(n6746), .B2(data_in[5]), 
        .ZN(n3653) );
  INV_X1 U2861 ( .A(n3654), .ZN(n5646) );
  AOI22_X1 U2862 ( .A1(\mem[122][6] ), .A2(n3648), .B1(n6746), .B2(data_in[6]), 
        .ZN(n3654) );
  INV_X1 U2863 ( .A(n3655), .ZN(n5645) );
  AOI22_X1 U2864 ( .A1(\mem[122][7] ), .A2(n3648), .B1(n6746), .B2(data_in[7]), 
        .ZN(n3655) );
  INV_X1 U2865 ( .A(n3656), .ZN(n5644) );
  AOI22_X1 U2866 ( .A1(\mem[123][0] ), .A2(n3657), .B1(n6745), .B2(data_in[0]), 
        .ZN(n3656) );
  INV_X1 U2867 ( .A(n3658), .ZN(n5643) );
  AOI22_X1 U2868 ( .A1(\mem[123][1] ), .A2(n3657), .B1(n6745), .B2(data_in[1]), 
        .ZN(n3658) );
  INV_X1 U2869 ( .A(n3659), .ZN(n5642) );
  AOI22_X1 U2870 ( .A1(\mem[123][2] ), .A2(n3657), .B1(n6745), .B2(data_in[2]), 
        .ZN(n3659) );
  INV_X1 U2871 ( .A(n3660), .ZN(n5641) );
  AOI22_X1 U2872 ( .A1(\mem[123][3] ), .A2(n3657), .B1(n6745), .B2(data_in[3]), 
        .ZN(n3660) );
  INV_X1 U2873 ( .A(n3661), .ZN(n5640) );
  AOI22_X1 U2874 ( .A1(\mem[123][4] ), .A2(n3657), .B1(n6745), .B2(data_in[4]), 
        .ZN(n3661) );
  INV_X1 U2875 ( .A(n3662), .ZN(n5639) );
  AOI22_X1 U2876 ( .A1(\mem[123][5] ), .A2(n3657), .B1(n6745), .B2(data_in[5]), 
        .ZN(n3662) );
  INV_X1 U2877 ( .A(n3663), .ZN(n5638) );
  AOI22_X1 U2878 ( .A1(\mem[123][6] ), .A2(n3657), .B1(n6745), .B2(data_in[6]), 
        .ZN(n3663) );
  INV_X1 U2879 ( .A(n3664), .ZN(n5637) );
  AOI22_X1 U2880 ( .A1(\mem[123][7] ), .A2(n3657), .B1(n6745), .B2(data_in[7]), 
        .ZN(n3664) );
  INV_X1 U2881 ( .A(n3665), .ZN(n5636) );
  AOI22_X1 U2882 ( .A1(\mem[124][0] ), .A2(n3666), .B1(n6744), .B2(data_in[0]), 
        .ZN(n3665) );
  INV_X1 U2883 ( .A(n3667), .ZN(n5635) );
  AOI22_X1 U2884 ( .A1(\mem[124][1] ), .A2(n3666), .B1(n6744), .B2(data_in[1]), 
        .ZN(n3667) );
  INV_X1 U2885 ( .A(n3668), .ZN(n5634) );
  AOI22_X1 U2886 ( .A1(\mem[124][2] ), .A2(n3666), .B1(n6744), .B2(data_in[2]), 
        .ZN(n3668) );
  INV_X1 U2887 ( .A(n3669), .ZN(n5633) );
  AOI22_X1 U2888 ( .A1(\mem[124][3] ), .A2(n3666), .B1(n6744), .B2(data_in[3]), 
        .ZN(n3669) );
  INV_X1 U2889 ( .A(n3670), .ZN(n5632) );
  AOI22_X1 U2890 ( .A1(\mem[124][4] ), .A2(n3666), .B1(n6744), .B2(data_in[4]), 
        .ZN(n3670) );
  INV_X1 U2891 ( .A(n3671), .ZN(n5631) );
  AOI22_X1 U2892 ( .A1(\mem[124][5] ), .A2(n3666), .B1(n6744), .B2(data_in[5]), 
        .ZN(n3671) );
  INV_X1 U2893 ( .A(n3672), .ZN(n5630) );
  AOI22_X1 U2894 ( .A1(\mem[124][6] ), .A2(n3666), .B1(n6744), .B2(data_in[6]), 
        .ZN(n3672) );
  INV_X1 U2895 ( .A(n3673), .ZN(n5629) );
  AOI22_X1 U2896 ( .A1(\mem[124][7] ), .A2(n3666), .B1(n6744), .B2(data_in[7]), 
        .ZN(n3673) );
  INV_X1 U2897 ( .A(n3674), .ZN(n5628) );
  AOI22_X1 U2898 ( .A1(\mem[125][0] ), .A2(n3675), .B1(n6743), .B2(data_in[0]), 
        .ZN(n3674) );
  INV_X1 U2899 ( .A(n3676), .ZN(n5627) );
  AOI22_X1 U2900 ( .A1(\mem[125][1] ), .A2(n3675), .B1(n6743), .B2(data_in[1]), 
        .ZN(n3676) );
  INV_X1 U2901 ( .A(n3677), .ZN(n5626) );
  AOI22_X1 U2902 ( .A1(\mem[125][2] ), .A2(n3675), .B1(n6743), .B2(data_in[2]), 
        .ZN(n3677) );
  INV_X1 U2903 ( .A(n3678), .ZN(n5625) );
  AOI22_X1 U2904 ( .A1(\mem[125][3] ), .A2(n3675), .B1(n6743), .B2(data_in[3]), 
        .ZN(n3678) );
  INV_X1 U2905 ( .A(n3679), .ZN(n5624) );
  AOI22_X1 U2906 ( .A1(\mem[125][4] ), .A2(n3675), .B1(n6743), .B2(data_in[4]), 
        .ZN(n3679) );
  INV_X1 U2907 ( .A(n3680), .ZN(n5623) );
  AOI22_X1 U2908 ( .A1(\mem[125][5] ), .A2(n3675), .B1(n6743), .B2(data_in[5]), 
        .ZN(n3680) );
  INV_X1 U2909 ( .A(n3681), .ZN(n5622) );
  AOI22_X1 U2910 ( .A1(\mem[125][6] ), .A2(n3675), .B1(n6743), .B2(data_in[6]), 
        .ZN(n3681) );
  INV_X1 U2911 ( .A(n3682), .ZN(n5621) );
  AOI22_X1 U2912 ( .A1(\mem[125][7] ), .A2(n3675), .B1(n6743), .B2(data_in[7]), 
        .ZN(n3682) );
  INV_X1 U2913 ( .A(n3683), .ZN(n5620) );
  AOI22_X1 U2914 ( .A1(\mem[126][0] ), .A2(n3684), .B1(n6742), .B2(data_in[0]), 
        .ZN(n3683) );
  INV_X1 U2915 ( .A(n3685), .ZN(n5619) );
  AOI22_X1 U2916 ( .A1(\mem[126][1] ), .A2(n3684), .B1(n6742), .B2(data_in[1]), 
        .ZN(n3685) );
  INV_X1 U2917 ( .A(n3686), .ZN(n5618) );
  AOI22_X1 U2918 ( .A1(\mem[126][2] ), .A2(n3684), .B1(n6742), .B2(data_in[2]), 
        .ZN(n3686) );
  INV_X1 U2919 ( .A(n3687), .ZN(n5617) );
  AOI22_X1 U2920 ( .A1(\mem[126][3] ), .A2(n3684), .B1(n6742), .B2(data_in[3]), 
        .ZN(n3687) );
  INV_X1 U2921 ( .A(n3688), .ZN(n5616) );
  AOI22_X1 U2922 ( .A1(\mem[126][4] ), .A2(n3684), .B1(n6742), .B2(data_in[4]), 
        .ZN(n3688) );
  INV_X1 U2923 ( .A(n3689), .ZN(n5615) );
  AOI22_X1 U2924 ( .A1(\mem[126][5] ), .A2(n3684), .B1(n6742), .B2(data_in[5]), 
        .ZN(n3689) );
  INV_X1 U2925 ( .A(n3690), .ZN(n5614) );
  AOI22_X1 U2926 ( .A1(\mem[126][6] ), .A2(n3684), .B1(n6742), .B2(data_in[6]), 
        .ZN(n3690) );
  INV_X1 U2927 ( .A(n3691), .ZN(n5613) );
  AOI22_X1 U2928 ( .A1(\mem[126][7] ), .A2(n3684), .B1(n6742), .B2(data_in[7]), 
        .ZN(n3691) );
  INV_X1 U2929 ( .A(n3692), .ZN(n5612) );
  AOI22_X1 U2930 ( .A1(\mem[127][0] ), .A2(n3693), .B1(n6741), .B2(data_in[0]), 
        .ZN(n3692) );
  INV_X1 U2931 ( .A(n3694), .ZN(n5611) );
  AOI22_X1 U2932 ( .A1(\mem[127][1] ), .A2(n3693), .B1(n6741), .B2(data_in[1]), 
        .ZN(n3694) );
  INV_X1 U2933 ( .A(n3695), .ZN(n5610) );
  AOI22_X1 U2934 ( .A1(\mem[127][2] ), .A2(n3693), .B1(n6741), .B2(data_in[2]), 
        .ZN(n3695) );
  INV_X1 U2935 ( .A(n3696), .ZN(n5609) );
  AOI22_X1 U2936 ( .A1(\mem[127][3] ), .A2(n3693), .B1(n6741), .B2(data_in[3]), 
        .ZN(n3696) );
  INV_X1 U2937 ( .A(n3697), .ZN(n5608) );
  AOI22_X1 U2938 ( .A1(\mem[127][4] ), .A2(n3693), .B1(n6741), .B2(data_in[4]), 
        .ZN(n3697) );
  INV_X1 U2939 ( .A(n3698), .ZN(n5607) );
  AOI22_X1 U2940 ( .A1(\mem[127][5] ), .A2(n3693), .B1(n6741), .B2(data_in[5]), 
        .ZN(n3698) );
  INV_X1 U2941 ( .A(n3699), .ZN(n5606) );
  AOI22_X1 U2942 ( .A1(\mem[127][6] ), .A2(n3693), .B1(n6741), .B2(data_in[6]), 
        .ZN(n3699) );
  INV_X1 U2943 ( .A(n3700), .ZN(n5605) );
  AOI22_X1 U2944 ( .A1(\mem[127][7] ), .A2(n3693), .B1(n6741), .B2(data_in[7]), 
        .ZN(n3700) );
  INV_X1 U2945 ( .A(n3701), .ZN(n5604) );
  AOI22_X1 U2946 ( .A1(\mem[128][0] ), .A2(n3702), .B1(n6740), .B2(data_in[0]), 
        .ZN(n3701) );
  INV_X1 U2947 ( .A(n3703), .ZN(n5603) );
  AOI22_X1 U2948 ( .A1(\mem[128][1] ), .A2(n3702), .B1(n6740), .B2(data_in[1]), 
        .ZN(n3703) );
  INV_X1 U2949 ( .A(n3704), .ZN(n5602) );
  AOI22_X1 U2950 ( .A1(\mem[128][2] ), .A2(n3702), .B1(n6740), .B2(data_in[2]), 
        .ZN(n3704) );
  INV_X1 U2951 ( .A(n3705), .ZN(n5601) );
  AOI22_X1 U2952 ( .A1(\mem[128][3] ), .A2(n3702), .B1(n6740), .B2(data_in[3]), 
        .ZN(n3705) );
  INV_X1 U2953 ( .A(n3706), .ZN(n5600) );
  AOI22_X1 U2954 ( .A1(\mem[128][4] ), .A2(n3702), .B1(n6740), .B2(data_in[4]), 
        .ZN(n3706) );
  INV_X1 U2955 ( .A(n3707), .ZN(n5599) );
  AOI22_X1 U2956 ( .A1(\mem[128][5] ), .A2(n3702), .B1(n6740), .B2(data_in[5]), 
        .ZN(n3707) );
  INV_X1 U2957 ( .A(n3708), .ZN(n5598) );
  AOI22_X1 U2958 ( .A1(\mem[128][6] ), .A2(n3702), .B1(n6740), .B2(data_in[6]), 
        .ZN(n3708) );
  INV_X1 U2959 ( .A(n3709), .ZN(n5597) );
  AOI22_X1 U2960 ( .A1(\mem[128][7] ), .A2(n3702), .B1(n6740), .B2(data_in[7]), 
        .ZN(n3709) );
  INV_X1 U2961 ( .A(n3711), .ZN(n5596) );
  AOI22_X1 U2962 ( .A1(\mem[129][0] ), .A2(n3712), .B1(n6739), .B2(data_in[0]), 
        .ZN(n3711) );
  INV_X1 U2963 ( .A(n3713), .ZN(n5595) );
  AOI22_X1 U2964 ( .A1(\mem[129][1] ), .A2(n3712), .B1(n6739), .B2(data_in[1]), 
        .ZN(n3713) );
  INV_X1 U2965 ( .A(n3714), .ZN(n5594) );
  AOI22_X1 U2966 ( .A1(\mem[129][2] ), .A2(n3712), .B1(n6739), .B2(data_in[2]), 
        .ZN(n3714) );
  INV_X1 U2967 ( .A(n3715), .ZN(n5593) );
  AOI22_X1 U2968 ( .A1(\mem[129][3] ), .A2(n3712), .B1(n6739), .B2(data_in[3]), 
        .ZN(n3715) );
  INV_X1 U2969 ( .A(n3716), .ZN(n5592) );
  AOI22_X1 U2970 ( .A1(\mem[129][4] ), .A2(n3712), .B1(n6739), .B2(data_in[4]), 
        .ZN(n3716) );
  INV_X1 U2971 ( .A(n3717), .ZN(n5591) );
  AOI22_X1 U2972 ( .A1(\mem[129][5] ), .A2(n3712), .B1(n6739), .B2(data_in[5]), 
        .ZN(n3717) );
  INV_X1 U2973 ( .A(n3718), .ZN(n5590) );
  AOI22_X1 U2974 ( .A1(\mem[129][6] ), .A2(n3712), .B1(n6739), .B2(data_in[6]), 
        .ZN(n3718) );
  INV_X1 U2975 ( .A(n3719), .ZN(n5589) );
  AOI22_X1 U2976 ( .A1(\mem[129][7] ), .A2(n3712), .B1(n6739), .B2(data_in[7]), 
        .ZN(n3719) );
  INV_X1 U2977 ( .A(n3720), .ZN(n5588) );
  AOI22_X1 U2978 ( .A1(\mem[130][0] ), .A2(n3721), .B1(n6738), .B2(data_in[0]), 
        .ZN(n3720) );
  INV_X1 U2979 ( .A(n3722), .ZN(n5587) );
  AOI22_X1 U2980 ( .A1(\mem[130][1] ), .A2(n3721), .B1(n6738), .B2(data_in[1]), 
        .ZN(n3722) );
  INV_X1 U2981 ( .A(n3723), .ZN(n5586) );
  AOI22_X1 U2982 ( .A1(\mem[130][2] ), .A2(n3721), .B1(n6738), .B2(data_in[2]), 
        .ZN(n3723) );
  INV_X1 U2983 ( .A(n3724), .ZN(n5585) );
  AOI22_X1 U2984 ( .A1(\mem[130][3] ), .A2(n3721), .B1(n6738), .B2(data_in[3]), 
        .ZN(n3724) );
  INV_X1 U2985 ( .A(n3725), .ZN(n5584) );
  AOI22_X1 U2986 ( .A1(\mem[130][4] ), .A2(n3721), .B1(n6738), .B2(data_in[4]), 
        .ZN(n3725) );
  INV_X1 U2987 ( .A(n3726), .ZN(n5583) );
  AOI22_X1 U2988 ( .A1(\mem[130][5] ), .A2(n3721), .B1(n6738), .B2(data_in[5]), 
        .ZN(n3726) );
  INV_X1 U2989 ( .A(n3727), .ZN(n5582) );
  AOI22_X1 U2990 ( .A1(\mem[130][6] ), .A2(n3721), .B1(n6738), .B2(data_in[6]), 
        .ZN(n3727) );
  INV_X1 U2991 ( .A(n3728), .ZN(n5581) );
  AOI22_X1 U2992 ( .A1(\mem[130][7] ), .A2(n3721), .B1(n6738), .B2(data_in[7]), 
        .ZN(n3728) );
  INV_X1 U2993 ( .A(n3729), .ZN(n5580) );
  AOI22_X1 U2994 ( .A1(\mem[131][0] ), .A2(n3730), .B1(n6737), .B2(data_in[0]), 
        .ZN(n3729) );
  INV_X1 U2995 ( .A(n3731), .ZN(n5579) );
  AOI22_X1 U2996 ( .A1(\mem[131][1] ), .A2(n3730), .B1(n6737), .B2(data_in[1]), 
        .ZN(n3731) );
  INV_X1 U2997 ( .A(n3732), .ZN(n5578) );
  AOI22_X1 U2998 ( .A1(\mem[131][2] ), .A2(n3730), .B1(n6737), .B2(data_in[2]), 
        .ZN(n3732) );
  INV_X1 U2999 ( .A(n3733), .ZN(n5577) );
  AOI22_X1 U3000 ( .A1(\mem[131][3] ), .A2(n3730), .B1(n6737), .B2(data_in[3]), 
        .ZN(n3733) );
  INV_X1 U3001 ( .A(n3734), .ZN(n5576) );
  AOI22_X1 U3002 ( .A1(\mem[131][4] ), .A2(n3730), .B1(n6737), .B2(data_in[4]), 
        .ZN(n3734) );
  INV_X1 U3003 ( .A(n3735), .ZN(n5575) );
  AOI22_X1 U3004 ( .A1(\mem[131][5] ), .A2(n3730), .B1(n6737), .B2(data_in[5]), 
        .ZN(n3735) );
  INV_X1 U3005 ( .A(n3736), .ZN(n5574) );
  AOI22_X1 U3006 ( .A1(\mem[131][6] ), .A2(n3730), .B1(n6737), .B2(data_in[6]), 
        .ZN(n3736) );
  INV_X1 U3007 ( .A(n3737), .ZN(n5573) );
  AOI22_X1 U3008 ( .A1(\mem[131][7] ), .A2(n3730), .B1(n6737), .B2(data_in[7]), 
        .ZN(n3737) );
  INV_X1 U3009 ( .A(n3738), .ZN(n5572) );
  AOI22_X1 U3010 ( .A1(\mem[132][0] ), .A2(n3739), .B1(n6736), .B2(data_in[0]), 
        .ZN(n3738) );
  INV_X1 U3011 ( .A(n3740), .ZN(n5571) );
  AOI22_X1 U3012 ( .A1(\mem[132][1] ), .A2(n3739), .B1(n6736), .B2(data_in[1]), 
        .ZN(n3740) );
  INV_X1 U3013 ( .A(n3741), .ZN(n5570) );
  AOI22_X1 U3014 ( .A1(\mem[132][2] ), .A2(n3739), .B1(n6736), .B2(data_in[2]), 
        .ZN(n3741) );
  INV_X1 U3015 ( .A(n3742), .ZN(n5569) );
  AOI22_X1 U3016 ( .A1(\mem[132][3] ), .A2(n3739), .B1(n6736), .B2(data_in[3]), 
        .ZN(n3742) );
  INV_X1 U3017 ( .A(n3743), .ZN(n5568) );
  AOI22_X1 U3018 ( .A1(\mem[132][4] ), .A2(n3739), .B1(n6736), .B2(data_in[4]), 
        .ZN(n3743) );
  INV_X1 U3019 ( .A(n3744), .ZN(n5567) );
  AOI22_X1 U3020 ( .A1(\mem[132][5] ), .A2(n3739), .B1(n6736), .B2(data_in[5]), 
        .ZN(n3744) );
  INV_X1 U3021 ( .A(n3745), .ZN(n5566) );
  AOI22_X1 U3022 ( .A1(\mem[132][6] ), .A2(n3739), .B1(n6736), .B2(data_in[6]), 
        .ZN(n3745) );
  INV_X1 U3023 ( .A(n3746), .ZN(n5565) );
  AOI22_X1 U3024 ( .A1(\mem[132][7] ), .A2(n3739), .B1(n6736), .B2(data_in[7]), 
        .ZN(n3746) );
  INV_X1 U3025 ( .A(n3747), .ZN(n5564) );
  AOI22_X1 U3026 ( .A1(\mem[133][0] ), .A2(n3748), .B1(n6735), .B2(data_in[0]), 
        .ZN(n3747) );
  INV_X1 U3027 ( .A(n3749), .ZN(n5563) );
  AOI22_X1 U3028 ( .A1(\mem[133][1] ), .A2(n3748), .B1(n6735), .B2(data_in[1]), 
        .ZN(n3749) );
  INV_X1 U3029 ( .A(n3750), .ZN(n5562) );
  AOI22_X1 U3030 ( .A1(\mem[133][2] ), .A2(n3748), .B1(n6735), .B2(data_in[2]), 
        .ZN(n3750) );
  INV_X1 U3031 ( .A(n3751), .ZN(n5561) );
  AOI22_X1 U3032 ( .A1(\mem[133][3] ), .A2(n3748), .B1(n6735), .B2(data_in[3]), 
        .ZN(n3751) );
  INV_X1 U3033 ( .A(n3752), .ZN(n5560) );
  AOI22_X1 U3034 ( .A1(\mem[133][4] ), .A2(n3748), .B1(n6735), .B2(data_in[4]), 
        .ZN(n3752) );
  INV_X1 U3035 ( .A(n3753), .ZN(n5559) );
  AOI22_X1 U3036 ( .A1(\mem[133][5] ), .A2(n3748), .B1(n6735), .B2(data_in[5]), 
        .ZN(n3753) );
  INV_X1 U3037 ( .A(n3754), .ZN(n5558) );
  AOI22_X1 U3038 ( .A1(\mem[133][6] ), .A2(n3748), .B1(n6735), .B2(data_in[6]), 
        .ZN(n3754) );
  INV_X1 U3039 ( .A(n3755), .ZN(n5557) );
  AOI22_X1 U3040 ( .A1(\mem[133][7] ), .A2(n3748), .B1(n6735), .B2(data_in[7]), 
        .ZN(n3755) );
  INV_X1 U3041 ( .A(n3756), .ZN(n5556) );
  AOI22_X1 U3042 ( .A1(\mem[134][0] ), .A2(n3757), .B1(n6734), .B2(data_in[0]), 
        .ZN(n3756) );
  INV_X1 U3043 ( .A(n3758), .ZN(n5555) );
  AOI22_X1 U3044 ( .A1(\mem[134][1] ), .A2(n3757), .B1(n6734), .B2(data_in[1]), 
        .ZN(n3758) );
  INV_X1 U3045 ( .A(n3759), .ZN(n5554) );
  AOI22_X1 U3046 ( .A1(\mem[134][2] ), .A2(n3757), .B1(n6734), .B2(data_in[2]), 
        .ZN(n3759) );
  INV_X1 U3047 ( .A(n3760), .ZN(n5553) );
  AOI22_X1 U3048 ( .A1(\mem[134][3] ), .A2(n3757), .B1(n6734), .B2(data_in[3]), 
        .ZN(n3760) );
  INV_X1 U3049 ( .A(n3761), .ZN(n5552) );
  AOI22_X1 U3050 ( .A1(\mem[134][4] ), .A2(n3757), .B1(n6734), .B2(data_in[4]), 
        .ZN(n3761) );
  INV_X1 U3051 ( .A(n3762), .ZN(n5551) );
  AOI22_X1 U3052 ( .A1(\mem[134][5] ), .A2(n3757), .B1(n6734), .B2(data_in[5]), 
        .ZN(n3762) );
  INV_X1 U3053 ( .A(n3763), .ZN(n5550) );
  AOI22_X1 U3054 ( .A1(\mem[134][6] ), .A2(n3757), .B1(n6734), .B2(data_in[6]), 
        .ZN(n3763) );
  INV_X1 U3055 ( .A(n3764), .ZN(n5549) );
  AOI22_X1 U3056 ( .A1(\mem[134][7] ), .A2(n3757), .B1(n6734), .B2(data_in[7]), 
        .ZN(n3764) );
  INV_X1 U3057 ( .A(n3765), .ZN(n5548) );
  AOI22_X1 U3058 ( .A1(\mem[135][0] ), .A2(n3766), .B1(n6733), .B2(data_in[0]), 
        .ZN(n3765) );
  INV_X1 U3059 ( .A(n3767), .ZN(n5547) );
  AOI22_X1 U3060 ( .A1(\mem[135][1] ), .A2(n3766), .B1(n6733), .B2(data_in[1]), 
        .ZN(n3767) );
  INV_X1 U3061 ( .A(n3768), .ZN(n5546) );
  AOI22_X1 U3062 ( .A1(\mem[135][2] ), .A2(n3766), .B1(n6733), .B2(data_in[2]), 
        .ZN(n3768) );
  INV_X1 U3063 ( .A(n3769), .ZN(n5545) );
  AOI22_X1 U3064 ( .A1(\mem[135][3] ), .A2(n3766), .B1(n6733), .B2(data_in[3]), 
        .ZN(n3769) );
  INV_X1 U3065 ( .A(n3770), .ZN(n5544) );
  AOI22_X1 U3066 ( .A1(\mem[135][4] ), .A2(n3766), .B1(n6733), .B2(data_in[4]), 
        .ZN(n3770) );
  INV_X1 U3067 ( .A(n3771), .ZN(n5543) );
  AOI22_X1 U3068 ( .A1(\mem[135][5] ), .A2(n3766), .B1(n6733), .B2(data_in[5]), 
        .ZN(n3771) );
  INV_X1 U3069 ( .A(n3772), .ZN(n5542) );
  AOI22_X1 U3070 ( .A1(\mem[135][6] ), .A2(n3766), .B1(n6733), .B2(data_in[6]), 
        .ZN(n3772) );
  INV_X1 U3071 ( .A(n3773), .ZN(n5541) );
  AOI22_X1 U3072 ( .A1(\mem[135][7] ), .A2(n3766), .B1(n6733), .B2(data_in[7]), 
        .ZN(n3773) );
  INV_X1 U3073 ( .A(n3774), .ZN(n5540) );
  AOI22_X1 U3074 ( .A1(\mem[136][0] ), .A2(n3775), .B1(n6732), .B2(data_in[0]), 
        .ZN(n3774) );
  INV_X1 U3075 ( .A(n3776), .ZN(n5539) );
  AOI22_X1 U3076 ( .A1(\mem[136][1] ), .A2(n3775), .B1(n6732), .B2(data_in[1]), 
        .ZN(n3776) );
  INV_X1 U3077 ( .A(n3777), .ZN(n5538) );
  AOI22_X1 U3078 ( .A1(\mem[136][2] ), .A2(n3775), .B1(n6732), .B2(data_in[2]), 
        .ZN(n3777) );
  INV_X1 U3079 ( .A(n3778), .ZN(n5537) );
  AOI22_X1 U3080 ( .A1(\mem[136][3] ), .A2(n3775), .B1(n6732), .B2(data_in[3]), 
        .ZN(n3778) );
  INV_X1 U3081 ( .A(n3779), .ZN(n5536) );
  AOI22_X1 U3082 ( .A1(\mem[136][4] ), .A2(n3775), .B1(n6732), .B2(data_in[4]), 
        .ZN(n3779) );
  INV_X1 U3083 ( .A(n3780), .ZN(n5535) );
  AOI22_X1 U3084 ( .A1(\mem[136][5] ), .A2(n3775), .B1(n6732), .B2(data_in[5]), 
        .ZN(n3780) );
  INV_X1 U3085 ( .A(n3781), .ZN(n5534) );
  AOI22_X1 U3086 ( .A1(\mem[136][6] ), .A2(n3775), .B1(n6732), .B2(data_in[6]), 
        .ZN(n3781) );
  INV_X1 U3087 ( .A(n3782), .ZN(n5533) );
  AOI22_X1 U3088 ( .A1(\mem[136][7] ), .A2(n3775), .B1(n6732), .B2(data_in[7]), 
        .ZN(n3782) );
  INV_X1 U3089 ( .A(n3783), .ZN(n5532) );
  AOI22_X1 U3090 ( .A1(\mem[137][0] ), .A2(n3784), .B1(n6731), .B2(data_in[0]), 
        .ZN(n3783) );
  INV_X1 U3091 ( .A(n3785), .ZN(n5531) );
  AOI22_X1 U3092 ( .A1(\mem[137][1] ), .A2(n3784), .B1(n6731), .B2(data_in[1]), 
        .ZN(n3785) );
  INV_X1 U3093 ( .A(n3786), .ZN(n5530) );
  AOI22_X1 U3094 ( .A1(\mem[137][2] ), .A2(n3784), .B1(n6731), .B2(data_in[2]), 
        .ZN(n3786) );
  INV_X1 U3095 ( .A(n3787), .ZN(n5529) );
  AOI22_X1 U3096 ( .A1(\mem[137][3] ), .A2(n3784), .B1(n6731), .B2(data_in[3]), 
        .ZN(n3787) );
  INV_X1 U3097 ( .A(n3788), .ZN(n5528) );
  AOI22_X1 U3098 ( .A1(\mem[137][4] ), .A2(n3784), .B1(n6731), .B2(data_in[4]), 
        .ZN(n3788) );
  INV_X1 U3099 ( .A(n3789), .ZN(n5527) );
  AOI22_X1 U3100 ( .A1(\mem[137][5] ), .A2(n3784), .B1(n6731), .B2(data_in[5]), 
        .ZN(n3789) );
  INV_X1 U3101 ( .A(n3790), .ZN(n5526) );
  AOI22_X1 U3102 ( .A1(\mem[137][6] ), .A2(n3784), .B1(n6731), .B2(data_in[6]), 
        .ZN(n3790) );
  INV_X1 U3103 ( .A(n3791), .ZN(n5525) );
  AOI22_X1 U3104 ( .A1(\mem[137][7] ), .A2(n3784), .B1(n6731), .B2(data_in[7]), 
        .ZN(n3791) );
  INV_X1 U3105 ( .A(n3792), .ZN(n5524) );
  AOI22_X1 U3106 ( .A1(\mem[138][0] ), .A2(n3793), .B1(n6730), .B2(data_in[0]), 
        .ZN(n3792) );
  INV_X1 U3107 ( .A(n3794), .ZN(n5523) );
  AOI22_X1 U3108 ( .A1(\mem[138][1] ), .A2(n3793), .B1(n6730), .B2(data_in[1]), 
        .ZN(n3794) );
  INV_X1 U3109 ( .A(n3795), .ZN(n5522) );
  AOI22_X1 U3110 ( .A1(\mem[138][2] ), .A2(n3793), .B1(n6730), .B2(data_in[2]), 
        .ZN(n3795) );
  INV_X1 U3111 ( .A(n3796), .ZN(n5521) );
  AOI22_X1 U3112 ( .A1(\mem[138][3] ), .A2(n3793), .B1(n6730), .B2(data_in[3]), 
        .ZN(n3796) );
  INV_X1 U3113 ( .A(n3797), .ZN(n5520) );
  AOI22_X1 U3114 ( .A1(\mem[138][4] ), .A2(n3793), .B1(n6730), .B2(data_in[4]), 
        .ZN(n3797) );
  INV_X1 U3115 ( .A(n3798), .ZN(n5519) );
  AOI22_X1 U3116 ( .A1(\mem[138][5] ), .A2(n3793), .B1(n6730), .B2(data_in[5]), 
        .ZN(n3798) );
  INV_X1 U3117 ( .A(n3799), .ZN(n5518) );
  AOI22_X1 U3118 ( .A1(\mem[138][6] ), .A2(n3793), .B1(n6730), .B2(data_in[6]), 
        .ZN(n3799) );
  INV_X1 U3119 ( .A(n3800), .ZN(n5517) );
  AOI22_X1 U3120 ( .A1(\mem[138][7] ), .A2(n3793), .B1(n6730), .B2(data_in[7]), 
        .ZN(n3800) );
  INV_X1 U3121 ( .A(n3801), .ZN(n5516) );
  AOI22_X1 U3122 ( .A1(\mem[139][0] ), .A2(n3802), .B1(n6729), .B2(data_in[0]), 
        .ZN(n3801) );
  INV_X1 U3123 ( .A(n3803), .ZN(n5515) );
  AOI22_X1 U3124 ( .A1(\mem[139][1] ), .A2(n3802), .B1(n6729), .B2(data_in[1]), 
        .ZN(n3803) );
  INV_X1 U3125 ( .A(n3804), .ZN(n5514) );
  AOI22_X1 U3126 ( .A1(\mem[139][2] ), .A2(n3802), .B1(n6729), .B2(data_in[2]), 
        .ZN(n3804) );
  INV_X1 U3127 ( .A(n3805), .ZN(n5513) );
  AOI22_X1 U3128 ( .A1(\mem[139][3] ), .A2(n3802), .B1(n6729), .B2(data_in[3]), 
        .ZN(n3805) );
  INV_X1 U3129 ( .A(n3806), .ZN(n5512) );
  AOI22_X1 U3130 ( .A1(\mem[139][4] ), .A2(n3802), .B1(n6729), .B2(data_in[4]), 
        .ZN(n3806) );
  INV_X1 U3131 ( .A(n3807), .ZN(n5511) );
  AOI22_X1 U3132 ( .A1(\mem[139][5] ), .A2(n3802), .B1(n6729), .B2(data_in[5]), 
        .ZN(n3807) );
  INV_X1 U3133 ( .A(n3808), .ZN(n5510) );
  AOI22_X1 U3134 ( .A1(\mem[139][6] ), .A2(n3802), .B1(n6729), .B2(data_in[6]), 
        .ZN(n3808) );
  INV_X1 U3135 ( .A(n3809), .ZN(n5509) );
  AOI22_X1 U3136 ( .A1(\mem[139][7] ), .A2(n3802), .B1(n6729), .B2(data_in[7]), 
        .ZN(n3809) );
  INV_X1 U3137 ( .A(n3810), .ZN(n5508) );
  AOI22_X1 U3138 ( .A1(\mem[140][0] ), .A2(n3811), .B1(n6728), .B2(data_in[0]), 
        .ZN(n3810) );
  INV_X1 U3139 ( .A(n3812), .ZN(n5507) );
  AOI22_X1 U3140 ( .A1(\mem[140][1] ), .A2(n3811), .B1(n6728), .B2(data_in[1]), 
        .ZN(n3812) );
  INV_X1 U3141 ( .A(n3813), .ZN(n5506) );
  AOI22_X1 U3142 ( .A1(\mem[140][2] ), .A2(n3811), .B1(n6728), .B2(data_in[2]), 
        .ZN(n3813) );
  INV_X1 U3143 ( .A(n3814), .ZN(n5505) );
  AOI22_X1 U3144 ( .A1(\mem[140][3] ), .A2(n3811), .B1(n6728), .B2(data_in[3]), 
        .ZN(n3814) );
  INV_X1 U3145 ( .A(n3815), .ZN(n5504) );
  AOI22_X1 U3146 ( .A1(\mem[140][4] ), .A2(n3811), .B1(n6728), .B2(data_in[4]), 
        .ZN(n3815) );
  INV_X1 U3147 ( .A(n3816), .ZN(n5503) );
  AOI22_X1 U3148 ( .A1(\mem[140][5] ), .A2(n3811), .B1(n6728), .B2(data_in[5]), 
        .ZN(n3816) );
  INV_X1 U3149 ( .A(n3817), .ZN(n5502) );
  AOI22_X1 U3150 ( .A1(\mem[140][6] ), .A2(n3811), .B1(n6728), .B2(data_in[6]), 
        .ZN(n3817) );
  INV_X1 U3151 ( .A(n3818), .ZN(n5501) );
  AOI22_X1 U3152 ( .A1(\mem[140][7] ), .A2(n3811), .B1(n6728), .B2(data_in[7]), 
        .ZN(n3818) );
  INV_X1 U3153 ( .A(n3819), .ZN(n5500) );
  AOI22_X1 U3154 ( .A1(\mem[141][0] ), .A2(n3820), .B1(n6727), .B2(data_in[0]), 
        .ZN(n3819) );
  INV_X1 U3155 ( .A(n3821), .ZN(n5499) );
  AOI22_X1 U3156 ( .A1(\mem[141][1] ), .A2(n3820), .B1(n6727), .B2(data_in[1]), 
        .ZN(n3821) );
  INV_X1 U3157 ( .A(n3822), .ZN(n5498) );
  AOI22_X1 U3158 ( .A1(\mem[141][2] ), .A2(n3820), .B1(n6727), .B2(data_in[2]), 
        .ZN(n3822) );
  INV_X1 U3159 ( .A(n3823), .ZN(n5497) );
  AOI22_X1 U3160 ( .A1(\mem[141][3] ), .A2(n3820), .B1(n6727), .B2(data_in[3]), 
        .ZN(n3823) );
  INV_X1 U3161 ( .A(n3824), .ZN(n5496) );
  AOI22_X1 U3162 ( .A1(\mem[141][4] ), .A2(n3820), .B1(n6727), .B2(data_in[4]), 
        .ZN(n3824) );
  INV_X1 U3163 ( .A(n3825), .ZN(n5495) );
  AOI22_X1 U3164 ( .A1(\mem[141][5] ), .A2(n3820), .B1(n6727), .B2(data_in[5]), 
        .ZN(n3825) );
  INV_X1 U3165 ( .A(n3826), .ZN(n5494) );
  AOI22_X1 U3166 ( .A1(\mem[141][6] ), .A2(n3820), .B1(n6727), .B2(data_in[6]), 
        .ZN(n3826) );
  INV_X1 U3167 ( .A(n3827), .ZN(n5493) );
  AOI22_X1 U3168 ( .A1(\mem[141][7] ), .A2(n3820), .B1(n6727), .B2(data_in[7]), 
        .ZN(n3827) );
  INV_X1 U3169 ( .A(n3828), .ZN(n5492) );
  AOI22_X1 U3170 ( .A1(\mem[142][0] ), .A2(n3829), .B1(n6726), .B2(data_in[0]), 
        .ZN(n3828) );
  INV_X1 U3171 ( .A(n3830), .ZN(n5491) );
  AOI22_X1 U3172 ( .A1(\mem[142][1] ), .A2(n3829), .B1(n6726), .B2(data_in[1]), 
        .ZN(n3830) );
  INV_X1 U3173 ( .A(n3831), .ZN(n5490) );
  AOI22_X1 U3174 ( .A1(\mem[142][2] ), .A2(n3829), .B1(n6726), .B2(data_in[2]), 
        .ZN(n3831) );
  INV_X1 U3175 ( .A(n3832), .ZN(n5489) );
  AOI22_X1 U3176 ( .A1(\mem[142][3] ), .A2(n3829), .B1(n6726), .B2(data_in[3]), 
        .ZN(n3832) );
  INV_X1 U3177 ( .A(n3833), .ZN(n5488) );
  AOI22_X1 U3178 ( .A1(\mem[142][4] ), .A2(n3829), .B1(n6726), .B2(data_in[4]), 
        .ZN(n3833) );
  INV_X1 U3179 ( .A(n3834), .ZN(n5487) );
  AOI22_X1 U3180 ( .A1(\mem[142][5] ), .A2(n3829), .B1(n6726), .B2(data_in[5]), 
        .ZN(n3834) );
  INV_X1 U3181 ( .A(n3835), .ZN(n5486) );
  AOI22_X1 U3182 ( .A1(\mem[142][6] ), .A2(n3829), .B1(n6726), .B2(data_in[6]), 
        .ZN(n3835) );
  INV_X1 U3183 ( .A(n3836), .ZN(n5485) );
  AOI22_X1 U3184 ( .A1(\mem[142][7] ), .A2(n3829), .B1(n6726), .B2(data_in[7]), 
        .ZN(n3836) );
  INV_X1 U3185 ( .A(n3837), .ZN(n5484) );
  AOI22_X1 U3186 ( .A1(\mem[143][0] ), .A2(n3838), .B1(n6725), .B2(data_in[0]), 
        .ZN(n3837) );
  INV_X1 U3187 ( .A(n3839), .ZN(n5483) );
  AOI22_X1 U3188 ( .A1(\mem[143][1] ), .A2(n3838), .B1(n6725), .B2(data_in[1]), 
        .ZN(n3839) );
  INV_X1 U3189 ( .A(n3840), .ZN(n5482) );
  AOI22_X1 U3190 ( .A1(\mem[143][2] ), .A2(n3838), .B1(n6725), .B2(data_in[2]), 
        .ZN(n3840) );
  INV_X1 U3191 ( .A(n3841), .ZN(n5481) );
  AOI22_X1 U3192 ( .A1(\mem[143][3] ), .A2(n3838), .B1(n6725), .B2(data_in[3]), 
        .ZN(n3841) );
  INV_X1 U3193 ( .A(n3842), .ZN(n5480) );
  AOI22_X1 U3194 ( .A1(\mem[143][4] ), .A2(n3838), .B1(n6725), .B2(data_in[4]), 
        .ZN(n3842) );
  INV_X1 U3195 ( .A(n3843), .ZN(n5479) );
  AOI22_X1 U3196 ( .A1(\mem[143][5] ), .A2(n3838), .B1(n6725), .B2(data_in[5]), 
        .ZN(n3843) );
  INV_X1 U3197 ( .A(n3844), .ZN(n5478) );
  AOI22_X1 U3198 ( .A1(\mem[143][6] ), .A2(n3838), .B1(n6725), .B2(data_in[6]), 
        .ZN(n3844) );
  INV_X1 U3199 ( .A(n3845), .ZN(n5477) );
  AOI22_X1 U3200 ( .A1(\mem[143][7] ), .A2(n3838), .B1(n6725), .B2(data_in[7]), 
        .ZN(n3845) );
  INV_X1 U3201 ( .A(n3847), .ZN(n5476) );
  AOI22_X1 U3202 ( .A1(\mem[144][0] ), .A2(n3848), .B1(n6724), .B2(data_in[0]), 
        .ZN(n3847) );
  INV_X1 U3203 ( .A(n3849), .ZN(n5475) );
  AOI22_X1 U3204 ( .A1(\mem[144][1] ), .A2(n3848), .B1(n6724), .B2(data_in[1]), 
        .ZN(n3849) );
  INV_X1 U3205 ( .A(n3850), .ZN(n5474) );
  AOI22_X1 U3206 ( .A1(\mem[144][2] ), .A2(n3848), .B1(n6724), .B2(data_in[2]), 
        .ZN(n3850) );
  INV_X1 U3207 ( .A(n3851), .ZN(n5473) );
  AOI22_X1 U3208 ( .A1(\mem[144][3] ), .A2(n3848), .B1(n6724), .B2(data_in[3]), 
        .ZN(n3851) );
  INV_X1 U3209 ( .A(n3852), .ZN(n5472) );
  AOI22_X1 U3210 ( .A1(\mem[144][4] ), .A2(n3848), .B1(n6724), .B2(data_in[4]), 
        .ZN(n3852) );
  INV_X1 U3211 ( .A(n3853), .ZN(n5471) );
  AOI22_X1 U3212 ( .A1(\mem[144][5] ), .A2(n3848), .B1(n6724), .B2(data_in[5]), 
        .ZN(n3853) );
  INV_X1 U3213 ( .A(n3854), .ZN(n5470) );
  AOI22_X1 U3214 ( .A1(\mem[144][6] ), .A2(n3848), .B1(n6724), .B2(data_in[6]), 
        .ZN(n3854) );
  INV_X1 U3215 ( .A(n3855), .ZN(n5469) );
  AOI22_X1 U3216 ( .A1(\mem[144][7] ), .A2(n3848), .B1(n6724), .B2(data_in[7]), 
        .ZN(n3855) );
  INV_X1 U3217 ( .A(n3857), .ZN(n5468) );
  AOI22_X1 U3218 ( .A1(\mem[145][0] ), .A2(n3858), .B1(n6723), .B2(data_in[0]), 
        .ZN(n3857) );
  INV_X1 U3219 ( .A(n3859), .ZN(n5467) );
  AOI22_X1 U3220 ( .A1(\mem[145][1] ), .A2(n3858), .B1(n6723), .B2(data_in[1]), 
        .ZN(n3859) );
  INV_X1 U3221 ( .A(n3860), .ZN(n5466) );
  AOI22_X1 U3222 ( .A1(\mem[145][2] ), .A2(n3858), .B1(n6723), .B2(data_in[2]), 
        .ZN(n3860) );
  INV_X1 U3223 ( .A(n3861), .ZN(n5465) );
  AOI22_X1 U3224 ( .A1(\mem[145][3] ), .A2(n3858), .B1(n6723), .B2(data_in[3]), 
        .ZN(n3861) );
  INV_X1 U3225 ( .A(n3862), .ZN(n5464) );
  AOI22_X1 U3226 ( .A1(\mem[145][4] ), .A2(n3858), .B1(n6723), .B2(data_in[4]), 
        .ZN(n3862) );
  INV_X1 U3227 ( .A(n3863), .ZN(n5463) );
  AOI22_X1 U3228 ( .A1(\mem[145][5] ), .A2(n3858), .B1(n6723), .B2(data_in[5]), 
        .ZN(n3863) );
  INV_X1 U3229 ( .A(n3864), .ZN(n5462) );
  AOI22_X1 U3230 ( .A1(\mem[145][6] ), .A2(n3858), .B1(n6723), .B2(data_in[6]), 
        .ZN(n3864) );
  INV_X1 U3231 ( .A(n3865), .ZN(n5461) );
  AOI22_X1 U3232 ( .A1(\mem[145][7] ), .A2(n3858), .B1(n6723), .B2(data_in[7]), 
        .ZN(n3865) );
  INV_X1 U3233 ( .A(n3866), .ZN(n5460) );
  AOI22_X1 U3234 ( .A1(\mem[146][0] ), .A2(n3867), .B1(n6722), .B2(data_in[0]), 
        .ZN(n3866) );
  INV_X1 U3235 ( .A(n3868), .ZN(n5459) );
  AOI22_X1 U3236 ( .A1(\mem[146][1] ), .A2(n3867), .B1(n6722), .B2(data_in[1]), 
        .ZN(n3868) );
  INV_X1 U3237 ( .A(n3869), .ZN(n5458) );
  AOI22_X1 U3238 ( .A1(\mem[146][2] ), .A2(n3867), .B1(n6722), .B2(data_in[2]), 
        .ZN(n3869) );
  INV_X1 U3239 ( .A(n3870), .ZN(n5457) );
  AOI22_X1 U3240 ( .A1(\mem[146][3] ), .A2(n3867), .B1(n6722), .B2(data_in[3]), 
        .ZN(n3870) );
  INV_X1 U3241 ( .A(n3871), .ZN(n5456) );
  AOI22_X1 U3242 ( .A1(\mem[146][4] ), .A2(n3867), .B1(n6722), .B2(data_in[4]), 
        .ZN(n3871) );
  INV_X1 U3243 ( .A(n3872), .ZN(n5455) );
  AOI22_X1 U3244 ( .A1(\mem[146][5] ), .A2(n3867), .B1(n6722), .B2(data_in[5]), 
        .ZN(n3872) );
  INV_X1 U3245 ( .A(n3873), .ZN(n5454) );
  AOI22_X1 U3246 ( .A1(\mem[146][6] ), .A2(n3867), .B1(n6722), .B2(data_in[6]), 
        .ZN(n3873) );
  INV_X1 U3247 ( .A(n3874), .ZN(n5453) );
  AOI22_X1 U3248 ( .A1(\mem[146][7] ), .A2(n3867), .B1(n6722), .B2(data_in[7]), 
        .ZN(n3874) );
  INV_X1 U3249 ( .A(n3875), .ZN(n5452) );
  AOI22_X1 U3250 ( .A1(\mem[147][0] ), .A2(n3876), .B1(n6721), .B2(data_in[0]), 
        .ZN(n3875) );
  INV_X1 U3251 ( .A(n3877), .ZN(n5451) );
  AOI22_X1 U3252 ( .A1(\mem[147][1] ), .A2(n3876), .B1(n6721), .B2(data_in[1]), 
        .ZN(n3877) );
  INV_X1 U3253 ( .A(n3878), .ZN(n5450) );
  AOI22_X1 U3254 ( .A1(\mem[147][2] ), .A2(n3876), .B1(n6721), .B2(data_in[2]), 
        .ZN(n3878) );
  INV_X1 U3255 ( .A(n3879), .ZN(n5449) );
  AOI22_X1 U3256 ( .A1(\mem[147][3] ), .A2(n3876), .B1(n6721), .B2(data_in[3]), 
        .ZN(n3879) );
  INV_X1 U3257 ( .A(n3880), .ZN(n5448) );
  AOI22_X1 U3258 ( .A1(\mem[147][4] ), .A2(n3876), .B1(n6721), .B2(data_in[4]), 
        .ZN(n3880) );
  INV_X1 U3259 ( .A(n3881), .ZN(n5447) );
  AOI22_X1 U3260 ( .A1(\mem[147][5] ), .A2(n3876), .B1(n6721), .B2(data_in[5]), 
        .ZN(n3881) );
  INV_X1 U3261 ( .A(n3882), .ZN(n5446) );
  AOI22_X1 U3262 ( .A1(\mem[147][6] ), .A2(n3876), .B1(n6721), .B2(data_in[6]), 
        .ZN(n3882) );
  INV_X1 U3263 ( .A(n3883), .ZN(n5445) );
  AOI22_X1 U3264 ( .A1(\mem[147][7] ), .A2(n3876), .B1(n6721), .B2(data_in[7]), 
        .ZN(n3883) );
  INV_X1 U3265 ( .A(n3884), .ZN(n5444) );
  AOI22_X1 U3266 ( .A1(\mem[148][0] ), .A2(n3885), .B1(n6720), .B2(data_in[0]), 
        .ZN(n3884) );
  INV_X1 U3267 ( .A(n3886), .ZN(n5443) );
  AOI22_X1 U3268 ( .A1(\mem[148][1] ), .A2(n3885), .B1(n6720), .B2(data_in[1]), 
        .ZN(n3886) );
  INV_X1 U3269 ( .A(n3887), .ZN(n5442) );
  AOI22_X1 U3270 ( .A1(\mem[148][2] ), .A2(n3885), .B1(n6720), .B2(data_in[2]), 
        .ZN(n3887) );
  INV_X1 U3271 ( .A(n3888), .ZN(n5441) );
  AOI22_X1 U3272 ( .A1(\mem[148][3] ), .A2(n3885), .B1(n6720), .B2(data_in[3]), 
        .ZN(n3888) );
  INV_X1 U3273 ( .A(n3889), .ZN(n5440) );
  AOI22_X1 U3274 ( .A1(\mem[148][4] ), .A2(n3885), .B1(n6720), .B2(data_in[4]), 
        .ZN(n3889) );
  INV_X1 U3275 ( .A(n3890), .ZN(n5439) );
  AOI22_X1 U3276 ( .A1(\mem[148][5] ), .A2(n3885), .B1(n6720), .B2(data_in[5]), 
        .ZN(n3890) );
  INV_X1 U3277 ( .A(n3891), .ZN(n5438) );
  AOI22_X1 U3278 ( .A1(\mem[148][6] ), .A2(n3885), .B1(n6720), .B2(data_in[6]), 
        .ZN(n3891) );
  INV_X1 U3279 ( .A(n3892), .ZN(n5437) );
  AOI22_X1 U3280 ( .A1(\mem[148][7] ), .A2(n3885), .B1(n6720), .B2(data_in[7]), 
        .ZN(n3892) );
  INV_X1 U3281 ( .A(n3893), .ZN(n5436) );
  AOI22_X1 U3282 ( .A1(\mem[149][0] ), .A2(n3894), .B1(n6719), .B2(data_in[0]), 
        .ZN(n3893) );
  INV_X1 U3283 ( .A(n3895), .ZN(n5435) );
  AOI22_X1 U3284 ( .A1(\mem[149][1] ), .A2(n3894), .B1(n6719), .B2(data_in[1]), 
        .ZN(n3895) );
  INV_X1 U3285 ( .A(n3896), .ZN(n5434) );
  AOI22_X1 U3286 ( .A1(\mem[149][2] ), .A2(n3894), .B1(n6719), .B2(data_in[2]), 
        .ZN(n3896) );
  INV_X1 U3287 ( .A(n3897), .ZN(n5433) );
  AOI22_X1 U3288 ( .A1(\mem[149][3] ), .A2(n3894), .B1(n6719), .B2(data_in[3]), 
        .ZN(n3897) );
  INV_X1 U3289 ( .A(n3898), .ZN(n5432) );
  AOI22_X1 U3290 ( .A1(\mem[149][4] ), .A2(n3894), .B1(n6719), .B2(data_in[4]), 
        .ZN(n3898) );
  INV_X1 U3291 ( .A(n3899), .ZN(n5431) );
  AOI22_X1 U3292 ( .A1(\mem[149][5] ), .A2(n3894), .B1(n6719), .B2(data_in[5]), 
        .ZN(n3899) );
  INV_X1 U3293 ( .A(n3900), .ZN(n5430) );
  AOI22_X1 U3294 ( .A1(\mem[149][6] ), .A2(n3894), .B1(n6719), .B2(data_in[6]), 
        .ZN(n3900) );
  INV_X1 U3295 ( .A(n3901), .ZN(n5429) );
  AOI22_X1 U3296 ( .A1(\mem[149][7] ), .A2(n3894), .B1(n6719), .B2(data_in[7]), 
        .ZN(n3901) );
  INV_X1 U3297 ( .A(n3902), .ZN(n5428) );
  AOI22_X1 U3298 ( .A1(\mem[150][0] ), .A2(n3903), .B1(n6718), .B2(data_in[0]), 
        .ZN(n3902) );
  INV_X1 U3299 ( .A(n3904), .ZN(n5427) );
  AOI22_X1 U3300 ( .A1(\mem[150][1] ), .A2(n3903), .B1(n6718), .B2(data_in[1]), 
        .ZN(n3904) );
  INV_X1 U3301 ( .A(n3905), .ZN(n5426) );
  AOI22_X1 U3302 ( .A1(\mem[150][2] ), .A2(n3903), .B1(n6718), .B2(data_in[2]), 
        .ZN(n3905) );
  INV_X1 U3303 ( .A(n3906), .ZN(n5425) );
  AOI22_X1 U3304 ( .A1(\mem[150][3] ), .A2(n3903), .B1(n6718), .B2(data_in[3]), 
        .ZN(n3906) );
  INV_X1 U3305 ( .A(n3907), .ZN(n5424) );
  AOI22_X1 U3306 ( .A1(\mem[150][4] ), .A2(n3903), .B1(n6718), .B2(data_in[4]), 
        .ZN(n3907) );
  INV_X1 U3307 ( .A(n3908), .ZN(n5423) );
  AOI22_X1 U3308 ( .A1(\mem[150][5] ), .A2(n3903), .B1(n6718), .B2(data_in[5]), 
        .ZN(n3908) );
  INV_X1 U3309 ( .A(n3909), .ZN(n5422) );
  AOI22_X1 U3310 ( .A1(\mem[150][6] ), .A2(n3903), .B1(n6718), .B2(data_in[6]), 
        .ZN(n3909) );
  INV_X1 U3311 ( .A(n3910), .ZN(n5421) );
  AOI22_X1 U3312 ( .A1(\mem[150][7] ), .A2(n3903), .B1(n6718), .B2(data_in[7]), 
        .ZN(n3910) );
  INV_X1 U3313 ( .A(n3911), .ZN(n5420) );
  AOI22_X1 U3314 ( .A1(\mem[151][0] ), .A2(n3912), .B1(n6717), .B2(data_in[0]), 
        .ZN(n3911) );
  INV_X1 U3315 ( .A(n3913), .ZN(n5419) );
  AOI22_X1 U3316 ( .A1(\mem[151][1] ), .A2(n3912), .B1(n6717), .B2(data_in[1]), 
        .ZN(n3913) );
  INV_X1 U3317 ( .A(n3914), .ZN(n5418) );
  AOI22_X1 U3318 ( .A1(\mem[151][2] ), .A2(n3912), .B1(n6717), .B2(data_in[2]), 
        .ZN(n3914) );
  INV_X1 U3319 ( .A(n3915), .ZN(n5417) );
  AOI22_X1 U3320 ( .A1(\mem[151][3] ), .A2(n3912), .B1(n6717), .B2(data_in[3]), 
        .ZN(n3915) );
  INV_X1 U3321 ( .A(n3916), .ZN(n5416) );
  AOI22_X1 U3322 ( .A1(\mem[151][4] ), .A2(n3912), .B1(n6717), .B2(data_in[4]), 
        .ZN(n3916) );
  INV_X1 U3323 ( .A(n3917), .ZN(n5415) );
  AOI22_X1 U3324 ( .A1(\mem[151][5] ), .A2(n3912), .B1(n6717), .B2(data_in[5]), 
        .ZN(n3917) );
  INV_X1 U3325 ( .A(n3918), .ZN(n5414) );
  AOI22_X1 U3326 ( .A1(\mem[151][6] ), .A2(n3912), .B1(n6717), .B2(data_in[6]), 
        .ZN(n3918) );
  INV_X1 U3327 ( .A(n3919), .ZN(n5413) );
  AOI22_X1 U3328 ( .A1(\mem[151][7] ), .A2(n3912), .B1(n6717), .B2(data_in[7]), 
        .ZN(n3919) );
  INV_X1 U3329 ( .A(n3920), .ZN(n5412) );
  AOI22_X1 U3330 ( .A1(\mem[152][0] ), .A2(n3921), .B1(n6716), .B2(data_in[0]), 
        .ZN(n3920) );
  INV_X1 U3331 ( .A(n3922), .ZN(n5411) );
  AOI22_X1 U3332 ( .A1(\mem[152][1] ), .A2(n3921), .B1(n6716), .B2(data_in[1]), 
        .ZN(n3922) );
  INV_X1 U3333 ( .A(n3923), .ZN(n5410) );
  AOI22_X1 U3334 ( .A1(\mem[152][2] ), .A2(n3921), .B1(n6716), .B2(data_in[2]), 
        .ZN(n3923) );
  INV_X1 U3335 ( .A(n3924), .ZN(n5409) );
  AOI22_X1 U3336 ( .A1(\mem[152][3] ), .A2(n3921), .B1(n6716), .B2(data_in[3]), 
        .ZN(n3924) );
  INV_X1 U3337 ( .A(n3925), .ZN(n5408) );
  AOI22_X1 U3338 ( .A1(\mem[152][4] ), .A2(n3921), .B1(n6716), .B2(data_in[4]), 
        .ZN(n3925) );
  INV_X1 U3339 ( .A(n3926), .ZN(n5407) );
  AOI22_X1 U3340 ( .A1(\mem[152][5] ), .A2(n3921), .B1(n6716), .B2(data_in[5]), 
        .ZN(n3926) );
  INV_X1 U3341 ( .A(n3927), .ZN(n5406) );
  AOI22_X1 U3342 ( .A1(\mem[152][6] ), .A2(n3921), .B1(n6716), .B2(data_in[6]), 
        .ZN(n3927) );
  INV_X1 U3343 ( .A(n3928), .ZN(n5405) );
  AOI22_X1 U3344 ( .A1(\mem[152][7] ), .A2(n3921), .B1(n6716), .B2(data_in[7]), 
        .ZN(n3928) );
  INV_X1 U3345 ( .A(n3929), .ZN(n5404) );
  AOI22_X1 U3346 ( .A1(\mem[153][0] ), .A2(n3930), .B1(n6715), .B2(data_in[0]), 
        .ZN(n3929) );
  INV_X1 U3347 ( .A(n3931), .ZN(n5403) );
  AOI22_X1 U3348 ( .A1(\mem[153][1] ), .A2(n3930), .B1(n6715), .B2(data_in[1]), 
        .ZN(n3931) );
  INV_X1 U3349 ( .A(n3932), .ZN(n5402) );
  AOI22_X1 U3350 ( .A1(\mem[153][2] ), .A2(n3930), .B1(n6715), .B2(data_in[2]), 
        .ZN(n3932) );
  INV_X1 U3351 ( .A(n3933), .ZN(n5401) );
  AOI22_X1 U3352 ( .A1(\mem[153][3] ), .A2(n3930), .B1(n6715), .B2(data_in[3]), 
        .ZN(n3933) );
  INV_X1 U3353 ( .A(n3934), .ZN(n5400) );
  AOI22_X1 U3354 ( .A1(\mem[153][4] ), .A2(n3930), .B1(n6715), .B2(data_in[4]), 
        .ZN(n3934) );
  INV_X1 U3355 ( .A(n3935), .ZN(n5399) );
  AOI22_X1 U3356 ( .A1(\mem[153][5] ), .A2(n3930), .B1(n6715), .B2(data_in[5]), 
        .ZN(n3935) );
  INV_X1 U3357 ( .A(n3936), .ZN(n5398) );
  AOI22_X1 U3358 ( .A1(\mem[153][6] ), .A2(n3930), .B1(n6715), .B2(data_in[6]), 
        .ZN(n3936) );
  INV_X1 U3359 ( .A(n3937), .ZN(n5397) );
  AOI22_X1 U3360 ( .A1(\mem[153][7] ), .A2(n3930), .B1(n6715), .B2(data_in[7]), 
        .ZN(n3937) );
  INV_X1 U3361 ( .A(n3938), .ZN(n5396) );
  AOI22_X1 U3362 ( .A1(\mem[154][0] ), .A2(n3939), .B1(n6714), .B2(data_in[0]), 
        .ZN(n3938) );
  INV_X1 U3363 ( .A(n3940), .ZN(n5395) );
  AOI22_X1 U3364 ( .A1(\mem[154][1] ), .A2(n3939), .B1(n6714), .B2(data_in[1]), 
        .ZN(n3940) );
  INV_X1 U3365 ( .A(n3941), .ZN(n5394) );
  AOI22_X1 U3366 ( .A1(\mem[154][2] ), .A2(n3939), .B1(n6714), .B2(data_in[2]), 
        .ZN(n3941) );
  INV_X1 U3367 ( .A(n3942), .ZN(n5393) );
  AOI22_X1 U3368 ( .A1(\mem[154][3] ), .A2(n3939), .B1(n6714), .B2(data_in[3]), 
        .ZN(n3942) );
  INV_X1 U3369 ( .A(n3943), .ZN(n5392) );
  AOI22_X1 U3370 ( .A1(\mem[154][4] ), .A2(n3939), .B1(n6714), .B2(data_in[4]), 
        .ZN(n3943) );
  INV_X1 U3371 ( .A(n3944), .ZN(n5391) );
  AOI22_X1 U3372 ( .A1(\mem[154][5] ), .A2(n3939), .B1(n6714), .B2(data_in[5]), 
        .ZN(n3944) );
  INV_X1 U3373 ( .A(n3945), .ZN(n5390) );
  AOI22_X1 U3374 ( .A1(\mem[154][6] ), .A2(n3939), .B1(n6714), .B2(data_in[6]), 
        .ZN(n3945) );
  INV_X1 U3375 ( .A(n3946), .ZN(n5389) );
  AOI22_X1 U3376 ( .A1(\mem[154][7] ), .A2(n3939), .B1(n6714), .B2(data_in[7]), 
        .ZN(n3946) );
  INV_X1 U3377 ( .A(n3947), .ZN(n5388) );
  AOI22_X1 U3378 ( .A1(\mem[155][0] ), .A2(n3948), .B1(n6713), .B2(data_in[0]), 
        .ZN(n3947) );
  INV_X1 U3379 ( .A(n3949), .ZN(n5387) );
  AOI22_X1 U3380 ( .A1(\mem[155][1] ), .A2(n3948), .B1(n6713), .B2(data_in[1]), 
        .ZN(n3949) );
  INV_X1 U3381 ( .A(n3950), .ZN(n5386) );
  AOI22_X1 U3382 ( .A1(\mem[155][2] ), .A2(n3948), .B1(n6713), .B2(data_in[2]), 
        .ZN(n3950) );
  INV_X1 U3383 ( .A(n3951), .ZN(n5385) );
  AOI22_X1 U3384 ( .A1(\mem[155][3] ), .A2(n3948), .B1(n6713), .B2(data_in[3]), 
        .ZN(n3951) );
  INV_X1 U3385 ( .A(n3952), .ZN(n5384) );
  AOI22_X1 U3386 ( .A1(\mem[155][4] ), .A2(n3948), .B1(n6713), .B2(data_in[4]), 
        .ZN(n3952) );
  INV_X1 U3387 ( .A(n3953), .ZN(n5383) );
  AOI22_X1 U3388 ( .A1(\mem[155][5] ), .A2(n3948), .B1(n6713), .B2(data_in[5]), 
        .ZN(n3953) );
  INV_X1 U3389 ( .A(n3954), .ZN(n5382) );
  AOI22_X1 U3390 ( .A1(\mem[155][6] ), .A2(n3948), .B1(n6713), .B2(data_in[6]), 
        .ZN(n3954) );
  INV_X1 U3391 ( .A(n3955), .ZN(n5381) );
  AOI22_X1 U3392 ( .A1(\mem[155][7] ), .A2(n3948), .B1(n6713), .B2(data_in[7]), 
        .ZN(n3955) );
  INV_X1 U3393 ( .A(n3956), .ZN(n5380) );
  AOI22_X1 U3394 ( .A1(\mem[156][0] ), .A2(n3957), .B1(n6712), .B2(data_in[0]), 
        .ZN(n3956) );
  INV_X1 U3395 ( .A(n3958), .ZN(n5379) );
  AOI22_X1 U3396 ( .A1(\mem[156][1] ), .A2(n3957), .B1(n6712), .B2(data_in[1]), 
        .ZN(n3958) );
  INV_X1 U3397 ( .A(n3959), .ZN(n5378) );
  AOI22_X1 U3398 ( .A1(\mem[156][2] ), .A2(n3957), .B1(n6712), .B2(data_in[2]), 
        .ZN(n3959) );
  INV_X1 U3399 ( .A(n3960), .ZN(n5377) );
  AOI22_X1 U3400 ( .A1(\mem[156][3] ), .A2(n3957), .B1(n6712), .B2(data_in[3]), 
        .ZN(n3960) );
  INV_X1 U3401 ( .A(n3961), .ZN(n5376) );
  AOI22_X1 U3402 ( .A1(\mem[156][4] ), .A2(n3957), .B1(n6712), .B2(data_in[4]), 
        .ZN(n3961) );
  INV_X1 U3403 ( .A(n3962), .ZN(n5375) );
  AOI22_X1 U3404 ( .A1(\mem[156][5] ), .A2(n3957), .B1(n6712), .B2(data_in[5]), 
        .ZN(n3962) );
  INV_X1 U3405 ( .A(n3963), .ZN(n5374) );
  AOI22_X1 U3406 ( .A1(\mem[156][6] ), .A2(n3957), .B1(n6712), .B2(data_in[6]), 
        .ZN(n3963) );
  INV_X1 U3407 ( .A(n3964), .ZN(n5373) );
  AOI22_X1 U3408 ( .A1(\mem[156][7] ), .A2(n3957), .B1(n6712), .B2(data_in[7]), 
        .ZN(n3964) );
  INV_X1 U3409 ( .A(n3965), .ZN(n5372) );
  AOI22_X1 U3410 ( .A1(\mem[157][0] ), .A2(n3966), .B1(n6711), .B2(data_in[0]), 
        .ZN(n3965) );
  INV_X1 U3411 ( .A(n3967), .ZN(n5371) );
  AOI22_X1 U3412 ( .A1(\mem[157][1] ), .A2(n3966), .B1(n6711), .B2(data_in[1]), 
        .ZN(n3967) );
  INV_X1 U3413 ( .A(n3968), .ZN(n5370) );
  AOI22_X1 U3414 ( .A1(\mem[157][2] ), .A2(n3966), .B1(n6711), .B2(data_in[2]), 
        .ZN(n3968) );
  INV_X1 U3415 ( .A(n3969), .ZN(n5369) );
  AOI22_X1 U3416 ( .A1(\mem[157][3] ), .A2(n3966), .B1(n6711), .B2(data_in[3]), 
        .ZN(n3969) );
  INV_X1 U3417 ( .A(n3970), .ZN(n5368) );
  AOI22_X1 U3418 ( .A1(\mem[157][4] ), .A2(n3966), .B1(n6711), .B2(data_in[4]), 
        .ZN(n3970) );
  INV_X1 U3419 ( .A(n3971), .ZN(n5367) );
  AOI22_X1 U3420 ( .A1(\mem[157][5] ), .A2(n3966), .B1(n6711), .B2(data_in[5]), 
        .ZN(n3971) );
  INV_X1 U3421 ( .A(n3972), .ZN(n5366) );
  AOI22_X1 U3422 ( .A1(\mem[157][6] ), .A2(n3966), .B1(n6711), .B2(data_in[6]), 
        .ZN(n3972) );
  INV_X1 U3423 ( .A(n3973), .ZN(n5365) );
  AOI22_X1 U3424 ( .A1(\mem[157][7] ), .A2(n3966), .B1(n6711), .B2(data_in[7]), 
        .ZN(n3973) );
  INV_X1 U3425 ( .A(n3974), .ZN(n5364) );
  AOI22_X1 U3426 ( .A1(\mem[158][0] ), .A2(n3975), .B1(n6710), .B2(data_in[0]), 
        .ZN(n3974) );
  INV_X1 U3427 ( .A(n3976), .ZN(n5363) );
  AOI22_X1 U3428 ( .A1(\mem[158][1] ), .A2(n3975), .B1(n6710), .B2(data_in[1]), 
        .ZN(n3976) );
  INV_X1 U3429 ( .A(n3977), .ZN(n5362) );
  AOI22_X1 U3430 ( .A1(\mem[158][2] ), .A2(n3975), .B1(n6710), .B2(data_in[2]), 
        .ZN(n3977) );
  INV_X1 U3431 ( .A(n3978), .ZN(n5361) );
  AOI22_X1 U3432 ( .A1(\mem[158][3] ), .A2(n3975), .B1(n6710), .B2(data_in[3]), 
        .ZN(n3978) );
  INV_X1 U3433 ( .A(n3979), .ZN(n5360) );
  AOI22_X1 U3434 ( .A1(\mem[158][4] ), .A2(n3975), .B1(n6710), .B2(data_in[4]), 
        .ZN(n3979) );
  INV_X1 U3435 ( .A(n3980), .ZN(n5359) );
  AOI22_X1 U3436 ( .A1(\mem[158][5] ), .A2(n3975), .B1(n6710), .B2(data_in[5]), 
        .ZN(n3980) );
  INV_X1 U3437 ( .A(n3981), .ZN(n5358) );
  AOI22_X1 U3438 ( .A1(\mem[158][6] ), .A2(n3975), .B1(n6710), .B2(data_in[6]), 
        .ZN(n3981) );
  INV_X1 U3439 ( .A(n3982), .ZN(n5357) );
  AOI22_X1 U3440 ( .A1(\mem[158][7] ), .A2(n3975), .B1(n6710), .B2(data_in[7]), 
        .ZN(n3982) );
  INV_X1 U3441 ( .A(n3983), .ZN(n5356) );
  AOI22_X1 U3442 ( .A1(\mem[159][0] ), .A2(n3984), .B1(n6709), .B2(data_in[0]), 
        .ZN(n3983) );
  INV_X1 U3443 ( .A(n3985), .ZN(n5355) );
  AOI22_X1 U3444 ( .A1(\mem[159][1] ), .A2(n3984), .B1(n6709), .B2(data_in[1]), 
        .ZN(n3985) );
  INV_X1 U3445 ( .A(n3986), .ZN(n5354) );
  AOI22_X1 U3446 ( .A1(\mem[159][2] ), .A2(n3984), .B1(n6709), .B2(data_in[2]), 
        .ZN(n3986) );
  INV_X1 U3447 ( .A(n3987), .ZN(n5353) );
  AOI22_X1 U3448 ( .A1(\mem[159][3] ), .A2(n3984), .B1(n6709), .B2(data_in[3]), 
        .ZN(n3987) );
  INV_X1 U3449 ( .A(n3988), .ZN(n5352) );
  AOI22_X1 U3450 ( .A1(\mem[159][4] ), .A2(n3984), .B1(n6709), .B2(data_in[4]), 
        .ZN(n3988) );
  INV_X1 U3451 ( .A(n3989), .ZN(n5351) );
  AOI22_X1 U3452 ( .A1(\mem[159][5] ), .A2(n3984), .B1(n6709), .B2(data_in[5]), 
        .ZN(n3989) );
  INV_X1 U3453 ( .A(n3990), .ZN(n5350) );
  AOI22_X1 U3454 ( .A1(\mem[159][6] ), .A2(n3984), .B1(n6709), .B2(data_in[6]), 
        .ZN(n3990) );
  INV_X1 U3455 ( .A(n3991), .ZN(n5349) );
  AOI22_X1 U3456 ( .A1(\mem[159][7] ), .A2(n3984), .B1(n6709), .B2(data_in[7]), 
        .ZN(n3991) );
  INV_X1 U3457 ( .A(n3992), .ZN(n5348) );
  AOI22_X1 U3458 ( .A1(\mem[160][0] ), .A2(n3993), .B1(n6708), .B2(data_in[0]), 
        .ZN(n3992) );
  INV_X1 U3459 ( .A(n3994), .ZN(n5347) );
  AOI22_X1 U3460 ( .A1(\mem[160][1] ), .A2(n3993), .B1(n6708), .B2(data_in[1]), 
        .ZN(n3994) );
  INV_X1 U3461 ( .A(n3995), .ZN(n5346) );
  AOI22_X1 U3462 ( .A1(\mem[160][2] ), .A2(n3993), .B1(n6708), .B2(data_in[2]), 
        .ZN(n3995) );
  INV_X1 U3463 ( .A(n3996), .ZN(n5345) );
  AOI22_X1 U3464 ( .A1(\mem[160][3] ), .A2(n3993), .B1(n6708), .B2(data_in[3]), 
        .ZN(n3996) );
  INV_X1 U3465 ( .A(n3997), .ZN(n5344) );
  AOI22_X1 U3466 ( .A1(\mem[160][4] ), .A2(n3993), .B1(n6708), .B2(data_in[4]), 
        .ZN(n3997) );
  INV_X1 U3467 ( .A(n3998), .ZN(n5343) );
  AOI22_X1 U3468 ( .A1(\mem[160][5] ), .A2(n3993), .B1(n6708), .B2(data_in[5]), 
        .ZN(n3998) );
  INV_X1 U3469 ( .A(n3999), .ZN(n5342) );
  AOI22_X1 U3470 ( .A1(\mem[160][6] ), .A2(n3993), .B1(n6708), .B2(data_in[6]), 
        .ZN(n3999) );
  INV_X1 U3471 ( .A(n4000), .ZN(n5341) );
  AOI22_X1 U3472 ( .A1(\mem[160][7] ), .A2(n3993), .B1(n6708), .B2(data_in[7]), 
        .ZN(n4000) );
  INV_X1 U3473 ( .A(n4002), .ZN(n5340) );
  AOI22_X1 U3474 ( .A1(\mem[161][0] ), .A2(n4003), .B1(n6707), .B2(data_in[0]), 
        .ZN(n4002) );
  INV_X1 U3475 ( .A(n4004), .ZN(n5339) );
  AOI22_X1 U3476 ( .A1(\mem[161][1] ), .A2(n4003), .B1(n6707), .B2(data_in[1]), 
        .ZN(n4004) );
  INV_X1 U3477 ( .A(n4005), .ZN(n5338) );
  AOI22_X1 U3478 ( .A1(\mem[161][2] ), .A2(n4003), .B1(n6707), .B2(data_in[2]), 
        .ZN(n4005) );
  INV_X1 U3479 ( .A(n4006), .ZN(n5337) );
  AOI22_X1 U3480 ( .A1(\mem[161][3] ), .A2(n4003), .B1(n6707), .B2(data_in[3]), 
        .ZN(n4006) );
  INV_X1 U3481 ( .A(n4007), .ZN(n5336) );
  AOI22_X1 U3482 ( .A1(\mem[161][4] ), .A2(n4003), .B1(n6707), .B2(data_in[4]), 
        .ZN(n4007) );
  INV_X1 U3483 ( .A(n4008), .ZN(n5335) );
  AOI22_X1 U3484 ( .A1(\mem[161][5] ), .A2(n4003), .B1(n6707), .B2(data_in[5]), 
        .ZN(n4008) );
  INV_X1 U3485 ( .A(n4009), .ZN(n5334) );
  AOI22_X1 U3486 ( .A1(\mem[161][6] ), .A2(n4003), .B1(n6707), .B2(data_in[6]), 
        .ZN(n4009) );
  INV_X1 U3487 ( .A(n4010), .ZN(n5333) );
  AOI22_X1 U3488 ( .A1(\mem[161][7] ), .A2(n4003), .B1(n6707), .B2(data_in[7]), 
        .ZN(n4010) );
  INV_X1 U3489 ( .A(n4011), .ZN(n5332) );
  AOI22_X1 U3490 ( .A1(\mem[162][0] ), .A2(n4012), .B1(n6706), .B2(data_in[0]), 
        .ZN(n4011) );
  INV_X1 U3491 ( .A(n4013), .ZN(n5331) );
  AOI22_X1 U3492 ( .A1(\mem[162][1] ), .A2(n4012), .B1(n6706), .B2(data_in[1]), 
        .ZN(n4013) );
  INV_X1 U3493 ( .A(n4014), .ZN(n5330) );
  AOI22_X1 U3494 ( .A1(\mem[162][2] ), .A2(n4012), .B1(n6706), .B2(data_in[2]), 
        .ZN(n4014) );
  INV_X1 U3495 ( .A(n4015), .ZN(n5329) );
  AOI22_X1 U3496 ( .A1(\mem[162][3] ), .A2(n4012), .B1(n6706), .B2(data_in[3]), 
        .ZN(n4015) );
  INV_X1 U3497 ( .A(n4016), .ZN(n5328) );
  AOI22_X1 U3498 ( .A1(\mem[162][4] ), .A2(n4012), .B1(n6706), .B2(data_in[4]), 
        .ZN(n4016) );
  INV_X1 U3499 ( .A(n4017), .ZN(n5327) );
  AOI22_X1 U3500 ( .A1(\mem[162][5] ), .A2(n4012), .B1(n6706), .B2(data_in[5]), 
        .ZN(n4017) );
  INV_X1 U3501 ( .A(n4018), .ZN(n5326) );
  AOI22_X1 U3502 ( .A1(\mem[162][6] ), .A2(n4012), .B1(n6706), .B2(data_in[6]), 
        .ZN(n4018) );
  INV_X1 U3503 ( .A(n4019), .ZN(n5325) );
  AOI22_X1 U3504 ( .A1(\mem[162][7] ), .A2(n4012), .B1(n6706), .B2(data_in[7]), 
        .ZN(n4019) );
  INV_X1 U3505 ( .A(n4020), .ZN(n5324) );
  AOI22_X1 U3506 ( .A1(\mem[163][0] ), .A2(n4021), .B1(n6705), .B2(data_in[0]), 
        .ZN(n4020) );
  INV_X1 U3507 ( .A(n4022), .ZN(n5323) );
  AOI22_X1 U3508 ( .A1(\mem[163][1] ), .A2(n4021), .B1(n6705), .B2(data_in[1]), 
        .ZN(n4022) );
  INV_X1 U3509 ( .A(n4023), .ZN(n5322) );
  AOI22_X1 U3510 ( .A1(\mem[163][2] ), .A2(n4021), .B1(n6705), .B2(data_in[2]), 
        .ZN(n4023) );
  INV_X1 U3511 ( .A(n4024), .ZN(n5321) );
  AOI22_X1 U3512 ( .A1(\mem[163][3] ), .A2(n4021), .B1(n6705), .B2(data_in[3]), 
        .ZN(n4024) );
  INV_X1 U3513 ( .A(n4025), .ZN(n5320) );
  AOI22_X1 U3514 ( .A1(\mem[163][4] ), .A2(n4021), .B1(n6705), .B2(data_in[4]), 
        .ZN(n4025) );
  INV_X1 U3515 ( .A(n4026), .ZN(n5319) );
  AOI22_X1 U3516 ( .A1(\mem[163][5] ), .A2(n4021), .B1(n6705), .B2(data_in[5]), 
        .ZN(n4026) );
  INV_X1 U3517 ( .A(n4027), .ZN(n5318) );
  AOI22_X1 U3518 ( .A1(\mem[163][6] ), .A2(n4021), .B1(n6705), .B2(data_in[6]), 
        .ZN(n4027) );
  INV_X1 U3519 ( .A(n4028), .ZN(n5317) );
  AOI22_X1 U3520 ( .A1(\mem[163][7] ), .A2(n4021), .B1(n6705), .B2(data_in[7]), 
        .ZN(n4028) );
  INV_X1 U3521 ( .A(n4029), .ZN(n5316) );
  AOI22_X1 U3522 ( .A1(\mem[164][0] ), .A2(n4030), .B1(n6704), .B2(data_in[0]), 
        .ZN(n4029) );
  INV_X1 U3523 ( .A(n4031), .ZN(n5315) );
  AOI22_X1 U3524 ( .A1(\mem[164][1] ), .A2(n4030), .B1(n6704), .B2(data_in[1]), 
        .ZN(n4031) );
  INV_X1 U3525 ( .A(n4032), .ZN(n5314) );
  AOI22_X1 U3526 ( .A1(\mem[164][2] ), .A2(n4030), .B1(n6704), .B2(data_in[2]), 
        .ZN(n4032) );
  INV_X1 U3527 ( .A(n4033), .ZN(n5313) );
  AOI22_X1 U3528 ( .A1(\mem[164][3] ), .A2(n4030), .B1(n6704), .B2(data_in[3]), 
        .ZN(n4033) );
  INV_X1 U3529 ( .A(n4034), .ZN(n5312) );
  AOI22_X1 U3530 ( .A1(\mem[164][4] ), .A2(n4030), .B1(n6704), .B2(data_in[4]), 
        .ZN(n4034) );
  INV_X1 U3531 ( .A(n4035), .ZN(n5311) );
  AOI22_X1 U3532 ( .A1(\mem[164][5] ), .A2(n4030), .B1(n6704), .B2(data_in[5]), 
        .ZN(n4035) );
  INV_X1 U3533 ( .A(n4036), .ZN(n5310) );
  AOI22_X1 U3534 ( .A1(\mem[164][6] ), .A2(n4030), .B1(n6704), .B2(data_in[6]), 
        .ZN(n4036) );
  INV_X1 U3535 ( .A(n4037), .ZN(n5309) );
  AOI22_X1 U3536 ( .A1(\mem[164][7] ), .A2(n4030), .B1(n6704), .B2(data_in[7]), 
        .ZN(n4037) );
  INV_X1 U3537 ( .A(n4038), .ZN(n5308) );
  AOI22_X1 U3538 ( .A1(\mem[165][0] ), .A2(n4039), .B1(n6703), .B2(data_in[0]), 
        .ZN(n4038) );
  INV_X1 U3539 ( .A(n4040), .ZN(n5307) );
  AOI22_X1 U3540 ( .A1(\mem[165][1] ), .A2(n4039), .B1(n6703), .B2(data_in[1]), 
        .ZN(n4040) );
  INV_X1 U3541 ( .A(n4041), .ZN(n5306) );
  AOI22_X1 U3542 ( .A1(\mem[165][2] ), .A2(n4039), .B1(n6703), .B2(data_in[2]), 
        .ZN(n4041) );
  INV_X1 U3543 ( .A(n4042), .ZN(n5305) );
  AOI22_X1 U3544 ( .A1(\mem[165][3] ), .A2(n4039), .B1(n6703), .B2(data_in[3]), 
        .ZN(n4042) );
  INV_X1 U3545 ( .A(n4043), .ZN(n5304) );
  AOI22_X1 U3546 ( .A1(\mem[165][4] ), .A2(n4039), .B1(n6703), .B2(data_in[4]), 
        .ZN(n4043) );
  INV_X1 U3547 ( .A(n4044), .ZN(n5303) );
  AOI22_X1 U3548 ( .A1(\mem[165][5] ), .A2(n4039), .B1(n6703), .B2(data_in[5]), 
        .ZN(n4044) );
  INV_X1 U3549 ( .A(n4045), .ZN(n5302) );
  AOI22_X1 U3550 ( .A1(\mem[165][6] ), .A2(n4039), .B1(n6703), .B2(data_in[6]), 
        .ZN(n4045) );
  INV_X1 U3551 ( .A(n4046), .ZN(n5301) );
  AOI22_X1 U3552 ( .A1(\mem[165][7] ), .A2(n4039), .B1(n6703), .B2(data_in[7]), 
        .ZN(n4046) );
  INV_X1 U3553 ( .A(n4047), .ZN(n5300) );
  AOI22_X1 U3554 ( .A1(\mem[166][0] ), .A2(n4048), .B1(n6702), .B2(data_in[0]), 
        .ZN(n4047) );
  INV_X1 U3555 ( .A(n4049), .ZN(n5299) );
  AOI22_X1 U3556 ( .A1(\mem[166][1] ), .A2(n4048), .B1(n6702), .B2(data_in[1]), 
        .ZN(n4049) );
  INV_X1 U3557 ( .A(n4050), .ZN(n5298) );
  AOI22_X1 U3558 ( .A1(\mem[166][2] ), .A2(n4048), .B1(n6702), .B2(data_in[2]), 
        .ZN(n4050) );
  INV_X1 U3559 ( .A(n4051), .ZN(n5297) );
  AOI22_X1 U3560 ( .A1(\mem[166][3] ), .A2(n4048), .B1(n6702), .B2(data_in[3]), 
        .ZN(n4051) );
  INV_X1 U3561 ( .A(n4052), .ZN(n5296) );
  AOI22_X1 U3562 ( .A1(\mem[166][4] ), .A2(n4048), .B1(n6702), .B2(data_in[4]), 
        .ZN(n4052) );
  INV_X1 U3563 ( .A(n4053), .ZN(n5295) );
  AOI22_X1 U3564 ( .A1(\mem[166][5] ), .A2(n4048), .B1(n6702), .B2(data_in[5]), 
        .ZN(n4053) );
  INV_X1 U3565 ( .A(n4054), .ZN(n5294) );
  AOI22_X1 U3566 ( .A1(\mem[166][6] ), .A2(n4048), .B1(n6702), .B2(data_in[6]), 
        .ZN(n4054) );
  INV_X1 U3567 ( .A(n4055), .ZN(n5293) );
  AOI22_X1 U3568 ( .A1(\mem[166][7] ), .A2(n4048), .B1(n6702), .B2(data_in[7]), 
        .ZN(n4055) );
  INV_X1 U3569 ( .A(n4056), .ZN(n5292) );
  AOI22_X1 U3570 ( .A1(\mem[167][0] ), .A2(n4057), .B1(n6701), .B2(data_in[0]), 
        .ZN(n4056) );
  INV_X1 U3571 ( .A(n4058), .ZN(n5291) );
  AOI22_X1 U3572 ( .A1(\mem[167][1] ), .A2(n4057), .B1(n6701), .B2(data_in[1]), 
        .ZN(n4058) );
  INV_X1 U3573 ( .A(n4059), .ZN(n5290) );
  AOI22_X1 U3574 ( .A1(\mem[167][2] ), .A2(n4057), .B1(n6701), .B2(data_in[2]), 
        .ZN(n4059) );
  INV_X1 U3575 ( .A(n4060), .ZN(n5289) );
  AOI22_X1 U3576 ( .A1(\mem[167][3] ), .A2(n4057), .B1(n6701), .B2(data_in[3]), 
        .ZN(n4060) );
  INV_X1 U3577 ( .A(n4061), .ZN(n5288) );
  AOI22_X1 U3578 ( .A1(\mem[167][4] ), .A2(n4057), .B1(n6701), .B2(data_in[4]), 
        .ZN(n4061) );
  INV_X1 U3579 ( .A(n4062), .ZN(n5287) );
  AOI22_X1 U3580 ( .A1(\mem[167][5] ), .A2(n4057), .B1(n6701), .B2(data_in[5]), 
        .ZN(n4062) );
  INV_X1 U3581 ( .A(n4063), .ZN(n5286) );
  AOI22_X1 U3582 ( .A1(\mem[167][6] ), .A2(n4057), .B1(n6701), .B2(data_in[6]), 
        .ZN(n4063) );
  INV_X1 U3583 ( .A(n4064), .ZN(n5285) );
  AOI22_X1 U3584 ( .A1(\mem[167][7] ), .A2(n4057), .B1(n6701), .B2(data_in[7]), 
        .ZN(n4064) );
  INV_X1 U3585 ( .A(n4065), .ZN(n5284) );
  AOI22_X1 U3586 ( .A1(\mem[168][0] ), .A2(n4066), .B1(n6700), .B2(data_in[0]), 
        .ZN(n4065) );
  INV_X1 U3587 ( .A(n4067), .ZN(n5283) );
  AOI22_X1 U3588 ( .A1(\mem[168][1] ), .A2(n4066), .B1(n6700), .B2(data_in[1]), 
        .ZN(n4067) );
  INV_X1 U3589 ( .A(n4068), .ZN(n5282) );
  AOI22_X1 U3590 ( .A1(\mem[168][2] ), .A2(n4066), .B1(n6700), .B2(data_in[2]), 
        .ZN(n4068) );
  INV_X1 U3591 ( .A(n4069), .ZN(n5281) );
  AOI22_X1 U3592 ( .A1(\mem[168][3] ), .A2(n4066), .B1(n6700), .B2(data_in[3]), 
        .ZN(n4069) );
  INV_X1 U3593 ( .A(n4070), .ZN(n5280) );
  AOI22_X1 U3594 ( .A1(\mem[168][4] ), .A2(n4066), .B1(n6700), .B2(data_in[4]), 
        .ZN(n4070) );
  INV_X1 U3595 ( .A(n4071), .ZN(n5279) );
  AOI22_X1 U3596 ( .A1(\mem[168][5] ), .A2(n4066), .B1(n6700), .B2(data_in[5]), 
        .ZN(n4071) );
  INV_X1 U3597 ( .A(n4072), .ZN(n5278) );
  AOI22_X1 U3598 ( .A1(\mem[168][6] ), .A2(n4066), .B1(n6700), .B2(data_in[6]), 
        .ZN(n4072) );
  INV_X1 U3599 ( .A(n4073), .ZN(n5277) );
  AOI22_X1 U3600 ( .A1(\mem[168][7] ), .A2(n4066), .B1(n6700), .B2(data_in[7]), 
        .ZN(n4073) );
  INV_X1 U3601 ( .A(n4074), .ZN(n5276) );
  AOI22_X1 U3602 ( .A1(\mem[169][0] ), .A2(n4075), .B1(n6699), .B2(data_in[0]), 
        .ZN(n4074) );
  INV_X1 U3603 ( .A(n4076), .ZN(n5275) );
  AOI22_X1 U3604 ( .A1(\mem[169][1] ), .A2(n4075), .B1(n6699), .B2(data_in[1]), 
        .ZN(n4076) );
  INV_X1 U3605 ( .A(n4077), .ZN(n5274) );
  AOI22_X1 U3606 ( .A1(\mem[169][2] ), .A2(n4075), .B1(n6699), .B2(data_in[2]), 
        .ZN(n4077) );
  INV_X1 U3607 ( .A(n4078), .ZN(n5273) );
  AOI22_X1 U3608 ( .A1(\mem[169][3] ), .A2(n4075), .B1(n6699), .B2(data_in[3]), 
        .ZN(n4078) );
  INV_X1 U3609 ( .A(n4079), .ZN(n5272) );
  AOI22_X1 U3610 ( .A1(\mem[169][4] ), .A2(n4075), .B1(n6699), .B2(data_in[4]), 
        .ZN(n4079) );
  INV_X1 U3611 ( .A(n4080), .ZN(n5271) );
  AOI22_X1 U3612 ( .A1(\mem[169][5] ), .A2(n4075), .B1(n6699), .B2(data_in[5]), 
        .ZN(n4080) );
  INV_X1 U3613 ( .A(n4081), .ZN(n5270) );
  AOI22_X1 U3614 ( .A1(\mem[169][6] ), .A2(n4075), .B1(n6699), .B2(data_in[6]), 
        .ZN(n4081) );
  INV_X1 U3615 ( .A(n4082), .ZN(n5269) );
  AOI22_X1 U3616 ( .A1(\mem[169][7] ), .A2(n4075), .B1(n6699), .B2(data_in[7]), 
        .ZN(n4082) );
  INV_X1 U3617 ( .A(n4083), .ZN(n5268) );
  AOI22_X1 U3618 ( .A1(\mem[170][0] ), .A2(n4084), .B1(n6698), .B2(data_in[0]), 
        .ZN(n4083) );
  INV_X1 U3619 ( .A(n4085), .ZN(n5267) );
  AOI22_X1 U3620 ( .A1(\mem[170][1] ), .A2(n4084), .B1(n6698), .B2(data_in[1]), 
        .ZN(n4085) );
  INV_X1 U3621 ( .A(n4086), .ZN(n5266) );
  AOI22_X1 U3622 ( .A1(\mem[170][2] ), .A2(n4084), .B1(n6698), .B2(data_in[2]), 
        .ZN(n4086) );
  INV_X1 U3623 ( .A(n4087), .ZN(n5265) );
  AOI22_X1 U3624 ( .A1(\mem[170][3] ), .A2(n4084), .B1(n6698), .B2(data_in[3]), 
        .ZN(n4087) );
  INV_X1 U3625 ( .A(n4088), .ZN(n5264) );
  AOI22_X1 U3626 ( .A1(\mem[170][4] ), .A2(n4084), .B1(n6698), .B2(data_in[4]), 
        .ZN(n4088) );
  INV_X1 U3627 ( .A(n4089), .ZN(n5263) );
  AOI22_X1 U3628 ( .A1(\mem[170][5] ), .A2(n4084), .B1(n6698), .B2(data_in[5]), 
        .ZN(n4089) );
  INV_X1 U3629 ( .A(n4090), .ZN(n5262) );
  AOI22_X1 U3630 ( .A1(\mem[170][6] ), .A2(n4084), .B1(n6698), .B2(data_in[6]), 
        .ZN(n4090) );
  INV_X1 U3631 ( .A(n4091), .ZN(n5261) );
  AOI22_X1 U3632 ( .A1(\mem[170][7] ), .A2(n4084), .B1(n6698), .B2(data_in[7]), 
        .ZN(n4091) );
  INV_X1 U3633 ( .A(n4092), .ZN(n5260) );
  AOI22_X1 U3634 ( .A1(\mem[171][0] ), .A2(n4093), .B1(n6697), .B2(data_in[0]), 
        .ZN(n4092) );
  INV_X1 U3635 ( .A(n4094), .ZN(n5259) );
  AOI22_X1 U3636 ( .A1(\mem[171][1] ), .A2(n4093), .B1(n6697), .B2(data_in[1]), 
        .ZN(n4094) );
  INV_X1 U3637 ( .A(n4095), .ZN(n5258) );
  AOI22_X1 U3638 ( .A1(\mem[171][2] ), .A2(n4093), .B1(n6697), .B2(data_in[2]), 
        .ZN(n4095) );
  INV_X1 U3639 ( .A(n4096), .ZN(n5257) );
  AOI22_X1 U3640 ( .A1(\mem[171][3] ), .A2(n4093), .B1(n6697), .B2(data_in[3]), 
        .ZN(n4096) );
  INV_X1 U3641 ( .A(n4097), .ZN(n5256) );
  AOI22_X1 U3642 ( .A1(\mem[171][4] ), .A2(n4093), .B1(n6697), .B2(data_in[4]), 
        .ZN(n4097) );
  INV_X1 U3643 ( .A(n4098), .ZN(n5255) );
  AOI22_X1 U3644 ( .A1(\mem[171][5] ), .A2(n4093), .B1(n6697), .B2(data_in[5]), 
        .ZN(n4098) );
  INV_X1 U3645 ( .A(n4099), .ZN(n5254) );
  AOI22_X1 U3646 ( .A1(\mem[171][6] ), .A2(n4093), .B1(n6697), .B2(data_in[6]), 
        .ZN(n4099) );
  INV_X1 U3647 ( .A(n4100), .ZN(n5253) );
  AOI22_X1 U3648 ( .A1(\mem[171][7] ), .A2(n4093), .B1(n6697), .B2(data_in[7]), 
        .ZN(n4100) );
  INV_X1 U3649 ( .A(n4101), .ZN(n5252) );
  AOI22_X1 U3650 ( .A1(\mem[172][0] ), .A2(n4102), .B1(n6696), .B2(data_in[0]), 
        .ZN(n4101) );
  INV_X1 U3651 ( .A(n4103), .ZN(n5251) );
  AOI22_X1 U3652 ( .A1(\mem[172][1] ), .A2(n4102), .B1(n6696), .B2(data_in[1]), 
        .ZN(n4103) );
  INV_X1 U3653 ( .A(n4104), .ZN(n5250) );
  AOI22_X1 U3654 ( .A1(\mem[172][2] ), .A2(n4102), .B1(n6696), .B2(data_in[2]), 
        .ZN(n4104) );
  INV_X1 U3655 ( .A(n4105), .ZN(n5249) );
  AOI22_X1 U3656 ( .A1(\mem[172][3] ), .A2(n4102), .B1(n6696), .B2(data_in[3]), 
        .ZN(n4105) );
  INV_X1 U3657 ( .A(n4106), .ZN(n5248) );
  AOI22_X1 U3658 ( .A1(\mem[172][4] ), .A2(n4102), .B1(n6696), .B2(data_in[4]), 
        .ZN(n4106) );
  INV_X1 U3659 ( .A(n4107), .ZN(n5247) );
  AOI22_X1 U3660 ( .A1(\mem[172][5] ), .A2(n4102), .B1(n6696), .B2(data_in[5]), 
        .ZN(n4107) );
  INV_X1 U3661 ( .A(n4108), .ZN(n5246) );
  AOI22_X1 U3662 ( .A1(\mem[172][6] ), .A2(n4102), .B1(n6696), .B2(data_in[6]), 
        .ZN(n4108) );
  INV_X1 U3663 ( .A(n4109), .ZN(n5245) );
  AOI22_X1 U3664 ( .A1(\mem[172][7] ), .A2(n4102), .B1(n6696), .B2(data_in[7]), 
        .ZN(n4109) );
  INV_X1 U3665 ( .A(n4110), .ZN(n5244) );
  AOI22_X1 U3666 ( .A1(\mem[173][0] ), .A2(n4111), .B1(n6695), .B2(data_in[0]), 
        .ZN(n4110) );
  INV_X1 U3667 ( .A(n4112), .ZN(n5243) );
  AOI22_X1 U3668 ( .A1(\mem[173][1] ), .A2(n4111), .B1(n6695), .B2(data_in[1]), 
        .ZN(n4112) );
  INV_X1 U3669 ( .A(n4113), .ZN(n5242) );
  AOI22_X1 U3670 ( .A1(\mem[173][2] ), .A2(n4111), .B1(n6695), .B2(data_in[2]), 
        .ZN(n4113) );
  INV_X1 U3671 ( .A(n4114), .ZN(n5241) );
  AOI22_X1 U3672 ( .A1(\mem[173][3] ), .A2(n4111), .B1(n6695), .B2(data_in[3]), 
        .ZN(n4114) );
  INV_X1 U3673 ( .A(n4115), .ZN(n5240) );
  AOI22_X1 U3674 ( .A1(\mem[173][4] ), .A2(n4111), .B1(n6695), .B2(data_in[4]), 
        .ZN(n4115) );
  INV_X1 U3675 ( .A(n4116), .ZN(n5239) );
  AOI22_X1 U3676 ( .A1(\mem[173][5] ), .A2(n4111), .B1(n6695), .B2(data_in[5]), 
        .ZN(n4116) );
  INV_X1 U3677 ( .A(n4117), .ZN(n5238) );
  AOI22_X1 U3678 ( .A1(\mem[173][6] ), .A2(n4111), .B1(n6695), .B2(data_in[6]), 
        .ZN(n4117) );
  INV_X1 U3679 ( .A(n4118), .ZN(n5237) );
  AOI22_X1 U3680 ( .A1(\mem[173][7] ), .A2(n4111), .B1(n6695), .B2(data_in[7]), 
        .ZN(n4118) );
  INV_X1 U3681 ( .A(n4119), .ZN(n5236) );
  AOI22_X1 U3682 ( .A1(\mem[174][0] ), .A2(n4120), .B1(n6694), .B2(data_in[0]), 
        .ZN(n4119) );
  INV_X1 U3683 ( .A(n4121), .ZN(n5235) );
  AOI22_X1 U3684 ( .A1(\mem[174][1] ), .A2(n4120), .B1(n6694), .B2(data_in[1]), 
        .ZN(n4121) );
  INV_X1 U3685 ( .A(n4122), .ZN(n5234) );
  AOI22_X1 U3686 ( .A1(\mem[174][2] ), .A2(n4120), .B1(n6694), .B2(data_in[2]), 
        .ZN(n4122) );
  INV_X1 U3687 ( .A(n4123), .ZN(n5233) );
  AOI22_X1 U3688 ( .A1(\mem[174][3] ), .A2(n4120), .B1(n6694), .B2(data_in[3]), 
        .ZN(n4123) );
  INV_X1 U3689 ( .A(n4124), .ZN(n5232) );
  AOI22_X1 U3690 ( .A1(\mem[174][4] ), .A2(n4120), .B1(n6694), .B2(data_in[4]), 
        .ZN(n4124) );
  INV_X1 U3691 ( .A(n4125), .ZN(n5231) );
  AOI22_X1 U3692 ( .A1(\mem[174][5] ), .A2(n4120), .B1(n6694), .B2(data_in[5]), 
        .ZN(n4125) );
  INV_X1 U3693 ( .A(n4126), .ZN(n5230) );
  AOI22_X1 U3694 ( .A1(\mem[174][6] ), .A2(n4120), .B1(n6694), .B2(data_in[6]), 
        .ZN(n4126) );
  INV_X1 U3695 ( .A(n4127), .ZN(n5229) );
  AOI22_X1 U3696 ( .A1(\mem[174][7] ), .A2(n4120), .B1(n6694), .B2(data_in[7]), 
        .ZN(n4127) );
  INV_X1 U3697 ( .A(n4128), .ZN(n5228) );
  AOI22_X1 U3698 ( .A1(\mem[175][0] ), .A2(n4129), .B1(n6693), .B2(data_in[0]), 
        .ZN(n4128) );
  INV_X1 U3699 ( .A(n4130), .ZN(n5227) );
  AOI22_X1 U3700 ( .A1(\mem[175][1] ), .A2(n4129), .B1(n6693), .B2(data_in[1]), 
        .ZN(n4130) );
  INV_X1 U3701 ( .A(n4131), .ZN(n5226) );
  AOI22_X1 U3702 ( .A1(\mem[175][2] ), .A2(n4129), .B1(n6693), .B2(data_in[2]), 
        .ZN(n4131) );
  INV_X1 U3703 ( .A(n4132), .ZN(n5225) );
  AOI22_X1 U3704 ( .A1(\mem[175][3] ), .A2(n4129), .B1(n6693), .B2(data_in[3]), 
        .ZN(n4132) );
  INV_X1 U3705 ( .A(n4133), .ZN(n5224) );
  AOI22_X1 U3706 ( .A1(\mem[175][4] ), .A2(n4129), .B1(n6693), .B2(data_in[4]), 
        .ZN(n4133) );
  INV_X1 U3707 ( .A(n4134), .ZN(n5223) );
  AOI22_X1 U3708 ( .A1(\mem[175][5] ), .A2(n4129), .B1(n6693), .B2(data_in[5]), 
        .ZN(n4134) );
  INV_X1 U3709 ( .A(n4135), .ZN(n5222) );
  AOI22_X1 U3710 ( .A1(\mem[175][6] ), .A2(n4129), .B1(n6693), .B2(data_in[6]), 
        .ZN(n4135) );
  INV_X1 U3711 ( .A(n4136), .ZN(n5221) );
  AOI22_X1 U3712 ( .A1(\mem[175][7] ), .A2(n4129), .B1(n6693), .B2(data_in[7]), 
        .ZN(n4136) );
  INV_X1 U3713 ( .A(n4137), .ZN(n5220) );
  AOI22_X1 U3714 ( .A1(\mem[176][0] ), .A2(n4138), .B1(n6692), .B2(data_in[0]), 
        .ZN(n4137) );
  INV_X1 U3715 ( .A(n4139), .ZN(n5219) );
  AOI22_X1 U3716 ( .A1(\mem[176][1] ), .A2(n4138), .B1(n6692), .B2(data_in[1]), 
        .ZN(n4139) );
  INV_X1 U3717 ( .A(n4140), .ZN(n5218) );
  AOI22_X1 U3718 ( .A1(\mem[176][2] ), .A2(n4138), .B1(n6692), .B2(data_in[2]), 
        .ZN(n4140) );
  INV_X1 U3719 ( .A(n4141), .ZN(n5217) );
  AOI22_X1 U3720 ( .A1(\mem[176][3] ), .A2(n4138), .B1(n6692), .B2(data_in[3]), 
        .ZN(n4141) );
  INV_X1 U3721 ( .A(n4142), .ZN(n5216) );
  AOI22_X1 U3722 ( .A1(\mem[176][4] ), .A2(n4138), .B1(n6692), .B2(data_in[4]), 
        .ZN(n4142) );
  INV_X1 U3723 ( .A(n4143), .ZN(n5215) );
  AOI22_X1 U3724 ( .A1(\mem[176][5] ), .A2(n4138), .B1(n6692), .B2(data_in[5]), 
        .ZN(n4143) );
  INV_X1 U3725 ( .A(n4144), .ZN(n5214) );
  AOI22_X1 U3726 ( .A1(\mem[176][6] ), .A2(n4138), .B1(n6692), .B2(data_in[6]), 
        .ZN(n4144) );
  INV_X1 U3727 ( .A(n4145), .ZN(n5213) );
  AOI22_X1 U3728 ( .A1(\mem[176][7] ), .A2(n4138), .B1(n6692), .B2(data_in[7]), 
        .ZN(n4145) );
  INV_X1 U3729 ( .A(n4147), .ZN(n5212) );
  AOI22_X1 U3730 ( .A1(\mem[177][0] ), .A2(n4148), .B1(n6691), .B2(data_in[0]), 
        .ZN(n4147) );
  INV_X1 U3731 ( .A(n4149), .ZN(n5211) );
  AOI22_X1 U3732 ( .A1(\mem[177][1] ), .A2(n4148), .B1(n6691), .B2(data_in[1]), 
        .ZN(n4149) );
  INV_X1 U3733 ( .A(n4150), .ZN(n5210) );
  AOI22_X1 U3734 ( .A1(\mem[177][2] ), .A2(n4148), .B1(n6691), .B2(data_in[2]), 
        .ZN(n4150) );
  INV_X1 U3735 ( .A(n4151), .ZN(n5209) );
  AOI22_X1 U3736 ( .A1(\mem[177][3] ), .A2(n4148), .B1(n6691), .B2(data_in[3]), 
        .ZN(n4151) );
  INV_X1 U3737 ( .A(n4152), .ZN(n5208) );
  AOI22_X1 U3738 ( .A1(\mem[177][4] ), .A2(n4148), .B1(n6691), .B2(data_in[4]), 
        .ZN(n4152) );
  INV_X1 U3739 ( .A(n4153), .ZN(n5207) );
  AOI22_X1 U3740 ( .A1(\mem[177][5] ), .A2(n4148), .B1(n6691), .B2(data_in[5]), 
        .ZN(n4153) );
  INV_X1 U3741 ( .A(n4154), .ZN(n5206) );
  AOI22_X1 U3742 ( .A1(\mem[177][6] ), .A2(n4148), .B1(n6691), .B2(data_in[6]), 
        .ZN(n4154) );
  INV_X1 U3743 ( .A(n4155), .ZN(n5205) );
  AOI22_X1 U3744 ( .A1(\mem[177][7] ), .A2(n4148), .B1(n6691), .B2(data_in[7]), 
        .ZN(n4155) );
  INV_X1 U3745 ( .A(n4156), .ZN(n5204) );
  AOI22_X1 U3746 ( .A1(\mem[178][0] ), .A2(n4157), .B1(n6690), .B2(data_in[0]), 
        .ZN(n4156) );
  INV_X1 U3747 ( .A(n4158), .ZN(n5203) );
  AOI22_X1 U3748 ( .A1(\mem[178][1] ), .A2(n4157), .B1(n6690), .B2(data_in[1]), 
        .ZN(n4158) );
  INV_X1 U3749 ( .A(n4159), .ZN(n5202) );
  AOI22_X1 U3750 ( .A1(\mem[178][2] ), .A2(n4157), .B1(n6690), .B2(data_in[2]), 
        .ZN(n4159) );
  INV_X1 U3751 ( .A(n4160), .ZN(n5201) );
  AOI22_X1 U3752 ( .A1(\mem[178][3] ), .A2(n4157), .B1(n6690), .B2(data_in[3]), 
        .ZN(n4160) );
  INV_X1 U3753 ( .A(n4161), .ZN(n5200) );
  AOI22_X1 U3754 ( .A1(\mem[178][4] ), .A2(n4157), .B1(n6690), .B2(data_in[4]), 
        .ZN(n4161) );
  INV_X1 U3755 ( .A(n4162), .ZN(n5199) );
  AOI22_X1 U3756 ( .A1(\mem[178][5] ), .A2(n4157), .B1(n6690), .B2(data_in[5]), 
        .ZN(n4162) );
  INV_X1 U3757 ( .A(n4163), .ZN(n5198) );
  AOI22_X1 U3758 ( .A1(\mem[178][6] ), .A2(n4157), .B1(n6690), .B2(data_in[6]), 
        .ZN(n4163) );
  INV_X1 U3759 ( .A(n4164), .ZN(n5197) );
  AOI22_X1 U3760 ( .A1(\mem[178][7] ), .A2(n4157), .B1(n6690), .B2(data_in[7]), 
        .ZN(n4164) );
  INV_X1 U3761 ( .A(n4165), .ZN(n5196) );
  AOI22_X1 U3762 ( .A1(\mem[179][0] ), .A2(n4166), .B1(n6689), .B2(data_in[0]), 
        .ZN(n4165) );
  INV_X1 U3763 ( .A(n4167), .ZN(n5195) );
  AOI22_X1 U3764 ( .A1(\mem[179][1] ), .A2(n4166), .B1(n6689), .B2(data_in[1]), 
        .ZN(n4167) );
  INV_X1 U3765 ( .A(n4168), .ZN(n5194) );
  AOI22_X1 U3766 ( .A1(\mem[179][2] ), .A2(n4166), .B1(n6689), .B2(data_in[2]), 
        .ZN(n4168) );
  INV_X1 U3767 ( .A(n4169), .ZN(n5193) );
  AOI22_X1 U3768 ( .A1(\mem[179][3] ), .A2(n4166), .B1(n6689), .B2(data_in[3]), 
        .ZN(n4169) );
  INV_X1 U3769 ( .A(n4170), .ZN(n5192) );
  AOI22_X1 U3770 ( .A1(\mem[179][4] ), .A2(n4166), .B1(n6689), .B2(data_in[4]), 
        .ZN(n4170) );
  INV_X1 U3771 ( .A(n4171), .ZN(n5191) );
  AOI22_X1 U3772 ( .A1(\mem[179][5] ), .A2(n4166), .B1(n6689), .B2(data_in[5]), 
        .ZN(n4171) );
  INV_X1 U3773 ( .A(n4172), .ZN(n5190) );
  AOI22_X1 U3774 ( .A1(\mem[179][6] ), .A2(n4166), .B1(n6689), .B2(data_in[6]), 
        .ZN(n4172) );
  INV_X1 U3775 ( .A(n4173), .ZN(n5189) );
  AOI22_X1 U3776 ( .A1(\mem[179][7] ), .A2(n4166), .B1(n6689), .B2(data_in[7]), 
        .ZN(n4173) );
  INV_X1 U3777 ( .A(n4174), .ZN(n5188) );
  AOI22_X1 U3778 ( .A1(\mem[180][0] ), .A2(n4175), .B1(n6688), .B2(data_in[0]), 
        .ZN(n4174) );
  INV_X1 U3779 ( .A(n4176), .ZN(n5187) );
  AOI22_X1 U3780 ( .A1(\mem[180][1] ), .A2(n4175), .B1(n6688), .B2(data_in[1]), 
        .ZN(n4176) );
  INV_X1 U3781 ( .A(n4177), .ZN(n5186) );
  AOI22_X1 U3782 ( .A1(\mem[180][2] ), .A2(n4175), .B1(n6688), .B2(data_in[2]), 
        .ZN(n4177) );
  INV_X1 U3783 ( .A(n4178), .ZN(n5185) );
  AOI22_X1 U3784 ( .A1(\mem[180][3] ), .A2(n4175), .B1(n6688), .B2(data_in[3]), 
        .ZN(n4178) );
  INV_X1 U3785 ( .A(n4179), .ZN(n5184) );
  AOI22_X1 U3786 ( .A1(\mem[180][4] ), .A2(n4175), .B1(n6688), .B2(data_in[4]), 
        .ZN(n4179) );
  INV_X1 U3787 ( .A(n4180), .ZN(n5183) );
  AOI22_X1 U3788 ( .A1(\mem[180][5] ), .A2(n4175), .B1(n6688), .B2(data_in[5]), 
        .ZN(n4180) );
  INV_X1 U3789 ( .A(n4181), .ZN(n5182) );
  AOI22_X1 U3790 ( .A1(\mem[180][6] ), .A2(n4175), .B1(n6688), .B2(data_in[6]), 
        .ZN(n4181) );
  INV_X1 U3791 ( .A(n4182), .ZN(n5181) );
  AOI22_X1 U3792 ( .A1(\mem[180][7] ), .A2(n4175), .B1(n6688), .B2(data_in[7]), 
        .ZN(n4182) );
  INV_X1 U3793 ( .A(n4183), .ZN(n5180) );
  AOI22_X1 U3794 ( .A1(\mem[181][0] ), .A2(n4184), .B1(n6687), .B2(data_in[0]), 
        .ZN(n4183) );
  INV_X1 U3795 ( .A(n4185), .ZN(n5179) );
  AOI22_X1 U3796 ( .A1(\mem[181][1] ), .A2(n4184), .B1(n6687), .B2(data_in[1]), 
        .ZN(n4185) );
  INV_X1 U3797 ( .A(n4186), .ZN(n5178) );
  AOI22_X1 U3798 ( .A1(\mem[181][2] ), .A2(n4184), .B1(n6687), .B2(data_in[2]), 
        .ZN(n4186) );
  INV_X1 U3799 ( .A(n4187), .ZN(n5177) );
  AOI22_X1 U3800 ( .A1(\mem[181][3] ), .A2(n4184), .B1(n6687), .B2(data_in[3]), 
        .ZN(n4187) );
  INV_X1 U3801 ( .A(n4188), .ZN(n5176) );
  AOI22_X1 U3802 ( .A1(\mem[181][4] ), .A2(n4184), .B1(n6687), .B2(data_in[4]), 
        .ZN(n4188) );
  INV_X1 U3803 ( .A(n4189), .ZN(n5175) );
  AOI22_X1 U3804 ( .A1(\mem[181][5] ), .A2(n4184), .B1(n6687), .B2(data_in[5]), 
        .ZN(n4189) );
  INV_X1 U3805 ( .A(n4190), .ZN(n5174) );
  AOI22_X1 U3806 ( .A1(\mem[181][6] ), .A2(n4184), .B1(n6687), .B2(data_in[6]), 
        .ZN(n4190) );
  INV_X1 U3807 ( .A(n4191), .ZN(n5173) );
  AOI22_X1 U3808 ( .A1(\mem[181][7] ), .A2(n4184), .B1(n6687), .B2(data_in[7]), 
        .ZN(n4191) );
  INV_X1 U3809 ( .A(n4192), .ZN(n5172) );
  AOI22_X1 U3810 ( .A1(\mem[182][0] ), .A2(n4193), .B1(n6686), .B2(data_in[0]), 
        .ZN(n4192) );
  INV_X1 U3811 ( .A(n4194), .ZN(n5171) );
  AOI22_X1 U3812 ( .A1(\mem[182][1] ), .A2(n4193), .B1(n6686), .B2(data_in[1]), 
        .ZN(n4194) );
  INV_X1 U3813 ( .A(n4195), .ZN(n5170) );
  AOI22_X1 U3814 ( .A1(\mem[182][2] ), .A2(n4193), .B1(n6686), .B2(data_in[2]), 
        .ZN(n4195) );
  INV_X1 U3815 ( .A(n4196), .ZN(n5169) );
  AOI22_X1 U3816 ( .A1(\mem[182][3] ), .A2(n4193), .B1(n6686), .B2(data_in[3]), 
        .ZN(n4196) );
  INV_X1 U3817 ( .A(n4197), .ZN(n5168) );
  AOI22_X1 U3818 ( .A1(\mem[182][4] ), .A2(n4193), .B1(n6686), .B2(data_in[4]), 
        .ZN(n4197) );
  INV_X1 U3819 ( .A(n4198), .ZN(n5167) );
  AOI22_X1 U3820 ( .A1(\mem[182][5] ), .A2(n4193), .B1(n6686), .B2(data_in[5]), 
        .ZN(n4198) );
  INV_X1 U3821 ( .A(n4199), .ZN(n5166) );
  AOI22_X1 U3822 ( .A1(\mem[182][6] ), .A2(n4193), .B1(n6686), .B2(data_in[6]), 
        .ZN(n4199) );
  INV_X1 U3823 ( .A(n4200), .ZN(n5165) );
  AOI22_X1 U3824 ( .A1(\mem[182][7] ), .A2(n4193), .B1(n6686), .B2(data_in[7]), 
        .ZN(n4200) );
  INV_X1 U3825 ( .A(n4201), .ZN(n5164) );
  AOI22_X1 U3826 ( .A1(\mem[183][0] ), .A2(n4202), .B1(n6685), .B2(data_in[0]), 
        .ZN(n4201) );
  INV_X1 U3827 ( .A(n4203), .ZN(n5163) );
  AOI22_X1 U3828 ( .A1(\mem[183][1] ), .A2(n4202), .B1(n6685), .B2(data_in[1]), 
        .ZN(n4203) );
  INV_X1 U3829 ( .A(n4204), .ZN(n5162) );
  AOI22_X1 U3830 ( .A1(\mem[183][2] ), .A2(n4202), .B1(n6685), .B2(data_in[2]), 
        .ZN(n4204) );
  INV_X1 U3831 ( .A(n4205), .ZN(n5161) );
  AOI22_X1 U3832 ( .A1(\mem[183][3] ), .A2(n4202), .B1(n6685), .B2(data_in[3]), 
        .ZN(n4205) );
  INV_X1 U3833 ( .A(n4206), .ZN(n5160) );
  AOI22_X1 U3834 ( .A1(\mem[183][4] ), .A2(n4202), .B1(n6685), .B2(data_in[4]), 
        .ZN(n4206) );
  INV_X1 U3835 ( .A(n4207), .ZN(n5159) );
  AOI22_X1 U3836 ( .A1(\mem[183][5] ), .A2(n4202), .B1(n6685), .B2(data_in[5]), 
        .ZN(n4207) );
  INV_X1 U3837 ( .A(n4208), .ZN(n5158) );
  AOI22_X1 U3838 ( .A1(\mem[183][6] ), .A2(n4202), .B1(n6685), .B2(data_in[6]), 
        .ZN(n4208) );
  INV_X1 U3839 ( .A(n4209), .ZN(n5157) );
  AOI22_X1 U3840 ( .A1(\mem[183][7] ), .A2(n4202), .B1(n6685), .B2(data_in[7]), 
        .ZN(n4209) );
  INV_X1 U3841 ( .A(n4210), .ZN(n5156) );
  AOI22_X1 U3842 ( .A1(\mem[184][0] ), .A2(n4211), .B1(n6684), .B2(data_in[0]), 
        .ZN(n4210) );
  INV_X1 U3843 ( .A(n4212), .ZN(n5155) );
  AOI22_X1 U3844 ( .A1(\mem[184][1] ), .A2(n4211), .B1(n6684), .B2(data_in[1]), 
        .ZN(n4212) );
  INV_X1 U3845 ( .A(n4213), .ZN(n5154) );
  AOI22_X1 U3846 ( .A1(\mem[184][2] ), .A2(n4211), .B1(n6684), .B2(data_in[2]), 
        .ZN(n4213) );
  INV_X1 U3847 ( .A(n4214), .ZN(n5153) );
  AOI22_X1 U3848 ( .A1(\mem[184][3] ), .A2(n4211), .B1(n6684), .B2(data_in[3]), 
        .ZN(n4214) );
  INV_X1 U3849 ( .A(n4215), .ZN(n5152) );
  AOI22_X1 U3850 ( .A1(\mem[184][4] ), .A2(n4211), .B1(n6684), .B2(data_in[4]), 
        .ZN(n4215) );
  INV_X1 U3851 ( .A(n4216), .ZN(n5151) );
  AOI22_X1 U3852 ( .A1(\mem[184][5] ), .A2(n4211), .B1(n6684), .B2(data_in[5]), 
        .ZN(n4216) );
  INV_X1 U3853 ( .A(n4217), .ZN(n5150) );
  AOI22_X1 U3854 ( .A1(\mem[184][6] ), .A2(n4211), .B1(n6684), .B2(data_in[6]), 
        .ZN(n4217) );
  INV_X1 U3855 ( .A(n4218), .ZN(n5149) );
  AOI22_X1 U3856 ( .A1(\mem[184][7] ), .A2(n4211), .B1(n6684), .B2(data_in[7]), 
        .ZN(n4218) );
  INV_X1 U3857 ( .A(n4219), .ZN(n5148) );
  AOI22_X1 U3858 ( .A1(\mem[185][0] ), .A2(n4220), .B1(n6683), .B2(data_in[0]), 
        .ZN(n4219) );
  INV_X1 U3859 ( .A(n4221), .ZN(n5147) );
  AOI22_X1 U3860 ( .A1(\mem[185][1] ), .A2(n4220), .B1(n6683), .B2(data_in[1]), 
        .ZN(n4221) );
  INV_X1 U3861 ( .A(n4222), .ZN(n5146) );
  AOI22_X1 U3862 ( .A1(\mem[185][2] ), .A2(n4220), .B1(n6683), .B2(data_in[2]), 
        .ZN(n4222) );
  INV_X1 U3863 ( .A(n4223), .ZN(n5145) );
  AOI22_X1 U3864 ( .A1(\mem[185][3] ), .A2(n4220), .B1(n6683), .B2(data_in[3]), 
        .ZN(n4223) );
  INV_X1 U3865 ( .A(n4224), .ZN(n5144) );
  AOI22_X1 U3866 ( .A1(\mem[185][4] ), .A2(n4220), .B1(n6683), .B2(data_in[4]), 
        .ZN(n4224) );
  INV_X1 U3867 ( .A(n4225), .ZN(n5143) );
  AOI22_X1 U3868 ( .A1(\mem[185][5] ), .A2(n4220), .B1(n6683), .B2(data_in[5]), 
        .ZN(n4225) );
  INV_X1 U3869 ( .A(n4226), .ZN(n5142) );
  AOI22_X1 U3870 ( .A1(\mem[185][6] ), .A2(n4220), .B1(n6683), .B2(data_in[6]), 
        .ZN(n4226) );
  INV_X1 U3871 ( .A(n4227), .ZN(n5141) );
  AOI22_X1 U3872 ( .A1(\mem[185][7] ), .A2(n4220), .B1(n6683), .B2(data_in[7]), 
        .ZN(n4227) );
  INV_X1 U3873 ( .A(n4228), .ZN(n5140) );
  AOI22_X1 U3874 ( .A1(\mem[186][0] ), .A2(n4229), .B1(n6682), .B2(data_in[0]), 
        .ZN(n4228) );
  INV_X1 U3875 ( .A(n4230), .ZN(n5139) );
  AOI22_X1 U3876 ( .A1(\mem[186][1] ), .A2(n4229), .B1(n6682), .B2(data_in[1]), 
        .ZN(n4230) );
  INV_X1 U3877 ( .A(n4231), .ZN(n5138) );
  AOI22_X1 U3878 ( .A1(\mem[186][2] ), .A2(n4229), .B1(n6682), .B2(data_in[2]), 
        .ZN(n4231) );
  INV_X1 U3879 ( .A(n4232), .ZN(n5137) );
  AOI22_X1 U3880 ( .A1(\mem[186][3] ), .A2(n4229), .B1(n6682), .B2(data_in[3]), 
        .ZN(n4232) );
  INV_X1 U3881 ( .A(n4233), .ZN(n5136) );
  AOI22_X1 U3882 ( .A1(\mem[186][4] ), .A2(n4229), .B1(n6682), .B2(data_in[4]), 
        .ZN(n4233) );
  INV_X1 U3883 ( .A(n4234), .ZN(n5135) );
  AOI22_X1 U3884 ( .A1(\mem[186][5] ), .A2(n4229), .B1(n6682), .B2(data_in[5]), 
        .ZN(n4234) );
  INV_X1 U3885 ( .A(n4235), .ZN(n5134) );
  AOI22_X1 U3886 ( .A1(\mem[186][6] ), .A2(n4229), .B1(n6682), .B2(data_in[6]), 
        .ZN(n4235) );
  INV_X1 U3887 ( .A(n4236), .ZN(n5133) );
  AOI22_X1 U3888 ( .A1(\mem[186][7] ), .A2(n4229), .B1(n6682), .B2(data_in[7]), 
        .ZN(n4236) );
  INV_X1 U3889 ( .A(n4237), .ZN(n5132) );
  AOI22_X1 U3890 ( .A1(\mem[187][0] ), .A2(n4238), .B1(n6681), .B2(data_in[0]), 
        .ZN(n4237) );
  INV_X1 U3891 ( .A(n4239), .ZN(n5131) );
  AOI22_X1 U3892 ( .A1(\mem[187][1] ), .A2(n4238), .B1(n6681), .B2(data_in[1]), 
        .ZN(n4239) );
  INV_X1 U3893 ( .A(n4240), .ZN(n5130) );
  AOI22_X1 U3894 ( .A1(\mem[187][2] ), .A2(n4238), .B1(n6681), .B2(data_in[2]), 
        .ZN(n4240) );
  INV_X1 U3895 ( .A(n4241), .ZN(n5129) );
  AOI22_X1 U3896 ( .A1(\mem[187][3] ), .A2(n4238), .B1(n6681), .B2(data_in[3]), 
        .ZN(n4241) );
  INV_X1 U3897 ( .A(n4242), .ZN(n5128) );
  AOI22_X1 U3898 ( .A1(\mem[187][4] ), .A2(n4238), .B1(n6681), .B2(data_in[4]), 
        .ZN(n4242) );
  INV_X1 U3899 ( .A(n4243), .ZN(n5127) );
  AOI22_X1 U3900 ( .A1(\mem[187][5] ), .A2(n4238), .B1(n6681), .B2(data_in[5]), 
        .ZN(n4243) );
  INV_X1 U3901 ( .A(n4244), .ZN(n5126) );
  AOI22_X1 U3902 ( .A1(\mem[187][6] ), .A2(n4238), .B1(n6681), .B2(data_in[6]), 
        .ZN(n4244) );
  INV_X1 U3903 ( .A(n4245), .ZN(n5125) );
  AOI22_X1 U3904 ( .A1(\mem[187][7] ), .A2(n4238), .B1(n6681), .B2(data_in[7]), 
        .ZN(n4245) );
  INV_X1 U3905 ( .A(n4246), .ZN(n5124) );
  AOI22_X1 U3906 ( .A1(\mem[188][0] ), .A2(n4247), .B1(n6680), .B2(data_in[0]), 
        .ZN(n4246) );
  INV_X1 U3907 ( .A(n4248), .ZN(n5123) );
  AOI22_X1 U3908 ( .A1(\mem[188][1] ), .A2(n4247), .B1(n6680), .B2(data_in[1]), 
        .ZN(n4248) );
  INV_X1 U3909 ( .A(n4249), .ZN(n5122) );
  AOI22_X1 U3910 ( .A1(\mem[188][2] ), .A2(n4247), .B1(n6680), .B2(data_in[2]), 
        .ZN(n4249) );
  INV_X1 U3911 ( .A(n4250), .ZN(n5121) );
  AOI22_X1 U3912 ( .A1(\mem[188][3] ), .A2(n4247), .B1(n6680), .B2(data_in[3]), 
        .ZN(n4250) );
  INV_X1 U3913 ( .A(n4251), .ZN(n5120) );
  AOI22_X1 U3914 ( .A1(\mem[188][4] ), .A2(n4247), .B1(n6680), .B2(data_in[4]), 
        .ZN(n4251) );
  INV_X1 U3915 ( .A(n4252), .ZN(n5119) );
  AOI22_X1 U3916 ( .A1(\mem[188][5] ), .A2(n4247), .B1(n6680), .B2(data_in[5]), 
        .ZN(n4252) );
  INV_X1 U3917 ( .A(n4253), .ZN(n5118) );
  AOI22_X1 U3918 ( .A1(\mem[188][6] ), .A2(n4247), .B1(n6680), .B2(data_in[6]), 
        .ZN(n4253) );
  INV_X1 U3919 ( .A(n4254), .ZN(n5117) );
  AOI22_X1 U3920 ( .A1(\mem[188][7] ), .A2(n4247), .B1(n6680), .B2(data_in[7]), 
        .ZN(n4254) );
  INV_X1 U3921 ( .A(n4255), .ZN(n5116) );
  AOI22_X1 U3922 ( .A1(\mem[189][0] ), .A2(n4256), .B1(n6679), .B2(data_in[0]), 
        .ZN(n4255) );
  INV_X1 U3923 ( .A(n4257), .ZN(n5115) );
  AOI22_X1 U3924 ( .A1(\mem[189][1] ), .A2(n4256), .B1(n6679), .B2(data_in[1]), 
        .ZN(n4257) );
  INV_X1 U3925 ( .A(n4258), .ZN(n5114) );
  AOI22_X1 U3926 ( .A1(\mem[189][2] ), .A2(n4256), .B1(n6679), .B2(data_in[2]), 
        .ZN(n4258) );
  INV_X1 U3927 ( .A(n4259), .ZN(n5113) );
  AOI22_X1 U3928 ( .A1(\mem[189][3] ), .A2(n4256), .B1(n6679), .B2(data_in[3]), 
        .ZN(n4259) );
  INV_X1 U3929 ( .A(n4260), .ZN(n5112) );
  AOI22_X1 U3930 ( .A1(\mem[189][4] ), .A2(n4256), .B1(n6679), .B2(data_in[4]), 
        .ZN(n4260) );
  INV_X1 U3931 ( .A(n4261), .ZN(n5111) );
  AOI22_X1 U3932 ( .A1(\mem[189][5] ), .A2(n4256), .B1(n6679), .B2(data_in[5]), 
        .ZN(n4261) );
  INV_X1 U3933 ( .A(n4262), .ZN(n5110) );
  AOI22_X1 U3934 ( .A1(\mem[189][6] ), .A2(n4256), .B1(n6679), .B2(data_in[6]), 
        .ZN(n4262) );
  INV_X1 U3935 ( .A(n4263), .ZN(n5109) );
  AOI22_X1 U3936 ( .A1(\mem[189][7] ), .A2(n4256), .B1(n6679), .B2(data_in[7]), 
        .ZN(n4263) );
  INV_X1 U3937 ( .A(n4264), .ZN(n5108) );
  AOI22_X1 U3938 ( .A1(\mem[190][0] ), .A2(n4265), .B1(n6678), .B2(data_in[0]), 
        .ZN(n4264) );
  INV_X1 U3939 ( .A(n4266), .ZN(n5107) );
  AOI22_X1 U3940 ( .A1(\mem[190][1] ), .A2(n4265), .B1(n6678), .B2(data_in[1]), 
        .ZN(n4266) );
  INV_X1 U3941 ( .A(n4267), .ZN(n5106) );
  AOI22_X1 U3942 ( .A1(\mem[190][2] ), .A2(n4265), .B1(n6678), .B2(data_in[2]), 
        .ZN(n4267) );
  INV_X1 U3943 ( .A(n4268), .ZN(n5105) );
  AOI22_X1 U3944 ( .A1(\mem[190][3] ), .A2(n4265), .B1(n6678), .B2(data_in[3]), 
        .ZN(n4268) );
  INV_X1 U3945 ( .A(n4269), .ZN(n5104) );
  AOI22_X1 U3946 ( .A1(\mem[190][4] ), .A2(n4265), .B1(n6678), .B2(data_in[4]), 
        .ZN(n4269) );
  INV_X1 U3947 ( .A(n4270), .ZN(n5103) );
  AOI22_X1 U3948 ( .A1(\mem[190][5] ), .A2(n4265), .B1(n6678), .B2(data_in[5]), 
        .ZN(n4270) );
  INV_X1 U3949 ( .A(n4271), .ZN(n5102) );
  AOI22_X1 U3950 ( .A1(\mem[190][6] ), .A2(n4265), .B1(n6678), .B2(data_in[6]), 
        .ZN(n4271) );
  INV_X1 U3951 ( .A(n4272), .ZN(n5101) );
  AOI22_X1 U3952 ( .A1(\mem[190][7] ), .A2(n4265), .B1(n6678), .B2(data_in[7]), 
        .ZN(n4272) );
  INV_X1 U3953 ( .A(n4273), .ZN(n5100) );
  AOI22_X1 U3954 ( .A1(\mem[191][0] ), .A2(n4274), .B1(n6677), .B2(data_in[0]), 
        .ZN(n4273) );
  INV_X1 U3955 ( .A(n4275), .ZN(n5099) );
  AOI22_X1 U3956 ( .A1(\mem[191][1] ), .A2(n4274), .B1(n6677), .B2(data_in[1]), 
        .ZN(n4275) );
  INV_X1 U3957 ( .A(n4276), .ZN(n5098) );
  AOI22_X1 U3958 ( .A1(\mem[191][2] ), .A2(n4274), .B1(n6677), .B2(data_in[2]), 
        .ZN(n4276) );
  INV_X1 U3959 ( .A(n4277), .ZN(n5097) );
  AOI22_X1 U3960 ( .A1(\mem[191][3] ), .A2(n4274), .B1(n6677), .B2(data_in[3]), 
        .ZN(n4277) );
  INV_X1 U3961 ( .A(n4278), .ZN(n5096) );
  AOI22_X1 U3962 ( .A1(\mem[191][4] ), .A2(n4274), .B1(n6677), .B2(data_in[4]), 
        .ZN(n4278) );
  INV_X1 U3963 ( .A(n4279), .ZN(n5095) );
  AOI22_X1 U3964 ( .A1(\mem[191][5] ), .A2(n4274), .B1(n6677), .B2(data_in[5]), 
        .ZN(n4279) );
  INV_X1 U3965 ( .A(n4280), .ZN(n5094) );
  AOI22_X1 U3966 ( .A1(\mem[191][6] ), .A2(n4274), .B1(n6677), .B2(data_in[6]), 
        .ZN(n4280) );
  INV_X1 U3967 ( .A(n4281), .ZN(n5093) );
  AOI22_X1 U3968 ( .A1(\mem[191][7] ), .A2(n4274), .B1(n6677), .B2(data_in[7]), 
        .ZN(n4281) );
  INV_X1 U3969 ( .A(n4282), .ZN(n5092) );
  AOI22_X1 U3970 ( .A1(\mem[192][0] ), .A2(n4283), .B1(n6676), .B2(data_in[0]), 
        .ZN(n4282) );
  INV_X1 U3971 ( .A(n4284), .ZN(n5091) );
  AOI22_X1 U3972 ( .A1(\mem[192][1] ), .A2(n4283), .B1(n6676), .B2(data_in[1]), 
        .ZN(n4284) );
  INV_X1 U3973 ( .A(n4285), .ZN(n5090) );
  AOI22_X1 U3974 ( .A1(\mem[192][2] ), .A2(n4283), .B1(n6676), .B2(data_in[2]), 
        .ZN(n4285) );
  INV_X1 U3975 ( .A(n4286), .ZN(n5089) );
  AOI22_X1 U3976 ( .A1(\mem[192][3] ), .A2(n4283), .B1(n6676), .B2(data_in[3]), 
        .ZN(n4286) );
  INV_X1 U3977 ( .A(n4287), .ZN(n5088) );
  AOI22_X1 U3978 ( .A1(\mem[192][4] ), .A2(n4283), .B1(n6676), .B2(data_in[4]), 
        .ZN(n4287) );
  INV_X1 U3979 ( .A(n4288), .ZN(n5087) );
  AOI22_X1 U3980 ( .A1(\mem[192][5] ), .A2(n4283), .B1(n6676), .B2(data_in[5]), 
        .ZN(n4288) );
  INV_X1 U3981 ( .A(n4289), .ZN(n5086) );
  AOI22_X1 U3982 ( .A1(\mem[192][6] ), .A2(n4283), .B1(n6676), .B2(data_in[6]), 
        .ZN(n4289) );
  INV_X1 U3983 ( .A(n4290), .ZN(n5085) );
  AOI22_X1 U3984 ( .A1(\mem[192][7] ), .A2(n4283), .B1(n6676), .B2(data_in[7]), 
        .ZN(n4290) );
  INV_X1 U3985 ( .A(n4292), .ZN(n5084) );
  AOI22_X1 U3986 ( .A1(\mem[193][0] ), .A2(n4293), .B1(n6675), .B2(data_in[0]), 
        .ZN(n4292) );
  INV_X1 U3987 ( .A(n4294), .ZN(n5083) );
  AOI22_X1 U3988 ( .A1(\mem[193][1] ), .A2(n4293), .B1(n6675), .B2(data_in[1]), 
        .ZN(n4294) );
  INV_X1 U3989 ( .A(n4295), .ZN(n5082) );
  AOI22_X1 U3990 ( .A1(\mem[193][2] ), .A2(n4293), .B1(n6675), .B2(data_in[2]), 
        .ZN(n4295) );
  INV_X1 U3991 ( .A(n4296), .ZN(n5081) );
  AOI22_X1 U3992 ( .A1(\mem[193][3] ), .A2(n4293), .B1(n6675), .B2(data_in[3]), 
        .ZN(n4296) );
  INV_X1 U3993 ( .A(n4297), .ZN(n5080) );
  AOI22_X1 U3994 ( .A1(\mem[193][4] ), .A2(n4293), .B1(n6675), .B2(data_in[4]), 
        .ZN(n4297) );
  INV_X1 U3995 ( .A(n4298), .ZN(n5079) );
  AOI22_X1 U3996 ( .A1(\mem[193][5] ), .A2(n4293), .B1(n6675), .B2(data_in[5]), 
        .ZN(n4298) );
  INV_X1 U3997 ( .A(n4299), .ZN(n5078) );
  AOI22_X1 U3998 ( .A1(\mem[193][6] ), .A2(n4293), .B1(n6675), .B2(data_in[6]), 
        .ZN(n4299) );
  INV_X1 U3999 ( .A(n4300), .ZN(n5077) );
  AOI22_X1 U4000 ( .A1(\mem[193][7] ), .A2(n4293), .B1(n6675), .B2(data_in[7]), 
        .ZN(n4300) );
  INV_X1 U4001 ( .A(n4301), .ZN(n5076) );
  AOI22_X1 U4002 ( .A1(\mem[194][0] ), .A2(n4302), .B1(n6674), .B2(data_in[0]), 
        .ZN(n4301) );
  INV_X1 U4003 ( .A(n4303), .ZN(n5075) );
  AOI22_X1 U4004 ( .A1(\mem[194][1] ), .A2(n4302), .B1(n6674), .B2(data_in[1]), 
        .ZN(n4303) );
  INV_X1 U4005 ( .A(n4304), .ZN(n5074) );
  AOI22_X1 U4006 ( .A1(\mem[194][2] ), .A2(n4302), .B1(n6674), .B2(data_in[2]), 
        .ZN(n4304) );
  INV_X1 U4007 ( .A(n4305), .ZN(n5073) );
  AOI22_X1 U4008 ( .A1(\mem[194][3] ), .A2(n4302), .B1(n6674), .B2(data_in[3]), 
        .ZN(n4305) );
  INV_X1 U4009 ( .A(n4306), .ZN(n5072) );
  AOI22_X1 U4010 ( .A1(\mem[194][4] ), .A2(n4302), .B1(n6674), .B2(data_in[4]), 
        .ZN(n4306) );
  INV_X1 U4011 ( .A(n4307), .ZN(n5071) );
  AOI22_X1 U4012 ( .A1(\mem[194][5] ), .A2(n4302), .B1(n6674), .B2(data_in[5]), 
        .ZN(n4307) );
  INV_X1 U4013 ( .A(n4308), .ZN(n5070) );
  AOI22_X1 U4014 ( .A1(\mem[194][6] ), .A2(n4302), .B1(n6674), .B2(data_in[6]), 
        .ZN(n4308) );
  INV_X1 U4015 ( .A(n4309), .ZN(n5069) );
  AOI22_X1 U4016 ( .A1(\mem[194][7] ), .A2(n4302), .B1(n6674), .B2(data_in[7]), 
        .ZN(n4309) );
  INV_X1 U4017 ( .A(n4310), .ZN(n5068) );
  AOI22_X1 U4018 ( .A1(\mem[195][0] ), .A2(n4311), .B1(n6673), .B2(data_in[0]), 
        .ZN(n4310) );
  INV_X1 U4019 ( .A(n4312), .ZN(n5067) );
  AOI22_X1 U4020 ( .A1(\mem[195][1] ), .A2(n4311), .B1(n6673), .B2(data_in[1]), 
        .ZN(n4312) );
  INV_X1 U4021 ( .A(n4313), .ZN(n5066) );
  AOI22_X1 U4022 ( .A1(\mem[195][2] ), .A2(n4311), .B1(n6673), .B2(data_in[2]), 
        .ZN(n4313) );
  INV_X1 U4023 ( .A(n4314), .ZN(n5065) );
  AOI22_X1 U4024 ( .A1(\mem[195][3] ), .A2(n4311), .B1(n6673), .B2(data_in[3]), 
        .ZN(n4314) );
  INV_X1 U4025 ( .A(n4315), .ZN(n5064) );
  AOI22_X1 U4026 ( .A1(\mem[195][4] ), .A2(n4311), .B1(n6673), .B2(data_in[4]), 
        .ZN(n4315) );
  INV_X1 U4027 ( .A(n4316), .ZN(n5063) );
  AOI22_X1 U4028 ( .A1(\mem[195][5] ), .A2(n4311), .B1(n6673), .B2(data_in[5]), 
        .ZN(n4316) );
  INV_X1 U4029 ( .A(n4317), .ZN(n5062) );
  AOI22_X1 U4030 ( .A1(\mem[195][6] ), .A2(n4311), .B1(n6673), .B2(data_in[6]), 
        .ZN(n4317) );
  INV_X1 U4031 ( .A(n4318), .ZN(n5061) );
  AOI22_X1 U4032 ( .A1(\mem[195][7] ), .A2(n4311), .B1(n6673), .B2(data_in[7]), 
        .ZN(n4318) );
  INV_X1 U4033 ( .A(n4319), .ZN(n5060) );
  AOI22_X1 U4034 ( .A1(\mem[196][0] ), .A2(n4320), .B1(n6672), .B2(data_in[0]), 
        .ZN(n4319) );
  INV_X1 U4035 ( .A(n4321), .ZN(n5059) );
  AOI22_X1 U4036 ( .A1(\mem[196][1] ), .A2(n4320), .B1(n6672), .B2(data_in[1]), 
        .ZN(n4321) );
  INV_X1 U4037 ( .A(n4322), .ZN(n5058) );
  AOI22_X1 U4038 ( .A1(\mem[196][2] ), .A2(n4320), .B1(n6672), .B2(data_in[2]), 
        .ZN(n4322) );
  INV_X1 U4039 ( .A(n4323), .ZN(n5057) );
  AOI22_X1 U4040 ( .A1(\mem[196][3] ), .A2(n4320), .B1(n6672), .B2(data_in[3]), 
        .ZN(n4323) );
  INV_X1 U4041 ( .A(n4324), .ZN(n5056) );
  AOI22_X1 U4042 ( .A1(\mem[196][4] ), .A2(n4320), .B1(n6672), .B2(data_in[4]), 
        .ZN(n4324) );
  INV_X1 U4043 ( .A(n4325), .ZN(n5055) );
  AOI22_X1 U4044 ( .A1(\mem[196][5] ), .A2(n4320), .B1(n6672), .B2(data_in[5]), 
        .ZN(n4325) );
  INV_X1 U4045 ( .A(n4326), .ZN(n5054) );
  AOI22_X1 U4046 ( .A1(\mem[196][6] ), .A2(n4320), .B1(n6672), .B2(data_in[6]), 
        .ZN(n4326) );
  INV_X1 U4047 ( .A(n4327), .ZN(n5053) );
  AOI22_X1 U4048 ( .A1(\mem[196][7] ), .A2(n4320), .B1(n6672), .B2(data_in[7]), 
        .ZN(n4327) );
  INV_X1 U4049 ( .A(n4328), .ZN(n5052) );
  AOI22_X1 U4050 ( .A1(\mem[197][0] ), .A2(n4329), .B1(n6671), .B2(data_in[0]), 
        .ZN(n4328) );
  INV_X1 U4051 ( .A(n4330), .ZN(n5051) );
  AOI22_X1 U4052 ( .A1(\mem[197][1] ), .A2(n4329), .B1(n6671), .B2(data_in[1]), 
        .ZN(n4330) );
  INV_X1 U4053 ( .A(n4331), .ZN(n5050) );
  AOI22_X1 U4054 ( .A1(\mem[197][2] ), .A2(n4329), .B1(n6671), .B2(data_in[2]), 
        .ZN(n4331) );
  INV_X1 U4055 ( .A(n4332), .ZN(n5049) );
  AOI22_X1 U4056 ( .A1(\mem[197][3] ), .A2(n4329), .B1(n6671), .B2(data_in[3]), 
        .ZN(n4332) );
  INV_X1 U4057 ( .A(n4333), .ZN(n5048) );
  AOI22_X1 U4058 ( .A1(\mem[197][4] ), .A2(n4329), .B1(n6671), .B2(data_in[4]), 
        .ZN(n4333) );
  INV_X1 U4059 ( .A(n4334), .ZN(n5047) );
  AOI22_X1 U4060 ( .A1(\mem[197][5] ), .A2(n4329), .B1(n6671), .B2(data_in[5]), 
        .ZN(n4334) );
  INV_X1 U4061 ( .A(n4335), .ZN(n5046) );
  AOI22_X1 U4062 ( .A1(\mem[197][6] ), .A2(n4329), .B1(n6671), .B2(data_in[6]), 
        .ZN(n4335) );
  INV_X1 U4063 ( .A(n4336), .ZN(n5045) );
  AOI22_X1 U4064 ( .A1(\mem[197][7] ), .A2(n4329), .B1(n6671), .B2(data_in[7]), 
        .ZN(n4336) );
  INV_X1 U4065 ( .A(n4337), .ZN(n5044) );
  AOI22_X1 U4066 ( .A1(\mem[198][0] ), .A2(n4338), .B1(n6670), .B2(data_in[0]), 
        .ZN(n4337) );
  INV_X1 U4067 ( .A(n4339), .ZN(n5043) );
  AOI22_X1 U4068 ( .A1(\mem[198][1] ), .A2(n4338), .B1(n6670), .B2(data_in[1]), 
        .ZN(n4339) );
  INV_X1 U4069 ( .A(n4340), .ZN(n5042) );
  AOI22_X1 U4070 ( .A1(\mem[198][2] ), .A2(n4338), .B1(n6670), .B2(data_in[2]), 
        .ZN(n4340) );
  INV_X1 U4071 ( .A(n4341), .ZN(n5041) );
  AOI22_X1 U4072 ( .A1(\mem[198][3] ), .A2(n4338), .B1(n6670), .B2(data_in[3]), 
        .ZN(n4341) );
  INV_X1 U4073 ( .A(n4342), .ZN(n5040) );
  AOI22_X1 U4074 ( .A1(\mem[198][4] ), .A2(n4338), .B1(n6670), .B2(data_in[4]), 
        .ZN(n4342) );
  INV_X1 U4075 ( .A(n4343), .ZN(n5039) );
  AOI22_X1 U4076 ( .A1(\mem[198][5] ), .A2(n4338), .B1(n6670), .B2(data_in[5]), 
        .ZN(n4343) );
  INV_X1 U4077 ( .A(n4344), .ZN(n5038) );
  AOI22_X1 U4078 ( .A1(\mem[198][6] ), .A2(n4338), .B1(n6670), .B2(data_in[6]), 
        .ZN(n4344) );
  INV_X1 U4079 ( .A(n4345), .ZN(n5037) );
  AOI22_X1 U4080 ( .A1(\mem[198][7] ), .A2(n4338), .B1(n6670), .B2(data_in[7]), 
        .ZN(n4345) );
  INV_X1 U4081 ( .A(n4346), .ZN(n5036) );
  AOI22_X1 U4082 ( .A1(\mem[199][0] ), .A2(n4347), .B1(n6669), .B2(data_in[0]), 
        .ZN(n4346) );
  INV_X1 U4083 ( .A(n4348), .ZN(n5035) );
  AOI22_X1 U4084 ( .A1(\mem[199][1] ), .A2(n4347), .B1(n6669), .B2(data_in[1]), 
        .ZN(n4348) );
  INV_X1 U4085 ( .A(n4349), .ZN(n5034) );
  AOI22_X1 U4086 ( .A1(\mem[199][2] ), .A2(n4347), .B1(n6669), .B2(data_in[2]), 
        .ZN(n4349) );
  INV_X1 U4087 ( .A(n4350), .ZN(n5033) );
  AOI22_X1 U4088 ( .A1(\mem[199][3] ), .A2(n4347), .B1(n6669), .B2(data_in[3]), 
        .ZN(n4350) );
  INV_X1 U4089 ( .A(n4351), .ZN(n5032) );
  AOI22_X1 U4090 ( .A1(\mem[199][4] ), .A2(n4347), .B1(n6669), .B2(data_in[4]), 
        .ZN(n4351) );
  INV_X1 U4091 ( .A(n4352), .ZN(n5031) );
  AOI22_X1 U4092 ( .A1(\mem[199][5] ), .A2(n4347), .B1(n6669), .B2(data_in[5]), 
        .ZN(n4352) );
  INV_X1 U4093 ( .A(n4353), .ZN(n5030) );
  AOI22_X1 U4094 ( .A1(\mem[199][6] ), .A2(n4347), .B1(n6669), .B2(data_in[6]), 
        .ZN(n4353) );
  INV_X1 U4095 ( .A(n4354), .ZN(n5029) );
  AOI22_X1 U4096 ( .A1(\mem[199][7] ), .A2(n4347), .B1(n6669), .B2(data_in[7]), 
        .ZN(n4354) );
  INV_X1 U4097 ( .A(n4355), .ZN(n5028) );
  AOI22_X1 U4098 ( .A1(\mem[200][0] ), .A2(n4356), .B1(n6668), .B2(data_in[0]), 
        .ZN(n4355) );
  INV_X1 U4099 ( .A(n4357), .ZN(n5027) );
  AOI22_X1 U4100 ( .A1(\mem[200][1] ), .A2(n4356), .B1(n6668), .B2(data_in[1]), 
        .ZN(n4357) );
  INV_X1 U4101 ( .A(n4358), .ZN(n5026) );
  AOI22_X1 U4102 ( .A1(\mem[200][2] ), .A2(n4356), .B1(n6668), .B2(data_in[2]), 
        .ZN(n4358) );
  INV_X1 U4103 ( .A(n4359), .ZN(n5025) );
  AOI22_X1 U4104 ( .A1(\mem[200][3] ), .A2(n4356), .B1(n6668), .B2(data_in[3]), 
        .ZN(n4359) );
  INV_X1 U4105 ( .A(n4360), .ZN(n5024) );
  AOI22_X1 U4106 ( .A1(\mem[200][4] ), .A2(n4356), .B1(n6668), .B2(data_in[4]), 
        .ZN(n4360) );
  INV_X1 U4107 ( .A(n4361), .ZN(n5023) );
  AOI22_X1 U4108 ( .A1(\mem[200][5] ), .A2(n4356), .B1(n6668), .B2(data_in[5]), 
        .ZN(n4361) );
  INV_X1 U4109 ( .A(n4362), .ZN(n5022) );
  AOI22_X1 U4110 ( .A1(\mem[200][6] ), .A2(n4356), .B1(n6668), .B2(data_in[6]), 
        .ZN(n4362) );
  INV_X1 U4111 ( .A(n4363), .ZN(n5021) );
  AOI22_X1 U4112 ( .A1(\mem[200][7] ), .A2(n4356), .B1(n6668), .B2(data_in[7]), 
        .ZN(n4363) );
  INV_X1 U4113 ( .A(n4364), .ZN(n5020) );
  AOI22_X1 U4114 ( .A1(\mem[201][0] ), .A2(n4365), .B1(n6667), .B2(data_in[0]), 
        .ZN(n4364) );
  INV_X1 U4115 ( .A(n4366), .ZN(n5019) );
  AOI22_X1 U4116 ( .A1(\mem[201][1] ), .A2(n4365), .B1(n6667), .B2(data_in[1]), 
        .ZN(n4366) );
  INV_X1 U4117 ( .A(n4367), .ZN(n5018) );
  AOI22_X1 U4118 ( .A1(\mem[201][2] ), .A2(n4365), .B1(n6667), .B2(data_in[2]), 
        .ZN(n4367) );
  INV_X1 U4119 ( .A(n4368), .ZN(n5017) );
  AOI22_X1 U4120 ( .A1(\mem[201][3] ), .A2(n4365), .B1(n6667), .B2(data_in[3]), 
        .ZN(n4368) );
  INV_X1 U4121 ( .A(n4369), .ZN(n5016) );
  AOI22_X1 U4122 ( .A1(\mem[201][4] ), .A2(n4365), .B1(n6667), .B2(data_in[4]), 
        .ZN(n4369) );
  INV_X1 U4123 ( .A(n4370), .ZN(n5015) );
  AOI22_X1 U4124 ( .A1(\mem[201][5] ), .A2(n4365), .B1(n6667), .B2(data_in[5]), 
        .ZN(n4370) );
  INV_X1 U4125 ( .A(n4371), .ZN(n5014) );
  AOI22_X1 U4126 ( .A1(\mem[201][6] ), .A2(n4365), .B1(n6667), .B2(data_in[6]), 
        .ZN(n4371) );
  INV_X1 U4127 ( .A(n4372), .ZN(n5013) );
  AOI22_X1 U4128 ( .A1(\mem[201][7] ), .A2(n4365), .B1(n6667), .B2(data_in[7]), 
        .ZN(n4372) );
  INV_X1 U4129 ( .A(n4373), .ZN(n5012) );
  AOI22_X1 U4130 ( .A1(\mem[202][0] ), .A2(n4374), .B1(n6666), .B2(data_in[0]), 
        .ZN(n4373) );
  INV_X1 U4131 ( .A(n4375), .ZN(n5011) );
  AOI22_X1 U4132 ( .A1(\mem[202][1] ), .A2(n4374), .B1(n6666), .B2(data_in[1]), 
        .ZN(n4375) );
  INV_X1 U4133 ( .A(n4376), .ZN(n5010) );
  AOI22_X1 U4134 ( .A1(\mem[202][2] ), .A2(n4374), .B1(n6666), .B2(data_in[2]), 
        .ZN(n4376) );
  INV_X1 U4135 ( .A(n4377), .ZN(n5009) );
  AOI22_X1 U4136 ( .A1(\mem[202][3] ), .A2(n4374), .B1(n6666), .B2(data_in[3]), 
        .ZN(n4377) );
  INV_X1 U4137 ( .A(n4378), .ZN(n5008) );
  AOI22_X1 U4138 ( .A1(\mem[202][4] ), .A2(n4374), .B1(n6666), .B2(data_in[4]), 
        .ZN(n4378) );
  INV_X1 U4139 ( .A(n4379), .ZN(n5007) );
  AOI22_X1 U4140 ( .A1(\mem[202][5] ), .A2(n4374), .B1(n6666), .B2(data_in[5]), 
        .ZN(n4379) );
  INV_X1 U4141 ( .A(n4380), .ZN(n5006) );
  AOI22_X1 U4142 ( .A1(\mem[202][6] ), .A2(n4374), .B1(n6666), .B2(data_in[6]), 
        .ZN(n4380) );
  INV_X1 U4143 ( .A(n4381), .ZN(n5005) );
  AOI22_X1 U4144 ( .A1(\mem[202][7] ), .A2(n4374), .B1(n6666), .B2(data_in[7]), 
        .ZN(n4381) );
  INV_X1 U4145 ( .A(n4382), .ZN(n5004) );
  AOI22_X1 U4146 ( .A1(\mem[203][0] ), .A2(n4383), .B1(n6665), .B2(data_in[0]), 
        .ZN(n4382) );
  INV_X1 U4147 ( .A(n4384), .ZN(n5003) );
  AOI22_X1 U4148 ( .A1(\mem[203][1] ), .A2(n4383), .B1(n6665), .B2(data_in[1]), 
        .ZN(n4384) );
  INV_X1 U4149 ( .A(n4385), .ZN(n5002) );
  AOI22_X1 U4150 ( .A1(\mem[203][2] ), .A2(n4383), .B1(n6665), .B2(data_in[2]), 
        .ZN(n4385) );
  INV_X1 U4151 ( .A(n4386), .ZN(n5001) );
  AOI22_X1 U4152 ( .A1(\mem[203][3] ), .A2(n4383), .B1(n6665), .B2(data_in[3]), 
        .ZN(n4386) );
  INV_X1 U4153 ( .A(n4387), .ZN(n5000) );
  AOI22_X1 U4154 ( .A1(\mem[203][4] ), .A2(n4383), .B1(n6665), .B2(data_in[4]), 
        .ZN(n4387) );
  INV_X1 U4155 ( .A(n4388), .ZN(n4999) );
  AOI22_X1 U4156 ( .A1(\mem[203][5] ), .A2(n4383), .B1(n6665), .B2(data_in[5]), 
        .ZN(n4388) );
  INV_X1 U4157 ( .A(n4389), .ZN(n4998) );
  AOI22_X1 U4158 ( .A1(\mem[203][6] ), .A2(n4383), .B1(n6665), .B2(data_in[6]), 
        .ZN(n4389) );
  INV_X1 U4159 ( .A(n4390), .ZN(n4997) );
  AOI22_X1 U4160 ( .A1(\mem[203][7] ), .A2(n4383), .B1(n6665), .B2(data_in[7]), 
        .ZN(n4390) );
  INV_X1 U4161 ( .A(n4391), .ZN(n4996) );
  AOI22_X1 U4162 ( .A1(\mem[204][0] ), .A2(n4392), .B1(n6664), .B2(data_in[0]), 
        .ZN(n4391) );
  INV_X1 U4163 ( .A(n4393), .ZN(n4995) );
  AOI22_X1 U4164 ( .A1(\mem[204][1] ), .A2(n4392), .B1(n6664), .B2(data_in[1]), 
        .ZN(n4393) );
  INV_X1 U4165 ( .A(n4394), .ZN(n4994) );
  AOI22_X1 U4166 ( .A1(\mem[204][2] ), .A2(n4392), .B1(n6664), .B2(data_in[2]), 
        .ZN(n4394) );
  INV_X1 U4167 ( .A(n4395), .ZN(n4993) );
  AOI22_X1 U4168 ( .A1(\mem[204][3] ), .A2(n4392), .B1(n6664), .B2(data_in[3]), 
        .ZN(n4395) );
  INV_X1 U4169 ( .A(n4396), .ZN(n4992) );
  AOI22_X1 U4170 ( .A1(\mem[204][4] ), .A2(n4392), .B1(n6664), .B2(data_in[4]), 
        .ZN(n4396) );
  INV_X1 U4171 ( .A(n4397), .ZN(n4991) );
  AOI22_X1 U4172 ( .A1(\mem[204][5] ), .A2(n4392), .B1(n6664), .B2(data_in[5]), 
        .ZN(n4397) );
  INV_X1 U4173 ( .A(n4398), .ZN(n4990) );
  AOI22_X1 U4174 ( .A1(\mem[204][6] ), .A2(n4392), .B1(n6664), .B2(data_in[6]), 
        .ZN(n4398) );
  INV_X1 U4175 ( .A(n4399), .ZN(n4989) );
  AOI22_X1 U4176 ( .A1(\mem[204][7] ), .A2(n4392), .B1(n6664), .B2(data_in[7]), 
        .ZN(n4399) );
  INV_X1 U4177 ( .A(n4400), .ZN(n4988) );
  AOI22_X1 U4178 ( .A1(\mem[205][0] ), .A2(n4401), .B1(n6663), .B2(data_in[0]), 
        .ZN(n4400) );
  INV_X1 U4179 ( .A(n4402), .ZN(n4987) );
  AOI22_X1 U4180 ( .A1(\mem[205][1] ), .A2(n4401), .B1(n6663), .B2(data_in[1]), 
        .ZN(n4402) );
  INV_X1 U4181 ( .A(n4403), .ZN(n4986) );
  AOI22_X1 U4182 ( .A1(\mem[205][2] ), .A2(n4401), .B1(n6663), .B2(data_in[2]), 
        .ZN(n4403) );
  INV_X1 U4183 ( .A(n4404), .ZN(n4985) );
  AOI22_X1 U4184 ( .A1(\mem[205][3] ), .A2(n4401), .B1(n6663), .B2(data_in[3]), 
        .ZN(n4404) );
  INV_X1 U4185 ( .A(n4405), .ZN(n4984) );
  AOI22_X1 U4186 ( .A1(\mem[205][4] ), .A2(n4401), .B1(n6663), .B2(data_in[4]), 
        .ZN(n4405) );
  INV_X1 U4187 ( .A(n4406), .ZN(n4983) );
  AOI22_X1 U4188 ( .A1(\mem[205][5] ), .A2(n4401), .B1(n6663), .B2(data_in[5]), 
        .ZN(n4406) );
  INV_X1 U4189 ( .A(n4407), .ZN(n4982) );
  AOI22_X1 U4190 ( .A1(\mem[205][6] ), .A2(n4401), .B1(n6663), .B2(data_in[6]), 
        .ZN(n4407) );
  INV_X1 U4191 ( .A(n4408), .ZN(n4981) );
  AOI22_X1 U4192 ( .A1(\mem[205][7] ), .A2(n4401), .B1(n6663), .B2(data_in[7]), 
        .ZN(n4408) );
  INV_X1 U4193 ( .A(n4409), .ZN(n4980) );
  AOI22_X1 U4194 ( .A1(\mem[206][0] ), .A2(n4410), .B1(n6662), .B2(data_in[0]), 
        .ZN(n4409) );
  INV_X1 U4195 ( .A(n4411), .ZN(n4979) );
  AOI22_X1 U4196 ( .A1(\mem[206][1] ), .A2(n4410), .B1(n6662), .B2(data_in[1]), 
        .ZN(n4411) );
  INV_X1 U4197 ( .A(n4412), .ZN(n4978) );
  AOI22_X1 U4198 ( .A1(\mem[206][2] ), .A2(n4410), .B1(n6662), .B2(data_in[2]), 
        .ZN(n4412) );
  INV_X1 U4199 ( .A(n4413), .ZN(n4977) );
  AOI22_X1 U4200 ( .A1(\mem[206][3] ), .A2(n4410), .B1(n6662), .B2(data_in[3]), 
        .ZN(n4413) );
  INV_X1 U4201 ( .A(n4414), .ZN(n4976) );
  AOI22_X1 U4202 ( .A1(\mem[206][4] ), .A2(n4410), .B1(n6662), .B2(data_in[4]), 
        .ZN(n4414) );
  INV_X1 U4203 ( .A(n4415), .ZN(n4975) );
  AOI22_X1 U4204 ( .A1(\mem[206][5] ), .A2(n4410), .B1(n6662), .B2(data_in[5]), 
        .ZN(n4415) );
  INV_X1 U4205 ( .A(n4416), .ZN(n4974) );
  AOI22_X1 U4206 ( .A1(\mem[206][6] ), .A2(n4410), .B1(n6662), .B2(data_in[6]), 
        .ZN(n4416) );
  INV_X1 U4207 ( .A(n4417), .ZN(n4973) );
  AOI22_X1 U4208 ( .A1(\mem[206][7] ), .A2(n4410), .B1(n6662), .B2(data_in[7]), 
        .ZN(n4417) );
  INV_X1 U4209 ( .A(n4418), .ZN(n4972) );
  AOI22_X1 U4210 ( .A1(\mem[207][0] ), .A2(n4419), .B1(n6661), .B2(data_in[0]), 
        .ZN(n4418) );
  INV_X1 U4211 ( .A(n4420), .ZN(n4971) );
  AOI22_X1 U4212 ( .A1(\mem[207][1] ), .A2(n4419), .B1(n6661), .B2(data_in[1]), 
        .ZN(n4420) );
  INV_X1 U4213 ( .A(n4421), .ZN(n4970) );
  AOI22_X1 U4214 ( .A1(\mem[207][2] ), .A2(n4419), .B1(n6661), .B2(data_in[2]), 
        .ZN(n4421) );
  INV_X1 U4215 ( .A(n4422), .ZN(n4969) );
  AOI22_X1 U4216 ( .A1(\mem[207][3] ), .A2(n4419), .B1(n6661), .B2(data_in[3]), 
        .ZN(n4422) );
  INV_X1 U4217 ( .A(n4423), .ZN(n4968) );
  AOI22_X1 U4218 ( .A1(\mem[207][4] ), .A2(n4419), .B1(n6661), .B2(data_in[4]), 
        .ZN(n4423) );
  INV_X1 U4219 ( .A(n4424), .ZN(n4967) );
  AOI22_X1 U4220 ( .A1(\mem[207][5] ), .A2(n4419), .B1(n6661), .B2(data_in[5]), 
        .ZN(n4424) );
  INV_X1 U4221 ( .A(n4425), .ZN(n4966) );
  AOI22_X1 U4222 ( .A1(\mem[207][6] ), .A2(n4419), .B1(n6661), .B2(data_in[6]), 
        .ZN(n4425) );
  INV_X1 U4223 ( .A(n4426), .ZN(n4965) );
  AOI22_X1 U4224 ( .A1(\mem[207][7] ), .A2(n4419), .B1(n6661), .B2(data_in[7]), 
        .ZN(n4426) );
  INV_X1 U4225 ( .A(n4427), .ZN(n4964) );
  AOI22_X1 U4226 ( .A1(\mem[208][0] ), .A2(n4428), .B1(n6660), .B2(data_in[0]), 
        .ZN(n4427) );
  INV_X1 U4227 ( .A(n4429), .ZN(n4963) );
  AOI22_X1 U4228 ( .A1(\mem[208][1] ), .A2(n4428), .B1(n6660), .B2(data_in[1]), 
        .ZN(n4429) );
  INV_X1 U4229 ( .A(n4430), .ZN(n4962) );
  AOI22_X1 U4230 ( .A1(\mem[208][2] ), .A2(n4428), .B1(n6660), .B2(data_in[2]), 
        .ZN(n4430) );
  INV_X1 U4231 ( .A(n4431), .ZN(n4961) );
  AOI22_X1 U4232 ( .A1(\mem[208][3] ), .A2(n4428), .B1(n6660), .B2(data_in[3]), 
        .ZN(n4431) );
  INV_X1 U4233 ( .A(n4432), .ZN(n4960) );
  AOI22_X1 U4234 ( .A1(\mem[208][4] ), .A2(n4428), .B1(n6660), .B2(data_in[4]), 
        .ZN(n4432) );
  INV_X1 U4235 ( .A(n4433), .ZN(n4959) );
  AOI22_X1 U4236 ( .A1(\mem[208][5] ), .A2(n4428), .B1(n6660), .B2(data_in[5]), 
        .ZN(n4433) );
  INV_X1 U4237 ( .A(n4434), .ZN(n4958) );
  AOI22_X1 U4238 ( .A1(\mem[208][6] ), .A2(n4428), .B1(n6660), .B2(data_in[6]), 
        .ZN(n4434) );
  INV_X1 U4239 ( .A(n4435), .ZN(n4957) );
  AOI22_X1 U4240 ( .A1(\mem[208][7] ), .A2(n4428), .B1(n6660), .B2(data_in[7]), 
        .ZN(n4435) );
  INV_X1 U4241 ( .A(n4437), .ZN(n4956) );
  AOI22_X1 U4242 ( .A1(\mem[209][0] ), .A2(n4438), .B1(n6659), .B2(data_in[0]), 
        .ZN(n4437) );
  INV_X1 U4243 ( .A(n4439), .ZN(n4955) );
  AOI22_X1 U4244 ( .A1(\mem[209][1] ), .A2(n4438), .B1(n6659), .B2(data_in[1]), 
        .ZN(n4439) );
  INV_X1 U4245 ( .A(n4440), .ZN(n4954) );
  AOI22_X1 U4246 ( .A1(\mem[209][2] ), .A2(n4438), .B1(n6659), .B2(data_in[2]), 
        .ZN(n4440) );
  INV_X1 U4247 ( .A(n4441), .ZN(n4953) );
  AOI22_X1 U4248 ( .A1(\mem[209][3] ), .A2(n4438), .B1(n6659), .B2(data_in[3]), 
        .ZN(n4441) );
  INV_X1 U4249 ( .A(n4442), .ZN(n4952) );
  AOI22_X1 U4250 ( .A1(\mem[209][4] ), .A2(n4438), .B1(n6659), .B2(data_in[4]), 
        .ZN(n4442) );
  INV_X1 U4251 ( .A(n4443), .ZN(n4951) );
  AOI22_X1 U4252 ( .A1(\mem[209][5] ), .A2(n4438), .B1(n6659), .B2(data_in[5]), 
        .ZN(n4443) );
  INV_X1 U4253 ( .A(n4444), .ZN(n4950) );
  AOI22_X1 U4254 ( .A1(\mem[209][6] ), .A2(n4438), .B1(n6659), .B2(data_in[6]), 
        .ZN(n4444) );
  INV_X1 U4255 ( .A(n4445), .ZN(n4949) );
  AOI22_X1 U4256 ( .A1(\mem[209][7] ), .A2(n4438), .B1(n6659), .B2(data_in[7]), 
        .ZN(n4445) );
  INV_X1 U4257 ( .A(n4446), .ZN(n4948) );
  AOI22_X1 U4258 ( .A1(\mem[210][0] ), .A2(n4447), .B1(n6658), .B2(data_in[0]), 
        .ZN(n4446) );
  INV_X1 U4259 ( .A(n4448), .ZN(n4947) );
  AOI22_X1 U4260 ( .A1(\mem[210][1] ), .A2(n4447), .B1(n6658), .B2(data_in[1]), 
        .ZN(n4448) );
  INV_X1 U4261 ( .A(n4449), .ZN(n4946) );
  AOI22_X1 U4262 ( .A1(\mem[210][2] ), .A2(n4447), .B1(n6658), .B2(data_in[2]), 
        .ZN(n4449) );
  INV_X1 U4263 ( .A(n4450), .ZN(n4945) );
  AOI22_X1 U4264 ( .A1(\mem[210][3] ), .A2(n4447), .B1(n6658), .B2(data_in[3]), 
        .ZN(n4450) );
  INV_X1 U4265 ( .A(n4451), .ZN(n4944) );
  AOI22_X1 U4266 ( .A1(\mem[210][4] ), .A2(n4447), .B1(n6658), .B2(data_in[4]), 
        .ZN(n4451) );
  INV_X1 U4267 ( .A(n4452), .ZN(n4943) );
  AOI22_X1 U4268 ( .A1(\mem[210][5] ), .A2(n4447), .B1(n6658), .B2(data_in[5]), 
        .ZN(n4452) );
  INV_X1 U4269 ( .A(n4453), .ZN(n4942) );
  AOI22_X1 U4270 ( .A1(\mem[210][6] ), .A2(n4447), .B1(n6658), .B2(data_in[6]), 
        .ZN(n4453) );
  INV_X1 U4271 ( .A(n4454), .ZN(n4941) );
  AOI22_X1 U4272 ( .A1(\mem[210][7] ), .A2(n4447), .B1(n6658), .B2(data_in[7]), 
        .ZN(n4454) );
  INV_X1 U4273 ( .A(n4455), .ZN(n4940) );
  AOI22_X1 U4274 ( .A1(\mem[211][0] ), .A2(n4456), .B1(n6657), .B2(data_in[0]), 
        .ZN(n4455) );
  INV_X1 U4275 ( .A(n4457), .ZN(n4939) );
  AOI22_X1 U4276 ( .A1(\mem[211][1] ), .A2(n4456), .B1(n6657), .B2(data_in[1]), 
        .ZN(n4457) );
  INV_X1 U4277 ( .A(n4458), .ZN(n4938) );
  AOI22_X1 U4278 ( .A1(\mem[211][2] ), .A2(n4456), .B1(n6657), .B2(data_in[2]), 
        .ZN(n4458) );
  INV_X1 U4279 ( .A(n4459), .ZN(n4937) );
  AOI22_X1 U4280 ( .A1(\mem[211][3] ), .A2(n4456), .B1(n6657), .B2(data_in[3]), 
        .ZN(n4459) );
  INV_X1 U4281 ( .A(n4460), .ZN(n4936) );
  AOI22_X1 U4282 ( .A1(\mem[211][4] ), .A2(n4456), .B1(n6657), .B2(data_in[4]), 
        .ZN(n4460) );
  INV_X1 U4283 ( .A(n4461), .ZN(n4935) );
  AOI22_X1 U4284 ( .A1(\mem[211][5] ), .A2(n4456), .B1(n6657), .B2(data_in[5]), 
        .ZN(n4461) );
  INV_X1 U4285 ( .A(n4462), .ZN(n4934) );
  AOI22_X1 U4286 ( .A1(\mem[211][6] ), .A2(n4456), .B1(n6657), .B2(data_in[6]), 
        .ZN(n4462) );
  INV_X1 U4287 ( .A(n4463), .ZN(n4933) );
  AOI22_X1 U4288 ( .A1(\mem[211][7] ), .A2(n4456), .B1(n6657), .B2(data_in[7]), 
        .ZN(n4463) );
  INV_X1 U4289 ( .A(n4464), .ZN(n4932) );
  AOI22_X1 U4290 ( .A1(\mem[212][0] ), .A2(n4465), .B1(n6656), .B2(data_in[0]), 
        .ZN(n4464) );
  INV_X1 U4291 ( .A(n4466), .ZN(n4931) );
  AOI22_X1 U4292 ( .A1(\mem[212][1] ), .A2(n4465), .B1(n6656), .B2(data_in[1]), 
        .ZN(n4466) );
  INV_X1 U4293 ( .A(n4467), .ZN(n4930) );
  AOI22_X1 U4294 ( .A1(\mem[212][2] ), .A2(n4465), .B1(n6656), .B2(data_in[2]), 
        .ZN(n4467) );
  INV_X1 U4295 ( .A(n4468), .ZN(n4929) );
  AOI22_X1 U4296 ( .A1(\mem[212][3] ), .A2(n4465), .B1(n6656), .B2(data_in[3]), 
        .ZN(n4468) );
  INV_X1 U4297 ( .A(n4469), .ZN(n4928) );
  AOI22_X1 U4298 ( .A1(\mem[212][4] ), .A2(n4465), .B1(n6656), .B2(data_in[4]), 
        .ZN(n4469) );
  INV_X1 U4299 ( .A(n4470), .ZN(n4927) );
  AOI22_X1 U4300 ( .A1(\mem[212][5] ), .A2(n4465), .B1(n6656), .B2(data_in[5]), 
        .ZN(n4470) );
  INV_X1 U4301 ( .A(n4471), .ZN(n4926) );
  AOI22_X1 U4302 ( .A1(\mem[212][6] ), .A2(n4465), .B1(n6656), .B2(data_in[6]), 
        .ZN(n4471) );
  INV_X1 U4303 ( .A(n4472), .ZN(n4925) );
  AOI22_X1 U4304 ( .A1(\mem[212][7] ), .A2(n4465), .B1(n6656), .B2(data_in[7]), 
        .ZN(n4472) );
  INV_X1 U4305 ( .A(n4473), .ZN(n4924) );
  AOI22_X1 U4306 ( .A1(\mem[213][0] ), .A2(n4474), .B1(n6655), .B2(data_in[0]), 
        .ZN(n4473) );
  INV_X1 U4307 ( .A(n4475), .ZN(n4923) );
  AOI22_X1 U4308 ( .A1(\mem[213][1] ), .A2(n4474), .B1(n6655), .B2(data_in[1]), 
        .ZN(n4475) );
  INV_X1 U4309 ( .A(n4476), .ZN(n4922) );
  AOI22_X1 U4310 ( .A1(\mem[213][2] ), .A2(n4474), .B1(n6655), .B2(data_in[2]), 
        .ZN(n4476) );
  INV_X1 U4311 ( .A(n4477), .ZN(n4921) );
  AOI22_X1 U4312 ( .A1(\mem[213][3] ), .A2(n4474), .B1(n6655), .B2(data_in[3]), 
        .ZN(n4477) );
  INV_X1 U4313 ( .A(n4478), .ZN(n4920) );
  AOI22_X1 U4314 ( .A1(\mem[213][4] ), .A2(n4474), .B1(n6655), .B2(data_in[4]), 
        .ZN(n4478) );
  INV_X1 U4315 ( .A(n4479), .ZN(n4919) );
  AOI22_X1 U4316 ( .A1(\mem[213][5] ), .A2(n4474), .B1(n6655), .B2(data_in[5]), 
        .ZN(n4479) );
  INV_X1 U4317 ( .A(n4480), .ZN(n4918) );
  AOI22_X1 U4318 ( .A1(\mem[213][6] ), .A2(n4474), .B1(n6655), .B2(data_in[6]), 
        .ZN(n4480) );
  INV_X1 U4319 ( .A(n4481), .ZN(n4917) );
  AOI22_X1 U4320 ( .A1(\mem[213][7] ), .A2(n4474), .B1(n6655), .B2(data_in[7]), 
        .ZN(n4481) );
  INV_X1 U4321 ( .A(n4482), .ZN(n4916) );
  AOI22_X1 U4322 ( .A1(\mem[214][0] ), .A2(n4483), .B1(n6654), .B2(data_in[0]), 
        .ZN(n4482) );
  INV_X1 U4323 ( .A(n4484), .ZN(n4915) );
  AOI22_X1 U4324 ( .A1(\mem[214][1] ), .A2(n4483), .B1(n6654), .B2(data_in[1]), 
        .ZN(n4484) );
  INV_X1 U4325 ( .A(n4485), .ZN(n4914) );
  AOI22_X1 U4326 ( .A1(\mem[214][2] ), .A2(n4483), .B1(n6654), .B2(data_in[2]), 
        .ZN(n4485) );
  INV_X1 U4327 ( .A(n4486), .ZN(n4913) );
  AOI22_X1 U4328 ( .A1(\mem[214][3] ), .A2(n4483), .B1(n6654), .B2(data_in[3]), 
        .ZN(n4486) );
  INV_X1 U4329 ( .A(n4487), .ZN(n4912) );
  AOI22_X1 U4330 ( .A1(\mem[214][4] ), .A2(n4483), .B1(n6654), .B2(data_in[4]), 
        .ZN(n4487) );
  INV_X1 U4331 ( .A(n4488), .ZN(n4911) );
  AOI22_X1 U4332 ( .A1(\mem[214][5] ), .A2(n4483), .B1(n6654), .B2(data_in[5]), 
        .ZN(n4488) );
  INV_X1 U4333 ( .A(n4489), .ZN(n4910) );
  AOI22_X1 U4334 ( .A1(\mem[214][6] ), .A2(n4483), .B1(n6654), .B2(data_in[6]), 
        .ZN(n4489) );
  INV_X1 U4335 ( .A(n4490), .ZN(n4909) );
  AOI22_X1 U4336 ( .A1(\mem[214][7] ), .A2(n4483), .B1(n6654), .B2(data_in[7]), 
        .ZN(n4490) );
  INV_X1 U4337 ( .A(n4491), .ZN(n4908) );
  AOI22_X1 U4338 ( .A1(\mem[215][0] ), .A2(n4492), .B1(n6653), .B2(data_in[0]), 
        .ZN(n4491) );
  INV_X1 U4339 ( .A(n4493), .ZN(n4907) );
  AOI22_X1 U4340 ( .A1(\mem[215][1] ), .A2(n4492), .B1(n6653), .B2(data_in[1]), 
        .ZN(n4493) );
  INV_X1 U4341 ( .A(n4494), .ZN(n4906) );
  AOI22_X1 U4342 ( .A1(\mem[215][2] ), .A2(n4492), .B1(n6653), .B2(data_in[2]), 
        .ZN(n4494) );
  INV_X1 U4343 ( .A(n4495), .ZN(n4905) );
  AOI22_X1 U4344 ( .A1(\mem[215][3] ), .A2(n4492), .B1(n6653), .B2(data_in[3]), 
        .ZN(n4495) );
  INV_X1 U4345 ( .A(n4496), .ZN(n4904) );
  AOI22_X1 U4346 ( .A1(\mem[215][4] ), .A2(n4492), .B1(n6653), .B2(data_in[4]), 
        .ZN(n4496) );
  INV_X1 U4347 ( .A(n4497), .ZN(n4903) );
  AOI22_X1 U4348 ( .A1(\mem[215][5] ), .A2(n4492), .B1(n6653), .B2(data_in[5]), 
        .ZN(n4497) );
  INV_X1 U4349 ( .A(n4498), .ZN(n4902) );
  AOI22_X1 U4350 ( .A1(\mem[215][6] ), .A2(n4492), .B1(n6653), .B2(data_in[6]), 
        .ZN(n4498) );
  INV_X1 U4351 ( .A(n4499), .ZN(n4901) );
  AOI22_X1 U4352 ( .A1(\mem[215][7] ), .A2(n4492), .B1(n6653), .B2(data_in[7]), 
        .ZN(n4499) );
  INV_X1 U4353 ( .A(n4500), .ZN(n4900) );
  AOI22_X1 U4354 ( .A1(\mem[216][0] ), .A2(n4501), .B1(n6652), .B2(data_in[0]), 
        .ZN(n4500) );
  INV_X1 U4355 ( .A(n4502), .ZN(n4899) );
  AOI22_X1 U4356 ( .A1(\mem[216][1] ), .A2(n4501), .B1(n6652), .B2(data_in[1]), 
        .ZN(n4502) );
  INV_X1 U4357 ( .A(n4503), .ZN(n4898) );
  AOI22_X1 U4358 ( .A1(\mem[216][2] ), .A2(n4501), .B1(n6652), .B2(data_in[2]), 
        .ZN(n4503) );
  INV_X1 U4359 ( .A(n4504), .ZN(n4897) );
  AOI22_X1 U4360 ( .A1(\mem[216][3] ), .A2(n4501), .B1(n6652), .B2(data_in[3]), 
        .ZN(n4504) );
  INV_X1 U4361 ( .A(n4505), .ZN(n4896) );
  AOI22_X1 U4362 ( .A1(\mem[216][4] ), .A2(n4501), .B1(n6652), .B2(data_in[4]), 
        .ZN(n4505) );
  INV_X1 U4363 ( .A(n4506), .ZN(n4895) );
  AOI22_X1 U4364 ( .A1(\mem[216][5] ), .A2(n4501), .B1(n6652), .B2(data_in[5]), 
        .ZN(n4506) );
  INV_X1 U4365 ( .A(n4507), .ZN(n4894) );
  AOI22_X1 U4366 ( .A1(\mem[216][6] ), .A2(n4501), .B1(n6652), .B2(data_in[6]), 
        .ZN(n4507) );
  INV_X1 U4367 ( .A(n4508), .ZN(n4893) );
  AOI22_X1 U4368 ( .A1(\mem[216][7] ), .A2(n4501), .B1(n6652), .B2(data_in[7]), 
        .ZN(n4508) );
  INV_X1 U4369 ( .A(n4509), .ZN(n4892) );
  AOI22_X1 U4370 ( .A1(\mem[217][0] ), .A2(n4510), .B1(n6651), .B2(data_in[0]), 
        .ZN(n4509) );
  INV_X1 U4371 ( .A(n4511), .ZN(n4891) );
  AOI22_X1 U4372 ( .A1(\mem[217][1] ), .A2(n4510), .B1(n6651), .B2(data_in[1]), 
        .ZN(n4511) );
  INV_X1 U4373 ( .A(n4512), .ZN(n4890) );
  AOI22_X1 U4374 ( .A1(\mem[217][2] ), .A2(n4510), .B1(n6651), .B2(data_in[2]), 
        .ZN(n4512) );
  INV_X1 U4375 ( .A(n4513), .ZN(n4889) );
  AOI22_X1 U4376 ( .A1(\mem[217][3] ), .A2(n4510), .B1(n6651), .B2(data_in[3]), 
        .ZN(n4513) );
  INV_X1 U4377 ( .A(n4514), .ZN(n4888) );
  AOI22_X1 U4378 ( .A1(\mem[217][4] ), .A2(n4510), .B1(n6651), .B2(data_in[4]), 
        .ZN(n4514) );
  INV_X1 U4379 ( .A(n4515), .ZN(n4887) );
  AOI22_X1 U4380 ( .A1(\mem[217][5] ), .A2(n4510), .B1(n6651), .B2(data_in[5]), 
        .ZN(n4515) );
  INV_X1 U4381 ( .A(n4516), .ZN(n4886) );
  AOI22_X1 U4382 ( .A1(\mem[217][6] ), .A2(n4510), .B1(n6651), .B2(data_in[6]), 
        .ZN(n4516) );
  INV_X1 U4383 ( .A(n4517), .ZN(n4885) );
  AOI22_X1 U4384 ( .A1(\mem[217][7] ), .A2(n4510), .B1(n6651), .B2(data_in[7]), 
        .ZN(n4517) );
  INV_X1 U4385 ( .A(n4518), .ZN(n4884) );
  AOI22_X1 U4386 ( .A1(\mem[218][0] ), .A2(n4519), .B1(n6650), .B2(data_in[0]), 
        .ZN(n4518) );
  INV_X1 U4387 ( .A(n4520), .ZN(n4883) );
  AOI22_X1 U4388 ( .A1(\mem[218][1] ), .A2(n4519), .B1(n6650), .B2(data_in[1]), 
        .ZN(n4520) );
  INV_X1 U4389 ( .A(n4521), .ZN(n4882) );
  AOI22_X1 U4390 ( .A1(\mem[218][2] ), .A2(n4519), .B1(n6650), .B2(data_in[2]), 
        .ZN(n4521) );
  INV_X1 U4391 ( .A(n4522), .ZN(n4881) );
  AOI22_X1 U4392 ( .A1(\mem[218][3] ), .A2(n4519), .B1(n6650), .B2(data_in[3]), 
        .ZN(n4522) );
  INV_X1 U4393 ( .A(n4523), .ZN(n4880) );
  AOI22_X1 U4394 ( .A1(\mem[218][4] ), .A2(n4519), .B1(n6650), .B2(data_in[4]), 
        .ZN(n4523) );
  INV_X1 U4395 ( .A(n4524), .ZN(n4879) );
  AOI22_X1 U4396 ( .A1(\mem[218][5] ), .A2(n4519), .B1(n6650), .B2(data_in[5]), 
        .ZN(n4524) );
  INV_X1 U4397 ( .A(n4525), .ZN(n4878) );
  AOI22_X1 U4398 ( .A1(\mem[218][6] ), .A2(n4519), .B1(n6650), .B2(data_in[6]), 
        .ZN(n4525) );
  INV_X1 U4399 ( .A(n4526), .ZN(n4877) );
  AOI22_X1 U4400 ( .A1(\mem[218][7] ), .A2(n4519), .B1(n6650), .B2(data_in[7]), 
        .ZN(n4526) );
  INV_X1 U4401 ( .A(n4529), .ZN(n4876) );
  AOI22_X1 U4402 ( .A1(\mem[219][0] ), .A2(n4530), .B1(n6649), .B2(data_in[0]), 
        .ZN(n4529) );
  INV_X1 U4403 ( .A(n4531), .ZN(n4875) );
  AOI22_X1 U4404 ( .A1(\mem[219][1] ), .A2(n4530), .B1(n6649), .B2(data_in[1]), 
        .ZN(n4531) );
  INV_X1 U4405 ( .A(n4532), .ZN(n4874) );
  AOI22_X1 U4406 ( .A1(\mem[219][2] ), .A2(n4530), .B1(n6649), .B2(data_in[2]), 
        .ZN(n4532) );
  INV_X1 U4407 ( .A(n4533), .ZN(n4873) );
  AOI22_X1 U4408 ( .A1(\mem[219][3] ), .A2(n4530), .B1(n6649), .B2(data_in[3]), 
        .ZN(n4533) );
  INV_X1 U4409 ( .A(n4534), .ZN(n4872) );
  AOI22_X1 U4410 ( .A1(\mem[219][4] ), .A2(n4530), .B1(n6649), .B2(data_in[4]), 
        .ZN(n4534) );
  INV_X1 U4411 ( .A(n4535), .ZN(n4871) );
  AOI22_X1 U4412 ( .A1(\mem[219][5] ), .A2(n4530), .B1(n6649), .B2(data_in[5]), 
        .ZN(n4535) );
  INV_X1 U4413 ( .A(n4536), .ZN(n4870) );
  AOI22_X1 U4414 ( .A1(\mem[219][6] ), .A2(n4530), .B1(n6649), .B2(data_in[6]), 
        .ZN(n4536) );
  INV_X1 U4415 ( .A(n4537), .ZN(n4869) );
  AOI22_X1 U4416 ( .A1(\mem[219][7] ), .A2(n4530), .B1(n6649), .B2(data_in[7]), 
        .ZN(n4537) );
  INV_X1 U4417 ( .A(n4539), .ZN(n4868) );
  AOI22_X1 U4418 ( .A1(\mem[220][0] ), .A2(n4540), .B1(n6648), .B2(data_in[0]), 
        .ZN(n4539) );
  INV_X1 U4419 ( .A(n4541), .ZN(n4867) );
  AOI22_X1 U4420 ( .A1(\mem[220][1] ), .A2(n4540), .B1(n6648), .B2(data_in[1]), 
        .ZN(n4541) );
  INV_X1 U4421 ( .A(n4542), .ZN(n4866) );
  AOI22_X1 U4422 ( .A1(\mem[220][2] ), .A2(n4540), .B1(n6648), .B2(data_in[2]), 
        .ZN(n4542) );
  INV_X1 U4423 ( .A(n4543), .ZN(n4865) );
  AOI22_X1 U4424 ( .A1(\mem[220][3] ), .A2(n4540), .B1(n6648), .B2(data_in[3]), 
        .ZN(n4543) );
  INV_X1 U4425 ( .A(n4544), .ZN(n4864) );
  AOI22_X1 U4426 ( .A1(\mem[220][4] ), .A2(n4540), .B1(n6648), .B2(data_in[4]), 
        .ZN(n4544) );
  INV_X1 U4427 ( .A(n4545), .ZN(n4863) );
  AOI22_X1 U4428 ( .A1(\mem[220][5] ), .A2(n4540), .B1(n6648), .B2(data_in[5]), 
        .ZN(n4545) );
  INV_X1 U4429 ( .A(n4546), .ZN(n4862) );
  AOI22_X1 U4430 ( .A1(\mem[220][6] ), .A2(n4540), .B1(n6648), .B2(data_in[6]), 
        .ZN(n4546) );
  INV_X1 U4431 ( .A(n4547), .ZN(n4861) );
  AOI22_X1 U4432 ( .A1(\mem[220][7] ), .A2(n4540), .B1(n6648), .B2(data_in[7]), 
        .ZN(n4547) );
  INV_X1 U4433 ( .A(n4550), .ZN(n4860) );
  AOI22_X1 U4434 ( .A1(\mem[221][0] ), .A2(n4551), .B1(n6647), .B2(data_in[0]), 
        .ZN(n4550) );
  INV_X1 U4435 ( .A(n4552), .ZN(n4859) );
  AOI22_X1 U4436 ( .A1(\mem[221][1] ), .A2(n4551), .B1(n6647), .B2(data_in[1]), 
        .ZN(n4552) );
  INV_X1 U4437 ( .A(n4553), .ZN(n4858) );
  AOI22_X1 U4438 ( .A1(\mem[221][2] ), .A2(n4551), .B1(n6647), .B2(data_in[2]), 
        .ZN(n4553) );
  INV_X1 U4439 ( .A(n4554), .ZN(n4857) );
  AOI22_X1 U4440 ( .A1(\mem[221][3] ), .A2(n4551), .B1(n6647), .B2(data_in[3]), 
        .ZN(n4554) );
  INV_X1 U4441 ( .A(n4555), .ZN(n4856) );
  AOI22_X1 U4442 ( .A1(\mem[221][4] ), .A2(n4551), .B1(n6647), .B2(data_in[4]), 
        .ZN(n4555) );
  INV_X1 U4443 ( .A(n4556), .ZN(n4855) );
  AOI22_X1 U4444 ( .A1(\mem[221][5] ), .A2(n4551), .B1(n6647), .B2(data_in[5]), 
        .ZN(n4556) );
  INV_X1 U4445 ( .A(n4557), .ZN(n4854) );
  AOI22_X1 U4446 ( .A1(\mem[221][6] ), .A2(n4551), .B1(n6647), .B2(data_in[6]), 
        .ZN(n4557) );
  INV_X1 U4447 ( .A(n4558), .ZN(n4853) );
  AOI22_X1 U4448 ( .A1(\mem[221][7] ), .A2(n4551), .B1(n6647), .B2(data_in[7]), 
        .ZN(n4558) );
  INV_X1 U4449 ( .A(n4560), .ZN(n4852) );
  AOI22_X1 U4450 ( .A1(\mem[222][0] ), .A2(n4561), .B1(n6646), .B2(data_in[0]), 
        .ZN(n4560) );
  INV_X1 U4451 ( .A(n4562), .ZN(n4851) );
  AOI22_X1 U4452 ( .A1(\mem[222][1] ), .A2(n4561), .B1(n6646), .B2(data_in[1]), 
        .ZN(n4562) );
  INV_X1 U4453 ( .A(n4563), .ZN(n4850) );
  AOI22_X1 U4454 ( .A1(\mem[222][2] ), .A2(n4561), .B1(n6646), .B2(data_in[2]), 
        .ZN(n4563) );
  INV_X1 U4455 ( .A(n4564), .ZN(n4849) );
  AOI22_X1 U4456 ( .A1(\mem[222][3] ), .A2(n4561), .B1(n6646), .B2(data_in[3]), 
        .ZN(n4564) );
  INV_X1 U4457 ( .A(n4565), .ZN(n4848) );
  AOI22_X1 U4458 ( .A1(\mem[222][4] ), .A2(n4561), .B1(n6646), .B2(data_in[4]), 
        .ZN(n4565) );
  INV_X1 U4459 ( .A(n4566), .ZN(n4847) );
  AOI22_X1 U4460 ( .A1(\mem[222][5] ), .A2(n4561), .B1(n6646), .B2(data_in[5]), 
        .ZN(n4566) );
  INV_X1 U4461 ( .A(n4567), .ZN(n4846) );
  AOI22_X1 U4462 ( .A1(\mem[222][6] ), .A2(n4561), .B1(n6646), .B2(data_in[6]), 
        .ZN(n4567) );
  INV_X1 U4463 ( .A(n4568), .ZN(n4845) );
  AOI22_X1 U4464 ( .A1(\mem[222][7] ), .A2(n4561), .B1(n6646), .B2(data_in[7]), 
        .ZN(n4568) );
  INV_X1 U4465 ( .A(n4569), .ZN(n4844) );
  AOI22_X1 U4466 ( .A1(\mem[223][0] ), .A2(n4570), .B1(n6645), .B2(data_in[0]), 
        .ZN(n4569) );
  INV_X1 U4467 ( .A(n4571), .ZN(n4843) );
  AOI22_X1 U4468 ( .A1(\mem[223][1] ), .A2(n4570), .B1(n6645), .B2(data_in[1]), 
        .ZN(n4571) );
  INV_X1 U4469 ( .A(n4572), .ZN(n4842) );
  AOI22_X1 U4470 ( .A1(\mem[223][2] ), .A2(n4570), .B1(n6645), .B2(data_in[2]), 
        .ZN(n4572) );
  INV_X1 U4471 ( .A(n4573), .ZN(n4841) );
  AOI22_X1 U4472 ( .A1(\mem[223][3] ), .A2(n4570), .B1(n6645), .B2(data_in[3]), 
        .ZN(n4573) );
  INV_X1 U4473 ( .A(n4574), .ZN(n4840) );
  AOI22_X1 U4474 ( .A1(\mem[223][4] ), .A2(n4570), .B1(n6645), .B2(data_in[4]), 
        .ZN(n4574) );
  INV_X1 U4475 ( .A(n4575), .ZN(n4839) );
  AOI22_X1 U4476 ( .A1(\mem[223][5] ), .A2(n4570), .B1(n6645), .B2(data_in[5]), 
        .ZN(n4575) );
  INV_X1 U4477 ( .A(n4576), .ZN(n4838) );
  AOI22_X1 U4478 ( .A1(\mem[223][6] ), .A2(n4570), .B1(n6645), .B2(data_in[6]), 
        .ZN(n4576) );
  INV_X1 U4479 ( .A(n4577), .ZN(n4837) );
  AOI22_X1 U4480 ( .A1(\mem[223][7] ), .A2(n4570), .B1(n6645), .B2(data_in[7]), 
        .ZN(n4577) );
  INV_X1 U4481 ( .A(n4578), .ZN(n4836) );
  AOI22_X1 U4482 ( .A1(\mem[224][0] ), .A2(n4579), .B1(n6638), .B2(data_in[0]), 
        .ZN(n4578) );
  INV_X1 U4483 ( .A(n4580), .ZN(n4835) );
  AOI22_X1 U4484 ( .A1(\mem[224][1] ), .A2(n4579), .B1(n6638), .B2(data_in[1]), 
        .ZN(n4580) );
  INV_X1 U4485 ( .A(n4581), .ZN(n4834) );
  AOI22_X1 U4486 ( .A1(\mem[224][2] ), .A2(n4579), .B1(n6638), .B2(data_in[2]), 
        .ZN(n4581) );
  INV_X1 U4487 ( .A(n4582), .ZN(n4833) );
  AOI22_X1 U4488 ( .A1(\mem[224][3] ), .A2(n4579), .B1(n6638), .B2(data_in[3]), 
        .ZN(n4582) );
  INV_X1 U4489 ( .A(n4583), .ZN(n4832) );
  AOI22_X1 U4490 ( .A1(\mem[224][4] ), .A2(n4579), .B1(n6638), .B2(data_in[4]), 
        .ZN(n4583) );
  INV_X1 U4491 ( .A(n4584), .ZN(n4831) );
  AOI22_X1 U4492 ( .A1(\mem[224][5] ), .A2(n4579), .B1(n6638), .B2(data_in[5]), 
        .ZN(n4584) );
  INV_X1 U4493 ( .A(n4585), .ZN(n4830) );
  AOI22_X1 U4494 ( .A1(\mem[224][6] ), .A2(n4579), .B1(n6638), .B2(data_in[6]), 
        .ZN(n4585) );
  INV_X1 U4495 ( .A(n4586), .ZN(n4829) );
  AOI22_X1 U4496 ( .A1(\mem[224][7] ), .A2(n4579), .B1(n6638), .B2(data_in[7]), 
        .ZN(n4586) );
  INV_X1 U4497 ( .A(n4588), .ZN(n4828) );
  AOI22_X1 U4498 ( .A1(\mem[225][0] ), .A2(n4589), .B1(n6637), .B2(data_in[0]), 
        .ZN(n4588) );
  INV_X1 U4499 ( .A(n4590), .ZN(n4827) );
  AOI22_X1 U4500 ( .A1(\mem[225][1] ), .A2(n4589), .B1(n6637), .B2(data_in[1]), 
        .ZN(n4590) );
  INV_X1 U4501 ( .A(n4591), .ZN(n4826) );
  AOI22_X1 U4502 ( .A1(\mem[225][2] ), .A2(n4589), .B1(n6637), .B2(data_in[2]), 
        .ZN(n4591) );
  INV_X1 U4503 ( .A(n4592), .ZN(n4825) );
  AOI22_X1 U4504 ( .A1(\mem[225][3] ), .A2(n4589), .B1(n6637), .B2(data_in[3]), 
        .ZN(n4592) );
  INV_X1 U4505 ( .A(n4593), .ZN(n4824) );
  AOI22_X1 U4506 ( .A1(\mem[225][4] ), .A2(n4589), .B1(n6637), .B2(data_in[4]), 
        .ZN(n4593) );
  INV_X1 U4507 ( .A(n4594), .ZN(n4823) );
  AOI22_X1 U4508 ( .A1(\mem[225][5] ), .A2(n4589), .B1(n6637), .B2(data_in[5]), 
        .ZN(n4594) );
  INV_X1 U4509 ( .A(n4595), .ZN(n4822) );
  AOI22_X1 U4510 ( .A1(\mem[225][6] ), .A2(n4589), .B1(n6637), .B2(data_in[6]), 
        .ZN(n4595) );
  INV_X1 U4511 ( .A(n4596), .ZN(n4821) );
  AOI22_X1 U4512 ( .A1(\mem[225][7] ), .A2(n4589), .B1(n6637), .B2(data_in[7]), 
        .ZN(n4596) );
  INV_X1 U4513 ( .A(n4597), .ZN(n4820) );
  AOI22_X1 U4514 ( .A1(\mem[226][0] ), .A2(n4598), .B1(n6636), .B2(data_in[0]), 
        .ZN(n4597) );
  INV_X1 U4515 ( .A(n4599), .ZN(n4819) );
  AOI22_X1 U4516 ( .A1(\mem[226][1] ), .A2(n4598), .B1(n6636), .B2(data_in[1]), 
        .ZN(n4599) );
  INV_X1 U4517 ( .A(n4600), .ZN(n4818) );
  AOI22_X1 U4518 ( .A1(\mem[226][2] ), .A2(n4598), .B1(n6636), .B2(data_in[2]), 
        .ZN(n4600) );
  INV_X1 U4519 ( .A(n4601), .ZN(n4817) );
  AOI22_X1 U4520 ( .A1(\mem[226][3] ), .A2(n4598), .B1(n6636), .B2(data_in[3]), 
        .ZN(n4601) );
  INV_X1 U4521 ( .A(n4602), .ZN(n4816) );
  AOI22_X1 U4522 ( .A1(\mem[226][4] ), .A2(n4598), .B1(n6636), .B2(data_in[4]), 
        .ZN(n4602) );
  INV_X1 U4523 ( .A(n4603), .ZN(n4815) );
  AOI22_X1 U4524 ( .A1(\mem[226][5] ), .A2(n4598), .B1(n6636), .B2(data_in[5]), 
        .ZN(n4603) );
  INV_X1 U4525 ( .A(n4604), .ZN(n4814) );
  AOI22_X1 U4526 ( .A1(\mem[226][6] ), .A2(n4598), .B1(n6636), .B2(data_in[6]), 
        .ZN(n4604) );
  INV_X1 U4527 ( .A(n4605), .ZN(n4813) );
  AOI22_X1 U4528 ( .A1(\mem[226][7] ), .A2(n4598), .B1(n6636), .B2(data_in[7]), 
        .ZN(n4605) );
  INV_X1 U4529 ( .A(n4606), .ZN(n4812) );
  AOI22_X1 U4530 ( .A1(\mem[227][0] ), .A2(n4607), .B1(n6635), .B2(data_in[0]), 
        .ZN(n4606) );
  INV_X1 U4531 ( .A(n4608), .ZN(n4811) );
  AOI22_X1 U4532 ( .A1(\mem[227][1] ), .A2(n4607), .B1(n6635), .B2(data_in[1]), 
        .ZN(n4608) );
  INV_X1 U4533 ( .A(n4609), .ZN(n4810) );
  AOI22_X1 U4534 ( .A1(\mem[227][2] ), .A2(n4607), .B1(n6635), .B2(data_in[2]), 
        .ZN(n4609) );
  INV_X1 U4535 ( .A(n4610), .ZN(n4809) );
  AOI22_X1 U4536 ( .A1(\mem[227][3] ), .A2(n4607), .B1(n6635), .B2(data_in[3]), 
        .ZN(n4610) );
  INV_X1 U4537 ( .A(n4611), .ZN(n4808) );
  AOI22_X1 U4538 ( .A1(\mem[227][4] ), .A2(n4607), .B1(n6635), .B2(data_in[4]), 
        .ZN(n4611) );
  INV_X1 U4539 ( .A(n4612), .ZN(n4807) );
  AOI22_X1 U4540 ( .A1(\mem[227][5] ), .A2(n4607), .B1(n6635), .B2(data_in[5]), 
        .ZN(n4612) );
  INV_X1 U4541 ( .A(n4613), .ZN(n4806) );
  AOI22_X1 U4542 ( .A1(\mem[227][6] ), .A2(n4607), .B1(n6635), .B2(data_in[6]), 
        .ZN(n4613) );
  INV_X1 U4543 ( .A(n4614), .ZN(n4805) );
  AOI22_X1 U4544 ( .A1(\mem[227][7] ), .A2(n4607), .B1(n6635), .B2(data_in[7]), 
        .ZN(n4614) );
  INV_X1 U4545 ( .A(n4615), .ZN(n4804) );
  AOI22_X1 U4546 ( .A1(\mem[228][0] ), .A2(n4616), .B1(n6634), .B2(data_in[0]), 
        .ZN(n4615) );
  INV_X1 U4547 ( .A(n4617), .ZN(n4803) );
  AOI22_X1 U4548 ( .A1(\mem[228][1] ), .A2(n4616), .B1(n6634), .B2(data_in[1]), 
        .ZN(n4617) );
  INV_X1 U4549 ( .A(n4618), .ZN(n4802) );
  AOI22_X1 U4550 ( .A1(\mem[228][2] ), .A2(n4616), .B1(n6634), .B2(data_in[2]), 
        .ZN(n4618) );
  INV_X1 U4551 ( .A(n4619), .ZN(n4801) );
  AOI22_X1 U4552 ( .A1(\mem[228][3] ), .A2(n4616), .B1(n6634), .B2(data_in[3]), 
        .ZN(n4619) );
  INV_X1 U4553 ( .A(n4620), .ZN(n4800) );
  AOI22_X1 U4554 ( .A1(\mem[228][4] ), .A2(n4616), .B1(n6634), .B2(data_in[4]), 
        .ZN(n4620) );
  INV_X1 U4555 ( .A(n4621), .ZN(n4799) );
  AOI22_X1 U4556 ( .A1(\mem[228][5] ), .A2(n4616), .B1(n6634), .B2(data_in[5]), 
        .ZN(n4621) );
  INV_X1 U4557 ( .A(n4622), .ZN(n4798) );
  AOI22_X1 U4558 ( .A1(\mem[228][6] ), .A2(n4616), .B1(n6634), .B2(data_in[6]), 
        .ZN(n4622) );
  INV_X1 U4559 ( .A(n4623), .ZN(n4797) );
  AOI22_X1 U4560 ( .A1(\mem[228][7] ), .A2(n4616), .B1(n6634), .B2(data_in[7]), 
        .ZN(n4623) );
  INV_X1 U4561 ( .A(n4625), .ZN(n4796) );
  AOI22_X1 U4562 ( .A1(\mem[229][0] ), .A2(n4626), .B1(n6633), .B2(data_in[0]), 
        .ZN(n4625) );
  INV_X1 U4563 ( .A(n4627), .ZN(n4795) );
  AOI22_X1 U4564 ( .A1(\mem[229][1] ), .A2(n4626), .B1(n6633), .B2(data_in[1]), 
        .ZN(n4627) );
  INV_X1 U4565 ( .A(n4628), .ZN(n4794) );
  AOI22_X1 U4566 ( .A1(\mem[229][2] ), .A2(n4626), .B1(n6633), .B2(data_in[2]), 
        .ZN(n4628) );
  INV_X1 U4567 ( .A(n4629), .ZN(n4793) );
  AOI22_X1 U4568 ( .A1(\mem[229][3] ), .A2(n4626), .B1(n6633), .B2(data_in[3]), 
        .ZN(n4629) );
  INV_X1 U4569 ( .A(n4630), .ZN(n4792) );
  AOI22_X1 U4570 ( .A1(\mem[229][4] ), .A2(n4626), .B1(n6633), .B2(data_in[4]), 
        .ZN(n4630) );
  INV_X1 U4571 ( .A(n4631), .ZN(n4791) );
  AOI22_X1 U4572 ( .A1(\mem[229][5] ), .A2(n4626), .B1(n6633), .B2(data_in[5]), 
        .ZN(n4631) );
  INV_X1 U4573 ( .A(n4632), .ZN(n4790) );
  AOI22_X1 U4574 ( .A1(\mem[229][6] ), .A2(n4626), .B1(n6633), .B2(data_in[6]), 
        .ZN(n4632) );
  INV_X1 U4575 ( .A(n4633), .ZN(n4789) );
  AOI22_X1 U4576 ( .A1(\mem[229][7] ), .A2(n4626), .B1(n6633), .B2(data_in[7]), 
        .ZN(n4633) );
  INV_X1 U4577 ( .A(n4634), .ZN(n4788) );
  AOI22_X1 U4578 ( .A1(\mem[230][0] ), .A2(n4635), .B1(n6632), .B2(data_in[0]), 
        .ZN(n4634) );
  INV_X1 U4579 ( .A(n4636), .ZN(n4787) );
  AOI22_X1 U4580 ( .A1(\mem[230][1] ), .A2(n4635), .B1(n6632), .B2(data_in[1]), 
        .ZN(n4636) );
  INV_X1 U4581 ( .A(n4637), .ZN(n4786) );
  AOI22_X1 U4582 ( .A1(\mem[230][2] ), .A2(n4635), .B1(n6632), .B2(data_in[2]), 
        .ZN(n4637) );
  INV_X1 U4583 ( .A(n4638), .ZN(n4785) );
  AOI22_X1 U4584 ( .A1(\mem[230][3] ), .A2(n4635), .B1(n6632), .B2(data_in[3]), 
        .ZN(n4638) );
  INV_X1 U4585 ( .A(n4639), .ZN(n4784) );
  AOI22_X1 U4586 ( .A1(\mem[230][4] ), .A2(n4635), .B1(n6632), .B2(data_in[4]), 
        .ZN(n4639) );
  INV_X1 U4587 ( .A(n4640), .ZN(n4783) );
  AOI22_X1 U4588 ( .A1(\mem[230][5] ), .A2(n4635), .B1(n6632), .B2(data_in[5]), 
        .ZN(n4640) );
  INV_X1 U4589 ( .A(n4641), .ZN(n4782) );
  AOI22_X1 U4590 ( .A1(\mem[230][6] ), .A2(n4635), .B1(n6632), .B2(data_in[6]), 
        .ZN(n4641) );
  INV_X1 U4591 ( .A(n4642), .ZN(n4781) );
  AOI22_X1 U4592 ( .A1(\mem[230][7] ), .A2(n4635), .B1(n6632), .B2(data_in[7]), 
        .ZN(n4642) );
  INV_X1 U4593 ( .A(n4643), .ZN(n4780) );
  AOI22_X1 U4594 ( .A1(\mem[231][0] ), .A2(n4644), .B1(n6631), .B2(data_in[0]), 
        .ZN(n4643) );
  INV_X1 U4595 ( .A(n4645), .ZN(n4779) );
  AOI22_X1 U4596 ( .A1(\mem[231][1] ), .A2(n4644), .B1(n6631), .B2(data_in[1]), 
        .ZN(n4645) );
  INV_X1 U4597 ( .A(n4646), .ZN(n4778) );
  AOI22_X1 U4598 ( .A1(\mem[231][2] ), .A2(n4644), .B1(n6631), .B2(data_in[2]), 
        .ZN(n4646) );
  INV_X1 U4599 ( .A(n4647), .ZN(n4777) );
  AOI22_X1 U4600 ( .A1(\mem[231][3] ), .A2(n4644), .B1(n6631), .B2(data_in[3]), 
        .ZN(n4647) );
  INV_X1 U4601 ( .A(n4648), .ZN(n4776) );
  AOI22_X1 U4602 ( .A1(\mem[231][4] ), .A2(n4644), .B1(n6631), .B2(data_in[4]), 
        .ZN(n4648) );
  INV_X1 U4603 ( .A(n4649), .ZN(n4775) );
  AOI22_X1 U4604 ( .A1(\mem[231][5] ), .A2(n4644), .B1(n6631), .B2(data_in[5]), 
        .ZN(n4649) );
  INV_X1 U4605 ( .A(n4650), .ZN(n4774) );
  AOI22_X1 U4606 ( .A1(\mem[231][6] ), .A2(n4644), .B1(n6631), .B2(data_in[6]), 
        .ZN(n4650) );
  INV_X1 U4607 ( .A(n4651), .ZN(n4773) );
  AOI22_X1 U4608 ( .A1(\mem[231][7] ), .A2(n4644), .B1(n6631), .B2(data_in[7]), 
        .ZN(n4651) );
  INV_X1 U4609 ( .A(n4652), .ZN(n4772) );
  AOI22_X1 U4610 ( .A1(\mem[232][0] ), .A2(n4653), .B1(n6630), .B2(data_in[0]), 
        .ZN(n4652) );
  INV_X1 U4611 ( .A(n4654), .ZN(n4771) );
  AOI22_X1 U4612 ( .A1(\mem[232][1] ), .A2(n4653), .B1(n6630), .B2(data_in[1]), 
        .ZN(n4654) );
  INV_X1 U4613 ( .A(n4655), .ZN(n4770) );
  AOI22_X1 U4614 ( .A1(\mem[232][2] ), .A2(n4653), .B1(n6630), .B2(data_in[2]), 
        .ZN(n4655) );
  INV_X1 U4615 ( .A(n4656), .ZN(n4769) );
  AOI22_X1 U4616 ( .A1(\mem[232][3] ), .A2(n4653), .B1(n6630), .B2(data_in[3]), 
        .ZN(n4656) );
  INV_X1 U4617 ( .A(n4657), .ZN(n4768) );
  AOI22_X1 U4618 ( .A1(\mem[232][4] ), .A2(n4653), .B1(n6630), .B2(data_in[4]), 
        .ZN(n4657) );
  INV_X1 U4619 ( .A(n4658), .ZN(n4767) );
  AOI22_X1 U4620 ( .A1(\mem[232][5] ), .A2(n4653), .B1(n6630), .B2(data_in[5]), 
        .ZN(n4658) );
  INV_X1 U4621 ( .A(n4659), .ZN(n4766) );
  AOI22_X1 U4622 ( .A1(\mem[232][6] ), .A2(n4653), .B1(n6630), .B2(data_in[6]), 
        .ZN(n4659) );
  INV_X1 U4623 ( .A(n4660), .ZN(n4765) );
  AOI22_X1 U4624 ( .A1(\mem[232][7] ), .A2(n4653), .B1(n6630), .B2(data_in[7]), 
        .ZN(n4660) );
  INV_X1 U4625 ( .A(n2329), .ZN(n4748) );
  AOI22_X1 U4626 ( .A1(\mem[235][0] ), .A2(n2330), .B1(n6643), .B2(data_in[0]), 
        .ZN(n2329) );
  INV_X1 U4627 ( .A(n2331), .ZN(n4747) );
  AOI22_X1 U4628 ( .A1(\mem[235][1] ), .A2(n2330), .B1(n6643), .B2(data_in[1]), 
        .ZN(n2331) );
  INV_X1 U4629 ( .A(n2332), .ZN(n4746) );
  AOI22_X1 U4630 ( .A1(\mem[235][2] ), .A2(n2330), .B1(n6643), .B2(data_in[2]), 
        .ZN(n2332) );
  INV_X1 U4631 ( .A(n2333), .ZN(n4745) );
  AOI22_X1 U4632 ( .A1(\mem[235][3] ), .A2(n2330), .B1(n6643), .B2(data_in[3]), 
        .ZN(n2333) );
  INV_X1 U4633 ( .A(n2334), .ZN(n4744) );
  AOI22_X1 U4634 ( .A1(\mem[235][4] ), .A2(n2330), .B1(n6643), .B2(data_in[4]), 
        .ZN(n2334) );
  INV_X1 U4635 ( .A(n2335), .ZN(n4743) );
  AOI22_X1 U4636 ( .A1(\mem[235][5] ), .A2(n2330), .B1(n6643), .B2(data_in[5]), 
        .ZN(n2335) );
  INV_X1 U4637 ( .A(n2336), .ZN(n4742) );
  AOI22_X1 U4638 ( .A1(\mem[235][6] ), .A2(n2330), .B1(n6643), .B2(data_in[6]), 
        .ZN(n2336) );
  INV_X1 U4639 ( .A(n2337), .ZN(n4741) );
  AOI22_X1 U4640 ( .A1(\mem[235][7] ), .A2(n2330), .B1(n6643), .B2(data_in[7]), 
        .ZN(n2337) );
  INV_X1 U4641 ( .A(n2339), .ZN(n4740) );
  AOI22_X1 U4642 ( .A1(\mem[236][0] ), .A2(n2340), .B1(n6642), .B2(data_in[0]), 
        .ZN(n2339) );
  INV_X1 U4643 ( .A(n2341), .ZN(n4739) );
  AOI22_X1 U4644 ( .A1(\mem[236][1] ), .A2(n2340), .B1(n6642), .B2(data_in[1]), 
        .ZN(n2341) );
  INV_X1 U4645 ( .A(n2342), .ZN(n4738) );
  AOI22_X1 U4646 ( .A1(\mem[236][2] ), .A2(n2340), .B1(n6642), .B2(data_in[2]), 
        .ZN(n2342) );
  INV_X1 U4647 ( .A(n2343), .ZN(n4737) );
  AOI22_X1 U4648 ( .A1(\mem[236][3] ), .A2(n2340), .B1(n6642), .B2(data_in[3]), 
        .ZN(n2343) );
  INV_X1 U4649 ( .A(n2344), .ZN(n4736) );
  AOI22_X1 U4650 ( .A1(\mem[236][4] ), .A2(n2340), .B1(n6642), .B2(data_in[4]), 
        .ZN(n2344) );
  INV_X1 U4651 ( .A(n2345), .ZN(n4735) );
  AOI22_X1 U4652 ( .A1(\mem[236][5] ), .A2(n2340), .B1(n6642), .B2(data_in[5]), 
        .ZN(n2345) );
  INV_X1 U4653 ( .A(n2346), .ZN(n4734) );
  AOI22_X1 U4654 ( .A1(\mem[236][6] ), .A2(n2340), .B1(n6642), .B2(data_in[6]), 
        .ZN(n2346) );
  INV_X1 U4655 ( .A(n2347), .ZN(n4733) );
  AOI22_X1 U4656 ( .A1(\mem[236][7] ), .A2(n2340), .B1(n6642), .B2(data_in[7]), 
        .ZN(n2347) );
  INV_X1 U4657 ( .A(n2349), .ZN(n4732) );
  AOI22_X1 U4658 ( .A1(\mem[237][0] ), .A2(n2350), .B1(n6641), .B2(data_in[0]), 
        .ZN(n2349) );
  INV_X1 U4659 ( .A(n2351), .ZN(n4731) );
  AOI22_X1 U4660 ( .A1(\mem[237][1] ), .A2(n2350), .B1(n6641), .B2(data_in[1]), 
        .ZN(n2351) );
  INV_X1 U4661 ( .A(n2352), .ZN(n4730) );
  AOI22_X1 U4662 ( .A1(\mem[237][2] ), .A2(n2350), .B1(n6641), .B2(data_in[2]), 
        .ZN(n2352) );
  INV_X1 U4663 ( .A(n2353), .ZN(n4729) );
  AOI22_X1 U4664 ( .A1(\mem[237][3] ), .A2(n2350), .B1(n6641), .B2(data_in[3]), 
        .ZN(n2353) );
  INV_X1 U4665 ( .A(n2354), .ZN(n4728) );
  AOI22_X1 U4666 ( .A1(\mem[237][4] ), .A2(n2350), .B1(n6641), .B2(data_in[4]), 
        .ZN(n2354) );
  INV_X1 U4667 ( .A(n2355), .ZN(n4727) );
  AOI22_X1 U4668 ( .A1(\mem[237][5] ), .A2(n2350), .B1(n6641), .B2(data_in[5]), 
        .ZN(n2355) );
  INV_X1 U4669 ( .A(n2356), .ZN(n4726) );
  AOI22_X1 U4670 ( .A1(\mem[237][6] ), .A2(n2350), .B1(n6641), .B2(data_in[6]), 
        .ZN(n2356) );
  INV_X1 U4671 ( .A(n2357), .ZN(n4725) );
  AOI22_X1 U4672 ( .A1(\mem[237][7] ), .A2(n2350), .B1(n6641), .B2(data_in[7]), 
        .ZN(n2357) );
  INV_X1 U4673 ( .A(n2359), .ZN(n4724) );
  AOI22_X1 U4674 ( .A1(\mem[238][0] ), .A2(n2360), .B1(n6640), .B2(data_in[0]), 
        .ZN(n2359) );
  INV_X1 U4675 ( .A(n2361), .ZN(n4723) );
  AOI22_X1 U4676 ( .A1(\mem[238][1] ), .A2(n2360), .B1(n6640), .B2(data_in[1]), 
        .ZN(n2361) );
  INV_X1 U4677 ( .A(n2362), .ZN(n4722) );
  AOI22_X1 U4678 ( .A1(\mem[238][2] ), .A2(n2360), .B1(n6640), .B2(data_in[2]), 
        .ZN(n2362) );
  INV_X1 U4679 ( .A(n2363), .ZN(n4721) );
  AOI22_X1 U4680 ( .A1(\mem[238][3] ), .A2(n2360), .B1(n6640), .B2(data_in[3]), 
        .ZN(n2363) );
  INV_X1 U4681 ( .A(n2364), .ZN(n4720) );
  AOI22_X1 U4682 ( .A1(\mem[238][4] ), .A2(n2360), .B1(n6640), .B2(data_in[4]), 
        .ZN(n2364) );
  INV_X1 U4683 ( .A(n2365), .ZN(n4719) );
  AOI22_X1 U4684 ( .A1(\mem[238][5] ), .A2(n2360), .B1(n6640), .B2(data_in[5]), 
        .ZN(n2365) );
  INV_X1 U4685 ( .A(n2366), .ZN(n4718) );
  AOI22_X1 U4686 ( .A1(\mem[238][6] ), .A2(n2360), .B1(n6640), .B2(data_in[6]), 
        .ZN(n2366) );
  INV_X1 U4687 ( .A(n2367), .ZN(n4717) );
  AOI22_X1 U4688 ( .A1(\mem[238][7] ), .A2(n2360), .B1(n6640), .B2(data_in[7]), 
        .ZN(n2367) );
  INV_X1 U4689 ( .A(n2369), .ZN(n4716) );
  AOI22_X1 U4690 ( .A1(\mem[239][0] ), .A2(n2370), .B1(n6639), .B2(data_in[0]), 
        .ZN(n2369) );
  INV_X1 U4691 ( .A(n2371), .ZN(n4715) );
  AOI22_X1 U4692 ( .A1(\mem[239][1] ), .A2(n2370), .B1(n6639), .B2(data_in[1]), 
        .ZN(n2371) );
  INV_X1 U4693 ( .A(n2372), .ZN(n4714) );
  AOI22_X1 U4694 ( .A1(\mem[239][2] ), .A2(n2370), .B1(n6639), .B2(data_in[2]), 
        .ZN(n2372) );
  INV_X1 U4695 ( .A(n2373), .ZN(n4713) );
  AOI22_X1 U4696 ( .A1(\mem[239][3] ), .A2(n2370), .B1(n6639), .B2(data_in[3]), 
        .ZN(n2373) );
  INV_X1 U4697 ( .A(n2374), .ZN(n4712) );
  AOI22_X1 U4698 ( .A1(\mem[239][4] ), .A2(n2370), .B1(n6639), .B2(data_in[4]), 
        .ZN(n2374) );
  INV_X1 U4699 ( .A(n2375), .ZN(n4711) );
  AOI22_X1 U4700 ( .A1(\mem[239][5] ), .A2(n2370), .B1(n6639), .B2(data_in[5]), 
        .ZN(n2375) );
  INV_X1 U4701 ( .A(n2376), .ZN(n4710) );
  AOI22_X1 U4702 ( .A1(\mem[239][6] ), .A2(n2370), .B1(n6639), .B2(data_in[6]), 
        .ZN(n2376) );
  INV_X1 U4703 ( .A(n2377), .ZN(n4709) );
  AOI22_X1 U4704 ( .A1(\mem[239][7] ), .A2(n2370), .B1(n6639), .B2(data_in[7]), 
        .ZN(n2377) );
  INV_X1 U4705 ( .A(n2379), .ZN(n4708) );
  AOI22_X1 U4706 ( .A1(\mem[240][0] ), .A2(n2380), .B1(n6884), .B2(data_in[0]), 
        .ZN(n2379) );
  INV_X1 U4707 ( .A(n2381), .ZN(n4707) );
  AOI22_X1 U4708 ( .A1(\mem[240][1] ), .A2(n2380), .B1(n6884), .B2(data_in[1]), 
        .ZN(n2381) );
  INV_X1 U4709 ( .A(n2382), .ZN(n4706) );
  AOI22_X1 U4710 ( .A1(\mem[240][2] ), .A2(n2380), .B1(n6884), .B2(data_in[2]), 
        .ZN(n2382) );
  INV_X1 U4711 ( .A(n2383), .ZN(n4705) );
  AOI22_X1 U4712 ( .A1(\mem[240][3] ), .A2(n2380), .B1(n6884), .B2(data_in[3]), 
        .ZN(n2383) );
  INV_X1 U4713 ( .A(n2384), .ZN(n4704) );
  AOI22_X1 U4714 ( .A1(\mem[240][4] ), .A2(n2380), .B1(n6884), .B2(data_in[4]), 
        .ZN(n2384) );
  INV_X1 U4715 ( .A(n2385), .ZN(n4703) );
  AOI22_X1 U4716 ( .A1(\mem[240][5] ), .A2(n2380), .B1(n6884), .B2(data_in[5]), 
        .ZN(n2385) );
  INV_X1 U4717 ( .A(n2386), .ZN(n4702) );
  AOI22_X1 U4718 ( .A1(\mem[240][6] ), .A2(n2380), .B1(n6884), .B2(data_in[6]), 
        .ZN(n2386) );
  INV_X1 U4719 ( .A(n2387), .ZN(n4701) );
  AOI22_X1 U4720 ( .A1(\mem[240][7] ), .A2(n2380), .B1(n6884), .B2(data_in[7]), 
        .ZN(n2387) );
  INV_X1 U4721 ( .A(n2390), .ZN(n4700) );
  AOI22_X1 U4722 ( .A1(\mem[241][0] ), .A2(n2391), .B1(n6883), .B2(data_in[0]), 
        .ZN(n2390) );
  INV_X1 U4723 ( .A(n2392), .ZN(n4699) );
  AOI22_X1 U4724 ( .A1(\mem[241][1] ), .A2(n2391), .B1(n6883), .B2(data_in[1]), 
        .ZN(n2392) );
  INV_X1 U4725 ( .A(n2393), .ZN(n4698) );
  AOI22_X1 U4726 ( .A1(\mem[241][2] ), .A2(n2391), .B1(n6883), .B2(data_in[2]), 
        .ZN(n2393) );
  INV_X1 U4727 ( .A(n2394), .ZN(n4697) );
  AOI22_X1 U4728 ( .A1(\mem[241][3] ), .A2(n2391), .B1(n6883), .B2(data_in[3]), 
        .ZN(n2394) );
  INV_X1 U4729 ( .A(n2395), .ZN(n4696) );
  AOI22_X1 U4730 ( .A1(\mem[241][4] ), .A2(n2391), .B1(n6883), .B2(data_in[4]), 
        .ZN(n2395) );
  INV_X1 U4731 ( .A(n2396), .ZN(n4695) );
  AOI22_X1 U4732 ( .A1(\mem[241][5] ), .A2(n2391), .B1(n6883), .B2(data_in[5]), 
        .ZN(n2396) );
  INV_X1 U4733 ( .A(n2397), .ZN(n4694) );
  AOI22_X1 U4734 ( .A1(\mem[241][6] ), .A2(n2391), .B1(n6883), .B2(data_in[6]), 
        .ZN(n2397) );
  INV_X1 U4735 ( .A(n2398), .ZN(n4693) );
  AOI22_X1 U4736 ( .A1(\mem[241][7] ), .A2(n2391), .B1(n6883), .B2(data_in[7]), 
        .ZN(n2398) );
  INV_X1 U4737 ( .A(n2400), .ZN(n4692) );
  AOI22_X1 U4738 ( .A1(\mem[242][0] ), .A2(n2401), .B1(n6882), .B2(data_in[0]), 
        .ZN(n2400) );
  INV_X1 U4739 ( .A(n2402), .ZN(n4691) );
  AOI22_X1 U4740 ( .A1(\mem[242][1] ), .A2(n2401), .B1(n6882), .B2(data_in[1]), 
        .ZN(n2402) );
  INV_X1 U4741 ( .A(n2403), .ZN(n4690) );
  AOI22_X1 U4742 ( .A1(\mem[242][2] ), .A2(n2401), .B1(n6882), .B2(data_in[2]), 
        .ZN(n2403) );
  INV_X1 U4743 ( .A(n2404), .ZN(n4689) );
  AOI22_X1 U4744 ( .A1(\mem[242][3] ), .A2(n2401), .B1(n6882), .B2(data_in[3]), 
        .ZN(n2404) );
  INV_X1 U4745 ( .A(n2405), .ZN(n4688) );
  AOI22_X1 U4746 ( .A1(\mem[242][4] ), .A2(n2401), .B1(n6882), .B2(data_in[4]), 
        .ZN(n2405) );
  INV_X1 U4747 ( .A(n2406), .ZN(n4687) );
  AOI22_X1 U4748 ( .A1(\mem[242][5] ), .A2(n2401), .B1(n6882), .B2(data_in[5]), 
        .ZN(n2406) );
  INV_X1 U4749 ( .A(n2407), .ZN(n4686) );
  AOI22_X1 U4750 ( .A1(\mem[242][6] ), .A2(n2401), .B1(n6882), .B2(data_in[6]), 
        .ZN(n2407) );
  INV_X1 U4751 ( .A(n2408), .ZN(n4685) );
  AOI22_X1 U4752 ( .A1(\mem[242][7] ), .A2(n2401), .B1(n6882), .B2(data_in[7]), 
        .ZN(n2408) );
  INV_X1 U4753 ( .A(n2410), .ZN(n4684) );
  AOI22_X1 U4754 ( .A1(\mem[243][0] ), .A2(n2411), .B1(n6881), .B2(data_in[0]), 
        .ZN(n2410) );
  INV_X1 U4755 ( .A(n2412), .ZN(n4683) );
  AOI22_X1 U4756 ( .A1(\mem[243][1] ), .A2(n2411), .B1(n6881), .B2(data_in[1]), 
        .ZN(n2412) );
  INV_X1 U4757 ( .A(n2413), .ZN(n4682) );
  AOI22_X1 U4758 ( .A1(\mem[243][2] ), .A2(n2411), .B1(n6881), .B2(data_in[2]), 
        .ZN(n2413) );
  INV_X1 U4759 ( .A(n2414), .ZN(n4681) );
  AOI22_X1 U4760 ( .A1(\mem[243][3] ), .A2(n2411), .B1(n6881), .B2(data_in[3]), 
        .ZN(n2414) );
  INV_X1 U4761 ( .A(n2415), .ZN(n4680) );
  AOI22_X1 U4762 ( .A1(\mem[243][4] ), .A2(n2411), .B1(n6881), .B2(data_in[4]), 
        .ZN(n2415) );
  INV_X1 U4763 ( .A(n2416), .ZN(n4679) );
  AOI22_X1 U4764 ( .A1(\mem[243][5] ), .A2(n2411), .B1(n6881), .B2(data_in[5]), 
        .ZN(n2416) );
  INV_X1 U4765 ( .A(n2417), .ZN(n4678) );
  AOI22_X1 U4766 ( .A1(\mem[243][6] ), .A2(n2411), .B1(n6881), .B2(data_in[6]), 
        .ZN(n2417) );
  INV_X1 U4767 ( .A(n2418), .ZN(n4677) );
  AOI22_X1 U4768 ( .A1(\mem[243][7] ), .A2(n2411), .B1(n6881), .B2(data_in[7]), 
        .ZN(n2418) );
  INV_X1 U4769 ( .A(n2420), .ZN(n4676) );
  AOI22_X1 U4770 ( .A1(\mem[244][0] ), .A2(n2421), .B1(n6880), .B2(data_in[0]), 
        .ZN(n2420) );
  INV_X1 U4771 ( .A(n2422), .ZN(n4675) );
  AOI22_X1 U4772 ( .A1(\mem[244][1] ), .A2(n2421), .B1(n6880), .B2(data_in[1]), 
        .ZN(n2422) );
  INV_X1 U4773 ( .A(n2423), .ZN(n4674) );
  AOI22_X1 U4774 ( .A1(\mem[244][2] ), .A2(n2421), .B1(n6880), .B2(data_in[2]), 
        .ZN(n2423) );
  INV_X1 U4775 ( .A(n2424), .ZN(n4673) );
  AOI22_X1 U4776 ( .A1(\mem[244][3] ), .A2(n2421), .B1(n6880), .B2(data_in[3]), 
        .ZN(n2424) );
  INV_X1 U4777 ( .A(n2425), .ZN(n4672) );
  AOI22_X1 U4778 ( .A1(\mem[244][4] ), .A2(n2421), .B1(n6880), .B2(data_in[4]), 
        .ZN(n2425) );
  INV_X1 U4779 ( .A(n2426), .ZN(n4671) );
  AOI22_X1 U4780 ( .A1(\mem[244][5] ), .A2(n2421), .B1(n6880), .B2(data_in[5]), 
        .ZN(n2426) );
  INV_X1 U4781 ( .A(n2427), .ZN(n4670) );
  AOI22_X1 U4782 ( .A1(\mem[244][6] ), .A2(n2421), .B1(n6880), .B2(data_in[6]), 
        .ZN(n2427) );
  INV_X1 U4783 ( .A(n2428), .ZN(n4669) );
  AOI22_X1 U4784 ( .A1(\mem[244][7] ), .A2(n2421), .B1(n6880), .B2(data_in[7]), 
        .ZN(n2428) );
  INV_X1 U4785 ( .A(n2430), .ZN(n4668) );
  AOI22_X1 U4786 ( .A1(\mem[245][0] ), .A2(n2431), .B1(n6879), .B2(data_in[0]), 
        .ZN(n2430) );
  INV_X1 U4787 ( .A(n2432), .ZN(n4667) );
  AOI22_X1 U4788 ( .A1(\mem[245][1] ), .A2(n2431), .B1(n6879), .B2(data_in[1]), 
        .ZN(n2432) );
  INV_X1 U4789 ( .A(n2433), .ZN(n4666) );
  AOI22_X1 U4790 ( .A1(\mem[245][2] ), .A2(n2431), .B1(n6879), .B2(data_in[2]), 
        .ZN(n2433) );
  INV_X1 U4791 ( .A(n2434), .ZN(n4665) );
  AOI22_X1 U4792 ( .A1(\mem[245][3] ), .A2(n2431), .B1(n6879), .B2(data_in[3]), 
        .ZN(n2434) );
  INV_X1 U4793 ( .A(n2435), .ZN(n2312) );
  AOI22_X1 U4794 ( .A1(\mem[245][4] ), .A2(n2431), .B1(n6879), .B2(data_in[4]), 
        .ZN(n2435) );
  INV_X1 U4795 ( .A(n2436), .ZN(n2311) );
  AOI22_X1 U4796 ( .A1(\mem[245][5] ), .A2(n2431), .B1(n6879), .B2(data_in[5]), 
        .ZN(n2436) );
  INV_X1 U4797 ( .A(n2437), .ZN(n2310) );
  AOI22_X1 U4798 ( .A1(\mem[245][6] ), .A2(n2431), .B1(n6879), .B2(data_in[6]), 
        .ZN(n2437) );
  INV_X1 U4799 ( .A(n2438), .ZN(n2309) );
  AOI22_X1 U4800 ( .A1(\mem[245][7] ), .A2(n2431), .B1(n6879), .B2(data_in[7]), 
        .ZN(n2438) );
  INV_X1 U4801 ( .A(n2440), .ZN(n2308) );
  AOI22_X1 U4802 ( .A1(\mem[246][0] ), .A2(n2441), .B1(n6878), .B2(data_in[0]), 
        .ZN(n2440) );
  INV_X1 U4803 ( .A(n2442), .ZN(n2307) );
  AOI22_X1 U4804 ( .A1(\mem[246][1] ), .A2(n2441), .B1(n6878), .B2(data_in[1]), 
        .ZN(n2442) );
  INV_X1 U4805 ( .A(n2443), .ZN(n2306) );
  AOI22_X1 U4806 ( .A1(\mem[246][2] ), .A2(n2441), .B1(n6878), .B2(data_in[2]), 
        .ZN(n2443) );
  INV_X1 U4807 ( .A(n2444), .ZN(n2305) );
  AOI22_X1 U4808 ( .A1(\mem[246][3] ), .A2(n2441), .B1(n6878), .B2(data_in[3]), 
        .ZN(n2444) );
  INV_X1 U4809 ( .A(n2445), .ZN(n2304) );
  AOI22_X1 U4810 ( .A1(\mem[246][4] ), .A2(n2441), .B1(n6878), .B2(data_in[4]), 
        .ZN(n2445) );
  INV_X1 U4811 ( .A(n2446), .ZN(n2303) );
  AOI22_X1 U4812 ( .A1(\mem[246][5] ), .A2(n2441), .B1(n6878), .B2(data_in[5]), 
        .ZN(n2446) );
  INV_X1 U4813 ( .A(n2447), .ZN(n2302) );
  AOI22_X1 U4814 ( .A1(\mem[246][6] ), .A2(n2441), .B1(n6878), .B2(data_in[6]), 
        .ZN(n2447) );
  INV_X1 U4815 ( .A(n2448), .ZN(n2301) );
  AOI22_X1 U4816 ( .A1(\mem[246][7] ), .A2(n2441), .B1(n6878), .B2(data_in[7]), 
        .ZN(n2448) );
  INV_X1 U4817 ( .A(n2450), .ZN(n2300) );
  AOI22_X1 U4818 ( .A1(\mem[247][0] ), .A2(n2451), .B1(n6877), .B2(data_in[0]), 
        .ZN(n2450) );
  INV_X1 U4819 ( .A(n2452), .ZN(n2299) );
  AOI22_X1 U4820 ( .A1(\mem[247][1] ), .A2(n2451), .B1(n6877), .B2(data_in[1]), 
        .ZN(n2452) );
  INV_X1 U4821 ( .A(n2453), .ZN(n2298) );
  AOI22_X1 U4822 ( .A1(\mem[247][2] ), .A2(n2451), .B1(n6877), .B2(data_in[2]), 
        .ZN(n2453) );
  INV_X1 U4823 ( .A(n2454), .ZN(n2297) );
  AOI22_X1 U4824 ( .A1(\mem[247][3] ), .A2(n2451), .B1(n6877), .B2(data_in[3]), 
        .ZN(n2454) );
  INV_X1 U4825 ( .A(n2455), .ZN(n2296) );
  AOI22_X1 U4826 ( .A1(\mem[247][4] ), .A2(n2451), .B1(n6877), .B2(data_in[4]), 
        .ZN(n2455) );
  INV_X1 U4827 ( .A(n2456), .ZN(n2295) );
  AOI22_X1 U4828 ( .A1(\mem[247][5] ), .A2(n2451), .B1(n6877), .B2(data_in[5]), 
        .ZN(n2456) );
  INV_X1 U4829 ( .A(n2457), .ZN(n2294) );
  AOI22_X1 U4830 ( .A1(\mem[247][6] ), .A2(n2451), .B1(n6877), .B2(data_in[6]), 
        .ZN(n2457) );
  INV_X1 U4831 ( .A(n2458), .ZN(n2293) );
  AOI22_X1 U4832 ( .A1(\mem[247][7] ), .A2(n2451), .B1(n6877), .B2(data_in[7]), 
        .ZN(n2458) );
  INV_X1 U4833 ( .A(n2460), .ZN(n2292) );
  AOI22_X1 U4834 ( .A1(\mem[248][0] ), .A2(n2461), .B1(n6876), .B2(data_in[0]), 
        .ZN(n2460) );
  INV_X1 U4835 ( .A(n2462), .ZN(n2291) );
  AOI22_X1 U4836 ( .A1(\mem[248][1] ), .A2(n2461), .B1(n6876), .B2(data_in[1]), 
        .ZN(n2462) );
  INV_X1 U4837 ( .A(n2463), .ZN(n2290) );
  AOI22_X1 U4838 ( .A1(\mem[248][2] ), .A2(n2461), .B1(n6876), .B2(data_in[2]), 
        .ZN(n2463) );
  INV_X1 U4839 ( .A(n2464), .ZN(n2289) );
  AOI22_X1 U4840 ( .A1(\mem[248][3] ), .A2(n2461), .B1(n6876), .B2(data_in[3]), 
        .ZN(n2464) );
  INV_X1 U4841 ( .A(n2465), .ZN(n2288) );
  AOI22_X1 U4842 ( .A1(\mem[248][4] ), .A2(n2461), .B1(n6876), .B2(data_in[4]), 
        .ZN(n2465) );
  INV_X1 U4843 ( .A(n2466), .ZN(n2287) );
  AOI22_X1 U4844 ( .A1(\mem[248][5] ), .A2(n2461), .B1(n6876), .B2(data_in[5]), 
        .ZN(n2466) );
  INV_X1 U4845 ( .A(n2467), .ZN(n2286) );
  AOI22_X1 U4846 ( .A1(\mem[248][6] ), .A2(n2461), .B1(n6876), .B2(data_in[6]), 
        .ZN(n2467) );
  INV_X1 U4847 ( .A(n2468), .ZN(n2285) );
  AOI22_X1 U4848 ( .A1(\mem[248][7] ), .A2(n2461), .B1(n6876), .B2(data_in[7]), 
        .ZN(n2468) );
  MUX2_X1 U4849 ( .A(\mem[254][0] ), .B(\mem[255][0] ), .S(n2165), .Z(n16) );
  MUX2_X1 U4850 ( .A(\mem[252][0] ), .B(\mem[253][0] ), .S(n2160), .Z(n17) );
  MUX2_X1 U4851 ( .A(n17), .B(n16), .S(n2100), .Z(n18) );
  MUX2_X1 U4852 ( .A(\mem[250][0] ), .B(\mem[251][0] ), .S(n2163), .Z(n19) );
  MUX2_X1 U4853 ( .A(\mem[248][0] ), .B(\mem[249][0] ), .S(n2163), .Z(n20) );
  MUX2_X1 U4854 ( .A(n20), .B(n19), .S(n2100), .Z(n21) );
  MUX2_X1 U4855 ( .A(n21), .B(n18), .S(n2070), .Z(n22) );
  MUX2_X1 U4856 ( .A(\mem[246][0] ), .B(\mem[247][0] ), .S(n2164), .Z(n23) );
  MUX2_X1 U4857 ( .A(\mem[244][0] ), .B(\mem[245][0] ), .S(n2165), .Z(n24) );
  MUX2_X1 U4858 ( .A(n24), .B(n23), .S(n2100), .Z(n25) );
  MUX2_X1 U4859 ( .A(\mem[242][0] ), .B(\mem[243][0] ), .S(n2162), .Z(n26) );
  MUX2_X1 U4860 ( .A(\mem[240][0] ), .B(\mem[241][0] ), .S(n2162), .Z(n27) );
  MUX2_X1 U4861 ( .A(n27), .B(n26), .S(n2100), .Z(n28) );
  MUX2_X1 U4862 ( .A(n28), .B(n25), .S(n2070), .Z(n29) );
  MUX2_X1 U4863 ( .A(n29), .B(n22), .S(n2057), .Z(n30) );
  MUX2_X1 U4864 ( .A(\mem[238][0] ), .B(\mem[239][0] ), .S(n8), .Z(n31) );
  MUX2_X1 U4865 ( .A(\mem[236][0] ), .B(\mem[237][0] ), .S(n8), .Z(n32) );
  MUX2_X1 U4866 ( .A(n32), .B(n31), .S(n2100), .Z(n33) );
  MUX2_X1 U4867 ( .A(\mem[234][0] ), .B(\mem[235][0] ), .S(n2160), .Z(n34) );
  MUX2_X1 U4868 ( .A(\mem[232][0] ), .B(\mem[233][0] ), .S(n2149), .Z(n35) );
  MUX2_X1 U4869 ( .A(n35), .B(n34), .S(n2100), .Z(n36) );
  MUX2_X1 U4870 ( .A(n36), .B(n33), .S(n2070), .Z(n37) );
  MUX2_X1 U4871 ( .A(\mem[230][0] ), .B(\mem[231][0] ), .S(n7), .Z(n38) );
  MUX2_X1 U4872 ( .A(\mem[228][0] ), .B(\mem[229][0] ), .S(n2148), .Z(n39) );
  MUX2_X1 U4873 ( .A(n39), .B(n38), .S(n2100), .Z(n40) );
  MUX2_X1 U4874 ( .A(\mem[226][0] ), .B(\mem[227][0] ), .S(n7), .Z(n41) );
  MUX2_X1 U4875 ( .A(\mem[224][0] ), .B(\mem[225][0] ), .S(n2148), .Z(n42) );
  MUX2_X1 U4876 ( .A(n42), .B(n41), .S(n2100), .Z(n43) );
  MUX2_X1 U4877 ( .A(n43), .B(n40), .S(n2070), .Z(n44) );
  MUX2_X1 U4878 ( .A(n44), .B(n37), .S(n2057), .Z(n45) );
  MUX2_X1 U4879 ( .A(n45), .B(n30), .S(n2051), .Z(n46) );
  MUX2_X1 U4880 ( .A(\mem[222][0] ), .B(\mem[223][0] ), .S(n2161), .Z(n47) );
  MUX2_X1 U4881 ( .A(\mem[220][0] ), .B(\mem[221][0] ), .S(n3), .Z(n48) );
  MUX2_X1 U4882 ( .A(n48), .B(n47), .S(n2101), .Z(n49) );
  MUX2_X1 U4883 ( .A(\mem[218][0] ), .B(\mem[219][0] ), .S(n4), .Z(n50) );
  MUX2_X1 U4884 ( .A(\mem[216][0] ), .B(\mem[217][0] ), .S(n2174), .Z(n51) );
  MUX2_X1 U4885 ( .A(n51), .B(n50), .S(n2101), .Z(n52) );
  MUX2_X1 U4886 ( .A(n52), .B(n49), .S(n2071), .Z(n53) );
  MUX2_X1 U4887 ( .A(\mem[214][0] ), .B(\mem[215][0] ), .S(n8), .Z(n54) );
  MUX2_X1 U4888 ( .A(\mem[212][0] ), .B(\mem[213][0] ), .S(n2152), .Z(n55) );
  MUX2_X1 U4889 ( .A(n55), .B(n54), .S(n2101), .Z(n56) );
  MUX2_X1 U4890 ( .A(\mem[210][0] ), .B(\mem[211][0] ), .S(n2175), .Z(n57) );
  MUX2_X1 U4891 ( .A(\mem[208][0] ), .B(\mem[209][0] ), .S(n2173), .Z(n58) );
  MUX2_X1 U4892 ( .A(n58), .B(n57), .S(n2101), .Z(n59) );
  MUX2_X1 U4893 ( .A(n59), .B(n56), .S(n2071), .Z(n60) );
  MUX2_X1 U4894 ( .A(n60), .B(n53), .S(n2057), .Z(n61) );
  MUX2_X1 U4895 ( .A(\mem[206][0] ), .B(\mem[207][0] ), .S(n2151), .Z(n62) );
  MUX2_X1 U4896 ( .A(\mem[204][0] ), .B(\mem[205][0] ), .S(n2172), .Z(n63) );
  MUX2_X1 U4897 ( .A(n63), .B(n62), .S(n2101), .Z(n64) );
  MUX2_X1 U4898 ( .A(\mem[202][0] ), .B(\mem[203][0] ), .S(n3), .Z(n65) );
  MUX2_X1 U4899 ( .A(\mem[200][0] ), .B(\mem[201][0] ), .S(n2150), .Z(n66) );
  MUX2_X1 U4900 ( .A(n66), .B(n65), .S(n2101), .Z(n67) );
  MUX2_X1 U4901 ( .A(n67), .B(n64), .S(n2071), .Z(n68) );
  MUX2_X1 U4902 ( .A(\mem[198][0] ), .B(\mem[199][0] ), .S(n2151), .Z(n69) );
  MUX2_X1 U4903 ( .A(\mem[196][0] ), .B(\mem[197][0] ), .S(n2151), .Z(n70) );
  MUX2_X1 U4904 ( .A(n70), .B(n69), .S(n2101), .Z(n71) );
  MUX2_X1 U4905 ( .A(\mem[194][0] ), .B(\mem[195][0] ), .S(n2152), .Z(n72) );
  MUX2_X1 U4906 ( .A(\mem[192][0] ), .B(\mem[193][0] ), .S(n2152), .Z(n73) );
  MUX2_X1 U4907 ( .A(n73), .B(n72), .S(n2101), .Z(n74) );
  MUX2_X1 U4908 ( .A(n74), .B(n71), .S(n2071), .Z(n75) );
  MUX2_X1 U4909 ( .A(n75), .B(n68), .S(n2057), .Z(n76) );
  MUX2_X1 U4910 ( .A(n76), .B(n61), .S(n2051), .Z(n77) );
  MUX2_X1 U4911 ( .A(n77), .B(n46), .S(n2048), .Z(n78) );
  MUX2_X1 U4912 ( .A(\mem[190][0] ), .B(\mem[191][0] ), .S(n2151), .Z(n79) );
  MUX2_X1 U4913 ( .A(\mem[188][0] ), .B(\mem[189][0] ), .S(n2151), .Z(n80) );
  MUX2_X1 U4914 ( .A(n80), .B(n79), .S(n2101), .Z(n81) );
  MUX2_X1 U4915 ( .A(\mem[186][0] ), .B(\mem[187][0] ), .S(n2161), .Z(n82) );
  MUX2_X1 U4916 ( .A(\mem[184][0] ), .B(\mem[185][0] ), .S(n2161), .Z(n83) );
  MUX2_X1 U4917 ( .A(n83), .B(n82), .S(n2101), .Z(n84) );
  MUX2_X1 U4918 ( .A(n84), .B(n81), .S(n2071), .Z(n85) );
  MUX2_X1 U4919 ( .A(\mem[182][0] ), .B(\mem[183][0] ), .S(n2152), .Z(n86) );
  MUX2_X1 U4920 ( .A(\mem[180][0] ), .B(\mem[181][0] ), .S(n2152), .Z(n87) );
  MUX2_X1 U4921 ( .A(n87), .B(n86), .S(n2101), .Z(n88) );
  MUX2_X1 U4922 ( .A(\mem[178][0] ), .B(\mem[179][0] ), .S(n2150), .Z(n89) );
  MUX2_X1 U4923 ( .A(\mem[176][0] ), .B(\mem[177][0] ), .S(n2152), .Z(n90) );
  MUX2_X1 U4924 ( .A(n90), .B(n89), .S(n2101), .Z(n91) );
  MUX2_X1 U4925 ( .A(n91), .B(n88), .S(n2071), .Z(n92) );
  MUX2_X1 U4926 ( .A(n92), .B(n85), .S(n2057), .Z(n93) );
  MUX2_X1 U4927 ( .A(\mem[174][0] ), .B(\mem[175][0] ), .S(n2150), .Z(n94) );
  MUX2_X1 U4928 ( .A(\mem[172][0] ), .B(\mem[173][0] ), .S(n2152), .Z(n95) );
  MUX2_X1 U4929 ( .A(n95), .B(n94), .S(n2102), .Z(n96) );
  MUX2_X1 U4930 ( .A(\mem[170][0] ), .B(\mem[171][0] ), .S(n2150), .Z(n97) );
  MUX2_X1 U4931 ( .A(\mem[168][0] ), .B(\mem[169][0] ), .S(n2173), .Z(n98) );
  MUX2_X1 U4932 ( .A(n98), .B(n97), .S(n2102), .Z(n99) );
  MUX2_X1 U4933 ( .A(n99), .B(n96), .S(n2071), .Z(n100) );
  MUX2_X1 U4934 ( .A(\mem[166][0] ), .B(\mem[167][0] ), .S(n2151), .Z(n101) );
  MUX2_X1 U4935 ( .A(\mem[164][0] ), .B(\mem[165][0] ), .S(n2152), .Z(n102) );
  MUX2_X1 U4936 ( .A(n102), .B(n101), .S(n2102), .Z(n103) );
  MUX2_X1 U4937 ( .A(\mem[162][0] ), .B(\mem[163][0] ), .S(n2173), .Z(n104) );
  MUX2_X1 U4938 ( .A(\mem[160][0] ), .B(\mem[161][0] ), .S(n4), .Z(n105) );
  MUX2_X1 U4939 ( .A(n105), .B(n104), .S(n2102), .Z(n106) );
  MUX2_X1 U4940 ( .A(n106), .B(n103), .S(n2071), .Z(n107) );
  MUX2_X1 U4941 ( .A(n107), .B(n100), .S(n2057), .Z(n108) );
  MUX2_X1 U4942 ( .A(n108), .B(n93), .S(n2051), .Z(n109) );
  MUX2_X1 U4943 ( .A(\mem[158][0] ), .B(\mem[159][0] ), .S(n7), .Z(n110) );
  MUX2_X1 U4944 ( .A(\mem[156][0] ), .B(\mem[157][0] ), .S(n2150), .Z(n111) );
  MUX2_X1 U4945 ( .A(n111), .B(n110), .S(n2102), .Z(n112) );
  MUX2_X1 U4946 ( .A(\mem[154][0] ), .B(\mem[155][0] ), .S(n2151), .Z(n113) );
  MUX2_X1 U4947 ( .A(\mem[152][0] ), .B(\mem[153][0] ), .S(n2150), .Z(n114) );
  MUX2_X1 U4948 ( .A(n114), .B(n113), .S(n2102), .Z(n115) );
  MUX2_X1 U4949 ( .A(n115), .B(n112), .S(n2071), .Z(n116) );
  MUX2_X1 U4950 ( .A(\mem[150][0] ), .B(\mem[151][0] ), .S(n2173), .Z(n117) );
  MUX2_X1 U4951 ( .A(\mem[148][0] ), .B(\mem[149][0] ), .S(n2151), .Z(n118) );
  MUX2_X1 U4952 ( .A(n118), .B(n117), .S(n2102), .Z(n119) );
  MUX2_X1 U4953 ( .A(\mem[146][0] ), .B(\mem[147][0] ), .S(n2151), .Z(n120) );
  MUX2_X1 U4954 ( .A(\mem[144][0] ), .B(\mem[145][0] ), .S(n2151), .Z(n121) );
  MUX2_X1 U4955 ( .A(n121), .B(n120), .S(n2102), .Z(n122) );
  MUX2_X1 U4956 ( .A(n122), .B(n119), .S(n2071), .Z(n123) );
  MUX2_X1 U4957 ( .A(n123), .B(n116), .S(n2057), .Z(n124) );
  MUX2_X1 U4958 ( .A(\mem[142][0] ), .B(\mem[143][0] ), .S(n2173), .Z(n125) );
  MUX2_X1 U4959 ( .A(\mem[140][0] ), .B(\mem[141][0] ), .S(n2150), .Z(n126) );
  MUX2_X1 U4960 ( .A(n126), .B(n125), .S(n2102), .Z(n127) );
  MUX2_X1 U4961 ( .A(\mem[138][0] ), .B(\mem[139][0] ), .S(n2150), .Z(n128) );
  MUX2_X1 U4962 ( .A(\mem[136][0] ), .B(\mem[137][0] ), .S(n2163), .Z(n129) );
  MUX2_X1 U4963 ( .A(n129), .B(n128), .S(n2102), .Z(n130) );
  MUX2_X1 U4964 ( .A(n130), .B(n127), .S(n2071), .Z(n131) );
  MUX2_X1 U4965 ( .A(\mem[134][0] ), .B(\mem[135][0] ), .S(n2151), .Z(n132) );
  MUX2_X1 U4966 ( .A(\mem[132][0] ), .B(\mem[133][0] ), .S(n2152), .Z(n133) );
  MUX2_X1 U4967 ( .A(n133), .B(n132), .S(n2102), .Z(n134) );
  MUX2_X1 U4968 ( .A(\mem[130][0] ), .B(\mem[131][0] ), .S(n2150), .Z(n135) );
  MUX2_X1 U4969 ( .A(\mem[128][0] ), .B(\mem[129][0] ), .S(n2161), .Z(n136) );
  MUX2_X1 U4970 ( .A(n136), .B(n135), .S(n2102), .Z(n137) );
  MUX2_X1 U4971 ( .A(n137), .B(n134), .S(n2071), .Z(n138) );
  MUX2_X1 U4972 ( .A(n138), .B(n131), .S(n2057), .Z(n139) );
  MUX2_X1 U4973 ( .A(n139), .B(n124), .S(n2051), .Z(n140) );
  MUX2_X1 U4974 ( .A(n140), .B(n109), .S(n2048), .Z(n141) );
  MUX2_X1 U4975 ( .A(n141), .B(n78), .S(N24), .Z(n142) );
  MUX2_X1 U4976 ( .A(\mem[126][0] ), .B(\mem[127][0] ), .S(n2154), .Z(n143) );
  MUX2_X1 U4977 ( .A(\mem[124][0] ), .B(\mem[125][0] ), .S(n2154), .Z(n144) );
  MUX2_X1 U4978 ( .A(n144), .B(n143), .S(n2103), .Z(n145) );
  MUX2_X1 U4979 ( .A(\mem[122][0] ), .B(\mem[123][0] ), .S(n2154), .Z(n146) );
  MUX2_X1 U4980 ( .A(\mem[120][0] ), .B(\mem[121][0] ), .S(n2154), .Z(n147) );
  MUX2_X1 U4981 ( .A(n147), .B(n146), .S(n2103), .Z(n148) );
  MUX2_X1 U4982 ( .A(n148), .B(n145), .S(n2072), .Z(n149) );
  MUX2_X1 U4983 ( .A(\mem[118][0] ), .B(\mem[119][0] ), .S(n2154), .Z(n150) );
  MUX2_X1 U4984 ( .A(\mem[116][0] ), .B(\mem[117][0] ), .S(n2154), .Z(n151) );
  MUX2_X1 U4985 ( .A(n151), .B(n150), .S(n2103), .Z(n152) );
  MUX2_X1 U4986 ( .A(\mem[114][0] ), .B(\mem[115][0] ), .S(n2154), .Z(n153) );
  MUX2_X1 U4987 ( .A(\mem[112][0] ), .B(\mem[113][0] ), .S(n2154), .Z(n154) );
  MUX2_X1 U4988 ( .A(n154), .B(n153), .S(n2103), .Z(n155) );
  MUX2_X1 U4989 ( .A(n155), .B(n152), .S(n2072), .Z(n156) );
  MUX2_X1 U4990 ( .A(n156), .B(n149), .S(n2058), .Z(n157) );
  MUX2_X1 U4991 ( .A(\mem[110][0] ), .B(\mem[111][0] ), .S(n2154), .Z(n158) );
  MUX2_X1 U4992 ( .A(\mem[108][0] ), .B(\mem[109][0] ), .S(n2154), .Z(n159) );
  MUX2_X1 U4993 ( .A(n159), .B(n158), .S(n2103), .Z(n160) );
  MUX2_X1 U4994 ( .A(\mem[106][0] ), .B(\mem[107][0] ), .S(n2154), .Z(n161) );
  MUX2_X1 U4995 ( .A(\mem[104][0] ), .B(\mem[105][0] ), .S(n2154), .Z(n162) );
  MUX2_X1 U4996 ( .A(n162), .B(n161), .S(n2103), .Z(n163) );
  MUX2_X1 U4997 ( .A(n163), .B(n160), .S(n2072), .Z(n164) );
  MUX2_X1 U4998 ( .A(\mem[102][0] ), .B(\mem[103][0] ), .S(n2155), .Z(n165) );
  MUX2_X1 U4999 ( .A(\mem[100][0] ), .B(\mem[101][0] ), .S(n2155), .Z(n166) );
  MUX2_X1 U5000 ( .A(n166), .B(n165), .S(n2103), .Z(n167) );
  MUX2_X1 U5001 ( .A(\mem[98][0] ), .B(\mem[99][0] ), .S(n2155), .Z(n168) );
  MUX2_X1 U5002 ( .A(\mem[96][0] ), .B(\mem[97][0] ), .S(n2155), .Z(n169) );
  MUX2_X1 U5003 ( .A(n169), .B(n168), .S(n2103), .Z(n170) );
  MUX2_X1 U5004 ( .A(n170), .B(n167), .S(n2072), .Z(n171) );
  MUX2_X1 U5005 ( .A(n171), .B(n164), .S(n2058), .Z(n172) );
  MUX2_X1 U5006 ( .A(n172), .B(n157), .S(n2052), .Z(n173) );
  MUX2_X1 U5007 ( .A(\mem[94][0] ), .B(\mem[95][0] ), .S(n2155), .Z(n174) );
  MUX2_X1 U5008 ( .A(\mem[92][0] ), .B(\mem[93][0] ), .S(n2155), .Z(n175) );
  MUX2_X1 U5009 ( .A(n175), .B(n174), .S(n2103), .Z(n176) );
  MUX2_X1 U5010 ( .A(\mem[90][0] ), .B(\mem[91][0] ), .S(n2155), .Z(n177) );
  MUX2_X1 U5011 ( .A(\mem[88][0] ), .B(\mem[89][0] ), .S(n2155), .Z(n178) );
  MUX2_X1 U5012 ( .A(n178), .B(n177), .S(n2103), .Z(n179) );
  MUX2_X1 U5013 ( .A(n179), .B(n176), .S(n2072), .Z(n180) );
  MUX2_X1 U5014 ( .A(\mem[86][0] ), .B(\mem[87][0] ), .S(n2155), .Z(n181) );
  MUX2_X1 U5015 ( .A(\mem[84][0] ), .B(\mem[85][0] ), .S(n2155), .Z(n182) );
  MUX2_X1 U5016 ( .A(n182), .B(n181), .S(n2103), .Z(n183) );
  MUX2_X1 U5017 ( .A(\mem[82][0] ), .B(\mem[83][0] ), .S(n2155), .Z(n184) );
  MUX2_X1 U5018 ( .A(\mem[80][0] ), .B(\mem[81][0] ), .S(n2155), .Z(n185) );
  MUX2_X1 U5019 ( .A(n185), .B(n184), .S(n2103), .Z(n186) );
  MUX2_X1 U5020 ( .A(n186), .B(n183), .S(n2072), .Z(n187) );
  MUX2_X1 U5021 ( .A(n187), .B(n180), .S(n2058), .Z(n188) );
  MUX2_X1 U5022 ( .A(\mem[78][0] ), .B(\mem[79][0] ), .S(n2156), .Z(n189) );
  MUX2_X1 U5023 ( .A(\mem[76][0] ), .B(\mem[77][0] ), .S(n2156), .Z(n190) );
  MUX2_X1 U5024 ( .A(n190), .B(n189), .S(n2104), .Z(n191) );
  MUX2_X1 U5025 ( .A(\mem[74][0] ), .B(\mem[75][0] ), .S(n2156), .Z(n192) );
  MUX2_X1 U5026 ( .A(\mem[72][0] ), .B(\mem[73][0] ), .S(n2156), .Z(n193) );
  MUX2_X1 U5027 ( .A(n193), .B(n192), .S(n2104), .Z(n194) );
  MUX2_X1 U5028 ( .A(n194), .B(n191), .S(n2072), .Z(n195) );
  MUX2_X1 U5029 ( .A(\mem[70][0] ), .B(\mem[71][0] ), .S(n2156), .Z(n196) );
  MUX2_X1 U5030 ( .A(\mem[68][0] ), .B(\mem[69][0] ), .S(n2156), .Z(n197) );
  MUX2_X1 U5031 ( .A(n197), .B(n196), .S(n2104), .Z(n198) );
  MUX2_X1 U5032 ( .A(\mem[66][0] ), .B(\mem[67][0] ), .S(n2156), .Z(n199) );
  MUX2_X1 U5033 ( .A(\mem[64][0] ), .B(\mem[65][0] ), .S(n2156), .Z(n200) );
  MUX2_X1 U5034 ( .A(n200), .B(n199), .S(n2104), .Z(n201) );
  MUX2_X1 U5035 ( .A(n201), .B(n198), .S(n2072), .Z(n202) );
  MUX2_X1 U5036 ( .A(n202), .B(n195), .S(n2058), .Z(n203) );
  MUX2_X1 U5037 ( .A(n203), .B(n188), .S(n2052), .Z(n204) );
  MUX2_X1 U5038 ( .A(n204), .B(n173), .S(n2048), .Z(n205) );
  MUX2_X1 U5039 ( .A(\mem[62][0] ), .B(\mem[63][0] ), .S(n2156), .Z(n206) );
  MUX2_X1 U5040 ( .A(\mem[60][0] ), .B(\mem[61][0] ), .S(n2156), .Z(n207) );
  MUX2_X1 U5041 ( .A(n207), .B(n206), .S(n2104), .Z(n208) );
  MUX2_X1 U5042 ( .A(\mem[58][0] ), .B(\mem[59][0] ), .S(n2156), .Z(n209) );
  MUX2_X1 U5043 ( .A(\mem[56][0] ), .B(\mem[57][0] ), .S(n2156), .Z(n210) );
  MUX2_X1 U5044 ( .A(n210), .B(n209), .S(n2104), .Z(n211) );
  MUX2_X1 U5045 ( .A(n211), .B(n208), .S(n2072), .Z(n212) );
  MUX2_X1 U5046 ( .A(\mem[54][0] ), .B(\mem[55][0] ), .S(n2157), .Z(n213) );
  MUX2_X1 U5047 ( .A(\mem[52][0] ), .B(\mem[53][0] ), .S(n2157), .Z(n214) );
  MUX2_X1 U5048 ( .A(n214), .B(n213), .S(n2104), .Z(n215) );
  MUX2_X1 U5049 ( .A(\mem[50][0] ), .B(\mem[51][0] ), .S(n2157), .Z(n216) );
  MUX2_X1 U5050 ( .A(\mem[48][0] ), .B(\mem[49][0] ), .S(n2157), .Z(n217) );
  MUX2_X1 U5051 ( .A(n217), .B(n216), .S(n2104), .Z(n218) );
  MUX2_X1 U5052 ( .A(n218), .B(n215), .S(n2072), .Z(n219) );
  MUX2_X1 U5053 ( .A(n219), .B(n212), .S(n2058), .Z(n220) );
  MUX2_X1 U5054 ( .A(\mem[46][0] ), .B(\mem[47][0] ), .S(n2157), .Z(n221) );
  MUX2_X1 U5055 ( .A(\mem[44][0] ), .B(\mem[45][0] ), .S(n2157), .Z(n222) );
  MUX2_X1 U5056 ( .A(n222), .B(n221), .S(n2104), .Z(n223) );
  MUX2_X1 U5057 ( .A(\mem[42][0] ), .B(\mem[43][0] ), .S(n2157), .Z(n224) );
  MUX2_X1 U5058 ( .A(\mem[40][0] ), .B(\mem[41][0] ), .S(n2157), .Z(n225) );
  MUX2_X1 U5059 ( .A(n225), .B(n224), .S(n2104), .Z(n226) );
  MUX2_X1 U5060 ( .A(n226), .B(n223), .S(n2072), .Z(n227) );
  MUX2_X1 U5061 ( .A(\mem[38][0] ), .B(\mem[39][0] ), .S(n2157), .Z(n228) );
  MUX2_X1 U5062 ( .A(\mem[36][0] ), .B(\mem[37][0] ), .S(n2157), .Z(n229) );
  MUX2_X1 U5063 ( .A(n229), .B(n228), .S(n2104), .Z(n230) );
  MUX2_X1 U5064 ( .A(\mem[34][0] ), .B(\mem[35][0] ), .S(n2157), .Z(n231) );
  MUX2_X1 U5065 ( .A(\mem[32][0] ), .B(\mem[33][0] ), .S(n2157), .Z(n232) );
  MUX2_X1 U5066 ( .A(n232), .B(n231), .S(n2104), .Z(n233) );
  MUX2_X1 U5067 ( .A(n233), .B(n230), .S(n2072), .Z(n234) );
  MUX2_X1 U5068 ( .A(n234), .B(n227), .S(n2058), .Z(n235) );
  MUX2_X1 U5069 ( .A(n235), .B(n220), .S(n2052), .Z(n236) );
  MUX2_X1 U5070 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n2158), .Z(n237) );
  MUX2_X1 U5071 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n2158), .Z(n238) );
  MUX2_X1 U5072 ( .A(n238), .B(n237), .S(n2105), .Z(n239) );
  MUX2_X1 U5073 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n2158), .Z(n240) );
  MUX2_X1 U5074 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n2158), .Z(n241) );
  MUX2_X1 U5075 ( .A(n241), .B(n240), .S(n2105), .Z(n242) );
  MUX2_X1 U5076 ( .A(n242), .B(n239), .S(n2073), .Z(n243) );
  MUX2_X1 U5077 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n2158), .Z(n244) );
  MUX2_X1 U5078 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n2158), .Z(n245) );
  MUX2_X1 U5079 ( .A(n245), .B(n244), .S(n2105), .Z(n246) );
  MUX2_X1 U5080 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n2158), .Z(n247) );
  MUX2_X1 U5081 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n2158), .Z(n248) );
  MUX2_X1 U5082 ( .A(n248), .B(n247), .S(n2105), .Z(n249) );
  MUX2_X1 U5083 ( .A(n249), .B(n246), .S(n2073), .Z(n250) );
  MUX2_X1 U5084 ( .A(n250), .B(n243), .S(n2058), .Z(n251) );
  MUX2_X1 U5085 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n2158), .Z(n252) );
  MUX2_X1 U5086 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n2158), .Z(n253) );
  MUX2_X1 U5087 ( .A(n253), .B(n252), .S(n2105), .Z(n254) );
  MUX2_X1 U5088 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n2158), .Z(n255) );
  MUX2_X1 U5089 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n2158), .Z(n256) );
  MUX2_X1 U5090 ( .A(n256), .B(n255), .S(n2105), .Z(n257) );
  MUX2_X1 U5091 ( .A(n257), .B(n254), .S(n2073), .Z(n258) );
  MUX2_X1 U5092 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n2159), .Z(n259) );
  MUX2_X1 U5093 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n2159), .Z(n260) );
  MUX2_X1 U5094 ( .A(n260), .B(n259), .S(n2105), .Z(n261) );
  MUX2_X1 U5095 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n2159), .Z(n262) );
  MUX2_X1 U5096 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n2159), .Z(n263) );
  MUX2_X1 U5097 ( .A(n263), .B(n262), .S(n2105), .Z(n264) );
  MUX2_X1 U5098 ( .A(n264), .B(n261), .S(n2073), .Z(n265) );
  MUX2_X1 U5099 ( .A(n265), .B(n258), .S(n2058), .Z(n266) );
  MUX2_X1 U5100 ( .A(n266), .B(n251), .S(n2052), .Z(n267) );
  MUX2_X1 U5101 ( .A(n267), .B(n236), .S(n2048), .Z(n268) );
  MUX2_X1 U5102 ( .A(n268), .B(n205), .S(N24), .Z(n269) );
  MUX2_X1 U5103 ( .A(n269), .B(n142), .S(N25), .Z(N33) );
  MUX2_X1 U5104 ( .A(\mem[254][1] ), .B(\mem[255][1] ), .S(n2159), .Z(n270) );
  MUX2_X1 U5105 ( .A(\mem[252][1] ), .B(\mem[253][1] ), .S(n2159), .Z(n271) );
  MUX2_X1 U5106 ( .A(n271), .B(n270), .S(n2105), .Z(n272) );
  MUX2_X1 U5107 ( .A(\mem[250][1] ), .B(\mem[251][1] ), .S(n2159), .Z(n273) );
  MUX2_X1 U5108 ( .A(\mem[248][1] ), .B(\mem[249][1] ), .S(n2159), .Z(n274) );
  MUX2_X1 U5109 ( .A(n274), .B(n273), .S(n2105), .Z(n275) );
  MUX2_X1 U5110 ( .A(n275), .B(n272), .S(n2073), .Z(n276) );
  MUX2_X1 U5111 ( .A(\mem[246][1] ), .B(\mem[247][1] ), .S(n2159), .Z(n277) );
  MUX2_X1 U5112 ( .A(\mem[244][1] ), .B(\mem[245][1] ), .S(n2159), .Z(n278) );
  MUX2_X1 U5113 ( .A(n278), .B(n277), .S(n2105), .Z(n279) );
  MUX2_X1 U5114 ( .A(\mem[242][1] ), .B(\mem[243][1] ), .S(n2159), .Z(n280) );
  MUX2_X1 U5115 ( .A(\mem[240][1] ), .B(\mem[241][1] ), .S(n2159), .Z(n281) );
  MUX2_X1 U5116 ( .A(n281), .B(n280), .S(n2105), .Z(n282) );
  MUX2_X1 U5117 ( .A(n282), .B(n279), .S(n2073), .Z(n283) );
  MUX2_X1 U5118 ( .A(n283), .B(n276), .S(n2058), .Z(n284) );
  MUX2_X1 U5119 ( .A(\mem[238][1] ), .B(\mem[239][1] ), .S(n3), .Z(n285) );
  MUX2_X1 U5120 ( .A(\mem[236][1] ), .B(\mem[237][1] ), .S(n2160), .Z(n286) );
  MUX2_X1 U5121 ( .A(n286), .B(n285), .S(n2106), .Z(n287) );
  MUX2_X1 U5122 ( .A(\mem[234][1] ), .B(\mem[235][1] ), .S(n2148), .Z(n288) );
  MUX2_X1 U5123 ( .A(\mem[232][1] ), .B(\mem[233][1] ), .S(n2162), .Z(n289) );
  MUX2_X1 U5124 ( .A(n289), .B(n288), .S(n2106), .Z(n290) );
  MUX2_X1 U5125 ( .A(n290), .B(n287), .S(n2073), .Z(n291) );
  MUX2_X1 U5126 ( .A(\mem[230][1] ), .B(\mem[231][1] ), .S(n7), .Z(n292) );
  MUX2_X1 U5127 ( .A(\mem[228][1] ), .B(\mem[229][1] ), .S(n8), .Z(n293) );
  MUX2_X1 U5128 ( .A(n293), .B(n292), .S(n2106), .Z(n294) );
  MUX2_X1 U5129 ( .A(\mem[226][1] ), .B(\mem[227][1] ), .S(n2163), .Z(n295) );
  MUX2_X1 U5130 ( .A(\mem[224][1] ), .B(\mem[225][1] ), .S(n2164), .Z(n296) );
  MUX2_X1 U5131 ( .A(n296), .B(n295), .S(n2106), .Z(n297) );
  MUX2_X1 U5132 ( .A(n297), .B(n294), .S(n2073), .Z(n298) );
  MUX2_X1 U5133 ( .A(n298), .B(n291), .S(n2058), .Z(n299) );
  MUX2_X1 U5134 ( .A(n299), .B(n284), .S(n2052), .Z(n300) );
  MUX2_X1 U5135 ( .A(\mem[222][1] ), .B(\mem[223][1] ), .S(n2149), .Z(n301) );
  MUX2_X1 U5136 ( .A(\mem[220][1] ), .B(\mem[221][1] ), .S(n8), .Z(n302) );
  MUX2_X1 U5137 ( .A(n302), .B(n301), .S(n2106), .Z(n303) );
  MUX2_X1 U5138 ( .A(\mem[218][1] ), .B(\mem[219][1] ), .S(n2152), .Z(n304) );
  MUX2_X1 U5139 ( .A(\mem[216][1] ), .B(\mem[217][1] ), .S(n2160), .Z(n305) );
  MUX2_X1 U5140 ( .A(n305), .B(n304), .S(n2106), .Z(n306) );
  MUX2_X1 U5141 ( .A(n306), .B(n303), .S(n2073), .Z(n307) );
  MUX2_X1 U5142 ( .A(\mem[214][1] ), .B(\mem[215][1] ), .S(n2162), .Z(n308) );
  MUX2_X1 U5143 ( .A(\mem[212][1] ), .B(\mem[213][1] ), .S(n2148), .Z(n309) );
  MUX2_X1 U5144 ( .A(n309), .B(n308), .S(n2106), .Z(n310) );
  MUX2_X1 U5145 ( .A(\mem[210][1] ), .B(\mem[211][1] ), .S(n2150), .Z(n311) );
  MUX2_X1 U5146 ( .A(\mem[208][1] ), .B(\mem[209][1] ), .S(n2165), .Z(n312) );
  MUX2_X1 U5147 ( .A(n312), .B(n311), .S(n2106), .Z(n313) );
  MUX2_X1 U5148 ( .A(n313), .B(n310), .S(n2073), .Z(n314) );
  MUX2_X1 U5149 ( .A(n314), .B(n307), .S(n2058), .Z(n315) );
  MUX2_X1 U5150 ( .A(\mem[206][1] ), .B(\mem[207][1] ), .S(n2162), .Z(n316) );
  MUX2_X1 U5151 ( .A(\mem[204][1] ), .B(\mem[205][1] ), .S(n2149), .Z(n317) );
  MUX2_X1 U5152 ( .A(n317), .B(n316), .S(n2106), .Z(n318) );
  MUX2_X1 U5153 ( .A(\mem[202][1] ), .B(\mem[203][1] ), .S(n2148), .Z(n319) );
  MUX2_X1 U5154 ( .A(\mem[200][1] ), .B(\mem[201][1] ), .S(n7), .Z(n320) );
  MUX2_X1 U5155 ( .A(n320), .B(n319), .S(n2106), .Z(n321) );
  MUX2_X1 U5156 ( .A(n321), .B(n318), .S(n2073), .Z(n322) );
  MUX2_X1 U5157 ( .A(\mem[198][1] ), .B(\mem[199][1] ), .S(n7), .Z(n323) );
  MUX2_X1 U5158 ( .A(\mem[196][1] ), .B(\mem[197][1] ), .S(n2152), .Z(n324) );
  MUX2_X1 U5159 ( .A(n324), .B(n323), .S(n2106), .Z(n325) );
  MUX2_X1 U5160 ( .A(\mem[194][1] ), .B(\mem[195][1] ), .S(n2148), .Z(n326) );
  MUX2_X1 U5161 ( .A(\mem[192][1] ), .B(\mem[193][1] ), .S(n2164), .Z(n327) );
  MUX2_X1 U5162 ( .A(n327), .B(n326), .S(n2106), .Z(n328) );
  MUX2_X1 U5163 ( .A(n328), .B(n325), .S(n2073), .Z(n329) );
  MUX2_X1 U5164 ( .A(n329), .B(n322), .S(n2058), .Z(n330) );
  MUX2_X1 U5165 ( .A(n330), .B(n315), .S(n2052), .Z(n331) );
  MUX2_X1 U5166 ( .A(n331), .B(n300), .S(n2048), .Z(n332) );
  MUX2_X1 U5167 ( .A(\mem[190][1] ), .B(\mem[191][1] ), .S(n2148), .Z(n333) );
  MUX2_X1 U5168 ( .A(\mem[188][1] ), .B(\mem[189][1] ), .S(n2174), .Z(n334) );
  MUX2_X1 U5169 ( .A(n334), .B(n333), .S(n2107), .Z(n335) );
  MUX2_X1 U5170 ( .A(\mem[186][1] ), .B(\mem[187][1] ), .S(n2163), .Z(n336) );
  MUX2_X1 U5171 ( .A(\mem[184][1] ), .B(\mem[185][1] ), .S(n2149), .Z(n337) );
  MUX2_X1 U5172 ( .A(n337), .B(n336), .S(n2107), .Z(n338) );
  MUX2_X1 U5173 ( .A(n338), .B(n335), .S(n2074), .Z(n339) );
  MUX2_X1 U5174 ( .A(\mem[182][1] ), .B(\mem[183][1] ), .S(n2164), .Z(n340) );
  MUX2_X1 U5175 ( .A(\mem[180][1] ), .B(\mem[181][1] ), .S(n2149), .Z(n341) );
  MUX2_X1 U5176 ( .A(n341), .B(n340), .S(n2107), .Z(n342) );
  MUX2_X1 U5177 ( .A(\mem[178][1] ), .B(\mem[179][1] ), .S(n2164), .Z(n343) );
  MUX2_X1 U5178 ( .A(\mem[176][1] ), .B(\mem[177][1] ), .S(n2148), .Z(n344) );
  MUX2_X1 U5179 ( .A(n344), .B(n343), .S(n2107), .Z(n345) );
  MUX2_X1 U5180 ( .A(n345), .B(n342), .S(n2074), .Z(n346) );
  MUX2_X1 U5181 ( .A(n346), .B(n339), .S(n2059), .Z(n347) );
  MUX2_X1 U5182 ( .A(\mem[174][1] ), .B(\mem[175][1] ), .S(n8), .Z(n348) );
  MUX2_X1 U5183 ( .A(\mem[172][1] ), .B(\mem[173][1] ), .S(n2149), .Z(n349) );
  MUX2_X1 U5184 ( .A(n349), .B(n348), .S(n2107), .Z(n350) );
  MUX2_X1 U5185 ( .A(\mem[170][1] ), .B(\mem[171][1] ), .S(n2164), .Z(n351) );
  MUX2_X1 U5186 ( .A(\mem[168][1] ), .B(\mem[169][1] ), .S(n2149), .Z(n352) );
  MUX2_X1 U5187 ( .A(n352), .B(n351), .S(n2107), .Z(n353) );
  MUX2_X1 U5188 ( .A(n353), .B(n350), .S(n2074), .Z(n354) );
  MUX2_X1 U5189 ( .A(\mem[166][1] ), .B(\mem[167][1] ), .S(n2149), .Z(n355) );
  MUX2_X1 U5190 ( .A(\mem[164][1] ), .B(\mem[165][1] ), .S(n2164), .Z(n356) );
  MUX2_X1 U5191 ( .A(n356), .B(n355), .S(n2107), .Z(n357) );
  MUX2_X1 U5192 ( .A(\mem[162][1] ), .B(\mem[163][1] ), .S(n2148), .Z(n358) );
  MUX2_X1 U5193 ( .A(\mem[160][1] ), .B(\mem[161][1] ), .S(n2165), .Z(n359) );
  MUX2_X1 U5194 ( .A(n359), .B(n358), .S(n2107), .Z(n360) );
  MUX2_X1 U5195 ( .A(n360), .B(n357), .S(n2074), .Z(n361) );
  MUX2_X1 U5196 ( .A(n361), .B(n354), .S(n2059), .Z(n362) );
  MUX2_X1 U5197 ( .A(n362), .B(n347), .S(n2052), .Z(n363) );
  MUX2_X1 U5198 ( .A(\mem[158][1] ), .B(\mem[159][1] ), .S(n2165), .Z(n364) );
  MUX2_X1 U5199 ( .A(\mem[156][1] ), .B(\mem[157][1] ), .S(n2148), .Z(n365) );
  MUX2_X1 U5200 ( .A(n365), .B(n364), .S(n2107), .Z(n366) );
  MUX2_X1 U5201 ( .A(\mem[154][1] ), .B(\mem[155][1] ), .S(n2165), .Z(n367) );
  MUX2_X1 U5202 ( .A(\mem[152][1] ), .B(\mem[153][1] ), .S(n2149), .Z(n368) );
  MUX2_X1 U5203 ( .A(n368), .B(n367), .S(n2107), .Z(n369) );
  MUX2_X1 U5204 ( .A(n369), .B(n366), .S(n2074), .Z(n370) );
  MUX2_X1 U5205 ( .A(\mem[150][1] ), .B(\mem[151][1] ), .S(n2160), .Z(n371) );
  MUX2_X1 U5206 ( .A(\mem[148][1] ), .B(\mem[149][1] ), .S(n2149), .Z(n372) );
  MUX2_X1 U5207 ( .A(n372), .B(n371), .S(n2107), .Z(n373) );
  MUX2_X1 U5208 ( .A(\mem[146][1] ), .B(\mem[147][1] ), .S(n2148), .Z(n374) );
  MUX2_X1 U5209 ( .A(\mem[144][1] ), .B(\mem[145][1] ), .S(n2164), .Z(n375) );
  MUX2_X1 U5210 ( .A(n375), .B(n374), .S(n2107), .Z(n376) );
  MUX2_X1 U5211 ( .A(n376), .B(n373), .S(n2074), .Z(n377) );
  MUX2_X1 U5212 ( .A(n377), .B(n370), .S(n2059), .Z(n378) );
  MUX2_X1 U5213 ( .A(\mem[142][1] ), .B(\mem[143][1] ), .S(n2148), .Z(n379) );
  MUX2_X1 U5214 ( .A(\mem[140][1] ), .B(\mem[141][1] ), .S(n2164), .Z(n380) );
  MUX2_X1 U5215 ( .A(n380), .B(n379), .S(n2108), .Z(n381) );
  MUX2_X1 U5216 ( .A(\mem[138][1] ), .B(\mem[139][1] ), .S(n2164), .Z(n382) );
  MUX2_X1 U5217 ( .A(\mem[136][1] ), .B(\mem[137][1] ), .S(n7), .Z(n383) );
  MUX2_X1 U5218 ( .A(n383), .B(n382), .S(n2108), .Z(n384) );
  MUX2_X1 U5219 ( .A(n384), .B(n381), .S(n2074), .Z(n385) );
  MUX2_X1 U5220 ( .A(\mem[134][1] ), .B(\mem[135][1] ), .S(n2149), .Z(n386) );
  MUX2_X1 U5221 ( .A(\mem[132][1] ), .B(\mem[133][1] ), .S(n2152), .Z(n387) );
  MUX2_X1 U5222 ( .A(n387), .B(n386), .S(n2108), .Z(n388) );
  MUX2_X1 U5223 ( .A(\mem[130][1] ), .B(\mem[131][1] ), .S(n2160), .Z(n389) );
  MUX2_X1 U5224 ( .A(\mem[128][1] ), .B(\mem[129][1] ), .S(n2163), .Z(n390) );
  MUX2_X1 U5225 ( .A(n390), .B(n389), .S(n2108), .Z(n391) );
  MUX2_X1 U5226 ( .A(n391), .B(n388), .S(n2074), .Z(n392) );
  MUX2_X1 U5227 ( .A(n392), .B(n385), .S(n2059), .Z(n393) );
  MUX2_X1 U5228 ( .A(n393), .B(n378), .S(n2052), .Z(n394) );
  MUX2_X1 U5229 ( .A(n394), .B(n363), .S(n2048), .Z(n395) );
  MUX2_X1 U5230 ( .A(n395), .B(n332), .S(N24), .Z(n396) );
  MUX2_X1 U5231 ( .A(\mem[126][1] ), .B(\mem[127][1] ), .S(n2149), .Z(n397) );
  MUX2_X1 U5232 ( .A(\mem[124][1] ), .B(\mem[125][1] ), .S(n2150), .Z(n398) );
  MUX2_X1 U5233 ( .A(n398), .B(n397), .S(n2108), .Z(n399) );
  MUX2_X1 U5234 ( .A(\mem[122][1] ), .B(\mem[123][1] ), .S(n2165), .Z(n400) );
  MUX2_X1 U5235 ( .A(\mem[120][1] ), .B(\mem[121][1] ), .S(n2164), .Z(n401) );
  MUX2_X1 U5236 ( .A(n401), .B(n400), .S(n2108), .Z(n402) );
  MUX2_X1 U5237 ( .A(n402), .B(n399), .S(n2074), .Z(n403) );
  MUX2_X1 U5238 ( .A(\mem[118][1] ), .B(\mem[119][1] ), .S(n2161), .Z(n404) );
  MUX2_X1 U5239 ( .A(\mem[116][1] ), .B(\mem[117][1] ), .S(n8), .Z(n405) );
  MUX2_X1 U5240 ( .A(n405), .B(n404), .S(n2108), .Z(n406) );
  MUX2_X1 U5241 ( .A(\mem[114][1] ), .B(\mem[115][1] ), .S(n2162), .Z(n407) );
  MUX2_X1 U5242 ( .A(\mem[112][1] ), .B(\mem[113][1] ), .S(n2163), .Z(n408) );
  MUX2_X1 U5243 ( .A(n408), .B(n407), .S(n2108), .Z(n409) );
  MUX2_X1 U5244 ( .A(n409), .B(n406), .S(n2074), .Z(n410) );
  MUX2_X1 U5245 ( .A(n410), .B(n403), .S(n2059), .Z(n411) );
  MUX2_X1 U5246 ( .A(\mem[110][1] ), .B(\mem[111][1] ), .S(n2164), .Z(n412) );
  MUX2_X1 U5247 ( .A(\mem[108][1] ), .B(\mem[109][1] ), .S(n2149), .Z(n413) );
  MUX2_X1 U5248 ( .A(n413), .B(n412), .S(n2108), .Z(n414) );
  MUX2_X1 U5249 ( .A(\mem[106][1] ), .B(\mem[107][1] ), .S(n2153), .Z(n415) );
  MUX2_X1 U5250 ( .A(\mem[104][1] ), .B(\mem[105][1] ), .S(n7), .Z(n416) );
  MUX2_X1 U5251 ( .A(n416), .B(n415), .S(n2108), .Z(n417) );
  MUX2_X1 U5252 ( .A(n417), .B(n414), .S(n2074), .Z(n418) );
  MUX2_X1 U5253 ( .A(\mem[102][1] ), .B(\mem[103][1] ), .S(n2160), .Z(n419) );
  MUX2_X1 U5254 ( .A(\mem[100][1] ), .B(\mem[101][1] ), .S(n2148), .Z(n420) );
  MUX2_X1 U5255 ( .A(n420), .B(n419), .S(n2108), .Z(n421) );
  MUX2_X1 U5256 ( .A(\mem[98][1] ), .B(\mem[99][1] ), .S(n2151), .Z(n422) );
  MUX2_X1 U5257 ( .A(\mem[96][1] ), .B(\mem[97][1] ), .S(n2150), .Z(n423) );
  MUX2_X1 U5258 ( .A(n423), .B(n422), .S(n2108), .Z(n424) );
  MUX2_X1 U5259 ( .A(n424), .B(n421), .S(n2074), .Z(n425) );
  MUX2_X1 U5260 ( .A(n425), .B(n418), .S(n2059), .Z(n426) );
  MUX2_X1 U5261 ( .A(n426), .B(n411), .S(n2052), .Z(n427) );
  MUX2_X1 U5262 ( .A(\mem[94][1] ), .B(\mem[95][1] ), .S(n2166), .Z(n428) );
  MUX2_X1 U5263 ( .A(\mem[92][1] ), .B(\mem[93][1] ), .S(n2166), .Z(n429) );
  MUX2_X1 U5264 ( .A(n429), .B(n428), .S(n2109), .Z(n430) );
  MUX2_X1 U5265 ( .A(\mem[90][1] ), .B(\mem[91][1] ), .S(n2166), .Z(n431) );
  MUX2_X1 U5266 ( .A(\mem[88][1] ), .B(\mem[89][1] ), .S(n2166), .Z(n432) );
  MUX2_X1 U5267 ( .A(n432), .B(n431), .S(n2109), .Z(n433) );
  MUX2_X1 U5268 ( .A(n433), .B(n430), .S(n2075), .Z(n434) );
  MUX2_X1 U5269 ( .A(\mem[86][1] ), .B(\mem[87][1] ), .S(n2166), .Z(n435) );
  MUX2_X1 U5270 ( .A(\mem[84][1] ), .B(\mem[85][1] ), .S(n2166), .Z(n436) );
  MUX2_X1 U5271 ( .A(n436), .B(n435), .S(n2109), .Z(n437) );
  MUX2_X1 U5272 ( .A(\mem[82][1] ), .B(\mem[83][1] ), .S(n2166), .Z(n438) );
  MUX2_X1 U5273 ( .A(\mem[80][1] ), .B(\mem[81][1] ), .S(n2166), .Z(n439) );
  MUX2_X1 U5274 ( .A(n439), .B(n438), .S(n2109), .Z(n440) );
  MUX2_X1 U5275 ( .A(n440), .B(n437), .S(n2075), .Z(n441) );
  MUX2_X1 U5276 ( .A(n441), .B(n434), .S(n2059), .Z(n442) );
  MUX2_X1 U5277 ( .A(\mem[78][1] ), .B(\mem[79][1] ), .S(n2166), .Z(n443) );
  MUX2_X1 U5278 ( .A(\mem[76][1] ), .B(\mem[77][1] ), .S(n2166), .Z(n444) );
  MUX2_X1 U5279 ( .A(n444), .B(n443), .S(n2109), .Z(n445) );
  MUX2_X1 U5280 ( .A(\mem[74][1] ), .B(\mem[75][1] ), .S(n2166), .Z(n446) );
  MUX2_X1 U5281 ( .A(\mem[72][1] ), .B(\mem[73][1] ), .S(n2166), .Z(n447) );
  MUX2_X1 U5282 ( .A(n447), .B(n446), .S(n2109), .Z(n448) );
  MUX2_X1 U5283 ( .A(n448), .B(n445), .S(n2075), .Z(n449) );
  MUX2_X1 U5284 ( .A(\mem[70][1] ), .B(\mem[71][1] ), .S(n2167), .Z(n450) );
  MUX2_X1 U5285 ( .A(\mem[68][1] ), .B(\mem[69][1] ), .S(n2167), .Z(n451) );
  MUX2_X1 U5286 ( .A(n451), .B(n450), .S(n2109), .Z(n452) );
  MUX2_X1 U5287 ( .A(\mem[66][1] ), .B(\mem[67][1] ), .S(n2167), .Z(n453) );
  MUX2_X1 U5288 ( .A(\mem[64][1] ), .B(\mem[65][1] ), .S(n2167), .Z(n454) );
  MUX2_X1 U5289 ( .A(n454), .B(n453), .S(n2109), .Z(n455) );
  MUX2_X1 U5290 ( .A(n455), .B(n452), .S(n2075), .Z(n456) );
  MUX2_X1 U5291 ( .A(n456), .B(n449), .S(n2059), .Z(n457) );
  MUX2_X1 U5292 ( .A(n457), .B(n442), .S(n2052), .Z(n458) );
  MUX2_X1 U5293 ( .A(n458), .B(n427), .S(n2048), .Z(n459) );
  MUX2_X1 U5294 ( .A(\mem[62][1] ), .B(\mem[63][1] ), .S(n2167), .Z(n460) );
  MUX2_X1 U5295 ( .A(\mem[60][1] ), .B(\mem[61][1] ), .S(n2167), .Z(n461) );
  MUX2_X1 U5296 ( .A(n461), .B(n460), .S(n2109), .Z(n462) );
  MUX2_X1 U5297 ( .A(\mem[58][1] ), .B(\mem[59][1] ), .S(n2167), .Z(n463) );
  MUX2_X1 U5298 ( .A(\mem[56][1] ), .B(\mem[57][1] ), .S(n2167), .Z(n464) );
  MUX2_X1 U5299 ( .A(n464), .B(n463), .S(n2109), .Z(n465) );
  MUX2_X1 U5300 ( .A(n465), .B(n462), .S(n2075), .Z(n466) );
  MUX2_X1 U5301 ( .A(\mem[54][1] ), .B(\mem[55][1] ), .S(n2167), .Z(n467) );
  MUX2_X1 U5302 ( .A(\mem[52][1] ), .B(\mem[53][1] ), .S(n2167), .Z(n468) );
  MUX2_X1 U5303 ( .A(n468), .B(n467), .S(n2109), .Z(n469) );
  MUX2_X1 U5304 ( .A(\mem[50][1] ), .B(\mem[51][1] ), .S(n2167), .Z(n470) );
  MUX2_X1 U5305 ( .A(\mem[48][1] ), .B(\mem[49][1] ), .S(n2167), .Z(n471) );
  MUX2_X1 U5306 ( .A(n471), .B(n470), .S(n2109), .Z(n472) );
  MUX2_X1 U5307 ( .A(n472), .B(n469), .S(n2075), .Z(n473) );
  MUX2_X1 U5308 ( .A(n473), .B(n466), .S(n2059), .Z(n474) );
  MUX2_X1 U5309 ( .A(\mem[46][1] ), .B(\mem[47][1] ), .S(n2168), .Z(n475) );
  MUX2_X1 U5310 ( .A(\mem[44][1] ), .B(\mem[45][1] ), .S(n2168), .Z(n476) );
  MUX2_X1 U5311 ( .A(n476), .B(n475), .S(n2110), .Z(n477) );
  MUX2_X1 U5312 ( .A(\mem[42][1] ), .B(\mem[43][1] ), .S(n2168), .Z(n478) );
  MUX2_X1 U5313 ( .A(\mem[40][1] ), .B(\mem[41][1] ), .S(n2168), .Z(n479) );
  MUX2_X1 U5314 ( .A(n479), .B(n478), .S(n2110), .Z(n480) );
  MUX2_X1 U5315 ( .A(n480), .B(n477), .S(n2075), .Z(n481) );
  MUX2_X1 U5316 ( .A(\mem[38][1] ), .B(\mem[39][1] ), .S(n2168), .Z(n482) );
  MUX2_X1 U5317 ( .A(\mem[36][1] ), .B(\mem[37][1] ), .S(n2168), .Z(n483) );
  MUX2_X1 U5318 ( .A(n483), .B(n482), .S(n2110), .Z(n484) );
  MUX2_X1 U5319 ( .A(\mem[34][1] ), .B(\mem[35][1] ), .S(n2168), .Z(n485) );
  MUX2_X1 U5320 ( .A(\mem[32][1] ), .B(\mem[33][1] ), .S(n2168), .Z(n486) );
  MUX2_X1 U5321 ( .A(n486), .B(n485), .S(n2110), .Z(n487) );
  MUX2_X1 U5322 ( .A(n487), .B(n484), .S(n2075), .Z(n488) );
  MUX2_X1 U5323 ( .A(n488), .B(n481), .S(n2059), .Z(n489) );
  MUX2_X1 U5324 ( .A(n489), .B(n474), .S(n2052), .Z(n490) );
  MUX2_X1 U5325 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n2168), .Z(n491) );
  MUX2_X1 U5326 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n2168), .Z(n492) );
  MUX2_X1 U5327 ( .A(n492), .B(n491), .S(n2110), .Z(n493) );
  MUX2_X1 U5328 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n2168), .Z(n494) );
  MUX2_X1 U5329 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n2168), .Z(n495) );
  MUX2_X1 U5330 ( .A(n495), .B(n494), .S(n2110), .Z(n496) );
  MUX2_X1 U5331 ( .A(n496), .B(n493), .S(n2075), .Z(n497) );
  MUX2_X1 U5332 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n2169), .Z(n498) );
  MUX2_X1 U5333 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n2169), .Z(n499) );
  MUX2_X1 U5334 ( .A(n499), .B(n498), .S(n2110), .Z(n500) );
  MUX2_X1 U5335 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n2169), .Z(n501) );
  MUX2_X1 U5336 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n2169), .Z(n502) );
  MUX2_X1 U5337 ( .A(n502), .B(n501), .S(n2110), .Z(n503) );
  MUX2_X1 U5338 ( .A(n503), .B(n500), .S(n2075), .Z(n504) );
  MUX2_X1 U5339 ( .A(n504), .B(n497), .S(n2059), .Z(n505) );
  MUX2_X1 U5340 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n2169), .Z(n506) );
  MUX2_X1 U5341 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n2169), .Z(n507) );
  MUX2_X1 U5342 ( .A(n507), .B(n506), .S(n2110), .Z(n508) );
  MUX2_X1 U5343 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n2169), .Z(n509) );
  MUX2_X1 U5344 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n2169), .Z(n510) );
  MUX2_X1 U5345 ( .A(n510), .B(n509), .S(n2110), .Z(n511) );
  MUX2_X1 U5346 ( .A(n511), .B(n508), .S(n2075), .Z(n512) );
  MUX2_X1 U5347 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n2169), .Z(n513) );
  MUX2_X1 U5348 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n2169), .Z(n514) );
  MUX2_X1 U5349 ( .A(n514), .B(n513), .S(n2110), .Z(n515) );
  MUX2_X1 U5350 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n2169), .Z(n516) );
  MUX2_X1 U5351 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n2169), .Z(n517) );
  MUX2_X1 U5352 ( .A(n517), .B(n516), .S(n2110), .Z(n518) );
  MUX2_X1 U5353 ( .A(n518), .B(n515), .S(n2075), .Z(n519) );
  MUX2_X1 U5354 ( .A(n519), .B(n512), .S(n2059), .Z(n520) );
  MUX2_X1 U5355 ( .A(n520), .B(n505), .S(n2052), .Z(n521) );
  MUX2_X1 U5356 ( .A(n521), .B(n490), .S(n2048), .Z(n522) );
  MUX2_X1 U5357 ( .A(n522), .B(n459), .S(N24), .Z(n523) );
  MUX2_X1 U5358 ( .A(\mem[254][2] ), .B(\mem[255][2] ), .S(n2170), .Z(n524) );
  MUX2_X1 U5359 ( .A(\mem[252][2] ), .B(\mem[253][2] ), .S(n2170), .Z(n525) );
  MUX2_X1 U5360 ( .A(n525), .B(n524), .S(n2111), .Z(n526) );
  MUX2_X1 U5361 ( .A(\mem[250][2] ), .B(\mem[251][2] ), .S(n2170), .Z(n527) );
  MUX2_X1 U5362 ( .A(\mem[248][2] ), .B(\mem[249][2] ), .S(n2170), .Z(n528) );
  MUX2_X1 U5363 ( .A(n528), .B(n527), .S(n2111), .Z(n529) );
  MUX2_X1 U5364 ( .A(n529), .B(n526), .S(n2076), .Z(n530) );
  MUX2_X1 U5365 ( .A(\mem[246][2] ), .B(\mem[247][2] ), .S(n2170), .Z(n531) );
  MUX2_X1 U5366 ( .A(\mem[244][2] ), .B(\mem[245][2] ), .S(n2170), .Z(n532) );
  MUX2_X1 U5367 ( .A(n532), .B(n531), .S(n2111), .Z(n533) );
  MUX2_X1 U5368 ( .A(\mem[242][2] ), .B(\mem[243][2] ), .S(n2170), .Z(n534) );
  MUX2_X1 U5369 ( .A(\mem[240][2] ), .B(\mem[241][2] ), .S(n2170), .Z(n535) );
  MUX2_X1 U5370 ( .A(n535), .B(n534), .S(n2111), .Z(n536) );
  MUX2_X1 U5371 ( .A(n536), .B(n533), .S(n2076), .Z(n537) );
  MUX2_X1 U5372 ( .A(n537), .B(n530), .S(n2060), .Z(n538) );
  MUX2_X1 U5373 ( .A(\mem[238][2] ), .B(\mem[239][2] ), .S(n2170), .Z(n539) );
  MUX2_X1 U5374 ( .A(\mem[236][2] ), .B(\mem[237][2] ), .S(n2170), .Z(n540) );
  MUX2_X1 U5375 ( .A(n540), .B(n539), .S(n2111), .Z(n541) );
  MUX2_X1 U5376 ( .A(\mem[234][2] ), .B(\mem[235][2] ), .S(n2170), .Z(n542) );
  MUX2_X1 U5377 ( .A(\mem[232][2] ), .B(\mem[233][2] ), .S(n2170), .Z(n543) );
  MUX2_X1 U5378 ( .A(n543), .B(n542), .S(n2111), .Z(n544) );
  MUX2_X1 U5379 ( .A(n544), .B(n541), .S(n2076), .Z(n545) );
  MUX2_X1 U5380 ( .A(\mem[230][2] ), .B(\mem[231][2] ), .S(n2171), .Z(n546) );
  MUX2_X1 U5381 ( .A(\mem[228][2] ), .B(\mem[229][2] ), .S(n2171), .Z(n547) );
  MUX2_X1 U5382 ( .A(n547), .B(n546), .S(n2111), .Z(n548) );
  MUX2_X1 U5383 ( .A(\mem[226][2] ), .B(\mem[227][2] ), .S(n2171), .Z(n549) );
  MUX2_X1 U5384 ( .A(\mem[224][2] ), .B(\mem[225][2] ), .S(n2171), .Z(n550) );
  MUX2_X1 U5385 ( .A(n550), .B(n549), .S(n2111), .Z(n551) );
  MUX2_X1 U5386 ( .A(n551), .B(n548), .S(n2076), .Z(n552) );
  MUX2_X1 U5387 ( .A(n552), .B(n545), .S(n2060), .Z(n553) );
  MUX2_X1 U5388 ( .A(n553), .B(n538), .S(n2053), .Z(n554) );
  MUX2_X1 U5389 ( .A(\mem[222][2] ), .B(\mem[223][2] ), .S(n2171), .Z(n555) );
  MUX2_X1 U5390 ( .A(\mem[220][2] ), .B(\mem[221][2] ), .S(n2171), .Z(n556) );
  MUX2_X1 U5391 ( .A(n556), .B(n555), .S(n2111), .Z(n557) );
  MUX2_X1 U5392 ( .A(\mem[218][2] ), .B(\mem[219][2] ), .S(n2171), .Z(n558) );
  MUX2_X1 U5393 ( .A(\mem[216][2] ), .B(\mem[217][2] ), .S(n2171), .Z(n559) );
  MUX2_X1 U5394 ( .A(n559), .B(n558), .S(n2111), .Z(n560) );
  MUX2_X1 U5395 ( .A(n560), .B(n557), .S(n2076), .Z(n561) );
  MUX2_X1 U5396 ( .A(\mem[214][2] ), .B(\mem[215][2] ), .S(n2171), .Z(n562) );
  MUX2_X1 U5397 ( .A(\mem[212][2] ), .B(\mem[213][2] ), .S(n2171), .Z(n563) );
  MUX2_X1 U5398 ( .A(n563), .B(n562), .S(n2111), .Z(n564) );
  MUX2_X1 U5399 ( .A(\mem[210][2] ), .B(\mem[211][2] ), .S(n2171), .Z(n565) );
  MUX2_X1 U5400 ( .A(\mem[208][2] ), .B(\mem[209][2] ), .S(n2171), .Z(n566) );
  MUX2_X1 U5401 ( .A(n566), .B(n565), .S(n2111), .Z(n567) );
  MUX2_X1 U5402 ( .A(n567), .B(n564), .S(n2076), .Z(n568) );
  MUX2_X1 U5403 ( .A(n568), .B(n561), .S(n2060), .Z(n569) );
  MUX2_X1 U5404 ( .A(\mem[206][2] ), .B(\mem[207][2] ), .S(n2205), .Z(n570) );
  MUX2_X1 U5405 ( .A(\mem[204][2] ), .B(\mem[205][2] ), .S(n1), .Z(n571) );
  MUX2_X1 U5406 ( .A(n571), .B(n570), .S(n2112), .Z(n572) );
  MUX2_X1 U5407 ( .A(\mem[202][2] ), .B(\mem[203][2] ), .S(n1), .Z(n573) );
  MUX2_X1 U5408 ( .A(\mem[200][2] ), .B(\mem[201][2] ), .S(n2161), .Z(n574) );
  MUX2_X1 U5409 ( .A(n574), .B(n573), .S(n2112), .Z(n575) );
  MUX2_X1 U5410 ( .A(n575), .B(n572), .S(n2076), .Z(n576) );
  MUX2_X1 U5411 ( .A(\mem[198][2] ), .B(\mem[199][2] ), .S(n1), .Z(n577) );
  MUX2_X1 U5412 ( .A(\mem[196][2] ), .B(\mem[197][2] ), .S(n3), .Z(n578) );
  MUX2_X1 U5413 ( .A(n578), .B(n577), .S(n2112), .Z(n579) );
  MUX2_X1 U5414 ( .A(\mem[194][2] ), .B(\mem[195][2] ), .S(n2174), .Z(n580) );
  MUX2_X1 U5415 ( .A(\mem[192][2] ), .B(\mem[193][2] ), .S(n2172), .Z(n581) );
  MUX2_X1 U5416 ( .A(n581), .B(n580), .S(n2112), .Z(n582) );
  MUX2_X1 U5417 ( .A(n582), .B(n579), .S(n2076), .Z(n583) );
  MUX2_X1 U5418 ( .A(n583), .B(n576), .S(n2060), .Z(n584) );
  MUX2_X1 U5419 ( .A(n584), .B(n569), .S(n2053), .Z(n585) );
  MUX2_X1 U5420 ( .A(n585), .B(n554), .S(n2049), .Z(n586) );
  MUX2_X1 U5421 ( .A(\mem[190][2] ), .B(\mem[191][2] ), .S(n2205), .Z(n587) );
  MUX2_X1 U5422 ( .A(\mem[188][2] ), .B(\mem[189][2] ), .S(n2205), .Z(n588) );
  MUX2_X1 U5423 ( .A(n588), .B(n587), .S(n2112), .Z(n589) );
  MUX2_X1 U5424 ( .A(\mem[186][2] ), .B(\mem[187][2] ), .S(n2205), .Z(n590) );
  MUX2_X1 U5425 ( .A(\mem[184][2] ), .B(\mem[185][2] ), .S(n2195), .Z(n591) );
  MUX2_X1 U5426 ( .A(n591), .B(n590), .S(n2112), .Z(n592) );
  MUX2_X1 U5427 ( .A(n592), .B(n589), .S(n2076), .Z(n593) );
  MUX2_X1 U5428 ( .A(\mem[182][2] ), .B(\mem[183][2] ), .S(n4), .Z(n594) );
  MUX2_X1 U5429 ( .A(\mem[180][2] ), .B(\mem[181][2] ), .S(n2173), .Z(n595) );
  MUX2_X1 U5430 ( .A(n595), .B(n594), .S(n2112), .Z(n596) );
  MUX2_X1 U5431 ( .A(\mem[178][2] ), .B(\mem[179][2] ), .S(n4), .Z(n597) );
  MUX2_X1 U5432 ( .A(\mem[176][2] ), .B(\mem[177][2] ), .S(n2173), .Z(n598) );
  MUX2_X1 U5433 ( .A(n598), .B(n597), .S(n2112), .Z(n599) );
  MUX2_X1 U5434 ( .A(n599), .B(n596), .S(n2076), .Z(n600) );
  MUX2_X1 U5435 ( .A(n600), .B(n593), .S(n2060), .Z(n601) );
  MUX2_X1 U5436 ( .A(\mem[174][2] ), .B(\mem[175][2] ), .S(n3), .Z(n602) );
  MUX2_X1 U5437 ( .A(\mem[172][2] ), .B(\mem[173][2] ), .S(n2172), .Z(n603) );
  MUX2_X1 U5438 ( .A(n603), .B(n602), .S(n2112), .Z(n604) );
  MUX2_X1 U5439 ( .A(\mem[170][2] ), .B(\mem[171][2] ), .S(n3), .Z(n605) );
  MUX2_X1 U5440 ( .A(\mem[168][2] ), .B(\mem[169][2] ), .S(n2165), .Z(n606) );
  MUX2_X1 U5441 ( .A(n606), .B(n605), .S(n2112), .Z(n607) );
  MUX2_X1 U5442 ( .A(n607), .B(n604), .S(n2076), .Z(n608) );
  MUX2_X1 U5443 ( .A(\mem[166][2] ), .B(\mem[167][2] ), .S(n2193), .Z(n609) );
  MUX2_X1 U5444 ( .A(\mem[164][2] ), .B(\mem[165][2] ), .S(n2172), .Z(n610) );
  MUX2_X1 U5445 ( .A(n610), .B(n609), .S(n2112), .Z(n611) );
  MUX2_X1 U5446 ( .A(\mem[162][2] ), .B(\mem[163][2] ), .S(n4), .Z(n612) );
  MUX2_X1 U5447 ( .A(\mem[160][2] ), .B(\mem[161][2] ), .S(n2172), .Z(n613) );
  MUX2_X1 U5448 ( .A(n613), .B(n612), .S(n2112), .Z(n614) );
  MUX2_X1 U5449 ( .A(n614), .B(n611), .S(n2076), .Z(n615) );
  MUX2_X1 U5450 ( .A(n615), .B(n608), .S(n2060), .Z(n616) );
  MUX2_X1 U5451 ( .A(n616), .B(n601), .S(n2053), .Z(n617) );
  MUX2_X1 U5452 ( .A(\mem[158][2] ), .B(\mem[159][2] ), .S(n2173), .Z(n618) );
  MUX2_X1 U5453 ( .A(\mem[156][2] ), .B(\mem[157][2] ), .S(n2173), .Z(n619) );
  MUX2_X1 U5454 ( .A(n619), .B(n618), .S(n2131), .Z(n620) );
  MUX2_X1 U5455 ( .A(\mem[154][2] ), .B(\mem[155][2] ), .S(n2175), .Z(n621) );
  MUX2_X1 U5456 ( .A(\mem[152][2] ), .B(\mem[153][2] ), .S(n2172), .Z(n622) );
  MUX2_X1 U5457 ( .A(n622), .B(n621), .S(n2093), .Z(n623) );
  MUX2_X1 U5458 ( .A(n623), .B(n620), .S(n2077), .Z(n624) );
  MUX2_X1 U5459 ( .A(\mem[150][2] ), .B(\mem[151][2] ), .S(n2172), .Z(n625) );
  MUX2_X1 U5460 ( .A(\mem[148][2] ), .B(\mem[149][2] ), .S(n2175), .Z(n626) );
  MUX2_X1 U5461 ( .A(n626), .B(n625), .S(n2093), .Z(n627) );
  MUX2_X1 U5462 ( .A(\mem[146][2] ), .B(\mem[147][2] ), .S(n2153), .Z(n628) );
  MUX2_X1 U5463 ( .A(\mem[144][2] ), .B(\mem[145][2] ), .S(n2172), .Z(n629) );
  MUX2_X1 U5464 ( .A(n629), .B(n628), .S(n2093), .Z(n630) );
  MUX2_X1 U5465 ( .A(n630), .B(n627), .S(n2077), .Z(n631) );
  MUX2_X1 U5466 ( .A(n631), .B(n624), .S(n2060), .Z(n632) );
  MUX2_X1 U5467 ( .A(\mem[142][2] ), .B(\mem[143][2] ), .S(n2153), .Z(n633) );
  MUX2_X1 U5468 ( .A(\mem[140][2] ), .B(\mem[141][2] ), .S(n2173), .Z(n634) );
  MUX2_X1 U5469 ( .A(n634), .B(n633), .S(n2093), .Z(n635) );
  MUX2_X1 U5470 ( .A(\mem[138][2] ), .B(\mem[139][2] ), .S(n2175), .Z(n636) );
  MUX2_X1 U5471 ( .A(\mem[136][2] ), .B(\mem[137][2] ), .S(n2172), .Z(n637) );
  MUX2_X1 U5472 ( .A(n637), .B(n636), .S(n2112), .Z(n638) );
  MUX2_X1 U5473 ( .A(n638), .B(n635), .S(n2077), .Z(n639) );
  MUX2_X1 U5474 ( .A(\mem[134][2] ), .B(\mem[135][2] ), .S(n2153), .Z(n640) );
  MUX2_X1 U5475 ( .A(\mem[132][2] ), .B(\mem[133][2] ), .S(n2173), .Z(n641) );
  MUX2_X1 U5476 ( .A(n641), .B(n640), .S(n2093), .Z(n642) );
  MUX2_X1 U5477 ( .A(\mem[130][2] ), .B(\mem[131][2] ), .S(n2175), .Z(n643) );
  MUX2_X1 U5478 ( .A(\mem[128][2] ), .B(\mem[129][2] ), .S(n2172), .Z(n644) );
  MUX2_X1 U5479 ( .A(n644), .B(n643), .S(n2111), .Z(n645) );
  MUX2_X1 U5480 ( .A(n645), .B(n642), .S(n2077), .Z(n646) );
  MUX2_X1 U5481 ( .A(n646), .B(n639), .S(n2060), .Z(n647) );
  MUX2_X1 U5482 ( .A(n647), .B(n632), .S(n2053), .Z(n648) );
  MUX2_X1 U5483 ( .A(n648), .B(n617), .S(n2049), .Z(n649) );
  MUX2_X1 U5484 ( .A(n649), .B(n586), .S(N24), .Z(n650) );
  MUX2_X1 U5485 ( .A(\mem[126][2] ), .B(\mem[127][2] ), .S(n2174), .Z(n651) );
  MUX2_X1 U5486 ( .A(\mem[124][2] ), .B(\mem[125][2] ), .S(n2172), .Z(n652) );
  MUX2_X1 U5487 ( .A(n652), .B(n651), .S(n2093), .Z(n653) );
  MUX2_X1 U5488 ( .A(\mem[122][2] ), .B(\mem[123][2] ), .S(n2175), .Z(n654) );
  MUX2_X1 U5489 ( .A(\mem[120][2] ), .B(\mem[121][2] ), .S(n2175), .Z(n655) );
  MUX2_X1 U5490 ( .A(n655), .B(n654), .S(n2125), .Z(n656) );
  MUX2_X1 U5491 ( .A(n656), .B(n653), .S(n2077), .Z(n657) );
  MUX2_X1 U5492 ( .A(\mem[118][2] ), .B(\mem[119][2] ), .S(n2153), .Z(n658) );
  MUX2_X1 U5493 ( .A(\mem[116][2] ), .B(\mem[117][2] ), .S(n2153), .Z(n659) );
  MUX2_X1 U5494 ( .A(n659), .B(n658), .S(n2120), .Z(n660) );
  MUX2_X1 U5495 ( .A(\mem[114][2] ), .B(\mem[115][2] ), .S(n2173), .Z(n661) );
  MUX2_X1 U5496 ( .A(\mem[112][2] ), .B(\mem[113][2] ), .S(n2172), .Z(n662) );
  MUX2_X1 U5497 ( .A(n662), .B(n661), .S(n2115), .Z(n663) );
  MUX2_X1 U5498 ( .A(n663), .B(n660), .S(n2077), .Z(n664) );
  MUX2_X1 U5499 ( .A(n664), .B(n657), .S(n2060), .Z(n665) );
  MUX2_X1 U5500 ( .A(\mem[110][2] ), .B(\mem[111][2] ), .S(n2173), .Z(n666) );
  MUX2_X1 U5501 ( .A(\mem[108][2] ), .B(\mem[109][2] ), .S(n4), .Z(n667) );
  MUX2_X1 U5502 ( .A(n667), .B(n666), .S(n2113), .Z(n668) );
  MUX2_X1 U5503 ( .A(\mem[106][2] ), .B(\mem[107][2] ), .S(n2188), .Z(n669) );
  MUX2_X1 U5504 ( .A(\mem[104][2] ), .B(\mem[105][2] ), .S(n2174), .Z(n670) );
  MUX2_X1 U5505 ( .A(n670), .B(n669), .S(n2113), .Z(n671) );
  MUX2_X1 U5506 ( .A(n671), .B(n668), .S(n2077), .Z(n672) );
  MUX2_X1 U5507 ( .A(\mem[102][2] ), .B(\mem[103][2] ), .S(n2160), .Z(n673) );
  MUX2_X1 U5508 ( .A(\mem[100][2] ), .B(\mem[101][2] ), .S(n2161), .Z(n674) );
  MUX2_X1 U5509 ( .A(n674), .B(n673), .S(n2113), .Z(n675) );
  MUX2_X1 U5510 ( .A(\mem[98][2] ), .B(\mem[99][2] ), .S(n3), .Z(n676) );
  MUX2_X1 U5511 ( .A(\mem[96][2] ), .B(\mem[97][2] ), .S(n2153), .Z(n677) );
  MUX2_X1 U5512 ( .A(n677), .B(n676), .S(n2113), .Z(n678) );
  MUX2_X1 U5513 ( .A(n678), .B(n675), .S(n2077), .Z(n679) );
  MUX2_X1 U5514 ( .A(n679), .B(n672), .S(n2060), .Z(n680) );
  MUX2_X1 U5515 ( .A(\mem[94][2] ), .B(\mem[95][2] ), .S(n2174), .Z(n682) );
  MUX2_X1 U5516 ( .A(\mem[92][2] ), .B(\mem[93][2] ), .S(n2155), .Z(n683) );
  MUX2_X1 U5517 ( .A(n683), .B(n682), .S(n2113), .Z(n684) );
  MUX2_X1 U5518 ( .A(\mem[90][2] ), .B(\mem[91][2] ), .S(n4), .Z(n685) );
  MUX2_X1 U5519 ( .A(\mem[88][2] ), .B(\mem[89][2] ), .S(n2174), .Z(n686) );
  MUX2_X1 U5520 ( .A(n686), .B(n685), .S(n2113), .Z(n687) );
  MUX2_X1 U5521 ( .A(n687), .B(n684), .S(n2077), .Z(n688) );
  MUX2_X1 U5522 ( .A(\mem[86][2] ), .B(\mem[87][2] ), .S(n2203), .Z(n689) );
  MUX2_X1 U5523 ( .A(\mem[84][2] ), .B(\mem[85][2] ), .S(n2153), .Z(n690) );
  MUX2_X1 U5524 ( .A(n690), .B(n689), .S(n2113), .Z(n691) );
  MUX2_X1 U5525 ( .A(\mem[82][2] ), .B(\mem[83][2] ), .S(n2175), .Z(n692) );
  MUX2_X1 U5526 ( .A(\mem[80][2] ), .B(\mem[81][2] ), .S(n2172), .Z(n693) );
  MUX2_X1 U5527 ( .A(n693), .B(n692), .S(n2113), .Z(n694) );
  MUX2_X1 U5528 ( .A(n694), .B(n691), .S(n2077), .Z(n695) );
  MUX2_X1 U5529 ( .A(n695), .B(n688), .S(n2060), .Z(n696) );
  MUX2_X1 U5530 ( .A(\mem[78][2] ), .B(\mem[79][2] ), .S(n2153), .Z(n697) );
  MUX2_X1 U5531 ( .A(\mem[76][2] ), .B(\mem[77][2] ), .S(n2153), .Z(n698) );
  MUX2_X1 U5532 ( .A(n698), .B(n697), .S(n2113), .Z(n699) );
  MUX2_X1 U5533 ( .A(\mem[74][2] ), .B(\mem[75][2] ), .S(n2175), .Z(n700) );
  MUX2_X1 U5534 ( .A(\mem[72][2] ), .B(\mem[73][2] ), .S(n2173), .Z(n701) );
  MUX2_X1 U5535 ( .A(n701), .B(n700), .S(n2113), .Z(n702) );
  MUX2_X1 U5536 ( .A(n702), .B(n699), .S(n2077), .Z(n703) );
  MUX2_X1 U5537 ( .A(\mem[70][2] ), .B(\mem[71][2] ), .S(n2175), .Z(n704) );
  MUX2_X1 U5538 ( .A(\mem[68][2] ), .B(\mem[69][2] ), .S(n2175), .Z(n705) );
  MUX2_X1 U5539 ( .A(n705), .B(n704), .S(n2113), .Z(n706) );
  MUX2_X1 U5540 ( .A(\mem[66][2] ), .B(\mem[67][2] ), .S(n2213), .Z(n707) );
  MUX2_X1 U5541 ( .A(\mem[64][2] ), .B(\mem[65][2] ), .S(n3), .Z(n708) );
  MUX2_X1 U5542 ( .A(n708), .B(n707), .S(n2113), .Z(n709) );
  MUX2_X1 U5543 ( .A(n709), .B(n706), .S(n2077), .Z(n710) );
  MUX2_X1 U5544 ( .A(n710), .B(n703), .S(n2060), .Z(n711) );
  MUX2_X1 U5545 ( .A(n711), .B(n696), .S(n2053), .Z(n712) );
  MUX2_X1 U5546 ( .A(n712), .B(n681), .S(n2049), .Z(n713) );
  MUX2_X1 U5547 ( .A(\mem[62][2] ), .B(\mem[63][2] ), .S(n2213), .Z(n714) );
  MUX2_X1 U5548 ( .A(\mem[60][2] ), .B(\mem[61][2] ), .S(n2176), .Z(n715) );
  MUX2_X1 U5549 ( .A(n715), .B(n714), .S(n2114), .Z(n716) );
  MUX2_X1 U5550 ( .A(\mem[58][2] ), .B(\mem[59][2] ), .S(n2176), .Z(n717) );
  MUX2_X1 U5551 ( .A(\mem[56][2] ), .B(\mem[57][2] ), .S(n2176), .Z(n718) );
  MUX2_X1 U5552 ( .A(n718), .B(n717), .S(n2114), .Z(n719) );
  MUX2_X1 U5553 ( .A(n719), .B(n716), .S(n2078), .Z(n720) );
  MUX2_X1 U5554 ( .A(\mem[54][2] ), .B(\mem[55][2] ), .S(n2176), .Z(n721) );
  MUX2_X1 U5555 ( .A(\mem[52][2] ), .B(\mem[53][2] ), .S(n2176), .Z(n722) );
  MUX2_X1 U5556 ( .A(n722), .B(n721), .S(n2114), .Z(n723) );
  MUX2_X1 U5557 ( .A(\mem[50][2] ), .B(\mem[51][2] ), .S(n2176), .Z(n724) );
  MUX2_X1 U5558 ( .A(\mem[48][2] ), .B(\mem[49][2] ), .S(n2176), .Z(n725) );
  MUX2_X1 U5559 ( .A(n725), .B(n724), .S(n2114), .Z(n726) );
  MUX2_X1 U5560 ( .A(n726), .B(n723), .S(n2078), .Z(n727) );
  MUX2_X1 U5561 ( .A(n727), .B(n720), .S(n2061), .Z(n728) );
  MUX2_X1 U5562 ( .A(\mem[46][2] ), .B(\mem[47][2] ), .S(n2176), .Z(n729) );
  MUX2_X1 U5563 ( .A(\mem[44][2] ), .B(\mem[45][2] ), .S(n2176), .Z(n730) );
  MUX2_X1 U5564 ( .A(n730), .B(n729), .S(n2114), .Z(n731) );
  MUX2_X1 U5565 ( .A(\mem[42][2] ), .B(\mem[43][2] ), .S(n2176), .Z(n732) );
  MUX2_X1 U5566 ( .A(\mem[40][2] ), .B(\mem[41][2] ), .S(n2176), .Z(n733) );
  MUX2_X1 U5567 ( .A(n733), .B(n732), .S(n2114), .Z(n734) );
  MUX2_X1 U5568 ( .A(n734), .B(n731), .S(n2078), .Z(n735) );
  MUX2_X1 U5569 ( .A(\mem[38][2] ), .B(\mem[39][2] ), .S(n2206), .Z(n736) );
  MUX2_X1 U5570 ( .A(\mem[36][2] ), .B(\mem[37][2] ), .S(n2177), .Z(n737) );
  MUX2_X1 U5571 ( .A(n737), .B(n736), .S(n2114), .Z(n738) );
  MUX2_X1 U5572 ( .A(\mem[34][2] ), .B(\mem[35][2] ), .S(n2206), .Z(n739) );
  MUX2_X1 U5573 ( .A(\mem[32][2] ), .B(\mem[33][2] ), .S(n2177), .Z(n740) );
  MUX2_X1 U5574 ( .A(n740), .B(n739), .S(n2114), .Z(n741) );
  MUX2_X1 U5575 ( .A(n741), .B(n738), .S(n2078), .Z(n742) );
  MUX2_X1 U5576 ( .A(n742), .B(n735), .S(n2061), .Z(n743) );
  MUX2_X1 U5577 ( .A(n743), .B(n728), .S(n2053), .Z(n744) );
  MUX2_X1 U5578 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n2206), .Z(n745) );
  MUX2_X1 U5579 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n2206), .Z(n746) );
  MUX2_X1 U5580 ( .A(n746), .B(n745), .S(n2114), .Z(n747) );
  MUX2_X1 U5581 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n2206), .Z(n748) );
  MUX2_X1 U5582 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n2177), .Z(n749) );
  MUX2_X1 U5583 ( .A(n749), .B(n748), .S(n2114), .Z(n750) );
  MUX2_X1 U5584 ( .A(n750), .B(n747), .S(n2078), .Z(n751) );
  MUX2_X1 U5585 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n2206), .Z(n752) );
  MUX2_X1 U5586 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n2177), .Z(n753) );
  MUX2_X1 U5587 ( .A(n753), .B(n752), .S(n2114), .Z(n754) );
  MUX2_X1 U5588 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n2206), .Z(n755) );
  MUX2_X1 U5589 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n2177), .Z(n756) );
  MUX2_X1 U5590 ( .A(n756), .B(n755), .S(n2114), .Z(n757) );
  MUX2_X1 U5591 ( .A(n757), .B(n754), .S(n2078), .Z(n758) );
  MUX2_X1 U5592 ( .A(n758), .B(n751), .S(n2061), .Z(n759) );
  MUX2_X1 U5593 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n2184), .Z(n760) );
  MUX2_X1 U5594 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n2178), .Z(n761) );
  MUX2_X1 U5595 ( .A(n761), .B(n760), .S(n2115), .Z(n762) );
  MUX2_X1 U5596 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n2178), .Z(n763) );
  MUX2_X1 U5597 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n2178), .Z(n764) );
  MUX2_X1 U5598 ( .A(n764), .B(n763), .S(n2115), .Z(n765) );
  MUX2_X1 U5599 ( .A(n765), .B(n762), .S(n2078), .Z(n766) );
  MUX2_X1 U5600 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n2178), .Z(n767) );
  MUX2_X1 U5601 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n2178), .Z(n768) );
  MUX2_X1 U5602 ( .A(n768), .B(n767), .S(n2115), .Z(n769) );
  MUX2_X1 U5603 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n2178), .Z(n770) );
  MUX2_X1 U5604 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n2178), .Z(n771) );
  MUX2_X1 U5605 ( .A(n771), .B(n770), .S(n2115), .Z(n772) );
  MUX2_X1 U5606 ( .A(n772), .B(n769), .S(n2078), .Z(n773) );
  MUX2_X1 U5607 ( .A(n773), .B(n766), .S(n2061), .Z(n774) );
  MUX2_X1 U5608 ( .A(n774), .B(n759), .S(n2053), .Z(n775) );
  MUX2_X1 U5609 ( .A(n775), .B(n744), .S(n2049), .Z(n776) );
  MUX2_X1 U5610 ( .A(\mem[254][3] ), .B(\mem[255][3] ), .S(n2178), .Z(n778) );
  MUX2_X1 U5611 ( .A(\mem[252][3] ), .B(\mem[253][3] ), .S(n2178), .Z(n779) );
  MUX2_X1 U5612 ( .A(n779), .B(n778), .S(n2115), .Z(n780) );
  MUX2_X1 U5613 ( .A(\mem[250][3] ), .B(\mem[251][3] ), .S(n2178), .Z(n781) );
  MUX2_X1 U5614 ( .A(\mem[248][3] ), .B(\mem[249][3] ), .S(n2178), .Z(n782) );
  MUX2_X1 U5615 ( .A(n782), .B(n781), .S(n2115), .Z(n783) );
  MUX2_X1 U5616 ( .A(n783), .B(n780), .S(n2078), .Z(n784) );
  MUX2_X1 U5617 ( .A(\mem[246][3] ), .B(\mem[247][3] ), .S(n2179), .Z(n785) );
  MUX2_X1 U5618 ( .A(\mem[244][3] ), .B(\mem[245][3] ), .S(n2179), .Z(n786) );
  MUX2_X1 U5619 ( .A(n786), .B(n785), .S(n2115), .Z(n787) );
  MUX2_X1 U5620 ( .A(\mem[242][3] ), .B(\mem[243][3] ), .S(n2179), .Z(n788) );
  MUX2_X1 U5621 ( .A(\mem[240][3] ), .B(\mem[241][3] ), .S(n2179), .Z(n789) );
  MUX2_X1 U5622 ( .A(n789), .B(n788), .S(n2115), .Z(n790) );
  MUX2_X1 U5623 ( .A(n790), .B(n787), .S(n2078), .Z(n791) );
  MUX2_X1 U5624 ( .A(n791), .B(n784), .S(n2061), .Z(n792) );
  MUX2_X1 U5625 ( .A(\mem[238][3] ), .B(\mem[239][3] ), .S(n2179), .Z(n793) );
  MUX2_X1 U5626 ( .A(\mem[236][3] ), .B(\mem[237][3] ), .S(n2179), .Z(n794) );
  MUX2_X1 U5627 ( .A(n794), .B(n793), .S(n2115), .Z(n795) );
  MUX2_X1 U5628 ( .A(\mem[234][3] ), .B(\mem[235][3] ), .S(n2179), .Z(n796) );
  MUX2_X1 U5629 ( .A(\mem[232][3] ), .B(\mem[233][3] ), .S(n2179), .Z(n797) );
  MUX2_X1 U5630 ( .A(n797), .B(n796), .S(n2115), .Z(n798) );
  MUX2_X1 U5631 ( .A(n798), .B(n795), .S(n2078), .Z(n799) );
  MUX2_X1 U5632 ( .A(\mem[230][3] ), .B(\mem[231][3] ), .S(n2179), .Z(n800) );
  MUX2_X1 U5633 ( .A(\mem[228][3] ), .B(\mem[229][3] ), .S(n2179), .Z(n801) );
  MUX2_X1 U5634 ( .A(n801), .B(n800), .S(n2115), .Z(n802) );
  MUX2_X1 U5635 ( .A(\mem[226][3] ), .B(\mem[227][3] ), .S(n2179), .Z(n803) );
  MUX2_X1 U5636 ( .A(\mem[224][3] ), .B(\mem[225][3] ), .S(n2179), .Z(n804) );
  MUX2_X1 U5637 ( .A(n804), .B(n803), .S(n2115), .Z(n805) );
  MUX2_X1 U5638 ( .A(n805), .B(n802), .S(n2078), .Z(n806) );
  MUX2_X1 U5639 ( .A(n806), .B(n799), .S(n2061), .Z(n807) );
  MUX2_X1 U5640 ( .A(n807), .B(n792), .S(n2053), .Z(n808) );
  MUX2_X1 U5641 ( .A(\mem[222][3] ), .B(\mem[223][3] ), .S(n2180), .Z(n809) );
  MUX2_X1 U5642 ( .A(\mem[220][3] ), .B(\mem[221][3] ), .S(n2180), .Z(n810) );
  MUX2_X1 U5643 ( .A(n810), .B(n809), .S(n2116), .Z(n811) );
  MUX2_X1 U5644 ( .A(\mem[218][3] ), .B(\mem[219][3] ), .S(n2180), .Z(n812) );
  MUX2_X1 U5645 ( .A(\mem[216][3] ), .B(\mem[217][3] ), .S(n2180), .Z(n813) );
  MUX2_X1 U5646 ( .A(n813), .B(n812), .S(n2116), .Z(n814) );
  MUX2_X1 U5647 ( .A(n814), .B(n811), .S(n2079), .Z(n815) );
  MUX2_X1 U5648 ( .A(\mem[214][3] ), .B(\mem[215][3] ), .S(n2180), .Z(n816) );
  MUX2_X1 U5649 ( .A(\mem[212][3] ), .B(\mem[213][3] ), .S(n2180), .Z(n817) );
  MUX2_X1 U5650 ( .A(n817), .B(n816), .S(n2116), .Z(n818) );
  MUX2_X1 U5651 ( .A(\mem[210][3] ), .B(\mem[211][3] ), .S(n2180), .Z(n819) );
  MUX2_X1 U5652 ( .A(\mem[208][3] ), .B(\mem[209][3] ), .S(n2180), .Z(n820) );
  MUX2_X1 U5653 ( .A(n820), .B(n819), .S(n2116), .Z(n821) );
  MUX2_X1 U5654 ( .A(n821), .B(n818), .S(n2079), .Z(n822) );
  MUX2_X1 U5655 ( .A(n822), .B(n815), .S(n2061), .Z(n823) );
  MUX2_X1 U5656 ( .A(\mem[206][3] ), .B(\mem[207][3] ), .S(n2180), .Z(n824) );
  MUX2_X1 U5657 ( .A(\mem[204][3] ), .B(\mem[205][3] ), .S(n2180), .Z(n825) );
  MUX2_X1 U5658 ( .A(n825), .B(n824), .S(n2116), .Z(n826) );
  MUX2_X1 U5659 ( .A(\mem[202][3] ), .B(\mem[203][3] ), .S(n2180), .Z(n827) );
  MUX2_X1 U5660 ( .A(\mem[200][3] ), .B(\mem[201][3] ), .S(n2180), .Z(n828) );
  MUX2_X1 U5661 ( .A(n828), .B(n827), .S(n2116), .Z(n829) );
  MUX2_X1 U5662 ( .A(n829), .B(n826), .S(n2079), .Z(n830) );
  MUX2_X1 U5663 ( .A(\mem[198][3] ), .B(\mem[199][3] ), .S(n2181), .Z(n831) );
  MUX2_X1 U5664 ( .A(\mem[196][3] ), .B(\mem[197][3] ), .S(n2181), .Z(n832) );
  MUX2_X1 U5665 ( .A(n832), .B(n831), .S(n2116), .Z(n833) );
  MUX2_X1 U5666 ( .A(\mem[194][3] ), .B(\mem[195][3] ), .S(n2181), .Z(n834) );
  MUX2_X1 U5667 ( .A(\mem[192][3] ), .B(\mem[193][3] ), .S(n2181), .Z(n835) );
  MUX2_X1 U5668 ( .A(n835), .B(n834), .S(n2116), .Z(n836) );
  MUX2_X1 U5669 ( .A(n836), .B(n833), .S(n2079), .Z(n837) );
  MUX2_X1 U5670 ( .A(n837), .B(n830), .S(n2061), .Z(n838) );
  MUX2_X1 U5671 ( .A(n838), .B(n823), .S(n2053), .Z(n839) );
  MUX2_X1 U5672 ( .A(n839), .B(n808), .S(n2049), .Z(n840) );
  MUX2_X1 U5673 ( .A(\mem[190][3] ), .B(\mem[191][3] ), .S(n2181), .Z(n841) );
  MUX2_X1 U5674 ( .A(\mem[188][3] ), .B(\mem[189][3] ), .S(n2181), .Z(n842) );
  MUX2_X1 U5675 ( .A(n842), .B(n841), .S(n2116), .Z(n843) );
  MUX2_X1 U5676 ( .A(\mem[186][3] ), .B(\mem[187][3] ), .S(n2181), .Z(n844) );
  MUX2_X1 U5677 ( .A(\mem[184][3] ), .B(\mem[185][3] ), .S(n2181), .Z(n845) );
  MUX2_X1 U5678 ( .A(n845), .B(n844), .S(n2116), .Z(n846) );
  MUX2_X1 U5679 ( .A(n846), .B(n843), .S(n2079), .Z(n847) );
  MUX2_X1 U5680 ( .A(\mem[182][3] ), .B(\mem[183][3] ), .S(n2181), .Z(n848) );
  MUX2_X1 U5681 ( .A(\mem[180][3] ), .B(\mem[181][3] ), .S(n2181), .Z(n849) );
  MUX2_X1 U5682 ( .A(n849), .B(n848), .S(n2116), .Z(n850) );
  MUX2_X1 U5683 ( .A(\mem[178][3] ), .B(\mem[179][3] ), .S(n2181), .Z(n851) );
  MUX2_X1 U5684 ( .A(\mem[176][3] ), .B(\mem[177][3] ), .S(n2181), .Z(n852) );
  MUX2_X1 U5685 ( .A(n852), .B(n851), .S(n2116), .Z(n853) );
  MUX2_X1 U5686 ( .A(n853), .B(n850), .S(n2079), .Z(n854) );
  MUX2_X1 U5687 ( .A(n854), .B(n847), .S(n2061), .Z(n855) );
  MUX2_X1 U5688 ( .A(\mem[174][3] ), .B(\mem[175][3] ), .S(n2182), .Z(n856) );
  MUX2_X1 U5689 ( .A(\mem[172][3] ), .B(\mem[173][3] ), .S(n2182), .Z(n857) );
  MUX2_X1 U5690 ( .A(n857), .B(n856), .S(n2117), .Z(n858) );
  MUX2_X1 U5691 ( .A(\mem[170][3] ), .B(\mem[171][3] ), .S(n2182), .Z(n859) );
  MUX2_X1 U5692 ( .A(\mem[168][3] ), .B(\mem[169][3] ), .S(n2182), .Z(n860) );
  MUX2_X1 U5693 ( .A(n860), .B(n859), .S(n2117), .Z(n861) );
  MUX2_X1 U5694 ( .A(n861), .B(n858), .S(n2079), .Z(n862) );
  MUX2_X1 U5695 ( .A(\mem[166][3] ), .B(\mem[167][3] ), .S(n2182), .Z(n863) );
  MUX2_X1 U5696 ( .A(\mem[164][3] ), .B(\mem[165][3] ), .S(n2182), .Z(n864) );
  MUX2_X1 U5697 ( .A(n864), .B(n863), .S(n2117), .Z(n865) );
  MUX2_X1 U5698 ( .A(\mem[162][3] ), .B(\mem[163][3] ), .S(n2182), .Z(n866) );
  MUX2_X1 U5699 ( .A(\mem[160][3] ), .B(\mem[161][3] ), .S(n2182), .Z(n867) );
  MUX2_X1 U5700 ( .A(n867), .B(n866), .S(n2117), .Z(n868) );
  MUX2_X1 U5701 ( .A(n868), .B(n865), .S(n2079), .Z(n869) );
  MUX2_X1 U5702 ( .A(n869), .B(n862), .S(n2061), .Z(n870) );
  MUX2_X1 U5703 ( .A(n870), .B(n855), .S(n2053), .Z(n871) );
  MUX2_X1 U5704 ( .A(\mem[158][3] ), .B(\mem[159][3] ), .S(n2182), .Z(n872) );
  MUX2_X1 U5705 ( .A(\mem[156][3] ), .B(\mem[157][3] ), .S(n2182), .Z(n873) );
  MUX2_X1 U5706 ( .A(n873), .B(n872), .S(n2117), .Z(n874) );
  MUX2_X1 U5707 ( .A(\mem[154][3] ), .B(\mem[155][3] ), .S(n2182), .Z(n875) );
  MUX2_X1 U5708 ( .A(\mem[152][3] ), .B(\mem[153][3] ), .S(n2182), .Z(n876) );
  MUX2_X1 U5709 ( .A(n876), .B(n875), .S(n2117), .Z(n877) );
  MUX2_X1 U5710 ( .A(n877), .B(n874), .S(n2079), .Z(n878) );
  MUX2_X1 U5711 ( .A(\mem[150][3] ), .B(\mem[151][3] ), .S(n2183), .Z(n879) );
  MUX2_X1 U5712 ( .A(\mem[148][3] ), .B(\mem[149][3] ), .S(n2183), .Z(n880) );
  MUX2_X1 U5713 ( .A(n880), .B(n879), .S(n2117), .Z(n881) );
  MUX2_X1 U5714 ( .A(\mem[146][3] ), .B(\mem[147][3] ), .S(n2183), .Z(n882) );
  MUX2_X1 U5715 ( .A(\mem[144][3] ), .B(\mem[145][3] ), .S(n2183), .Z(n883) );
  MUX2_X1 U5716 ( .A(n883), .B(n882), .S(n2117), .Z(n884) );
  MUX2_X1 U5717 ( .A(n884), .B(n881), .S(n2079), .Z(n885) );
  MUX2_X1 U5718 ( .A(n885), .B(n878), .S(n2061), .Z(n886) );
  MUX2_X1 U5719 ( .A(\mem[142][3] ), .B(\mem[143][3] ), .S(n2183), .Z(n887) );
  MUX2_X1 U5720 ( .A(\mem[140][3] ), .B(\mem[141][3] ), .S(n2183), .Z(n888) );
  MUX2_X1 U5721 ( .A(n888), .B(n887), .S(n2117), .Z(n889) );
  MUX2_X1 U5722 ( .A(\mem[138][3] ), .B(\mem[139][3] ), .S(n2183), .Z(n890) );
  MUX2_X1 U5723 ( .A(\mem[136][3] ), .B(\mem[137][3] ), .S(n2183), .Z(n891) );
  MUX2_X1 U5724 ( .A(n891), .B(n890), .S(n2117), .Z(n892) );
  MUX2_X1 U5725 ( .A(n892), .B(n889), .S(n2079), .Z(n893) );
  MUX2_X1 U5726 ( .A(\mem[134][3] ), .B(\mem[135][3] ), .S(n2183), .Z(n894) );
  MUX2_X1 U5727 ( .A(\mem[132][3] ), .B(\mem[133][3] ), .S(n2183), .Z(n895) );
  MUX2_X1 U5728 ( .A(n895), .B(n894), .S(n2117), .Z(n896) );
  MUX2_X1 U5729 ( .A(\mem[130][3] ), .B(\mem[131][3] ), .S(n2183), .Z(n897) );
  MUX2_X1 U5730 ( .A(\mem[128][3] ), .B(\mem[129][3] ), .S(n2183), .Z(n898) );
  MUX2_X1 U5731 ( .A(n898), .B(n897), .S(n2117), .Z(n899) );
  MUX2_X1 U5732 ( .A(n899), .B(n896), .S(n2079), .Z(n900) );
  MUX2_X1 U5733 ( .A(n900), .B(n893), .S(n2061), .Z(n901) );
  MUX2_X1 U5734 ( .A(n901), .B(n886), .S(n2053), .Z(n902) );
  MUX2_X1 U5735 ( .A(n902), .B(n871), .S(n2049), .Z(n903) );
  MUX2_X1 U5736 ( .A(n903), .B(n840), .S(N24), .Z(n904) );
  MUX2_X1 U5737 ( .A(\mem[126][3] ), .B(\mem[127][3] ), .S(n2184), .Z(n905) );
  MUX2_X1 U5738 ( .A(\mem[124][3] ), .B(\mem[125][3] ), .S(n2184), .Z(n906) );
  MUX2_X1 U5739 ( .A(n906), .B(n905), .S(n2118), .Z(n907) );
  MUX2_X1 U5740 ( .A(\mem[122][3] ), .B(\mem[123][3] ), .S(n2184), .Z(n908) );
  MUX2_X1 U5741 ( .A(\mem[120][3] ), .B(\mem[121][3] ), .S(n2184), .Z(n909) );
  MUX2_X1 U5742 ( .A(n909), .B(n908), .S(n2118), .Z(n910) );
  MUX2_X1 U5743 ( .A(n910), .B(n907), .S(n2080), .Z(n911) );
  MUX2_X1 U5744 ( .A(\mem[118][3] ), .B(\mem[119][3] ), .S(n2184), .Z(n912) );
  MUX2_X1 U5745 ( .A(\mem[116][3] ), .B(\mem[117][3] ), .S(n2184), .Z(n913) );
  MUX2_X1 U5746 ( .A(n913), .B(n912), .S(n2118), .Z(n914) );
  MUX2_X1 U5747 ( .A(\mem[114][3] ), .B(\mem[115][3] ), .S(n2184), .Z(n915) );
  MUX2_X1 U5748 ( .A(\mem[112][3] ), .B(\mem[113][3] ), .S(n2184), .Z(n916) );
  MUX2_X1 U5749 ( .A(n916), .B(n915), .S(n2118), .Z(n917) );
  MUX2_X1 U5750 ( .A(n917), .B(n914), .S(n2080), .Z(n918) );
  MUX2_X1 U5751 ( .A(n918), .B(n911), .S(n2062), .Z(n919) );
  MUX2_X1 U5752 ( .A(\mem[110][3] ), .B(\mem[111][3] ), .S(n2184), .Z(n920) );
  MUX2_X1 U5753 ( .A(\mem[108][3] ), .B(\mem[109][3] ), .S(n2184), .Z(n921) );
  MUX2_X1 U5754 ( .A(n921), .B(n920), .S(n2118), .Z(n922) );
  MUX2_X1 U5755 ( .A(\mem[106][3] ), .B(\mem[107][3] ), .S(n2184), .Z(n923) );
  MUX2_X1 U5756 ( .A(\mem[104][3] ), .B(\mem[105][3] ), .S(n2184), .Z(n924) );
  MUX2_X1 U5757 ( .A(n924), .B(n923), .S(n2118), .Z(n925) );
  MUX2_X1 U5758 ( .A(n925), .B(n922), .S(n2080), .Z(n926) );
  MUX2_X1 U5759 ( .A(\mem[102][3] ), .B(\mem[103][3] ), .S(n2185), .Z(n927) );
  MUX2_X1 U5760 ( .A(\mem[100][3] ), .B(\mem[101][3] ), .S(n2185), .Z(n928) );
  MUX2_X1 U5761 ( .A(n928), .B(n927), .S(n2118), .Z(n929) );
  MUX2_X1 U5762 ( .A(\mem[98][3] ), .B(\mem[99][3] ), .S(n2185), .Z(n930) );
  MUX2_X1 U5763 ( .A(\mem[96][3] ), .B(\mem[97][3] ), .S(n2185), .Z(n931) );
  MUX2_X1 U5764 ( .A(n931), .B(n930), .S(n2118), .Z(n932) );
  MUX2_X1 U5765 ( .A(n932), .B(n929), .S(n2080), .Z(n933) );
  MUX2_X1 U5766 ( .A(n933), .B(n926), .S(n2062), .Z(n934) );
  MUX2_X1 U5767 ( .A(n934), .B(n919), .S(n2054), .Z(n935) );
  MUX2_X1 U5768 ( .A(\mem[94][3] ), .B(\mem[95][3] ), .S(n2185), .Z(n936) );
  MUX2_X1 U5769 ( .A(\mem[92][3] ), .B(\mem[93][3] ), .S(n2185), .Z(n937) );
  MUX2_X1 U5770 ( .A(n937), .B(n936), .S(n2118), .Z(n938) );
  MUX2_X1 U5771 ( .A(\mem[90][3] ), .B(\mem[91][3] ), .S(n2185), .Z(n939) );
  MUX2_X1 U5772 ( .A(\mem[88][3] ), .B(\mem[89][3] ), .S(n2185), .Z(n940) );
  MUX2_X1 U5773 ( .A(n940), .B(n939), .S(n2118), .Z(n941) );
  MUX2_X1 U5774 ( .A(n941), .B(n938), .S(n2080), .Z(n942) );
  MUX2_X1 U5775 ( .A(\mem[86][3] ), .B(\mem[87][3] ), .S(n2185), .Z(n943) );
  MUX2_X1 U5776 ( .A(\mem[84][3] ), .B(\mem[85][3] ), .S(n2185), .Z(n944) );
  MUX2_X1 U5777 ( .A(n944), .B(n943), .S(n2118), .Z(n945) );
  MUX2_X1 U5778 ( .A(\mem[82][3] ), .B(\mem[83][3] ), .S(n2185), .Z(n946) );
  MUX2_X1 U5779 ( .A(\mem[80][3] ), .B(\mem[81][3] ), .S(n2185), .Z(n947) );
  MUX2_X1 U5780 ( .A(n947), .B(n946), .S(n2118), .Z(n948) );
  MUX2_X1 U5781 ( .A(n948), .B(n945), .S(n2080), .Z(n949) );
  MUX2_X1 U5782 ( .A(n949), .B(n942), .S(n2062), .Z(n950) );
  MUX2_X1 U5783 ( .A(\mem[78][3] ), .B(\mem[79][3] ), .S(n2186), .Z(n951) );
  MUX2_X1 U5784 ( .A(\mem[76][3] ), .B(\mem[77][3] ), .S(n2186), .Z(n952) );
  MUX2_X1 U5785 ( .A(n952), .B(n951), .S(n2119), .Z(n953) );
  MUX2_X1 U5786 ( .A(\mem[74][3] ), .B(\mem[75][3] ), .S(n2186), .Z(n954) );
  MUX2_X1 U5787 ( .A(\mem[72][3] ), .B(\mem[73][3] ), .S(n2186), .Z(n955) );
  MUX2_X1 U5788 ( .A(n955), .B(n954), .S(n2119), .Z(n956) );
  MUX2_X1 U5789 ( .A(n956), .B(n953), .S(n2080), .Z(n957) );
  MUX2_X1 U5790 ( .A(\mem[70][3] ), .B(\mem[71][3] ), .S(n2186), .Z(n958) );
  MUX2_X1 U5791 ( .A(\mem[68][3] ), .B(\mem[69][3] ), .S(n2186), .Z(n959) );
  MUX2_X1 U5792 ( .A(n959), .B(n958), .S(n2119), .Z(n960) );
  MUX2_X1 U5793 ( .A(\mem[66][3] ), .B(\mem[67][3] ), .S(n2186), .Z(n961) );
  MUX2_X1 U5794 ( .A(\mem[64][3] ), .B(\mem[65][3] ), .S(n2186), .Z(n962) );
  MUX2_X1 U5795 ( .A(n962), .B(n961), .S(n2119), .Z(n963) );
  MUX2_X1 U5796 ( .A(n963), .B(n960), .S(n2080), .Z(n964) );
  MUX2_X1 U5797 ( .A(n964), .B(n957), .S(n2062), .Z(n965) );
  MUX2_X1 U5798 ( .A(n965), .B(n950), .S(n2054), .Z(n966) );
  MUX2_X1 U5799 ( .A(n966), .B(n935), .S(n2049), .Z(n967) );
  MUX2_X1 U5800 ( .A(\mem[62][3] ), .B(\mem[63][3] ), .S(n2186), .Z(n968) );
  MUX2_X1 U5801 ( .A(\mem[60][3] ), .B(\mem[61][3] ), .S(n2186), .Z(n969) );
  MUX2_X1 U5802 ( .A(n969), .B(n968), .S(n2119), .Z(n970) );
  MUX2_X1 U5803 ( .A(\mem[58][3] ), .B(\mem[59][3] ), .S(n2186), .Z(n971) );
  MUX2_X1 U5804 ( .A(\mem[56][3] ), .B(\mem[57][3] ), .S(n2186), .Z(n972) );
  MUX2_X1 U5805 ( .A(n972), .B(n971), .S(n2119), .Z(n973) );
  MUX2_X1 U5806 ( .A(n973), .B(n970), .S(n2080), .Z(n974) );
  MUX2_X1 U5807 ( .A(\mem[54][3] ), .B(\mem[55][3] ), .S(n2187), .Z(n975) );
  MUX2_X1 U5808 ( .A(\mem[52][3] ), .B(\mem[53][3] ), .S(n2187), .Z(n976) );
  MUX2_X1 U5809 ( .A(n976), .B(n975), .S(n2119), .Z(n977) );
  MUX2_X1 U5810 ( .A(\mem[50][3] ), .B(\mem[51][3] ), .S(n2187), .Z(n978) );
  MUX2_X1 U5811 ( .A(\mem[48][3] ), .B(\mem[49][3] ), .S(n2187), .Z(n979) );
  MUX2_X1 U5812 ( .A(n979), .B(n978), .S(n2119), .Z(n980) );
  MUX2_X1 U5813 ( .A(n980), .B(n977), .S(n2080), .Z(n981) );
  MUX2_X1 U5814 ( .A(n981), .B(n974), .S(n2062), .Z(n982) );
  MUX2_X1 U5815 ( .A(\mem[46][3] ), .B(\mem[47][3] ), .S(n2187), .Z(n983) );
  MUX2_X1 U5816 ( .A(\mem[44][3] ), .B(\mem[45][3] ), .S(n2187), .Z(n984) );
  MUX2_X1 U5817 ( .A(n984), .B(n983), .S(n2119), .Z(n985) );
  MUX2_X1 U5818 ( .A(\mem[42][3] ), .B(\mem[43][3] ), .S(n2187), .Z(n986) );
  MUX2_X1 U5819 ( .A(\mem[40][3] ), .B(\mem[41][3] ), .S(n2187), .Z(n987) );
  MUX2_X1 U5820 ( .A(n987), .B(n986), .S(n2119), .Z(n988) );
  MUX2_X1 U5821 ( .A(n988), .B(n985), .S(n2080), .Z(n989) );
  MUX2_X1 U5822 ( .A(\mem[38][3] ), .B(\mem[39][3] ), .S(n2187), .Z(n990) );
  MUX2_X1 U5823 ( .A(\mem[36][3] ), .B(\mem[37][3] ), .S(n2187), .Z(n991) );
  MUX2_X1 U5824 ( .A(n991), .B(n990), .S(n2119), .Z(n992) );
  MUX2_X1 U5825 ( .A(\mem[34][3] ), .B(\mem[35][3] ), .S(n2187), .Z(n993) );
  MUX2_X1 U5826 ( .A(\mem[32][3] ), .B(\mem[33][3] ), .S(n2187), .Z(n994) );
  MUX2_X1 U5827 ( .A(n994), .B(n993), .S(n2119), .Z(n995) );
  MUX2_X1 U5828 ( .A(n995), .B(n992), .S(n2080), .Z(n996) );
  MUX2_X1 U5829 ( .A(n996), .B(n989), .S(n2062), .Z(n997) );
  MUX2_X1 U5830 ( .A(n997), .B(n982), .S(n2054), .Z(n998) );
  MUX2_X1 U5831 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n2142), .Z(n999) );
  MUX2_X1 U5832 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n2148), .Z(n1000) );
  MUX2_X1 U5833 ( .A(n1000), .B(n999), .S(n2120), .Z(n1001) );
  MUX2_X1 U5834 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n2201), .Z(n1002) );
  MUX2_X1 U5835 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n2164), .Z(n1003) );
  MUX2_X1 U5836 ( .A(n1003), .B(n1002), .S(n2120), .Z(n1004) );
  MUX2_X1 U5837 ( .A(n1004), .B(n1001), .S(n2081), .Z(n1005) );
  MUX2_X1 U5838 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n2198), .Z(n1006) );
  MUX2_X1 U5839 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n2200), .Z(n1007) );
  MUX2_X1 U5840 ( .A(n1007), .B(n1006), .S(n2120), .Z(n1008) );
  MUX2_X1 U5841 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n2149), .Z(n1009) );
  MUX2_X1 U5842 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n2199), .Z(n1010) );
  MUX2_X1 U5843 ( .A(n1010), .B(n1009), .S(n2120), .Z(n1011) );
  MUX2_X1 U5844 ( .A(n1011), .B(n1008), .S(n2081), .Z(n1012) );
  MUX2_X1 U5845 ( .A(n1012), .B(n1005), .S(n2062), .Z(n1013) );
  MUX2_X1 U5846 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n2177), .Z(n1014) );
  MUX2_X1 U5847 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n2214), .Z(n1015) );
  MUX2_X1 U5848 ( .A(n1015), .B(n1014), .S(n2120), .Z(n1016) );
  MUX2_X1 U5849 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n2153), .Z(n1017) );
  MUX2_X1 U5850 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n2202), .Z(n1018) );
  MUX2_X1 U5851 ( .A(n1018), .B(n1017), .S(n2120), .Z(n1019) );
  MUX2_X1 U5852 ( .A(n1019), .B(n1016), .S(n2081), .Z(n1020) );
  MUX2_X1 U5853 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n2200), .Z(n1021) );
  MUX2_X1 U5854 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n2200), .Z(n1022) );
  MUX2_X1 U5855 ( .A(n1022), .B(n1021), .S(n2120), .Z(n1023) );
  MUX2_X1 U5856 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n2200), .Z(n1024) );
  MUX2_X1 U5857 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n2200), .Z(n1025) );
  MUX2_X1 U5858 ( .A(n1025), .B(n1024), .S(n2120), .Z(n1026) );
  MUX2_X1 U5859 ( .A(n1026), .B(n1023), .S(n2081), .Z(n1027) );
  MUX2_X1 U5860 ( .A(n1027), .B(n1020), .S(n2062), .Z(n1028) );
  MUX2_X1 U5861 ( .A(n1028), .B(n1013), .S(n2054), .Z(n1029) );
  MUX2_X1 U5862 ( .A(n1029), .B(n998), .S(n2049), .Z(n1030) );
  MUX2_X1 U5863 ( .A(n1030), .B(n967), .S(N24), .Z(n1031) );
  MUX2_X1 U5864 ( .A(\mem[254][4] ), .B(\mem[255][4] ), .S(n2147), .Z(n1032)
         );
  MUX2_X1 U5865 ( .A(\mem[252][4] ), .B(\mem[253][4] ), .S(n2200), .Z(n1033)
         );
  MUX2_X1 U5866 ( .A(n1033), .B(n1032), .S(n2120), .Z(n1034) );
  MUX2_X1 U5867 ( .A(\mem[250][4] ), .B(\mem[251][4] ), .S(n2200), .Z(n1035)
         );
  MUX2_X1 U5868 ( .A(\mem[248][4] ), .B(\mem[249][4] ), .S(n2184), .Z(n1036)
         );
  MUX2_X1 U5869 ( .A(n1036), .B(n1035), .S(n2120), .Z(n1037) );
  MUX2_X1 U5870 ( .A(n1037), .B(n1034), .S(n2081), .Z(n1038) );
  MUX2_X1 U5871 ( .A(\mem[246][4] ), .B(\mem[247][4] ), .S(n2200), .Z(n1039)
         );
  MUX2_X1 U5872 ( .A(\mem[244][4] ), .B(\mem[245][4] ), .S(n2200), .Z(n1040)
         );
  MUX2_X1 U5873 ( .A(n1040), .B(n1039), .S(n2120), .Z(n1041) );
  MUX2_X1 U5874 ( .A(\mem[242][4] ), .B(\mem[243][4] ), .S(n2184), .Z(n1042)
         );
  MUX2_X1 U5875 ( .A(\mem[240][4] ), .B(\mem[241][4] ), .S(n2200), .Z(n1043)
         );
  MUX2_X1 U5876 ( .A(n1043), .B(n1042), .S(n2120), .Z(n1044) );
  MUX2_X1 U5877 ( .A(n1044), .B(n1041), .S(n2081), .Z(n1045) );
  MUX2_X1 U5878 ( .A(n1045), .B(n1038), .S(n2062), .Z(n1046) );
  MUX2_X1 U5879 ( .A(\mem[238][4] ), .B(\mem[239][4] ), .S(n2175), .Z(n1047)
         );
  MUX2_X1 U5880 ( .A(\mem[236][4] ), .B(\mem[237][4] ), .S(n2188), .Z(n1048)
         );
  MUX2_X1 U5881 ( .A(n1048), .B(n1047), .S(n2121), .Z(n1049) );
  MUX2_X1 U5882 ( .A(\mem[234][4] ), .B(\mem[235][4] ), .S(n2172), .Z(n1050)
         );
  MUX2_X1 U5883 ( .A(\mem[232][4] ), .B(\mem[233][4] ), .S(n2188), .Z(n1051)
         );
  MUX2_X1 U5884 ( .A(n1051), .B(n1050), .S(n2121), .Z(n1052) );
  MUX2_X1 U5885 ( .A(n1052), .B(n1049), .S(n2081), .Z(n1053) );
  MUX2_X1 U5886 ( .A(\mem[230][4] ), .B(\mem[231][4] ), .S(n2175), .Z(n1054)
         );
  MUX2_X1 U5887 ( .A(\mem[228][4] ), .B(\mem[229][4] ), .S(n2188), .Z(n1055)
         );
  MUX2_X1 U5888 ( .A(n1055), .B(n1054), .S(n2121), .Z(n1056) );
  MUX2_X1 U5889 ( .A(\mem[226][4] ), .B(\mem[227][4] ), .S(n2188), .Z(n1057)
         );
  MUX2_X1 U5890 ( .A(\mem[224][4] ), .B(\mem[225][4] ), .S(n2188), .Z(n1058)
         );
  MUX2_X1 U5891 ( .A(n1058), .B(n1057), .S(n2121), .Z(n1059) );
  MUX2_X1 U5892 ( .A(n1059), .B(n1056), .S(n2081), .Z(n1060) );
  MUX2_X1 U5893 ( .A(n1060), .B(n1053), .S(n2062), .Z(n1061) );
  MUX2_X1 U5894 ( .A(n1061), .B(n1046), .S(n2054), .Z(n1062) );
  MUX2_X1 U5895 ( .A(\mem[222][4] ), .B(\mem[223][4] ), .S(n2153), .Z(n1063)
         );
  MUX2_X1 U5896 ( .A(\mem[220][4] ), .B(\mem[221][4] ), .S(n2188), .Z(n1064)
         );
  MUX2_X1 U5897 ( .A(n1064), .B(n1063), .S(n2121), .Z(n1065) );
  MUX2_X1 U5898 ( .A(\mem[218][4] ), .B(\mem[219][4] ), .S(n2188), .Z(n1066)
         );
  MUX2_X1 U5899 ( .A(\mem[216][4] ), .B(\mem[217][4] ), .S(n2188), .Z(n1067)
         );
  MUX2_X1 U5900 ( .A(n1067), .B(n1066), .S(n2121), .Z(n1068) );
  MUX2_X1 U5901 ( .A(n1068), .B(n1065), .S(n2081), .Z(n1069) );
  MUX2_X1 U5902 ( .A(\mem[214][4] ), .B(\mem[215][4] ), .S(n2177), .Z(n1070)
         );
  MUX2_X1 U5903 ( .A(\mem[212][4] ), .B(\mem[213][4] ), .S(n2177), .Z(n1071)
         );
  MUX2_X1 U5904 ( .A(n1071), .B(n1070), .S(n2121), .Z(n1072) );
  MUX2_X1 U5905 ( .A(\mem[210][4] ), .B(\mem[211][4] ), .S(n2177), .Z(n1073)
         );
  MUX2_X1 U5906 ( .A(\mem[208][4] ), .B(\mem[209][4] ), .S(n2190), .Z(n1074)
         );
  MUX2_X1 U5907 ( .A(n1074), .B(n1073), .S(n2121), .Z(n1075) );
  MUX2_X1 U5908 ( .A(n1075), .B(n1072), .S(n2081), .Z(n1076) );
  MUX2_X1 U5909 ( .A(n1076), .B(n1069), .S(n2062), .Z(n1077) );
  MUX2_X1 U5910 ( .A(\mem[206][4] ), .B(\mem[207][4] ), .S(n2177), .Z(n1078)
         );
  MUX2_X1 U5911 ( .A(\mem[204][4] ), .B(\mem[205][4] ), .S(n2177), .Z(n1079)
         );
  MUX2_X1 U5912 ( .A(n1079), .B(n1078), .S(n2121), .Z(n1080) );
  MUX2_X1 U5913 ( .A(\mem[202][4] ), .B(\mem[203][4] ), .S(n2177), .Z(n1081)
         );
  MUX2_X1 U5914 ( .A(\mem[200][4] ), .B(\mem[201][4] ), .S(n2189), .Z(n1082)
         );
  MUX2_X1 U5915 ( .A(n1082), .B(n1081), .S(n2121), .Z(n1083) );
  MUX2_X1 U5916 ( .A(n1083), .B(n1080), .S(n2081), .Z(n1084) );
  MUX2_X1 U5917 ( .A(\mem[198][4] ), .B(\mem[199][4] ), .S(n2177), .Z(n1085)
         );
  MUX2_X1 U5918 ( .A(\mem[196][4] ), .B(\mem[197][4] ), .S(n2177), .Z(n1086)
         );
  MUX2_X1 U5919 ( .A(n1086), .B(n1085), .S(n2121), .Z(n1087) );
  MUX2_X1 U5920 ( .A(\mem[194][4] ), .B(\mem[195][4] ), .S(n2177), .Z(n1088)
         );
  MUX2_X1 U5921 ( .A(\mem[192][4] ), .B(\mem[193][4] ), .S(n2209), .Z(n1089)
         );
  MUX2_X1 U5922 ( .A(n1089), .B(n1088), .S(n2121), .Z(n1090) );
  MUX2_X1 U5923 ( .A(n1090), .B(n1087), .S(n2081), .Z(n1091) );
  MUX2_X1 U5924 ( .A(n1091), .B(n1084), .S(n2062), .Z(n1092) );
  MUX2_X1 U5925 ( .A(n1092), .B(n1077), .S(n2054), .Z(n1093) );
  MUX2_X1 U5926 ( .A(n1093), .B(n1062), .S(n2049), .Z(n1094) );
  MUX2_X1 U5927 ( .A(\mem[190][4] ), .B(\mem[191][4] ), .S(n2173), .Z(n1095)
         );
  MUX2_X1 U5928 ( .A(\mem[188][4] ), .B(\mem[189][4] ), .S(n2189), .Z(n1096)
         );
  MUX2_X1 U5929 ( .A(n1096), .B(n1095), .S(n2122), .Z(n1097) );
  MUX2_X1 U5930 ( .A(\mem[186][4] ), .B(\mem[187][4] ), .S(n2161), .Z(n1098)
         );
  MUX2_X1 U5931 ( .A(\mem[184][4] ), .B(\mem[185][4] ), .S(n2189), .Z(n1099)
         );
  MUX2_X1 U5932 ( .A(n1099), .B(n1098), .S(n2122), .Z(n1100) );
  MUX2_X1 U5933 ( .A(n1100), .B(n1097), .S(n2082), .Z(n1101) );
  MUX2_X1 U5934 ( .A(\mem[182][4] ), .B(\mem[183][4] ), .S(n2194), .Z(n1102)
         );
  MUX2_X1 U5935 ( .A(\mem[180][4] ), .B(\mem[181][4] ), .S(n2189), .Z(n1103)
         );
  MUX2_X1 U5936 ( .A(n1103), .B(n1102), .S(n2122), .Z(n1104) );
  MUX2_X1 U5937 ( .A(\mem[178][4] ), .B(\mem[179][4] ), .S(n2189), .Z(n1105)
         );
  MUX2_X1 U5938 ( .A(\mem[176][4] ), .B(\mem[177][4] ), .S(n2189), .Z(n1106)
         );
  MUX2_X1 U5939 ( .A(n1106), .B(n1105), .S(n2122), .Z(n1107) );
  MUX2_X1 U5940 ( .A(n1107), .B(n1104), .S(n2082), .Z(n1108) );
  MUX2_X1 U5941 ( .A(n1108), .B(n1101), .S(n2063), .Z(n1109) );
  MUX2_X1 U5942 ( .A(\mem[174][4] ), .B(\mem[175][4] ), .S(n2171), .Z(n1110)
         );
  MUX2_X1 U5943 ( .A(\mem[172][4] ), .B(\mem[173][4] ), .S(n2189), .Z(n1111)
         );
  MUX2_X1 U5944 ( .A(n1111), .B(n1110), .S(n2122), .Z(n1112) );
  MUX2_X1 U5945 ( .A(\mem[170][4] ), .B(\mem[171][4] ), .S(n2189), .Z(n1113)
         );
  MUX2_X1 U5946 ( .A(\mem[168][4] ), .B(\mem[169][4] ), .S(n2189), .Z(n1114)
         );
  MUX2_X1 U5947 ( .A(n1114), .B(n1113), .S(n2122), .Z(n1115) );
  MUX2_X1 U5948 ( .A(n1115), .B(n1112), .S(n2082), .Z(n1116) );
  MUX2_X1 U5949 ( .A(\mem[166][4] ), .B(\mem[167][4] ), .S(n2153), .Z(n1117)
         );
  MUX2_X1 U5950 ( .A(\mem[164][4] ), .B(\mem[165][4] ), .S(n2190), .Z(n1118)
         );
  MUX2_X1 U5951 ( .A(n1118), .B(n1117), .S(n2122), .Z(n1119) );
  MUX2_X1 U5952 ( .A(\mem[162][4] ), .B(\mem[163][4] ), .S(n2190), .Z(n1120)
         );
  MUX2_X1 U5953 ( .A(\mem[160][4] ), .B(\mem[161][4] ), .S(n2190), .Z(n1121)
         );
  MUX2_X1 U5954 ( .A(n1121), .B(n1120), .S(n2122), .Z(n1122) );
  MUX2_X1 U5955 ( .A(n1122), .B(n1119), .S(n2082), .Z(n1123) );
  MUX2_X1 U5956 ( .A(n1123), .B(n1116), .S(n2063), .Z(n1124) );
  MUX2_X1 U5957 ( .A(n1124), .B(n1109), .S(n2054), .Z(n1125) );
  MUX2_X1 U5958 ( .A(\mem[158][4] ), .B(\mem[159][4] ), .S(n2153), .Z(n1126)
         );
  MUX2_X1 U5959 ( .A(\mem[156][4] ), .B(\mem[157][4] ), .S(n2190), .Z(n1127)
         );
  MUX2_X1 U5960 ( .A(n1127), .B(n1126), .S(n2122), .Z(n1128) );
  MUX2_X1 U5961 ( .A(\mem[154][4] ), .B(\mem[155][4] ), .S(n2175), .Z(n1129)
         );
  MUX2_X1 U5962 ( .A(\mem[152][4] ), .B(\mem[153][4] ), .S(n2190), .Z(n1130)
         );
  MUX2_X1 U5963 ( .A(n1130), .B(n1129), .S(n2122), .Z(n1131) );
  MUX2_X1 U5964 ( .A(n1131), .B(n1128), .S(n2082), .Z(n1132) );
  MUX2_X1 U5965 ( .A(\mem[150][4] ), .B(\mem[151][4] ), .S(n2174), .Z(n1133)
         );
  MUX2_X1 U5966 ( .A(\mem[148][4] ), .B(\mem[149][4] ), .S(n2190), .Z(n1134)
         );
  MUX2_X1 U5967 ( .A(n1134), .B(n1133), .S(n2122), .Z(n1135) );
  MUX2_X1 U5968 ( .A(\mem[146][4] ), .B(\mem[147][4] ), .S(n2190), .Z(n1136)
         );
  MUX2_X1 U5969 ( .A(\mem[144][4] ), .B(\mem[145][4] ), .S(n2190), .Z(n1137)
         );
  MUX2_X1 U5970 ( .A(n1137), .B(n1136), .S(n2122), .Z(n1138) );
  MUX2_X1 U5971 ( .A(n1138), .B(n1135), .S(n2082), .Z(n1139) );
  MUX2_X1 U5972 ( .A(n1139), .B(n1132), .S(n2063), .Z(n1140) );
  MUX2_X1 U5973 ( .A(\mem[142][4] ), .B(\mem[143][4] ), .S(n2174), .Z(n1141)
         );
  MUX2_X1 U5974 ( .A(\mem[140][4] ), .B(\mem[141][4] ), .S(n2174), .Z(n1142)
         );
  MUX2_X1 U5975 ( .A(n1142), .B(n1141), .S(n2123), .Z(n1143) );
  MUX2_X1 U5976 ( .A(\mem[138][4] ), .B(\mem[139][4] ), .S(n2174), .Z(n1144)
         );
  MUX2_X1 U5977 ( .A(\mem[136][4] ), .B(\mem[137][4] ), .S(n2191), .Z(n1145)
         );
  MUX2_X1 U5978 ( .A(n1145), .B(n1144), .S(n2123), .Z(n1146) );
  MUX2_X1 U5979 ( .A(n1146), .B(n1143), .S(n2082), .Z(n1147) );
  MUX2_X1 U5980 ( .A(\mem[134][4] ), .B(\mem[135][4] ), .S(n2174), .Z(n1148)
         );
  MUX2_X1 U5981 ( .A(\mem[132][4] ), .B(\mem[133][4] ), .S(n2191), .Z(n1149)
         );
  MUX2_X1 U5982 ( .A(n1149), .B(n1148), .S(n2123), .Z(n1150) );
  MUX2_X1 U5983 ( .A(\mem[130][4] ), .B(\mem[131][4] ), .S(n2191), .Z(n1151)
         );
  MUX2_X1 U5984 ( .A(\mem[128][4] ), .B(\mem[129][4] ), .S(n2191), .Z(n1152)
         );
  MUX2_X1 U5985 ( .A(n1152), .B(n1151), .S(n2123), .Z(n1153) );
  MUX2_X1 U5986 ( .A(n1153), .B(n1150), .S(n2082), .Z(n1154) );
  MUX2_X1 U5987 ( .A(n1154), .B(n1147), .S(n2063), .Z(n1155) );
  MUX2_X1 U5988 ( .A(n1155), .B(n1140), .S(n2054), .Z(n1156) );
  MUX2_X1 U5989 ( .A(n1156), .B(n1125), .S(n2049), .Z(n1157) );
  MUX2_X1 U5990 ( .A(n1157), .B(n1094), .S(N24), .Z(n1158) );
  MUX2_X1 U5991 ( .A(\mem[126][4] ), .B(\mem[127][4] ), .S(n2174), .Z(n1159)
         );
  MUX2_X1 U5992 ( .A(\mem[124][4] ), .B(\mem[125][4] ), .S(n2174), .Z(n1160)
         );
  MUX2_X1 U5993 ( .A(n1160), .B(n1159), .S(n2123), .Z(n1161) );
  MUX2_X1 U5994 ( .A(\mem[122][4] ), .B(\mem[123][4] ), .S(n2174), .Z(n1162)
         );
  MUX2_X1 U5995 ( .A(\mem[120][4] ), .B(\mem[121][4] ), .S(n2174), .Z(n1163)
         );
  MUX2_X1 U5996 ( .A(n1163), .B(n1162), .S(n2123), .Z(n1164) );
  MUX2_X1 U5997 ( .A(n1164), .B(n1161), .S(n2082), .Z(n1165) );
  MUX2_X1 U5998 ( .A(\mem[118][4] ), .B(\mem[119][4] ), .S(n2192), .Z(n1166)
         );
  MUX2_X1 U5999 ( .A(\mem[116][4] ), .B(\mem[117][4] ), .S(n2192), .Z(n1167)
         );
  MUX2_X1 U6000 ( .A(n1167), .B(n1166), .S(n2123), .Z(n1168) );
  MUX2_X1 U6001 ( .A(\mem[114][4] ), .B(\mem[115][4] ), .S(n2192), .Z(n1169)
         );
  MUX2_X1 U6002 ( .A(\mem[112][4] ), .B(\mem[113][4] ), .S(n2192), .Z(n1170)
         );
  MUX2_X1 U6003 ( .A(n1170), .B(n1169), .S(n2123), .Z(n1171) );
  MUX2_X1 U6004 ( .A(n1171), .B(n1168), .S(n2082), .Z(n1172) );
  MUX2_X1 U6005 ( .A(n1172), .B(n1165), .S(n2063), .Z(n1173) );
  MUX2_X1 U6006 ( .A(\mem[110][4] ), .B(\mem[111][4] ), .S(n2192), .Z(n1174)
         );
  MUX2_X1 U6007 ( .A(\mem[108][4] ), .B(\mem[109][4] ), .S(n2192), .Z(n1175)
         );
  MUX2_X1 U6008 ( .A(n1175), .B(n1174), .S(n2123), .Z(n1176) );
  MUX2_X1 U6009 ( .A(\mem[106][4] ), .B(\mem[107][4] ), .S(n2192), .Z(n1177)
         );
  MUX2_X1 U6010 ( .A(\mem[104][4] ), .B(\mem[105][4] ), .S(n2192), .Z(n1178)
         );
  MUX2_X1 U6011 ( .A(n1178), .B(n1177), .S(n2123), .Z(n1179) );
  MUX2_X1 U6012 ( .A(n1179), .B(n1176), .S(n2082), .Z(n1180) );
  MUX2_X1 U6013 ( .A(\mem[102][4] ), .B(\mem[103][4] ), .S(n2192), .Z(n1181)
         );
  MUX2_X1 U6014 ( .A(\mem[100][4] ), .B(\mem[101][4] ), .S(n2192), .Z(n1182)
         );
  MUX2_X1 U6015 ( .A(n1182), .B(n1181), .S(n2123), .Z(n1183) );
  MUX2_X1 U6016 ( .A(\mem[98][4] ), .B(\mem[99][4] ), .S(n2192), .Z(n1184) );
  MUX2_X1 U6017 ( .A(\mem[96][4] ), .B(\mem[97][4] ), .S(n2192), .Z(n1185) );
  MUX2_X1 U6018 ( .A(n1185), .B(n1184), .S(n2123), .Z(n1186) );
  MUX2_X1 U6019 ( .A(n1186), .B(n1183), .S(n2082), .Z(n1187) );
  MUX2_X1 U6020 ( .A(n1187), .B(n1180), .S(n2063), .Z(n1188) );
  MUX2_X1 U6021 ( .A(n1188), .B(n1173), .S(n2054), .Z(n1189) );
  MUX2_X1 U6022 ( .A(\mem[94][4] ), .B(\mem[95][4] ), .S(n2193), .Z(n1190) );
  MUX2_X1 U6023 ( .A(\mem[92][4] ), .B(\mem[93][4] ), .S(n2193), .Z(n1191) );
  MUX2_X1 U6024 ( .A(n1191), .B(n1190), .S(n2124), .Z(n1192) );
  MUX2_X1 U6025 ( .A(\mem[90][4] ), .B(\mem[91][4] ), .S(n2193), .Z(n1193) );
  MUX2_X1 U6026 ( .A(\mem[88][4] ), .B(\mem[89][4] ), .S(n2193), .Z(n1194) );
  MUX2_X1 U6027 ( .A(n1194), .B(n1193), .S(n2124), .Z(n1195) );
  MUX2_X1 U6028 ( .A(n1195), .B(n1192), .S(n2083), .Z(n1196) );
  MUX2_X1 U6029 ( .A(\mem[86][4] ), .B(\mem[87][4] ), .S(n2193), .Z(n1197) );
  MUX2_X1 U6030 ( .A(\mem[84][4] ), .B(\mem[85][4] ), .S(n2193), .Z(n1198) );
  MUX2_X1 U6031 ( .A(n1198), .B(n1197), .S(n2124), .Z(n1199) );
  MUX2_X1 U6032 ( .A(\mem[82][4] ), .B(\mem[83][4] ), .S(n2193), .Z(n1200) );
  MUX2_X1 U6033 ( .A(\mem[80][4] ), .B(\mem[81][4] ), .S(n2193), .Z(n1201) );
  MUX2_X1 U6034 ( .A(n1201), .B(n1200), .S(n2124), .Z(n1202) );
  MUX2_X1 U6035 ( .A(n1202), .B(n1199), .S(n2083), .Z(n1203) );
  MUX2_X1 U6036 ( .A(n1203), .B(n1196), .S(n2063), .Z(n1204) );
  MUX2_X1 U6037 ( .A(\mem[78][4] ), .B(\mem[79][4] ), .S(n2193), .Z(n1205) );
  MUX2_X1 U6038 ( .A(\mem[76][4] ), .B(\mem[77][4] ), .S(n2193), .Z(n1206) );
  MUX2_X1 U6039 ( .A(n1206), .B(n1205), .S(n2124), .Z(n1207) );
  MUX2_X1 U6040 ( .A(\mem[74][4] ), .B(\mem[75][4] ), .S(n2193), .Z(n1208) );
  MUX2_X1 U6041 ( .A(\mem[72][4] ), .B(\mem[73][4] ), .S(n2193), .Z(n1209) );
  MUX2_X1 U6042 ( .A(n1209), .B(n1208), .S(n2124), .Z(n1210) );
  MUX2_X1 U6043 ( .A(n1210), .B(n1207), .S(n2083), .Z(n1211) );
  MUX2_X1 U6044 ( .A(\mem[70][4] ), .B(\mem[71][4] ), .S(n2194), .Z(n1212) );
  MUX2_X1 U6045 ( .A(\mem[68][4] ), .B(\mem[69][4] ), .S(n2194), .Z(n1213) );
  MUX2_X1 U6046 ( .A(n1213), .B(n1212), .S(n2124), .Z(n1214) );
  MUX2_X1 U6047 ( .A(\mem[66][4] ), .B(\mem[67][4] ), .S(n2194), .Z(n1215) );
  MUX2_X1 U6048 ( .A(\mem[64][4] ), .B(\mem[65][4] ), .S(n2194), .Z(n1216) );
  MUX2_X1 U6049 ( .A(n1216), .B(n1215), .S(n2124), .Z(n1217) );
  MUX2_X1 U6050 ( .A(n1217), .B(n1214), .S(n2083), .Z(n1218) );
  MUX2_X1 U6051 ( .A(n1218), .B(n1211), .S(n2063), .Z(n1219) );
  MUX2_X1 U6052 ( .A(n1219), .B(n1204), .S(n2054), .Z(n1220) );
  MUX2_X1 U6053 ( .A(n1220), .B(n1189), .S(n2049), .Z(n1221) );
  MUX2_X1 U6054 ( .A(\mem[62][4] ), .B(\mem[63][4] ), .S(n2194), .Z(n1222) );
  MUX2_X1 U6055 ( .A(\mem[60][4] ), .B(\mem[61][4] ), .S(n2194), .Z(n1223) );
  MUX2_X1 U6056 ( .A(n1223), .B(n1222), .S(n2124), .Z(n1224) );
  MUX2_X1 U6057 ( .A(\mem[58][4] ), .B(\mem[59][4] ), .S(n2194), .Z(n1225) );
  MUX2_X1 U6058 ( .A(\mem[56][4] ), .B(\mem[57][4] ), .S(n2194), .Z(n1226) );
  MUX2_X1 U6059 ( .A(n1226), .B(n1225), .S(n2124), .Z(n1227) );
  MUX2_X1 U6060 ( .A(n1227), .B(n1224), .S(n2083), .Z(n1228) );
  MUX2_X1 U6061 ( .A(\mem[54][4] ), .B(\mem[55][4] ), .S(n2194), .Z(n1229) );
  MUX2_X1 U6062 ( .A(\mem[52][4] ), .B(\mem[53][4] ), .S(n2194), .Z(n1230) );
  MUX2_X1 U6063 ( .A(n1230), .B(n1229), .S(n2124), .Z(n1231) );
  MUX2_X1 U6064 ( .A(\mem[50][4] ), .B(\mem[51][4] ), .S(n2194), .Z(n1232) );
  MUX2_X1 U6065 ( .A(\mem[48][4] ), .B(\mem[49][4] ), .S(n2194), .Z(n1233) );
  MUX2_X1 U6066 ( .A(n1233), .B(n1232), .S(n2124), .Z(n1234) );
  MUX2_X1 U6067 ( .A(n1234), .B(n1231), .S(n2083), .Z(n1235) );
  MUX2_X1 U6068 ( .A(n1235), .B(n1228), .S(n2063), .Z(n1236) );
  MUX2_X1 U6069 ( .A(\mem[46][4] ), .B(\mem[47][4] ), .S(n2195), .Z(n1237) );
  MUX2_X1 U6070 ( .A(\mem[44][4] ), .B(\mem[45][4] ), .S(n2195), .Z(n1238) );
  MUX2_X1 U6071 ( .A(n1238), .B(n1237), .S(n2125), .Z(n1239) );
  MUX2_X1 U6072 ( .A(\mem[42][4] ), .B(\mem[43][4] ), .S(n2195), .Z(n1240) );
  MUX2_X1 U6073 ( .A(\mem[40][4] ), .B(\mem[41][4] ), .S(n2195), .Z(n1241) );
  MUX2_X1 U6074 ( .A(n1241), .B(n1240), .S(n2125), .Z(n1242) );
  MUX2_X1 U6075 ( .A(n1242), .B(n1239), .S(n2083), .Z(n1243) );
  MUX2_X1 U6076 ( .A(\mem[38][4] ), .B(\mem[39][4] ), .S(n2195), .Z(n1244) );
  MUX2_X1 U6077 ( .A(\mem[36][4] ), .B(\mem[37][4] ), .S(n2195), .Z(n1245) );
  MUX2_X1 U6078 ( .A(n1245), .B(n1244), .S(n2125), .Z(n1246) );
  MUX2_X1 U6079 ( .A(\mem[34][4] ), .B(\mem[35][4] ), .S(n2195), .Z(n1247) );
  MUX2_X1 U6080 ( .A(\mem[32][4] ), .B(\mem[33][4] ), .S(n2195), .Z(n1248) );
  MUX2_X1 U6081 ( .A(n1248), .B(n1247), .S(n2125), .Z(n1249) );
  MUX2_X1 U6082 ( .A(n1249), .B(n1246), .S(n2083), .Z(n1250) );
  MUX2_X1 U6083 ( .A(n1250), .B(n1243), .S(n2063), .Z(n1251) );
  MUX2_X1 U6084 ( .A(n1251), .B(n1236), .S(n2054), .Z(n1252) );
  MUX2_X1 U6085 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n2195), .Z(n1253) );
  MUX2_X1 U6086 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n2195), .Z(n1254) );
  MUX2_X1 U6087 ( .A(n1254), .B(n1253), .S(n2125), .Z(n1255) );
  MUX2_X1 U6088 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n2195), .Z(n1256) );
  MUX2_X1 U6089 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n2195), .Z(n1257) );
  MUX2_X1 U6090 ( .A(n1257), .B(n1256), .S(n2125), .Z(n1258) );
  MUX2_X1 U6091 ( .A(n1258), .B(n1255), .S(n2083), .Z(n1259) );
  MUX2_X1 U6092 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n2196), .Z(n1260) );
  MUX2_X1 U6093 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n2196), .Z(n1261) );
  MUX2_X1 U6094 ( .A(n1261), .B(n1260), .S(n2125), .Z(n1262) );
  MUX2_X1 U6095 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n2196), .Z(n1263) );
  MUX2_X1 U6096 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n2196), .Z(n1264) );
  MUX2_X1 U6097 ( .A(n1264), .B(n1263), .S(n2125), .Z(n1265) );
  MUX2_X1 U6098 ( .A(n1265), .B(n1262), .S(n2083), .Z(n1266) );
  MUX2_X1 U6099 ( .A(n1266), .B(n1259), .S(n2063), .Z(n1267) );
  MUX2_X1 U6100 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n2196), .Z(n1268) );
  MUX2_X1 U6101 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n2196), .Z(n1269) );
  MUX2_X1 U6102 ( .A(n1269), .B(n1268), .S(n2125), .Z(n1270) );
  MUX2_X1 U6103 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n2196), .Z(n1271) );
  MUX2_X1 U6104 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n2196), .Z(n1272) );
  MUX2_X1 U6105 ( .A(n1272), .B(n1271), .S(n2125), .Z(n1273) );
  MUX2_X1 U6106 ( .A(n1273), .B(n1270), .S(n2083), .Z(n1274) );
  MUX2_X1 U6107 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n2196), .Z(n1275) );
  MUX2_X1 U6108 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n2196), .Z(n1276) );
  MUX2_X1 U6109 ( .A(n1276), .B(n1275), .S(n2125), .Z(n1277) );
  MUX2_X1 U6110 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n2196), .Z(n1278) );
  MUX2_X1 U6111 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n2196), .Z(n1279) );
  MUX2_X1 U6112 ( .A(n1279), .B(n1278), .S(n2125), .Z(n1280) );
  MUX2_X1 U6113 ( .A(n1280), .B(n1277), .S(n2083), .Z(n1281) );
  MUX2_X1 U6114 ( .A(n1281), .B(n1274), .S(n2063), .Z(n1282) );
  MUX2_X1 U6115 ( .A(n1282), .B(n1267), .S(n2054), .Z(n1283) );
  MUX2_X1 U6116 ( .A(n1283), .B(n1252), .S(n2049), .Z(n1284) );
  MUX2_X1 U6117 ( .A(n1284), .B(n1221), .S(N24), .Z(n1285) );
  MUX2_X1 U6118 ( .A(\mem[254][5] ), .B(\mem[255][5] ), .S(n2155), .Z(n1286)
         );
  MUX2_X1 U6119 ( .A(\mem[252][5] ), .B(\mem[253][5] ), .S(n2155), .Z(n1287)
         );
  MUX2_X1 U6120 ( .A(n1287), .B(n1286), .S(n2126), .Z(n1288) );
  MUX2_X1 U6121 ( .A(\mem[250][5] ), .B(\mem[251][5] ), .S(n2155), .Z(n1289)
         );
  MUX2_X1 U6122 ( .A(\mem[248][5] ), .B(\mem[249][5] ), .S(n2155), .Z(n1290)
         );
  MUX2_X1 U6123 ( .A(n1290), .B(n1289), .S(n2126), .Z(n1291) );
  MUX2_X1 U6124 ( .A(n1291), .B(n1288), .S(n2079), .Z(n1292) );
  MUX2_X1 U6125 ( .A(\mem[246][5] ), .B(\mem[247][5] ), .S(n2155), .Z(n1293)
         );
  MUX2_X1 U6126 ( .A(\mem[244][5] ), .B(\mem[245][5] ), .S(n2155), .Z(n1294)
         );
  MUX2_X1 U6127 ( .A(n1294), .B(n1293), .S(n2126), .Z(n1295) );
  MUX2_X1 U6128 ( .A(\mem[242][5] ), .B(\mem[243][5] ), .S(n2155), .Z(n1296)
         );
  MUX2_X1 U6129 ( .A(\mem[240][5] ), .B(\mem[241][5] ), .S(n2155), .Z(n1297)
         );
  MUX2_X1 U6130 ( .A(n1297), .B(n1296), .S(n2126), .Z(n1298) );
  MUX2_X1 U6131 ( .A(n1298), .B(n1295), .S(n2075), .Z(n1299) );
  MUX2_X1 U6132 ( .A(n1299), .B(n1292), .S(n2064), .Z(n1300) );
  MUX2_X1 U6133 ( .A(\mem[238][5] ), .B(\mem[239][5] ), .S(n2155), .Z(n1301)
         );
  MUX2_X1 U6134 ( .A(\mem[236][5] ), .B(\mem[237][5] ), .S(n2155), .Z(n1302)
         );
  MUX2_X1 U6135 ( .A(n1302), .B(n1301), .S(n2126), .Z(n1303) );
  MUX2_X1 U6136 ( .A(\mem[234][5] ), .B(\mem[235][5] ), .S(n2155), .Z(n1304)
         );
  MUX2_X1 U6137 ( .A(\mem[232][5] ), .B(\mem[233][5] ), .S(n2206), .Z(n1305)
         );
  MUX2_X1 U6138 ( .A(n1305), .B(n1304), .S(n2126), .Z(n1306) );
  MUX2_X1 U6139 ( .A(n1306), .B(n1303), .S(n2089), .Z(n1307) );
  MUX2_X1 U6140 ( .A(\mem[230][5] ), .B(\mem[231][5] ), .S(n1), .Z(n1308) );
  MUX2_X1 U6141 ( .A(\mem[228][5] ), .B(\mem[229][5] ), .S(n2144), .Z(n1309)
         );
  MUX2_X1 U6142 ( .A(n1309), .B(n1308), .S(n2126), .Z(n1310) );
  MUX2_X1 U6143 ( .A(\mem[226][5] ), .B(\mem[227][5] ), .S(n2196), .Z(n1311)
         );
  MUX2_X1 U6144 ( .A(\mem[224][5] ), .B(\mem[225][5] ), .S(n1), .Z(n1312) );
  MUX2_X1 U6145 ( .A(n1312), .B(n1311), .S(n2126), .Z(n1313) );
  MUX2_X1 U6146 ( .A(n1313), .B(n1310), .S(n2088), .Z(n1314) );
  MUX2_X1 U6147 ( .A(n1314), .B(n1307), .S(n2064), .Z(n1315) );
  MUX2_X1 U6148 ( .A(n1315), .B(n1300), .S(n2055), .Z(n1316) );
  MUX2_X1 U6149 ( .A(\mem[222][5] ), .B(\mem[223][5] ), .S(n2205), .Z(n1317)
         );
  MUX2_X1 U6150 ( .A(\mem[220][5] ), .B(\mem[221][5] ), .S(n2172), .Z(n1318)
         );
  MUX2_X1 U6151 ( .A(n1318), .B(n1317), .S(n2126), .Z(n1319) );
  MUX2_X1 U6152 ( .A(\mem[218][5] ), .B(\mem[219][5] ), .S(n2175), .Z(n1320)
         );
  MUX2_X1 U6153 ( .A(\mem[216][5] ), .B(\mem[217][5] ), .S(n2205), .Z(n1321)
         );
  MUX2_X1 U6154 ( .A(n1321), .B(n1320), .S(n2126), .Z(n1322) );
  MUX2_X1 U6155 ( .A(n1322), .B(n1319), .S(n2088), .Z(n1323) );
  MUX2_X1 U6156 ( .A(\mem[214][5] ), .B(\mem[215][5] ), .S(n2170), .Z(n1324)
         );
  MUX2_X1 U6157 ( .A(\mem[212][5] ), .B(\mem[213][5] ), .S(n2212), .Z(n1325)
         );
  MUX2_X1 U6158 ( .A(n1325), .B(n1324), .S(n2126), .Z(n1326) );
  MUX2_X1 U6159 ( .A(\mem[210][5] ), .B(\mem[211][5] ), .S(n2206), .Z(n1327)
         );
  MUX2_X1 U6160 ( .A(\mem[208][5] ), .B(\mem[209][5] ), .S(n1), .Z(n1328) );
  MUX2_X1 U6161 ( .A(n1328), .B(n1327), .S(n2126), .Z(n1329) );
  MUX2_X1 U6162 ( .A(n1329), .B(n1326), .S(n2088), .Z(n1330) );
  MUX2_X1 U6163 ( .A(n1330), .B(n1323), .S(n2064), .Z(n1331) );
  MUX2_X1 U6164 ( .A(\mem[206][5] ), .B(\mem[207][5] ), .S(n2163), .Z(n1332)
         );
  MUX2_X1 U6165 ( .A(\mem[204][5] ), .B(\mem[205][5] ), .S(n2140), .Z(n1333)
         );
  MUX2_X1 U6166 ( .A(n1333), .B(n1332), .S(n2127), .Z(n1334) );
  MUX2_X1 U6167 ( .A(\mem[202][5] ), .B(\mem[203][5] ), .S(n2140), .Z(n1335)
         );
  MUX2_X1 U6168 ( .A(\mem[200][5] ), .B(\mem[201][5] ), .S(n2177), .Z(n1336)
         );
  MUX2_X1 U6169 ( .A(n1336), .B(n1335), .S(n2127), .Z(n1337) );
  MUX2_X1 U6170 ( .A(n1337), .B(n1334), .S(n2088), .Z(n1338) );
  MUX2_X1 U6171 ( .A(\mem[198][5] ), .B(\mem[199][5] ), .S(n2140), .Z(n1339)
         );
  MUX2_X1 U6172 ( .A(\mem[196][5] ), .B(\mem[197][5] ), .S(n2172), .Z(n1340)
         );
  MUX2_X1 U6173 ( .A(n1340), .B(n1339), .S(n2127), .Z(n1341) );
  MUX2_X1 U6174 ( .A(\mem[194][5] ), .B(\mem[195][5] ), .S(n2140), .Z(n1342)
         );
  MUX2_X1 U6175 ( .A(\mem[192][5] ), .B(\mem[193][5] ), .S(n2190), .Z(n1343)
         );
  MUX2_X1 U6176 ( .A(n1343), .B(n1342), .S(n2127), .Z(n1344) );
  MUX2_X1 U6177 ( .A(n1344), .B(n1341), .S(n2088), .Z(n1345) );
  MUX2_X1 U6178 ( .A(n1345), .B(n1338), .S(n2064), .Z(n1346) );
  MUX2_X1 U6179 ( .A(n1346), .B(n1331), .S(n2055), .Z(n1347) );
  MUX2_X1 U6180 ( .A(n1347), .B(n1316), .S(n2050), .Z(n1348) );
  MUX2_X1 U6181 ( .A(\mem[190][5] ), .B(\mem[191][5] ), .S(n2164), .Z(n1349)
         );
  MUX2_X1 U6182 ( .A(\mem[188][5] ), .B(\mem[189][5] ), .S(n2140), .Z(n1350)
         );
  MUX2_X1 U6183 ( .A(n1350), .B(n1349), .S(n2127), .Z(n1351) );
  MUX2_X1 U6184 ( .A(\mem[186][5] ), .B(\mem[187][5] ), .S(n8), .Z(n1352) );
  MUX2_X1 U6185 ( .A(\mem[184][5] ), .B(\mem[185][5] ), .S(n2140), .Z(n1353)
         );
  MUX2_X1 U6186 ( .A(n1353), .B(n1352), .S(n2127), .Z(n1354) );
  MUX2_X1 U6187 ( .A(n1354), .B(n1351), .S(n2076), .Z(n1355) );
  MUX2_X1 U6188 ( .A(\mem[182][5] ), .B(\mem[183][5] ), .S(n2189), .Z(n1356)
         );
  MUX2_X1 U6189 ( .A(\mem[180][5] ), .B(\mem[181][5] ), .S(n2190), .Z(n1357)
         );
  MUX2_X1 U6190 ( .A(n1357), .B(n1356), .S(n2127), .Z(n1358) );
  MUX2_X1 U6191 ( .A(\mem[178][5] ), .B(\mem[179][5] ), .S(n2150), .Z(n1359)
         );
  MUX2_X1 U6192 ( .A(\mem[176][5] ), .B(\mem[177][5] ), .S(n2204), .Z(n1360)
         );
  MUX2_X1 U6193 ( .A(n1360), .B(n1359), .S(n2127), .Z(n1361) );
  MUX2_X1 U6194 ( .A(n1361), .B(n1358), .S(n2089), .Z(n1362) );
  MUX2_X1 U6195 ( .A(n1362), .B(n1355), .S(n2064), .Z(n1363) );
  MUX2_X1 U6196 ( .A(\mem[174][5] ), .B(\mem[175][5] ), .S(n2140), .Z(n1364)
         );
  MUX2_X1 U6197 ( .A(\mem[172][5] ), .B(\mem[173][5] ), .S(n2190), .Z(n1365)
         );
  MUX2_X1 U6198 ( .A(n1365), .B(n1364), .S(n2127), .Z(n1366) );
  MUX2_X1 U6199 ( .A(\mem[170][5] ), .B(\mem[171][5] ), .S(n2151), .Z(n1367)
         );
  MUX2_X1 U6200 ( .A(\mem[168][5] ), .B(\mem[169][5] ), .S(n2188), .Z(n1368)
         );
  MUX2_X1 U6201 ( .A(n1368), .B(n1367), .S(n2127), .Z(n1369) );
  MUX2_X1 U6202 ( .A(n1369), .B(n1366), .S(n2089), .Z(n1370) );
  MUX2_X1 U6203 ( .A(\mem[166][5] ), .B(\mem[167][5] ), .S(n2188), .Z(n1371)
         );
  MUX2_X1 U6204 ( .A(\mem[164][5] ), .B(\mem[165][5] ), .S(n2160), .Z(n1372)
         );
  MUX2_X1 U6205 ( .A(n1372), .B(n1371), .S(n2127), .Z(n1373) );
  MUX2_X1 U6206 ( .A(\mem[162][5] ), .B(\mem[163][5] ), .S(n2207), .Z(n1374)
         );
  MUX2_X1 U6207 ( .A(\mem[160][5] ), .B(\mem[161][5] ), .S(n2197), .Z(n1375)
         );
  MUX2_X1 U6208 ( .A(n1375), .B(n1374), .S(n2127), .Z(n1376) );
  MUX2_X1 U6209 ( .A(n1376), .B(n1373), .S(n2089), .Z(n1377) );
  MUX2_X1 U6210 ( .A(n1377), .B(n1370), .S(n2064), .Z(n1378) );
  MUX2_X1 U6211 ( .A(n1378), .B(n1363), .S(n2055), .Z(n1379) );
  MUX2_X1 U6212 ( .A(\mem[158][5] ), .B(\mem[159][5] ), .S(n2177), .Z(n1380)
         );
  MUX2_X1 U6213 ( .A(\mem[156][5] ), .B(\mem[157][5] ), .S(n2153), .Z(n1381)
         );
  MUX2_X1 U6214 ( .A(n1381), .B(n1380), .S(n2128), .Z(n1382) );
  MUX2_X1 U6215 ( .A(\mem[154][5] ), .B(\mem[155][5] ), .S(n4), .Z(n1383) );
  MUX2_X1 U6216 ( .A(\mem[152][5] ), .B(\mem[153][5] ), .S(n2152), .Z(n1384)
         );
  MUX2_X1 U6217 ( .A(n1384), .B(n1383), .S(n2128), .Z(n1385) );
  MUX2_X1 U6218 ( .A(n1385), .B(n1382), .S(n2079), .Z(n1386) );
  MUX2_X1 U6219 ( .A(\mem[150][5] ), .B(\mem[151][5] ), .S(n2192), .Z(n1387)
         );
  MUX2_X1 U6220 ( .A(\mem[148][5] ), .B(\mem[149][5] ), .S(n2177), .Z(n1388)
         );
  MUX2_X1 U6221 ( .A(n1388), .B(n1387), .S(n2128), .Z(n1389) );
  MUX2_X1 U6222 ( .A(\mem[146][5] ), .B(\mem[147][5] ), .S(n2153), .Z(n1390)
         );
  MUX2_X1 U6223 ( .A(\mem[144][5] ), .B(\mem[145][5] ), .S(n2150), .Z(n1391)
         );
  MUX2_X1 U6224 ( .A(n1391), .B(n1390), .S(n2128), .Z(n1392) );
  MUX2_X1 U6225 ( .A(n1392), .B(n1389), .S(n2082), .Z(n1393) );
  MUX2_X1 U6226 ( .A(n1393), .B(n1386), .S(n2064), .Z(n1394) );
  MUX2_X1 U6227 ( .A(\mem[142][5] ), .B(\mem[143][5] ), .S(n2177), .Z(n1395)
         );
  MUX2_X1 U6228 ( .A(\mem[140][5] ), .B(\mem[141][5] ), .S(n2151), .Z(n1396)
         );
  MUX2_X1 U6229 ( .A(n1396), .B(n1395), .S(n2128), .Z(n1397) );
  MUX2_X1 U6230 ( .A(\mem[138][5] ), .B(\mem[139][5] ), .S(n2210), .Z(n1398)
         );
  MUX2_X1 U6231 ( .A(\mem[136][5] ), .B(\mem[137][5] ), .S(n2214), .Z(n1399)
         );
  MUX2_X1 U6232 ( .A(n1399), .B(n1398), .S(n2128), .Z(n1400) );
  MUX2_X1 U6233 ( .A(n1400), .B(n1397), .S(n2076), .Z(n1401) );
  MUX2_X1 U6234 ( .A(\mem[134][5] ), .B(\mem[135][5] ), .S(n2154), .Z(n1402)
         );
  MUX2_X1 U6235 ( .A(\mem[132][5] ), .B(\mem[133][5] ), .S(n2154), .Z(n1403)
         );
  MUX2_X1 U6236 ( .A(n1403), .B(n1402), .S(n2128), .Z(n1404) );
  MUX2_X1 U6237 ( .A(\mem[130][5] ), .B(\mem[131][5] ), .S(n2154), .Z(n1405)
         );
  MUX2_X1 U6238 ( .A(\mem[128][5] ), .B(\mem[129][5] ), .S(n2197), .Z(n1406)
         );
  MUX2_X1 U6239 ( .A(n1406), .B(n1405), .S(n2128), .Z(n1407) );
  MUX2_X1 U6240 ( .A(n1407), .B(n1404), .S(n2089), .Z(n1408) );
  MUX2_X1 U6241 ( .A(n1408), .B(n1401), .S(n2064), .Z(n1409) );
  MUX2_X1 U6242 ( .A(n1409), .B(n1394), .S(n2055), .Z(n1410) );
  MUX2_X1 U6243 ( .A(n1410), .B(n1379), .S(n2050), .Z(n1411) );
  MUX2_X1 U6244 ( .A(n1411), .B(n1348), .S(N24), .Z(n1412) );
  MUX2_X1 U6245 ( .A(\mem[126][5] ), .B(\mem[127][5] ), .S(n2154), .Z(n1413)
         );
  MUX2_X1 U6246 ( .A(\mem[124][5] ), .B(\mem[125][5] ), .S(n2154), .Z(n1414)
         );
  MUX2_X1 U6247 ( .A(n1414), .B(n1413), .S(n2128), .Z(n1415) );
  MUX2_X1 U6248 ( .A(\mem[122][5] ), .B(\mem[123][5] ), .S(n2154), .Z(n1416)
         );
  MUX2_X1 U6249 ( .A(\mem[120][5] ), .B(\mem[121][5] ), .S(n2154), .Z(n1417)
         );
  MUX2_X1 U6250 ( .A(n1417), .B(n1416), .S(n2128), .Z(n1418) );
  MUX2_X1 U6251 ( .A(n1418), .B(n1415), .S(n2070), .Z(n1419) );
  MUX2_X1 U6252 ( .A(\mem[118][5] ), .B(\mem[119][5] ), .S(n2154), .Z(n1420)
         );
  MUX2_X1 U6253 ( .A(\mem[116][5] ), .B(\mem[117][5] ), .S(n2154), .Z(n1421)
         );
  MUX2_X1 U6254 ( .A(n1421), .B(n1420), .S(n2128), .Z(n1422) );
  MUX2_X1 U6255 ( .A(\mem[114][5] ), .B(\mem[115][5] ), .S(n2154), .Z(n1423)
         );
  MUX2_X1 U6256 ( .A(\mem[112][5] ), .B(\mem[113][5] ), .S(n2154), .Z(n1424)
         );
  MUX2_X1 U6257 ( .A(n1424), .B(n1423), .S(n2128), .Z(n1425) );
  MUX2_X1 U6258 ( .A(n1425), .B(n1422), .S(n2070), .Z(n1426) );
  MUX2_X1 U6259 ( .A(n1426), .B(n1419), .S(n2064), .Z(n1427) );
  MUX2_X1 U6260 ( .A(\mem[110][5] ), .B(\mem[111][5] ), .S(n2198), .Z(n1428)
         );
  MUX2_X1 U6261 ( .A(\mem[108][5] ), .B(\mem[109][5] ), .S(n2198), .Z(n1429)
         );
  MUX2_X1 U6262 ( .A(n1429), .B(n1428), .S(n2100), .Z(n1430) );
  MUX2_X1 U6263 ( .A(\mem[106][5] ), .B(\mem[107][5] ), .S(n2198), .Z(n1431)
         );
  MUX2_X1 U6264 ( .A(\mem[104][5] ), .B(\mem[105][5] ), .S(n2163), .Z(n1432)
         );
  MUX2_X1 U6265 ( .A(n1432), .B(n1431), .S(n2110), .Z(n1433) );
  MUX2_X1 U6266 ( .A(n1433), .B(n1430), .S(n2070), .Z(n1434) );
  MUX2_X1 U6267 ( .A(\mem[102][5] ), .B(\mem[103][5] ), .S(n2198), .Z(n1435)
         );
  MUX2_X1 U6268 ( .A(\mem[100][5] ), .B(\mem[101][5] ), .S(n2198), .Z(n1436)
         );
  MUX2_X1 U6269 ( .A(n1436), .B(n1435), .S(n2092), .Z(n1437) );
  MUX2_X1 U6270 ( .A(\mem[98][5] ), .B(\mem[99][5] ), .S(n2201), .Z(n1438) );
  MUX2_X1 U6271 ( .A(\mem[96][5] ), .B(\mem[97][5] ), .S(n2197), .Z(n1439) );
  MUX2_X1 U6272 ( .A(n1439), .B(n1438), .S(n2106), .Z(n1440) );
  MUX2_X1 U6273 ( .A(n1440), .B(n1437), .S(n2070), .Z(n1441) );
  MUX2_X1 U6274 ( .A(n1441), .B(n1434), .S(n2064), .Z(n1442) );
  MUX2_X1 U6275 ( .A(n1442), .B(n1427), .S(n2055), .Z(n1443) );
  MUX2_X1 U6276 ( .A(\mem[94][5] ), .B(\mem[95][5] ), .S(n2198), .Z(n1444) );
  MUX2_X1 U6277 ( .A(\mem[92][5] ), .B(\mem[93][5] ), .S(n2198), .Z(n1445) );
  MUX2_X1 U6278 ( .A(n1445), .B(n1444), .S(n2129), .Z(n1446) );
  MUX2_X1 U6279 ( .A(\mem[90][5] ), .B(\mem[91][5] ), .S(n2198), .Z(n1447) );
  MUX2_X1 U6280 ( .A(\mem[88][5] ), .B(\mem[89][5] ), .S(n2165), .Z(n1448) );
  MUX2_X1 U6281 ( .A(n1448), .B(n1447), .S(n2093), .Z(n1449) );
  MUX2_X1 U6282 ( .A(n1449), .B(n1446), .S(n2070), .Z(n1450) );
  MUX2_X1 U6283 ( .A(\mem[86][5] ), .B(\mem[87][5] ), .S(n2198), .Z(n1451) );
  MUX2_X1 U6284 ( .A(\mem[84][5] ), .B(\mem[85][5] ), .S(n2198), .Z(n1452) );
  MUX2_X1 U6285 ( .A(n1452), .B(n1451), .S(n2092), .Z(n1453) );
  MUX2_X1 U6286 ( .A(\mem[82][5] ), .B(\mem[83][5] ), .S(n2198), .Z(n1454) );
  MUX2_X1 U6287 ( .A(\mem[80][5] ), .B(\mem[81][5] ), .S(n2198), .Z(n1455) );
  MUX2_X1 U6288 ( .A(n1455), .B(n1454), .S(n2109), .Z(n1456) );
  MUX2_X1 U6289 ( .A(n1456), .B(n1453), .S(n2090), .Z(n1457) );
  MUX2_X1 U6290 ( .A(n1457), .B(n1450), .S(n2064), .Z(n1458) );
  MUX2_X1 U6291 ( .A(\mem[78][5] ), .B(\mem[79][5] ), .S(n2198), .Z(n1459) );
  MUX2_X1 U6292 ( .A(\mem[76][5] ), .B(\mem[77][5] ), .S(n2198), .Z(n1460) );
  MUX2_X1 U6293 ( .A(n1460), .B(n1459), .S(n2113), .Z(n1461) );
  MUX2_X1 U6294 ( .A(\mem[74][5] ), .B(\mem[75][5] ), .S(n2198), .Z(n1462) );
  MUX2_X1 U6295 ( .A(\mem[72][5] ), .B(\mem[73][5] ), .S(n2198), .Z(n1463) );
  MUX2_X1 U6296 ( .A(n1463), .B(n1462), .S(n2108), .Z(n1464) );
  MUX2_X1 U6297 ( .A(n1464), .B(n1461), .S(n2070), .Z(n1465) );
  MUX2_X1 U6298 ( .A(\mem[70][5] ), .B(\mem[71][5] ), .S(n2198), .Z(n1466) );
  MUX2_X1 U6299 ( .A(\mem[68][5] ), .B(\mem[69][5] ), .S(n2198), .Z(n1467) );
  MUX2_X1 U6300 ( .A(n1467), .B(n1466), .S(n2107), .Z(n1468) );
  MUX2_X1 U6301 ( .A(\mem[66][5] ), .B(\mem[67][5] ), .S(n2198), .Z(n1469) );
  MUX2_X1 U6302 ( .A(\mem[64][5] ), .B(\mem[65][5] ), .S(n2198), .Z(n1470) );
  MUX2_X1 U6303 ( .A(n1470), .B(n1469), .S(n2097), .Z(n1471) );
  MUX2_X1 U6304 ( .A(n1471), .B(n1468), .S(n2070), .Z(n1472) );
  MUX2_X1 U6305 ( .A(n1472), .B(n1465), .S(n2064), .Z(n1473) );
  MUX2_X1 U6306 ( .A(n1473), .B(n1458), .S(n2055), .Z(n1474) );
  MUX2_X1 U6307 ( .A(n1474), .B(n1443), .S(n2050), .Z(n1475) );
  MUX2_X1 U6308 ( .A(\mem[62][5] ), .B(\mem[63][5] ), .S(n2198), .Z(n1476) );
  MUX2_X1 U6309 ( .A(\mem[60][5] ), .B(\mem[61][5] ), .S(n2153), .Z(n1477) );
  MUX2_X1 U6310 ( .A(n1477), .B(n1476), .S(n2129), .Z(n1478) );
  MUX2_X1 U6311 ( .A(\mem[58][5] ), .B(\mem[59][5] ), .S(n2178), .Z(n1479) );
  MUX2_X1 U6312 ( .A(\mem[56][5] ), .B(\mem[57][5] ), .S(n2201), .Z(n1480) );
  MUX2_X1 U6313 ( .A(n1480), .B(n1479), .S(n2129), .Z(n1481) );
  MUX2_X1 U6314 ( .A(n1481), .B(n1478), .S(n2091), .Z(n1482) );
  MUX2_X1 U6315 ( .A(\mem[54][5] ), .B(\mem[55][5] ), .S(n8), .Z(n1483) );
  MUX2_X1 U6316 ( .A(\mem[52][5] ), .B(\mem[53][5] ), .S(n2204), .Z(n1484) );
  MUX2_X1 U6317 ( .A(n1484), .B(n1483), .S(n2129), .Z(n1485) );
  MUX2_X1 U6318 ( .A(\mem[50][5] ), .B(\mem[51][5] ), .S(n2176), .Z(n1486) );
  MUX2_X1 U6319 ( .A(\mem[48][5] ), .B(\mem[49][5] ), .S(n1), .Z(n1487) );
  MUX2_X1 U6320 ( .A(n1487), .B(n1486), .S(n2129), .Z(n1488) );
  MUX2_X1 U6321 ( .A(n1488), .B(n1485), .S(n2087), .Z(n1489) );
  MUX2_X1 U6322 ( .A(n1489), .B(n1482), .S(n2065), .Z(n1490) );
  MUX2_X1 U6323 ( .A(\mem[46][5] ), .B(\mem[47][5] ), .S(n2200), .Z(n1491) );
  MUX2_X1 U6324 ( .A(\mem[44][5] ), .B(\mem[45][5] ), .S(n2201), .Z(n1492) );
  MUX2_X1 U6325 ( .A(n1492), .B(n1491), .S(n2129), .Z(n1493) );
  MUX2_X1 U6326 ( .A(\mem[42][5] ), .B(\mem[43][5] ), .S(n2182), .Z(n1494) );
  MUX2_X1 U6327 ( .A(\mem[40][5] ), .B(\mem[41][5] ), .S(n7), .Z(n1495) );
  MUX2_X1 U6328 ( .A(n1495), .B(n1494), .S(n2129), .Z(n1496) );
  MUX2_X1 U6329 ( .A(n1496), .B(n1493), .S(n2091), .Z(n1497) );
  MUX2_X1 U6330 ( .A(\mem[38][5] ), .B(\mem[39][5] ), .S(n2214), .Z(n1498) );
  MUX2_X1 U6331 ( .A(\mem[36][5] ), .B(\mem[37][5] ), .S(n2198), .Z(n1499) );
  MUX2_X1 U6332 ( .A(n1499), .B(n1498), .S(n2129), .Z(n1500) );
  MUX2_X1 U6333 ( .A(\mem[34][5] ), .B(\mem[35][5] ), .S(n2140), .Z(n1501) );
  MUX2_X1 U6334 ( .A(\mem[32][5] ), .B(\mem[33][5] ), .S(n2153), .Z(n1502) );
  MUX2_X1 U6335 ( .A(n1502), .B(n1501), .S(n2129), .Z(n1503) );
  MUX2_X1 U6336 ( .A(n1503), .B(n1500), .S(n2087), .Z(n1504) );
  MUX2_X1 U6337 ( .A(n1504), .B(n1497), .S(n2065), .Z(n1505) );
  MUX2_X1 U6338 ( .A(n1505), .B(n1490), .S(n2055), .Z(n1506) );
  MUX2_X1 U6339 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n2213), .Z(n1507) );
  MUX2_X1 U6340 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n2201), .Z(n1508) );
  MUX2_X1 U6341 ( .A(n1508), .B(n1507), .S(n2129), .Z(n1509) );
  MUX2_X1 U6342 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n2137), .Z(n1510) );
  MUX2_X1 U6343 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n2199), .Z(n1511) );
  MUX2_X1 U6344 ( .A(n1511), .B(n1510), .S(n2129), .Z(n1512) );
  MUX2_X1 U6345 ( .A(n1512), .B(n1509), .S(n2089), .Z(n1513) );
  MUX2_X1 U6346 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n2213), .Z(n1514) );
  MUX2_X1 U6347 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n2201), .Z(n1515) );
  MUX2_X1 U6348 ( .A(n1515), .B(n1514), .S(n2129), .Z(n1516) );
  MUX2_X1 U6349 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n2182), .Z(n1517) );
  MUX2_X1 U6350 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n2184), .Z(n1518) );
  MUX2_X1 U6351 ( .A(n1518), .B(n1517), .S(n2129), .Z(n1519) );
  MUX2_X1 U6352 ( .A(n1519), .B(n1516), .S(n2073), .Z(n1520) );
  MUX2_X1 U6353 ( .A(n1520), .B(n1513), .S(n2065), .Z(n1521) );
  MUX2_X1 U6354 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n2199), .Z(n1522) );
  MUX2_X1 U6355 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n2199), .Z(n1523) );
  MUX2_X1 U6356 ( .A(n1523), .B(n1522), .S(n2124), .Z(n1524) );
  MUX2_X1 U6357 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n2199), .Z(n1525) );
  MUX2_X1 U6358 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n2199), .Z(n1526) );
  MUX2_X1 U6359 ( .A(n1526), .B(n1525), .S(n2128), .Z(n1527) );
  MUX2_X1 U6360 ( .A(n1527), .B(n1524), .S(n2089), .Z(n1528) );
  MUX2_X1 U6361 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n2199), .Z(n1529) );
  MUX2_X1 U6362 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n2199), .Z(n1530) );
  MUX2_X1 U6363 ( .A(n1530), .B(n1529), .S(n2123), .Z(n1531) );
  MUX2_X1 U6364 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n2199), .Z(n1532) );
  MUX2_X1 U6365 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n2199), .Z(n1533) );
  MUX2_X1 U6366 ( .A(n1533), .B(n1532), .S(n2118), .Z(n1534) );
  MUX2_X1 U6367 ( .A(n1534), .B(n1531), .S(n2072), .Z(n1535) );
  MUX2_X1 U6368 ( .A(n1535), .B(n1528), .S(n2065), .Z(n1536) );
  MUX2_X1 U6369 ( .A(n1536), .B(n1521), .S(n2055), .Z(n1537) );
  MUX2_X1 U6370 ( .A(n1537), .B(n1506), .S(n2050), .Z(n1538) );
  MUX2_X1 U6371 ( .A(n1538), .B(n1475), .S(N24), .Z(n1539) );
  MUX2_X1 U6372 ( .A(\mem[254][6] ), .B(\mem[255][6] ), .S(n2199), .Z(n1540)
         );
  MUX2_X1 U6373 ( .A(\mem[252][6] ), .B(\mem[253][6] ), .S(n2199), .Z(n1541)
         );
  MUX2_X1 U6374 ( .A(n1541), .B(n1540), .S(n2114), .Z(n1542) );
  MUX2_X1 U6375 ( .A(\mem[250][6] ), .B(\mem[251][6] ), .S(n2199), .Z(n1543)
         );
  MUX2_X1 U6376 ( .A(\mem[248][6] ), .B(\mem[249][6] ), .S(n2199), .Z(n1544)
         );
  MUX2_X1 U6377 ( .A(n1544), .B(n1543), .S(n2113), .Z(n1545) );
  MUX2_X1 U6378 ( .A(n1545), .B(n1542), .S(n2071), .Z(n1546) );
  MUX2_X1 U6379 ( .A(\mem[246][6] ), .B(\mem[247][6] ), .S(n2140), .Z(n1547)
         );
  MUX2_X1 U6380 ( .A(\mem[244][6] ), .B(\mem[245][6] ), .S(n2191), .Z(n1548)
         );
  MUX2_X1 U6381 ( .A(n1548), .B(n1547), .S(n2132), .Z(n1549) );
  MUX2_X1 U6382 ( .A(\mem[242][6] ), .B(\mem[243][6] ), .S(n2188), .Z(n1550)
         );
  MUX2_X1 U6383 ( .A(\mem[240][6] ), .B(\mem[241][6] ), .S(n2197), .Z(n1551)
         );
  MUX2_X1 U6384 ( .A(n1551), .B(n1550), .S(n2117), .Z(n1552) );
  MUX2_X1 U6385 ( .A(n1552), .B(n1549), .S(n2088), .Z(n1553) );
  MUX2_X1 U6386 ( .A(n1553), .B(n1546), .S(n2065), .Z(n1554) );
  MUX2_X1 U6387 ( .A(\mem[238][6] ), .B(\mem[239][6] ), .S(n2197), .Z(n1555)
         );
  MUX2_X1 U6388 ( .A(\mem[236][6] ), .B(\mem[237][6] ), .S(n2205), .Z(n1556)
         );
  MUX2_X1 U6389 ( .A(n1556), .B(n1555), .S(n2110), .Z(n1557) );
  MUX2_X1 U6390 ( .A(\mem[234][6] ), .B(\mem[235][6] ), .S(n2207), .Z(n1558)
         );
  MUX2_X1 U6391 ( .A(\mem[232][6] ), .B(\mem[233][6] ), .S(n2140), .Z(n1559)
         );
  MUX2_X1 U6392 ( .A(n1559), .B(n1558), .S(n2121), .Z(n1560) );
  MUX2_X1 U6393 ( .A(n1560), .B(n1557), .S(n2089), .Z(n1561) );
  MUX2_X1 U6394 ( .A(\mem[230][6] ), .B(\mem[231][6] ), .S(n2197), .Z(n1562)
         );
  MUX2_X1 U6395 ( .A(\mem[228][6] ), .B(\mem[229][6] ), .S(n2152), .Z(n1563)
         );
  MUX2_X1 U6396 ( .A(n1563), .B(n1562), .S(n2127), .Z(n1564) );
  MUX2_X1 U6397 ( .A(\mem[226][6] ), .B(\mem[227][6] ), .S(n2191), .Z(n1565)
         );
  MUX2_X1 U6398 ( .A(\mem[224][6] ), .B(\mem[225][6] ), .S(n2211), .Z(n1566)
         );
  MUX2_X1 U6399 ( .A(n1566), .B(n1565), .S(n2116), .Z(n1567) );
  MUX2_X1 U6400 ( .A(n1567), .B(n1564), .S(n2083), .Z(n1568) );
  MUX2_X1 U6401 ( .A(n1568), .B(n1561), .S(n2065), .Z(n1569) );
  MUX2_X1 U6402 ( .A(n1569), .B(n1554), .S(n2055), .Z(n1570) );
  MUX2_X1 U6403 ( .A(\mem[222][6] ), .B(\mem[223][6] ), .S(n2200), .Z(n1571)
         );
  MUX2_X1 U6404 ( .A(\mem[220][6] ), .B(\mem[221][6] ), .S(n2201), .Z(n1572)
         );
  MUX2_X1 U6405 ( .A(n1572), .B(n1571), .S(n2122), .Z(n1573) );
  MUX2_X1 U6406 ( .A(\mem[218][6] ), .B(\mem[219][6] ), .S(n2183), .Z(n1574)
         );
  MUX2_X1 U6407 ( .A(\mem[216][6] ), .B(\mem[217][6] ), .S(n2201), .Z(n1575)
         );
  MUX2_X1 U6408 ( .A(n1575), .B(n1574), .S(n2100), .Z(n1576) );
  MUX2_X1 U6409 ( .A(n1576), .B(n1573), .S(n2070), .Z(n1577) );
  MUX2_X1 U6410 ( .A(\mem[214][6] ), .B(\mem[215][6] ), .S(n2189), .Z(n1578)
         );
  MUX2_X1 U6411 ( .A(\mem[212][6] ), .B(\mem[213][6] ), .S(n2201), .Z(n1579)
         );
  MUX2_X1 U6412 ( .A(n1579), .B(n1578), .S(n2116), .Z(n1580) );
  MUX2_X1 U6413 ( .A(\mem[210][6] ), .B(\mem[211][6] ), .S(n2180), .Z(n1581)
         );
  MUX2_X1 U6414 ( .A(\mem[208][6] ), .B(\mem[209][6] ), .S(n2190), .Z(n1582)
         );
  MUX2_X1 U6415 ( .A(n1582), .B(n1581), .S(n2129), .Z(n1583) );
  MUX2_X1 U6416 ( .A(n1583), .B(n1580), .S(n2089), .Z(n1584) );
  MUX2_X1 U6417 ( .A(n1584), .B(n1577), .S(n2065), .Z(n1585) );
  MUX2_X1 U6418 ( .A(\mem[206][6] ), .B(\mem[207][6] ), .S(n2140), .Z(n1586)
         );
  MUX2_X1 U6419 ( .A(\mem[204][6] ), .B(\mem[205][6] ), .S(n2189), .Z(n1587)
         );
  MUX2_X1 U6420 ( .A(n1587), .B(n1586), .S(n2121), .Z(n1588) );
  MUX2_X1 U6421 ( .A(\mem[202][6] ), .B(\mem[203][6] ), .S(n2181), .Z(n1589)
         );
  MUX2_X1 U6422 ( .A(\mem[200][6] ), .B(\mem[201][6] ), .S(n1), .Z(n1590) );
  MUX2_X1 U6423 ( .A(n1590), .B(n1589), .S(n2135), .Z(n1591) );
  MUX2_X1 U6424 ( .A(n1591), .B(n1588), .S(n2078), .Z(n1592) );
  MUX2_X1 U6425 ( .A(\mem[198][6] ), .B(\mem[199][6] ), .S(n2140), .Z(n1593)
         );
  MUX2_X1 U6426 ( .A(\mem[196][6] ), .B(\mem[197][6] ), .S(n2200), .Z(n1594)
         );
  MUX2_X1 U6427 ( .A(n1594), .B(n1593), .S(n2092), .Z(n1595) );
  MUX2_X1 U6428 ( .A(\mem[194][6] ), .B(\mem[195][6] ), .S(n2200), .Z(n1596)
         );
  MUX2_X1 U6429 ( .A(\mem[192][6] ), .B(\mem[193][6] ), .S(n2200), .Z(n1597)
         );
  MUX2_X1 U6430 ( .A(n1597), .B(n1596), .S(n2106), .Z(n1598) );
  MUX2_X1 U6431 ( .A(n1598), .B(n1595), .S(n2080), .Z(n1599) );
  MUX2_X1 U6432 ( .A(n1599), .B(n1592), .S(n2065), .Z(n1600) );
  MUX2_X1 U6433 ( .A(n1600), .B(n1585), .S(n2055), .Z(n1601) );
  MUX2_X1 U6434 ( .A(n1601), .B(n1570), .S(n2050), .Z(n1602) );
  MUX2_X1 U6435 ( .A(\mem[190][6] ), .B(\mem[191][6] ), .S(n2200), .Z(n1603)
         );
  MUX2_X1 U6436 ( .A(\mem[188][6] ), .B(\mem[189][6] ), .S(n2201), .Z(n1604)
         );
  MUX2_X1 U6437 ( .A(n1604), .B(n1603), .S(n2126), .Z(n1605) );
  MUX2_X1 U6438 ( .A(\mem[186][6] ), .B(\mem[187][6] ), .S(n2201), .Z(n1606)
         );
  MUX2_X1 U6439 ( .A(\mem[184][6] ), .B(\mem[185][6] ), .S(n2200), .Z(n1607)
         );
  MUX2_X1 U6440 ( .A(n1607), .B(n1606), .S(n2117), .Z(n1608) );
  MUX2_X1 U6441 ( .A(n1608), .B(n1605), .S(n2091), .Z(n1609) );
  MUX2_X1 U6442 ( .A(\mem[182][6] ), .B(\mem[183][6] ), .S(n2200), .Z(n1610)
         );
  MUX2_X1 U6443 ( .A(\mem[180][6] ), .B(\mem[181][6] ), .S(n2200), .Z(n1611)
         );
  MUX2_X1 U6444 ( .A(n1611), .B(n1610), .S(n2127), .Z(n1612) );
  MUX2_X1 U6445 ( .A(\mem[178][6] ), .B(\mem[179][6] ), .S(n2188), .Z(n1613)
         );
  MUX2_X1 U6446 ( .A(\mem[176][6] ), .B(\mem[177][6] ), .S(n2201), .Z(n1614)
         );
  MUX2_X1 U6447 ( .A(n1614), .B(n1613), .S(n2122), .Z(n1615) );
  MUX2_X1 U6448 ( .A(n1615), .B(n1612), .S(n2074), .Z(n1616) );
  MUX2_X1 U6449 ( .A(n1616), .B(n1609), .S(n2065), .Z(n1617) );
  MUX2_X1 U6450 ( .A(\mem[174][6] ), .B(\mem[175][6] ), .S(n2162), .Z(n1618)
         );
  MUX2_X1 U6451 ( .A(\mem[172][6] ), .B(\mem[173][6] ), .S(n2201), .Z(n1619)
         );
  MUX2_X1 U6452 ( .A(n1619), .B(n1618), .S(n2108), .Z(n1620) );
  MUX2_X1 U6453 ( .A(\mem[170][6] ), .B(\mem[171][6] ), .S(n2179), .Z(n1621)
         );
  MUX2_X1 U6454 ( .A(\mem[168][6] ), .B(\mem[169][6] ), .S(n2189), .Z(n1622)
         );
  MUX2_X1 U6455 ( .A(n1622), .B(n1621), .S(n2130), .Z(n1623) );
  MUX2_X1 U6456 ( .A(n1623), .B(n1620), .S(n2077), .Z(n1624) );
  MUX2_X1 U6457 ( .A(\mem[166][6] ), .B(\mem[167][6] ), .S(n2201), .Z(n1625)
         );
  MUX2_X1 U6458 ( .A(\mem[164][6] ), .B(\mem[165][6] ), .S(n2184), .Z(n1626)
         );
  MUX2_X1 U6459 ( .A(n1626), .B(n1625), .S(n2112), .Z(n1627) );
  MUX2_X1 U6460 ( .A(\mem[162][6] ), .B(\mem[163][6] ), .S(n2201), .Z(n1628)
         );
  MUX2_X1 U6461 ( .A(\mem[160][6] ), .B(\mem[161][6] ), .S(n2189), .Z(n1629)
         );
  MUX2_X1 U6462 ( .A(n1629), .B(n1628), .S(n2125), .Z(n1630) );
  MUX2_X1 U6463 ( .A(n1630), .B(n1627), .S(n2081), .Z(n1631) );
  MUX2_X1 U6464 ( .A(n1631), .B(n1624), .S(n2065), .Z(n1632) );
  MUX2_X1 U6465 ( .A(n1632), .B(n1617), .S(n2055), .Z(n1633) );
  MUX2_X1 U6466 ( .A(\mem[158][6] ), .B(\mem[159][6] ), .S(n2200), .Z(n1634)
         );
  MUX2_X1 U6467 ( .A(\mem[156][6] ), .B(\mem[157][6] ), .S(n2197), .Z(n1635)
         );
  MUX2_X1 U6468 ( .A(n1635), .B(n1634), .S(n2099), .Z(n1636) );
  MUX2_X1 U6469 ( .A(\mem[154][6] ), .B(\mem[155][6] ), .S(n2183), .Z(n1637)
         );
  MUX2_X1 U6470 ( .A(\mem[152][6] ), .B(\mem[153][6] ), .S(n2201), .Z(n1638)
         );
  MUX2_X1 U6471 ( .A(n1638), .B(n1637), .S(n2093), .Z(n1639) );
  MUX2_X1 U6472 ( .A(n1639), .B(n1636), .S(n2075), .Z(n1640) );
  MUX2_X1 U6473 ( .A(\mem[150][6] ), .B(\mem[151][6] ), .S(n2188), .Z(n1641)
         );
  MUX2_X1 U6474 ( .A(\mem[148][6] ), .B(\mem[149][6] ), .S(n2197), .Z(n1642)
         );
  MUX2_X1 U6475 ( .A(n1642), .B(n1641), .S(n2111), .Z(n1643) );
  MUX2_X1 U6476 ( .A(\mem[146][6] ), .B(\mem[147][6] ), .S(n2201), .Z(n1644)
         );
  MUX2_X1 U6477 ( .A(\mem[144][6] ), .B(\mem[145][6] ), .S(n2175), .Z(n1645)
         );
  MUX2_X1 U6478 ( .A(n1645), .B(n1644), .S(n2115), .Z(n1646) );
  MUX2_X1 U6479 ( .A(n1646), .B(n1643), .S(n2083), .Z(n1647) );
  MUX2_X1 U6480 ( .A(n1647), .B(n1640), .S(n2065), .Z(n1648) );
  MUX2_X1 U6481 ( .A(\mem[142][6] ), .B(\mem[143][6] ), .S(n2200), .Z(n1649)
         );
  MUX2_X1 U6482 ( .A(\mem[140][6] ), .B(\mem[141][6] ), .S(n2184), .Z(n1650)
         );
  MUX2_X1 U6483 ( .A(n1650), .B(n1649), .S(n2105), .Z(n1651) );
  MUX2_X1 U6484 ( .A(\mem[138][6] ), .B(\mem[139][6] ), .S(n2197), .Z(n1652)
         );
  MUX2_X1 U6485 ( .A(\mem[136][6] ), .B(\mem[137][6] ), .S(n2173), .Z(n1653)
         );
  MUX2_X1 U6486 ( .A(n1653), .B(n1652), .S(n2098), .Z(n1654) );
  MUX2_X1 U6487 ( .A(n1654), .B(n1651), .S(n2091), .Z(n1655) );
  MUX2_X1 U6488 ( .A(\mem[134][6] ), .B(\mem[135][6] ), .S(n2200), .Z(n1656)
         );
  MUX2_X1 U6489 ( .A(\mem[132][6] ), .B(\mem[133][6] ), .S(n2205), .Z(n1657)
         );
  MUX2_X1 U6490 ( .A(n1657), .B(n1656), .S(n2120), .Z(n1658) );
  MUX2_X1 U6491 ( .A(\mem[130][6] ), .B(\mem[131][6] ), .S(n2197), .Z(n1659)
         );
  MUX2_X1 U6492 ( .A(\mem[128][6] ), .B(\mem[129][6] ), .S(n2201), .Z(n1660)
         );
  MUX2_X1 U6493 ( .A(n1660), .B(n1659), .S(n2119), .Z(n1661) );
  MUX2_X1 U6494 ( .A(n1661), .B(n1658), .S(n2087), .Z(n1662) );
  MUX2_X1 U6495 ( .A(n1662), .B(n1655), .S(n2065), .Z(n1663) );
  MUX2_X1 U6496 ( .A(n1663), .B(n1648), .S(n2055), .Z(n1664) );
  MUX2_X1 U6497 ( .A(n1664), .B(n1633), .S(n2050), .Z(n1665) );
  MUX2_X1 U6498 ( .A(n1665), .B(n1602), .S(N24), .Z(n1666) );
  MUX2_X1 U6499 ( .A(\mem[126][6] ), .B(\mem[127][6] ), .S(n2140), .Z(n1667)
         );
  MUX2_X1 U6500 ( .A(\mem[124][6] ), .B(\mem[125][6] ), .S(n2140), .Z(n1668)
         );
  MUX2_X1 U6501 ( .A(n1668), .B(n1667), .S(n2130), .Z(n1669) );
  MUX2_X1 U6502 ( .A(\mem[122][6] ), .B(\mem[123][6] ), .S(n2200), .Z(n1670)
         );
  MUX2_X1 U6503 ( .A(\mem[120][6] ), .B(\mem[121][6] ), .S(n2203), .Z(n1671)
         );
  MUX2_X1 U6504 ( .A(n1671), .B(n1670), .S(n2130), .Z(n1672) );
  MUX2_X1 U6505 ( .A(n1672), .B(n1669), .S(n2070), .Z(n1673) );
  MUX2_X1 U6506 ( .A(\mem[118][6] ), .B(\mem[119][6] ), .S(n2201), .Z(n1674)
         );
  MUX2_X1 U6507 ( .A(\mem[116][6] ), .B(\mem[117][6] ), .S(n2201), .Z(n1675)
         );
  MUX2_X1 U6508 ( .A(n1675), .B(n1674), .S(n2130), .Z(n1676) );
  MUX2_X1 U6509 ( .A(\mem[114][6] ), .B(\mem[115][6] ), .S(n2202), .Z(n1677)
         );
  MUX2_X1 U6510 ( .A(\mem[112][6] ), .B(\mem[113][6] ), .S(n2200), .Z(n1678)
         );
  MUX2_X1 U6511 ( .A(n1678), .B(n1677), .S(n2130), .Z(n1679) );
  MUX2_X1 U6512 ( .A(n1679), .B(n1676), .S(n2081), .Z(n1680) );
  MUX2_X1 U6513 ( .A(n1680), .B(n1673), .S(n2066), .Z(n1681) );
  MUX2_X1 U6514 ( .A(\mem[110][6] ), .B(\mem[111][6] ), .S(n2201), .Z(n1682)
         );
  MUX2_X1 U6515 ( .A(\mem[108][6] ), .B(\mem[109][6] ), .S(n2201), .Z(n1683)
         );
  MUX2_X1 U6516 ( .A(n1683), .B(n1682), .S(n2130), .Z(n1684) );
  MUX2_X1 U6517 ( .A(\mem[106][6] ), .B(\mem[107][6] ), .S(n2201), .Z(n1685)
         );
  MUX2_X1 U6518 ( .A(\mem[104][6] ), .B(\mem[105][6] ), .S(n2201), .Z(n1686)
         );
  MUX2_X1 U6519 ( .A(n1686), .B(n1685), .S(n2130), .Z(n1687) );
  MUX2_X1 U6520 ( .A(n1687), .B(n1684), .S(n2088), .Z(n1688) );
  MUX2_X1 U6521 ( .A(\mem[102][6] ), .B(\mem[103][6] ), .S(n2201), .Z(n1689)
         );
  MUX2_X1 U6522 ( .A(\mem[100][6] ), .B(\mem[101][6] ), .S(n2201), .Z(n1690)
         );
  MUX2_X1 U6523 ( .A(n1690), .B(n1689), .S(n2130), .Z(n1691) );
  MUX2_X1 U6524 ( .A(\mem[98][6] ), .B(\mem[99][6] ), .S(n2200), .Z(n1692) );
  MUX2_X1 U6525 ( .A(\mem[96][6] ), .B(\mem[97][6] ), .S(n2201), .Z(n1693) );
  MUX2_X1 U6526 ( .A(n1693), .B(n1692), .S(n2130), .Z(n1694) );
  MUX2_X1 U6527 ( .A(n1694), .B(n1691), .S(N20), .Z(n1695) );
  MUX2_X1 U6528 ( .A(n1695), .B(n1688), .S(n2066), .Z(n1696) );
  MUX2_X1 U6529 ( .A(n1696), .B(n1681), .S(n2056), .Z(n1697) );
  MUX2_X1 U6530 ( .A(\mem[94][6] ), .B(\mem[95][6] ), .S(n2214), .Z(n1698) );
  MUX2_X1 U6531 ( .A(\mem[92][6] ), .B(\mem[93][6] ), .S(n2183), .Z(n1699) );
  MUX2_X1 U6532 ( .A(n1699), .B(n1698), .S(n2130), .Z(n1700) );
  MUX2_X1 U6533 ( .A(\mem[90][6] ), .B(\mem[91][6] ), .S(n2190), .Z(n1701) );
  MUX2_X1 U6534 ( .A(\mem[88][6] ), .B(\mem[89][6] ), .S(n2190), .Z(n1702) );
  MUX2_X1 U6535 ( .A(n1702), .B(n1701), .S(n2130), .Z(n1703) );
  MUX2_X1 U6536 ( .A(n1703), .B(n1700), .S(N20), .Z(n1704) );
  MUX2_X1 U6537 ( .A(\mem[86][6] ), .B(\mem[87][6] ), .S(n2197), .Z(n1705) );
  MUX2_X1 U6538 ( .A(\mem[84][6] ), .B(\mem[85][6] ), .S(n2201), .Z(n1706) );
  MUX2_X1 U6539 ( .A(n1706), .B(n1705), .S(n2130), .Z(n1707) );
  MUX2_X1 U6540 ( .A(\mem[82][6] ), .B(\mem[83][6] ), .S(n2207), .Z(n1708) );
  MUX2_X1 U6541 ( .A(\mem[80][6] ), .B(\mem[81][6] ), .S(n2188), .Z(n1709) );
  MUX2_X1 U6542 ( .A(n1709), .B(n1708), .S(n2130), .Z(n1710) );
  MUX2_X1 U6543 ( .A(n1710), .B(n1707), .S(N20), .Z(n1711) );
  MUX2_X1 U6544 ( .A(n1711), .B(n1704), .S(n2066), .Z(n1712) );
  MUX2_X1 U6545 ( .A(\mem[78][6] ), .B(\mem[79][6] ), .S(n2202), .Z(n1713) );
  MUX2_X1 U6546 ( .A(\mem[76][6] ), .B(\mem[77][6] ), .S(n2202), .Z(n1714) );
  MUX2_X1 U6547 ( .A(n1714), .B(n1713), .S(n2106), .Z(n1715) );
  MUX2_X1 U6548 ( .A(\mem[74][6] ), .B(\mem[75][6] ), .S(n2202), .Z(n1716) );
  MUX2_X1 U6549 ( .A(\mem[72][6] ), .B(\mem[73][6] ), .S(n2202), .Z(n1717) );
  MUX2_X1 U6550 ( .A(n1717), .B(n1716), .S(n2131), .Z(n1718) );
  MUX2_X1 U6551 ( .A(n1718), .B(n1715), .S(N20), .Z(n1719) );
  MUX2_X1 U6552 ( .A(\mem[70][6] ), .B(\mem[71][6] ), .S(n2202), .Z(n1720) );
  MUX2_X1 U6553 ( .A(\mem[68][6] ), .B(\mem[69][6] ), .S(n2202), .Z(n1721) );
  MUX2_X1 U6554 ( .A(n1721), .B(n1720), .S(n2107), .Z(n1722) );
  MUX2_X1 U6555 ( .A(\mem[66][6] ), .B(\mem[67][6] ), .S(n2202), .Z(n1723) );
  MUX2_X1 U6556 ( .A(\mem[64][6] ), .B(\mem[65][6] ), .S(n2202), .Z(n1724) );
  MUX2_X1 U6557 ( .A(n1724), .B(n1723), .S(n2132), .Z(n1725) );
  MUX2_X1 U6558 ( .A(n1725), .B(n1722), .S(N20), .Z(n1726) );
  MUX2_X1 U6559 ( .A(n1726), .B(n1719), .S(n2066), .Z(n1727) );
  MUX2_X1 U6560 ( .A(n1728), .B(n1697), .S(n2050), .Z(n1729) );
  MUX2_X1 U6561 ( .A(\mem[62][6] ), .B(\mem[63][6] ), .S(n2202), .Z(n1730) );
  MUX2_X1 U6562 ( .A(\mem[60][6] ), .B(\mem[61][6] ), .S(n2202), .Z(n1731) );
  MUX2_X1 U6563 ( .A(n1731), .B(n1730), .S(n2092), .Z(n1732) );
  MUX2_X1 U6564 ( .A(\mem[58][6] ), .B(\mem[59][6] ), .S(n2202), .Z(n1733) );
  MUX2_X1 U6565 ( .A(\mem[56][6] ), .B(\mem[57][6] ), .S(n2202), .Z(n1734) );
  MUX2_X1 U6566 ( .A(n1734), .B(n1733), .S(n2097), .Z(n1735) );
  MUX2_X1 U6567 ( .A(n1735), .B(n1732), .S(n2088), .Z(n1736) );
  MUX2_X1 U6568 ( .A(\mem[54][6] ), .B(\mem[55][6] ), .S(n2203), .Z(n1737) );
  MUX2_X1 U6569 ( .A(\mem[52][6] ), .B(\mem[53][6] ), .S(n2203), .Z(n1738) );
  MUX2_X1 U6570 ( .A(n1738), .B(n1737), .S(n2093), .Z(n1739) );
  MUX2_X1 U6571 ( .A(\mem[50][6] ), .B(\mem[51][6] ), .S(n2203), .Z(n1740) );
  MUX2_X1 U6572 ( .A(\mem[48][6] ), .B(\mem[49][6] ), .S(n2203), .Z(n1741) );
  MUX2_X1 U6573 ( .A(n1741), .B(n1740), .S(n2094), .Z(n1742) );
  MUX2_X1 U6574 ( .A(n1742), .B(n1739), .S(N20), .Z(n1743) );
  MUX2_X1 U6575 ( .A(n1743), .B(n1736), .S(n2066), .Z(n1744) );
  MUX2_X1 U6576 ( .A(\mem[46][6] ), .B(\mem[47][6] ), .S(n2203), .Z(n1745) );
  MUX2_X1 U6577 ( .A(\mem[44][6] ), .B(\mem[45][6] ), .S(n2203), .Z(n1746) );
  MUX2_X1 U6578 ( .A(n1746), .B(n1745), .S(n2092), .Z(n1747) );
  MUX2_X1 U6579 ( .A(\mem[42][6] ), .B(\mem[43][6] ), .S(n2203), .Z(n1748) );
  MUX2_X1 U6580 ( .A(\mem[40][6] ), .B(\mem[41][6] ), .S(n2203), .Z(n1749) );
  MUX2_X1 U6581 ( .A(n1749), .B(n1748), .S(n2096), .Z(n1750) );
  MUX2_X1 U6582 ( .A(n1750), .B(n1747), .S(N20), .Z(n1751) );
  MUX2_X1 U6583 ( .A(\mem[38][6] ), .B(\mem[39][6] ), .S(n2203), .Z(n1752) );
  MUX2_X1 U6584 ( .A(\mem[36][6] ), .B(\mem[37][6] ), .S(n2203), .Z(n1753) );
  MUX2_X1 U6585 ( .A(n1753), .B(n1752), .S(n2095), .Z(n1754) );
  MUX2_X1 U6586 ( .A(\mem[34][6] ), .B(\mem[35][6] ), .S(n2203), .Z(n1755) );
  MUX2_X1 U6587 ( .A(\mem[32][6] ), .B(\mem[33][6] ), .S(n2203), .Z(n1756) );
  MUX2_X1 U6588 ( .A(n1756), .B(n1755), .S(n2126), .Z(n1757) );
  MUX2_X1 U6589 ( .A(n1757), .B(n1754), .S(n2090), .Z(n1758) );
  MUX2_X1 U6590 ( .A(n1758), .B(n1751), .S(n2066), .Z(n1759) );
  MUX2_X1 U6591 ( .A(n1759), .B(n1744), .S(n2056), .Z(n1760) );
  MUX2_X1 U6592 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n2204), .Z(n1761) );
  MUX2_X1 U6593 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n2204), .Z(n1762) );
  MUX2_X1 U6594 ( .A(n1762), .B(n1761), .S(n2093), .Z(n1763) );
  MUX2_X1 U6595 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n2204), .Z(n1764) );
  MUX2_X1 U6596 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n2204), .Z(n1765) );
  MUX2_X1 U6597 ( .A(n1765), .B(n1764), .S(n2100), .Z(n1766) );
  MUX2_X1 U6598 ( .A(n1766), .B(n1763), .S(n2084), .Z(n1767) );
  MUX2_X1 U6599 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n2204), .Z(n1768) );
  MUX2_X1 U6600 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n2204), .Z(n1769) );
  MUX2_X1 U6601 ( .A(n1769), .B(n1768), .S(n2109), .Z(n1770) );
  MUX2_X1 U6602 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n2204), .Z(n1771) );
  MUX2_X1 U6603 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n2204), .Z(n1772) );
  MUX2_X1 U6604 ( .A(n1772), .B(n1771), .S(n2093), .Z(n1773) );
  MUX2_X1 U6605 ( .A(n1773), .B(n1770), .S(n2084), .Z(n1774) );
  MUX2_X1 U6606 ( .A(n1774), .B(n1767), .S(n2066), .Z(n1775) );
  MUX2_X1 U6607 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n2204), .Z(n1776) );
  MUX2_X1 U6608 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n2204), .Z(n1777) );
  MUX2_X1 U6609 ( .A(n1777), .B(n1776), .S(n2108), .Z(n1778) );
  MUX2_X1 U6610 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n2204), .Z(n1779) );
  MUX2_X1 U6611 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n2204), .Z(n1780) );
  MUX2_X1 U6612 ( .A(n1780), .B(n1779), .S(n2100), .Z(n1781) );
  MUX2_X1 U6613 ( .A(n1781), .B(n1778), .S(n2084), .Z(n1782) );
  MUX2_X1 U6614 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n1), .Z(n1783) );
  MUX2_X1 U6615 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n1), .Z(n1784) );
  MUX2_X1 U6616 ( .A(n1784), .B(n1783), .S(n2092), .Z(n1785) );
  MUX2_X1 U6617 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n1), .Z(n1786) );
  MUX2_X1 U6618 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n1), .Z(n1787) );
  MUX2_X1 U6619 ( .A(n1787), .B(n1786), .S(n2135), .Z(n1788) );
  MUX2_X1 U6620 ( .A(n1788), .B(n1785), .S(n2084), .Z(n1789) );
  MUX2_X1 U6621 ( .A(n1789), .B(n1782), .S(n2066), .Z(n1790) );
  MUX2_X1 U6622 ( .A(n1790), .B(n1775), .S(n2056), .Z(n1791) );
  MUX2_X1 U6623 ( .A(n1791), .B(n1760), .S(n2050), .Z(n1792) );
  MUX2_X1 U6624 ( .A(n1792), .B(n1729), .S(N24), .Z(n1793) );
  MUX2_X1 U6625 ( .A(\mem[254][7] ), .B(\mem[255][7] ), .S(n2189), .Z(n1794)
         );
  MUX2_X1 U6626 ( .A(\mem[252][7] ), .B(\mem[253][7] ), .S(n2205), .Z(n1795)
         );
  MUX2_X1 U6627 ( .A(n1795), .B(n1794), .S(n2107), .Z(n1796) );
  MUX2_X1 U6628 ( .A(\mem[250][7] ), .B(\mem[251][7] ), .S(n2205), .Z(n1797)
         );
  MUX2_X1 U6629 ( .A(\mem[248][7] ), .B(\mem[249][7] ), .S(n2205), .Z(n1798)
         );
  MUX2_X1 U6630 ( .A(n1798), .B(n1797), .S(n2111), .Z(n1799) );
  MUX2_X1 U6631 ( .A(n1799), .B(n1796), .S(n2084), .Z(n1800) );
  MUX2_X1 U6632 ( .A(\mem[246][7] ), .B(\mem[247][7] ), .S(n2205), .Z(n1801)
         );
  MUX2_X1 U6633 ( .A(\mem[244][7] ), .B(\mem[245][7] ), .S(n2205), .Z(n1802)
         );
  MUX2_X1 U6634 ( .A(n1802), .B(n1801), .S(n2109), .Z(n1803) );
  MUX2_X1 U6635 ( .A(\mem[242][7] ), .B(\mem[243][7] ), .S(n2205), .Z(n1804)
         );
  MUX2_X1 U6636 ( .A(\mem[240][7] ), .B(\mem[241][7] ), .S(n1), .Z(n1805) );
  MUX2_X1 U6637 ( .A(n1805), .B(n1804), .S(n2112), .Z(n1806) );
  MUX2_X1 U6638 ( .A(n1806), .B(n1803), .S(n2084), .Z(n1807) );
  MUX2_X1 U6639 ( .A(n1807), .B(n1800), .S(n2066), .Z(n1808) );
  MUX2_X1 U6640 ( .A(\mem[238][7] ), .B(\mem[239][7] ), .S(n2206), .Z(n1809)
         );
  MUX2_X1 U6641 ( .A(\mem[236][7] ), .B(\mem[237][7] ), .S(n2206), .Z(n1810)
         );
  MUX2_X1 U6642 ( .A(n1810), .B(n1809), .S(n2131), .Z(n1811) );
  MUX2_X1 U6643 ( .A(\mem[234][7] ), .B(\mem[235][7] ), .S(n2206), .Z(n1812)
         );
  MUX2_X1 U6644 ( .A(\mem[232][7] ), .B(\mem[233][7] ), .S(n2206), .Z(n1813)
         );
  MUX2_X1 U6645 ( .A(n1813), .B(n1812), .S(n2131), .Z(n1814) );
  MUX2_X1 U6646 ( .A(n1814), .B(n1811), .S(n2084), .Z(n1815) );
  MUX2_X1 U6647 ( .A(\mem[230][7] ), .B(\mem[231][7] ), .S(n2206), .Z(n1816)
         );
  MUX2_X1 U6648 ( .A(\mem[228][7] ), .B(\mem[229][7] ), .S(n2206), .Z(n1817)
         );
  MUX2_X1 U6649 ( .A(n1817), .B(n1816), .S(n2131), .Z(n1818) );
  MUX2_X1 U6650 ( .A(\mem[226][7] ), .B(\mem[227][7] ), .S(n2206), .Z(n1819)
         );
  MUX2_X1 U6651 ( .A(\mem[224][7] ), .B(\mem[225][7] ), .S(n2206), .Z(n1820)
         );
  MUX2_X1 U6652 ( .A(n1820), .B(n1819), .S(n2131), .Z(n1821) );
  MUX2_X1 U6653 ( .A(n1821), .B(n1818), .S(n2084), .Z(n1822) );
  MUX2_X1 U6654 ( .A(n1822), .B(n1815), .S(n2066), .Z(n1823) );
  MUX2_X1 U6655 ( .A(n1823), .B(n1808), .S(n2056), .Z(n1824) );
  MUX2_X1 U6656 ( .A(\mem[222][7] ), .B(\mem[223][7] ), .S(n2206), .Z(n1825)
         );
  MUX2_X1 U6657 ( .A(\mem[220][7] ), .B(\mem[221][7] ), .S(n2206), .Z(n1826)
         );
  MUX2_X1 U6658 ( .A(n1826), .B(n1825), .S(n2131), .Z(n1827) );
  MUX2_X1 U6659 ( .A(\mem[218][7] ), .B(\mem[219][7] ), .S(n2206), .Z(n1828)
         );
  MUX2_X1 U6660 ( .A(\mem[216][7] ), .B(\mem[217][7] ), .S(n2206), .Z(n1829)
         );
  MUX2_X1 U6661 ( .A(n1829), .B(n1828), .S(n2131), .Z(n1830) );
  MUX2_X1 U6662 ( .A(n1830), .B(n1827), .S(n2084), .Z(n1831) );
  MUX2_X1 U6663 ( .A(\mem[214][7] ), .B(\mem[215][7] ), .S(n2207), .Z(n1832)
         );
  MUX2_X1 U6664 ( .A(\mem[212][7] ), .B(\mem[213][7] ), .S(n2207), .Z(n1833)
         );
  MUX2_X1 U6665 ( .A(n1833), .B(n1832), .S(n2131), .Z(n1834) );
  MUX2_X1 U6666 ( .A(\mem[210][7] ), .B(\mem[211][7] ), .S(n2207), .Z(n1835)
         );
  MUX2_X1 U6667 ( .A(\mem[208][7] ), .B(\mem[209][7] ), .S(n2207), .Z(n1836)
         );
  MUX2_X1 U6668 ( .A(n1836), .B(n1835), .S(n2131), .Z(n1837) );
  MUX2_X1 U6669 ( .A(n1837), .B(n1834), .S(n2084), .Z(n1838) );
  MUX2_X1 U6670 ( .A(n1838), .B(n1831), .S(n2066), .Z(n1839) );
  MUX2_X1 U6671 ( .A(\mem[206][7] ), .B(\mem[207][7] ), .S(n2207), .Z(n1840)
         );
  MUX2_X1 U6672 ( .A(\mem[204][7] ), .B(\mem[205][7] ), .S(n2207), .Z(n1841)
         );
  MUX2_X1 U6673 ( .A(n1841), .B(n1840), .S(n2131), .Z(n1842) );
  MUX2_X1 U6674 ( .A(\mem[202][7] ), .B(\mem[203][7] ), .S(n2207), .Z(n1843)
         );
  MUX2_X1 U6675 ( .A(\mem[200][7] ), .B(\mem[201][7] ), .S(n2207), .Z(n1844)
         );
  MUX2_X1 U6676 ( .A(n1844), .B(n1843), .S(n2131), .Z(n1845) );
  MUX2_X1 U6677 ( .A(n1845), .B(n1842), .S(n2084), .Z(n1846) );
  MUX2_X1 U6678 ( .A(\mem[198][7] ), .B(\mem[199][7] ), .S(n2207), .Z(n1847)
         );
  MUX2_X1 U6679 ( .A(\mem[196][7] ), .B(\mem[197][7] ), .S(n2207), .Z(n1848)
         );
  MUX2_X1 U6680 ( .A(n1848), .B(n1847), .S(n2131), .Z(n1849) );
  MUX2_X1 U6681 ( .A(\mem[194][7] ), .B(\mem[195][7] ), .S(n2207), .Z(n1850)
         );
  MUX2_X1 U6682 ( .A(\mem[192][7] ), .B(\mem[193][7] ), .S(n2207), .Z(n1851)
         );
  MUX2_X1 U6683 ( .A(n1851), .B(n1850), .S(n2131), .Z(n1852) );
  MUX2_X1 U6684 ( .A(n1852), .B(n1849), .S(n2084), .Z(n1853) );
  MUX2_X1 U6685 ( .A(n1853), .B(n1846), .S(n2066), .Z(n1854) );
  MUX2_X1 U6686 ( .A(n1854), .B(n1839), .S(n2056), .Z(n1855) );
  MUX2_X1 U6687 ( .A(n1855), .B(n1824), .S(n2050), .Z(n1856) );
  MUX2_X1 U6688 ( .A(\mem[190][7] ), .B(\mem[191][7] ), .S(n2212), .Z(n1857)
         );
  MUX2_X1 U6689 ( .A(\mem[188][7] ), .B(\mem[189][7] ), .S(n2208), .Z(n1858)
         );
  MUX2_X1 U6690 ( .A(n1858), .B(n1857), .S(n2132), .Z(n1859) );
  MUX2_X1 U6691 ( .A(\mem[186][7] ), .B(\mem[187][7] ), .S(n2209), .Z(n1860)
         );
  MUX2_X1 U6692 ( .A(\mem[184][7] ), .B(\mem[185][7] ), .S(n2209), .Z(n1861)
         );
  MUX2_X1 U6693 ( .A(n1861), .B(n1860), .S(n2132), .Z(n1862) );
  MUX2_X1 U6694 ( .A(n1862), .B(n1859), .S(n2085), .Z(n1863) );
  MUX2_X1 U6695 ( .A(\mem[182][7] ), .B(\mem[183][7] ), .S(n2170), .Z(n1864)
         );
  MUX2_X1 U6696 ( .A(\mem[180][7] ), .B(\mem[181][7] ), .S(n2209), .Z(n1865)
         );
  MUX2_X1 U6697 ( .A(n1865), .B(n1864), .S(n2132), .Z(n1866) );
  MUX2_X1 U6698 ( .A(\mem[178][7] ), .B(\mem[179][7] ), .S(n2208), .Z(n1867)
         );
  MUX2_X1 U6699 ( .A(\mem[176][7] ), .B(\mem[177][7] ), .S(n2209), .Z(n1868)
         );
  MUX2_X1 U6700 ( .A(n1868), .B(n1867), .S(n2132), .Z(n1869) );
  MUX2_X1 U6701 ( .A(n1869), .B(n1866), .S(n2085), .Z(n1870) );
  MUX2_X1 U6702 ( .A(n1870), .B(n1863), .S(n2067), .Z(n1871) );
  MUX2_X1 U6703 ( .A(\mem[174][7] ), .B(\mem[175][7] ), .S(n2211), .Z(n1872)
         );
  MUX2_X1 U6704 ( .A(\mem[172][7] ), .B(\mem[173][7] ), .S(n2211), .Z(n1873)
         );
  MUX2_X1 U6705 ( .A(n1873), .B(n1872), .S(n2132), .Z(n1874) );
  MUX2_X1 U6706 ( .A(\mem[170][7] ), .B(\mem[171][7] ), .S(n2210), .Z(n1875)
         );
  MUX2_X1 U6707 ( .A(\mem[168][7] ), .B(\mem[169][7] ), .S(n2212), .Z(n1876)
         );
  MUX2_X1 U6708 ( .A(n1876), .B(n1875), .S(n2132), .Z(n1877) );
  MUX2_X1 U6709 ( .A(n1877), .B(n1874), .S(n2085), .Z(n1878) );
  MUX2_X1 U6710 ( .A(\mem[166][7] ), .B(\mem[167][7] ), .S(n2209), .Z(n1879)
         );
  MUX2_X1 U6711 ( .A(\mem[164][7] ), .B(\mem[165][7] ), .S(n2210), .Z(n1880)
         );
  MUX2_X1 U6712 ( .A(n1880), .B(n1879), .S(n2132), .Z(n1881) );
  MUX2_X1 U6713 ( .A(\mem[162][7] ), .B(\mem[163][7] ), .S(n2212), .Z(n1882)
         );
  MUX2_X1 U6714 ( .A(\mem[160][7] ), .B(\mem[161][7] ), .S(n2184), .Z(n1883)
         );
  MUX2_X1 U6715 ( .A(n1883), .B(n1882), .S(n2132), .Z(n1884) );
  MUX2_X1 U6716 ( .A(n1884), .B(n1881), .S(n2085), .Z(n1885) );
  MUX2_X1 U6717 ( .A(n1885), .B(n1878), .S(n2067), .Z(n1886) );
  MUX2_X1 U6718 ( .A(n1886), .B(n1871), .S(n2056), .Z(n1887) );
  MUX2_X1 U6719 ( .A(\mem[158][7] ), .B(\mem[159][7] ), .S(n2211), .Z(n1888)
         );
  MUX2_X1 U6720 ( .A(\mem[156][7] ), .B(\mem[157][7] ), .S(n2210), .Z(n1889)
         );
  MUX2_X1 U6721 ( .A(n1889), .B(n1888), .S(n2132), .Z(n1890) );
  MUX2_X1 U6722 ( .A(\mem[154][7] ), .B(\mem[155][7] ), .S(n2210), .Z(n1891)
         );
  MUX2_X1 U6723 ( .A(\mem[152][7] ), .B(\mem[153][7] ), .S(n2211), .Z(n1892)
         );
  MUX2_X1 U6724 ( .A(n1892), .B(n1891), .S(n2132), .Z(n1893) );
  MUX2_X1 U6725 ( .A(n1893), .B(n1890), .S(n2085), .Z(n1894) );
  MUX2_X1 U6726 ( .A(\mem[150][7] ), .B(\mem[151][7] ), .S(n2212), .Z(n1895)
         );
  MUX2_X1 U6727 ( .A(\mem[148][7] ), .B(\mem[149][7] ), .S(n2208), .Z(n1896)
         );
  MUX2_X1 U6728 ( .A(n1896), .B(n1895), .S(n2132), .Z(n1897) );
  MUX2_X1 U6729 ( .A(\mem[146][7] ), .B(\mem[147][7] ), .S(n2210), .Z(n1898)
         );
  MUX2_X1 U6730 ( .A(\mem[144][7] ), .B(\mem[145][7] ), .S(n2211), .Z(n1899)
         );
  MUX2_X1 U6731 ( .A(n1899), .B(n1898), .S(n2132), .Z(n1900) );
  MUX2_X1 U6732 ( .A(n1900), .B(n1897), .S(n2085), .Z(n1901) );
  MUX2_X1 U6733 ( .A(n1901), .B(n1894), .S(n2067), .Z(n1902) );
  MUX2_X1 U6734 ( .A(\mem[142][7] ), .B(\mem[143][7] ), .S(n2211), .Z(n1903)
         );
  MUX2_X1 U6735 ( .A(\mem[140][7] ), .B(\mem[141][7] ), .S(n2212), .Z(n1904)
         );
  MUX2_X1 U6736 ( .A(n1904), .B(n1903), .S(n2117), .Z(n1905) );
  MUX2_X1 U6737 ( .A(\mem[138][7] ), .B(\mem[139][7] ), .S(n2210), .Z(n1906)
         );
  MUX2_X1 U6738 ( .A(\mem[136][7] ), .B(\mem[137][7] ), .S(n2211), .Z(n1907)
         );
  MUX2_X1 U6739 ( .A(n1907), .B(n1906), .S(n2122), .Z(n1908) );
  MUX2_X1 U6740 ( .A(n1908), .B(n1905), .S(n2085), .Z(n1909) );
  MUX2_X1 U6741 ( .A(\mem[134][7] ), .B(\mem[135][7] ), .S(n2209), .Z(n1910)
         );
  MUX2_X1 U6742 ( .A(\mem[132][7] ), .B(\mem[133][7] ), .S(n2208), .Z(n1911)
         );
  MUX2_X1 U6743 ( .A(n1911), .B(n1910), .S(n2121), .Z(n1912) );
  MUX2_X1 U6744 ( .A(\mem[130][7] ), .B(\mem[131][7] ), .S(n2208), .Z(n1913)
         );
  MUX2_X1 U6745 ( .A(\mem[128][7] ), .B(\mem[129][7] ), .S(n2209), .Z(n1914)
         );
  MUX2_X1 U6746 ( .A(n1914), .B(n1913), .S(n2127), .Z(n1915) );
  MUX2_X1 U6747 ( .A(n1915), .B(n1912), .S(n2085), .Z(n1916) );
  MUX2_X1 U6748 ( .A(n1916), .B(n1909), .S(n2067), .Z(n1917) );
  MUX2_X1 U6749 ( .A(n1917), .B(n1902), .S(n2056), .Z(n1918) );
  MUX2_X1 U6750 ( .A(n1918), .B(n1887), .S(n2050), .Z(n1919) );
  MUX2_X1 U6751 ( .A(n1919), .B(n1856), .S(N24), .Z(n1920) );
  MUX2_X1 U6752 ( .A(\mem[126][7] ), .B(\mem[127][7] ), .S(n2212), .Z(n1921)
         );
  MUX2_X1 U6753 ( .A(\mem[124][7] ), .B(\mem[125][7] ), .S(n2210), .Z(n1922)
         );
  MUX2_X1 U6754 ( .A(n1922), .B(n1921), .S(n2119), .Z(n1923) );
  MUX2_X1 U6755 ( .A(\mem[122][7] ), .B(\mem[123][7] ), .S(n2208), .Z(n1924)
         );
  MUX2_X1 U6756 ( .A(\mem[120][7] ), .B(\mem[121][7] ), .S(n2184), .Z(n1925)
         );
  MUX2_X1 U6757 ( .A(n1925), .B(n1924), .S(n2128), .Z(n1926) );
  MUX2_X1 U6758 ( .A(n1926), .B(n1923), .S(n2085), .Z(n1927) );
  MUX2_X1 U6759 ( .A(\mem[118][7] ), .B(\mem[119][7] ), .S(n2210), .Z(n1928)
         );
  MUX2_X1 U6760 ( .A(\mem[116][7] ), .B(\mem[117][7] ), .S(n2208), .Z(n1929)
         );
  MUX2_X1 U6761 ( .A(n1929), .B(n1928), .S(n2124), .Z(n1930) );
  MUX2_X1 U6762 ( .A(\mem[114][7] ), .B(\mem[115][7] ), .S(n2209), .Z(n1931)
         );
  MUX2_X1 U6763 ( .A(\mem[112][7] ), .B(\mem[113][7] ), .S(n2200), .Z(n1932)
         );
  MUX2_X1 U6764 ( .A(n1932), .B(n1931), .S(n2114), .Z(n1933) );
  MUX2_X1 U6765 ( .A(n1933), .B(n1930), .S(n2085), .Z(n1934) );
  MUX2_X1 U6766 ( .A(n1934), .B(n1927), .S(n2067), .Z(n1935) );
  MUX2_X1 U6767 ( .A(\mem[110][7] ), .B(\mem[111][7] ), .S(n2208), .Z(n1936)
         );
  MUX2_X1 U6768 ( .A(\mem[108][7] ), .B(\mem[109][7] ), .S(n2200), .Z(n1937)
         );
  MUX2_X1 U6769 ( .A(n1937), .B(n1936), .S(n2123), .Z(n1938) );
  MUX2_X1 U6770 ( .A(\mem[106][7] ), .B(\mem[107][7] ), .S(n2212), .Z(n1939)
         );
  MUX2_X1 U6771 ( .A(\mem[104][7] ), .B(\mem[105][7] ), .S(n2211), .Z(n1940)
         );
  MUX2_X1 U6772 ( .A(n1940), .B(n1939), .S(n2110), .Z(n1941) );
  MUX2_X1 U6773 ( .A(n1941), .B(n1938), .S(n2085), .Z(n1942) );
  MUX2_X1 U6774 ( .A(\mem[102][7] ), .B(\mem[103][7] ), .S(n2208), .Z(n1943)
         );
  MUX2_X1 U6775 ( .A(\mem[100][7] ), .B(\mem[101][7] ), .S(n2210), .Z(n1944)
         );
  MUX2_X1 U6776 ( .A(n1944), .B(n1943), .S(n2118), .Z(n1945) );
  MUX2_X1 U6777 ( .A(\mem[98][7] ), .B(\mem[99][7] ), .S(n2211), .Z(n1946) );
  MUX2_X1 U6778 ( .A(\mem[96][7] ), .B(\mem[97][7] ), .S(n2210), .Z(n1947) );
  MUX2_X1 U6779 ( .A(n1947), .B(n1946), .S(n2113), .Z(n1948) );
  MUX2_X1 U6780 ( .A(n1948), .B(n1945), .S(n2085), .Z(n1949) );
  MUX2_X1 U6781 ( .A(n1949), .B(n1942), .S(n2067), .Z(n1950) );
  MUX2_X1 U6782 ( .A(n1950), .B(n1935), .S(n2056), .Z(n1951) );
  MUX2_X1 U6783 ( .A(\mem[94][7] ), .B(\mem[95][7] ), .S(n2212), .Z(n1952) );
  MUX2_X1 U6784 ( .A(\mem[92][7] ), .B(\mem[93][7] ), .S(n2210), .Z(n1953) );
  MUX2_X1 U6785 ( .A(n1953), .B(n1952), .S(n2133), .Z(n1954) );
  MUX2_X1 U6786 ( .A(\mem[90][7] ), .B(\mem[91][7] ), .S(n2211), .Z(n1955) );
  MUX2_X1 U6787 ( .A(\mem[88][7] ), .B(\mem[89][7] ), .S(n2208), .Z(n1956) );
  MUX2_X1 U6788 ( .A(n1956), .B(n1955), .S(n2133), .Z(n1957) );
  MUX2_X1 U6789 ( .A(n1957), .B(n1954), .S(n2086), .Z(n1958) );
  MUX2_X1 U6790 ( .A(\mem[86][7] ), .B(\mem[87][7] ), .S(n2210), .Z(n1959) );
  MUX2_X1 U6791 ( .A(\mem[84][7] ), .B(\mem[85][7] ), .S(n2210), .Z(n1960) );
  MUX2_X1 U6792 ( .A(n1960), .B(n1959), .S(n2133), .Z(n1961) );
  MUX2_X1 U6793 ( .A(\mem[82][7] ), .B(\mem[83][7] ), .S(n2209), .Z(n1962) );
  MUX2_X1 U6794 ( .A(\mem[80][7] ), .B(\mem[81][7] ), .S(n2210), .Z(n1963) );
  MUX2_X1 U6795 ( .A(n1963), .B(n1962), .S(n2133), .Z(n1964) );
  MUX2_X1 U6796 ( .A(n1964), .B(n1961), .S(n2086), .Z(n1965) );
  MUX2_X1 U6797 ( .A(n1965), .B(n1958), .S(n2067), .Z(n1966) );
  MUX2_X1 U6798 ( .A(\mem[78][7] ), .B(\mem[79][7] ), .S(n2210), .Z(n1967) );
  MUX2_X1 U6799 ( .A(\mem[76][7] ), .B(\mem[77][7] ), .S(n2210), .Z(n1968) );
  MUX2_X1 U6800 ( .A(n1968), .B(n1967), .S(n2133), .Z(n1969) );
  MUX2_X1 U6801 ( .A(\mem[74][7] ), .B(\mem[75][7] ), .S(n2212), .Z(n1970) );
  MUX2_X1 U6802 ( .A(\mem[72][7] ), .B(\mem[73][7] ), .S(n2212), .Z(n1971) );
  MUX2_X1 U6803 ( .A(n1971), .B(n1970), .S(n2133), .Z(n1972) );
  MUX2_X1 U6804 ( .A(n1972), .B(n1969), .S(n2086), .Z(n1973) );
  MUX2_X1 U6805 ( .A(\mem[70][7] ), .B(\mem[71][7] ), .S(n2208), .Z(n1974) );
  MUX2_X1 U6806 ( .A(\mem[68][7] ), .B(\mem[69][7] ), .S(n2209), .Z(n1975) );
  MUX2_X1 U6807 ( .A(n1975), .B(n1974), .S(n2133), .Z(n1976) );
  MUX2_X1 U6808 ( .A(\mem[66][7] ), .B(\mem[67][7] ), .S(n2211), .Z(n1977) );
  MUX2_X1 U6809 ( .A(\mem[64][7] ), .B(\mem[65][7] ), .S(n2209), .Z(n1978) );
  MUX2_X1 U6810 ( .A(n1978), .B(n1977), .S(n2133), .Z(n1979) );
  MUX2_X1 U6811 ( .A(n1979), .B(n1976), .S(n2086), .Z(n1980) );
  MUX2_X1 U6812 ( .A(n1980), .B(n1973), .S(n2067), .Z(n1981) );
  MUX2_X1 U6813 ( .A(n1981), .B(n1966), .S(n2056), .Z(n1982) );
  MUX2_X1 U6814 ( .A(n1982), .B(n1951), .S(n2050), .Z(n1983) );
  MUX2_X1 U6815 ( .A(\mem[62][7] ), .B(\mem[63][7] ), .S(n2200), .Z(n1984) );
  MUX2_X1 U6816 ( .A(\mem[60][7] ), .B(\mem[61][7] ), .S(n2211), .Z(n1985) );
  MUX2_X1 U6817 ( .A(n1985), .B(n1984), .S(n2133), .Z(n1986) );
  MUX2_X1 U6818 ( .A(\mem[58][7] ), .B(\mem[59][7] ), .S(n2210), .Z(n1987) );
  MUX2_X1 U6819 ( .A(\mem[56][7] ), .B(\mem[57][7] ), .S(n2209), .Z(n1988) );
  MUX2_X1 U6820 ( .A(n1988), .B(n1987), .S(n2133), .Z(n1989) );
  MUX2_X1 U6821 ( .A(n1989), .B(n1986), .S(n2086), .Z(n1990) );
  MUX2_X1 U6822 ( .A(\mem[54][7] ), .B(\mem[55][7] ), .S(n2184), .Z(n1991) );
  MUX2_X1 U6823 ( .A(\mem[52][7] ), .B(\mem[53][7] ), .S(n2210), .Z(n1992) );
  MUX2_X1 U6824 ( .A(n1992), .B(n1991), .S(n2133), .Z(n1993) );
  MUX2_X1 U6825 ( .A(\mem[50][7] ), .B(\mem[51][7] ), .S(n2212), .Z(n1994) );
  MUX2_X1 U6826 ( .A(\mem[48][7] ), .B(\mem[49][7] ), .S(n2208), .Z(n1995) );
  MUX2_X1 U6827 ( .A(n1995), .B(n1994), .S(n2133), .Z(n1996) );
  MUX2_X1 U6828 ( .A(n1996), .B(n1993), .S(n2086), .Z(n1997) );
  MUX2_X1 U6829 ( .A(n1997), .B(n1990), .S(n2067), .Z(n1998) );
  MUX2_X1 U6830 ( .A(\mem[46][7] ), .B(\mem[47][7] ), .S(n2213), .Z(n1999) );
  MUX2_X1 U6831 ( .A(\mem[44][7] ), .B(\mem[45][7] ), .S(n2213), .Z(n2000) );
  MUX2_X1 U6832 ( .A(n2000), .B(n1999), .S(n2134), .Z(n2001) );
  MUX2_X1 U6833 ( .A(\mem[42][7] ), .B(\mem[43][7] ), .S(n2213), .Z(n2002) );
  MUX2_X1 U6834 ( .A(\mem[40][7] ), .B(\mem[41][7] ), .S(n2213), .Z(n2003) );
  MUX2_X1 U6835 ( .A(n2003), .B(n2002), .S(n2134), .Z(n2004) );
  MUX2_X1 U6836 ( .A(n2004), .B(n2001), .S(n2086), .Z(n2005) );
  MUX2_X1 U6837 ( .A(\mem[38][7] ), .B(\mem[39][7] ), .S(n2213), .Z(n2006) );
  MUX2_X1 U6838 ( .A(\mem[36][7] ), .B(\mem[37][7] ), .S(n2213), .Z(n2007) );
  MUX2_X1 U6839 ( .A(n2007), .B(n2006), .S(n2134), .Z(n2008) );
  MUX2_X1 U6840 ( .A(\mem[34][7] ), .B(\mem[35][7] ), .S(n2213), .Z(n2009) );
  MUX2_X1 U6841 ( .A(\mem[32][7] ), .B(\mem[33][7] ), .S(n2213), .Z(n2010) );
  MUX2_X1 U6842 ( .A(n2010), .B(n2009), .S(n2134), .Z(n2011) );
  MUX2_X1 U6843 ( .A(n2011), .B(n2008), .S(n2086), .Z(n2012) );
  MUX2_X1 U6844 ( .A(n2012), .B(n2005), .S(n2067), .Z(n2013) );
  MUX2_X1 U6845 ( .A(n2013), .B(n1998), .S(n2056), .Z(n2014) );
  MUX2_X1 U6846 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n2213), .Z(n2015) );
  MUX2_X1 U6847 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n2213), .Z(n2016) );
  MUX2_X1 U6848 ( .A(n2016), .B(n2015), .S(n2134), .Z(n2017) );
  MUX2_X1 U6849 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n2213), .Z(n2018) );
  MUX2_X1 U6850 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n2213), .Z(n2019) );
  MUX2_X1 U6851 ( .A(n2019), .B(n2018), .S(n2134), .Z(n2020) );
  MUX2_X1 U6852 ( .A(n2020), .B(n2017), .S(n2086), .Z(n2021) );
  MUX2_X1 U6853 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n2214), .Z(n2022) );
  MUX2_X1 U6854 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n2214), .Z(n2023) );
  MUX2_X1 U6855 ( .A(n2023), .B(n2022), .S(n2134), .Z(n2024) );
  MUX2_X1 U6856 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n2214), .Z(n2025) );
  MUX2_X1 U6857 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n2214), .Z(n2026) );
  MUX2_X1 U6858 ( .A(n2026), .B(n2025), .S(n2134), .Z(n2027) );
  MUX2_X1 U6859 ( .A(n2027), .B(n2024), .S(n2086), .Z(n2028) );
  MUX2_X1 U6860 ( .A(n2028), .B(n2021), .S(n2067), .Z(n2029) );
  MUX2_X1 U6861 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n2214), .Z(n2030) );
  MUX2_X1 U6862 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n2214), .Z(n2031) );
  MUX2_X1 U6863 ( .A(n2031), .B(n2030), .S(n2134), .Z(n2032) );
  MUX2_X1 U6864 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n2214), .Z(n2033) );
  MUX2_X1 U6865 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n2214), .Z(n2034) );
  MUX2_X1 U6866 ( .A(n2034), .B(n2033), .S(n2134), .Z(n2035) );
  MUX2_X1 U6867 ( .A(n2035), .B(n2032), .S(n2086), .Z(n2036) );
  MUX2_X1 U6868 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n2214), .Z(n2037) );
  MUX2_X1 U6869 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n2214), .Z(n2038) );
  MUX2_X1 U6870 ( .A(n2038), .B(n2037), .S(n2134), .Z(n2039) );
  MUX2_X1 U6871 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n2214), .Z(n2040) );
  MUX2_X1 U6872 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n2214), .Z(n2041) );
  MUX2_X1 U6873 ( .A(n2041), .B(n2040), .S(n2134), .Z(n2042) );
  MUX2_X1 U6874 ( .A(n2042), .B(n2039), .S(n2086), .Z(n2043) );
  MUX2_X1 U6875 ( .A(n2043), .B(n2036), .S(n2067), .Z(n2044) );
  MUX2_X1 U6876 ( .A(n2044), .B(n2029), .S(n2056), .Z(n2045) );
  MUX2_X1 U6877 ( .A(n2045), .B(n2014), .S(n2050), .Z(n2046) );
  MUX2_X1 U6878 ( .A(n2046), .B(n1983), .S(N24), .Z(n2047) );
  CLKBUF_X1 U6879 ( .A(N22), .Z(n2051) );
  CLKBUF_X1 U6880 ( .A(n2068), .Z(n2057) );
  NOR2_X1 U6881 ( .A1(n13), .A2(N19), .ZN(n4549) );
  NOR2_X1 U6882 ( .A1(n2224), .A2(n2222), .ZN(n4527) );
  INV_X1 U6883 ( .A(N18), .ZN(n2223) );
  AND2_X4 U6884 ( .A1(n4549), .A2(n4528), .ZN(n2469) );
  AND2_X4 U6885 ( .A1(n4527), .A2(n4528), .ZN(n2327) );
endmodule


module memory_WIDTH16_SIZE16_LOGSIZE4 ( clk, data_in, data_out, addr, wr_en );
  input [15:0] data_in;
  output [15:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][15] , \mem[15][14] , \mem[15][13] ,
         \mem[15][12] , \mem[15][11] , \mem[15][10] , \mem[15][9] ,
         \mem[15][8] , \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] ,
         \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][15] ,
         \mem[14][14] , \mem[14][13] , \mem[14][12] , \mem[14][11] ,
         \mem[14][10] , \mem[14][9] , \mem[14][8] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][15] , \mem[13][14] , \mem[13][13] ,
         \mem[13][12] , \mem[13][11] , \mem[13][10] , \mem[13][9] ,
         \mem[13][8] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][15] ,
         \mem[12][14] , \mem[12][13] , \mem[12][12] , \mem[12][11] ,
         \mem[12][10] , \mem[12][9] , \mem[12][8] , \mem[12][7] , \mem[12][6] ,
         \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] , \mem[12][1] ,
         \mem[12][0] , \mem[11][15] , \mem[11][14] , \mem[11][13] ,
         \mem[11][12] , \mem[11][11] , \mem[11][10] , \mem[11][9] ,
         \mem[11][8] , \mem[11][7] , \mem[11][6] , \mem[11][5] , \mem[11][4] ,
         \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] , \mem[10][15] ,
         \mem[10][14] , \mem[10][13] , \mem[10][12] , \mem[10][11] ,
         \mem[10][10] , \mem[10][9] , \mem[10][8] , \mem[10][7] , \mem[10][6] ,
         \mem[10][5] , \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] ,
         \mem[10][0] , \mem[9][15] , \mem[9][14] , \mem[9][13] , \mem[9][12] ,
         \mem[9][11] , \mem[9][10] , \mem[9][9] , \mem[9][8] , \mem[9][7] ,
         \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] ,
         \mem[9][1] , \mem[9][0] , \mem[8][15] , \mem[8][14] , \mem[8][13] ,
         \mem[8][12] , \mem[8][11] , \mem[8][10] , \mem[8][9] , \mem[8][8] ,
         \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] , \mem[8][3] ,
         \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][15] , \mem[7][14] ,
         \mem[7][13] , \mem[7][12] , \mem[7][11] , \mem[7][10] , \mem[7][9] ,
         \mem[7][8] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][15] ,
         \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] ,
         \mem[4][11] , \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] ,
         \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] ,
         \mem[4][1] , \mem[4][0] , \mem[3][15] , \mem[3][14] , \mem[3][13] ,
         \mem[3][12] , \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] ,
         \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] ,
         \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][15] , \mem[2][14] ,
         \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] ,
         \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][15] ,
         \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[15]  ( .D(N14), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N15), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(N16), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(N17), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(N18), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N19), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N20), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N21), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N22), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N23), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N24), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N25), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N26), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N27), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N28), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N29), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][15]  ( .D(n557), .CK(clk), .Q(\mem[15][15] ) );
  DFF_X1 \mem_reg[15][14]  ( .D(n556), .CK(clk), .Q(\mem[15][14] ) );
  DFF_X1 \mem_reg[15][13]  ( .D(n555), .CK(clk), .Q(\mem[15][13] ) );
  DFF_X1 \mem_reg[15][12]  ( .D(n554), .CK(clk), .Q(\mem[15][12] ) );
  DFF_X1 \mem_reg[15][11]  ( .D(n553), .CK(clk), .Q(\mem[15][11] ) );
  DFF_X1 \mem_reg[15][10]  ( .D(n552), .CK(clk), .Q(\mem[15][10] ) );
  DFF_X1 \mem_reg[15][9]  ( .D(n551), .CK(clk), .Q(\mem[15][9] ) );
  DFF_X1 \mem_reg[15][8]  ( .D(n550), .CK(clk), .Q(\mem[15][8] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n549), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n548), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n547), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n546), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n545), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n544), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n543), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n542), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][15]  ( .D(n541), .CK(clk), .Q(\mem[14][15] ) );
  DFF_X1 \mem_reg[14][14]  ( .D(n540), .CK(clk), .Q(\mem[14][14] ) );
  DFF_X1 \mem_reg[14][13]  ( .D(n539), .CK(clk), .Q(\mem[14][13] ) );
  DFF_X1 \mem_reg[14][12]  ( .D(n538), .CK(clk), .Q(\mem[14][12] ) );
  DFF_X1 \mem_reg[14][11]  ( .D(n537), .CK(clk), .Q(\mem[14][11] ) );
  DFF_X1 \mem_reg[14][10]  ( .D(n536), .CK(clk), .Q(\mem[14][10] ) );
  DFF_X1 \mem_reg[14][9]  ( .D(n535), .CK(clk), .Q(\mem[14][9] ) );
  DFF_X1 \mem_reg[14][8]  ( .D(n534), .CK(clk), .Q(\mem[14][8] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n533), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n532), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n531), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n530), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n529), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n528), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n527), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n526), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][15]  ( .D(n525), .CK(clk), .Q(\mem[13][15] ) );
  DFF_X1 \mem_reg[13][14]  ( .D(n524), .CK(clk), .Q(\mem[13][14] ) );
  DFF_X1 \mem_reg[13][13]  ( .D(n523), .CK(clk), .Q(\mem[13][13] ) );
  DFF_X1 \mem_reg[13][12]  ( .D(n522), .CK(clk), .Q(\mem[13][12] ) );
  DFF_X1 \mem_reg[13][11]  ( .D(n521), .CK(clk), .Q(\mem[13][11] ) );
  DFF_X1 \mem_reg[13][10]  ( .D(n520), .CK(clk), .Q(\mem[13][10] ) );
  DFF_X1 \mem_reg[13][9]  ( .D(n519), .CK(clk), .Q(\mem[13][9] ) );
  DFF_X1 \mem_reg[13][8]  ( .D(n518), .CK(clk), .Q(\mem[13][8] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n517), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n516), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n515), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n514), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n513), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n512), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n511), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n510), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][15]  ( .D(n509), .CK(clk), .Q(\mem[12][15] ) );
  DFF_X1 \mem_reg[12][14]  ( .D(n508), .CK(clk), .Q(\mem[12][14] ) );
  DFF_X1 \mem_reg[12][13]  ( .D(n507), .CK(clk), .Q(\mem[12][13] ) );
  DFF_X1 \mem_reg[12][12]  ( .D(n506), .CK(clk), .Q(\mem[12][12] ) );
  DFF_X1 \mem_reg[12][11]  ( .D(n505), .CK(clk), .Q(\mem[12][11] ) );
  DFF_X1 \mem_reg[12][10]  ( .D(n504), .CK(clk), .Q(\mem[12][10] ) );
  DFF_X1 \mem_reg[12][9]  ( .D(n503), .CK(clk), .Q(\mem[12][9] ) );
  DFF_X1 \mem_reg[12][8]  ( .D(n502), .CK(clk), .Q(\mem[12][8] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n501), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n500), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n499), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n498), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n497), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n496), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n495), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n494), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][15]  ( .D(n493), .CK(clk), .Q(\mem[11][15] ) );
  DFF_X1 \mem_reg[11][14]  ( .D(n492), .CK(clk), .Q(\mem[11][14] ) );
  DFF_X1 \mem_reg[11][13]  ( .D(n491), .CK(clk), .Q(\mem[11][13] ) );
  DFF_X1 \mem_reg[11][12]  ( .D(n490), .CK(clk), .Q(\mem[11][12] ) );
  DFF_X1 \mem_reg[11][11]  ( .D(n489), .CK(clk), .Q(\mem[11][11] ) );
  DFF_X1 \mem_reg[11][10]  ( .D(n488), .CK(clk), .Q(\mem[11][10] ) );
  DFF_X1 \mem_reg[11][9]  ( .D(n487), .CK(clk), .Q(\mem[11][9] ) );
  DFF_X1 \mem_reg[11][8]  ( .D(n486), .CK(clk), .Q(\mem[11][8] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n485), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n484), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n483), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n482), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n481), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n480), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n479), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n478), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][15]  ( .D(n477), .CK(clk), .Q(\mem[10][15] ) );
  DFF_X1 \mem_reg[10][14]  ( .D(n476), .CK(clk), .Q(\mem[10][14] ) );
  DFF_X1 \mem_reg[10][13]  ( .D(n475), .CK(clk), .Q(\mem[10][13] ) );
  DFF_X1 \mem_reg[10][12]  ( .D(n474), .CK(clk), .Q(\mem[10][12] ) );
  DFF_X1 \mem_reg[10][11]  ( .D(n473), .CK(clk), .Q(\mem[10][11] ) );
  DFF_X1 \mem_reg[10][10]  ( .D(n472), .CK(clk), .Q(\mem[10][10] ) );
  DFF_X1 \mem_reg[10][9]  ( .D(n471), .CK(clk), .Q(\mem[10][9] ) );
  DFF_X1 \mem_reg[10][8]  ( .D(n470), .CK(clk), .Q(\mem[10][8] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n469), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n468), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n467), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n466), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n465), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n464), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n463), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n462), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][15]  ( .D(n461), .CK(clk), .Q(\mem[9][15] ) );
  DFF_X1 \mem_reg[9][14]  ( .D(n460), .CK(clk), .Q(\mem[9][14] ) );
  DFF_X1 \mem_reg[9][13]  ( .D(n459), .CK(clk), .Q(\mem[9][13] ) );
  DFF_X1 \mem_reg[9][12]  ( .D(n458), .CK(clk), .Q(\mem[9][12] ) );
  DFF_X1 \mem_reg[9][11]  ( .D(n457), .CK(clk), .Q(\mem[9][11] ) );
  DFF_X1 \mem_reg[9][10]  ( .D(n456), .CK(clk), .Q(\mem[9][10] ) );
  DFF_X1 \mem_reg[9][9]  ( .D(n455), .CK(clk), .Q(\mem[9][9] ) );
  DFF_X1 \mem_reg[9][8]  ( .D(n454), .CK(clk), .Q(\mem[9][8] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n453), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n452), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n451), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n450), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n449), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n448), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n447), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n446), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][15]  ( .D(n445), .CK(clk), .Q(\mem[8][15] ) );
  DFF_X1 \mem_reg[8][14]  ( .D(n444), .CK(clk), .Q(\mem[8][14] ) );
  DFF_X1 \mem_reg[8][13]  ( .D(n443), .CK(clk), .Q(\mem[8][13] ) );
  DFF_X1 \mem_reg[8][12]  ( .D(n442), .CK(clk), .Q(\mem[8][12] ) );
  DFF_X1 \mem_reg[8][11]  ( .D(n441), .CK(clk), .Q(\mem[8][11] ) );
  DFF_X1 \mem_reg[8][10]  ( .D(n440), .CK(clk), .Q(\mem[8][10] ) );
  DFF_X1 \mem_reg[8][9]  ( .D(n439), .CK(clk), .Q(\mem[8][9] ) );
  DFF_X1 \mem_reg[8][8]  ( .D(n438), .CK(clk), .Q(\mem[8][8] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n437), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n436), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n435), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n434), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n433), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n432), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n431), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n430), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n429), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n428), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n427), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n426), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n425), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n424), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n423), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n422), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n421), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n420), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n419), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n418), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n417), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n416), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n415), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n414), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n413), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n412), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n411), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n410), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n409), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n408), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n407), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n406), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n405), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n404), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n403), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n402), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n401), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n400), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n399), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n398), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n397), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n396), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n395), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n394), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n393), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n392), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n391), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n390), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n389), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n388), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n387), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n386), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n385), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n384), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n383), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n382), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n381), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n380), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n379), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n378), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n377), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n376), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n375), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n374), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n373), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n372), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n371), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n370), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n369), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n368), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n367), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n366), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n365), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n364), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n363), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n362), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n361), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n360), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n359), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n358), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n357), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n356), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n355), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n354), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n353), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n352), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n351), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n350), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n349), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n348), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n347), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n346), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n345), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n344), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n343), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n342), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n341), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n340), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n339), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n338), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n337), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n336), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n335), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n334), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n333), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n332), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n331), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n330), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n329), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n328), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n327), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n326), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n325), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n324), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n323), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n322), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n321), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n320), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n319), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n318), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n317), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n316), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n315), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n314), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n313), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n312), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n311), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n310), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n309), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n308), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n307), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n306), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n305), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n304), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n303), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n302), .CK(clk), .Q(\mem[0][0] ) );
  BUF_X1 U3 ( .A(N10), .Z(n770) );
  BUF_X1 U4 ( .A(n777), .Z(n774) );
  BUF_X1 U5 ( .A(n777), .Z(n775) );
  BUF_X1 U6 ( .A(n777), .Z(n776) );
  BUF_X1 U7 ( .A(n777), .Z(n773) );
  BUF_X1 U8 ( .A(n777), .Z(n771) );
  BUF_X1 U9 ( .A(n777), .Z(n772) );
  BUF_X1 U10 ( .A(n20), .Z(n793) );
  BUF_X1 U11 ( .A(n39), .Z(n792) );
  BUF_X1 U12 ( .A(n57), .Z(n791) );
  BUF_X1 U13 ( .A(n75), .Z(n790) );
  BUF_X1 U14 ( .A(n92), .Z(n789) );
  BUF_X1 U15 ( .A(n127), .Z(n787) );
  BUF_X1 U16 ( .A(n146), .Z(n786) );
  BUF_X1 U17 ( .A(n163), .Z(n785) );
  BUF_X1 U18 ( .A(n181), .Z(n784) );
  BUF_X1 U19 ( .A(n199), .Z(n783) );
  BUF_X1 U20 ( .A(n216), .Z(n782) );
  BUF_X1 U21 ( .A(n233), .Z(n781) );
  BUF_X1 U22 ( .A(n250), .Z(n780) );
  BUF_X1 U23 ( .A(n267), .Z(n779) );
  BUF_X1 U24 ( .A(n285), .Z(n778) );
  BUF_X1 U25 ( .A(n110), .Z(n788) );
  BUF_X1 U26 ( .A(N11), .Z(n765) );
  BUF_X1 U27 ( .A(N11), .Z(n766) );
  BUF_X1 U28 ( .A(N11), .Z(n767) );
  BUF_X1 U29 ( .A(N11), .Z(n768) );
  BUF_X1 U30 ( .A(N11), .Z(n769) );
  BUF_X1 U31 ( .A(N10), .Z(n777) );
  AND2_X1 U32 ( .A1(n145), .A2(n794), .ZN(n38) );
  AND2_X1 U33 ( .A1(N10), .A2(n145), .ZN(n56) );
  AND2_X1 U34 ( .A1(n284), .A2(N10), .ZN(n198) );
  AND2_X1 U35 ( .A1(n284), .A2(n794), .ZN(n180) );
  NAND2_X1 U36 ( .A1(n37), .A2(n38), .ZN(n20) );
  NAND2_X1 U37 ( .A1(n74), .A2(n38), .ZN(n57) );
  NAND2_X1 U38 ( .A1(n74), .A2(n56), .ZN(n75) );
  NAND2_X1 U39 ( .A1(n56), .A2(n37), .ZN(n39) );
  NAND2_X1 U40 ( .A1(n180), .A2(n37), .ZN(n163) );
  NAND2_X1 U41 ( .A1(n198), .A2(n37), .ZN(n181) );
  NAND2_X1 U42 ( .A1(n180), .A2(n74), .ZN(n199) );
  NAND2_X1 U43 ( .A1(n198), .A2(n74), .ZN(n216) );
  NAND2_X1 U44 ( .A1(n109), .A2(n38), .ZN(n92) );
  NAND2_X1 U45 ( .A1(n109), .A2(n56), .ZN(n110) );
  NAND2_X1 U46 ( .A1(n144), .A2(n38), .ZN(n127) );
  NAND2_X1 U47 ( .A1(n144), .A2(n56), .ZN(n146) );
  NAND2_X1 U48 ( .A1(n180), .A2(n144), .ZN(n267) );
  NAND2_X1 U49 ( .A1(n198), .A2(n144), .ZN(n285) );
  NAND2_X1 U50 ( .A1(n180), .A2(n109), .ZN(n233) );
  NAND2_X1 U51 ( .A1(n198), .A2(n109), .ZN(n250) );
  INV_X1 U52 ( .A(data_in[4]), .ZN(n801) );
  INV_X1 U53 ( .A(data_in[5]), .ZN(n802) );
  INV_X1 U54 ( .A(data_in[6]), .ZN(n803) );
  INV_X1 U55 ( .A(data_in[7]), .ZN(n804) );
  INV_X1 U56 ( .A(data_in[8]), .ZN(n805) );
  INV_X1 U57 ( .A(data_in[9]), .ZN(n806) );
  INV_X1 U58 ( .A(data_in[10]), .ZN(n807) );
  INV_X1 U59 ( .A(data_in[11]), .ZN(n808) );
  INV_X1 U60 ( .A(data_in[12]), .ZN(n809) );
  INV_X1 U61 ( .A(data_in[13]), .ZN(n810) );
  INV_X1 U62 ( .A(data_in[15]), .ZN(n812) );
  INV_X1 U63 ( .A(data_in[3]), .ZN(n800) );
  NOR2_X1 U64 ( .A1(N11), .A2(N12), .ZN(n37) );
  NOR2_X1 U65 ( .A1(n795), .A2(N12), .ZN(n74) );
  INV_X1 U66 ( .A(data_in[14]), .ZN(n811) );
  OAI21_X1 U67 ( .B1(n793), .B2(n797), .A(n21), .ZN(n302) );
  NAND2_X1 U68 ( .A1(\mem[0][0] ), .A2(n20), .ZN(n21) );
  OAI21_X1 U69 ( .B1(n793), .B2(n798), .A(n22), .ZN(n303) );
  NAND2_X1 U70 ( .A1(\mem[0][1] ), .A2(n20), .ZN(n22) );
  OAI21_X1 U71 ( .B1(n793), .B2(n799), .A(n23), .ZN(n304) );
  NAND2_X1 U72 ( .A1(\mem[0][2] ), .A2(n20), .ZN(n23) );
  OAI21_X1 U73 ( .B1(n797), .B2(n39), .A(n40), .ZN(n318) );
  NAND2_X1 U74 ( .A1(\mem[1][0] ), .A2(n792), .ZN(n40) );
  OAI21_X1 U75 ( .B1(n798), .B2(n39), .A(n41), .ZN(n319) );
  NAND2_X1 U76 ( .A1(\mem[1][1] ), .A2(n792), .ZN(n41) );
  OAI21_X1 U77 ( .B1(n799), .B2(n39), .A(n42), .ZN(n320) );
  NAND2_X1 U78 ( .A1(\mem[1][2] ), .A2(n792), .ZN(n42) );
  OAI21_X1 U79 ( .B1(n797), .B2(n57), .A(n58), .ZN(n334) );
  NAND2_X1 U80 ( .A1(\mem[2][0] ), .A2(n791), .ZN(n58) );
  OAI21_X1 U81 ( .B1(n798), .B2(n57), .A(n59), .ZN(n335) );
  NAND2_X1 U82 ( .A1(\mem[2][1] ), .A2(n791), .ZN(n59) );
  OAI21_X1 U83 ( .B1(n799), .B2(n57), .A(n60), .ZN(n336) );
  NAND2_X1 U84 ( .A1(\mem[2][2] ), .A2(n791), .ZN(n60) );
  OAI21_X1 U85 ( .B1(n797), .B2(n75), .A(n76), .ZN(n350) );
  NAND2_X1 U86 ( .A1(\mem[3][0] ), .A2(n790), .ZN(n76) );
  OAI21_X1 U87 ( .B1(n798), .B2(n75), .A(n77), .ZN(n351) );
  NAND2_X1 U88 ( .A1(\mem[3][1] ), .A2(n790), .ZN(n77) );
  OAI21_X1 U89 ( .B1(n799), .B2(n75), .A(n78), .ZN(n352) );
  NAND2_X1 U90 ( .A1(\mem[3][2] ), .A2(n790), .ZN(n78) );
  OAI21_X1 U91 ( .B1(n797), .B2(n92), .A(n93), .ZN(n366) );
  NAND2_X1 U92 ( .A1(\mem[4][0] ), .A2(n789), .ZN(n93) );
  OAI21_X1 U93 ( .B1(n798), .B2(n92), .A(n94), .ZN(n367) );
  NAND2_X1 U94 ( .A1(\mem[4][1] ), .A2(n789), .ZN(n94) );
  OAI21_X1 U95 ( .B1(n799), .B2(n92), .A(n95), .ZN(n368) );
  NAND2_X1 U96 ( .A1(\mem[4][2] ), .A2(n789), .ZN(n95) );
  OAI21_X1 U97 ( .B1(n797), .B2(n110), .A(n111), .ZN(n382) );
  NAND2_X1 U98 ( .A1(\mem[5][0] ), .A2(n110), .ZN(n111) );
  OAI21_X1 U99 ( .B1(n798), .B2(n110), .A(n112), .ZN(n383) );
  NAND2_X1 U100 ( .A1(\mem[5][1] ), .A2(n110), .ZN(n112) );
  OAI21_X1 U101 ( .B1(n799), .B2(n110), .A(n113), .ZN(n384) );
  NAND2_X1 U102 ( .A1(\mem[5][2] ), .A2(n110), .ZN(n113) );
  OAI21_X1 U103 ( .B1(n797), .B2(n127), .A(n128), .ZN(n398) );
  NAND2_X1 U104 ( .A1(\mem[6][0] ), .A2(n787), .ZN(n128) );
  OAI21_X1 U105 ( .B1(n798), .B2(n127), .A(n129), .ZN(n399) );
  NAND2_X1 U106 ( .A1(\mem[6][1] ), .A2(n787), .ZN(n129) );
  OAI21_X1 U107 ( .B1(n799), .B2(n127), .A(n130), .ZN(n400) );
  NAND2_X1 U108 ( .A1(\mem[6][2] ), .A2(n787), .ZN(n130) );
  OAI21_X1 U109 ( .B1(n797), .B2(n146), .A(n147), .ZN(n414) );
  NAND2_X1 U110 ( .A1(\mem[7][0] ), .A2(n786), .ZN(n147) );
  OAI21_X1 U111 ( .B1(n798), .B2(n146), .A(n148), .ZN(n415) );
  NAND2_X1 U112 ( .A1(\mem[7][1] ), .A2(n786), .ZN(n148) );
  OAI21_X1 U113 ( .B1(n799), .B2(n146), .A(n149), .ZN(n416) );
  NAND2_X1 U114 ( .A1(\mem[7][2] ), .A2(n786), .ZN(n149) );
  OAI21_X1 U115 ( .B1(n797), .B2(n163), .A(n164), .ZN(n430) );
  NAND2_X1 U116 ( .A1(\mem[8][0] ), .A2(n785), .ZN(n164) );
  OAI21_X1 U117 ( .B1(n798), .B2(n163), .A(n165), .ZN(n431) );
  NAND2_X1 U118 ( .A1(\mem[8][1] ), .A2(n785), .ZN(n165) );
  OAI21_X1 U119 ( .B1(n799), .B2(n163), .A(n166), .ZN(n432) );
  NAND2_X1 U120 ( .A1(\mem[8][2] ), .A2(n785), .ZN(n166) );
  OAI21_X1 U121 ( .B1(n797), .B2(n181), .A(n182), .ZN(n446) );
  NAND2_X1 U122 ( .A1(\mem[9][0] ), .A2(n784), .ZN(n182) );
  OAI21_X1 U123 ( .B1(n798), .B2(n181), .A(n183), .ZN(n447) );
  NAND2_X1 U124 ( .A1(\mem[9][1] ), .A2(n784), .ZN(n183) );
  OAI21_X1 U125 ( .B1(n799), .B2(n181), .A(n184), .ZN(n448) );
  NAND2_X1 U126 ( .A1(\mem[9][2] ), .A2(n784), .ZN(n184) );
  OAI21_X1 U127 ( .B1(n797), .B2(n199), .A(n200), .ZN(n462) );
  NAND2_X1 U128 ( .A1(\mem[10][0] ), .A2(n783), .ZN(n200) );
  OAI21_X1 U129 ( .B1(n798), .B2(n199), .A(n201), .ZN(n463) );
  NAND2_X1 U130 ( .A1(\mem[10][1] ), .A2(n783), .ZN(n201) );
  OAI21_X1 U131 ( .B1(n799), .B2(n199), .A(n202), .ZN(n464) );
  NAND2_X1 U132 ( .A1(\mem[10][2] ), .A2(n783), .ZN(n202) );
  OAI21_X1 U133 ( .B1(n797), .B2(n216), .A(n217), .ZN(n478) );
  NAND2_X1 U134 ( .A1(\mem[11][0] ), .A2(n782), .ZN(n217) );
  OAI21_X1 U135 ( .B1(n798), .B2(n216), .A(n218), .ZN(n479) );
  NAND2_X1 U136 ( .A1(\mem[11][1] ), .A2(n782), .ZN(n218) );
  OAI21_X1 U137 ( .B1(n799), .B2(n216), .A(n219), .ZN(n480) );
  NAND2_X1 U138 ( .A1(\mem[11][2] ), .A2(n782), .ZN(n219) );
  OAI21_X1 U139 ( .B1(n797), .B2(n233), .A(n234), .ZN(n494) );
  NAND2_X1 U140 ( .A1(\mem[12][0] ), .A2(n781), .ZN(n234) );
  OAI21_X1 U141 ( .B1(n798), .B2(n233), .A(n235), .ZN(n495) );
  NAND2_X1 U142 ( .A1(\mem[12][1] ), .A2(n781), .ZN(n235) );
  OAI21_X1 U143 ( .B1(n799), .B2(n233), .A(n236), .ZN(n496) );
  NAND2_X1 U144 ( .A1(\mem[12][2] ), .A2(n781), .ZN(n236) );
  OAI21_X1 U145 ( .B1(n797), .B2(n250), .A(n251), .ZN(n510) );
  NAND2_X1 U146 ( .A1(\mem[13][0] ), .A2(n780), .ZN(n251) );
  OAI21_X1 U147 ( .B1(n798), .B2(n250), .A(n252), .ZN(n511) );
  NAND2_X1 U148 ( .A1(\mem[13][1] ), .A2(n780), .ZN(n252) );
  OAI21_X1 U149 ( .B1(n799), .B2(n250), .A(n253), .ZN(n512) );
  NAND2_X1 U150 ( .A1(\mem[13][2] ), .A2(n780), .ZN(n253) );
  OAI21_X1 U151 ( .B1(n797), .B2(n267), .A(n268), .ZN(n526) );
  NAND2_X1 U152 ( .A1(\mem[14][0] ), .A2(n779), .ZN(n268) );
  OAI21_X1 U153 ( .B1(n798), .B2(n267), .A(n269), .ZN(n527) );
  NAND2_X1 U154 ( .A1(\mem[14][1] ), .A2(n779), .ZN(n269) );
  OAI21_X1 U155 ( .B1(n799), .B2(n267), .A(n270), .ZN(n528) );
  NAND2_X1 U156 ( .A1(\mem[14][2] ), .A2(n779), .ZN(n270) );
  OAI21_X1 U157 ( .B1(n797), .B2(n285), .A(n286), .ZN(n542) );
  NAND2_X1 U158 ( .A1(\mem[15][0] ), .A2(n778), .ZN(n286) );
  OAI21_X1 U159 ( .B1(n798), .B2(n285), .A(n287), .ZN(n543) );
  NAND2_X1 U160 ( .A1(\mem[15][1] ), .A2(n778), .ZN(n287) );
  OAI21_X1 U161 ( .B1(n799), .B2(n285), .A(n288), .ZN(n544) );
  NAND2_X1 U162 ( .A1(\mem[15][2] ), .A2(n778), .ZN(n288) );
  NOR2_X1 U163 ( .A1(n796), .A2(N13), .ZN(n145) );
  INV_X1 U164 ( .A(wr_en), .ZN(n796) );
  AND2_X1 U165 ( .A1(N12), .A2(n795), .ZN(n109) );
  AND2_X1 U166 ( .A1(N12), .A2(N11), .ZN(n144) );
  BUF_X1 U167 ( .A(N12), .Z(n763) );
  OAI21_X1 U168 ( .B1(n793), .B2(n801), .A(n25), .ZN(n306) );
  NAND2_X1 U169 ( .A1(\mem[0][4] ), .A2(n793), .ZN(n25) );
  OAI21_X1 U170 ( .B1(n793), .B2(n802), .A(n26), .ZN(n307) );
  NAND2_X1 U171 ( .A1(\mem[0][5] ), .A2(n793), .ZN(n26) );
  OAI21_X1 U172 ( .B1(n793), .B2(n803), .A(n27), .ZN(n308) );
  NAND2_X1 U173 ( .A1(\mem[0][6] ), .A2(n793), .ZN(n27) );
  OAI21_X1 U174 ( .B1(n793), .B2(n804), .A(n28), .ZN(n309) );
  NAND2_X1 U175 ( .A1(\mem[0][7] ), .A2(n793), .ZN(n28) );
  OAI21_X1 U176 ( .B1(n20), .B2(n805), .A(n29), .ZN(n310) );
  NAND2_X1 U177 ( .A1(\mem[0][8] ), .A2(n20), .ZN(n29) );
  OAI21_X1 U178 ( .B1(n20), .B2(n806), .A(n30), .ZN(n311) );
  NAND2_X1 U179 ( .A1(\mem[0][9] ), .A2(n20), .ZN(n30) );
  OAI21_X1 U180 ( .B1(n20), .B2(n807), .A(n31), .ZN(n312) );
  NAND2_X1 U181 ( .A1(\mem[0][10] ), .A2(n20), .ZN(n31) );
  OAI21_X1 U182 ( .B1(n20), .B2(n808), .A(n32), .ZN(n313) );
  NAND2_X1 U183 ( .A1(\mem[0][11] ), .A2(n20), .ZN(n32) );
  OAI21_X1 U184 ( .B1(n793), .B2(n809), .A(n33), .ZN(n314) );
  NAND2_X1 U185 ( .A1(\mem[0][12] ), .A2(n20), .ZN(n33) );
  OAI21_X1 U186 ( .B1(n20), .B2(n810), .A(n34), .ZN(n315) );
  NAND2_X1 U187 ( .A1(\mem[0][13] ), .A2(n20), .ZN(n34) );
  OAI21_X1 U188 ( .B1(n793), .B2(n812), .A(n36), .ZN(n317) );
  NAND2_X1 U189 ( .A1(\mem[0][15] ), .A2(n20), .ZN(n36) );
  OAI21_X1 U190 ( .B1(n793), .B2(n800), .A(n24), .ZN(n305) );
  NAND2_X1 U191 ( .A1(\mem[0][3] ), .A2(n793), .ZN(n24) );
  OAI21_X1 U192 ( .B1(n801), .B2(n39), .A(n44), .ZN(n322) );
  NAND2_X1 U193 ( .A1(\mem[1][4] ), .A2(n792), .ZN(n44) );
  OAI21_X1 U194 ( .B1(n802), .B2(n39), .A(n45), .ZN(n323) );
  NAND2_X1 U195 ( .A1(\mem[1][5] ), .A2(n39), .ZN(n45) );
  OAI21_X1 U196 ( .B1(n803), .B2(n39), .A(n46), .ZN(n324) );
  NAND2_X1 U197 ( .A1(\mem[1][6] ), .A2(n39), .ZN(n46) );
  OAI21_X1 U198 ( .B1(n804), .B2(n39), .A(n47), .ZN(n325) );
  NAND2_X1 U199 ( .A1(\mem[1][7] ), .A2(n39), .ZN(n47) );
  OAI21_X1 U200 ( .B1(n805), .B2(n39), .A(n48), .ZN(n326) );
  NAND2_X1 U201 ( .A1(\mem[1][8] ), .A2(n792), .ZN(n48) );
  OAI21_X1 U202 ( .B1(n806), .B2(n39), .A(n49), .ZN(n327) );
  NAND2_X1 U203 ( .A1(\mem[1][9] ), .A2(n792), .ZN(n49) );
  OAI21_X1 U204 ( .B1(n807), .B2(n792), .A(n50), .ZN(n328) );
  NAND2_X1 U205 ( .A1(\mem[1][10] ), .A2(n792), .ZN(n50) );
  OAI21_X1 U206 ( .B1(n808), .B2(n39), .A(n51), .ZN(n329) );
  NAND2_X1 U207 ( .A1(\mem[1][11] ), .A2(n792), .ZN(n51) );
  OAI21_X1 U208 ( .B1(n809), .B2(n39), .A(n52), .ZN(n330) );
  NAND2_X1 U209 ( .A1(\mem[1][12] ), .A2(n792), .ZN(n52) );
  OAI21_X1 U210 ( .B1(n810), .B2(n39), .A(n53), .ZN(n331) );
  NAND2_X1 U211 ( .A1(\mem[1][13] ), .A2(n792), .ZN(n53) );
  OAI21_X1 U212 ( .B1(n812), .B2(n39), .A(n55), .ZN(n333) );
  NAND2_X1 U213 ( .A1(\mem[1][15] ), .A2(n792), .ZN(n55) );
  OAI21_X1 U214 ( .B1(n801), .B2(n57), .A(n62), .ZN(n338) );
  NAND2_X1 U215 ( .A1(\mem[2][4] ), .A2(n791), .ZN(n62) );
  OAI21_X1 U216 ( .B1(n802), .B2(n57), .A(n63), .ZN(n339) );
  NAND2_X1 U217 ( .A1(\mem[2][5] ), .A2(n57), .ZN(n63) );
  OAI21_X1 U218 ( .B1(n803), .B2(n57), .A(n64), .ZN(n340) );
  NAND2_X1 U219 ( .A1(\mem[2][6] ), .A2(n57), .ZN(n64) );
  OAI21_X1 U220 ( .B1(n804), .B2(n57), .A(n65), .ZN(n341) );
  NAND2_X1 U221 ( .A1(\mem[2][7] ), .A2(n57), .ZN(n65) );
  OAI21_X1 U222 ( .B1(n805), .B2(n57), .A(n66), .ZN(n342) );
  NAND2_X1 U223 ( .A1(\mem[2][8] ), .A2(n791), .ZN(n66) );
  OAI21_X1 U224 ( .B1(n806), .B2(n57), .A(n67), .ZN(n343) );
  NAND2_X1 U225 ( .A1(\mem[2][9] ), .A2(n791), .ZN(n67) );
  OAI21_X1 U226 ( .B1(n807), .B2(n791), .A(n68), .ZN(n344) );
  NAND2_X1 U227 ( .A1(\mem[2][10] ), .A2(n791), .ZN(n68) );
  OAI21_X1 U228 ( .B1(n808), .B2(n57), .A(n69), .ZN(n345) );
  NAND2_X1 U229 ( .A1(\mem[2][11] ), .A2(n791), .ZN(n69) );
  OAI21_X1 U230 ( .B1(n809), .B2(n57), .A(n70), .ZN(n346) );
  NAND2_X1 U231 ( .A1(\mem[2][12] ), .A2(n791), .ZN(n70) );
  OAI21_X1 U232 ( .B1(n810), .B2(n57), .A(n71), .ZN(n347) );
  NAND2_X1 U233 ( .A1(\mem[2][13] ), .A2(n791), .ZN(n71) );
  OAI21_X1 U234 ( .B1(n812), .B2(n57), .A(n73), .ZN(n349) );
  NAND2_X1 U235 ( .A1(\mem[2][15] ), .A2(n791), .ZN(n73) );
  OAI21_X1 U236 ( .B1(n801), .B2(n75), .A(n80), .ZN(n354) );
  NAND2_X1 U237 ( .A1(\mem[3][4] ), .A2(n790), .ZN(n80) );
  OAI21_X1 U238 ( .B1(n802), .B2(n75), .A(n81), .ZN(n355) );
  NAND2_X1 U239 ( .A1(\mem[3][5] ), .A2(n75), .ZN(n81) );
  OAI21_X1 U240 ( .B1(n803), .B2(n75), .A(n82), .ZN(n356) );
  NAND2_X1 U241 ( .A1(\mem[3][6] ), .A2(n75), .ZN(n82) );
  OAI21_X1 U242 ( .B1(n804), .B2(n75), .A(n83), .ZN(n357) );
  NAND2_X1 U243 ( .A1(\mem[3][7] ), .A2(n75), .ZN(n83) );
  OAI21_X1 U244 ( .B1(n805), .B2(n75), .A(n84), .ZN(n358) );
  NAND2_X1 U245 ( .A1(\mem[3][8] ), .A2(n790), .ZN(n84) );
  OAI21_X1 U246 ( .B1(n806), .B2(n75), .A(n85), .ZN(n359) );
  NAND2_X1 U247 ( .A1(\mem[3][9] ), .A2(n790), .ZN(n85) );
  OAI21_X1 U248 ( .B1(n807), .B2(n790), .A(n86), .ZN(n360) );
  NAND2_X1 U249 ( .A1(\mem[3][10] ), .A2(n790), .ZN(n86) );
  OAI21_X1 U250 ( .B1(n808), .B2(n75), .A(n87), .ZN(n361) );
  NAND2_X1 U251 ( .A1(\mem[3][11] ), .A2(n790), .ZN(n87) );
  OAI21_X1 U252 ( .B1(n809), .B2(n75), .A(n88), .ZN(n362) );
  NAND2_X1 U253 ( .A1(\mem[3][12] ), .A2(n790), .ZN(n88) );
  OAI21_X1 U254 ( .B1(n810), .B2(n75), .A(n89), .ZN(n363) );
  NAND2_X1 U255 ( .A1(\mem[3][13] ), .A2(n790), .ZN(n89) );
  OAI21_X1 U256 ( .B1(n812), .B2(n75), .A(n91), .ZN(n365) );
  NAND2_X1 U257 ( .A1(\mem[3][15] ), .A2(n790), .ZN(n91) );
  OAI21_X1 U258 ( .B1(n801), .B2(n92), .A(n97), .ZN(n370) );
  NAND2_X1 U259 ( .A1(\mem[4][4] ), .A2(n789), .ZN(n97) );
  OAI21_X1 U260 ( .B1(n802), .B2(n92), .A(n98), .ZN(n371) );
  NAND2_X1 U261 ( .A1(\mem[4][5] ), .A2(n92), .ZN(n98) );
  OAI21_X1 U262 ( .B1(n803), .B2(n92), .A(n99), .ZN(n372) );
  NAND2_X1 U263 ( .A1(\mem[4][6] ), .A2(n92), .ZN(n99) );
  OAI21_X1 U264 ( .B1(n804), .B2(n92), .A(n100), .ZN(n373) );
  NAND2_X1 U265 ( .A1(\mem[4][7] ), .A2(n92), .ZN(n100) );
  OAI21_X1 U266 ( .B1(n805), .B2(n92), .A(n101), .ZN(n374) );
  NAND2_X1 U267 ( .A1(\mem[4][8] ), .A2(n789), .ZN(n101) );
  OAI21_X1 U268 ( .B1(n806), .B2(n92), .A(n102), .ZN(n375) );
  NAND2_X1 U269 ( .A1(\mem[4][9] ), .A2(n789), .ZN(n102) );
  OAI21_X1 U270 ( .B1(n807), .B2(n789), .A(n103), .ZN(n376) );
  NAND2_X1 U271 ( .A1(\mem[4][10] ), .A2(n789), .ZN(n103) );
  OAI21_X1 U272 ( .B1(n808), .B2(n92), .A(n104), .ZN(n377) );
  NAND2_X1 U273 ( .A1(\mem[4][11] ), .A2(n789), .ZN(n104) );
  OAI21_X1 U274 ( .B1(n809), .B2(n92), .A(n105), .ZN(n378) );
  NAND2_X1 U275 ( .A1(\mem[4][12] ), .A2(n789), .ZN(n105) );
  OAI21_X1 U276 ( .B1(n810), .B2(n92), .A(n106), .ZN(n379) );
  NAND2_X1 U277 ( .A1(\mem[4][13] ), .A2(n789), .ZN(n106) );
  OAI21_X1 U278 ( .B1(n812), .B2(n92), .A(n108), .ZN(n381) );
  NAND2_X1 U279 ( .A1(\mem[4][15] ), .A2(n789), .ZN(n108) );
  OAI21_X1 U280 ( .B1(n801), .B2(n110), .A(n115), .ZN(n386) );
  NAND2_X1 U281 ( .A1(\mem[5][4] ), .A2(n788), .ZN(n115) );
  OAI21_X1 U282 ( .B1(n802), .B2(n110), .A(n116), .ZN(n387) );
  NAND2_X1 U283 ( .A1(\mem[5][5] ), .A2(n788), .ZN(n116) );
  OAI21_X1 U284 ( .B1(n803), .B2(n110), .A(n117), .ZN(n388) );
  NAND2_X1 U285 ( .A1(\mem[5][6] ), .A2(n788), .ZN(n117) );
  OAI21_X1 U286 ( .B1(n804), .B2(n788), .A(n118), .ZN(n389) );
  NAND2_X1 U287 ( .A1(\mem[5][7] ), .A2(n788), .ZN(n118) );
  OAI21_X1 U288 ( .B1(n805), .B2(n788), .A(n119), .ZN(n390) );
  NAND2_X1 U289 ( .A1(\mem[5][8] ), .A2(n110), .ZN(n119) );
  OAI21_X1 U290 ( .B1(n806), .B2(n788), .A(n120), .ZN(n391) );
  NAND2_X1 U291 ( .A1(\mem[5][9] ), .A2(n110), .ZN(n120) );
  OAI21_X1 U292 ( .B1(n807), .B2(n788), .A(n121), .ZN(n392) );
  NAND2_X1 U293 ( .A1(\mem[5][10] ), .A2(n110), .ZN(n121) );
  OAI21_X1 U294 ( .B1(n808), .B2(n788), .A(n122), .ZN(n393) );
  NAND2_X1 U295 ( .A1(\mem[5][11] ), .A2(n110), .ZN(n122) );
  OAI21_X1 U296 ( .B1(n809), .B2(n788), .A(n123), .ZN(n394) );
  NAND2_X1 U297 ( .A1(\mem[5][12] ), .A2(n110), .ZN(n123) );
  OAI21_X1 U298 ( .B1(n810), .B2(n788), .A(n124), .ZN(n395) );
  NAND2_X1 U299 ( .A1(\mem[5][13] ), .A2(n110), .ZN(n124) );
  OAI21_X1 U300 ( .B1(n812), .B2(n110), .A(n126), .ZN(n397) );
  NAND2_X1 U301 ( .A1(\mem[5][15] ), .A2(n110), .ZN(n126) );
  OAI21_X1 U302 ( .B1(n801), .B2(n127), .A(n132), .ZN(n402) );
  NAND2_X1 U303 ( .A1(\mem[6][4] ), .A2(n787), .ZN(n132) );
  OAI21_X1 U304 ( .B1(n802), .B2(n127), .A(n133), .ZN(n403) );
  NAND2_X1 U305 ( .A1(\mem[6][5] ), .A2(n127), .ZN(n133) );
  OAI21_X1 U306 ( .B1(n803), .B2(n127), .A(n134), .ZN(n404) );
  NAND2_X1 U307 ( .A1(\mem[6][6] ), .A2(n127), .ZN(n134) );
  OAI21_X1 U308 ( .B1(n804), .B2(n127), .A(n135), .ZN(n405) );
  NAND2_X1 U309 ( .A1(\mem[6][7] ), .A2(n127), .ZN(n135) );
  OAI21_X1 U310 ( .B1(n805), .B2(n127), .A(n136), .ZN(n406) );
  NAND2_X1 U311 ( .A1(\mem[6][8] ), .A2(n787), .ZN(n136) );
  OAI21_X1 U312 ( .B1(n806), .B2(n127), .A(n137), .ZN(n407) );
  NAND2_X1 U313 ( .A1(\mem[6][9] ), .A2(n787), .ZN(n137) );
  OAI21_X1 U314 ( .B1(n807), .B2(n787), .A(n138), .ZN(n408) );
  NAND2_X1 U315 ( .A1(\mem[6][10] ), .A2(n787), .ZN(n138) );
  OAI21_X1 U316 ( .B1(n808), .B2(n127), .A(n139), .ZN(n409) );
  NAND2_X1 U317 ( .A1(\mem[6][11] ), .A2(n787), .ZN(n139) );
  OAI21_X1 U318 ( .B1(n809), .B2(n127), .A(n140), .ZN(n410) );
  NAND2_X1 U319 ( .A1(\mem[6][12] ), .A2(n787), .ZN(n140) );
  OAI21_X1 U320 ( .B1(n810), .B2(n127), .A(n141), .ZN(n411) );
  NAND2_X1 U321 ( .A1(\mem[6][13] ), .A2(n787), .ZN(n141) );
  OAI21_X1 U322 ( .B1(n812), .B2(n127), .A(n143), .ZN(n413) );
  NAND2_X1 U323 ( .A1(\mem[6][15] ), .A2(n787), .ZN(n143) );
  OAI21_X1 U324 ( .B1(n801), .B2(n146), .A(n151), .ZN(n418) );
  NAND2_X1 U325 ( .A1(\mem[7][4] ), .A2(n786), .ZN(n151) );
  OAI21_X1 U326 ( .B1(n802), .B2(n146), .A(n152), .ZN(n419) );
  NAND2_X1 U327 ( .A1(\mem[7][5] ), .A2(n146), .ZN(n152) );
  OAI21_X1 U328 ( .B1(n803), .B2(n146), .A(n153), .ZN(n420) );
  NAND2_X1 U329 ( .A1(\mem[7][6] ), .A2(n146), .ZN(n153) );
  OAI21_X1 U330 ( .B1(n804), .B2(n146), .A(n154), .ZN(n421) );
  NAND2_X1 U331 ( .A1(\mem[7][7] ), .A2(n146), .ZN(n154) );
  OAI21_X1 U332 ( .B1(n805), .B2(n146), .A(n155), .ZN(n422) );
  NAND2_X1 U333 ( .A1(\mem[7][8] ), .A2(n786), .ZN(n155) );
  OAI21_X1 U334 ( .B1(n806), .B2(n146), .A(n156), .ZN(n423) );
  NAND2_X1 U335 ( .A1(\mem[7][9] ), .A2(n786), .ZN(n156) );
  OAI21_X1 U336 ( .B1(n807), .B2(n786), .A(n157), .ZN(n424) );
  NAND2_X1 U337 ( .A1(\mem[7][10] ), .A2(n786), .ZN(n157) );
  OAI21_X1 U338 ( .B1(n808), .B2(n146), .A(n158), .ZN(n425) );
  NAND2_X1 U339 ( .A1(\mem[7][11] ), .A2(n786), .ZN(n158) );
  OAI21_X1 U340 ( .B1(n809), .B2(n146), .A(n159), .ZN(n426) );
  NAND2_X1 U341 ( .A1(\mem[7][12] ), .A2(n786), .ZN(n159) );
  OAI21_X1 U342 ( .B1(n810), .B2(n146), .A(n160), .ZN(n427) );
  NAND2_X1 U343 ( .A1(\mem[7][13] ), .A2(n786), .ZN(n160) );
  OAI21_X1 U344 ( .B1(n812), .B2(n146), .A(n162), .ZN(n429) );
  NAND2_X1 U345 ( .A1(\mem[7][15] ), .A2(n786), .ZN(n162) );
  OAI21_X1 U346 ( .B1(n801), .B2(n163), .A(n168), .ZN(n434) );
  NAND2_X1 U347 ( .A1(\mem[8][4] ), .A2(n785), .ZN(n168) );
  OAI21_X1 U348 ( .B1(n802), .B2(n163), .A(n169), .ZN(n435) );
  NAND2_X1 U349 ( .A1(\mem[8][5] ), .A2(n163), .ZN(n169) );
  OAI21_X1 U350 ( .B1(n803), .B2(n163), .A(n170), .ZN(n436) );
  NAND2_X1 U351 ( .A1(\mem[8][6] ), .A2(n163), .ZN(n170) );
  OAI21_X1 U352 ( .B1(n804), .B2(n163), .A(n171), .ZN(n437) );
  NAND2_X1 U353 ( .A1(\mem[8][7] ), .A2(n163), .ZN(n171) );
  OAI21_X1 U354 ( .B1(n805), .B2(n163), .A(n172), .ZN(n438) );
  NAND2_X1 U355 ( .A1(\mem[8][8] ), .A2(n785), .ZN(n172) );
  OAI21_X1 U356 ( .B1(n806), .B2(n163), .A(n173), .ZN(n439) );
  NAND2_X1 U357 ( .A1(\mem[8][9] ), .A2(n785), .ZN(n173) );
  OAI21_X1 U358 ( .B1(n807), .B2(n785), .A(n174), .ZN(n440) );
  NAND2_X1 U359 ( .A1(\mem[8][10] ), .A2(n785), .ZN(n174) );
  OAI21_X1 U360 ( .B1(n808), .B2(n163), .A(n175), .ZN(n441) );
  NAND2_X1 U361 ( .A1(\mem[8][11] ), .A2(n785), .ZN(n175) );
  OAI21_X1 U362 ( .B1(n809), .B2(n163), .A(n176), .ZN(n442) );
  NAND2_X1 U363 ( .A1(\mem[8][12] ), .A2(n785), .ZN(n176) );
  OAI21_X1 U364 ( .B1(n810), .B2(n163), .A(n177), .ZN(n443) );
  NAND2_X1 U365 ( .A1(\mem[8][13] ), .A2(n785), .ZN(n177) );
  OAI21_X1 U366 ( .B1(n812), .B2(n163), .A(n179), .ZN(n445) );
  NAND2_X1 U367 ( .A1(\mem[8][15] ), .A2(n785), .ZN(n179) );
  OAI21_X1 U368 ( .B1(n801), .B2(n181), .A(n186), .ZN(n450) );
  NAND2_X1 U369 ( .A1(\mem[9][4] ), .A2(n784), .ZN(n186) );
  OAI21_X1 U370 ( .B1(n802), .B2(n181), .A(n187), .ZN(n451) );
  NAND2_X1 U371 ( .A1(\mem[9][5] ), .A2(n181), .ZN(n187) );
  OAI21_X1 U372 ( .B1(n803), .B2(n181), .A(n188), .ZN(n452) );
  NAND2_X1 U373 ( .A1(\mem[9][6] ), .A2(n181), .ZN(n188) );
  OAI21_X1 U374 ( .B1(n804), .B2(n181), .A(n189), .ZN(n453) );
  NAND2_X1 U375 ( .A1(\mem[9][7] ), .A2(n181), .ZN(n189) );
  OAI21_X1 U376 ( .B1(n805), .B2(n181), .A(n190), .ZN(n454) );
  NAND2_X1 U377 ( .A1(\mem[9][8] ), .A2(n784), .ZN(n190) );
  OAI21_X1 U378 ( .B1(n806), .B2(n181), .A(n191), .ZN(n455) );
  NAND2_X1 U379 ( .A1(\mem[9][9] ), .A2(n784), .ZN(n191) );
  OAI21_X1 U380 ( .B1(n807), .B2(n784), .A(n192), .ZN(n456) );
  NAND2_X1 U381 ( .A1(\mem[9][10] ), .A2(n784), .ZN(n192) );
  OAI21_X1 U382 ( .B1(n808), .B2(n181), .A(n193), .ZN(n457) );
  NAND2_X1 U383 ( .A1(\mem[9][11] ), .A2(n784), .ZN(n193) );
  OAI21_X1 U384 ( .B1(n809), .B2(n181), .A(n194), .ZN(n458) );
  NAND2_X1 U385 ( .A1(\mem[9][12] ), .A2(n784), .ZN(n194) );
  OAI21_X1 U386 ( .B1(n810), .B2(n181), .A(n195), .ZN(n459) );
  NAND2_X1 U387 ( .A1(\mem[9][13] ), .A2(n784), .ZN(n195) );
  OAI21_X1 U388 ( .B1(n812), .B2(n181), .A(n197), .ZN(n461) );
  NAND2_X1 U389 ( .A1(\mem[9][15] ), .A2(n784), .ZN(n197) );
  OAI21_X1 U390 ( .B1(n801), .B2(n199), .A(n204), .ZN(n466) );
  NAND2_X1 U391 ( .A1(\mem[10][4] ), .A2(n783), .ZN(n204) );
  OAI21_X1 U392 ( .B1(n802), .B2(n199), .A(n205), .ZN(n467) );
  NAND2_X1 U393 ( .A1(\mem[10][5] ), .A2(n199), .ZN(n205) );
  OAI21_X1 U394 ( .B1(n803), .B2(n199), .A(n206), .ZN(n468) );
  NAND2_X1 U395 ( .A1(\mem[10][6] ), .A2(n199), .ZN(n206) );
  OAI21_X1 U396 ( .B1(n804), .B2(n199), .A(n207), .ZN(n469) );
  NAND2_X1 U397 ( .A1(\mem[10][7] ), .A2(n199), .ZN(n207) );
  OAI21_X1 U398 ( .B1(n805), .B2(n199), .A(n208), .ZN(n470) );
  NAND2_X1 U399 ( .A1(\mem[10][8] ), .A2(n783), .ZN(n208) );
  OAI21_X1 U400 ( .B1(n806), .B2(n199), .A(n209), .ZN(n471) );
  NAND2_X1 U401 ( .A1(\mem[10][9] ), .A2(n783), .ZN(n209) );
  OAI21_X1 U402 ( .B1(n807), .B2(n783), .A(n210), .ZN(n472) );
  NAND2_X1 U403 ( .A1(\mem[10][10] ), .A2(n783), .ZN(n210) );
  OAI21_X1 U404 ( .B1(n808), .B2(n199), .A(n211), .ZN(n473) );
  NAND2_X1 U405 ( .A1(\mem[10][11] ), .A2(n783), .ZN(n211) );
  OAI21_X1 U406 ( .B1(n809), .B2(n199), .A(n212), .ZN(n474) );
  NAND2_X1 U407 ( .A1(\mem[10][12] ), .A2(n783), .ZN(n212) );
  OAI21_X1 U408 ( .B1(n810), .B2(n199), .A(n213), .ZN(n475) );
  NAND2_X1 U409 ( .A1(\mem[10][13] ), .A2(n783), .ZN(n213) );
  OAI21_X1 U410 ( .B1(n812), .B2(n199), .A(n215), .ZN(n477) );
  NAND2_X1 U411 ( .A1(\mem[10][15] ), .A2(n783), .ZN(n215) );
  OAI21_X1 U412 ( .B1(n801), .B2(n216), .A(n221), .ZN(n482) );
  NAND2_X1 U413 ( .A1(\mem[11][4] ), .A2(n782), .ZN(n221) );
  OAI21_X1 U414 ( .B1(n802), .B2(n216), .A(n222), .ZN(n483) );
  NAND2_X1 U415 ( .A1(\mem[11][5] ), .A2(n216), .ZN(n222) );
  OAI21_X1 U416 ( .B1(n803), .B2(n216), .A(n223), .ZN(n484) );
  NAND2_X1 U417 ( .A1(\mem[11][6] ), .A2(n216), .ZN(n223) );
  OAI21_X1 U418 ( .B1(n804), .B2(n216), .A(n224), .ZN(n485) );
  NAND2_X1 U419 ( .A1(\mem[11][7] ), .A2(n216), .ZN(n224) );
  OAI21_X1 U420 ( .B1(n805), .B2(n216), .A(n225), .ZN(n486) );
  NAND2_X1 U421 ( .A1(\mem[11][8] ), .A2(n782), .ZN(n225) );
  OAI21_X1 U422 ( .B1(n806), .B2(n216), .A(n226), .ZN(n487) );
  NAND2_X1 U423 ( .A1(\mem[11][9] ), .A2(n782), .ZN(n226) );
  OAI21_X1 U424 ( .B1(n807), .B2(n782), .A(n227), .ZN(n488) );
  NAND2_X1 U425 ( .A1(\mem[11][10] ), .A2(n782), .ZN(n227) );
  OAI21_X1 U426 ( .B1(n808), .B2(n216), .A(n228), .ZN(n489) );
  NAND2_X1 U427 ( .A1(\mem[11][11] ), .A2(n782), .ZN(n228) );
  OAI21_X1 U428 ( .B1(n809), .B2(n216), .A(n229), .ZN(n490) );
  NAND2_X1 U429 ( .A1(\mem[11][12] ), .A2(n782), .ZN(n229) );
  OAI21_X1 U430 ( .B1(n810), .B2(n216), .A(n230), .ZN(n491) );
  NAND2_X1 U431 ( .A1(\mem[11][13] ), .A2(n782), .ZN(n230) );
  OAI21_X1 U432 ( .B1(n812), .B2(n216), .A(n232), .ZN(n493) );
  NAND2_X1 U433 ( .A1(\mem[11][15] ), .A2(n782), .ZN(n232) );
  OAI21_X1 U434 ( .B1(n801), .B2(n233), .A(n238), .ZN(n498) );
  NAND2_X1 U435 ( .A1(\mem[12][4] ), .A2(n781), .ZN(n238) );
  OAI21_X1 U436 ( .B1(n802), .B2(n233), .A(n239), .ZN(n499) );
  NAND2_X1 U437 ( .A1(\mem[12][5] ), .A2(n233), .ZN(n239) );
  OAI21_X1 U438 ( .B1(n803), .B2(n233), .A(n240), .ZN(n500) );
  NAND2_X1 U439 ( .A1(\mem[12][6] ), .A2(n233), .ZN(n240) );
  OAI21_X1 U440 ( .B1(n804), .B2(n233), .A(n241), .ZN(n501) );
  NAND2_X1 U441 ( .A1(\mem[12][7] ), .A2(n233), .ZN(n241) );
  OAI21_X1 U442 ( .B1(n805), .B2(n233), .A(n242), .ZN(n502) );
  NAND2_X1 U443 ( .A1(\mem[12][8] ), .A2(n781), .ZN(n242) );
  OAI21_X1 U444 ( .B1(n806), .B2(n233), .A(n243), .ZN(n503) );
  NAND2_X1 U445 ( .A1(\mem[12][9] ), .A2(n781), .ZN(n243) );
  OAI21_X1 U446 ( .B1(n807), .B2(n781), .A(n244), .ZN(n504) );
  NAND2_X1 U447 ( .A1(\mem[12][10] ), .A2(n781), .ZN(n244) );
  OAI21_X1 U448 ( .B1(n808), .B2(n233), .A(n245), .ZN(n505) );
  NAND2_X1 U449 ( .A1(\mem[12][11] ), .A2(n781), .ZN(n245) );
  OAI21_X1 U450 ( .B1(n809), .B2(n233), .A(n246), .ZN(n506) );
  NAND2_X1 U451 ( .A1(\mem[12][12] ), .A2(n781), .ZN(n246) );
  OAI21_X1 U452 ( .B1(n810), .B2(n233), .A(n247), .ZN(n507) );
  NAND2_X1 U453 ( .A1(\mem[12][13] ), .A2(n781), .ZN(n247) );
  OAI21_X1 U454 ( .B1(n812), .B2(n233), .A(n249), .ZN(n509) );
  NAND2_X1 U455 ( .A1(\mem[12][15] ), .A2(n781), .ZN(n249) );
  OAI21_X1 U456 ( .B1(n801), .B2(n250), .A(n255), .ZN(n514) );
  NAND2_X1 U457 ( .A1(\mem[13][4] ), .A2(n780), .ZN(n255) );
  OAI21_X1 U458 ( .B1(n802), .B2(n250), .A(n256), .ZN(n515) );
  NAND2_X1 U459 ( .A1(\mem[13][5] ), .A2(n250), .ZN(n256) );
  OAI21_X1 U460 ( .B1(n803), .B2(n250), .A(n257), .ZN(n516) );
  NAND2_X1 U461 ( .A1(\mem[13][6] ), .A2(n250), .ZN(n257) );
  OAI21_X1 U462 ( .B1(n804), .B2(n250), .A(n258), .ZN(n517) );
  NAND2_X1 U463 ( .A1(\mem[13][7] ), .A2(n250), .ZN(n258) );
  OAI21_X1 U464 ( .B1(n805), .B2(n250), .A(n259), .ZN(n518) );
  NAND2_X1 U465 ( .A1(\mem[13][8] ), .A2(n780), .ZN(n259) );
  OAI21_X1 U466 ( .B1(n806), .B2(n250), .A(n260), .ZN(n519) );
  NAND2_X1 U467 ( .A1(\mem[13][9] ), .A2(n780), .ZN(n260) );
  OAI21_X1 U468 ( .B1(n807), .B2(n780), .A(n261), .ZN(n520) );
  NAND2_X1 U469 ( .A1(\mem[13][10] ), .A2(n780), .ZN(n261) );
  OAI21_X1 U470 ( .B1(n808), .B2(n250), .A(n262), .ZN(n521) );
  NAND2_X1 U471 ( .A1(\mem[13][11] ), .A2(n780), .ZN(n262) );
  OAI21_X1 U472 ( .B1(n809), .B2(n250), .A(n263), .ZN(n522) );
  NAND2_X1 U473 ( .A1(\mem[13][12] ), .A2(n780), .ZN(n263) );
  OAI21_X1 U474 ( .B1(n810), .B2(n250), .A(n264), .ZN(n523) );
  NAND2_X1 U475 ( .A1(\mem[13][13] ), .A2(n780), .ZN(n264) );
  OAI21_X1 U476 ( .B1(n812), .B2(n250), .A(n266), .ZN(n525) );
  NAND2_X1 U477 ( .A1(\mem[13][15] ), .A2(n780), .ZN(n266) );
  OAI21_X1 U478 ( .B1(n801), .B2(n267), .A(n272), .ZN(n530) );
  NAND2_X1 U479 ( .A1(\mem[14][4] ), .A2(n779), .ZN(n272) );
  OAI21_X1 U480 ( .B1(n802), .B2(n267), .A(n273), .ZN(n531) );
  NAND2_X1 U481 ( .A1(\mem[14][5] ), .A2(n267), .ZN(n273) );
  OAI21_X1 U482 ( .B1(n803), .B2(n267), .A(n274), .ZN(n532) );
  NAND2_X1 U483 ( .A1(\mem[14][6] ), .A2(n267), .ZN(n274) );
  OAI21_X1 U484 ( .B1(n804), .B2(n267), .A(n275), .ZN(n533) );
  NAND2_X1 U485 ( .A1(\mem[14][7] ), .A2(n267), .ZN(n275) );
  OAI21_X1 U486 ( .B1(n805), .B2(n267), .A(n276), .ZN(n534) );
  NAND2_X1 U487 ( .A1(\mem[14][8] ), .A2(n779), .ZN(n276) );
  OAI21_X1 U488 ( .B1(n806), .B2(n267), .A(n277), .ZN(n535) );
  NAND2_X1 U489 ( .A1(\mem[14][9] ), .A2(n779), .ZN(n277) );
  OAI21_X1 U490 ( .B1(n807), .B2(n779), .A(n278), .ZN(n536) );
  NAND2_X1 U491 ( .A1(\mem[14][10] ), .A2(n779), .ZN(n278) );
  OAI21_X1 U492 ( .B1(n808), .B2(n267), .A(n279), .ZN(n537) );
  NAND2_X1 U493 ( .A1(\mem[14][11] ), .A2(n779), .ZN(n279) );
  OAI21_X1 U494 ( .B1(n809), .B2(n267), .A(n280), .ZN(n538) );
  NAND2_X1 U495 ( .A1(\mem[14][12] ), .A2(n779), .ZN(n280) );
  OAI21_X1 U496 ( .B1(n810), .B2(n267), .A(n281), .ZN(n539) );
  NAND2_X1 U497 ( .A1(\mem[14][13] ), .A2(n779), .ZN(n281) );
  OAI21_X1 U498 ( .B1(n812), .B2(n267), .A(n283), .ZN(n541) );
  NAND2_X1 U499 ( .A1(\mem[14][15] ), .A2(n779), .ZN(n283) );
  OAI21_X1 U500 ( .B1(n801), .B2(n285), .A(n290), .ZN(n546) );
  NAND2_X1 U501 ( .A1(\mem[15][4] ), .A2(n778), .ZN(n290) );
  OAI21_X1 U502 ( .B1(n802), .B2(n285), .A(n291), .ZN(n547) );
  NAND2_X1 U503 ( .A1(\mem[15][5] ), .A2(n285), .ZN(n291) );
  OAI21_X1 U504 ( .B1(n803), .B2(n285), .A(n292), .ZN(n548) );
  NAND2_X1 U505 ( .A1(\mem[15][6] ), .A2(n285), .ZN(n292) );
  OAI21_X1 U506 ( .B1(n804), .B2(n285), .A(n293), .ZN(n549) );
  NAND2_X1 U507 ( .A1(\mem[15][7] ), .A2(n285), .ZN(n293) );
  OAI21_X1 U508 ( .B1(n805), .B2(n285), .A(n294), .ZN(n550) );
  NAND2_X1 U509 ( .A1(\mem[15][8] ), .A2(n778), .ZN(n294) );
  OAI21_X1 U510 ( .B1(n806), .B2(n285), .A(n295), .ZN(n551) );
  NAND2_X1 U511 ( .A1(\mem[15][9] ), .A2(n778), .ZN(n295) );
  OAI21_X1 U512 ( .B1(n807), .B2(n778), .A(n296), .ZN(n552) );
  NAND2_X1 U513 ( .A1(\mem[15][10] ), .A2(n778), .ZN(n296) );
  OAI21_X1 U514 ( .B1(n808), .B2(n285), .A(n297), .ZN(n553) );
  NAND2_X1 U515 ( .A1(\mem[15][11] ), .A2(n778), .ZN(n297) );
  OAI21_X1 U516 ( .B1(n809), .B2(n285), .A(n298), .ZN(n554) );
  NAND2_X1 U517 ( .A1(\mem[15][12] ), .A2(n778), .ZN(n298) );
  OAI21_X1 U518 ( .B1(n810), .B2(n285), .A(n299), .ZN(n555) );
  NAND2_X1 U519 ( .A1(\mem[15][13] ), .A2(n778), .ZN(n299) );
  OAI21_X1 U520 ( .B1(n812), .B2(n285), .A(n301), .ZN(n557) );
  NAND2_X1 U521 ( .A1(\mem[15][15] ), .A2(n778), .ZN(n301) );
  OAI21_X1 U522 ( .B1(n800), .B2(n39), .A(n43), .ZN(n321) );
  NAND2_X1 U523 ( .A1(\mem[1][3] ), .A2(n792), .ZN(n43) );
  OAI21_X1 U524 ( .B1(n800), .B2(n57), .A(n61), .ZN(n337) );
  NAND2_X1 U525 ( .A1(\mem[2][3] ), .A2(n791), .ZN(n61) );
  OAI21_X1 U526 ( .B1(n800), .B2(n75), .A(n79), .ZN(n353) );
  NAND2_X1 U527 ( .A1(\mem[3][3] ), .A2(n790), .ZN(n79) );
  OAI21_X1 U528 ( .B1(n800), .B2(n92), .A(n96), .ZN(n369) );
  NAND2_X1 U529 ( .A1(\mem[4][3] ), .A2(n789), .ZN(n96) );
  OAI21_X1 U530 ( .B1(n800), .B2(n788), .A(n114), .ZN(n385) );
  NAND2_X1 U531 ( .A1(\mem[5][3] ), .A2(n788), .ZN(n114) );
  OAI21_X1 U532 ( .B1(n800), .B2(n127), .A(n131), .ZN(n401) );
  NAND2_X1 U533 ( .A1(\mem[6][3] ), .A2(n787), .ZN(n131) );
  OAI21_X1 U534 ( .B1(n800), .B2(n146), .A(n150), .ZN(n417) );
  NAND2_X1 U535 ( .A1(\mem[7][3] ), .A2(n786), .ZN(n150) );
  OAI21_X1 U536 ( .B1(n800), .B2(n163), .A(n167), .ZN(n433) );
  NAND2_X1 U537 ( .A1(\mem[8][3] ), .A2(n785), .ZN(n167) );
  OAI21_X1 U538 ( .B1(n800), .B2(n181), .A(n185), .ZN(n449) );
  NAND2_X1 U539 ( .A1(\mem[9][3] ), .A2(n784), .ZN(n185) );
  OAI21_X1 U540 ( .B1(n800), .B2(n199), .A(n203), .ZN(n465) );
  NAND2_X1 U541 ( .A1(\mem[10][3] ), .A2(n783), .ZN(n203) );
  OAI21_X1 U542 ( .B1(n800), .B2(n216), .A(n220), .ZN(n481) );
  NAND2_X1 U543 ( .A1(\mem[11][3] ), .A2(n782), .ZN(n220) );
  OAI21_X1 U544 ( .B1(n800), .B2(n233), .A(n237), .ZN(n497) );
  NAND2_X1 U545 ( .A1(\mem[12][3] ), .A2(n781), .ZN(n237) );
  OAI21_X1 U546 ( .B1(n800), .B2(n250), .A(n254), .ZN(n513) );
  NAND2_X1 U547 ( .A1(\mem[13][3] ), .A2(n780), .ZN(n254) );
  OAI21_X1 U548 ( .B1(n800), .B2(n267), .A(n271), .ZN(n529) );
  NAND2_X1 U549 ( .A1(\mem[14][3] ), .A2(n779), .ZN(n271) );
  OAI21_X1 U550 ( .B1(n800), .B2(n285), .A(n289), .ZN(n545) );
  NAND2_X1 U551 ( .A1(\mem[15][3] ), .A2(n778), .ZN(n289) );
  OAI21_X1 U552 ( .B1(n811), .B2(n57), .A(n72), .ZN(n348) );
  NAND2_X1 U553 ( .A1(\mem[2][14] ), .A2(n791), .ZN(n72) );
  OAI21_X1 U554 ( .B1(n811), .B2(n75), .A(n90), .ZN(n364) );
  NAND2_X1 U555 ( .A1(\mem[3][14] ), .A2(n790), .ZN(n90) );
  OAI21_X1 U556 ( .B1(n811), .B2(n39), .A(n54), .ZN(n332) );
  NAND2_X1 U557 ( .A1(\mem[1][14] ), .A2(n792), .ZN(n54) );
  OAI21_X1 U558 ( .B1(n811), .B2(n92), .A(n107), .ZN(n380) );
  NAND2_X1 U559 ( .A1(\mem[4][14] ), .A2(n789), .ZN(n107) );
  OAI21_X1 U560 ( .B1(n811), .B2(n788), .A(n125), .ZN(n396) );
  NAND2_X1 U561 ( .A1(\mem[5][14] ), .A2(n110), .ZN(n125) );
  OAI21_X1 U562 ( .B1(n811), .B2(n127), .A(n142), .ZN(n412) );
  NAND2_X1 U563 ( .A1(\mem[6][14] ), .A2(n787), .ZN(n142) );
  OAI21_X1 U564 ( .B1(n811), .B2(n146), .A(n161), .ZN(n428) );
  NAND2_X1 U565 ( .A1(\mem[7][14] ), .A2(n786), .ZN(n161) );
  OAI21_X1 U566 ( .B1(n811), .B2(n163), .A(n178), .ZN(n444) );
  NAND2_X1 U567 ( .A1(\mem[8][14] ), .A2(n785), .ZN(n178) );
  OAI21_X1 U568 ( .B1(n811), .B2(n181), .A(n196), .ZN(n460) );
  NAND2_X1 U569 ( .A1(\mem[9][14] ), .A2(n784), .ZN(n196) );
  OAI21_X1 U570 ( .B1(n811), .B2(n199), .A(n214), .ZN(n476) );
  NAND2_X1 U571 ( .A1(\mem[10][14] ), .A2(n783), .ZN(n214) );
  OAI21_X1 U572 ( .B1(n811), .B2(n216), .A(n231), .ZN(n492) );
  NAND2_X1 U573 ( .A1(\mem[11][14] ), .A2(n782), .ZN(n231) );
  OAI21_X1 U574 ( .B1(n811), .B2(n233), .A(n248), .ZN(n508) );
  NAND2_X1 U575 ( .A1(\mem[12][14] ), .A2(n781), .ZN(n248) );
  OAI21_X1 U576 ( .B1(n811), .B2(n250), .A(n265), .ZN(n524) );
  NAND2_X1 U577 ( .A1(\mem[13][14] ), .A2(n780), .ZN(n265) );
  OAI21_X1 U578 ( .B1(n811), .B2(n267), .A(n282), .ZN(n540) );
  NAND2_X1 U579 ( .A1(\mem[14][14] ), .A2(n779), .ZN(n282) );
  OAI21_X1 U580 ( .B1(n811), .B2(n285), .A(n300), .ZN(n556) );
  NAND2_X1 U581 ( .A1(\mem[15][14] ), .A2(n778), .ZN(n300) );
  OAI21_X1 U582 ( .B1(n20), .B2(n811), .A(n35), .ZN(n316) );
  NAND2_X1 U583 ( .A1(\mem[0][14] ), .A2(n20), .ZN(n35) );
  AND2_X1 U584 ( .A1(N13), .A2(wr_en), .ZN(n284) );
  MUX2_X1 U585 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n770), .Z(n1) );
  MUX2_X1 U586 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n770), .Z(n2) );
  MUX2_X1 U587 ( .A(n2), .B(n1), .S(n764), .Z(n3) );
  MUX2_X1 U588 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n770), .Z(n4) );
  MUX2_X1 U589 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n770), .Z(n5) );
  MUX2_X1 U590 ( .A(n5), .B(n4), .S(n764), .Z(n6) );
  MUX2_X1 U591 ( .A(n6), .B(n3), .S(n763), .Z(n7) );
  MUX2_X1 U592 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n770), .Z(n8) );
  MUX2_X1 U593 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n770), .Z(n9) );
  MUX2_X1 U594 ( .A(n9), .B(n8), .S(n764), .Z(n10) );
  MUX2_X1 U595 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n770), .Z(n11) );
  MUX2_X1 U596 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n770), .Z(n12) );
  MUX2_X1 U597 ( .A(n12), .B(n11), .S(n764), .Z(n13) );
  MUX2_X1 U598 ( .A(n13), .B(n10), .S(n763), .Z(n14) );
  MUX2_X1 U599 ( .A(n14), .B(n7), .S(N13), .Z(N29) );
  MUX2_X1 U600 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n777), .Z(n15) );
  MUX2_X1 U601 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(N10), .Z(n16) );
  MUX2_X1 U602 ( .A(n16), .B(n15), .S(n765), .Z(n17) );
  MUX2_X1 U603 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(N10), .Z(n18) );
  MUX2_X1 U604 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(N10), .Z(n19) );
  MUX2_X1 U605 ( .A(n19), .B(n18), .S(n765), .Z(n558) );
  MUX2_X1 U606 ( .A(n558), .B(n17), .S(n763), .Z(n559) );
  MUX2_X1 U607 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(N10), .Z(n560) );
  MUX2_X1 U608 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(N10), .Z(n561) );
  MUX2_X1 U609 ( .A(n561), .B(n560), .S(n765), .Z(n562) );
  MUX2_X1 U610 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(N10), .Z(n563) );
  MUX2_X1 U611 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n777), .Z(n564) );
  MUX2_X1 U612 ( .A(n564), .B(n563), .S(n765), .Z(n565) );
  MUX2_X1 U613 ( .A(n565), .B(n562), .S(n763), .Z(n566) );
  MUX2_X1 U614 ( .A(n566), .B(n559), .S(N13), .Z(N28) );
  MUX2_X1 U615 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n777), .Z(n567) );
  MUX2_X1 U616 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(N10), .Z(n568) );
  MUX2_X1 U617 ( .A(n568), .B(n567), .S(n765), .Z(n569) );
  MUX2_X1 U618 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(N10), .Z(n570) );
  MUX2_X1 U619 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(N10), .Z(n571) );
  MUX2_X1 U620 ( .A(n571), .B(n570), .S(n765), .Z(n572) );
  MUX2_X1 U621 ( .A(n572), .B(n569), .S(n763), .Z(n573) );
  MUX2_X1 U622 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n770), .Z(n574) );
  MUX2_X1 U623 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(N10), .Z(n575) );
  MUX2_X1 U624 ( .A(n575), .B(n574), .S(n765), .Z(n576) );
  MUX2_X1 U625 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(N10), .Z(n577) );
  MUX2_X1 U626 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(N10), .Z(n578) );
  MUX2_X1 U627 ( .A(n578), .B(n577), .S(n765), .Z(n579) );
  MUX2_X1 U628 ( .A(n579), .B(n576), .S(n763), .Z(n580) );
  MUX2_X1 U629 ( .A(n580), .B(n573), .S(N13), .Z(N27) );
  MUX2_X1 U630 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n770), .Z(n581) );
  MUX2_X1 U631 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n777), .Z(n582) );
  MUX2_X1 U632 ( .A(n582), .B(n581), .S(n765), .Z(n583) );
  MUX2_X1 U633 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n777), .Z(n584) );
  MUX2_X1 U634 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n585) );
  MUX2_X1 U635 ( .A(n585), .B(n584), .S(n765), .Z(n586) );
  MUX2_X1 U636 ( .A(n586), .B(n583), .S(n763), .Z(n587) );
  MUX2_X1 U637 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n770), .Z(n588) );
  MUX2_X1 U638 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n589) );
  MUX2_X1 U639 ( .A(n589), .B(n588), .S(n765), .Z(n590) );
  MUX2_X1 U640 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n591) );
  MUX2_X1 U641 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n592) );
  MUX2_X1 U642 ( .A(n592), .B(n591), .S(n765), .Z(n593) );
  MUX2_X1 U643 ( .A(n593), .B(n590), .S(n763), .Z(n594) );
  MUX2_X1 U644 ( .A(n594), .B(n587), .S(N13), .Z(N26) );
  MUX2_X1 U645 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n771), .Z(n595) );
  MUX2_X1 U646 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n771), .Z(n596) );
  MUX2_X1 U647 ( .A(n596), .B(n595), .S(n766), .Z(n597) );
  MUX2_X1 U648 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n771), .Z(n598) );
  MUX2_X1 U649 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n771), .Z(n599) );
  MUX2_X1 U650 ( .A(n599), .B(n598), .S(n766), .Z(n600) );
  MUX2_X1 U651 ( .A(n600), .B(n597), .S(n763), .Z(n601) );
  MUX2_X1 U652 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n771), .Z(n602) );
  MUX2_X1 U653 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n771), .Z(n603) );
  MUX2_X1 U654 ( .A(n603), .B(n602), .S(n766), .Z(n604) );
  MUX2_X1 U655 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n771), .Z(n605) );
  MUX2_X1 U656 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n771), .Z(n606) );
  MUX2_X1 U657 ( .A(n606), .B(n605), .S(n766), .Z(n607) );
  MUX2_X1 U658 ( .A(n607), .B(n604), .S(N12), .Z(n608) );
  MUX2_X1 U659 ( .A(n608), .B(n601), .S(N13), .Z(N25) );
  MUX2_X1 U660 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n771), .Z(n609) );
  MUX2_X1 U661 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n771), .Z(n610) );
  MUX2_X1 U662 ( .A(n610), .B(n609), .S(n766), .Z(n611) );
  MUX2_X1 U663 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n771), .Z(n612) );
  MUX2_X1 U664 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n771), .Z(n613) );
  MUX2_X1 U665 ( .A(n613), .B(n612), .S(n766), .Z(n614) );
  MUX2_X1 U666 ( .A(n614), .B(n611), .S(n763), .Z(n615) );
  MUX2_X1 U667 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n772), .Z(n616) );
  MUX2_X1 U668 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n772), .Z(n617) );
  MUX2_X1 U669 ( .A(n617), .B(n616), .S(n766), .Z(n618) );
  MUX2_X1 U670 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n772), .Z(n619) );
  MUX2_X1 U671 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n772), .Z(n620) );
  MUX2_X1 U672 ( .A(n620), .B(n619), .S(n766), .Z(n621) );
  MUX2_X1 U673 ( .A(n621), .B(n618), .S(n763), .Z(n622) );
  MUX2_X1 U674 ( .A(n622), .B(n615), .S(N13), .Z(N24) );
  MUX2_X1 U675 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n772), .Z(n623) );
  MUX2_X1 U676 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n772), .Z(n624) );
  MUX2_X1 U677 ( .A(n624), .B(n623), .S(n766), .Z(n625) );
  MUX2_X1 U678 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n772), .Z(n626) );
  MUX2_X1 U679 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n772), .Z(n627) );
  MUX2_X1 U680 ( .A(n627), .B(n626), .S(n766), .Z(n628) );
  MUX2_X1 U681 ( .A(n628), .B(n625), .S(n763), .Z(n629) );
  MUX2_X1 U682 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n772), .Z(n630) );
  MUX2_X1 U683 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n772), .Z(n631) );
  MUX2_X1 U684 ( .A(n631), .B(n630), .S(n766), .Z(n632) );
  MUX2_X1 U685 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n772), .Z(n633) );
  MUX2_X1 U686 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n772), .Z(n634) );
  MUX2_X1 U687 ( .A(n634), .B(n633), .S(n766), .Z(n635) );
  MUX2_X1 U688 ( .A(n635), .B(n632), .S(N12), .Z(n636) );
  MUX2_X1 U689 ( .A(n636), .B(n629), .S(N13), .Z(N23) );
  MUX2_X1 U690 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n773), .Z(n637) );
  MUX2_X1 U691 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n773), .Z(n638) );
  MUX2_X1 U692 ( .A(n638), .B(n637), .S(n767), .Z(n639) );
  MUX2_X1 U693 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n773), .Z(n640) );
  MUX2_X1 U694 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n773), .Z(n641) );
  MUX2_X1 U695 ( .A(n641), .B(n640), .S(n767), .Z(n642) );
  MUX2_X1 U696 ( .A(n642), .B(n639), .S(n763), .Z(n643) );
  MUX2_X1 U697 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n773), .Z(n644) );
  MUX2_X1 U698 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n773), .Z(n645) );
  MUX2_X1 U699 ( .A(n645), .B(n644), .S(n767), .Z(n646) );
  MUX2_X1 U700 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n773), .Z(n647) );
  MUX2_X1 U701 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n773), .Z(n648) );
  MUX2_X1 U702 ( .A(n648), .B(n647), .S(n767), .Z(n649) );
  MUX2_X1 U703 ( .A(n649), .B(n646), .S(n763), .Z(n650) );
  MUX2_X1 U704 ( .A(n650), .B(n643), .S(N13), .Z(N22) );
  MUX2_X1 U705 ( .A(\mem[14][8] ), .B(\mem[15][8] ), .S(n773), .Z(n651) );
  MUX2_X1 U706 ( .A(\mem[12][8] ), .B(\mem[13][8] ), .S(n773), .Z(n652) );
  MUX2_X1 U707 ( .A(n652), .B(n651), .S(n767), .Z(n653) );
  MUX2_X1 U708 ( .A(\mem[10][8] ), .B(\mem[11][8] ), .S(n773), .Z(n654) );
  MUX2_X1 U709 ( .A(\mem[8][8] ), .B(\mem[9][8] ), .S(n773), .Z(n655) );
  MUX2_X1 U710 ( .A(n655), .B(n654), .S(n767), .Z(n656) );
  MUX2_X1 U711 ( .A(n656), .B(n653), .S(n763), .Z(n657) );
  MUX2_X1 U712 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n777), .Z(n658) );
  MUX2_X1 U713 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n777), .Z(n659) );
  MUX2_X1 U714 ( .A(n659), .B(n658), .S(n767), .Z(n660) );
  MUX2_X1 U715 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n777), .Z(n661) );
  MUX2_X1 U716 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n777), .Z(n662) );
  MUX2_X1 U717 ( .A(n662), .B(n661), .S(n767), .Z(n663) );
  MUX2_X1 U718 ( .A(n663), .B(n660), .S(N12), .Z(n664) );
  MUX2_X1 U719 ( .A(n664), .B(n657), .S(N13), .Z(N21) );
  MUX2_X1 U720 ( .A(\mem[14][9] ), .B(\mem[15][9] ), .S(n777), .Z(n665) );
  MUX2_X1 U721 ( .A(\mem[12][9] ), .B(\mem[13][9] ), .S(n777), .Z(n666) );
  MUX2_X1 U722 ( .A(n666), .B(n665), .S(n767), .Z(n667) );
  MUX2_X1 U723 ( .A(\mem[10][9] ), .B(\mem[11][9] ), .S(n777), .Z(n668) );
  MUX2_X1 U724 ( .A(\mem[8][9] ), .B(\mem[9][9] ), .S(n777), .Z(n669) );
  MUX2_X1 U725 ( .A(n669), .B(n668), .S(n767), .Z(n670) );
  MUX2_X1 U726 ( .A(n670), .B(n667), .S(n763), .Z(n671) );
  MUX2_X1 U727 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n777), .Z(n672) );
  MUX2_X1 U728 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n777), .Z(n673) );
  MUX2_X1 U729 ( .A(n673), .B(n672), .S(n767), .Z(n674) );
  MUX2_X1 U730 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n777), .Z(n675) );
  MUX2_X1 U731 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n777), .Z(n676) );
  MUX2_X1 U732 ( .A(n676), .B(n675), .S(n767), .Z(n677) );
  MUX2_X1 U733 ( .A(n677), .B(n674), .S(n763), .Z(n678) );
  MUX2_X1 U734 ( .A(n678), .B(n671), .S(N13), .Z(N20) );
  MUX2_X1 U735 ( .A(\mem[14][10] ), .B(\mem[15][10] ), .S(n770), .Z(n679) );
  MUX2_X1 U736 ( .A(\mem[12][10] ), .B(\mem[13][10] ), .S(n770), .Z(n680) );
  MUX2_X1 U737 ( .A(n680), .B(n679), .S(n768), .Z(n681) );
  MUX2_X1 U738 ( .A(\mem[10][10] ), .B(\mem[11][10] ), .S(n770), .Z(n682) );
  MUX2_X1 U739 ( .A(\mem[8][10] ), .B(\mem[9][10] ), .S(n770), .Z(n683) );
  MUX2_X1 U740 ( .A(n683), .B(n682), .S(n768), .Z(n684) );
  MUX2_X1 U741 ( .A(n684), .B(n681), .S(n763), .Z(n685) );
  MUX2_X1 U742 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n770), .Z(n686) );
  MUX2_X1 U743 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n770), .Z(n687) );
  MUX2_X1 U744 ( .A(n687), .B(n686), .S(n768), .Z(n688) );
  MUX2_X1 U745 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n770), .Z(n689) );
  MUX2_X1 U746 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n770), .Z(n690) );
  MUX2_X1 U747 ( .A(n690), .B(n689), .S(n768), .Z(n691) );
  MUX2_X1 U748 ( .A(n691), .B(n688), .S(N12), .Z(n692) );
  MUX2_X1 U749 ( .A(n692), .B(n685), .S(N13), .Z(N19) );
  MUX2_X1 U750 ( .A(\mem[14][11] ), .B(\mem[15][11] ), .S(n770), .Z(n693) );
  MUX2_X1 U751 ( .A(\mem[12][11] ), .B(\mem[13][11] ), .S(n770), .Z(n694) );
  MUX2_X1 U752 ( .A(n694), .B(n693), .S(n768), .Z(n695) );
  MUX2_X1 U753 ( .A(\mem[10][11] ), .B(\mem[11][11] ), .S(n770), .Z(n696) );
  MUX2_X1 U754 ( .A(\mem[8][11] ), .B(\mem[9][11] ), .S(n770), .Z(n697) );
  MUX2_X1 U755 ( .A(n697), .B(n696), .S(n768), .Z(n698) );
  MUX2_X1 U756 ( .A(n698), .B(n695), .S(n763), .Z(n699) );
  MUX2_X1 U757 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n774), .Z(n700) );
  MUX2_X1 U758 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n774), .Z(n701) );
  MUX2_X1 U759 ( .A(n701), .B(n700), .S(n768), .Z(n702) );
  MUX2_X1 U760 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n774), .Z(n703) );
  MUX2_X1 U761 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n774), .Z(n704) );
  MUX2_X1 U762 ( .A(n704), .B(n703), .S(n768), .Z(n705) );
  MUX2_X1 U763 ( .A(n705), .B(n702), .S(N12), .Z(n706) );
  MUX2_X1 U764 ( .A(n706), .B(n699), .S(N13), .Z(N18) );
  MUX2_X1 U765 ( .A(\mem[14][12] ), .B(\mem[15][12] ), .S(n774), .Z(n707) );
  MUX2_X1 U766 ( .A(\mem[12][12] ), .B(\mem[13][12] ), .S(n774), .Z(n708) );
  MUX2_X1 U767 ( .A(n708), .B(n707), .S(n768), .Z(n709) );
  MUX2_X1 U768 ( .A(\mem[10][12] ), .B(\mem[11][12] ), .S(n774), .Z(n710) );
  MUX2_X1 U769 ( .A(\mem[8][12] ), .B(\mem[9][12] ), .S(n774), .Z(n711) );
  MUX2_X1 U770 ( .A(n711), .B(n710), .S(n768), .Z(n712) );
  MUX2_X1 U771 ( .A(n712), .B(n709), .S(n763), .Z(n713) );
  MUX2_X1 U772 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n774), .Z(n714) );
  MUX2_X1 U773 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n774), .Z(n715) );
  MUX2_X1 U774 ( .A(n715), .B(n714), .S(n768), .Z(n716) );
  MUX2_X1 U775 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n774), .Z(n717) );
  MUX2_X1 U776 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n774), .Z(n718) );
  MUX2_X1 U777 ( .A(n718), .B(n717), .S(n768), .Z(n719) );
  MUX2_X1 U778 ( .A(n719), .B(n716), .S(N12), .Z(n720) );
  MUX2_X1 U779 ( .A(n720), .B(n713), .S(N13), .Z(N17) );
  MUX2_X1 U780 ( .A(\mem[14][13] ), .B(\mem[15][13] ), .S(n775), .Z(n721) );
  MUX2_X1 U781 ( .A(\mem[12][13] ), .B(\mem[13][13] ), .S(n775), .Z(n722) );
  MUX2_X1 U782 ( .A(n722), .B(n721), .S(n769), .Z(n723) );
  MUX2_X1 U783 ( .A(\mem[10][13] ), .B(\mem[11][13] ), .S(n775), .Z(n724) );
  MUX2_X1 U784 ( .A(\mem[8][13] ), .B(\mem[9][13] ), .S(n775), .Z(n725) );
  MUX2_X1 U785 ( .A(n725), .B(n724), .S(n769), .Z(n726) );
  MUX2_X1 U786 ( .A(n726), .B(n723), .S(n763), .Z(n727) );
  MUX2_X1 U787 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n775), .Z(n728) );
  MUX2_X1 U788 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n775), .Z(n729) );
  MUX2_X1 U789 ( .A(n729), .B(n728), .S(n769), .Z(n730) );
  MUX2_X1 U790 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n775), .Z(n731) );
  MUX2_X1 U791 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n775), .Z(n732) );
  MUX2_X1 U792 ( .A(n732), .B(n731), .S(n769), .Z(n733) );
  MUX2_X1 U793 ( .A(n733), .B(n730), .S(N12), .Z(n734) );
  MUX2_X1 U794 ( .A(n734), .B(n727), .S(N13), .Z(N16) );
  MUX2_X1 U795 ( .A(\mem[14][14] ), .B(\mem[15][14] ), .S(n775), .Z(n735) );
  MUX2_X1 U796 ( .A(\mem[12][14] ), .B(\mem[13][14] ), .S(n775), .Z(n736) );
  MUX2_X1 U797 ( .A(n736), .B(n735), .S(n769), .Z(n737) );
  MUX2_X1 U798 ( .A(\mem[10][14] ), .B(\mem[11][14] ), .S(n775), .Z(n738) );
  MUX2_X1 U799 ( .A(\mem[8][14] ), .B(\mem[9][14] ), .S(n775), .Z(n739) );
  MUX2_X1 U800 ( .A(n739), .B(n738), .S(n769), .Z(n740) );
  MUX2_X1 U801 ( .A(n740), .B(n737), .S(n763), .Z(n741) );
  MUX2_X1 U802 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n776), .Z(n742) );
  MUX2_X1 U803 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n776), .Z(n743) );
  MUX2_X1 U804 ( .A(n743), .B(n742), .S(n769), .Z(n744) );
  MUX2_X1 U805 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n776), .Z(n745) );
  MUX2_X1 U806 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n776), .Z(n746) );
  MUX2_X1 U807 ( .A(n746), .B(n745), .S(n769), .Z(n747) );
  MUX2_X1 U808 ( .A(n747), .B(n744), .S(N12), .Z(n748) );
  MUX2_X1 U809 ( .A(n748), .B(n741), .S(N13), .Z(N15) );
  MUX2_X1 U810 ( .A(\mem[14][15] ), .B(\mem[15][15] ), .S(n776), .Z(n749) );
  MUX2_X1 U811 ( .A(\mem[12][15] ), .B(\mem[13][15] ), .S(n776), .Z(n750) );
  MUX2_X1 U812 ( .A(n750), .B(n749), .S(n769), .Z(n751) );
  MUX2_X1 U813 ( .A(\mem[10][15] ), .B(\mem[11][15] ), .S(n776), .Z(n752) );
  MUX2_X1 U814 ( .A(\mem[8][15] ), .B(\mem[9][15] ), .S(n776), .Z(n753) );
  MUX2_X1 U815 ( .A(n753), .B(n752), .S(n769), .Z(n754) );
  MUX2_X1 U816 ( .A(n754), .B(n751), .S(n763), .Z(n755) );
  MUX2_X1 U817 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n776), .Z(n756) );
  MUX2_X1 U818 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n776), .Z(n757) );
  MUX2_X1 U819 ( .A(n757), .B(n756), .S(n769), .Z(n758) );
  MUX2_X1 U820 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n776), .Z(n759) );
  MUX2_X1 U821 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n776), .Z(n760) );
  MUX2_X1 U822 ( .A(n760), .B(n759), .S(n769), .Z(n761) );
  MUX2_X1 U823 ( .A(n761), .B(n758), .S(N12), .Z(n762) );
  MUX2_X1 U824 ( .A(n762), .B(n755), .S(N13), .Z(N14) );
  CLKBUF_X1 U825 ( .A(N11), .Z(n764) );
  INV_X1 U826 ( .A(data_in[2]), .ZN(n799) );
  INV_X1 U827 ( .A(data_in[1]), .ZN(n798) );
  INV_X1 U828 ( .A(data_in[0]), .ZN(n797) );
  INV_X1 U829 ( .A(N10), .ZN(n794) );
  INV_X1 U830 ( .A(N11), .ZN(n795) );
endmodule


module datapath_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n17, n18,
         n19, n21, n23, n24, n25, n26, n27, n29, n31, n32, n33, n34, n35, n37,
         n39, n40, n41, n42, n43, n45, n47, n48, n49, n50, n51, n53, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n72, n73, n76, n78, n80, n82, n84, n85, n86, n87, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n154, n155, n156, n157,
         n158, n159;

  FA_X1 U6 ( .A(A[14]), .B(B[14]), .CI(n73), .CO(n18), .S(SUM[14]) );
  OR2_X1 U107 ( .A1(A[0]), .A2(B[0]), .ZN(n143) );
  CLKBUF_X1 U108 ( .A(n40), .Z(n144) );
  AOI21_X1 U109 ( .B1(n144), .B2(n155), .A(n37), .ZN(n145) );
  CLKBUF_X1 U110 ( .A(n59), .Z(n146) );
  CLKBUF_X1 U111 ( .A(n43), .Z(n147) );
  CLKBUF_X1 U112 ( .A(n56), .Z(n148) );
  CLKBUF_X1 U113 ( .A(n32), .Z(n149) );
  AOI21_X1 U114 ( .B1(n56), .B2(n156), .A(n53), .ZN(n150) );
  AOI21_X1 U115 ( .B1(n32), .B2(n157), .A(n29), .ZN(n151) );
  NOR2_X1 U116 ( .A1(A[3]), .A2(B[3]), .ZN(n152) );
  INV_X1 U117 ( .A(n68), .ZN(n67) );
  INV_X1 U118 ( .A(n39), .ZN(n37) );
  INV_X1 U119 ( .A(n31), .ZN(n29) );
  INV_X1 U120 ( .A(n55), .ZN(n53) );
  INV_X1 U121 ( .A(n47), .ZN(n45) );
  OAI21_X1 U122 ( .B1(n69), .B2(n72), .A(n70), .ZN(n68) );
  AOI21_X1 U123 ( .B1(n60), .B2(n68), .A(n61), .ZN(n59) );
  NAND2_X1 U124 ( .A1(n82), .A2(n50), .ZN(n9) );
  INV_X1 U125 ( .A(n49), .ZN(n82) );
  XOR2_X1 U126 ( .A(n14), .B(n72), .Z(SUM[1]) );
  NAND2_X1 U127 ( .A1(n87), .A2(n70), .ZN(n14) );
  NAND2_X1 U128 ( .A1(n156), .A2(n55), .ZN(n10) );
  XNOR2_X1 U129 ( .A(n64), .B(n12), .ZN(SUM[3]) );
  NAND2_X1 U130 ( .A1(n85), .A2(n63), .ZN(n12) );
  OAI21_X1 U131 ( .B1(n67), .B2(n65), .A(n66), .ZN(n64) );
  AND2_X1 U132 ( .A1(n143), .A2(n72), .ZN(SUM[0]) );
  NAND2_X1 U133 ( .A1(n84), .A2(n58), .ZN(n11) );
  INV_X1 U134 ( .A(n57), .ZN(n84) );
  NAND2_X1 U135 ( .A1(n76), .A2(n26), .ZN(n3) );
  INV_X1 U136 ( .A(n25), .ZN(n76) );
  NAND2_X1 U137 ( .A1(n78), .A2(n34), .ZN(n5) );
  INV_X1 U138 ( .A(n33), .ZN(n78) );
  NAND2_X1 U139 ( .A1(n80), .A2(n42), .ZN(n7) );
  INV_X1 U140 ( .A(n41), .ZN(n80) );
  XOR2_X1 U141 ( .A(n67), .B(n13), .Z(SUM[2]) );
  NAND2_X1 U142 ( .A1(n86), .A2(n66), .ZN(n13) );
  INV_X1 U143 ( .A(n65), .ZN(n86) );
  NAND2_X1 U144 ( .A1(n158), .A2(n23), .ZN(n2) );
  NAND2_X1 U145 ( .A1(n157), .A2(n31), .ZN(n4) );
  NAND2_X1 U146 ( .A1(n155), .A2(n39), .ZN(n6) );
  NAND2_X1 U147 ( .A1(n154), .A2(n47), .ZN(n8) );
  NOR2_X1 U148 ( .A1(A[2]), .A2(B[2]), .ZN(n65) );
  NAND2_X1 U149 ( .A1(A[2]), .A2(B[2]), .ZN(n66) );
  NAND2_X1 U150 ( .A1(A[0]), .A2(B[0]), .ZN(n72) );
  NOR2_X1 U151 ( .A1(A[1]), .A2(B[1]), .ZN(n69) );
  INV_X1 U152 ( .A(n23), .ZN(n21) );
  NOR2_X1 U153 ( .A1(A[8]), .A2(B[8]), .ZN(n41) );
  NOR2_X1 U154 ( .A1(A[6]), .A2(B[6]), .ZN(n49) );
  NOR2_X1 U155 ( .A1(A[4]), .A2(B[4]), .ZN(n57) );
  NOR2_X1 U156 ( .A1(A[12]), .A2(B[12]), .ZN(n25) );
  NOR2_X1 U157 ( .A1(A[10]), .A2(B[10]), .ZN(n33) );
  NAND2_X1 U158 ( .A1(A[7]), .A2(B[7]), .ZN(n47) );
  NAND2_X1 U159 ( .A1(A[9]), .A2(B[9]), .ZN(n39) );
  NAND2_X1 U160 ( .A1(A[5]), .A2(B[5]), .ZN(n55) );
  NAND2_X1 U161 ( .A1(A[11]), .A2(B[11]), .ZN(n31) );
  NAND2_X1 U162 ( .A1(A[13]), .A2(B[13]), .ZN(n23) );
  NAND2_X1 U163 ( .A1(A[8]), .A2(B[8]), .ZN(n42) );
  NAND2_X1 U164 ( .A1(A[6]), .A2(B[6]), .ZN(n50) );
  NAND2_X1 U165 ( .A1(A[4]), .A2(B[4]), .ZN(n58) );
  NAND2_X1 U166 ( .A1(A[12]), .A2(B[12]), .ZN(n26) );
  NAND2_X1 U167 ( .A1(A[10]), .A2(B[10]), .ZN(n34) );
  OR2_X1 U168 ( .A1(A[7]), .A2(B[7]), .ZN(n154) );
  OR2_X1 U169 ( .A1(A[9]), .A2(B[9]), .ZN(n155) );
  OR2_X1 U170 ( .A1(A[5]), .A2(B[5]), .ZN(n156) );
  OR2_X1 U171 ( .A1(A[11]), .A2(B[11]), .ZN(n157) );
  OR2_X1 U172 ( .A1(A[13]), .A2(B[13]), .ZN(n158) );
  NAND2_X1 U173 ( .A1(A[3]), .A2(B[3]), .ZN(n63) );
  OR2_X1 U174 ( .A1(A[15]), .A2(B[15]), .ZN(n159) );
  XNOR2_X1 U175 ( .A(n18), .B(n1), .ZN(SUM[15]) );
  NAND2_X1 U176 ( .A1(n159), .A2(n17), .ZN(n1) );
  NAND2_X1 U177 ( .A1(A[15]), .A2(B[15]), .ZN(n17) );
  INV_X1 U178 ( .A(n152), .ZN(n85) );
  OAI21_X1 U179 ( .B1(n43), .B2(n41), .A(n42), .ZN(n40) );
  AOI21_X1 U180 ( .B1(n48), .B2(n154), .A(n45), .ZN(n43) );
  XNOR2_X1 U181 ( .A(n48), .B(n8), .ZN(SUM[7]) );
  INV_X1 U182 ( .A(n69), .ZN(n87) );
  OAI21_X1 U183 ( .B1(n150), .B2(n49), .A(n50), .ZN(n48) );
  XNOR2_X1 U184 ( .A(n149), .B(n4), .ZN(SUM[11]) );
  AOI21_X1 U185 ( .B1(n149), .B2(n157), .A(n29), .ZN(n27) );
  OAI21_X1 U186 ( .B1(n35), .B2(n33), .A(n34), .ZN(n32) );
  XNOR2_X1 U187 ( .A(n144), .B(n6), .ZN(SUM[9]) );
  XOR2_X1 U188 ( .A(n145), .B(n5), .Z(SUM[10]) );
  XOR2_X1 U189 ( .A(n51), .B(n9), .Z(SUM[6]) );
  AOI21_X1 U190 ( .B1(n40), .B2(n155), .A(n37), .ZN(n35) );
  AOI21_X1 U191 ( .B1(n148), .B2(n156), .A(n53), .ZN(n51) );
  XOR2_X1 U192 ( .A(n27), .B(n3), .Z(SUM[12]) );
  XOR2_X1 U193 ( .A(n147), .B(n7), .Z(SUM[8]) );
  XNOR2_X1 U194 ( .A(n148), .B(n10), .ZN(SUM[5]) );
  NAND2_X1 U195 ( .A1(A[1]), .A2(B[1]), .ZN(n70) );
  OAI21_X1 U196 ( .B1(n59), .B2(n57), .A(n58), .ZN(n56) );
  XOR2_X1 U197 ( .A(n146), .B(n11), .Z(SUM[4]) );
  XNOR2_X1 U198 ( .A(n24), .B(n2), .ZN(SUM[13]) );
  INV_X1 U199 ( .A(n19), .ZN(n73) );
  OAI21_X1 U200 ( .B1(n62), .B2(n66), .A(n63), .ZN(n61) );
  NOR2_X1 U201 ( .A1(n65), .A2(n152), .ZN(n60) );
  OAI21_X1 U202 ( .B1(n151), .B2(n25), .A(n26), .ZN(n24) );
  AOI21_X1 U203 ( .B1(n24), .B2(n158), .A(n21), .ZN(n19) );
  NOR2_X1 U204 ( .A1(A[3]), .A2(B[3]), .ZN(n62) );
endmodule


module datapath_DW_mult_tc_1 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n16,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n44, n45, n46, n47, n50,
         n56, n57, n58, n62, n63, n64, n65, n66, n67, n68, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n83, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n95, n97, n100, n101, n102, n103, n105, n108,
         n109, n111, n112, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n160, n161, n163, n164, n166, n167, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n258, n259, n261, n262, n263, n264, n265, n266, n267,
         n268, n276, n306, n307, n308, n309, n310, n311, n312, n313, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398;
  assign n167 = a[0];
  assign n248 = b[0];
  assign n265 = a[7];
  assign n266 = a[5];
  assign n267 = a[3];
  assign n268 = a[1];

  FA_X1 U131 ( .A(n174), .B(n181), .CI(n121), .CO(n117), .S(n118) );
  FA_X1 U134 ( .A(n129), .B(n176), .CI(n126), .CO(n123), .S(n124) );
  FA_X1 U135 ( .A(n335), .B(n182), .CI(n189), .CO(n125), .S(n126) );
  FA_X1 U136 ( .A(n135), .B(n137), .CI(n130), .CO(n127), .S(n128) );
  FA_X1 U137 ( .A(n177), .B(n183), .CI(n132), .CO(n129), .S(n130) );
  FA_X1 U140 ( .A(n197), .B(n184), .CI(n143), .CO(n135), .S(n136) );
  FA_X1 U144 ( .A(n185), .B(n198), .CI(n191), .CO(n141), .S(n142) );
  HA_X1 U145 ( .A(n179), .B(n169), .CO(n143), .S(n144) );
  FA_X1 U147 ( .A(n199), .B(n180), .CI(n192), .CO(n147), .S(n148) );
  HA_X1 U149 ( .A(n187), .B(n170), .CO(n151), .S(n152) );
  FA_X1 U150 ( .A(n201), .B(n188), .CI(n194), .CO(n153), .S(n154) );
  HA_X1 U151 ( .A(n195), .B(n202), .CO(n155), .S(n156) );
  BUF_X1 U271 ( .A(n266), .Z(n388) );
  AND2_X1 U272 ( .A1(n204), .A2(n172), .ZN(n326) );
  BUF_X1 U273 ( .A(n268), .Z(n383) );
  AND2_X1 U274 ( .A1(n120), .A2(n123), .ZN(n313) );
  INV_X1 U275 ( .A(n326), .ZN(n100) );
  OR2_X1 U276 ( .A1(n204), .A2(n172), .ZN(n306) );
  INV_X1 U277 ( .A(n276), .ZN(n307) );
  NAND2_X1 U278 ( .A1(n259), .A2(n251), .ZN(n308) );
  BUF_X1 U279 ( .A(n265), .Z(n309) );
  BUF_X1 U280 ( .A(n265), .Z(n310) );
  CLKBUF_X1 U281 ( .A(n41), .Z(n311) );
  OR2_X1 U282 ( .A1(n123), .A2(n120), .ZN(n312) );
  AND2_X1 U283 ( .A1(n340), .A2(n20), .ZN(product[15]) );
  CLKBUF_X1 U284 ( .A(n141), .Z(n315) );
  NAND2_X1 U285 ( .A1(n338), .A2(n339), .ZN(n316) );
  CLKBUF_X1 U286 ( .A(n267), .Z(n317) );
  NOR2_X1 U287 ( .A1(n41), .A2(n34), .ZN(n318) );
  OAI21_X1 U288 ( .B1(n354), .B2(n81), .A(n80), .ZN(n319) );
  OAI21_X1 U289 ( .B1(n87), .B2(n89), .A(n88), .ZN(n320) );
  NOR2_X2 U290 ( .A1(n154), .A2(n155), .ZN(n87) );
  AOI21_X1 U291 ( .B1(n380), .B2(n320), .A(n83), .ZN(n321) );
  OAI21_X1 U292 ( .B1(n72), .B2(n76), .A(n73), .ZN(n322) );
  INV_X1 U293 ( .A(n313), .ZN(n323) );
  XNOR2_X1 U294 ( .A(n148), .B(n324), .ZN(n146) );
  XNOR2_X1 U295 ( .A(n151), .B(n186), .ZN(n324) );
  XNOR2_X1 U296 ( .A(n325), .B(n142), .ZN(n140) );
  XNOR2_X1 U297 ( .A(n147), .B(n144), .ZN(n325) );
  BUF_X1 U298 ( .A(n136), .Z(n329) );
  BUF_X1 U299 ( .A(n152), .Z(n327) );
  NAND2_X1 U300 ( .A1(n128), .A2(n133), .ZN(n328) );
  CLKBUF_X3 U301 ( .A(n268), .Z(n349) );
  INV_X1 U302 ( .A(n39), .ZN(n330) );
  NAND2_X1 U303 ( .A1(n64), .A2(n331), .ZN(n37) );
  NOR2_X1 U304 ( .A1(n386), .A2(n330), .ZN(n331) );
  CLKBUF_X1 U305 ( .A(n267), .Z(n332) );
  CLKBUF_X1 U306 ( .A(n266), .Z(n333) );
  XNOR2_X2 U307 ( .A(n383), .B(a[2]), .ZN(n375) );
  OAI21_X1 U308 ( .B1(n354), .B2(n81), .A(n80), .ZN(n370) );
  INV_X1 U309 ( .A(n65), .ZN(n334) );
  OAI22_X1 U310 ( .A1(n395), .A2(n224), .B1(n375), .B2(n223), .ZN(n335) );
  NAND2_X1 U311 ( .A1(n267), .A2(n337), .ZN(n338) );
  NAND2_X1 U312 ( .A1(n336), .A2(a[2]), .ZN(n339) );
  NAND2_X1 U313 ( .A1(n338), .A2(n339), .ZN(n251) );
  INV_X1 U314 ( .A(n267), .ZN(n336) );
  INV_X1 U315 ( .A(a[2]), .ZN(n337) );
  OAI22_X1 U316 ( .A1(n308), .A2(n224), .B1(n375), .B2(n223), .ZN(n131) );
  OR2_X1 U317 ( .A1(n358), .A2(n19), .ZN(n340) );
  CLKBUF_X1 U318 ( .A(n267), .Z(n341) );
  CLKBUF_X1 U319 ( .A(n75), .Z(n342) );
  CLKBUF_X1 U320 ( .A(n321), .Z(n343) );
  NAND2_X1 U321 ( .A1(n142), .A2(n147), .ZN(n344) );
  NAND2_X1 U322 ( .A1(n142), .A2(n144), .ZN(n345) );
  NAND2_X1 U323 ( .A1(n147), .A2(n144), .ZN(n346) );
  NAND3_X1 U324 ( .A1(n344), .A2(n345), .A3(n346), .ZN(n139) );
  NOR2_X1 U325 ( .A1(n66), .A2(n386), .ZN(n347) );
  NOR2_X1 U326 ( .A1(n124), .A2(n127), .ZN(n348) );
  NOR2_X1 U327 ( .A1(n66), .A2(n386), .ZN(n3) );
  NOR2_X1 U328 ( .A1(n124), .A2(n127), .ZN(n386) );
  XNOR2_X2 U329 ( .A(n266), .B(a[6]), .ZN(n372) );
  NAND2_X1 U330 ( .A1(n148), .A2(n151), .ZN(n350) );
  NAND2_X1 U331 ( .A1(n148), .A2(n186), .ZN(n351) );
  NAND2_X1 U332 ( .A1(n151), .A2(n186), .ZN(n352) );
  NAND3_X1 U333 ( .A1(n350), .A2(n351), .A3(n352), .ZN(n145) );
  CLKBUF_X1 U334 ( .A(n2), .Z(n353) );
  NOR2_X1 U335 ( .A1(n146), .A2(n149), .ZN(n354) );
  NOR2_X1 U336 ( .A1(n146), .A2(n149), .ZN(n79) );
  XNOR2_X1 U337 ( .A(n355), .B(n136), .ZN(n134) );
  XNOR2_X1 U338 ( .A(n141), .B(n138), .ZN(n355) );
  BUF_X1 U339 ( .A(n312), .Z(n356) );
  CLKBUF_X1 U340 ( .A(n76), .Z(n357) );
  AOI21_X1 U341 ( .B1(n370), .B2(n70), .A(n322), .ZN(n358) );
  AOI21_X1 U342 ( .B1(n70), .B2(n319), .A(n322), .ZN(n376) );
  AOI21_X1 U343 ( .B1(n32), .B2(n313), .A(n33), .ZN(n359) );
  NAND2_X1 U344 ( .A1(n258), .A2(n250), .ZN(n360) );
  NAND2_X1 U345 ( .A1(n250), .A2(n258), .ZN(n254) );
  XOR2_X1 U346 ( .A(n122), .B(n175), .Z(n361) );
  XOR2_X1 U347 ( .A(n125), .B(n361), .Z(n120) );
  NAND2_X1 U348 ( .A1(n125), .A2(n122), .ZN(n362) );
  NAND2_X1 U349 ( .A1(n125), .A2(n175), .ZN(n363) );
  NAND2_X1 U350 ( .A1(n122), .A2(n175), .ZN(n364) );
  NAND3_X1 U351 ( .A1(n362), .A2(n363), .A3(n364), .ZN(n119) );
  NAND2_X1 U352 ( .A1(n329), .A2(n315), .ZN(n365) );
  NAND2_X1 U353 ( .A1(n329), .A2(n138), .ZN(n366) );
  NAND2_X1 U354 ( .A1(n315), .A2(n138), .ZN(n367) );
  NAND3_X1 U355 ( .A1(n365), .A2(n366), .A3(n367), .ZN(n133) );
  BUF_X2 U356 ( .A(n384), .Z(n368) );
  BUF_X1 U357 ( .A(n384), .Z(n369) );
  XNOR2_X1 U358 ( .A(n267), .B(a[4]), .ZN(n384) );
  NAND2_X1 U359 ( .A1(n249), .A2(n387), .ZN(n371) );
  BUF_X1 U360 ( .A(n256), .Z(n381) );
  OAI21_X1 U361 ( .B1(n328), .B2(n348), .A(n62), .ZN(n373) );
  OAI21_X1 U362 ( .B1(n67), .B2(n348), .A(n62), .ZN(n2) );
  XNOR2_X1 U363 ( .A(n349), .B(a[2]), .ZN(n374) );
  XNOR2_X1 U364 ( .A(n383), .B(a[2]), .ZN(n259) );
  XNOR2_X1 U365 ( .A(n68), .B(n9), .ZN(product[9]) );
  XOR2_X1 U366 ( .A(n265), .B(a[6]), .Z(n249) );
  NOR2_X1 U367 ( .A1(n134), .A2(n139), .ZN(n377) );
  AOI21_X1 U368 ( .B1(n70), .B2(n78), .A(n71), .ZN(n1) );
  INV_X1 U369 ( .A(n30), .ZN(n28) );
  INV_X1 U370 ( .A(n66), .ZN(n64) );
  OAI21_X1 U371 ( .B1(n359), .B2(n23), .A(n24), .ZN(n22) );
  NOR2_X1 U372 ( .A1(n30), .A2(n23), .ZN(n21) );
  INV_X1 U373 ( .A(n23), .ZN(n101) );
  INV_X1 U374 ( .A(n34), .ZN(n102) );
  INV_X1 U375 ( .A(n386), .ZN(n105) );
  INV_X1 U376 ( .A(n97), .ZN(n95) );
  INV_X1 U377 ( .A(n115), .ZN(n116) );
  NOR2_X1 U378 ( .A1(n173), .A2(n115), .ZN(n23) );
  NOR2_X1 U379 ( .A1(n140), .A2(n145), .ZN(n75) );
  NAND2_X1 U380 ( .A1(n112), .A2(n92), .ZN(n15) );
  INV_X1 U381 ( .A(n91), .ZN(n112) );
  NAND2_X1 U382 ( .A1(n111), .A2(n88), .ZN(n14) );
  NAND2_X1 U383 ( .A1(n173), .A2(n115), .ZN(n24) );
  NOR2_X1 U384 ( .A1(n117), .A2(n116), .ZN(n34) );
  NAND2_X1 U385 ( .A1(n119), .A2(n118), .ZN(n44) );
  NAND2_X1 U386 ( .A1(n117), .A2(n116), .ZN(n35) );
  NAND2_X1 U387 ( .A1(n109), .A2(n80), .ZN(n12) );
  INV_X1 U388 ( .A(n354), .ZN(n109) );
  XOR2_X1 U389 ( .A(n77), .B(n11), .Z(product[7]) );
  INV_X1 U390 ( .A(n342), .ZN(n108) );
  NAND2_X1 U391 ( .A1(n101), .A2(n24), .ZN(n4) );
  NAND2_X1 U392 ( .A1(n102), .A2(n35), .ZN(n5) );
  XNOR2_X1 U393 ( .A(n56), .B(n7), .ZN(product[11]) );
  XNOR2_X1 U394 ( .A(n45), .B(n6), .ZN(product[12]) );
  XNOR2_X1 U395 ( .A(n74), .B(n10), .ZN(product[8]) );
  XNOR2_X1 U396 ( .A(n16), .B(n326), .ZN(product[2]) );
  NAND2_X1 U397 ( .A1(n379), .A2(n97), .ZN(n16) );
  AND2_X1 U398 ( .A1(n306), .A2(n100), .ZN(product[1]) );
  BUF_X1 U399 ( .A(n253), .Z(n393) );
  INV_X1 U400 ( .A(n157), .ZN(n173) );
  OR2_X1 U401 ( .A1(n203), .A2(n196), .ZN(n379) );
  OR2_X1 U402 ( .A1(n150), .A2(n153), .ZN(n380) );
  NAND2_X1 U403 ( .A1(n154), .A2(n155), .ZN(n88) );
  OR2_X1 U404 ( .A1(n248), .A2(n262), .ZN(n222) );
  OR2_X1 U405 ( .A1(n248), .A2(n264), .ZN(n240) );
  XNOR2_X1 U406 ( .A(n267), .B(a[4]), .ZN(n258) );
  AND2_X1 U407 ( .A1(n248), .A2(n158), .ZN(n180) );
  AND2_X1 U408 ( .A1(n248), .A2(n164), .ZN(n196) );
  AND2_X1 U409 ( .A1(n248), .A2(n307), .ZN(product[0]) );
  OR2_X1 U410 ( .A1(n248), .A2(n261), .ZN(n213) );
  NAND2_X1 U411 ( .A1(n64), .A2(n334), .ZN(n9) );
  INV_X1 U412 ( .A(n328), .ZN(n65) );
  AOI21_X1 U413 ( .B1(n313), .B2(n318), .A(n33), .ZN(n31) );
  BUF_X2 U414 ( .A(n256), .Z(n382) );
  NAND2_X1 U415 ( .A1(n252), .A2(n276), .ZN(n256) );
  NAND2_X1 U416 ( .A1(n124), .A2(n127), .ZN(n62) );
  XNOR2_X1 U417 ( .A(n36), .B(n5), .ZN(product[13]) );
  XNOR2_X1 U418 ( .A(n13), .B(n320), .ZN(product[5]) );
  INV_X1 U419 ( .A(n87), .ZN(n111) );
  OAI21_X1 U420 ( .B1(n87), .B2(n89), .A(n88), .ZN(n86) );
  XNOR2_X1 U421 ( .A(n152), .B(n385), .ZN(n150) );
  XNOR2_X1 U422 ( .A(n193), .B(n200), .ZN(n385) );
  XNOR2_X1 U423 ( .A(n266), .B(a[6]), .ZN(n387) );
  INV_X1 U424 ( .A(n166), .ZN(n197) );
  NAND2_X1 U425 ( .A1(n396), .A2(n73), .ZN(n10) );
  NAND2_X1 U426 ( .A1(n103), .A2(n44), .ZN(n6) );
  OAI21_X1 U427 ( .B1(n44), .B2(n34), .A(n35), .ZN(n33) );
  NAND2_X1 U428 ( .A1(n134), .A2(n139), .ZN(n73) );
  OAI21_X1 U429 ( .B1(n77), .B2(n342), .A(n357), .ZN(n74) );
  NAND2_X1 U430 ( .A1(n108), .A2(n357), .ZN(n11) );
  XNOR2_X1 U431 ( .A(n310), .B(b[4]), .ZN(n208) );
  XNOR2_X1 U432 ( .A(n310), .B(b[5]), .ZN(n207) );
  XNOR2_X1 U433 ( .A(n310), .B(b[6]), .ZN(n206) );
  XNOR2_X1 U434 ( .A(n310), .B(b[2]), .ZN(n210) );
  XNOR2_X1 U435 ( .A(n309), .B(b[7]), .ZN(n205) );
  XNOR2_X1 U436 ( .A(n310), .B(b[3]), .ZN(n209) );
  XNOR2_X1 U437 ( .A(n309), .B(n248), .ZN(n212) );
  XNOR2_X1 U438 ( .A(n309), .B(b[1]), .ZN(n211) );
  INV_X1 U439 ( .A(n265), .ZN(n261) );
  NOR2_X1 U440 ( .A1(n156), .A2(n171), .ZN(n91) );
  XNOR2_X1 U441 ( .A(n25), .B(n4), .ZN(product[14]) );
  XOR2_X1 U442 ( .A(n15), .B(n93), .Z(product[3]) );
  NAND2_X1 U443 ( .A1(n203), .A2(n196), .ZN(n97) );
  NAND2_X1 U444 ( .A1(n140), .A2(n145), .ZN(n76) );
  AOI21_X1 U445 ( .B1(n353), .B2(n21), .A(n22), .ZN(n20) );
  INV_X1 U446 ( .A(n373), .ZN(n58) );
  NOR2_X1 U447 ( .A1(n133), .A2(n128), .ZN(n66) );
  NAND2_X1 U448 ( .A1(n128), .A2(n133), .ZN(n67) );
  XOR2_X1 U449 ( .A(n14), .B(n89), .Z(product[4]) );
  NAND2_X1 U450 ( .A1(n327), .A2(n193), .ZN(n389) );
  NAND2_X1 U451 ( .A1(n327), .A2(n200), .ZN(n390) );
  NAND2_X1 U452 ( .A1(n193), .A2(n200), .ZN(n391) );
  NAND3_X1 U453 ( .A1(n389), .A2(n390), .A3(n391), .ZN(n149) );
  NAND2_X1 U454 ( .A1(n146), .A2(n149), .ZN(n80) );
  XNOR2_X1 U455 ( .A(n63), .B(n392), .ZN(product[10]) );
  AND2_X1 U456 ( .A1(n105), .A2(n62), .ZN(n392) );
  OR2_X1 U457 ( .A1(n190), .A2(n178), .ZN(n137) );
  XNOR2_X1 U458 ( .A(n190), .B(n178), .ZN(n138) );
  INV_X1 U459 ( .A(n163), .ZN(n189) );
  INV_X1 U460 ( .A(n121), .ZN(n122) );
  AND2_X1 U461 ( .A1(n248), .A2(n161), .ZN(n188) );
  INV_X1 U462 ( .A(n160), .ZN(n181) );
  OR2_X1 U463 ( .A1(n248), .A2(n263), .ZN(n231) );
  NAND2_X1 U464 ( .A1(n387), .A2(n249), .ZN(n253) );
  OAI22_X1 U465 ( .A1(n382), .A2(n235), .B1(n234), .B2(n276), .ZN(n200) );
  OAI22_X1 U466 ( .A1(n382), .A2(n236), .B1(n235), .B2(n276), .ZN(n201) );
  OAI22_X1 U467 ( .A1(n381), .A2(n234), .B1(n233), .B2(n276), .ZN(n199) );
  OAI22_X1 U468 ( .A1(n381), .A2(n233), .B1(n232), .B2(n276), .ZN(n198) );
  OAI22_X1 U469 ( .A1(n381), .A2(n239), .B1(n238), .B2(n276), .ZN(n204) );
  OAI22_X1 U470 ( .A1(n382), .A2(n237), .B1(n236), .B2(n276), .ZN(n202) );
  OAI22_X1 U471 ( .A1(n232), .A2(n382), .B1(n232), .B2(n276), .ZN(n166) );
  OAI22_X1 U472 ( .A1(n381), .A2(n238), .B1(n237), .B2(n276), .ZN(n203) );
  NAND2_X1 U473 ( .A1(n316), .A2(n374), .ZN(n394) );
  NAND2_X1 U474 ( .A1(n259), .A2(n251), .ZN(n395) );
  NAND2_X1 U475 ( .A1(n316), .A2(n259), .ZN(n255) );
  INV_X1 U476 ( .A(n90), .ZN(n89) );
  OR2_X1 U477 ( .A1(n134), .A2(n139), .ZN(n396) );
  NAND2_X1 U478 ( .A1(n380), .A2(n85), .ZN(n13) );
  INV_X1 U479 ( .A(n85), .ZN(n83) );
  INV_X1 U480 ( .A(n31), .ZN(n29) );
  NOR2_X1 U481 ( .A1(n254), .A2(n221), .ZN(n397) );
  NOR2_X1 U482 ( .A1(n368), .A2(n220), .ZN(n398) );
  OR2_X1 U483 ( .A1(n397), .A2(n398), .ZN(n187) );
  AOI21_X1 U484 ( .B1(n379), .B2(n326), .A(n95), .ZN(n93) );
  OAI21_X1 U485 ( .B1(n91), .B2(n93), .A(n92), .ZN(n90) );
  OAI22_X1 U486 ( .A1(n382), .A2(n264), .B1(n240), .B2(n276), .ZN(n172) );
  OAI21_X1 U487 ( .B1(n377), .B2(n76), .A(n73), .ZN(n71) );
  NOR2_X1 U488 ( .A1(n72), .A2(n75), .ZN(n70) );
  NOR2_X1 U489 ( .A1(n134), .A2(n139), .ZN(n72) );
  INV_X1 U490 ( .A(n131), .ZN(n132) );
  AOI21_X1 U491 ( .B1(n373), .B2(n39), .A(n40), .ZN(n38) );
  AOI21_X1 U492 ( .B1(n2), .B2(n28), .A(n29), .ZN(n27) );
  NAND2_X1 U493 ( .A1(n3), .A2(n28), .ZN(n26) );
  INV_X1 U494 ( .A(n347), .ZN(n57) );
  NAND2_X1 U495 ( .A1(n347), .A2(n21), .ZN(n19) );
  NAND2_X1 U496 ( .A1(n150), .A2(n153), .ZN(n85) );
  INV_X1 U497 ( .A(n319), .ZN(n77) );
  NAND2_X1 U498 ( .A1(n156), .A2(n171), .ZN(n92) );
  INV_X1 U499 ( .A(n311), .ZN(n103) );
  OAI21_X1 U500 ( .B1(n323), .B2(n311), .A(n44), .ZN(n40) );
  NOR2_X1 U501 ( .A1(n50), .A2(n41), .ZN(n39) );
  NOR2_X1 U502 ( .A1(n41), .A2(n34), .ZN(n32) );
  NOR2_X2 U503 ( .A1(n119), .A2(n118), .ZN(n41) );
  OAI22_X1 U504 ( .A1(n395), .A2(n263), .B1(n231), .B2(n375), .ZN(n171) );
  OAI22_X1 U505 ( .A1(n394), .A2(n228), .B1(n375), .B2(n227), .ZN(n193) );
  OAI22_X1 U506 ( .A1(n394), .A2(n229), .B1(n375), .B2(n228), .ZN(n194) );
  OAI22_X1 U507 ( .A1(n308), .A2(n225), .B1(n375), .B2(n224), .ZN(n190) );
  OAI22_X1 U508 ( .A1(n394), .A2(n227), .B1(n375), .B2(n226), .ZN(n192) );
  OAI22_X1 U509 ( .A1(n395), .A2(n226), .B1(n375), .B2(n225), .ZN(n191) );
  XNOR2_X1 U510 ( .A(n349), .B(b[4]), .ZN(n235) );
  XNOR2_X1 U511 ( .A(n349), .B(b[5]), .ZN(n234) );
  OAI22_X1 U512 ( .A1(n255), .A2(n230), .B1(n375), .B2(n229), .ZN(n195) );
  INV_X1 U513 ( .A(n374), .ZN(n164) );
  XNOR2_X1 U514 ( .A(n349), .B(b[6]), .ZN(n233) );
  OAI22_X1 U515 ( .A1(n255), .A2(n223), .B1(n223), .B2(n375), .ZN(n163) );
  XNOR2_X1 U516 ( .A(n349), .B(b[3]), .ZN(n236) );
  XNOR2_X1 U517 ( .A(n349), .B(b[2]), .ZN(n237) );
  XNOR2_X1 U518 ( .A(n349), .B(n248), .ZN(n239) );
  XNOR2_X1 U519 ( .A(n349), .B(b[1]), .ZN(n238) );
  XNOR2_X1 U520 ( .A(n349), .B(b[7]), .ZN(n232) );
  INV_X1 U521 ( .A(n349), .ZN(n264) );
  XOR2_X1 U522 ( .A(n268), .B(n167), .Z(n252) );
  AOI21_X1 U523 ( .B1(n2), .B2(n356), .A(n313), .ZN(n47) );
  NAND2_X1 U524 ( .A1(n3), .A2(n356), .ZN(n46) );
  NAND2_X1 U525 ( .A1(n356), .A2(n323), .ZN(n7) );
  NAND2_X1 U526 ( .A1(n312), .A2(n32), .ZN(n30) );
  NOR2_X1 U527 ( .A1(n123), .A2(n120), .ZN(n50) );
  XOR2_X1 U528 ( .A(n12), .B(n343), .Z(product[6]) );
  OAI21_X1 U529 ( .B1(n321), .B2(n79), .A(n80), .ZN(n78) );
  OAI22_X1 U530 ( .A1(n360), .A2(n220), .B1(n368), .B2(n219), .ZN(n186) );
  OAI22_X1 U531 ( .A1(n360), .A2(n215), .B1(n368), .B2(n214), .ZN(n121) );
  OAI22_X1 U532 ( .A1(n360), .A2(n217), .B1(n369), .B2(n216), .ZN(n183) );
  INV_X1 U533 ( .A(n368), .ZN(n161) );
  OAI22_X1 U534 ( .A1(n254), .A2(n219), .B1(n368), .B2(n218), .ZN(n185) );
  OAI22_X1 U535 ( .A1(n218), .A2(n360), .B1(n369), .B2(n217), .ZN(n184) );
  OAI22_X1 U536 ( .A1(n214), .A2(n360), .B1(n214), .B2(n369), .ZN(n160) );
  OAI22_X1 U537 ( .A1(n254), .A2(n216), .B1(n368), .B2(n215), .ZN(n182) );
  INV_X1 U538 ( .A(n332), .ZN(n263) );
  OAI22_X1 U539 ( .A1(n360), .A2(n262), .B1(n222), .B2(n369), .ZN(n170) );
  XNOR2_X1 U540 ( .A(n341), .B(b[3]), .ZN(n227) );
  XNOR2_X1 U541 ( .A(n332), .B(b[4]), .ZN(n226) );
  XNOR2_X1 U542 ( .A(n332), .B(b[2]), .ZN(n228) );
  XNOR2_X1 U543 ( .A(n341), .B(b[5]), .ZN(n225) );
  XNOR2_X1 U544 ( .A(n317), .B(b[6]), .ZN(n224) );
  XNOR2_X1 U545 ( .A(n317), .B(n248), .ZN(n230) );
  XNOR2_X1 U546 ( .A(n341), .B(b[1]), .ZN(n229) );
  XNOR2_X1 U547 ( .A(n267), .B(b[7]), .ZN(n223) );
  OAI22_X1 U548 ( .A1(n205), .A2(n393), .B1(n205), .B2(n372), .ZN(n157) );
  OAI22_X1 U549 ( .A1(n393), .A2(n209), .B1(n372), .B2(n208), .ZN(n176) );
  OAI22_X1 U550 ( .A1(n393), .A2(n206), .B1(n372), .B2(n205), .ZN(n115) );
  OAI22_X1 U551 ( .A1(n393), .A2(n208), .B1(n372), .B2(n207), .ZN(n175) );
  OAI22_X1 U552 ( .A1(n393), .A2(n207), .B1(n372), .B2(n206), .ZN(n174) );
  OAI22_X1 U553 ( .A1(n371), .A2(n210), .B1(n372), .B2(n209), .ZN(n177) );
  INV_X1 U554 ( .A(n372), .ZN(n158) );
  OAI22_X1 U555 ( .A1(n393), .A2(n211), .B1(n372), .B2(n210), .ZN(n178) );
  OAI22_X1 U556 ( .A1(n371), .A2(n261), .B1(n213), .B2(n372), .ZN(n169) );
  OAI22_X1 U557 ( .A1(n253), .A2(n212), .B1(n372), .B2(n211), .ZN(n179) );
  XNOR2_X1 U558 ( .A(n388), .B(b[7]), .ZN(n214) );
  XNOR2_X1 U559 ( .A(n388), .B(b[2]), .ZN(n219) );
  XNOR2_X1 U560 ( .A(n388), .B(b[5]), .ZN(n216) );
  XNOR2_X1 U561 ( .A(n333), .B(b[6]), .ZN(n215) );
  XNOR2_X1 U562 ( .A(n333), .B(b[3]), .ZN(n218) );
  XNOR2_X1 U563 ( .A(n333), .B(b[4]), .ZN(n217) );
  XNOR2_X1 U564 ( .A(n388), .B(n248), .ZN(n221) );
  INV_X1 U565 ( .A(n333), .ZN(n262) );
  XNOR2_X1 U566 ( .A(n388), .B(b[1]), .ZN(n220) );
  XOR2_X1 U567 ( .A(n266), .B(a[4]), .Z(n250) );
  INV_X1 U568 ( .A(n1), .ZN(n68) );
  OAI21_X1 U569 ( .B1(n376), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U570 ( .B1(n46), .B2(n358), .A(n47), .ZN(n45) );
  OAI21_X1 U571 ( .B1(n376), .B2(n37), .A(n38), .ZN(n36) );
  OAI21_X1 U572 ( .B1(n26), .B2(n358), .A(n27), .ZN(n25) );
  AOI21_X1 U573 ( .B1(n68), .B2(n64), .A(n65), .ZN(n63) );
  AOI21_X1 U574 ( .B1(n380), .B2(n86), .A(n83), .ZN(n81) );
  INV_X2 U575 ( .A(n167), .ZN(n276) );
endmodule


module datapath ( clk, data_in, addr_x, wr_en_x, addr_a, wr_en_a, addr_y, 
        wr_en_y, clear_acc, data_out );
  input [7:0] data_in;
  input [3:0] addr_x;
  input [7:0] addr_a;
  input [3:0] addr_y;
  output [15:0] data_out;
  input clk, wr_en_x, wr_en_a, wr_en_y, clear_acc;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, n2;
  wire   [7:0] data_out_x;
  wire   [7:0] data_out_a;
  wire   [15:0] f;
  wire   [15:0] mul_out_r;
  wire   [15:0] add_r;
  wire   [15:0] mul_out;

  DFF_X1 \mul_out_r_reg[15]  ( .D(N34), .CK(clk), .Q(mul_out_r[15]) );
  DFF_X1 \mul_out_r_reg[14]  ( .D(N33), .CK(clk), .Q(mul_out_r[14]) );
  DFF_X1 \mul_out_r_reg[9]  ( .D(N28), .CK(clk), .Q(mul_out_r[9]) );
  DFF_X1 \mul_out_r_reg[8]  ( .D(N27), .CK(clk), .Q(mul_out_r[8]) );
  DFF_X1 \mul_out_r_reg[7]  ( .D(N26), .CK(clk), .Q(mul_out_r[7]) );
  DFF_X1 \mul_out_r_reg[6]  ( .D(N25), .CK(clk), .Q(mul_out_r[6]) );
  DFF_X1 \mul_out_r_reg[5]  ( .D(N24), .CK(clk), .Q(mul_out_r[5]) );
  DFF_X1 \mul_out_r_reg[4]  ( .D(N23), .CK(clk), .Q(mul_out_r[4]) );
  DFF_X1 \mul_out_r_reg[3]  ( .D(N22), .CK(clk), .Q(mul_out_r[3]) );
  DFF_X1 \mul_out_r_reg[2]  ( .D(N21), .CK(clk), .Q(mul_out_r[2]) );
  DFF_X1 \mul_out_r_reg[1]  ( .D(N20), .CK(clk), .Q(mul_out_r[1]) );
  DFF_X1 \mul_out_r_reg[0]  ( .D(N19), .CK(clk), .Q(mul_out_r[0]) );
  DFF_X1 \f_reg[0]  ( .D(N3), .CK(clk), .Q(f[0]) );
  DFF_X1 \f_reg[1]  ( .D(N4), .CK(clk), .Q(f[1]) );
  DFF_X1 \f_reg[2]  ( .D(N5), .CK(clk), .Q(f[2]) );
  DFF_X1 \f_reg[3]  ( .D(N6), .CK(clk), .Q(f[3]) );
  DFF_X1 \f_reg[4]  ( .D(N7), .CK(clk), .Q(f[4]) );
  DFF_X1 \f_reg[5]  ( .D(N8), .CK(clk), .Q(f[5]) );
  DFF_X1 \f_reg[6]  ( .D(N9), .CK(clk), .Q(f[6]) );
  DFF_X1 \f_reg[7]  ( .D(N10), .CK(clk), .Q(f[7]) );
  DFF_X1 \f_reg[8]  ( .D(N11), .CK(clk), .Q(f[8]) );
  DFF_X1 \f_reg[9]  ( .D(N12), .CK(clk), .Q(f[9]) );
  DFF_X1 \f_reg[10]  ( .D(N13), .CK(clk), .Q(f[10]) );
  DFF_X1 \f_reg[11]  ( .D(N14), .CK(clk), .Q(f[11]) );
  DFF_X1 \f_reg[12]  ( .D(N15), .CK(clk), .Q(f[12]) );
  DFF_X1 \f_reg[13]  ( .D(N16), .CK(clk), .Q(f[13]) );
  DFF_X1 \f_reg[14]  ( .D(N17), .CK(clk), .Q(f[14]) );
  memory_WIDTH8_SIZE16_LOGSIZE4 mem_x ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_x), .addr(addr_x), .wr_en(wr_en_x) );
  memory_WIDTH8_SIZE256_LOGSIZE8 mem_a ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a), .addr(addr_a), .wr_en(wr_en_a) );
  memory_WIDTH16_SIZE16_LOGSIZE4 mem_y ( .clk(clk), .data_in(f), .data_out(
        data_out), .addr(addr_y), .wr_en(wr_en_y) );
  datapath_DW01_add_1 add_68 ( .A(f), .B(mul_out_r), .CI(1'b0), .SUM(add_r) );
  datapath_DW_mult_tc_1 mult_67 ( .a(data_out_a), .b(data_out_x), .product(
        mul_out) );
  DFF_X1 \mul_out_r_reg[10]  ( .D(N29), .CK(clk), .Q(mul_out_r[10]) );
  DFF_X1 \mul_out_r_reg[12]  ( .D(N31), .CK(clk), .Q(mul_out_r[12]) );
  DFF_X2 \f_reg[15]  ( .D(N18), .CK(clk), .Q(f[15]) );
  DFF_X1 \mul_out_r_reg[13]  ( .D(N32), .CK(clk), .Q(mul_out_r[13]) );
  DFF_X1 \mul_out_r_reg[11]  ( .D(N30), .CK(clk), .Q(mul_out_r[11]) );
  INV_X1 U3 ( .A(clear_acc), .ZN(n2) );
  AND2_X1 U4 ( .A1(add_r[14]), .A2(n2), .ZN(N17) );
  AND2_X1 U5 ( .A1(add_r[13]), .A2(n2), .ZN(N16) );
  AND2_X1 U7 ( .A1(add_r[12]), .A2(n2), .ZN(N15) );
  AND2_X1 U8 ( .A1(add_r[11]), .A2(n2), .ZN(N14) );
  AND2_X1 U9 ( .A1(add_r[10]), .A2(n2), .ZN(N13) );
  AND2_X1 U10 ( .A1(add_r[9]), .A2(n2), .ZN(N12) );
  AND2_X1 U11 ( .A1(add_r[8]), .A2(n2), .ZN(N11) );
  AND2_X1 U12 ( .A1(add_r[7]), .A2(n2), .ZN(N10) );
  AND2_X1 U13 ( .A1(add_r[6]), .A2(n2), .ZN(N9) );
  AND2_X1 U14 ( .A1(add_r[5]), .A2(n2), .ZN(N8) );
  AND2_X1 U15 ( .A1(add_r[4]), .A2(n2), .ZN(N7) );
  AND2_X1 U16 ( .A1(add_r[3]), .A2(n2), .ZN(N6) );
  AND2_X1 U17 ( .A1(add_r[2]), .A2(n2), .ZN(N5) );
  AND2_X1 U18 ( .A1(add_r[1]), .A2(n2), .ZN(N4) );
  AND2_X1 U19 ( .A1(add_r[0]), .A2(n2), .ZN(N3) );
  AND2_X1 U20 ( .A1(mul_out[15]), .A2(n2), .ZN(N34) );
  AND2_X1 U21 ( .A1(mul_out[14]), .A2(n2), .ZN(N33) );
  AND2_X1 U22 ( .A1(mul_out[13]), .A2(n2), .ZN(N32) );
  AND2_X1 U23 ( .A1(mul_out[12]), .A2(n2), .ZN(N31) );
  AND2_X1 U24 ( .A1(mul_out[11]), .A2(n2), .ZN(N30) );
  AND2_X1 U25 ( .A1(mul_out[10]), .A2(n2), .ZN(N29) );
  AND2_X1 U26 ( .A1(mul_out[9]), .A2(n2), .ZN(N28) );
  AND2_X1 U27 ( .A1(mul_out[8]), .A2(n2), .ZN(N27) );
  AND2_X1 U28 ( .A1(mul_out[7]), .A2(n2), .ZN(N26) );
  AND2_X1 U29 ( .A1(mul_out[6]), .A2(n2), .ZN(N25) );
  AND2_X1 U30 ( .A1(mul_out[5]), .A2(n2), .ZN(N24) );
  AND2_X1 U31 ( .A1(mul_out[4]), .A2(n2), .ZN(N23) );
  AND2_X1 U32 ( .A1(mul_out[3]), .A2(n2), .ZN(N22) );
  AND2_X1 U33 ( .A1(mul_out[2]), .A2(n2), .ZN(N21) );
  AND2_X1 U34 ( .A1(mul_out[1]), .A2(n2), .ZN(N20) );
  AND2_X1 U35 ( .A1(mul_out[0]), .A2(n2), .ZN(N19) );
  AND2_X1 U36 ( .A1(add_r[15]), .A2(n2), .ZN(N18) );
endmodule


module ctrlpath_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[0]), .ZN(SUM[0]) );
  XOR2_X1 U2 ( .A(carry[7]), .B(A[7]), .Z(SUM[7]) );
endmodule


module ctrlpath ( clk, reset, start, addr_x, wr_en_x, addr_a, wr_en_a, 
        clear_acc, addr_y, wr_en_y, done, loadMatrix, loadVector );
  output [3:0] addr_x;
  output [7:0] addr_a;
  output [3:0] addr_y;
  input clk, reset, start, loadMatrix, loadVector;
  output wr_en_x, wr_en_a, clear_acc, wr_en_y, done;
  wire   N17, N18, N19, N20, N21, N25, N26, N27, N28, N29, N30, N31, N32, N49,
         N50, N51, N52, N61, N62, N63, N64, N67, N74, n42, n43, n44, n46, n47,
         n48, n49, n51, n52, n53, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32;
  wire   [3:0] state;

  DFF_X1 \addr_y_reg[0]  ( .D(N61), .CK(clk), .Q(addr_y[0]), .QN(n53) );
  DFF_X1 \addr_y_reg[2]  ( .D(N63), .CK(clk), .Q(addr_y[2]), .QN(n51) );
  DFF_X1 \state_reg[0]  ( .D(N17), .CK(clk), .Q(state[0]), .QN(n44) );
  DFF_X1 \state_reg[3]  ( .D(N20), .CK(clk), .Q(state[3]) );
  DFF_X1 \addr_x_reg[0]  ( .D(N49), .CK(clk), .Q(addr_x[0]) );
  DFF_X1 \addr_x_reg[1]  ( .D(N50), .CK(clk), .Q(addr_x[1]), .QN(n48) );
  DFF_X1 \addr_x_reg[2]  ( .D(N51), .CK(clk), .Q(addr_x[2]), .QN(n47) );
  DFF_X1 \addr_x_reg[3]  ( .D(N52), .CK(clk), .Q(addr_x[3]), .QN(n46) );
  DFF_X1 \state_reg[1]  ( .D(N18), .CK(clk), .Q(state[1]), .QN(n43) );
  DFF_X1 done_reg ( .D(N21), .CK(clk), .Q(done) );
  DFF_X1 \state_reg[2]  ( .D(N19), .CK(clk), .Q(state[2]), .QN(n42) );
  DFF_X1 \addr_y_reg[1]  ( .D(N62), .CK(clk), .Q(addr_y[1]), .QN(n52) );
  DFF_X1 \addr_y_reg[3]  ( .D(N64), .CK(clk), .Q(addr_y[3]), .QN(n49) );
  DFF_X1 \addr_a_reg[0]  ( .D(n10), .CK(clk), .Q(addr_a[0]), .QN(n1) );
  DFF_X1 \addr_a_reg[1]  ( .D(n11), .CK(clk), .Q(addr_a[1]) );
  DFF_X1 \addr_a_reg[2]  ( .D(n12), .CK(clk), .Q(addr_a[2]) );
  DFF_X1 \addr_a_reg[3]  ( .D(n13), .CK(clk), .Q(addr_a[3]) );
  DFF_X1 \addr_a_reg[4]  ( .D(n14), .CK(clk), .Q(addr_a[4]) );
  DFF_X1 \addr_a_reg[5]  ( .D(n15), .CK(clk), .Q(addr_a[5]) );
  DFF_X1 \addr_a_reg[7]  ( .D(n17), .CK(clk), .Q(addr_a[7]) );
  DFF_X1 clear_acc_reg ( .D(N67), .CK(clk), .Q(clear_acc) );
  NOR2_X2 U35 ( .A1(n91), .A2(reset), .ZN(wr_en_a) );
  NAND3_X1 U95 ( .A1(n57), .A2(n49), .A3(n28), .ZN(n56) );
  NAND3_X1 U96 ( .A1(addr_y[0]), .A2(n52), .A3(n28), .ZN(n62) );
  NAND3_X1 U97 ( .A1(n63), .A2(n60), .A3(addr_y[0]), .ZN(n64) );
  XOR2_X1 U98 ( .A(addr_x[0]), .B(n48), .Z(n70) );
  NAND3_X1 U100 ( .A1(n89), .A2(n90), .A3(N74), .ZN(n88) );
  NAND3_X1 U101 ( .A1(n91), .A2(n29), .A3(n89), .ZN(n73) );
  NAND3_X1 U102 ( .A1(n72), .A2(n87), .A3(n95), .ZN(N67) );
  XOR2_X1 U103 ( .A(n44), .B(state[1]), .Z(n99) );
  NAND3_X1 U104 ( .A1(n44), .A2(n43), .A3(n65), .ZN(n86) );
  NAND3_X1 U105 ( .A1(n114), .A2(n42), .A3(state[3]), .ZN(n85) );
  NAND3_X1 U106 ( .A1(n113), .A2(n42), .A3(state[3]), .ZN(n95) );
  NAND3_X1 U107 ( .A1(n44), .A2(n43), .A3(n112), .ZN(n63) );
  NAND3_X1 U108 ( .A1(state[1]), .A2(state[0]), .A3(n112), .ZN(n90) );
  NAND3_X1 U109 ( .A1(addr_x[1]), .A2(addr_x[0]), .A3(addr_x[2]), .ZN(n66) );
  ctrlpath_DW01_inc_0 add_103 ( .A({addr_a[7:1], n2}), .SUM({N32, N31, N30, 
        N29, N28, N27, N26, N25}) );
  DFF_X2 \addr_a_reg[6]  ( .D(n16), .CK(clk), .Q(addr_a[6]) );
  NOR2_X1 U3 ( .A1(n42), .A2(state[3]), .ZN(n65) );
  INV_X1 U4 ( .A(n1), .ZN(n2) );
  INV_X1 U5 ( .A(n69), .ZN(n19) );
  INV_X1 U6 ( .A(n72), .ZN(n26) );
  INV_X1 U7 ( .A(n110), .ZN(n23) );
  INV_X1 U8 ( .A(n96), .ZN(n29) );
  INV_X1 U9 ( .A(n107), .ZN(n6) );
  NOR2_X1 U10 ( .A1(n76), .A2(n84), .ZN(n75) );
  AND4_X1 U11 ( .A1(n85), .A2(n86), .A3(n87), .A4(n29), .ZN(n84) );
  NAND3_X1 U12 ( .A1(n73), .A2(n18), .A3(n88), .ZN(n76) );
  INV_X1 U13 ( .A(wr_en_y), .ZN(n18) );
  OAI21_X1 U14 ( .B1(n71), .B2(n72), .A(n73), .ZN(n69) );
  AOI22_X1 U15 ( .A1(n65), .A2(n114), .B1(n102), .B2(n30), .ZN(n107) );
  INV_X1 U16 ( .A(n94), .ZN(n30) );
  NAND2_X1 U17 ( .A1(n65), .A2(n113), .ZN(n87) );
  NOR2_X1 U18 ( .A1(n31), .A2(n90), .ZN(n96) );
  NOR2_X1 U19 ( .A1(n102), .A2(n87), .ZN(N21) );
  INV_X1 U20 ( .A(n60), .ZN(n28) );
  NAND2_X1 U21 ( .A1(n112), .A2(n114), .ZN(n72) );
  NAND2_X1 U22 ( .A1(n63), .A2(n95), .ZN(n110) );
  NAND2_X1 U23 ( .A1(n107), .A2(n85), .ZN(n101) );
  NAND2_X1 U24 ( .A1(n112), .A2(n113), .ZN(n91) );
  INV_X1 U25 ( .A(n71), .ZN(n31) );
  INV_X1 U26 ( .A(n86), .ZN(n25) );
  AND4_X1 U27 ( .A1(n92), .A2(n20), .A3(n63), .A4(n93), .ZN(n89) );
  AND3_X1 U28 ( .A1(n94), .A2(n86), .A3(n85), .ZN(n93) );
  INV_X1 U29 ( .A(N67), .ZN(n20) );
  INV_X1 U30 ( .A(n92), .ZN(n24) );
  OAI21_X1 U31 ( .B1(state[1]), .B2(state[0]), .A(n65), .ZN(n60) );
  NOR4_X1 U32 ( .A1(start), .A2(loadVector), .A3(loadMatrix), .A4(n95), .ZN(
        n98) );
  OAI222_X1 U33 ( .A1(n31), .A2(n27), .B1(reset), .B2(n97), .C1(N74), .C2(n22), 
        .ZN(N20) );
  INV_X1 U34 ( .A(wr_en_x), .ZN(n27) );
  NOR3_X1 U36 ( .A1(n98), .A2(n24), .A3(n25), .ZN(n97) );
  INV_X1 U37 ( .A(wr_en_a), .ZN(n22) );
  NOR2_X1 U38 ( .A1(n46), .A2(n66), .ZN(n71) );
  OAI22_X1 U39 ( .A1(n71), .A2(n90), .B1(n23), .B2(n32), .ZN(n106) );
  INV_X1 U40 ( .A(start), .ZN(n32) );
  AOI21_X1 U41 ( .B1(n103), .B2(n104), .A(reset), .ZN(N18) );
  AOI211_X1 U42 ( .C1(n105), .C2(loadVector), .A(n9), .B(n25), .ZN(n104) );
  AOI211_X1 U43 ( .C1(n26), .C2(n31), .A(n106), .B(n6), .ZN(n103) );
  INV_X1 U44 ( .A(n87), .ZN(n9) );
  NOR3_X1 U45 ( .A1(n52), .A2(n53), .A3(n51), .ZN(n57) );
  AOI22_X1 U46 ( .A1(n53), .A2(n28), .B1(n60), .B2(n63), .ZN(n61) );
  NOR2_X1 U47 ( .A1(state[3]), .A2(state[2]), .ZN(n112) );
  NAND2_X1 U48 ( .A1(addr_y[3]), .A2(n57), .ZN(n102) );
  OAI22_X1 U49 ( .A1(loadVector), .A2(n95), .B1(n5), .B2(n87), .ZN(n111) );
  INV_X1 U50 ( .A(n102), .ZN(n5) );
  NOR2_X1 U51 ( .A1(n44), .A2(state[1]), .ZN(n113) );
  NOR2_X1 U52 ( .A1(n87), .A2(reset), .ZN(wr_en_y) );
  NOR2_X1 U53 ( .A1(n43), .A2(state[0]), .ZN(n114) );
  NOR2_X1 U54 ( .A1(n72), .A2(reset), .ZN(wr_en_x) );
  OAI21_X1 U55 ( .B1(addr_y[1]), .B2(n60), .A(n61), .ZN(n58) );
  OAI21_X1 U56 ( .B1(state[2]), .B2(n99), .A(state[3]), .ZN(n92) );
  OAI22_X1 U57 ( .A1(n19), .A2(n46), .B1(n19), .B2(n66), .ZN(N52) );
  NOR2_X1 U58 ( .A1(n19), .A2(addr_x[0]), .ZN(N49) );
  OAI21_X1 U59 ( .B1(addr_y[0]), .B2(n60), .A(n64), .ZN(N61) );
  AOI21_X1 U60 ( .B1(n100), .B2(n7), .A(reset), .ZN(N19) );
  INV_X1 U61 ( .A(n101), .ZN(n7) );
  NOR2_X1 U62 ( .A1(N21), .A2(n96), .ZN(n100) );
  AOI21_X1 U63 ( .B1(n108), .B2(n109), .A(reset), .ZN(N17) );
  AOI211_X1 U64 ( .C1(loadMatrix), .C2(n110), .A(n111), .B(n21), .ZN(n109) );
  AOI211_X1 U65 ( .C1(n71), .C2(n26), .A(n106), .B(n101), .ZN(n108) );
  INV_X1 U66 ( .A(n91), .ZN(n21) );
  NOR2_X1 U67 ( .A1(loadMatrix), .A2(n23), .ZN(n105) );
  OAI21_X1 U68 ( .B1(n61), .B2(n52), .A(n62), .ZN(N62) );
  NAND2_X1 U69 ( .A1(state[1]), .A2(n65), .ZN(n94) );
  OAI21_X1 U70 ( .B1(n67), .B2(n47), .A(n68), .ZN(N51) );
  NAND4_X1 U71 ( .A1(addr_x[1]), .A2(addr_x[0]), .A3(n69), .A4(n47), .ZN(n68)
         );
  AOI21_X1 U72 ( .B1(n69), .B2(n48), .A(N49), .ZN(n67) );
  OAI21_X1 U73 ( .B1(n55), .B2(n49), .A(n56), .ZN(N64) );
  AOI21_X1 U74 ( .B1(n28), .B2(n51), .A(n58), .ZN(n55) );
  NOR2_X1 U75 ( .A1(n19), .A2(n70), .ZN(N50) );
  INV_X1 U76 ( .A(n77), .ZN(n16) );
  AOI22_X1 U77 ( .A1(addr_a[6]), .A2(n75), .B1(N31), .B2(n76), .ZN(n77) );
  OAI21_X1 U78 ( .B1(n8), .B2(n51), .A(n59), .ZN(N63) );
  NAND4_X1 U79 ( .A1(n28), .A2(addr_y[1]), .A3(addr_y[0]), .A4(n51), .ZN(n59)
         );
  INV_X1 U80 ( .A(n58), .ZN(n8) );
  INV_X1 U81 ( .A(n74), .ZN(n17) );
  AOI22_X1 U82 ( .A1(addr_a[7]), .A2(n75), .B1(N32), .B2(n76), .ZN(n74) );
  INV_X1 U83 ( .A(n83), .ZN(n10) );
  INV_X1 U84 ( .A(n78), .ZN(n15) );
  AOI22_X1 U85 ( .A1(addr_a[5]), .A2(n75), .B1(N30), .B2(n76), .ZN(n78) );
  INV_X1 U86 ( .A(n79), .ZN(n14) );
  AOI22_X1 U87 ( .A1(addr_a[4]), .A2(n75), .B1(N29), .B2(n76), .ZN(n79) );
  INV_X1 U88 ( .A(n80), .ZN(n13) );
  AOI22_X1 U89 ( .A1(addr_a[3]), .A2(n75), .B1(N28), .B2(n76), .ZN(n80) );
  INV_X1 U90 ( .A(n81), .ZN(n12) );
  AOI22_X1 U91 ( .A1(addr_a[2]), .A2(n75), .B1(N27), .B2(n76), .ZN(n81) );
  INV_X1 U92 ( .A(n82), .ZN(n11) );
  AOI22_X1 U93 ( .A1(addr_a[1]), .A2(n75), .B1(N26), .B2(n76), .ZN(n82) );
  AOI22_X1 U94 ( .A1(n2), .A2(n75), .B1(N25), .B2(n76), .ZN(n83) );
  NAND4_X1 U99 ( .A1(addr_a[3]), .A2(addr_a[2]), .A3(addr_a[1]), .A4(n2), .ZN(
        n4) );
  NAND4_X1 U110 ( .A1(addr_a[7]), .A2(addr_a[6]), .A3(addr_a[5]), .A4(
        addr_a[4]), .ZN(n3) );
  OR2_X1 U111 ( .A1(n4), .A2(n3), .ZN(N74) );
endmodule


module mvm_16_1_8_1 ( clk, reset, loadMatrix, loadVector, start, done, data_in, 
        data_out );
  input [7:0] data_in;
  output [15:0] data_out;
  input clk, reset, loadMatrix, loadVector, start;
  output done;
  wire   wr_en_x, wr_en_a, wr_en_y, clear_acc;
  wire   [3:0] addr_x;
  wire   [7:0] addr_a;
  wire   [3:0] addr_y;

  datapath d ( .clk(clk), .data_in(data_in), .addr_x(addr_x), .wr_en_x(wr_en_x), .addr_a(addr_a), .wr_en_a(wr_en_a), .addr_y(addr_y), .wr_en_y(wr_en_y), 
        .clear_acc(clear_acc), .data_out(data_out) );
  ctrlpath c ( .clk(clk), .reset(reset), .start(start), .addr_x(addr_x), 
        .wr_en_x(wr_en_x), .addr_a(addr_a), .wr_en_a(wr_en_a), .clear_acc(
        clear_acc), .addr_y(addr_y), .wr_en_y(wr_en_y), .done(done), 
        .loadMatrix(loadMatrix), .loadVector(loadVector) );
endmodule

