
module memory_WIDTH20_SIZE8_LOGSIZE3_0 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \mem_reg[7][19]  ( .D(n353), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n352), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n351), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n350), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n349), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n348), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n347), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n346), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n345), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n344), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n343), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n342), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n341), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n340), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n339), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n338), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n337), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n336), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n335), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n334), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n333), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n332), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n331), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n330), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n329), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n328), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n327), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n326), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n325), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n324), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n323), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n322), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n321), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n320), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n319), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n318), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n317), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n316), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n315), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n314), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n313), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n312), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n311), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n310), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n309), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n308), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n307), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n306), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n305), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n304), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n303), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n302), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n301), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n300), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n299), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n298), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n297), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n296), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n295), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n294), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n293), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n292), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n291), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n290), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n289), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n288), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n287), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n286), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n285), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n284), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n283), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n282), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n281), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n280), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n279), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n278), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n277), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n276), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n275), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n274), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n273), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n272), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n271), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n270), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n269), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n268), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n267), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n266), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n265), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n264), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n263), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n262), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n261), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n260), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n259), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n258), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n257), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n256), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n255), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n254), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n253), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n252), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n251), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n250), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n249), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n248), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n247), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n246), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n245), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n244), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n243), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n242), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n241), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n240), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n239), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n238), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n237), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n236), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n235), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n234), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n233), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n232), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n231), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n230), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n229), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n228), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n227), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n226), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n225), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n224), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n223), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n222), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n221), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n220), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n219), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n218), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n217), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n216), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n215), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n214), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n213), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n212), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n211), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n210), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n209), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n208), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n207), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n206), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n205), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n204), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n203), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n202), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n201), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n200), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n199), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n198), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n197), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n196), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n195), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n194), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U348 ( .A1(n468), .A2(n469), .A3(n45), .ZN(n24) );
  NAND3_X1 U349 ( .A1(n45), .A2(n469), .A3(N10), .ZN(n46) );
  NAND3_X1 U350 ( .A1(n45), .A2(n468), .A3(N11), .ZN(n67) );
  NAND3_X1 U351 ( .A1(N10), .A2(n45), .A3(N11), .ZN(n88) );
  NAND3_X1 U352 ( .A1(n468), .A2(n469), .A3(n130), .ZN(n109) );
  NAND3_X1 U353 ( .A1(N10), .A2(n469), .A3(n130), .ZN(n131) );
  NAND3_X1 U354 ( .A1(N11), .A2(n468), .A3(n130), .ZN(n152) );
  NAND3_X1 U355 ( .A1(N11), .A2(N10), .A3(n130), .ZN(n173) );
  SDFF_X1 \data_out_reg[4]  ( .D(n364), .SI(n361), .SE(N12), .CK(clk), .Q(
        data_out[4]) );
  SDFF_X1 \data_out_reg[2]  ( .D(n22), .SI(n19), .SE(N12), .CK(clk), .Q(
        data_out[2]) );
  SDFF_X1 \data_out_reg[12]  ( .D(n412), .SI(n409), .SE(N12), .CK(clk), .Q(
        data_out[12]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n16), .SI(n13), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[18]  ( .D(n448), .SI(n445), .SE(N12), .CK(clk), .Q(
        data_out[18]) );
  SDFF_X1 \data_out_reg[10]  ( .D(n400), .SI(n397), .SE(N12), .CK(clk), .Q(
        data_out[10]) );
  SDFF_X1 \data_out_reg[16]  ( .D(n436), .SI(n433), .SE(N12), .CK(clk), .Q(
        data_out[16]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n394), .SI(n391), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[6]  ( .D(n376), .SI(n373), .SE(N12), .CK(clk), .Q(
        data_out[6]) );
  SDFF_X1 \data_out_reg[14]  ( .D(n424), .SI(n421), .SE(N12), .CK(clk), .Q(
        data_out[14]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n418), .SI(n415), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[19]  ( .D(n454), .SI(n451), .SE(N12), .CK(clk), .Q(
        data_out[19]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n430), .SI(n427), .SE(N12), .CK(clk), .Q(
        data_out[15]) );
  SDFF_X1 \data_out_reg[8]  ( .D(n388), .SI(n385), .SE(N12), .CK(clk), .Q(
        data_out[8]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n358), .SI(n355), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n10), .SI(n7), .SE(N12), .CK(clk), .Q(
        data_out[0]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n370), .SI(n367), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n382), .SI(n379), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n406), .SI(n403), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[17]  ( .D(n442), .SI(n439), .SE(N12), .CK(clk), .Q(
        data_out[17]) );
  BUF_X1 U3 ( .A(n67), .Z(n465) );
  BUF_X1 U4 ( .A(n88), .Z(n464) );
  BUF_X1 U5 ( .A(n173), .Z(n460) );
  BUF_X1 U6 ( .A(n109), .Z(n463) );
  BUF_X1 U7 ( .A(n456), .Z(n455) );
  BUF_X1 U8 ( .A(n24), .Z(n467) );
  BUF_X1 U9 ( .A(n46), .Z(n466) );
  BUF_X1 U10 ( .A(n131), .Z(n462) );
  BUF_X1 U11 ( .A(n152), .Z(n461) );
  BUF_X1 U12 ( .A(N10), .Z(n457) );
  BUF_X1 U13 ( .A(N10), .Z(n458) );
  BUF_X1 U14 ( .A(N10), .Z(n459) );
  BUF_X1 U15 ( .A(N11), .Z(n456) );
  NOR2_X1 U16 ( .A1(n470), .A2(N12), .ZN(n45) );
  INV_X1 U17 ( .A(wr_en), .ZN(n470) );
  AND2_X1 U18 ( .A1(N12), .A2(wr_en), .ZN(n130) );
  OAI21_X1 U19 ( .B1(n490), .B2(n46), .A(n47), .ZN(n214) );
  NAND2_X1 U20 ( .A1(\mem[1][0] ), .A2(n466), .ZN(n47) );
  OAI21_X1 U21 ( .B1(n489), .B2(n46), .A(n48), .ZN(n215) );
  NAND2_X1 U22 ( .A1(\mem[1][1] ), .A2(n466), .ZN(n48) );
  OAI21_X1 U23 ( .B1(n488), .B2(n46), .A(n49), .ZN(n216) );
  NAND2_X1 U24 ( .A1(\mem[1][2] ), .A2(n466), .ZN(n49) );
  OAI21_X1 U25 ( .B1(n487), .B2(n46), .A(n50), .ZN(n217) );
  NAND2_X1 U26 ( .A1(\mem[1][3] ), .A2(n466), .ZN(n50) );
  OAI21_X1 U27 ( .B1(n486), .B2(n466), .A(n51), .ZN(n218) );
  NAND2_X1 U28 ( .A1(\mem[1][4] ), .A2(n466), .ZN(n51) );
  OAI21_X1 U29 ( .B1(n485), .B2(n466), .A(n52), .ZN(n219) );
  NAND2_X1 U30 ( .A1(\mem[1][5] ), .A2(n466), .ZN(n52) );
  OAI21_X1 U31 ( .B1(n484), .B2(n46), .A(n53), .ZN(n220) );
  NAND2_X1 U32 ( .A1(\mem[1][6] ), .A2(n466), .ZN(n53) );
  OAI21_X1 U33 ( .B1(n483), .B2(n46), .A(n54), .ZN(n221) );
  NAND2_X1 U34 ( .A1(\mem[1][7] ), .A2(n466), .ZN(n54) );
  OAI21_X1 U35 ( .B1(n482), .B2(n46), .A(n55), .ZN(n222) );
  NAND2_X1 U36 ( .A1(\mem[1][8] ), .A2(n466), .ZN(n55) );
  OAI21_X1 U37 ( .B1(n481), .B2(n46), .A(n56), .ZN(n223) );
  NAND2_X1 U38 ( .A1(\mem[1][9] ), .A2(n466), .ZN(n56) );
  OAI21_X1 U39 ( .B1(n480), .B2(n46), .A(n57), .ZN(n224) );
  NAND2_X1 U40 ( .A1(\mem[1][10] ), .A2(n466), .ZN(n57) );
  OAI21_X1 U41 ( .B1(n479), .B2(n46), .A(n58), .ZN(n225) );
  NAND2_X1 U42 ( .A1(\mem[1][11] ), .A2(n466), .ZN(n58) );
  OAI21_X1 U43 ( .B1(n478), .B2(n46), .A(n59), .ZN(n226) );
  NAND2_X1 U44 ( .A1(\mem[1][12] ), .A2(n46), .ZN(n59) );
  OAI21_X1 U45 ( .B1(n477), .B2(n46), .A(n60), .ZN(n227) );
  NAND2_X1 U46 ( .A1(\mem[1][13] ), .A2(n46), .ZN(n60) );
  OAI21_X1 U47 ( .B1(n476), .B2(n46), .A(n61), .ZN(n228) );
  NAND2_X1 U48 ( .A1(\mem[1][14] ), .A2(n46), .ZN(n61) );
  OAI21_X1 U49 ( .B1(n475), .B2(n46), .A(n62), .ZN(n229) );
  NAND2_X1 U50 ( .A1(\mem[1][15] ), .A2(n466), .ZN(n62) );
  OAI21_X1 U51 ( .B1(n474), .B2(n46), .A(n63), .ZN(n230) );
  NAND2_X1 U52 ( .A1(\mem[1][16] ), .A2(n46), .ZN(n63) );
  OAI21_X1 U53 ( .B1(n473), .B2(n46), .A(n64), .ZN(n231) );
  NAND2_X1 U54 ( .A1(\mem[1][17] ), .A2(n46), .ZN(n64) );
  OAI21_X1 U55 ( .B1(n472), .B2(n46), .A(n65), .ZN(n232) );
  NAND2_X1 U56 ( .A1(\mem[1][18] ), .A2(n46), .ZN(n65) );
  OAI21_X1 U57 ( .B1(n471), .B2(n46), .A(n66), .ZN(n233) );
  NAND2_X1 U58 ( .A1(\mem[1][19] ), .A2(n466), .ZN(n66) );
  OAI21_X1 U59 ( .B1(n490), .B2(n465), .A(n68), .ZN(n234) );
  NAND2_X1 U60 ( .A1(\mem[2][0] ), .A2(n465), .ZN(n68) );
  OAI21_X1 U61 ( .B1(n489), .B2(n465), .A(n69), .ZN(n235) );
  NAND2_X1 U62 ( .A1(\mem[2][1] ), .A2(n465), .ZN(n69) );
  OAI21_X1 U63 ( .B1(n488), .B2(n465), .A(n70), .ZN(n236) );
  NAND2_X1 U64 ( .A1(\mem[2][2] ), .A2(n67), .ZN(n70) );
  OAI21_X1 U65 ( .B1(n487), .B2(n67), .A(n71), .ZN(n237) );
  NAND2_X1 U66 ( .A1(\mem[2][3] ), .A2(n465), .ZN(n71) );
  OAI21_X1 U67 ( .B1(n486), .B2(n67), .A(n72), .ZN(n238) );
  NAND2_X1 U68 ( .A1(\mem[2][4] ), .A2(n465), .ZN(n72) );
  OAI21_X1 U69 ( .B1(n485), .B2(n67), .A(n73), .ZN(n239) );
  NAND2_X1 U70 ( .A1(\mem[2][5] ), .A2(n67), .ZN(n73) );
  OAI21_X1 U71 ( .B1(n484), .B2(n67), .A(n74), .ZN(n240) );
  NAND2_X1 U72 ( .A1(\mem[2][6] ), .A2(n67), .ZN(n74) );
  OAI21_X1 U73 ( .B1(n483), .B2(n67), .A(n75), .ZN(n241) );
  NAND2_X1 U74 ( .A1(\mem[2][7] ), .A2(n67), .ZN(n75) );
  OAI21_X1 U75 ( .B1(n482), .B2(n67), .A(n76), .ZN(n242) );
  NAND2_X1 U76 ( .A1(\mem[2][8] ), .A2(n67), .ZN(n76) );
  OAI21_X1 U77 ( .B1(n481), .B2(n465), .A(n77), .ZN(n243) );
  NAND2_X1 U78 ( .A1(\mem[2][9] ), .A2(n67), .ZN(n77) );
  OAI21_X1 U79 ( .B1(n480), .B2(n67), .A(n78), .ZN(n244) );
  NAND2_X1 U80 ( .A1(\mem[2][10] ), .A2(n67), .ZN(n78) );
  OAI21_X1 U81 ( .B1(n479), .B2(n67), .A(n79), .ZN(n245) );
  NAND2_X1 U82 ( .A1(\mem[2][11] ), .A2(n67), .ZN(n79) );
  OAI21_X1 U83 ( .B1(n478), .B2(n465), .A(n80), .ZN(n246) );
  NAND2_X1 U84 ( .A1(\mem[2][12] ), .A2(n465), .ZN(n80) );
  OAI21_X1 U85 ( .B1(n477), .B2(n465), .A(n81), .ZN(n247) );
  NAND2_X1 U86 ( .A1(\mem[2][13] ), .A2(n465), .ZN(n81) );
  OAI21_X1 U87 ( .B1(n476), .B2(n465), .A(n82), .ZN(n248) );
  NAND2_X1 U88 ( .A1(\mem[2][14] ), .A2(n465), .ZN(n82) );
  OAI21_X1 U89 ( .B1(n475), .B2(n67), .A(n83), .ZN(n249) );
  NAND2_X1 U90 ( .A1(\mem[2][15] ), .A2(n465), .ZN(n83) );
  OAI21_X1 U91 ( .B1(n474), .B2(n67), .A(n84), .ZN(n250) );
  NAND2_X1 U92 ( .A1(\mem[2][16] ), .A2(n465), .ZN(n84) );
  OAI21_X1 U93 ( .B1(n473), .B2(n67), .A(n85), .ZN(n251) );
  NAND2_X1 U94 ( .A1(\mem[2][17] ), .A2(n465), .ZN(n85) );
  OAI21_X1 U95 ( .B1(n472), .B2(n465), .A(n86), .ZN(n252) );
  NAND2_X1 U96 ( .A1(\mem[2][18] ), .A2(n465), .ZN(n86) );
  OAI21_X1 U97 ( .B1(n471), .B2(n465), .A(n87), .ZN(n253) );
  NAND2_X1 U98 ( .A1(\mem[2][19] ), .A2(n465), .ZN(n87) );
  OAI21_X1 U99 ( .B1(n490), .B2(n464), .A(n89), .ZN(n254) );
  NAND2_X1 U100 ( .A1(\mem[3][0] ), .A2(n464), .ZN(n89) );
  OAI21_X1 U101 ( .B1(n489), .B2(n464), .A(n90), .ZN(n255) );
  NAND2_X1 U102 ( .A1(\mem[3][1] ), .A2(n464), .ZN(n90) );
  OAI21_X1 U103 ( .B1(n488), .B2(n464), .A(n91), .ZN(n256) );
  NAND2_X1 U104 ( .A1(\mem[3][2] ), .A2(n88), .ZN(n91) );
  OAI21_X1 U105 ( .B1(n487), .B2(n88), .A(n92), .ZN(n257) );
  NAND2_X1 U106 ( .A1(\mem[3][3] ), .A2(n464), .ZN(n92) );
  OAI21_X1 U107 ( .B1(n486), .B2(n88), .A(n93), .ZN(n258) );
  NAND2_X1 U108 ( .A1(\mem[3][4] ), .A2(n464), .ZN(n93) );
  OAI21_X1 U109 ( .B1(n485), .B2(n88), .A(n94), .ZN(n259) );
  NAND2_X1 U110 ( .A1(\mem[3][5] ), .A2(n88), .ZN(n94) );
  OAI21_X1 U111 ( .B1(n484), .B2(n88), .A(n95), .ZN(n260) );
  NAND2_X1 U112 ( .A1(\mem[3][6] ), .A2(n88), .ZN(n95) );
  OAI21_X1 U113 ( .B1(n483), .B2(n88), .A(n96), .ZN(n261) );
  NAND2_X1 U114 ( .A1(\mem[3][7] ), .A2(n88), .ZN(n96) );
  OAI21_X1 U115 ( .B1(n482), .B2(n88), .A(n97), .ZN(n262) );
  NAND2_X1 U116 ( .A1(\mem[3][8] ), .A2(n88), .ZN(n97) );
  OAI21_X1 U117 ( .B1(n481), .B2(n464), .A(n98), .ZN(n263) );
  NAND2_X1 U118 ( .A1(\mem[3][9] ), .A2(n88), .ZN(n98) );
  OAI21_X1 U119 ( .B1(n480), .B2(n88), .A(n99), .ZN(n264) );
  NAND2_X1 U120 ( .A1(\mem[3][10] ), .A2(n88), .ZN(n99) );
  OAI21_X1 U121 ( .B1(n479), .B2(n88), .A(n100), .ZN(n265) );
  NAND2_X1 U122 ( .A1(\mem[3][11] ), .A2(n88), .ZN(n100) );
  OAI21_X1 U123 ( .B1(n478), .B2(n464), .A(n101), .ZN(n266) );
  NAND2_X1 U124 ( .A1(\mem[3][12] ), .A2(n464), .ZN(n101) );
  OAI21_X1 U125 ( .B1(n477), .B2(n464), .A(n102), .ZN(n267) );
  NAND2_X1 U126 ( .A1(\mem[3][13] ), .A2(n464), .ZN(n102) );
  OAI21_X1 U127 ( .B1(n476), .B2(n464), .A(n103), .ZN(n268) );
  NAND2_X1 U128 ( .A1(\mem[3][14] ), .A2(n464), .ZN(n103) );
  OAI21_X1 U129 ( .B1(n475), .B2(n88), .A(n104), .ZN(n269) );
  NAND2_X1 U130 ( .A1(\mem[3][15] ), .A2(n464), .ZN(n104) );
  OAI21_X1 U131 ( .B1(n474), .B2(n88), .A(n105), .ZN(n270) );
  NAND2_X1 U132 ( .A1(\mem[3][16] ), .A2(n464), .ZN(n105) );
  OAI21_X1 U133 ( .B1(n473), .B2(n88), .A(n106), .ZN(n271) );
  NAND2_X1 U134 ( .A1(\mem[3][17] ), .A2(n464), .ZN(n106) );
  OAI21_X1 U135 ( .B1(n472), .B2(n464), .A(n107), .ZN(n272) );
  NAND2_X1 U136 ( .A1(\mem[3][18] ), .A2(n464), .ZN(n107) );
  OAI21_X1 U137 ( .B1(n471), .B2(n464), .A(n108), .ZN(n273) );
  NAND2_X1 U138 ( .A1(\mem[3][19] ), .A2(n464), .ZN(n108) );
  OAI21_X1 U139 ( .B1(n490), .B2(n109), .A(n110), .ZN(n274) );
  NAND2_X1 U140 ( .A1(\mem[4][0] ), .A2(n109), .ZN(n110) );
  OAI21_X1 U141 ( .B1(n489), .B2(n463), .A(n111), .ZN(n275) );
  NAND2_X1 U142 ( .A1(\mem[4][1] ), .A2(n109), .ZN(n111) );
  OAI21_X1 U143 ( .B1(n488), .B2(n463), .A(n112), .ZN(n276) );
  NAND2_X1 U144 ( .A1(\mem[4][2] ), .A2(n109), .ZN(n112) );
  OAI21_X1 U145 ( .B1(n487), .B2(n463), .A(n113), .ZN(n277) );
  NAND2_X1 U146 ( .A1(\mem[4][3] ), .A2(n109), .ZN(n113) );
  OAI21_X1 U147 ( .B1(n486), .B2(n463), .A(n114), .ZN(n278) );
  NAND2_X1 U148 ( .A1(\mem[4][4] ), .A2(n109), .ZN(n114) );
  OAI21_X1 U149 ( .B1(n485), .B2(n463), .A(n115), .ZN(n279) );
  NAND2_X1 U150 ( .A1(\mem[4][5] ), .A2(n109), .ZN(n115) );
  OAI21_X1 U151 ( .B1(n484), .B2(n463), .A(n116), .ZN(n280) );
  NAND2_X1 U152 ( .A1(\mem[4][6] ), .A2(n109), .ZN(n116) );
  OAI21_X1 U153 ( .B1(n483), .B2(n463), .A(n117), .ZN(n281) );
  NAND2_X1 U154 ( .A1(\mem[4][7] ), .A2(n109), .ZN(n117) );
  OAI21_X1 U155 ( .B1(n482), .B2(n463), .A(n118), .ZN(n282) );
  NAND2_X1 U156 ( .A1(\mem[4][8] ), .A2(n109), .ZN(n118) );
  OAI21_X1 U157 ( .B1(n481), .B2(n109), .A(n119), .ZN(n283) );
  NAND2_X1 U158 ( .A1(\mem[4][9] ), .A2(n109), .ZN(n119) );
  OAI21_X1 U159 ( .B1(n480), .B2(n463), .A(n120), .ZN(n284) );
  NAND2_X1 U160 ( .A1(\mem[4][10] ), .A2(n109), .ZN(n120) );
  OAI21_X1 U161 ( .B1(n479), .B2(n463), .A(n121), .ZN(n285) );
  NAND2_X1 U162 ( .A1(\mem[4][11] ), .A2(n109), .ZN(n121) );
  OAI21_X1 U163 ( .B1(n478), .B2(n109), .A(n122), .ZN(n286) );
  NAND2_X1 U164 ( .A1(\mem[4][12] ), .A2(n109), .ZN(n122) );
  OAI21_X1 U165 ( .B1(n477), .B2(n463), .A(n123), .ZN(n287) );
  NAND2_X1 U166 ( .A1(\mem[4][13] ), .A2(n109), .ZN(n123) );
  OAI21_X1 U167 ( .B1(n476), .B2(n109), .A(n124), .ZN(n288) );
  NAND2_X1 U168 ( .A1(\mem[4][14] ), .A2(n109), .ZN(n124) );
  OAI21_X1 U169 ( .B1(n475), .B2(n463), .A(n125), .ZN(n289) );
  NAND2_X1 U170 ( .A1(\mem[4][15] ), .A2(n109), .ZN(n125) );
  OAI21_X1 U171 ( .B1(n474), .B2(n463), .A(n126), .ZN(n290) );
  NAND2_X1 U172 ( .A1(\mem[4][16] ), .A2(n109), .ZN(n126) );
  OAI21_X1 U173 ( .B1(n473), .B2(n463), .A(n127), .ZN(n291) );
  NAND2_X1 U174 ( .A1(\mem[4][17] ), .A2(n109), .ZN(n127) );
  OAI21_X1 U175 ( .B1(n472), .B2(n463), .A(n128), .ZN(n292) );
  NAND2_X1 U176 ( .A1(\mem[4][18] ), .A2(n109), .ZN(n128) );
  OAI21_X1 U177 ( .B1(n471), .B2(n463), .A(n129), .ZN(n293) );
  NAND2_X1 U178 ( .A1(\mem[4][19] ), .A2(n109), .ZN(n129) );
  OAI21_X1 U179 ( .B1(n490), .B2(n131), .A(n132), .ZN(n294) );
  NAND2_X1 U180 ( .A1(\mem[5][0] ), .A2(n462), .ZN(n132) );
  OAI21_X1 U181 ( .B1(n489), .B2(n131), .A(n133), .ZN(n295) );
  NAND2_X1 U182 ( .A1(\mem[5][1] ), .A2(n462), .ZN(n133) );
  OAI21_X1 U183 ( .B1(n488), .B2(n131), .A(n134), .ZN(n296) );
  NAND2_X1 U184 ( .A1(\mem[5][2] ), .A2(n462), .ZN(n134) );
  OAI21_X1 U185 ( .B1(n487), .B2(n131), .A(n135), .ZN(n297) );
  NAND2_X1 U186 ( .A1(\mem[5][3] ), .A2(n462), .ZN(n135) );
  OAI21_X1 U187 ( .B1(n486), .B2(n462), .A(n136), .ZN(n298) );
  NAND2_X1 U188 ( .A1(\mem[5][4] ), .A2(n462), .ZN(n136) );
  OAI21_X1 U189 ( .B1(n485), .B2(n131), .A(n137), .ZN(n299) );
  NAND2_X1 U190 ( .A1(\mem[5][5] ), .A2(n462), .ZN(n137) );
  OAI21_X1 U191 ( .B1(n484), .B2(n131), .A(n138), .ZN(n300) );
  NAND2_X1 U192 ( .A1(\mem[5][6] ), .A2(n462), .ZN(n138) );
  OAI21_X1 U193 ( .B1(n483), .B2(n131), .A(n139), .ZN(n301) );
  NAND2_X1 U194 ( .A1(\mem[5][7] ), .A2(n462), .ZN(n139) );
  OAI21_X1 U195 ( .B1(n482), .B2(n131), .A(n140), .ZN(n302) );
  NAND2_X1 U196 ( .A1(\mem[5][8] ), .A2(n462), .ZN(n140) );
  OAI21_X1 U197 ( .B1(n481), .B2(n131), .A(n141), .ZN(n303) );
  NAND2_X1 U198 ( .A1(\mem[5][9] ), .A2(n462), .ZN(n141) );
  OAI21_X1 U199 ( .B1(n480), .B2(n131), .A(n142), .ZN(n304) );
  NAND2_X1 U200 ( .A1(\mem[5][10] ), .A2(n462), .ZN(n142) );
  OAI21_X1 U201 ( .B1(n479), .B2(n131), .A(n143), .ZN(n305) );
  NAND2_X1 U202 ( .A1(\mem[5][11] ), .A2(n462), .ZN(n143) );
  OAI21_X1 U203 ( .B1(n478), .B2(n131), .A(n144), .ZN(n306) );
  NAND2_X1 U204 ( .A1(\mem[5][12] ), .A2(n131), .ZN(n144) );
  OAI21_X1 U205 ( .B1(n477), .B2(n462), .A(n145), .ZN(n307) );
  NAND2_X1 U206 ( .A1(\mem[5][13] ), .A2(n131), .ZN(n145) );
  OAI21_X1 U207 ( .B1(n476), .B2(n462), .A(n146), .ZN(n308) );
  NAND2_X1 U208 ( .A1(\mem[5][14] ), .A2(n131), .ZN(n146) );
  OAI21_X1 U209 ( .B1(n475), .B2(n131), .A(n147), .ZN(n309) );
  NAND2_X1 U210 ( .A1(\mem[5][15] ), .A2(n131), .ZN(n147) );
  OAI21_X1 U211 ( .B1(n474), .B2(n131), .A(n148), .ZN(n310) );
  NAND2_X1 U212 ( .A1(\mem[5][16] ), .A2(n131), .ZN(n148) );
  OAI21_X1 U213 ( .B1(n473), .B2(n131), .A(n149), .ZN(n311) );
  NAND2_X1 U214 ( .A1(\mem[5][17] ), .A2(n131), .ZN(n149) );
  OAI21_X1 U215 ( .B1(n472), .B2(n131), .A(n150), .ZN(n312) );
  NAND2_X1 U216 ( .A1(\mem[5][18] ), .A2(n131), .ZN(n150) );
  OAI21_X1 U217 ( .B1(n471), .B2(n131), .A(n151), .ZN(n313) );
  NAND2_X1 U218 ( .A1(\mem[5][19] ), .A2(n462), .ZN(n151) );
  OAI21_X1 U219 ( .B1(n490), .B2(n152), .A(n153), .ZN(n314) );
  NAND2_X1 U220 ( .A1(\mem[6][0] ), .A2(n461), .ZN(n153) );
  OAI21_X1 U221 ( .B1(n489), .B2(n152), .A(n154), .ZN(n315) );
  NAND2_X1 U222 ( .A1(\mem[6][1] ), .A2(n461), .ZN(n154) );
  OAI21_X1 U223 ( .B1(n488), .B2(n152), .A(n155), .ZN(n316) );
  NAND2_X1 U224 ( .A1(\mem[6][2] ), .A2(n461), .ZN(n155) );
  OAI21_X1 U225 ( .B1(n487), .B2(n152), .A(n156), .ZN(n317) );
  NAND2_X1 U226 ( .A1(\mem[6][3] ), .A2(n461), .ZN(n156) );
  OAI21_X1 U227 ( .B1(n486), .B2(n461), .A(n157), .ZN(n318) );
  NAND2_X1 U228 ( .A1(\mem[6][4] ), .A2(n461), .ZN(n157) );
  OAI21_X1 U229 ( .B1(n485), .B2(n152), .A(n158), .ZN(n319) );
  NAND2_X1 U230 ( .A1(\mem[6][5] ), .A2(n461), .ZN(n158) );
  OAI21_X1 U231 ( .B1(n484), .B2(n152), .A(n159), .ZN(n320) );
  NAND2_X1 U232 ( .A1(\mem[6][6] ), .A2(n461), .ZN(n159) );
  OAI21_X1 U233 ( .B1(n483), .B2(n152), .A(n160), .ZN(n321) );
  NAND2_X1 U234 ( .A1(\mem[6][7] ), .A2(n461), .ZN(n160) );
  OAI21_X1 U235 ( .B1(n482), .B2(n152), .A(n161), .ZN(n322) );
  NAND2_X1 U236 ( .A1(\mem[6][8] ), .A2(n461), .ZN(n161) );
  OAI21_X1 U237 ( .B1(n481), .B2(n152), .A(n162), .ZN(n323) );
  NAND2_X1 U238 ( .A1(\mem[6][9] ), .A2(n461), .ZN(n162) );
  OAI21_X1 U239 ( .B1(n480), .B2(n152), .A(n163), .ZN(n324) );
  NAND2_X1 U240 ( .A1(\mem[6][10] ), .A2(n461), .ZN(n163) );
  OAI21_X1 U241 ( .B1(n479), .B2(n152), .A(n164), .ZN(n325) );
  NAND2_X1 U242 ( .A1(\mem[6][11] ), .A2(n461), .ZN(n164) );
  OAI21_X1 U243 ( .B1(n478), .B2(n152), .A(n165), .ZN(n326) );
  NAND2_X1 U244 ( .A1(\mem[6][12] ), .A2(n152), .ZN(n165) );
  OAI21_X1 U245 ( .B1(n477), .B2(n461), .A(n166), .ZN(n327) );
  NAND2_X1 U246 ( .A1(\mem[6][13] ), .A2(n152), .ZN(n166) );
  OAI21_X1 U247 ( .B1(n476), .B2(n461), .A(n167), .ZN(n328) );
  NAND2_X1 U248 ( .A1(\mem[6][14] ), .A2(n152), .ZN(n167) );
  OAI21_X1 U249 ( .B1(n475), .B2(n152), .A(n168), .ZN(n329) );
  NAND2_X1 U250 ( .A1(\mem[6][15] ), .A2(n152), .ZN(n168) );
  OAI21_X1 U251 ( .B1(n474), .B2(n152), .A(n169), .ZN(n330) );
  NAND2_X1 U252 ( .A1(\mem[6][16] ), .A2(n152), .ZN(n169) );
  OAI21_X1 U253 ( .B1(n473), .B2(n152), .A(n170), .ZN(n331) );
  NAND2_X1 U254 ( .A1(\mem[6][17] ), .A2(n152), .ZN(n170) );
  OAI21_X1 U255 ( .B1(n472), .B2(n152), .A(n171), .ZN(n332) );
  NAND2_X1 U256 ( .A1(\mem[6][18] ), .A2(n152), .ZN(n171) );
  OAI21_X1 U257 ( .B1(n471), .B2(n152), .A(n172), .ZN(n333) );
  NAND2_X1 U258 ( .A1(\mem[6][19] ), .A2(n461), .ZN(n172) );
  OAI21_X1 U259 ( .B1(n490), .B2(n460), .A(n174), .ZN(n334) );
  NAND2_X1 U260 ( .A1(\mem[7][0] ), .A2(n460), .ZN(n174) );
  OAI21_X1 U261 ( .B1(n489), .B2(n460), .A(n175), .ZN(n335) );
  NAND2_X1 U262 ( .A1(\mem[7][1] ), .A2(n460), .ZN(n175) );
  OAI21_X1 U263 ( .B1(n488), .B2(n460), .A(n176), .ZN(n336) );
  NAND2_X1 U264 ( .A1(\mem[7][2] ), .A2(n173), .ZN(n176) );
  OAI21_X1 U265 ( .B1(n487), .B2(n173), .A(n177), .ZN(n337) );
  NAND2_X1 U266 ( .A1(\mem[7][3] ), .A2(n460), .ZN(n177) );
  OAI21_X1 U267 ( .B1(n486), .B2(n173), .A(n178), .ZN(n338) );
  NAND2_X1 U268 ( .A1(\mem[7][4] ), .A2(n173), .ZN(n178) );
  OAI21_X1 U269 ( .B1(n485), .B2(n173), .A(n179), .ZN(n339) );
  NAND2_X1 U270 ( .A1(\mem[7][5] ), .A2(n173), .ZN(n179) );
  OAI21_X1 U271 ( .B1(n484), .B2(n173), .A(n180), .ZN(n340) );
  NAND2_X1 U272 ( .A1(\mem[7][6] ), .A2(n173), .ZN(n180) );
  OAI21_X1 U273 ( .B1(n483), .B2(n173), .A(n181), .ZN(n341) );
  NAND2_X1 U274 ( .A1(\mem[7][7] ), .A2(n173), .ZN(n181) );
  OAI21_X1 U275 ( .B1(n482), .B2(n173), .A(n182), .ZN(n342) );
  NAND2_X1 U276 ( .A1(\mem[7][8] ), .A2(n173), .ZN(n182) );
  OAI21_X1 U277 ( .B1(n481), .B2(n460), .A(n183), .ZN(n343) );
  NAND2_X1 U278 ( .A1(\mem[7][9] ), .A2(n173), .ZN(n183) );
  OAI21_X1 U279 ( .B1(n480), .B2(n173), .A(n184), .ZN(n344) );
  NAND2_X1 U280 ( .A1(\mem[7][10] ), .A2(n173), .ZN(n184) );
  OAI21_X1 U281 ( .B1(n479), .B2(n173), .A(n185), .ZN(n345) );
  NAND2_X1 U282 ( .A1(\mem[7][11] ), .A2(n173), .ZN(n185) );
  OAI21_X1 U283 ( .B1(n478), .B2(n460), .A(n186), .ZN(n346) );
  NAND2_X1 U284 ( .A1(\mem[7][12] ), .A2(n460), .ZN(n186) );
  OAI21_X1 U285 ( .B1(n477), .B2(n460), .A(n187), .ZN(n347) );
  NAND2_X1 U286 ( .A1(\mem[7][13] ), .A2(n460), .ZN(n187) );
  OAI21_X1 U287 ( .B1(n476), .B2(n460), .A(n188), .ZN(n348) );
  NAND2_X1 U288 ( .A1(\mem[7][14] ), .A2(n460), .ZN(n188) );
  OAI21_X1 U289 ( .B1(n475), .B2(n173), .A(n189), .ZN(n349) );
  NAND2_X1 U290 ( .A1(\mem[7][15] ), .A2(n460), .ZN(n189) );
  OAI21_X1 U291 ( .B1(n474), .B2(n173), .A(n190), .ZN(n350) );
  NAND2_X1 U292 ( .A1(\mem[7][16] ), .A2(n460), .ZN(n190) );
  OAI21_X1 U293 ( .B1(n473), .B2(n173), .A(n191), .ZN(n351) );
  NAND2_X1 U294 ( .A1(\mem[7][17] ), .A2(n460), .ZN(n191) );
  OAI21_X1 U295 ( .B1(n472), .B2(n460), .A(n192), .ZN(n352) );
  NAND2_X1 U296 ( .A1(\mem[7][18] ), .A2(n460), .ZN(n192) );
  OAI21_X1 U297 ( .B1(n471), .B2(n460), .A(n193), .ZN(n353) );
  NAND2_X1 U298 ( .A1(\mem[7][19] ), .A2(n460), .ZN(n193) );
  OAI21_X1 U299 ( .B1(n24), .B2(n488), .A(n27), .ZN(n196) );
  NAND2_X1 U300 ( .A1(\mem[0][2] ), .A2(n467), .ZN(n27) );
  OAI21_X1 U301 ( .B1(n24), .B2(n487), .A(n28), .ZN(n197) );
  NAND2_X1 U302 ( .A1(\mem[0][3] ), .A2(n467), .ZN(n28) );
  OAI21_X1 U303 ( .B1(n24), .B2(n486), .A(n29), .ZN(n198) );
  NAND2_X1 U304 ( .A1(\mem[0][4] ), .A2(n467), .ZN(n29) );
  OAI21_X1 U305 ( .B1(n24), .B2(n485), .A(n30), .ZN(n199) );
  NAND2_X1 U306 ( .A1(\mem[0][5] ), .A2(n467), .ZN(n30) );
  OAI21_X1 U307 ( .B1(n24), .B2(n484), .A(n31), .ZN(n200) );
  NAND2_X1 U308 ( .A1(\mem[0][6] ), .A2(n467), .ZN(n31) );
  OAI21_X1 U309 ( .B1(n24), .B2(n483), .A(n32), .ZN(n201) );
  NAND2_X1 U310 ( .A1(\mem[0][7] ), .A2(n467), .ZN(n32) );
  OAI21_X1 U311 ( .B1(n24), .B2(n482), .A(n33), .ZN(n202) );
  NAND2_X1 U312 ( .A1(\mem[0][8] ), .A2(n467), .ZN(n33) );
  OAI21_X1 U313 ( .B1(n24), .B2(n481), .A(n34), .ZN(n203) );
  NAND2_X1 U314 ( .A1(\mem[0][9] ), .A2(n467), .ZN(n34) );
  OAI21_X1 U315 ( .B1(n24), .B2(n480), .A(n35), .ZN(n204) );
  NAND2_X1 U316 ( .A1(\mem[0][10] ), .A2(n467), .ZN(n35) );
  OAI21_X1 U317 ( .B1(n24), .B2(n479), .A(n36), .ZN(n205) );
  NAND2_X1 U318 ( .A1(\mem[0][11] ), .A2(n467), .ZN(n36) );
  OAI21_X1 U319 ( .B1(n24), .B2(n478), .A(n37), .ZN(n206) );
  NAND2_X1 U320 ( .A1(\mem[0][12] ), .A2(n24), .ZN(n37) );
  OAI21_X1 U321 ( .B1(n24), .B2(n477), .A(n38), .ZN(n207) );
  NAND2_X1 U322 ( .A1(\mem[0][13] ), .A2(n24), .ZN(n38) );
  OAI21_X1 U323 ( .B1(n467), .B2(n476), .A(n39), .ZN(n208) );
  NAND2_X1 U324 ( .A1(\mem[0][14] ), .A2(n24), .ZN(n39) );
  OAI21_X1 U325 ( .B1(n24), .B2(n475), .A(n40), .ZN(n209) );
  NAND2_X1 U326 ( .A1(\mem[0][15] ), .A2(n467), .ZN(n40) );
  OAI21_X1 U327 ( .B1(n24), .B2(n474), .A(n41), .ZN(n210) );
  NAND2_X1 U328 ( .A1(\mem[0][16] ), .A2(n24), .ZN(n41) );
  OAI21_X1 U329 ( .B1(n24), .B2(n473), .A(n42), .ZN(n211) );
  NAND2_X1 U330 ( .A1(\mem[0][17] ), .A2(n24), .ZN(n42) );
  OAI21_X1 U331 ( .B1(n24), .B2(n472), .A(n43), .ZN(n212) );
  NAND2_X1 U332 ( .A1(\mem[0][18] ), .A2(n24), .ZN(n43) );
  OAI21_X1 U333 ( .B1(n467), .B2(n490), .A(n25), .ZN(n194) );
  NAND2_X1 U334 ( .A1(\mem[0][0] ), .A2(n467), .ZN(n25) );
  OAI21_X1 U335 ( .B1(n24), .B2(n489), .A(n26), .ZN(n195) );
  NAND2_X1 U336 ( .A1(\mem[0][1] ), .A2(n467), .ZN(n26) );
  OAI21_X1 U337 ( .B1(n24), .B2(n471), .A(n44), .ZN(n213) );
  NAND2_X1 U338 ( .A1(\mem[0][19] ), .A2(n467), .ZN(n44) );
  INV_X1 U339 ( .A(N10), .ZN(n468) );
  INV_X1 U340 ( .A(N11), .ZN(n469) );
  INV_X1 U341 ( .A(data_in[0]), .ZN(n490) );
  INV_X1 U342 ( .A(data_in[1]), .ZN(n489) );
  INV_X1 U343 ( .A(data_in[2]), .ZN(n488) );
  INV_X1 U344 ( .A(data_in[3]), .ZN(n487) );
  INV_X1 U345 ( .A(data_in[4]), .ZN(n486) );
  INV_X1 U346 ( .A(data_in[5]), .ZN(n485) );
  INV_X1 U347 ( .A(data_in[6]), .ZN(n484) );
  INV_X1 U356 ( .A(data_in[7]), .ZN(n483) );
  INV_X1 U357 ( .A(data_in[8]), .ZN(n482) );
  INV_X1 U358 ( .A(data_in[9]), .ZN(n481) );
  INV_X1 U359 ( .A(data_in[10]), .ZN(n480) );
  INV_X1 U360 ( .A(data_in[11]), .ZN(n479) );
  INV_X1 U361 ( .A(data_in[12]), .ZN(n478) );
  INV_X1 U362 ( .A(data_in[13]), .ZN(n477) );
  INV_X1 U363 ( .A(data_in[14]), .ZN(n476) );
  INV_X1 U364 ( .A(data_in[15]), .ZN(n475) );
  INV_X1 U365 ( .A(data_in[16]), .ZN(n474) );
  INV_X1 U366 ( .A(data_in[17]), .ZN(n473) );
  INV_X1 U367 ( .A(data_in[18]), .ZN(n472) );
  INV_X1 U368 ( .A(data_in[19]), .ZN(n471) );
  MUX2_X1 U369 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n457), .Z(n5) );
  MUX2_X1 U370 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n459), .Z(n6) );
  MUX2_X1 U371 ( .A(n6), .B(n5), .S(n456), .Z(n7) );
  MUX2_X1 U372 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n459), .Z(n8) );
  MUX2_X1 U373 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n457), .Z(n9) );
  MUX2_X1 U374 ( .A(n9), .B(n8), .S(n456), .Z(n10) );
  MUX2_X1 U375 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n458), .Z(n11) );
  MUX2_X1 U376 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n458), .Z(n12) );
  MUX2_X1 U377 ( .A(n12), .B(n11), .S(n456), .Z(n13) );
  MUX2_X1 U378 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n457), .Z(n14) );
  MUX2_X1 U379 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n458), .Z(n15) );
  MUX2_X1 U380 ( .A(n15), .B(n14), .S(n456), .Z(n16) );
  MUX2_X1 U381 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n459), .Z(n17) );
  MUX2_X1 U382 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n459), .Z(n18) );
  MUX2_X1 U383 ( .A(n18), .B(n17), .S(n456), .Z(n19) );
  MUX2_X1 U384 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n458), .Z(n20) );
  MUX2_X1 U385 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n458), .Z(n21) );
  MUX2_X1 U386 ( .A(n21), .B(n20), .S(n455), .Z(n22) );
  MUX2_X1 U387 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n457), .Z(n23) );
  MUX2_X1 U388 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n354) );
  MUX2_X1 U389 ( .A(n354), .B(n23), .S(n456), .Z(n355) );
  MUX2_X1 U390 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n459), .Z(n356) );
  MUX2_X1 U391 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n457), .Z(n357) );
  MUX2_X1 U392 ( .A(n357), .B(n356), .S(n455), .Z(n358) );
  MUX2_X1 U393 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n458), .Z(n359) );
  MUX2_X1 U394 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n458), .Z(n360) );
  MUX2_X1 U395 ( .A(n360), .B(n359), .S(n456), .Z(n361) );
  MUX2_X1 U396 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(N10), .Z(n362) );
  MUX2_X1 U397 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n458), .Z(n363) );
  MUX2_X1 U398 ( .A(n363), .B(n362), .S(n455), .Z(n364) );
  MUX2_X1 U399 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n457), .Z(n365) );
  MUX2_X1 U400 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n457), .Z(n366) );
  MUX2_X1 U401 ( .A(n366), .B(n365), .S(n456), .Z(n367) );
  MUX2_X1 U402 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n457), .Z(n368) );
  MUX2_X1 U403 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n457), .Z(n369) );
  MUX2_X1 U404 ( .A(n369), .B(n368), .S(n455), .Z(n370) );
  MUX2_X1 U405 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n457), .Z(n371) );
  MUX2_X1 U406 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n457), .Z(n372) );
  MUX2_X1 U407 ( .A(n372), .B(n371), .S(n456), .Z(n373) );
  MUX2_X1 U408 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n457), .Z(n374) );
  MUX2_X1 U409 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n457), .Z(n375) );
  MUX2_X1 U410 ( .A(n375), .B(n374), .S(N11), .Z(n376) );
  MUX2_X1 U411 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n457), .Z(n377) );
  MUX2_X1 U412 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n457), .Z(n378) );
  MUX2_X1 U413 ( .A(n378), .B(n377), .S(n456), .Z(n379) );
  MUX2_X1 U414 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n457), .Z(n380) );
  MUX2_X1 U415 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n457), .Z(n381) );
  MUX2_X1 U416 ( .A(n381), .B(n380), .S(N11), .Z(n382) );
  MUX2_X1 U417 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n458), .Z(n383) );
  MUX2_X1 U418 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n458), .Z(n384) );
  MUX2_X1 U419 ( .A(n384), .B(n383), .S(n456), .Z(n385) );
  MUX2_X1 U420 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n458), .Z(n386) );
  MUX2_X1 U421 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n458), .Z(n387) );
  MUX2_X1 U422 ( .A(n387), .B(n386), .S(n456), .Z(n388) );
  MUX2_X1 U423 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n458), .Z(n389) );
  MUX2_X1 U424 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n458), .Z(n390) );
  MUX2_X1 U425 ( .A(n390), .B(n389), .S(n456), .Z(n391) );
  MUX2_X1 U426 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n458), .Z(n392) );
  MUX2_X1 U427 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n458), .Z(n393) );
  MUX2_X1 U428 ( .A(n393), .B(n392), .S(n456), .Z(n394) );
  MUX2_X1 U429 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n458), .Z(n395) );
  MUX2_X1 U430 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n458), .Z(n396) );
  MUX2_X1 U431 ( .A(n396), .B(n395), .S(n456), .Z(n397) );
  MUX2_X1 U432 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n458), .Z(n398) );
  MUX2_X1 U433 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n458), .Z(n399) );
  MUX2_X1 U434 ( .A(n399), .B(n398), .S(n456), .Z(n400) );
  MUX2_X1 U435 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n459), .Z(n401) );
  MUX2_X1 U436 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n459), .Z(n402) );
  MUX2_X1 U437 ( .A(n402), .B(n401), .S(n456), .Z(n403) );
  MUX2_X1 U438 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n459), .Z(n404) );
  MUX2_X1 U439 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n459), .Z(n405) );
  MUX2_X1 U440 ( .A(n405), .B(n404), .S(n456), .Z(n406) );
  MUX2_X1 U441 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n459), .Z(n407) );
  MUX2_X1 U442 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n459), .Z(n408) );
  MUX2_X1 U443 ( .A(n408), .B(n407), .S(n456), .Z(n409) );
  MUX2_X1 U444 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n459), .Z(n410) );
  MUX2_X1 U445 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n459), .Z(n411) );
  MUX2_X1 U446 ( .A(n411), .B(n410), .S(n456), .Z(n412) );
  MUX2_X1 U447 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n459), .Z(n413) );
  MUX2_X1 U448 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n459), .Z(n414) );
  MUX2_X1 U449 ( .A(n414), .B(n413), .S(n456), .Z(n415) );
  MUX2_X1 U450 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n459), .Z(n416) );
  MUX2_X1 U451 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n459), .Z(n417) );
  MUX2_X1 U452 ( .A(n417), .B(n416), .S(n456), .Z(n418) );
  MUX2_X1 U453 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n459), .Z(n419) );
  MUX2_X1 U454 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n459), .Z(n420) );
  MUX2_X1 U455 ( .A(n420), .B(n419), .S(n455), .Z(n421) );
  MUX2_X1 U456 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(N10), .Z(n422) );
  MUX2_X1 U457 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(N10), .Z(n423) );
  MUX2_X1 U458 ( .A(n423), .B(n422), .S(n455), .Z(n424) );
  MUX2_X1 U459 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n457), .Z(n425) );
  MUX2_X1 U460 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n457), .Z(n426) );
  MUX2_X1 U461 ( .A(n426), .B(n425), .S(n455), .Z(n427) );
  MUX2_X1 U462 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(N10), .Z(n428) );
  MUX2_X1 U463 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(N10), .Z(n429) );
  MUX2_X1 U464 ( .A(n429), .B(n428), .S(n455), .Z(n430) );
  MUX2_X1 U465 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n458), .Z(n431) );
  MUX2_X1 U466 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n458), .Z(n432) );
  MUX2_X1 U467 ( .A(n432), .B(n431), .S(n455), .Z(n433) );
  MUX2_X1 U468 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(N10), .Z(n434) );
  MUX2_X1 U469 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(N10), .Z(n435) );
  MUX2_X1 U470 ( .A(n435), .B(n434), .S(n455), .Z(n436) );
  MUX2_X1 U471 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n459), .Z(n437) );
  MUX2_X1 U472 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n459), .Z(n438) );
  MUX2_X1 U473 ( .A(n438), .B(n437), .S(n455), .Z(n439) );
  MUX2_X1 U474 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(N10), .Z(n440) );
  MUX2_X1 U475 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n459), .Z(n441) );
  MUX2_X1 U476 ( .A(n441), .B(n440), .S(n455), .Z(n442) );
  MUX2_X1 U477 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n459), .Z(n443) );
  MUX2_X1 U478 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(N10), .Z(n444) );
  MUX2_X1 U479 ( .A(n444), .B(n443), .S(n455), .Z(n445) );
  MUX2_X1 U480 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n457), .Z(n446) );
  MUX2_X1 U481 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(N10), .Z(n447) );
  MUX2_X1 U482 ( .A(n447), .B(n446), .S(n455), .Z(n448) );
  MUX2_X1 U483 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n457), .Z(n449) );
  MUX2_X1 U484 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n457), .Z(n450) );
  MUX2_X1 U485 ( .A(n450), .B(n449), .S(n455), .Z(n451) );
  MUX2_X1 U486 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n458), .Z(n452) );
  MUX2_X1 U487 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n457), .Z(n453) );
  MUX2_X1 U488 ( .A(n453), .B(n452), .S(n455), .Z(n454) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE3_8 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N15, N16, N18, N20, N22, N23, N26, N30, N32, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[16]  ( .D(N16), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N20), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N22), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N23), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[6]  ( .D(N26), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[2]  ( .D(N30), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N32), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n486), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n487), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n488), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n489), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n490), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n491), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n492), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n493), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n494), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n495), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n496), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n497), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n498), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n499), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n500), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n501), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n502), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n503), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n504), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n505), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n506), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n507), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n508), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n509), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n510), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n511), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n512), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n513), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n514), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n515), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n516), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n517), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n518), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n519), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n520), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n521), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n522), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n523), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n524), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n525), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n526), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n527), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n528), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n529), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n530), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n531), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n532), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n533), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n534), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n535), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n536), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n537), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n538), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n539), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n540), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n541), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n542), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n543), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n544), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n545), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n546), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n547), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n548), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n549), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n550), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n551), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n552), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n553), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n554), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n555), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n556), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n557), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n558), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n559), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n560), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n561), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n562), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n563), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n564), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n565), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n566), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n567), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n568), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n569), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n570), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n571), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n572), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n573), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n574), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n575), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n576), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n577), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n578), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n579), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n580), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n581), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n582), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n583), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n584), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n585), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n586), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n587), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n588), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n589), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n590), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n591), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n592), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n593), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n594), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n595), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n596), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n597), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n598), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n599), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n600), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n601), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n602), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n603), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n604), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n605), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n606), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n607), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n608), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n609), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n610), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n611), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n612), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n613), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n614), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n615), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n616), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n617), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n618), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n619), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n620), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n621), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n622), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n623), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n624), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n625), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n626), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n627), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n628), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n629), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n630), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n631), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n632), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n633), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n634), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n635), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n636), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n637), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n638), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n639), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n640), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n641), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n642), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n643), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n644), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n645), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U348 ( .A1(n463), .A2(n464), .A3(n794), .ZN(n815) );
  NAND3_X1 U349 ( .A1(n794), .A2(n464), .A3(N10), .ZN(n793) );
  NAND3_X1 U350 ( .A1(n794), .A2(n463), .A3(N11), .ZN(n772) );
  NAND3_X1 U351 ( .A1(N10), .A2(n794), .A3(N11), .ZN(n751) );
  NAND3_X1 U352 ( .A1(n463), .A2(n464), .A3(n709), .ZN(n730) );
  NAND3_X1 U353 ( .A1(N10), .A2(n464), .A3(n709), .ZN(n708) );
  NAND3_X1 U354 ( .A1(N11), .A2(n463), .A3(n709), .ZN(n687) );
  NAND3_X1 U355 ( .A1(N11), .A2(N10), .A3(n709), .ZN(n666) );
  DFF_X1 \data_out_reg[17]  ( .D(N15), .CK(clk), .Q(data_out[17]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n402), .SI(n399), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n366), .SI(n363), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n354), .SI(n21), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[19]  ( .D(n450), .SI(n447), .SE(N12), .CK(clk), .Q(
        data_out[19]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n12), .SI(n9), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n414), .SI(n411), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n378), .SI(n375), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n426), .SI(n423), .SE(N12), .CK(clk), .Q(
        data_out[15]) );
  SDFF_X1 \data_out_reg[18]  ( .D(n444), .SI(n441), .SE(N12), .CK(clk), .Q(
        data_out[18]) );
  SDFF_X1 \data_out_reg[8]  ( .D(n384), .SI(n381), .SE(N12), .CK(clk), .Q(
        data_out[8]) );
  SDFF_X1 \data_out_reg[4]  ( .D(n360), .SI(n357), .SE(N12), .CK(clk), .Q(
        data_out[4]) );
  BUF_X1 U3 ( .A(n815), .Z(n462) );
  BUF_X1 U4 ( .A(n793), .Z(n461) );
  BUF_X1 U5 ( .A(n751), .Z(n459) );
  BUF_X1 U6 ( .A(n666), .Z(n455) );
  BUF_X1 U7 ( .A(n772), .Z(n460) );
  BUF_X1 U8 ( .A(n730), .Z(n458) );
  BUF_X1 U9 ( .A(n708), .Z(n457) );
  BUF_X1 U10 ( .A(n687), .Z(n456) );
  BUF_X1 U11 ( .A(N10), .Z(n453) );
  BUF_X1 U12 ( .A(N10), .Z(n454) );
  BUF_X1 U13 ( .A(N11), .Z(n451) );
  NOR2_X1 U14 ( .A1(n465), .A2(N12), .ZN(n794) );
  INV_X1 U15 ( .A(wr_en), .ZN(n465) );
  AND2_X1 U16 ( .A1(N12), .A2(wr_en), .ZN(n709) );
  OAI21_X1 U17 ( .B1(n485), .B2(n461), .A(n792), .ZN(n625) );
  NAND2_X1 U18 ( .A1(\mem[1][0] ), .A2(n461), .ZN(n792) );
  OAI21_X1 U19 ( .B1(n484), .B2(n461), .A(n791), .ZN(n624) );
  NAND2_X1 U20 ( .A1(\mem[1][1] ), .A2(n461), .ZN(n791) );
  OAI21_X1 U21 ( .B1(n483), .B2(n461), .A(n790), .ZN(n623) );
  NAND2_X1 U22 ( .A1(\mem[1][2] ), .A2(n793), .ZN(n790) );
  OAI21_X1 U23 ( .B1(n482), .B2(n793), .A(n789), .ZN(n622) );
  NAND2_X1 U24 ( .A1(\mem[1][3] ), .A2(n461), .ZN(n789) );
  OAI21_X1 U25 ( .B1(n481), .B2(n793), .A(n788), .ZN(n621) );
  NAND2_X1 U26 ( .A1(\mem[1][4] ), .A2(n461), .ZN(n788) );
  OAI21_X1 U27 ( .B1(n480), .B2(n793), .A(n787), .ZN(n620) );
  NAND2_X1 U28 ( .A1(\mem[1][5] ), .A2(n793), .ZN(n787) );
  OAI21_X1 U29 ( .B1(n479), .B2(n793), .A(n786), .ZN(n619) );
  NAND2_X1 U30 ( .A1(\mem[1][6] ), .A2(n793), .ZN(n786) );
  OAI21_X1 U31 ( .B1(n478), .B2(n793), .A(n785), .ZN(n618) );
  NAND2_X1 U32 ( .A1(\mem[1][7] ), .A2(n793), .ZN(n785) );
  OAI21_X1 U33 ( .B1(n477), .B2(n793), .A(n784), .ZN(n617) );
  NAND2_X1 U34 ( .A1(\mem[1][8] ), .A2(n793), .ZN(n784) );
  OAI21_X1 U35 ( .B1(n476), .B2(n461), .A(n783), .ZN(n616) );
  NAND2_X1 U36 ( .A1(\mem[1][9] ), .A2(n793), .ZN(n783) );
  OAI21_X1 U37 ( .B1(n475), .B2(n793), .A(n782), .ZN(n615) );
  NAND2_X1 U38 ( .A1(\mem[1][10] ), .A2(n793), .ZN(n782) );
  OAI21_X1 U39 ( .B1(n474), .B2(n793), .A(n781), .ZN(n614) );
  NAND2_X1 U40 ( .A1(\mem[1][11] ), .A2(n793), .ZN(n781) );
  OAI21_X1 U41 ( .B1(n473), .B2(n461), .A(n780), .ZN(n613) );
  NAND2_X1 U42 ( .A1(\mem[1][12] ), .A2(n461), .ZN(n780) );
  OAI21_X1 U43 ( .B1(n472), .B2(n461), .A(n779), .ZN(n612) );
  NAND2_X1 U44 ( .A1(\mem[1][13] ), .A2(n461), .ZN(n779) );
  OAI21_X1 U45 ( .B1(n471), .B2(n461), .A(n778), .ZN(n611) );
  NAND2_X1 U46 ( .A1(\mem[1][14] ), .A2(n461), .ZN(n778) );
  OAI21_X1 U47 ( .B1(n470), .B2(n793), .A(n777), .ZN(n610) );
  NAND2_X1 U48 ( .A1(\mem[1][15] ), .A2(n461), .ZN(n777) );
  OAI21_X1 U49 ( .B1(n469), .B2(n793), .A(n776), .ZN(n609) );
  NAND2_X1 U50 ( .A1(\mem[1][16] ), .A2(n461), .ZN(n776) );
  OAI21_X1 U51 ( .B1(n468), .B2(n793), .A(n775), .ZN(n608) );
  NAND2_X1 U52 ( .A1(\mem[1][17] ), .A2(n461), .ZN(n775) );
  OAI21_X1 U53 ( .B1(n467), .B2(n461), .A(n774), .ZN(n607) );
  NAND2_X1 U54 ( .A1(\mem[1][18] ), .A2(n461), .ZN(n774) );
  OAI21_X1 U55 ( .B1(n466), .B2(n461), .A(n773), .ZN(n606) );
  NAND2_X1 U56 ( .A1(\mem[1][19] ), .A2(n461), .ZN(n773) );
  OAI21_X1 U57 ( .B1(n485), .B2(n772), .A(n771), .ZN(n605) );
  NAND2_X1 U58 ( .A1(\mem[2][0] ), .A2(n460), .ZN(n771) );
  OAI21_X1 U59 ( .B1(n484), .B2(n772), .A(n770), .ZN(n604) );
  NAND2_X1 U60 ( .A1(\mem[2][1] ), .A2(n460), .ZN(n770) );
  OAI21_X1 U61 ( .B1(n483), .B2(n772), .A(n769), .ZN(n603) );
  NAND2_X1 U62 ( .A1(\mem[2][2] ), .A2(n460), .ZN(n769) );
  OAI21_X1 U63 ( .B1(n482), .B2(n772), .A(n768), .ZN(n602) );
  NAND2_X1 U64 ( .A1(\mem[2][3] ), .A2(n460), .ZN(n768) );
  OAI21_X1 U65 ( .B1(n481), .B2(n460), .A(n767), .ZN(n601) );
  NAND2_X1 U66 ( .A1(\mem[2][4] ), .A2(n460), .ZN(n767) );
  OAI21_X1 U67 ( .B1(n480), .B2(n460), .A(n766), .ZN(n600) );
  NAND2_X1 U68 ( .A1(\mem[2][5] ), .A2(n460), .ZN(n766) );
  OAI21_X1 U69 ( .B1(n479), .B2(n772), .A(n765), .ZN(n599) );
  NAND2_X1 U70 ( .A1(\mem[2][6] ), .A2(n460), .ZN(n765) );
  OAI21_X1 U71 ( .B1(n478), .B2(n772), .A(n764), .ZN(n598) );
  NAND2_X1 U72 ( .A1(\mem[2][7] ), .A2(n460), .ZN(n764) );
  OAI21_X1 U73 ( .B1(n477), .B2(n772), .A(n763), .ZN(n597) );
  NAND2_X1 U74 ( .A1(\mem[2][8] ), .A2(n460), .ZN(n763) );
  OAI21_X1 U75 ( .B1(n476), .B2(n772), .A(n762), .ZN(n596) );
  NAND2_X1 U76 ( .A1(\mem[2][9] ), .A2(n460), .ZN(n762) );
  OAI21_X1 U77 ( .B1(n475), .B2(n772), .A(n761), .ZN(n595) );
  NAND2_X1 U78 ( .A1(\mem[2][10] ), .A2(n460), .ZN(n761) );
  OAI21_X1 U79 ( .B1(n474), .B2(n772), .A(n760), .ZN(n594) );
  NAND2_X1 U80 ( .A1(\mem[2][11] ), .A2(n460), .ZN(n760) );
  OAI21_X1 U81 ( .B1(n473), .B2(n772), .A(n759), .ZN(n593) );
  NAND2_X1 U82 ( .A1(\mem[2][12] ), .A2(n772), .ZN(n759) );
  OAI21_X1 U83 ( .B1(n472), .B2(n772), .A(n758), .ZN(n592) );
  NAND2_X1 U84 ( .A1(\mem[2][13] ), .A2(n772), .ZN(n758) );
  OAI21_X1 U85 ( .B1(n471), .B2(n772), .A(n757), .ZN(n591) );
  NAND2_X1 U86 ( .A1(\mem[2][14] ), .A2(n772), .ZN(n757) );
  OAI21_X1 U87 ( .B1(n470), .B2(n772), .A(n756), .ZN(n590) );
  NAND2_X1 U88 ( .A1(\mem[2][15] ), .A2(n460), .ZN(n756) );
  OAI21_X1 U89 ( .B1(n469), .B2(n772), .A(n755), .ZN(n589) );
  NAND2_X1 U90 ( .A1(\mem[2][16] ), .A2(n772), .ZN(n755) );
  OAI21_X1 U91 ( .B1(n468), .B2(n772), .A(n754), .ZN(n588) );
  NAND2_X1 U92 ( .A1(\mem[2][17] ), .A2(n772), .ZN(n754) );
  OAI21_X1 U93 ( .B1(n467), .B2(n772), .A(n753), .ZN(n587) );
  NAND2_X1 U94 ( .A1(\mem[2][18] ), .A2(n772), .ZN(n753) );
  OAI21_X1 U95 ( .B1(n466), .B2(n772), .A(n752), .ZN(n586) );
  NAND2_X1 U96 ( .A1(\mem[2][19] ), .A2(n460), .ZN(n752) );
  OAI21_X1 U97 ( .B1(n485), .B2(n459), .A(n750), .ZN(n585) );
  NAND2_X1 U98 ( .A1(\mem[3][0] ), .A2(n459), .ZN(n750) );
  OAI21_X1 U99 ( .B1(n484), .B2(n459), .A(n749), .ZN(n584) );
  NAND2_X1 U100 ( .A1(\mem[3][1] ), .A2(n459), .ZN(n749) );
  OAI21_X1 U101 ( .B1(n483), .B2(n459), .A(n748), .ZN(n583) );
  NAND2_X1 U102 ( .A1(\mem[3][2] ), .A2(n751), .ZN(n748) );
  OAI21_X1 U103 ( .B1(n482), .B2(n751), .A(n747), .ZN(n582) );
  NAND2_X1 U104 ( .A1(\mem[3][3] ), .A2(n459), .ZN(n747) );
  OAI21_X1 U105 ( .B1(n481), .B2(n751), .A(n746), .ZN(n581) );
  NAND2_X1 U106 ( .A1(\mem[3][4] ), .A2(n459), .ZN(n746) );
  OAI21_X1 U107 ( .B1(n480), .B2(n751), .A(n745), .ZN(n580) );
  NAND2_X1 U108 ( .A1(\mem[3][5] ), .A2(n751), .ZN(n745) );
  OAI21_X1 U109 ( .B1(n479), .B2(n751), .A(n744), .ZN(n579) );
  NAND2_X1 U110 ( .A1(\mem[3][6] ), .A2(n751), .ZN(n744) );
  OAI21_X1 U111 ( .B1(n478), .B2(n751), .A(n743), .ZN(n578) );
  NAND2_X1 U112 ( .A1(\mem[3][7] ), .A2(n751), .ZN(n743) );
  OAI21_X1 U113 ( .B1(n477), .B2(n751), .A(n742), .ZN(n577) );
  NAND2_X1 U114 ( .A1(\mem[3][8] ), .A2(n751), .ZN(n742) );
  OAI21_X1 U115 ( .B1(n476), .B2(n459), .A(n741), .ZN(n576) );
  NAND2_X1 U116 ( .A1(\mem[3][9] ), .A2(n751), .ZN(n741) );
  OAI21_X1 U117 ( .B1(n475), .B2(n751), .A(n740), .ZN(n575) );
  NAND2_X1 U118 ( .A1(\mem[3][10] ), .A2(n751), .ZN(n740) );
  OAI21_X1 U119 ( .B1(n474), .B2(n751), .A(n739), .ZN(n574) );
  NAND2_X1 U120 ( .A1(\mem[3][11] ), .A2(n751), .ZN(n739) );
  OAI21_X1 U121 ( .B1(n473), .B2(n459), .A(n738), .ZN(n573) );
  NAND2_X1 U122 ( .A1(\mem[3][12] ), .A2(n459), .ZN(n738) );
  OAI21_X1 U123 ( .B1(n472), .B2(n459), .A(n737), .ZN(n572) );
  NAND2_X1 U124 ( .A1(\mem[3][13] ), .A2(n459), .ZN(n737) );
  OAI21_X1 U125 ( .B1(n471), .B2(n459), .A(n736), .ZN(n571) );
  NAND2_X1 U126 ( .A1(\mem[3][14] ), .A2(n459), .ZN(n736) );
  OAI21_X1 U127 ( .B1(n470), .B2(n751), .A(n735), .ZN(n570) );
  NAND2_X1 U128 ( .A1(\mem[3][15] ), .A2(n459), .ZN(n735) );
  OAI21_X1 U129 ( .B1(n469), .B2(n751), .A(n734), .ZN(n569) );
  NAND2_X1 U130 ( .A1(\mem[3][16] ), .A2(n459), .ZN(n734) );
  OAI21_X1 U131 ( .B1(n468), .B2(n751), .A(n733), .ZN(n568) );
  NAND2_X1 U132 ( .A1(\mem[3][17] ), .A2(n459), .ZN(n733) );
  OAI21_X1 U133 ( .B1(n467), .B2(n459), .A(n732), .ZN(n567) );
  NAND2_X1 U134 ( .A1(\mem[3][18] ), .A2(n459), .ZN(n732) );
  OAI21_X1 U135 ( .B1(n466), .B2(n459), .A(n731), .ZN(n566) );
  NAND2_X1 U136 ( .A1(\mem[3][19] ), .A2(n459), .ZN(n731) );
  OAI21_X1 U137 ( .B1(n485), .B2(n730), .A(n729), .ZN(n565) );
  NAND2_X1 U138 ( .A1(\mem[4][0] ), .A2(n458), .ZN(n729) );
  OAI21_X1 U139 ( .B1(n484), .B2(n730), .A(n728), .ZN(n564) );
  NAND2_X1 U140 ( .A1(\mem[4][1] ), .A2(n458), .ZN(n728) );
  OAI21_X1 U141 ( .B1(n483), .B2(n730), .A(n727), .ZN(n563) );
  NAND2_X1 U142 ( .A1(\mem[4][2] ), .A2(n458), .ZN(n727) );
  OAI21_X1 U143 ( .B1(n482), .B2(n730), .A(n726), .ZN(n562) );
  NAND2_X1 U144 ( .A1(\mem[4][3] ), .A2(n458), .ZN(n726) );
  OAI21_X1 U145 ( .B1(n481), .B2(n458), .A(n725), .ZN(n561) );
  NAND2_X1 U146 ( .A1(\mem[4][4] ), .A2(n458), .ZN(n725) );
  OAI21_X1 U147 ( .B1(n480), .B2(n730), .A(n724), .ZN(n560) );
  NAND2_X1 U148 ( .A1(\mem[4][5] ), .A2(n458), .ZN(n724) );
  OAI21_X1 U149 ( .B1(n479), .B2(n730), .A(n723), .ZN(n559) );
  NAND2_X1 U150 ( .A1(\mem[4][6] ), .A2(n458), .ZN(n723) );
  OAI21_X1 U151 ( .B1(n478), .B2(n730), .A(n722), .ZN(n558) );
  NAND2_X1 U152 ( .A1(\mem[4][7] ), .A2(n458), .ZN(n722) );
  OAI21_X1 U153 ( .B1(n477), .B2(n730), .A(n721), .ZN(n557) );
  NAND2_X1 U154 ( .A1(\mem[4][8] ), .A2(n458), .ZN(n721) );
  OAI21_X1 U155 ( .B1(n476), .B2(n730), .A(n720), .ZN(n556) );
  NAND2_X1 U156 ( .A1(\mem[4][9] ), .A2(n458), .ZN(n720) );
  OAI21_X1 U157 ( .B1(n475), .B2(n730), .A(n719), .ZN(n555) );
  NAND2_X1 U158 ( .A1(\mem[4][10] ), .A2(n458), .ZN(n719) );
  OAI21_X1 U159 ( .B1(n474), .B2(n730), .A(n718), .ZN(n554) );
  NAND2_X1 U160 ( .A1(\mem[4][11] ), .A2(n458), .ZN(n718) );
  OAI21_X1 U161 ( .B1(n473), .B2(n730), .A(n717), .ZN(n553) );
  NAND2_X1 U162 ( .A1(\mem[4][12] ), .A2(n730), .ZN(n717) );
  OAI21_X1 U163 ( .B1(n472), .B2(n458), .A(n716), .ZN(n552) );
  NAND2_X1 U164 ( .A1(\mem[4][13] ), .A2(n730), .ZN(n716) );
  OAI21_X1 U165 ( .B1(n471), .B2(n458), .A(n715), .ZN(n551) );
  NAND2_X1 U166 ( .A1(\mem[4][14] ), .A2(n730), .ZN(n715) );
  OAI21_X1 U167 ( .B1(n470), .B2(n730), .A(n714), .ZN(n550) );
  NAND2_X1 U168 ( .A1(\mem[4][15] ), .A2(n730), .ZN(n714) );
  OAI21_X1 U169 ( .B1(n469), .B2(n730), .A(n713), .ZN(n549) );
  NAND2_X1 U170 ( .A1(\mem[4][16] ), .A2(n730), .ZN(n713) );
  OAI21_X1 U171 ( .B1(n468), .B2(n730), .A(n712), .ZN(n548) );
  NAND2_X1 U172 ( .A1(\mem[4][17] ), .A2(n730), .ZN(n712) );
  OAI21_X1 U173 ( .B1(n467), .B2(n730), .A(n711), .ZN(n547) );
  NAND2_X1 U174 ( .A1(\mem[4][18] ), .A2(n730), .ZN(n711) );
  OAI21_X1 U175 ( .B1(n466), .B2(n730), .A(n710), .ZN(n546) );
  NAND2_X1 U176 ( .A1(\mem[4][19] ), .A2(n458), .ZN(n710) );
  OAI21_X1 U177 ( .B1(n485), .B2(n708), .A(n707), .ZN(n545) );
  NAND2_X1 U178 ( .A1(\mem[5][0] ), .A2(n457), .ZN(n707) );
  OAI21_X1 U179 ( .B1(n484), .B2(n708), .A(n706), .ZN(n544) );
  NAND2_X1 U180 ( .A1(\mem[5][1] ), .A2(n457), .ZN(n706) );
  OAI21_X1 U181 ( .B1(n483), .B2(n708), .A(n705), .ZN(n543) );
  NAND2_X1 U182 ( .A1(\mem[5][2] ), .A2(n457), .ZN(n705) );
  OAI21_X1 U183 ( .B1(n482), .B2(n708), .A(n704), .ZN(n542) );
  NAND2_X1 U184 ( .A1(\mem[5][3] ), .A2(n457), .ZN(n704) );
  OAI21_X1 U185 ( .B1(n481), .B2(n457), .A(n703), .ZN(n541) );
  NAND2_X1 U186 ( .A1(\mem[5][4] ), .A2(n457), .ZN(n703) );
  OAI21_X1 U187 ( .B1(n480), .B2(n708), .A(n702), .ZN(n540) );
  NAND2_X1 U188 ( .A1(\mem[5][5] ), .A2(n457), .ZN(n702) );
  OAI21_X1 U189 ( .B1(n479), .B2(n708), .A(n701), .ZN(n539) );
  NAND2_X1 U190 ( .A1(\mem[5][6] ), .A2(n457), .ZN(n701) );
  OAI21_X1 U191 ( .B1(n478), .B2(n708), .A(n700), .ZN(n538) );
  NAND2_X1 U192 ( .A1(\mem[5][7] ), .A2(n457), .ZN(n700) );
  OAI21_X1 U193 ( .B1(n477), .B2(n708), .A(n699), .ZN(n537) );
  NAND2_X1 U194 ( .A1(\mem[5][8] ), .A2(n457), .ZN(n699) );
  OAI21_X1 U195 ( .B1(n476), .B2(n708), .A(n698), .ZN(n536) );
  NAND2_X1 U196 ( .A1(\mem[5][9] ), .A2(n457), .ZN(n698) );
  OAI21_X1 U197 ( .B1(n475), .B2(n708), .A(n697), .ZN(n535) );
  NAND2_X1 U198 ( .A1(\mem[5][10] ), .A2(n457), .ZN(n697) );
  OAI21_X1 U199 ( .B1(n474), .B2(n708), .A(n696), .ZN(n534) );
  NAND2_X1 U200 ( .A1(\mem[5][11] ), .A2(n457), .ZN(n696) );
  OAI21_X1 U201 ( .B1(n473), .B2(n708), .A(n695), .ZN(n533) );
  NAND2_X1 U202 ( .A1(\mem[5][12] ), .A2(n708), .ZN(n695) );
  OAI21_X1 U203 ( .B1(n472), .B2(n457), .A(n694), .ZN(n532) );
  NAND2_X1 U204 ( .A1(\mem[5][13] ), .A2(n708), .ZN(n694) );
  OAI21_X1 U205 ( .B1(n471), .B2(n457), .A(n693), .ZN(n531) );
  NAND2_X1 U206 ( .A1(\mem[5][14] ), .A2(n708), .ZN(n693) );
  OAI21_X1 U207 ( .B1(n470), .B2(n708), .A(n692), .ZN(n530) );
  NAND2_X1 U208 ( .A1(\mem[5][15] ), .A2(n708), .ZN(n692) );
  OAI21_X1 U209 ( .B1(n469), .B2(n708), .A(n691), .ZN(n529) );
  NAND2_X1 U210 ( .A1(\mem[5][16] ), .A2(n708), .ZN(n691) );
  OAI21_X1 U211 ( .B1(n468), .B2(n708), .A(n690), .ZN(n528) );
  NAND2_X1 U212 ( .A1(\mem[5][17] ), .A2(n708), .ZN(n690) );
  OAI21_X1 U213 ( .B1(n467), .B2(n708), .A(n689), .ZN(n527) );
  NAND2_X1 U214 ( .A1(\mem[5][18] ), .A2(n708), .ZN(n689) );
  OAI21_X1 U215 ( .B1(n466), .B2(n708), .A(n688), .ZN(n526) );
  NAND2_X1 U216 ( .A1(\mem[5][19] ), .A2(n457), .ZN(n688) );
  OAI21_X1 U217 ( .B1(n485), .B2(n687), .A(n686), .ZN(n525) );
  NAND2_X1 U218 ( .A1(\mem[6][0] ), .A2(n456), .ZN(n686) );
  OAI21_X1 U219 ( .B1(n484), .B2(n687), .A(n685), .ZN(n524) );
  NAND2_X1 U220 ( .A1(\mem[6][1] ), .A2(n456), .ZN(n685) );
  OAI21_X1 U221 ( .B1(n483), .B2(n687), .A(n684), .ZN(n523) );
  NAND2_X1 U222 ( .A1(\mem[6][2] ), .A2(n456), .ZN(n684) );
  OAI21_X1 U223 ( .B1(n482), .B2(n687), .A(n683), .ZN(n522) );
  NAND2_X1 U224 ( .A1(\mem[6][3] ), .A2(n456), .ZN(n683) );
  OAI21_X1 U225 ( .B1(n481), .B2(n456), .A(n682), .ZN(n521) );
  NAND2_X1 U226 ( .A1(\mem[6][4] ), .A2(n456), .ZN(n682) );
  OAI21_X1 U227 ( .B1(n480), .B2(n687), .A(n681), .ZN(n520) );
  NAND2_X1 U228 ( .A1(\mem[6][5] ), .A2(n456), .ZN(n681) );
  OAI21_X1 U229 ( .B1(n479), .B2(n687), .A(n680), .ZN(n519) );
  NAND2_X1 U230 ( .A1(\mem[6][6] ), .A2(n456), .ZN(n680) );
  OAI21_X1 U231 ( .B1(n478), .B2(n687), .A(n679), .ZN(n518) );
  NAND2_X1 U232 ( .A1(\mem[6][7] ), .A2(n456), .ZN(n679) );
  OAI21_X1 U233 ( .B1(n477), .B2(n687), .A(n678), .ZN(n517) );
  NAND2_X1 U234 ( .A1(\mem[6][8] ), .A2(n456), .ZN(n678) );
  OAI21_X1 U235 ( .B1(n476), .B2(n687), .A(n677), .ZN(n516) );
  NAND2_X1 U236 ( .A1(\mem[6][9] ), .A2(n456), .ZN(n677) );
  OAI21_X1 U237 ( .B1(n475), .B2(n687), .A(n676), .ZN(n515) );
  NAND2_X1 U238 ( .A1(\mem[6][10] ), .A2(n456), .ZN(n676) );
  OAI21_X1 U239 ( .B1(n474), .B2(n687), .A(n675), .ZN(n514) );
  NAND2_X1 U240 ( .A1(\mem[6][11] ), .A2(n456), .ZN(n675) );
  OAI21_X1 U241 ( .B1(n473), .B2(n687), .A(n674), .ZN(n513) );
  NAND2_X1 U242 ( .A1(\mem[6][12] ), .A2(n687), .ZN(n674) );
  OAI21_X1 U243 ( .B1(n472), .B2(n456), .A(n673), .ZN(n512) );
  NAND2_X1 U244 ( .A1(\mem[6][13] ), .A2(n687), .ZN(n673) );
  OAI21_X1 U245 ( .B1(n471), .B2(n456), .A(n672), .ZN(n511) );
  NAND2_X1 U246 ( .A1(\mem[6][14] ), .A2(n687), .ZN(n672) );
  OAI21_X1 U247 ( .B1(n470), .B2(n687), .A(n671), .ZN(n510) );
  NAND2_X1 U248 ( .A1(\mem[6][15] ), .A2(n687), .ZN(n671) );
  OAI21_X1 U249 ( .B1(n469), .B2(n687), .A(n670), .ZN(n509) );
  NAND2_X1 U250 ( .A1(\mem[6][16] ), .A2(n687), .ZN(n670) );
  OAI21_X1 U251 ( .B1(n468), .B2(n687), .A(n669), .ZN(n508) );
  NAND2_X1 U252 ( .A1(\mem[6][17] ), .A2(n687), .ZN(n669) );
  OAI21_X1 U253 ( .B1(n467), .B2(n687), .A(n668), .ZN(n507) );
  NAND2_X1 U254 ( .A1(\mem[6][18] ), .A2(n687), .ZN(n668) );
  OAI21_X1 U255 ( .B1(n466), .B2(n687), .A(n667), .ZN(n506) );
  NAND2_X1 U256 ( .A1(\mem[6][19] ), .A2(n456), .ZN(n667) );
  OAI21_X1 U257 ( .B1(n485), .B2(n666), .A(n665), .ZN(n505) );
  NAND2_X1 U258 ( .A1(\mem[7][0] ), .A2(n666), .ZN(n665) );
  OAI21_X1 U259 ( .B1(n484), .B2(n455), .A(n664), .ZN(n504) );
  NAND2_X1 U260 ( .A1(\mem[7][1] ), .A2(n666), .ZN(n664) );
  OAI21_X1 U261 ( .B1(n483), .B2(n455), .A(n663), .ZN(n503) );
  NAND2_X1 U262 ( .A1(\mem[7][2] ), .A2(n666), .ZN(n663) );
  OAI21_X1 U263 ( .B1(n482), .B2(n455), .A(n662), .ZN(n502) );
  NAND2_X1 U264 ( .A1(\mem[7][3] ), .A2(n666), .ZN(n662) );
  OAI21_X1 U265 ( .B1(n481), .B2(n455), .A(n661), .ZN(n501) );
  NAND2_X1 U266 ( .A1(\mem[7][4] ), .A2(n666), .ZN(n661) );
  OAI21_X1 U267 ( .B1(n480), .B2(n455), .A(n660), .ZN(n500) );
  NAND2_X1 U268 ( .A1(\mem[7][5] ), .A2(n666), .ZN(n660) );
  OAI21_X1 U269 ( .B1(n479), .B2(n455), .A(n659), .ZN(n499) );
  NAND2_X1 U270 ( .A1(\mem[7][6] ), .A2(n666), .ZN(n659) );
  OAI21_X1 U271 ( .B1(n478), .B2(n455), .A(n658), .ZN(n498) );
  NAND2_X1 U272 ( .A1(\mem[7][7] ), .A2(n666), .ZN(n658) );
  OAI21_X1 U273 ( .B1(n477), .B2(n455), .A(n657), .ZN(n497) );
  NAND2_X1 U274 ( .A1(\mem[7][8] ), .A2(n666), .ZN(n657) );
  OAI21_X1 U275 ( .B1(n476), .B2(n666), .A(n656), .ZN(n496) );
  NAND2_X1 U276 ( .A1(\mem[7][9] ), .A2(n666), .ZN(n656) );
  OAI21_X1 U277 ( .B1(n475), .B2(n455), .A(n655), .ZN(n495) );
  NAND2_X1 U278 ( .A1(\mem[7][10] ), .A2(n666), .ZN(n655) );
  OAI21_X1 U279 ( .B1(n474), .B2(n455), .A(n654), .ZN(n494) );
  NAND2_X1 U280 ( .A1(\mem[7][11] ), .A2(n666), .ZN(n654) );
  OAI21_X1 U281 ( .B1(n473), .B2(n666), .A(n653), .ZN(n493) );
  NAND2_X1 U282 ( .A1(\mem[7][12] ), .A2(n666), .ZN(n653) );
  OAI21_X1 U283 ( .B1(n472), .B2(n455), .A(n652), .ZN(n492) );
  NAND2_X1 U284 ( .A1(\mem[7][13] ), .A2(n666), .ZN(n652) );
  OAI21_X1 U285 ( .B1(n471), .B2(n666), .A(n651), .ZN(n491) );
  NAND2_X1 U286 ( .A1(\mem[7][14] ), .A2(n666), .ZN(n651) );
  OAI21_X1 U287 ( .B1(n470), .B2(n455), .A(n650), .ZN(n490) );
  NAND2_X1 U288 ( .A1(\mem[7][15] ), .A2(n666), .ZN(n650) );
  OAI21_X1 U289 ( .B1(n469), .B2(n455), .A(n649), .ZN(n489) );
  NAND2_X1 U290 ( .A1(\mem[7][16] ), .A2(n666), .ZN(n649) );
  OAI21_X1 U291 ( .B1(n468), .B2(n455), .A(n648), .ZN(n488) );
  NAND2_X1 U292 ( .A1(\mem[7][17] ), .A2(n666), .ZN(n648) );
  OAI21_X1 U293 ( .B1(n467), .B2(n455), .A(n647), .ZN(n487) );
  NAND2_X1 U294 ( .A1(\mem[7][18] ), .A2(n666), .ZN(n647) );
  OAI21_X1 U295 ( .B1(n466), .B2(n455), .A(n646), .ZN(n486) );
  NAND2_X1 U296 ( .A1(\mem[7][19] ), .A2(n666), .ZN(n646) );
  OAI21_X1 U297 ( .B1(n462), .B2(n483), .A(n812), .ZN(n643) );
  NAND2_X1 U298 ( .A1(\mem[0][2] ), .A2(n462), .ZN(n812) );
  OAI21_X1 U299 ( .B1(n815), .B2(n482), .A(n811), .ZN(n642) );
  NAND2_X1 U300 ( .A1(\mem[0][3] ), .A2(n462), .ZN(n811) );
  OAI21_X1 U301 ( .B1(n815), .B2(n481), .A(n810), .ZN(n641) );
  NAND2_X1 U302 ( .A1(\mem[0][4] ), .A2(n462), .ZN(n810) );
  OAI21_X1 U303 ( .B1(n815), .B2(n480), .A(n809), .ZN(n640) );
  NAND2_X1 U304 ( .A1(\mem[0][5] ), .A2(n462), .ZN(n809) );
  OAI21_X1 U305 ( .B1(n815), .B2(n479), .A(n808), .ZN(n639) );
  NAND2_X1 U306 ( .A1(\mem[0][6] ), .A2(n462), .ZN(n808) );
  OAI21_X1 U307 ( .B1(n815), .B2(n478), .A(n807), .ZN(n638) );
  NAND2_X1 U308 ( .A1(\mem[0][7] ), .A2(n462), .ZN(n807) );
  OAI21_X1 U309 ( .B1(n815), .B2(n477), .A(n806), .ZN(n637) );
  NAND2_X1 U310 ( .A1(\mem[0][8] ), .A2(n462), .ZN(n806) );
  OAI21_X1 U311 ( .B1(n815), .B2(n476), .A(n805), .ZN(n636) );
  NAND2_X1 U312 ( .A1(\mem[0][9] ), .A2(n462), .ZN(n805) );
  OAI21_X1 U313 ( .B1(n815), .B2(n475), .A(n804), .ZN(n635) );
  NAND2_X1 U314 ( .A1(\mem[0][10] ), .A2(n462), .ZN(n804) );
  OAI21_X1 U315 ( .B1(n815), .B2(n474), .A(n803), .ZN(n634) );
  NAND2_X1 U316 ( .A1(\mem[0][11] ), .A2(n462), .ZN(n803) );
  OAI21_X1 U317 ( .B1(n815), .B2(n473), .A(n802), .ZN(n633) );
  NAND2_X1 U318 ( .A1(\mem[0][12] ), .A2(n815), .ZN(n802) );
  OAI21_X1 U319 ( .B1(n815), .B2(n472), .A(n801), .ZN(n632) );
  NAND2_X1 U320 ( .A1(\mem[0][13] ), .A2(n815), .ZN(n801) );
  OAI21_X1 U321 ( .B1(n462), .B2(n471), .A(n800), .ZN(n631) );
  NAND2_X1 U322 ( .A1(\mem[0][14] ), .A2(n815), .ZN(n800) );
  OAI21_X1 U323 ( .B1(n815), .B2(n470), .A(n799), .ZN(n630) );
  NAND2_X1 U324 ( .A1(\mem[0][15] ), .A2(n815), .ZN(n799) );
  OAI21_X1 U325 ( .B1(n815), .B2(n469), .A(n798), .ZN(n629) );
  NAND2_X1 U326 ( .A1(\mem[0][16] ), .A2(n815), .ZN(n798) );
  OAI21_X1 U327 ( .B1(n815), .B2(n468), .A(n797), .ZN(n628) );
  NAND2_X1 U328 ( .A1(\mem[0][17] ), .A2(n815), .ZN(n797) );
  OAI21_X1 U329 ( .B1(n815), .B2(n467), .A(n796), .ZN(n627) );
  NAND2_X1 U330 ( .A1(\mem[0][18] ), .A2(n815), .ZN(n796) );
  OAI21_X1 U331 ( .B1(n815), .B2(n485), .A(n814), .ZN(n645) );
  NAND2_X1 U332 ( .A1(\mem[0][0] ), .A2(n462), .ZN(n814) );
  OAI21_X1 U333 ( .B1(n462), .B2(n484), .A(n813), .ZN(n644) );
  NAND2_X1 U334 ( .A1(\mem[0][1] ), .A2(n462), .ZN(n813) );
  OAI21_X1 U335 ( .B1(n815), .B2(n466), .A(n795), .ZN(n626) );
  NAND2_X1 U336 ( .A1(\mem[0][19] ), .A2(n462), .ZN(n795) );
  INV_X1 U337 ( .A(N10), .ZN(n463) );
  INV_X1 U338 ( .A(N11), .ZN(n464) );
  INV_X1 U339 ( .A(data_in[0]), .ZN(n485) );
  INV_X1 U340 ( .A(data_in[1]), .ZN(n484) );
  INV_X1 U341 ( .A(data_in[2]), .ZN(n483) );
  INV_X1 U342 ( .A(data_in[3]), .ZN(n482) );
  INV_X1 U343 ( .A(data_in[4]), .ZN(n481) );
  INV_X1 U344 ( .A(data_in[5]), .ZN(n480) );
  INV_X1 U345 ( .A(data_in[6]), .ZN(n479) );
  INV_X1 U346 ( .A(data_in[7]), .ZN(n478) );
  INV_X1 U347 ( .A(data_in[8]), .ZN(n477) );
  INV_X1 U356 ( .A(data_in[9]), .ZN(n476) );
  INV_X1 U357 ( .A(data_in[10]), .ZN(n475) );
  INV_X1 U358 ( .A(data_in[11]), .ZN(n474) );
  INV_X1 U359 ( .A(data_in[12]), .ZN(n473) );
  INV_X1 U360 ( .A(data_in[13]), .ZN(n472) );
  INV_X1 U361 ( .A(data_in[14]), .ZN(n471) );
  INV_X1 U362 ( .A(data_in[15]), .ZN(n470) );
  INV_X1 U363 ( .A(data_in[16]), .ZN(n469) );
  INV_X1 U364 ( .A(data_in[17]), .ZN(n468) );
  INV_X1 U365 ( .A(data_in[18]), .ZN(n467) );
  INV_X1 U366 ( .A(data_in[19]), .ZN(n466) );
  MUX2_X1 U367 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n452), .Z(n1) );
  MUX2_X1 U368 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n452), .Z(n2) );
  MUX2_X1 U369 ( .A(n2), .B(n1), .S(n451), .Z(n3) );
  MUX2_X1 U370 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n452), .Z(n4) );
  MUX2_X1 U371 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n452), .Z(n5) );
  MUX2_X1 U372 ( .A(n5), .B(n4), .S(n451), .Z(n6) );
  MUX2_X1 U373 ( .A(n6), .B(n3), .S(N12), .Z(N32) );
  MUX2_X1 U374 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n452), .Z(n7) );
  MUX2_X1 U375 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n452), .Z(n8) );
  MUX2_X1 U376 ( .A(n8), .B(n7), .S(N11), .Z(n9) );
  MUX2_X1 U377 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n452), .Z(n10) );
  MUX2_X1 U378 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n452), .Z(n11) );
  MUX2_X1 U379 ( .A(n11), .B(n10), .S(n451), .Z(n12) );
  MUX2_X1 U380 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n452), .Z(n13) );
  MUX2_X1 U381 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n452), .Z(n14) );
  MUX2_X1 U382 ( .A(n14), .B(n13), .S(n451), .Z(n15) );
  MUX2_X1 U383 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n452), .Z(n16) );
  MUX2_X1 U384 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n453), .Z(n17) );
  MUX2_X1 U385 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U386 ( .A(n18), .B(n15), .S(N12), .Z(N30) );
  MUX2_X1 U387 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n454), .Z(n19) );
  MUX2_X1 U388 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n454), .Z(n20) );
  MUX2_X1 U389 ( .A(n20), .B(n19), .S(N11), .Z(n21) );
  MUX2_X1 U390 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n452), .Z(n22) );
  MUX2_X1 U391 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n454), .Z(n23) );
  MUX2_X1 U392 ( .A(n23), .B(n22), .S(N11), .Z(n354) );
  MUX2_X1 U393 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(N10), .Z(n355) );
  MUX2_X1 U394 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n453), .Z(n356) );
  MUX2_X1 U395 ( .A(n356), .B(n355), .S(N11), .Z(n357) );
  MUX2_X1 U396 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n453), .Z(n358) );
  MUX2_X1 U397 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n359) );
  MUX2_X1 U398 ( .A(n359), .B(n358), .S(N11), .Z(n360) );
  MUX2_X1 U399 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n453), .Z(n361) );
  MUX2_X1 U400 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n453), .Z(n362) );
  MUX2_X1 U401 ( .A(n362), .B(n361), .S(N11), .Z(n363) );
  MUX2_X1 U402 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n453), .Z(n364) );
  MUX2_X1 U403 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n453), .Z(n365) );
  MUX2_X1 U404 ( .A(n365), .B(n364), .S(N11), .Z(n366) );
  MUX2_X1 U405 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n453), .Z(n367) );
  MUX2_X1 U406 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n453), .Z(n368) );
  MUX2_X1 U407 ( .A(n368), .B(n367), .S(n451), .Z(n369) );
  MUX2_X1 U408 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n453), .Z(n370) );
  MUX2_X1 U409 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n453), .Z(n371) );
  MUX2_X1 U410 ( .A(n371), .B(n370), .S(N11), .Z(n372) );
  MUX2_X1 U411 ( .A(n372), .B(n369), .S(N12), .Z(N26) );
  MUX2_X1 U412 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n453), .Z(n373) );
  MUX2_X1 U413 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n453), .Z(n374) );
  MUX2_X1 U414 ( .A(n374), .B(n373), .S(N11), .Z(n375) );
  MUX2_X1 U415 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n453), .Z(n376) );
  MUX2_X1 U416 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n453), .Z(n377) );
  MUX2_X1 U417 ( .A(n377), .B(n376), .S(N11), .Z(n378) );
  MUX2_X1 U418 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n454), .Z(n379) );
  MUX2_X1 U419 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n454), .Z(n380) );
  MUX2_X1 U420 ( .A(n380), .B(n379), .S(n451), .Z(n381) );
  MUX2_X1 U421 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n454), .Z(n382) );
  MUX2_X1 U422 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n454), .Z(n383) );
  MUX2_X1 U423 ( .A(n383), .B(n382), .S(n451), .Z(n384) );
  MUX2_X1 U424 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n454), .Z(n385) );
  MUX2_X1 U425 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n454), .Z(n386) );
  MUX2_X1 U426 ( .A(n386), .B(n385), .S(n451), .Z(n387) );
  MUX2_X1 U427 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n454), .Z(n388) );
  MUX2_X1 U428 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n454), .Z(n389) );
  MUX2_X1 U429 ( .A(n389), .B(n388), .S(n451), .Z(n390) );
  MUX2_X1 U430 ( .A(n390), .B(n387), .S(N12), .Z(N23) );
  MUX2_X1 U431 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n454), .Z(n391) );
  MUX2_X1 U432 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n454), .Z(n392) );
  MUX2_X1 U433 ( .A(n392), .B(n391), .S(n451), .Z(n393) );
  MUX2_X1 U434 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n454), .Z(n394) );
  MUX2_X1 U435 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n454), .Z(n395) );
  MUX2_X1 U436 ( .A(n395), .B(n394), .S(n451), .Z(n396) );
  MUX2_X1 U437 ( .A(n396), .B(n393), .S(N12), .Z(N22) );
  MUX2_X1 U438 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n452), .Z(n397) );
  MUX2_X1 U439 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(N10), .Z(n398) );
  MUX2_X1 U440 ( .A(n398), .B(n397), .S(n451), .Z(n399) );
  MUX2_X1 U441 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(N10), .Z(n400) );
  MUX2_X1 U442 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(N10), .Z(n401) );
  MUX2_X1 U443 ( .A(n401), .B(n400), .S(n451), .Z(n402) );
  MUX2_X1 U444 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n454), .Z(n403) );
  MUX2_X1 U445 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n452), .Z(n404) );
  MUX2_X1 U446 ( .A(n404), .B(n403), .S(n451), .Z(n405) );
  MUX2_X1 U447 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n453), .Z(n406) );
  MUX2_X1 U448 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n453), .Z(n407) );
  MUX2_X1 U449 ( .A(n407), .B(n406), .S(n451), .Z(n408) );
  MUX2_X1 U450 ( .A(n408), .B(n405), .S(N12), .Z(N20) );
  MUX2_X1 U451 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n452), .Z(n409) );
  MUX2_X1 U452 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(N10), .Z(n410) );
  MUX2_X1 U453 ( .A(n410), .B(n409), .S(n451), .Z(n411) );
  MUX2_X1 U454 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(N10), .Z(n412) );
  MUX2_X1 U455 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(N10), .Z(n413) );
  MUX2_X1 U456 ( .A(n413), .B(n412), .S(n451), .Z(n414) );
  MUX2_X1 U457 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n453), .Z(n415) );
  MUX2_X1 U458 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n454), .Z(n416) );
  MUX2_X1 U459 ( .A(n416), .B(n415), .S(n451), .Z(n417) );
  MUX2_X1 U460 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n453), .Z(n418) );
  MUX2_X1 U461 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n454), .Z(n419) );
  MUX2_X1 U462 ( .A(n419), .B(n418), .S(n451), .Z(n420) );
  MUX2_X1 U463 ( .A(n420), .B(n417), .S(N12), .Z(N18) );
  MUX2_X1 U464 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n452), .Z(n421) );
  MUX2_X1 U465 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n452), .Z(n422) );
  MUX2_X1 U466 ( .A(n422), .B(n421), .S(N11), .Z(n423) );
  MUX2_X1 U467 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(N10), .Z(n424) );
  MUX2_X1 U468 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n452), .Z(n425) );
  MUX2_X1 U469 ( .A(n425), .B(n424), .S(N11), .Z(n426) );
  MUX2_X1 U470 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n454), .Z(n427) );
  MUX2_X1 U471 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n454), .Z(n428) );
  MUX2_X1 U472 ( .A(n428), .B(n427), .S(n451), .Z(n429) );
  MUX2_X1 U473 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n452), .Z(n430) );
  MUX2_X1 U474 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n453), .Z(n431) );
  MUX2_X1 U475 ( .A(n431), .B(n430), .S(N11), .Z(n432) );
  MUX2_X1 U476 ( .A(n432), .B(n429), .S(N12), .Z(N16) );
  MUX2_X1 U477 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n454), .Z(n433) );
  MUX2_X1 U478 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n452), .Z(n434) );
  MUX2_X1 U479 ( .A(n434), .B(n433), .S(n451), .Z(n435) );
  MUX2_X1 U480 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n452), .Z(n436) );
  MUX2_X1 U481 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n453), .Z(n437) );
  MUX2_X1 U482 ( .A(n437), .B(n436), .S(N11), .Z(n438) );
  MUX2_X1 U483 ( .A(n438), .B(n435), .S(N12), .Z(N15) );
  MUX2_X1 U484 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n454), .Z(n439) );
  MUX2_X1 U485 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n452), .Z(n440) );
  MUX2_X1 U486 ( .A(n440), .B(n439), .S(N11), .Z(n441) );
  MUX2_X1 U487 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n454), .Z(n442) );
  MUX2_X1 U488 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n452), .Z(n443) );
  MUX2_X1 U489 ( .A(n443), .B(n442), .S(n451), .Z(n444) );
  MUX2_X1 U490 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(N10), .Z(n445) );
  MUX2_X1 U491 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n453), .Z(n446) );
  MUX2_X1 U492 ( .A(n446), .B(n445), .S(N11), .Z(n447) );
  MUX2_X1 U493 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(N10), .Z(n448) );
  MUX2_X1 U494 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n453), .Z(n449) );
  MUX2_X1 U495 ( .A(n449), .B(n448), .S(n451), .Z(n450) );
  CLKBUF_X1 U496 ( .A(N10), .Z(n452) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE3_7 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N14, N16, N18, N20, N22, N24, N26, N28, N32, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[18]  ( .D(N14), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[16]  ( .D(N16), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N20), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N22), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[8]  ( .D(N24), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N26), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N28), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[0]  ( .D(N32), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n486), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n487), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n488), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n489), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n490), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n491), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n492), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n493), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n494), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n495), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n496), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n497), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n498), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n499), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n500), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n501), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n502), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n503), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n504), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n505), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n506), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n507), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n508), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n509), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n510), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n511), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n512), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n513), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n514), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n515), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n516), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n517), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n518), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n519), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n520), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n521), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n522), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n523), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n524), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n525), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n526), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n527), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n528), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n529), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n530), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n531), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n532), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n533), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n534), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n535), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n536), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n537), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n538), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n539), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n540), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n541), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n542), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n543), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n544), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n545), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n546), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n547), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n548), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n549), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n550), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n551), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n552), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n553), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n554), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n555), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n556), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n557), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n558), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n559), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n560), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n561), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n562), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n563), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n564), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n565), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n566), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n567), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n568), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n569), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n570), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n571), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n572), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n573), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n574), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n575), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n576), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n577), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n578), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n579), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n580), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n581), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n582), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n583), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n584), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n585), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n586), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n587), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n588), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n589), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n590), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n591), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n592), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n593), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n594), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n595), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n596), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n597), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n598), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n599), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n600), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n601), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n602), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n603), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n604), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n605), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n606), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n607), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n608), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n609), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n610), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n611), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n612), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n613), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n614), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n615), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n616), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n617), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n618), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n619), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n620), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n621), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n622), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n623), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n624), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n625), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n626), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n627), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n628), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n629), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n630), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n631), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n632), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n633), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n634), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n635), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n636), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n637), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n638), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n639), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n640), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n641), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n642), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n643), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n644), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n645), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U348 ( .A1(n463), .A2(n464), .A3(n794), .ZN(n815) );
  NAND3_X1 U349 ( .A1(n794), .A2(n464), .A3(N10), .ZN(n793) );
  NAND3_X1 U350 ( .A1(n794), .A2(n463), .A3(N11), .ZN(n772) );
  NAND3_X1 U351 ( .A1(N10), .A2(n794), .A3(N11), .ZN(n751) );
  NAND3_X1 U352 ( .A1(n463), .A2(n464), .A3(n709), .ZN(n730) );
  NAND3_X1 U353 ( .A1(N10), .A2(n464), .A3(n709), .ZN(n708) );
  NAND3_X1 U354 ( .A1(N11), .A2(n463), .A3(n709), .ZN(n687) );
  NAND3_X1 U355 ( .A1(N11), .A2(N10), .A3(n709), .ZN(n666) );
  SDFF_X1 \data_out_reg[11]  ( .D(n402), .SI(n399), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n414), .SI(n411), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n426), .SI(n423), .SE(N12), .CK(clk), .Q(
        data_out[15]) );
  SDFF_X1 \data_out_reg[19]  ( .D(n450), .SI(n447), .SE(N12), .CK(clk), .Q(
        data_out[19]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n354), .SI(n21), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n12), .SI(n9), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[17]  ( .D(n438), .SI(n435), .SE(N12), .CK(clk), .Q(
        data_out[17]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n366), .SI(n363), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n378), .SI(n375), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n390), .SI(n387), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[2]  ( .D(n18), .SI(n15), .SE(N12), .CK(clk), .Q(
        data_out[2]) );
  BUF_X1 U3 ( .A(n666), .Z(n455) );
  BUF_X1 U4 ( .A(n772), .Z(n460) );
  BUF_X1 U5 ( .A(n730), .Z(n458) );
  BUF_X1 U6 ( .A(n815), .Z(n462) );
  BUF_X1 U7 ( .A(n751), .Z(n459) );
  BUF_X1 U8 ( .A(n793), .Z(n461) );
  BUF_X1 U9 ( .A(n687), .Z(n456) );
  BUF_X1 U10 ( .A(n708), .Z(n457) );
  BUF_X1 U11 ( .A(N10), .Z(n454) );
  BUF_X1 U12 ( .A(N10), .Z(n453) );
  BUF_X1 U13 ( .A(N11), .Z(n451) );
  AND2_X1 U14 ( .A1(N12), .A2(wr_en), .ZN(n709) );
  OAI21_X1 U15 ( .B1(n485), .B2(n793), .A(n792), .ZN(n625) );
  NAND2_X1 U16 ( .A1(\mem[1][0] ), .A2(n461), .ZN(n792) );
  OAI21_X1 U17 ( .B1(n484), .B2(n793), .A(n791), .ZN(n624) );
  NAND2_X1 U18 ( .A1(\mem[1][1] ), .A2(n461), .ZN(n791) );
  OAI21_X1 U19 ( .B1(n483), .B2(n793), .A(n790), .ZN(n623) );
  NAND2_X1 U20 ( .A1(\mem[1][2] ), .A2(n461), .ZN(n790) );
  OAI21_X1 U21 ( .B1(n482), .B2(n793), .A(n789), .ZN(n622) );
  NAND2_X1 U22 ( .A1(\mem[1][3] ), .A2(n461), .ZN(n789) );
  OAI21_X1 U23 ( .B1(n481), .B2(n461), .A(n788), .ZN(n621) );
  NAND2_X1 U24 ( .A1(\mem[1][4] ), .A2(n461), .ZN(n788) );
  OAI21_X1 U25 ( .B1(n480), .B2(n461), .A(n787), .ZN(n620) );
  NAND2_X1 U26 ( .A1(\mem[1][5] ), .A2(n461), .ZN(n787) );
  OAI21_X1 U27 ( .B1(n479), .B2(n793), .A(n786), .ZN(n619) );
  NAND2_X1 U28 ( .A1(\mem[1][6] ), .A2(n461), .ZN(n786) );
  OAI21_X1 U29 ( .B1(n478), .B2(n793), .A(n785), .ZN(n618) );
  NAND2_X1 U30 ( .A1(\mem[1][7] ), .A2(n461), .ZN(n785) );
  OAI21_X1 U31 ( .B1(n477), .B2(n793), .A(n784), .ZN(n617) );
  NAND2_X1 U32 ( .A1(\mem[1][8] ), .A2(n461), .ZN(n784) );
  OAI21_X1 U33 ( .B1(n476), .B2(n793), .A(n783), .ZN(n616) );
  NAND2_X1 U34 ( .A1(\mem[1][9] ), .A2(n461), .ZN(n783) );
  OAI21_X1 U35 ( .B1(n475), .B2(n793), .A(n782), .ZN(n615) );
  NAND2_X1 U36 ( .A1(\mem[1][10] ), .A2(n461), .ZN(n782) );
  OAI21_X1 U37 ( .B1(n474), .B2(n793), .A(n781), .ZN(n614) );
  NAND2_X1 U38 ( .A1(\mem[1][11] ), .A2(n461), .ZN(n781) );
  OAI21_X1 U39 ( .B1(n473), .B2(n793), .A(n780), .ZN(n613) );
  NAND2_X1 U40 ( .A1(\mem[1][12] ), .A2(n793), .ZN(n780) );
  OAI21_X1 U41 ( .B1(n472), .B2(n793), .A(n779), .ZN(n612) );
  NAND2_X1 U42 ( .A1(\mem[1][13] ), .A2(n793), .ZN(n779) );
  OAI21_X1 U43 ( .B1(n471), .B2(n793), .A(n778), .ZN(n611) );
  NAND2_X1 U44 ( .A1(\mem[1][14] ), .A2(n793), .ZN(n778) );
  OAI21_X1 U45 ( .B1(n470), .B2(n793), .A(n777), .ZN(n610) );
  NAND2_X1 U46 ( .A1(\mem[1][15] ), .A2(n461), .ZN(n777) );
  OAI21_X1 U47 ( .B1(n469), .B2(n793), .A(n776), .ZN(n609) );
  NAND2_X1 U48 ( .A1(\mem[1][16] ), .A2(n793), .ZN(n776) );
  OAI21_X1 U49 ( .B1(n468), .B2(n793), .A(n775), .ZN(n608) );
  NAND2_X1 U50 ( .A1(\mem[1][17] ), .A2(n793), .ZN(n775) );
  OAI21_X1 U51 ( .B1(n467), .B2(n793), .A(n774), .ZN(n607) );
  NAND2_X1 U52 ( .A1(\mem[1][18] ), .A2(n793), .ZN(n774) );
  OAI21_X1 U53 ( .B1(n466), .B2(n793), .A(n773), .ZN(n606) );
  NAND2_X1 U54 ( .A1(\mem[1][19] ), .A2(n461), .ZN(n773) );
  OAI21_X1 U55 ( .B1(n485), .B2(n772), .A(n771), .ZN(n605) );
  NAND2_X1 U56 ( .A1(\mem[2][0] ), .A2(n772), .ZN(n771) );
  OAI21_X1 U57 ( .B1(n484), .B2(n772), .A(n770), .ZN(n604) );
  NAND2_X1 U58 ( .A1(\mem[2][1] ), .A2(n772), .ZN(n770) );
  OAI21_X1 U59 ( .B1(n483), .B2(n772), .A(n769), .ZN(n603) );
  NAND2_X1 U60 ( .A1(\mem[2][2] ), .A2(n772), .ZN(n769) );
  OAI21_X1 U61 ( .B1(n482), .B2(n460), .A(n768), .ZN(n602) );
  NAND2_X1 U62 ( .A1(\mem[2][3] ), .A2(n772), .ZN(n768) );
  OAI21_X1 U63 ( .B1(n481), .B2(n460), .A(n767), .ZN(n601) );
  NAND2_X1 U64 ( .A1(\mem[2][4] ), .A2(n772), .ZN(n767) );
  OAI21_X1 U65 ( .B1(n480), .B2(n460), .A(n766), .ZN(n600) );
  NAND2_X1 U66 ( .A1(\mem[2][5] ), .A2(n772), .ZN(n766) );
  OAI21_X1 U67 ( .B1(n479), .B2(n460), .A(n765), .ZN(n599) );
  NAND2_X1 U68 ( .A1(\mem[2][6] ), .A2(n772), .ZN(n765) );
  OAI21_X1 U69 ( .B1(n478), .B2(n460), .A(n764), .ZN(n598) );
  NAND2_X1 U70 ( .A1(\mem[2][7] ), .A2(n772), .ZN(n764) );
  OAI21_X1 U71 ( .B1(n477), .B2(n460), .A(n763), .ZN(n597) );
  NAND2_X1 U72 ( .A1(\mem[2][8] ), .A2(n772), .ZN(n763) );
  OAI21_X1 U73 ( .B1(n476), .B2(n460), .A(n762), .ZN(n596) );
  NAND2_X1 U74 ( .A1(\mem[2][9] ), .A2(n772), .ZN(n762) );
  OAI21_X1 U75 ( .B1(n475), .B2(n460), .A(n761), .ZN(n595) );
  NAND2_X1 U76 ( .A1(\mem[2][10] ), .A2(n772), .ZN(n761) );
  OAI21_X1 U77 ( .B1(n474), .B2(n460), .A(n760), .ZN(n594) );
  NAND2_X1 U78 ( .A1(\mem[2][11] ), .A2(n772), .ZN(n760) );
  OAI21_X1 U79 ( .B1(n473), .B2(n460), .A(n759), .ZN(n593) );
  NAND2_X1 U80 ( .A1(\mem[2][12] ), .A2(n772), .ZN(n759) );
  OAI21_X1 U81 ( .B1(n472), .B2(n460), .A(n758), .ZN(n592) );
  NAND2_X1 U82 ( .A1(\mem[2][13] ), .A2(n772), .ZN(n758) );
  OAI21_X1 U83 ( .B1(n471), .B2(n460), .A(n757), .ZN(n591) );
  NAND2_X1 U84 ( .A1(\mem[2][14] ), .A2(n772), .ZN(n757) );
  OAI21_X1 U85 ( .B1(n470), .B2(n460), .A(n756), .ZN(n590) );
  NAND2_X1 U86 ( .A1(\mem[2][15] ), .A2(n772), .ZN(n756) );
  OAI21_X1 U87 ( .B1(n469), .B2(n460), .A(n755), .ZN(n589) );
  NAND2_X1 U88 ( .A1(\mem[2][16] ), .A2(n772), .ZN(n755) );
  OAI21_X1 U89 ( .B1(n468), .B2(n460), .A(n754), .ZN(n588) );
  NAND2_X1 U90 ( .A1(\mem[2][17] ), .A2(n772), .ZN(n754) );
  OAI21_X1 U91 ( .B1(n467), .B2(n460), .A(n753), .ZN(n587) );
  NAND2_X1 U92 ( .A1(\mem[2][18] ), .A2(n772), .ZN(n753) );
  OAI21_X1 U93 ( .B1(n466), .B2(n772), .A(n752), .ZN(n586) );
  NAND2_X1 U94 ( .A1(\mem[2][19] ), .A2(n772), .ZN(n752) );
  OAI21_X1 U95 ( .B1(n485), .B2(n751), .A(n750), .ZN(n585) );
  NAND2_X1 U96 ( .A1(\mem[3][0] ), .A2(n459), .ZN(n750) );
  OAI21_X1 U97 ( .B1(n484), .B2(n751), .A(n749), .ZN(n584) );
  NAND2_X1 U98 ( .A1(\mem[3][1] ), .A2(n459), .ZN(n749) );
  OAI21_X1 U99 ( .B1(n483), .B2(n751), .A(n748), .ZN(n583) );
  NAND2_X1 U100 ( .A1(\mem[3][2] ), .A2(n459), .ZN(n748) );
  OAI21_X1 U101 ( .B1(n482), .B2(n751), .A(n747), .ZN(n582) );
  NAND2_X1 U102 ( .A1(\mem[3][3] ), .A2(n459), .ZN(n747) );
  OAI21_X1 U103 ( .B1(n481), .B2(n459), .A(n746), .ZN(n581) );
  NAND2_X1 U104 ( .A1(\mem[3][4] ), .A2(n459), .ZN(n746) );
  OAI21_X1 U105 ( .B1(n480), .B2(n459), .A(n745), .ZN(n580) );
  NAND2_X1 U106 ( .A1(\mem[3][5] ), .A2(n459), .ZN(n745) );
  OAI21_X1 U107 ( .B1(n479), .B2(n751), .A(n744), .ZN(n579) );
  NAND2_X1 U108 ( .A1(\mem[3][6] ), .A2(n459), .ZN(n744) );
  OAI21_X1 U109 ( .B1(n478), .B2(n751), .A(n743), .ZN(n578) );
  NAND2_X1 U110 ( .A1(\mem[3][7] ), .A2(n459), .ZN(n743) );
  OAI21_X1 U111 ( .B1(n477), .B2(n751), .A(n742), .ZN(n577) );
  NAND2_X1 U112 ( .A1(\mem[3][8] ), .A2(n459), .ZN(n742) );
  OAI21_X1 U113 ( .B1(n476), .B2(n751), .A(n741), .ZN(n576) );
  NAND2_X1 U114 ( .A1(\mem[3][9] ), .A2(n459), .ZN(n741) );
  OAI21_X1 U115 ( .B1(n475), .B2(n751), .A(n740), .ZN(n575) );
  NAND2_X1 U116 ( .A1(\mem[3][10] ), .A2(n459), .ZN(n740) );
  OAI21_X1 U117 ( .B1(n474), .B2(n751), .A(n739), .ZN(n574) );
  NAND2_X1 U118 ( .A1(\mem[3][11] ), .A2(n459), .ZN(n739) );
  OAI21_X1 U119 ( .B1(n473), .B2(n751), .A(n738), .ZN(n573) );
  NAND2_X1 U120 ( .A1(\mem[3][12] ), .A2(n751), .ZN(n738) );
  OAI21_X1 U121 ( .B1(n472), .B2(n751), .A(n737), .ZN(n572) );
  NAND2_X1 U122 ( .A1(\mem[3][13] ), .A2(n751), .ZN(n737) );
  OAI21_X1 U123 ( .B1(n471), .B2(n751), .A(n736), .ZN(n571) );
  NAND2_X1 U124 ( .A1(\mem[3][14] ), .A2(n751), .ZN(n736) );
  OAI21_X1 U125 ( .B1(n470), .B2(n751), .A(n735), .ZN(n570) );
  NAND2_X1 U126 ( .A1(\mem[3][15] ), .A2(n459), .ZN(n735) );
  OAI21_X1 U127 ( .B1(n469), .B2(n751), .A(n734), .ZN(n569) );
  NAND2_X1 U128 ( .A1(\mem[3][16] ), .A2(n751), .ZN(n734) );
  OAI21_X1 U129 ( .B1(n468), .B2(n751), .A(n733), .ZN(n568) );
  NAND2_X1 U130 ( .A1(\mem[3][17] ), .A2(n751), .ZN(n733) );
  OAI21_X1 U131 ( .B1(n467), .B2(n751), .A(n732), .ZN(n567) );
  NAND2_X1 U132 ( .A1(\mem[3][18] ), .A2(n751), .ZN(n732) );
  OAI21_X1 U133 ( .B1(n466), .B2(n751), .A(n731), .ZN(n566) );
  NAND2_X1 U134 ( .A1(\mem[3][19] ), .A2(n459), .ZN(n731) );
  OAI21_X1 U135 ( .B1(n485), .B2(n730), .A(n729), .ZN(n565) );
  NAND2_X1 U136 ( .A1(\mem[4][0] ), .A2(n730), .ZN(n729) );
  OAI21_X1 U137 ( .B1(n484), .B2(n458), .A(n728), .ZN(n564) );
  NAND2_X1 U138 ( .A1(\mem[4][1] ), .A2(n730), .ZN(n728) );
  OAI21_X1 U139 ( .B1(n483), .B2(n458), .A(n727), .ZN(n563) );
  NAND2_X1 U140 ( .A1(\mem[4][2] ), .A2(n730), .ZN(n727) );
  OAI21_X1 U141 ( .B1(n482), .B2(n458), .A(n726), .ZN(n562) );
  NAND2_X1 U142 ( .A1(\mem[4][3] ), .A2(n730), .ZN(n726) );
  OAI21_X1 U143 ( .B1(n481), .B2(n458), .A(n725), .ZN(n561) );
  NAND2_X1 U144 ( .A1(\mem[4][4] ), .A2(n730), .ZN(n725) );
  OAI21_X1 U145 ( .B1(n480), .B2(n458), .A(n724), .ZN(n560) );
  NAND2_X1 U146 ( .A1(\mem[4][5] ), .A2(n730), .ZN(n724) );
  OAI21_X1 U147 ( .B1(n479), .B2(n458), .A(n723), .ZN(n559) );
  NAND2_X1 U148 ( .A1(\mem[4][6] ), .A2(n730), .ZN(n723) );
  OAI21_X1 U149 ( .B1(n478), .B2(n458), .A(n722), .ZN(n558) );
  NAND2_X1 U150 ( .A1(\mem[4][7] ), .A2(n730), .ZN(n722) );
  OAI21_X1 U151 ( .B1(n477), .B2(n458), .A(n721), .ZN(n557) );
  NAND2_X1 U152 ( .A1(\mem[4][8] ), .A2(n730), .ZN(n721) );
  OAI21_X1 U153 ( .B1(n476), .B2(n730), .A(n720), .ZN(n556) );
  NAND2_X1 U154 ( .A1(\mem[4][9] ), .A2(n730), .ZN(n720) );
  OAI21_X1 U155 ( .B1(n475), .B2(n458), .A(n719), .ZN(n555) );
  NAND2_X1 U156 ( .A1(\mem[4][10] ), .A2(n730), .ZN(n719) );
  OAI21_X1 U157 ( .B1(n474), .B2(n458), .A(n718), .ZN(n554) );
  NAND2_X1 U158 ( .A1(\mem[4][11] ), .A2(n730), .ZN(n718) );
  OAI21_X1 U159 ( .B1(n473), .B2(n730), .A(n717), .ZN(n553) );
  NAND2_X1 U160 ( .A1(\mem[4][12] ), .A2(n730), .ZN(n717) );
  OAI21_X1 U161 ( .B1(n472), .B2(n458), .A(n716), .ZN(n552) );
  NAND2_X1 U162 ( .A1(\mem[4][13] ), .A2(n730), .ZN(n716) );
  OAI21_X1 U163 ( .B1(n471), .B2(n730), .A(n715), .ZN(n551) );
  NAND2_X1 U164 ( .A1(\mem[4][14] ), .A2(n730), .ZN(n715) );
  OAI21_X1 U165 ( .B1(n470), .B2(n458), .A(n714), .ZN(n550) );
  NAND2_X1 U166 ( .A1(\mem[4][15] ), .A2(n730), .ZN(n714) );
  OAI21_X1 U167 ( .B1(n469), .B2(n458), .A(n713), .ZN(n549) );
  NAND2_X1 U168 ( .A1(\mem[4][16] ), .A2(n730), .ZN(n713) );
  OAI21_X1 U169 ( .B1(n468), .B2(n458), .A(n712), .ZN(n548) );
  NAND2_X1 U170 ( .A1(\mem[4][17] ), .A2(n730), .ZN(n712) );
  OAI21_X1 U171 ( .B1(n467), .B2(n458), .A(n711), .ZN(n547) );
  NAND2_X1 U172 ( .A1(\mem[4][18] ), .A2(n730), .ZN(n711) );
  OAI21_X1 U173 ( .B1(n466), .B2(n458), .A(n710), .ZN(n546) );
  NAND2_X1 U174 ( .A1(\mem[4][19] ), .A2(n730), .ZN(n710) );
  OAI21_X1 U175 ( .B1(n485), .B2(n708), .A(n707), .ZN(n545) );
  NAND2_X1 U176 ( .A1(\mem[5][0] ), .A2(n708), .ZN(n707) );
  OAI21_X1 U177 ( .B1(n484), .B2(n708), .A(n706), .ZN(n544) );
  NAND2_X1 U178 ( .A1(\mem[5][1] ), .A2(n708), .ZN(n706) );
  OAI21_X1 U179 ( .B1(n483), .B2(n708), .A(n705), .ZN(n543) );
  NAND2_X1 U180 ( .A1(\mem[5][2] ), .A2(n708), .ZN(n705) );
  OAI21_X1 U181 ( .B1(n482), .B2(n457), .A(n704), .ZN(n542) );
  NAND2_X1 U182 ( .A1(\mem[5][3] ), .A2(n457), .ZN(n704) );
  OAI21_X1 U183 ( .B1(n481), .B2(n708), .A(n703), .ZN(n541) );
  NAND2_X1 U184 ( .A1(\mem[5][4] ), .A2(n457), .ZN(n703) );
  OAI21_X1 U185 ( .B1(n480), .B2(n708), .A(n702), .ZN(n540) );
  NAND2_X1 U186 ( .A1(\mem[5][5] ), .A2(n708), .ZN(n702) );
  OAI21_X1 U187 ( .B1(n479), .B2(n708), .A(n701), .ZN(n539) );
  NAND2_X1 U188 ( .A1(\mem[5][6] ), .A2(n708), .ZN(n701) );
  OAI21_X1 U189 ( .B1(n478), .B2(n457), .A(n700), .ZN(n538) );
  NAND2_X1 U190 ( .A1(\mem[5][7] ), .A2(n708), .ZN(n700) );
  OAI21_X1 U191 ( .B1(n477), .B2(n457), .A(n699), .ZN(n537) );
  NAND2_X1 U192 ( .A1(\mem[5][8] ), .A2(n708), .ZN(n699) );
  OAI21_X1 U193 ( .B1(n476), .B2(n457), .A(n698), .ZN(n536) );
  NAND2_X1 U194 ( .A1(\mem[5][9] ), .A2(n708), .ZN(n698) );
  OAI21_X1 U195 ( .B1(n475), .B2(n457), .A(n697), .ZN(n535) );
  NAND2_X1 U196 ( .A1(\mem[5][10] ), .A2(n708), .ZN(n697) );
  OAI21_X1 U197 ( .B1(n474), .B2(n457), .A(n696), .ZN(n534) );
  NAND2_X1 U198 ( .A1(\mem[5][11] ), .A2(n708), .ZN(n696) );
  OAI21_X1 U199 ( .B1(n473), .B2(n708), .A(n695), .ZN(n533) );
  NAND2_X1 U200 ( .A1(\mem[5][12] ), .A2(n457), .ZN(n695) );
  OAI21_X1 U201 ( .B1(n472), .B2(n708), .A(n694), .ZN(n532) );
  NAND2_X1 U202 ( .A1(\mem[5][13] ), .A2(n457), .ZN(n694) );
  OAI21_X1 U203 ( .B1(n471), .B2(n708), .A(n693), .ZN(n531) );
  NAND2_X1 U204 ( .A1(\mem[5][14] ), .A2(n457), .ZN(n693) );
  OAI21_X1 U205 ( .B1(n470), .B2(n708), .A(n692), .ZN(n530) );
  NAND2_X1 U206 ( .A1(\mem[5][15] ), .A2(n457), .ZN(n692) );
  OAI21_X1 U207 ( .B1(n469), .B2(n708), .A(n691), .ZN(n529) );
  NAND2_X1 U208 ( .A1(\mem[5][16] ), .A2(n457), .ZN(n691) );
  OAI21_X1 U209 ( .B1(n468), .B2(n708), .A(n690), .ZN(n528) );
  NAND2_X1 U210 ( .A1(\mem[5][17] ), .A2(n457), .ZN(n690) );
  OAI21_X1 U211 ( .B1(n467), .B2(n708), .A(n689), .ZN(n527) );
  NAND2_X1 U212 ( .A1(\mem[5][18] ), .A2(n457), .ZN(n689) );
  OAI21_X1 U213 ( .B1(n466), .B2(n708), .A(n688), .ZN(n526) );
  NAND2_X1 U214 ( .A1(\mem[5][19] ), .A2(n457), .ZN(n688) );
  OAI21_X1 U215 ( .B1(n485), .B2(n687), .A(n686), .ZN(n525) );
  NAND2_X1 U216 ( .A1(\mem[6][0] ), .A2(n456), .ZN(n686) );
  OAI21_X1 U217 ( .B1(n484), .B2(n687), .A(n685), .ZN(n524) );
  NAND2_X1 U218 ( .A1(\mem[6][1] ), .A2(n456), .ZN(n685) );
  OAI21_X1 U219 ( .B1(n483), .B2(n687), .A(n684), .ZN(n523) );
  NAND2_X1 U220 ( .A1(\mem[6][2] ), .A2(n456), .ZN(n684) );
  OAI21_X1 U221 ( .B1(n482), .B2(n687), .A(n683), .ZN(n522) );
  NAND2_X1 U222 ( .A1(\mem[6][3] ), .A2(n456), .ZN(n683) );
  OAI21_X1 U223 ( .B1(n481), .B2(n456), .A(n682), .ZN(n521) );
  NAND2_X1 U224 ( .A1(\mem[6][4] ), .A2(n456), .ZN(n682) );
  OAI21_X1 U225 ( .B1(n480), .B2(n687), .A(n681), .ZN(n520) );
  NAND2_X1 U226 ( .A1(\mem[6][5] ), .A2(n456), .ZN(n681) );
  OAI21_X1 U227 ( .B1(n479), .B2(n687), .A(n680), .ZN(n519) );
  NAND2_X1 U228 ( .A1(\mem[6][6] ), .A2(n456), .ZN(n680) );
  OAI21_X1 U229 ( .B1(n478), .B2(n687), .A(n679), .ZN(n518) );
  NAND2_X1 U230 ( .A1(\mem[6][7] ), .A2(n456), .ZN(n679) );
  OAI21_X1 U231 ( .B1(n477), .B2(n687), .A(n678), .ZN(n517) );
  NAND2_X1 U232 ( .A1(\mem[6][8] ), .A2(n456), .ZN(n678) );
  OAI21_X1 U233 ( .B1(n476), .B2(n687), .A(n677), .ZN(n516) );
  NAND2_X1 U234 ( .A1(\mem[6][9] ), .A2(n456), .ZN(n677) );
  OAI21_X1 U235 ( .B1(n475), .B2(n687), .A(n676), .ZN(n515) );
  NAND2_X1 U236 ( .A1(\mem[6][10] ), .A2(n456), .ZN(n676) );
  OAI21_X1 U237 ( .B1(n474), .B2(n687), .A(n675), .ZN(n514) );
  NAND2_X1 U238 ( .A1(\mem[6][11] ), .A2(n456), .ZN(n675) );
  OAI21_X1 U239 ( .B1(n473), .B2(n687), .A(n674), .ZN(n513) );
  NAND2_X1 U240 ( .A1(\mem[6][12] ), .A2(n687), .ZN(n674) );
  OAI21_X1 U241 ( .B1(n472), .B2(n456), .A(n673), .ZN(n512) );
  NAND2_X1 U242 ( .A1(\mem[6][13] ), .A2(n687), .ZN(n673) );
  OAI21_X1 U243 ( .B1(n471), .B2(n456), .A(n672), .ZN(n511) );
  NAND2_X1 U244 ( .A1(\mem[6][14] ), .A2(n687), .ZN(n672) );
  OAI21_X1 U245 ( .B1(n470), .B2(n687), .A(n671), .ZN(n510) );
  NAND2_X1 U246 ( .A1(\mem[6][15] ), .A2(n687), .ZN(n671) );
  OAI21_X1 U247 ( .B1(n469), .B2(n687), .A(n670), .ZN(n509) );
  NAND2_X1 U248 ( .A1(\mem[6][16] ), .A2(n687), .ZN(n670) );
  OAI21_X1 U249 ( .B1(n468), .B2(n687), .A(n669), .ZN(n508) );
  NAND2_X1 U250 ( .A1(\mem[6][17] ), .A2(n687), .ZN(n669) );
  OAI21_X1 U251 ( .B1(n467), .B2(n687), .A(n668), .ZN(n507) );
  NAND2_X1 U252 ( .A1(\mem[6][18] ), .A2(n687), .ZN(n668) );
  OAI21_X1 U253 ( .B1(n466), .B2(n687), .A(n667), .ZN(n506) );
  NAND2_X1 U254 ( .A1(\mem[6][19] ), .A2(n456), .ZN(n667) );
  OAI21_X1 U255 ( .B1(n485), .B2(n455), .A(n665), .ZN(n505) );
  NAND2_X1 U256 ( .A1(\mem[7][0] ), .A2(n455), .ZN(n665) );
  OAI21_X1 U257 ( .B1(n484), .B2(n455), .A(n664), .ZN(n504) );
  NAND2_X1 U258 ( .A1(\mem[7][1] ), .A2(n455), .ZN(n664) );
  OAI21_X1 U259 ( .B1(n483), .B2(n455), .A(n663), .ZN(n503) );
  NAND2_X1 U260 ( .A1(\mem[7][2] ), .A2(n666), .ZN(n663) );
  OAI21_X1 U261 ( .B1(n482), .B2(n666), .A(n662), .ZN(n502) );
  NAND2_X1 U262 ( .A1(\mem[7][3] ), .A2(n455), .ZN(n662) );
  OAI21_X1 U263 ( .B1(n481), .B2(n666), .A(n661), .ZN(n501) );
  NAND2_X1 U264 ( .A1(\mem[7][4] ), .A2(n666), .ZN(n661) );
  OAI21_X1 U265 ( .B1(n480), .B2(n666), .A(n660), .ZN(n500) );
  NAND2_X1 U266 ( .A1(\mem[7][5] ), .A2(n666), .ZN(n660) );
  OAI21_X1 U267 ( .B1(n479), .B2(n666), .A(n659), .ZN(n499) );
  NAND2_X1 U268 ( .A1(\mem[7][6] ), .A2(n666), .ZN(n659) );
  OAI21_X1 U269 ( .B1(n478), .B2(n666), .A(n658), .ZN(n498) );
  NAND2_X1 U270 ( .A1(\mem[7][7] ), .A2(n666), .ZN(n658) );
  OAI21_X1 U271 ( .B1(n477), .B2(n666), .A(n657), .ZN(n497) );
  NAND2_X1 U272 ( .A1(\mem[7][8] ), .A2(n666), .ZN(n657) );
  OAI21_X1 U273 ( .B1(n476), .B2(n455), .A(n656), .ZN(n496) );
  NAND2_X1 U274 ( .A1(\mem[7][9] ), .A2(n666), .ZN(n656) );
  OAI21_X1 U275 ( .B1(n475), .B2(n666), .A(n655), .ZN(n495) );
  NAND2_X1 U276 ( .A1(\mem[7][10] ), .A2(n666), .ZN(n655) );
  OAI21_X1 U277 ( .B1(n474), .B2(n666), .A(n654), .ZN(n494) );
  NAND2_X1 U278 ( .A1(\mem[7][11] ), .A2(n666), .ZN(n654) );
  OAI21_X1 U279 ( .B1(n473), .B2(n455), .A(n653), .ZN(n493) );
  NAND2_X1 U280 ( .A1(\mem[7][12] ), .A2(n455), .ZN(n653) );
  OAI21_X1 U281 ( .B1(n472), .B2(n455), .A(n652), .ZN(n492) );
  NAND2_X1 U282 ( .A1(\mem[7][13] ), .A2(n455), .ZN(n652) );
  OAI21_X1 U283 ( .B1(n471), .B2(n455), .A(n651), .ZN(n491) );
  NAND2_X1 U284 ( .A1(\mem[7][14] ), .A2(n455), .ZN(n651) );
  OAI21_X1 U285 ( .B1(n470), .B2(n666), .A(n650), .ZN(n490) );
  NAND2_X1 U286 ( .A1(\mem[7][15] ), .A2(n455), .ZN(n650) );
  OAI21_X1 U287 ( .B1(n469), .B2(n666), .A(n649), .ZN(n489) );
  NAND2_X1 U288 ( .A1(\mem[7][16] ), .A2(n455), .ZN(n649) );
  OAI21_X1 U289 ( .B1(n468), .B2(n666), .A(n648), .ZN(n488) );
  NAND2_X1 U290 ( .A1(\mem[7][17] ), .A2(n455), .ZN(n648) );
  OAI21_X1 U291 ( .B1(n467), .B2(n455), .A(n647), .ZN(n487) );
  NAND2_X1 U292 ( .A1(\mem[7][18] ), .A2(n455), .ZN(n647) );
  OAI21_X1 U293 ( .B1(n466), .B2(n455), .A(n646), .ZN(n486) );
  NAND2_X1 U294 ( .A1(\mem[7][19] ), .A2(n455), .ZN(n646) );
  OAI21_X1 U295 ( .B1(n815), .B2(n483), .A(n812), .ZN(n643) );
  NAND2_X1 U296 ( .A1(\mem[0][2] ), .A2(n462), .ZN(n812) );
  OAI21_X1 U297 ( .B1(n815), .B2(n482), .A(n811), .ZN(n642) );
  NAND2_X1 U298 ( .A1(\mem[0][3] ), .A2(n462), .ZN(n811) );
  OAI21_X1 U299 ( .B1(n815), .B2(n481), .A(n810), .ZN(n641) );
  NAND2_X1 U300 ( .A1(\mem[0][4] ), .A2(n462), .ZN(n810) );
  OAI21_X1 U301 ( .B1(n815), .B2(n480), .A(n809), .ZN(n640) );
  NAND2_X1 U302 ( .A1(\mem[0][5] ), .A2(n462), .ZN(n809) );
  OAI21_X1 U303 ( .B1(n815), .B2(n479), .A(n808), .ZN(n639) );
  NAND2_X1 U304 ( .A1(\mem[0][6] ), .A2(n462), .ZN(n808) );
  OAI21_X1 U305 ( .B1(n815), .B2(n478), .A(n807), .ZN(n638) );
  NAND2_X1 U306 ( .A1(\mem[0][7] ), .A2(n462), .ZN(n807) );
  OAI21_X1 U307 ( .B1(n815), .B2(n477), .A(n806), .ZN(n637) );
  NAND2_X1 U308 ( .A1(\mem[0][8] ), .A2(n462), .ZN(n806) );
  OAI21_X1 U309 ( .B1(n815), .B2(n476), .A(n805), .ZN(n636) );
  NAND2_X1 U310 ( .A1(\mem[0][9] ), .A2(n462), .ZN(n805) );
  OAI21_X1 U311 ( .B1(n815), .B2(n475), .A(n804), .ZN(n635) );
  NAND2_X1 U312 ( .A1(\mem[0][10] ), .A2(n462), .ZN(n804) );
  OAI21_X1 U313 ( .B1(n815), .B2(n474), .A(n803), .ZN(n634) );
  NAND2_X1 U314 ( .A1(\mem[0][11] ), .A2(n462), .ZN(n803) );
  OAI21_X1 U315 ( .B1(n815), .B2(n473), .A(n802), .ZN(n633) );
  NAND2_X1 U316 ( .A1(\mem[0][12] ), .A2(n815), .ZN(n802) );
  OAI21_X1 U317 ( .B1(n815), .B2(n472), .A(n801), .ZN(n632) );
  NAND2_X1 U318 ( .A1(\mem[0][13] ), .A2(n815), .ZN(n801) );
  OAI21_X1 U319 ( .B1(n462), .B2(n471), .A(n800), .ZN(n631) );
  NAND2_X1 U320 ( .A1(\mem[0][14] ), .A2(n815), .ZN(n800) );
  OAI21_X1 U321 ( .B1(n815), .B2(n470), .A(n799), .ZN(n630) );
  NAND2_X1 U322 ( .A1(\mem[0][15] ), .A2(n462), .ZN(n799) );
  OAI21_X1 U323 ( .B1(n815), .B2(n469), .A(n798), .ZN(n629) );
  NAND2_X1 U324 ( .A1(\mem[0][16] ), .A2(n815), .ZN(n798) );
  OAI21_X1 U325 ( .B1(n815), .B2(n468), .A(n797), .ZN(n628) );
  NAND2_X1 U326 ( .A1(\mem[0][17] ), .A2(n815), .ZN(n797) );
  OAI21_X1 U327 ( .B1(n815), .B2(n467), .A(n796), .ZN(n627) );
  NAND2_X1 U328 ( .A1(\mem[0][18] ), .A2(n815), .ZN(n796) );
  OAI21_X1 U329 ( .B1(n462), .B2(n485), .A(n814), .ZN(n645) );
  NAND2_X1 U330 ( .A1(\mem[0][0] ), .A2(n462), .ZN(n814) );
  OAI21_X1 U331 ( .B1(n815), .B2(n484), .A(n813), .ZN(n644) );
  NAND2_X1 U332 ( .A1(\mem[0][1] ), .A2(n462), .ZN(n813) );
  OAI21_X1 U333 ( .B1(n815), .B2(n466), .A(n795), .ZN(n626) );
  NAND2_X1 U334 ( .A1(\mem[0][19] ), .A2(n462), .ZN(n795) );
  NOR2_X1 U335 ( .A1(n465), .A2(N12), .ZN(n794) );
  INV_X1 U336 ( .A(wr_en), .ZN(n465) );
  INV_X1 U337 ( .A(N10), .ZN(n463) );
  INV_X1 U338 ( .A(N11), .ZN(n464) );
  INV_X1 U339 ( .A(data_in[0]), .ZN(n485) );
  INV_X1 U340 ( .A(data_in[1]), .ZN(n484) );
  INV_X1 U341 ( .A(data_in[2]), .ZN(n483) );
  INV_X1 U342 ( .A(data_in[3]), .ZN(n482) );
  INV_X1 U343 ( .A(data_in[4]), .ZN(n481) );
  INV_X1 U344 ( .A(data_in[5]), .ZN(n480) );
  INV_X1 U345 ( .A(data_in[6]), .ZN(n479) );
  INV_X1 U346 ( .A(data_in[7]), .ZN(n478) );
  INV_X1 U347 ( .A(data_in[8]), .ZN(n477) );
  INV_X1 U356 ( .A(data_in[9]), .ZN(n476) );
  INV_X1 U357 ( .A(data_in[10]), .ZN(n475) );
  INV_X1 U358 ( .A(data_in[11]), .ZN(n474) );
  INV_X1 U359 ( .A(data_in[12]), .ZN(n473) );
  INV_X1 U360 ( .A(data_in[13]), .ZN(n472) );
  INV_X1 U361 ( .A(data_in[14]), .ZN(n471) );
  INV_X1 U362 ( .A(data_in[15]), .ZN(n470) );
  INV_X1 U363 ( .A(data_in[16]), .ZN(n469) );
  INV_X1 U364 ( .A(data_in[17]), .ZN(n468) );
  INV_X1 U365 ( .A(data_in[18]), .ZN(n467) );
  INV_X1 U366 ( .A(data_in[19]), .ZN(n466) );
  MUX2_X1 U367 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n452), .Z(n1) );
  MUX2_X1 U368 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n452), .Z(n2) );
  MUX2_X1 U369 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U370 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n452), .Z(n4) );
  MUX2_X1 U371 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n452), .Z(n5) );
  MUX2_X1 U372 ( .A(n5), .B(n4), .S(N11), .Z(n6) );
  MUX2_X1 U373 ( .A(n6), .B(n3), .S(N12), .Z(N32) );
  MUX2_X1 U374 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n452), .Z(n7) );
  MUX2_X1 U375 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n452), .Z(n8) );
  MUX2_X1 U376 ( .A(n8), .B(n7), .S(N11), .Z(n9) );
  MUX2_X1 U377 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n452), .Z(n10) );
  MUX2_X1 U378 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n452), .Z(n11) );
  MUX2_X1 U379 ( .A(n11), .B(n10), .S(N11), .Z(n12) );
  MUX2_X1 U380 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n453), .Z(n13) );
  MUX2_X1 U381 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n453), .Z(n14) );
  MUX2_X1 U382 ( .A(n14), .B(n13), .S(N11), .Z(n15) );
  MUX2_X1 U383 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n453), .Z(n16) );
  MUX2_X1 U384 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n453), .Z(n17) );
  MUX2_X1 U385 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U386 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n453), .Z(n19) );
  MUX2_X1 U387 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n453), .Z(n20) );
  MUX2_X1 U388 ( .A(n20), .B(n19), .S(N11), .Z(n21) );
  MUX2_X1 U389 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n453), .Z(n22) );
  MUX2_X1 U390 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n453), .Z(n23) );
  MUX2_X1 U391 ( .A(n23), .B(n22), .S(N11), .Z(n354) );
  MUX2_X1 U392 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n453), .Z(n355) );
  MUX2_X1 U393 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n453), .Z(n356) );
  MUX2_X1 U394 ( .A(n356), .B(n355), .S(N11), .Z(n357) );
  MUX2_X1 U395 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n453), .Z(n358) );
  MUX2_X1 U396 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n453), .Z(n359) );
  MUX2_X1 U397 ( .A(n359), .B(n358), .S(N11), .Z(n360) );
  MUX2_X1 U398 ( .A(n360), .B(n357), .S(N12), .Z(N28) );
  MUX2_X1 U399 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n452), .Z(n361) );
  MUX2_X1 U400 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(N10), .Z(n362) );
  MUX2_X1 U401 ( .A(n362), .B(n361), .S(N11), .Z(n363) );
  MUX2_X1 U402 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n364) );
  MUX2_X1 U403 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(N10), .Z(n365) );
  MUX2_X1 U404 ( .A(n365), .B(n364), .S(N11), .Z(n366) );
  MUX2_X1 U405 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n454), .Z(n367) );
  MUX2_X1 U406 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n453), .Z(n368) );
  MUX2_X1 U407 ( .A(n368), .B(n367), .S(n451), .Z(n369) );
  MUX2_X1 U408 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n454), .Z(n370) );
  MUX2_X1 U409 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n452), .Z(n371) );
  MUX2_X1 U410 ( .A(n371), .B(n370), .S(N11), .Z(n372) );
  MUX2_X1 U411 ( .A(n372), .B(n369), .S(N12), .Z(N26) );
  MUX2_X1 U412 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n373) );
  MUX2_X1 U413 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n374) );
  MUX2_X1 U414 ( .A(n374), .B(n373), .S(N11), .Z(n375) );
  MUX2_X1 U415 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n376) );
  MUX2_X1 U416 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n377) );
  MUX2_X1 U417 ( .A(n377), .B(n376), .S(N11), .Z(n378) );
  MUX2_X1 U418 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n453), .Z(n379) );
  MUX2_X1 U419 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n454), .Z(n380) );
  MUX2_X1 U420 ( .A(n380), .B(n379), .S(n451), .Z(n381) );
  MUX2_X1 U421 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n453), .Z(n382) );
  MUX2_X1 U422 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n453), .Z(n383) );
  MUX2_X1 U423 ( .A(n383), .B(n382), .S(n451), .Z(n384) );
  MUX2_X1 U424 ( .A(n384), .B(n381), .S(N12), .Z(N24) );
  MUX2_X1 U425 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n453), .Z(n385) );
  MUX2_X1 U426 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(N10), .Z(n386) );
  MUX2_X1 U427 ( .A(n386), .B(n385), .S(n451), .Z(n387) );
  MUX2_X1 U428 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n454), .Z(n388) );
  MUX2_X1 U429 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n453), .Z(n389) );
  MUX2_X1 U430 ( .A(n389), .B(n388), .S(n451), .Z(n390) );
  MUX2_X1 U431 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n454), .Z(n391) );
  MUX2_X1 U432 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n452), .Z(n392) );
  MUX2_X1 U433 ( .A(n392), .B(n391), .S(n451), .Z(n393) );
  MUX2_X1 U434 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n452), .Z(n394) );
  MUX2_X1 U435 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n452), .Z(n395) );
  MUX2_X1 U436 ( .A(n395), .B(n394), .S(n451), .Z(n396) );
  MUX2_X1 U437 ( .A(n396), .B(n393), .S(N12), .Z(N22) );
  MUX2_X1 U438 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(N10), .Z(n397) );
  MUX2_X1 U439 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n453), .Z(n398) );
  MUX2_X1 U440 ( .A(n398), .B(n397), .S(n451), .Z(n399) );
  MUX2_X1 U441 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n452), .Z(n400) );
  MUX2_X1 U442 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n452), .Z(n401) );
  MUX2_X1 U443 ( .A(n401), .B(n400), .S(n451), .Z(n402) );
  MUX2_X1 U444 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n452), .Z(n403) );
  MUX2_X1 U445 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n453), .Z(n404) );
  MUX2_X1 U446 ( .A(n404), .B(n403), .S(n451), .Z(n405) );
  MUX2_X1 U447 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n452), .Z(n406) );
  MUX2_X1 U448 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n454), .Z(n407) );
  MUX2_X1 U449 ( .A(n407), .B(n406), .S(n451), .Z(n408) );
  MUX2_X1 U450 ( .A(n408), .B(n405), .S(N12), .Z(N20) );
  MUX2_X1 U451 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n452), .Z(n409) );
  MUX2_X1 U452 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n454), .Z(n410) );
  MUX2_X1 U453 ( .A(n410), .B(n409), .S(n451), .Z(n411) );
  MUX2_X1 U454 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(N10), .Z(n412) );
  MUX2_X1 U455 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n453), .Z(n413) );
  MUX2_X1 U456 ( .A(n413), .B(n412), .S(n451), .Z(n414) );
  MUX2_X1 U457 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n452), .Z(n415) );
  MUX2_X1 U458 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n454), .Z(n416) );
  MUX2_X1 U459 ( .A(n416), .B(n415), .S(n451), .Z(n417) );
  MUX2_X1 U460 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n452), .Z(n418) );
  MUX2_X1 U461 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n454), .Z(n419) );
  MUX2_X1 U462 ( .A(n419), .B(n418), .S(n451), .Z(n420) );
  MUX2_X1 U463 ( .A(n420), .B(n417), .S(N12), .Z(N18) );
  MUX2_X1 U464 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n452), .Z(n421) );
  MUX2_X1 U465 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n453), .Z(n422) );
  MUX2_X1 U466 ( .A(n422), .B(n421), .S(n451), .Z(n423) );
  MUX2_X1 U467 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n454), .Z(n424) );
  MUX2_X1 U468 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(N10), .Z(n425) );
  MUX2_X1 U469 ( .A(n425), .B(n424), .S(n451), .Z(n426) );
  MUX2_X1 U470 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n452), .Z(n427) );
  MUX2_X1 U471 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n453), .Z(n428) );
  MUX2_X1 U472 ( .A(n428), .B(n427), .S(N11), .Z(n429) );
  MUX2_X1 U473 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n454), .Z(n430) );
  MUX2_X1 U474 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n452), .Z(n431) );
  MUX2_X1 U475 ( .A(n431), .B(n430), .S(n451), .Z(n432) );
  MUX2_X1 U476 ( .A(n432), .B(n429), .S(N12), .Z(N16) );
  MUX2_X1 U477 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n454), .Z(n433) );
  MUX2_X1 U478 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n454), .Z(n434) );
  MUX2_X1 U479 ( .A(n434), .B(n433), .S(n451), .Z(n435) );
  MUX2_X1 U480 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n454), .Z(n436) );
  MUX2_X1 U481 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n454), .Z(n437) );
  MUX2_X1 U482 ( .A(n437), .B(n436), .S(n451), .Z(n438) );
  MUX2_X1 U483 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n454), .Z(n439) );
  MUX2_X1 U484 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n454), .Z(n440) );
  MUX2_X1 U485 ( .A(n440), .B(n439), .S(N11), .Z(n441) );
  MUX2_X1 U486 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n454), .Z(n442) );
  MUX2_X1 U487 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n454), .Z(n443) );
  MUX2_X1 U488 ( .A(n443), .B(n442), .S(n451), .Z(n444) );
  MUX2_X1 U489 ( .A(n444), .B(n441), .S(N12), .Z(N14) );
  MUX2_X1 U490 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n454), .Z(n445) );
  MUX2_X1 U491 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n454), .Z(n446) );
  MUX2_X1 U492 ( .A(n446), .B(n445), .S(n451), .Z(n447) );
  MUX2_X1 U493 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n454), .Z(n448) );
  MUX2_X1 U494 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n454), .Z(n449) );
  MUX2_X1 U495 ( .A(n449), .B(n448), .S(n451), .Z(n450) );
  CLKBUF_X1 U496 ( .A(N10), .Z(n452) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE3_6 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N13, N14, N16, N18, N20, N22, N24, N26, N28, N30, N31,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[19]  ( .D(N13), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \data_out_reg[18]  ( .D(N14), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[16]  ( .D(N16), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N20), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N22), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[8]  ( .D(N24), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N26), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N28), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N30), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N31), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n486), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n487), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n488), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n489), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n490), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n491), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n492), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n493), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n494), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n495), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n496), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n497), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n498), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n499), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n500), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n501), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n502), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n503), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n504), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n505), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n506), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n507), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n508), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n509), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n510), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n511), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n512), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n513), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n514), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n515), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n516), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n517), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n518), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n519), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n520), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n521), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n522), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n523), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n524), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n525), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n526), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n527), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n528), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n529), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n530), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n531), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n532), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n533), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n534), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n535), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n536), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n537), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n538), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n539), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n540), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n541), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n542), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n543), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n544), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n545), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n546), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n547), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n548), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n549), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n550), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n551), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n552), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n553), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n554), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n555), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n556), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n557), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n558), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n559), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n560), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n561), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n562), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n563), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n564), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n565), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n566), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n567), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n568), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n569), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n570), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n571), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n572), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n573), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n574), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n575), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n576), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n577), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n578), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n579), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n580), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n581), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n582), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n583), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n584), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n585), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n586), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n587), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n588), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n589), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n590), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n591), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n592), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n593), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n594), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n595), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n596), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n597), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n598), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n599), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n600), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n601), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n602), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n603), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n604), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n605), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n606), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n607), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n608), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n609), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n610), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n611), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n612), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n613), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n614), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n615), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n616), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n617), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n618), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n619), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n620), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n621), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n622), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n623), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n624), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n625), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n626), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n627), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n628), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n629), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n630), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n631), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n632), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n633), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n634), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n635), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n636), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n637), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n638), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n639), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n640), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n641), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n642), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n643), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n644), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n645), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U348 ( .A1(n463), .A2(n464), .A3(n794), .ZN(n815) );
  NAND3_X1 U349 ( .A1(n794), .A2(n464), .A3(N10), .ZN(n793) );
  NAND3_X1 U350 ( .A1(n794), .A2(n463), .A3(N11), .ZN(n772) );
  NAND3_X1 U351 ( .A1(N10), .A2(n794), .A3(N11), .ZN(n751) );
  NAND3_X1 U352 ( .A1(n463), .A2(n464), .A3(n709), .ZN(n730) );
  NAND3_X1 U353 ( .A1(N10), .A2(n464), .A3(n709), .ZN(n708) );
  NAND3_X1 U354 ( .A1(N11), .A2(n463), .A3(n709), .ZN(n687) );
  NAND3_X1 U355 ( .A1(N11), .A2(N10), .A3(n709), .ZN(n666) );
  SDFF_X1 \data_out_reg[15]  ( .D(n426), .SI(n423), .SE(N12), .CK(clk), .Q(
        data_out[15]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n354), .SI(n21), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n390), .SI(n387), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n366), .SI(n363), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n378), .SI(n375), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[17]  ( .D(n438), .SI(n435), .SE(N12), .CK(clk), .Q(
        data_out[17]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n402), .SI(n399), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n414), .SI(n411), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n6), .SI(n3), .SE(N12), .CK(clk), .Q(
        data_out[0]) );
  BUF_X1 U3 ( .A(n793), .Z(n461) );
  BUF_X1 U4 ( .A(n751), .Z(n459) );
  BUF_X1 U5 ( .A(n666), .Z(n455) );
  BUF_X1 U6 ( .A(n815), .Z(n462) );
  BUF_X1 U7 ( .A(n772), .Z(n460) );
  BUF_X1 U8 ( .A(n730), .Z(n458) );
  BUF_X1 U9 ( .A(n708), .Z(n457) );
  BUF_X1 U10 ( .A(n687), .Z(n456) );
  BUF_X1 U11 ( .A(N10), .Z(n452) );
  BUF_X1 U12 ( .A(N10), .Z(n453) );
  BUF_X1 U13 ( .A(N10), .Z(n454) );
  BUF_X1 U14 ( .A(N11), .Z(n451) );
  NOR2_X1 U15 ( .A1(n465), .A2(N12), .ZN(n794) );
  INV_X1 U16 ( .A(wr_en), .ZN(n465) );
  AND2_X1 U17 ( .A1(N12), .A2(wr_en), .ZN(n709) );
  OAI21_X1 U18 ( .B1(n485), .B2(n461), .A(n792), .ZN(n625) );
  NAND2_X1 U19 ( .A1(\mem[1][0] ), .A2(n461), .ZN(n792) );
  OAI21_X1 U20 ( .B1(n484), .B2(n461), .A(n791), .ZN(n624) );
  NAND2_X1 U21 ( .A1(\mem[1][1] ), .A2(n461), .ZN(n791) );
  OAI21_X1 U22 ( .B1(n483), .B2(n461), .A(n790), .ZN(n623) );
  NAND2_X1 U23 ( .A1(\mem[1][2] ), .A2(n793), .ZN(n790) );
  OAI21_X1 U24 ( .B1(n482), .B2(n793), .A(n789), .ZN(n622) );
  NAND2_X1 U25 ( .A1(\mem[1][3] ), .A2(n461), .ZN(n789) );
  OAI21_X1 U26 ( .B1(n481), .B2(n793), .A(n788), .ZN(n621) );
  NAND2_X1 U27 ( .A1(\mem[1][4] ), .A2(n461), .ZN(n788) );
  OAI21_X1 U28 ( .B1(n480), .B2(n793), .A(n787), .ZN(n620) );
  NAND2_X1 U29 ( .A1(\mem[1][5] ), .A2(n793), .ZN(n787) );
  OAI21_X1 U30 ( .B1(n479), .B2(n793), .A(n786), .ZN(n619) );
  NAND2_X1 U31 ( .A1(\mem[1][6] ), .A2(n793), .ZN(n786) );
  OAI21_X1 U32 ( .B1(n478), .B2(n793), .A(n785), .ZN(n618) );
  NAND2_X1 U33 ( .A1(\mem[1][7] ), .A2(n793), .ZN(n785) );
  OAI21_X1 U34 ( .B1(n477), .B2(n793), .A(n784), .ZN(n617) );
  NAND2_X1 U35 ( .A1(\mem[1][8] ), .A2(n793), .ZN(n784) );
  OAI21_X1 U36 ( .B1(n476), .B2(n461), .A(n783), .ZN(n616) );
  NAND2_X1 U37 ( .A1(\mem[1][9] ), .A2(n793), .ZN(n783) );
  OAI21_X1 U38 ( .B1(n475), .B2(n793), .A(n782), .ZN(n615) );
  NAND2_X1 U39 ( .A1(\mem[1][10] ), .A2(n793), .ZN(n782) );
  OAI21_X1 U40 ( .B1(n474), .B2(n793), .A(n781), .ZN(n614) );
  NAND2_X1 U41 ( .A1(\mem[1][11] ), .A2(n793), .ZN(n781) );
  OAI21_X1 U42 ( .B1(n473), .B2(n461), .A(n780), .ZN(n613) );
  NAND2_X1 U43 ( .A1(\mem[1][12] ), .A2(n461), .ZN(n780) );
  OAI21_X1 U44 ( .B1(n472), .B2(n461), .A(n779), .ZN(n612) );
  NAND2_X1 U45 ( .A1(\mem[1][13] ), .A2(n461), .ZN(n779) );
  OAI21_X1 U46 ( .B1(n471), .B2(n461), .A(n778), .ZN(n611) );
  NAND2_X1 U47 ( .A1(\mem[1][14] ), .A2(n461), .ZN(n778) );
  OAI21_X1 U48 ( .B1(n470), .B2(n793), .A(n777), .ZN(n610) );
  NAND2_X1 U49 ( .A1(\mem[1][15] ), .A2(n461), .ZN(n777) );
  OAI21_X1 U50 ( .B1(n469), .B2(n793), .A(n776), .ZN(n609) );
  NAND2_X1 U51 ( .A1(\mem[1][16] ), .A2(n461), .ZN(n776) );
  OAI21_X1 U52 ( .B1(n468), .B2(n793), .A(n775), .ZN(n608) );
  NAND2_X1 U53 ( .A1(\mem[1][17] ), .A2(n461), .ZN(n775) );
  OAI21_X1 U54 ( .B1(n467), .B2(n461), .A(n774), .ZN(n607) );
  NAND2_X1 U55 ( .A1(\mem[1][18] ), .A2(n461), .ZN(n774) );
  OAI21_X1 U56 ( .B1(n466), .B2(n461), .A(n773), .ZN(n606) );
  NAND2_X1 U57 ( .A1(\mem[1][19] ), .A2(n461), .ZN(n773) );
  OAI21_X1 U58 ( .B1(n485), .B2(n772), .A(n771), .ZN(n605) );
  NAND2_X1 U59 ( .A1(\mem[2][0] ), .A2(n460), .ZN(n771) );
  OAI21_X1 U60 ( .B1(n484), .B2(n772), .A(n770), .ZN(n604) );
  NAND2_X1 U61 ( .A1(\mem[2][1] ), .A2(n460), .ZN(n770) );
  OAI21_X1 U62 ( .B1(n483), .B2(n772), .A(n769), .ZN(n603) );
  NAND2_X1 U63 ( .A1(\mem[2][2] ), .A2(n460), .ZN(n769) );
  OAI21_X1 U64 ( .B1(n482), .B2(n772), .A(n768), .ZN(n602) );
  NAND2_X1 U65 ( .A1(\mem[2][3] ), .A2(n460), .ZN(n768) );
  OAI21_X1 U66 ( .B1(n481), .B2(n460), .A(n767), .ZN(n601) );
  NAND2_X1 U67 ( .A1(\mem[2][4] ), .A2(n460), .ZN(n767) );
  OAI21_X1 U68 ( .B1(n480), .B2(n460), .A(n766), .ZN(n600) );
  NAND2_X1 U69 ( .A1(\mem[2][5] ), .A2(n460), .ZN(n766) );
  OAI21_X1 U70 ( .B1(n479), .B2(n772), .A(n765), .ZN(n599) );
  NAND2_X1 U71 ( .A1(\mem[2][6] ), .A2(n460), .ZN(n765) );
  OAI21_X1 U72 ( .B1(n478), .B2(n772), .A(n764), .ZN(n598) );
  NAND2_X1 U73 ( .A1(\mem[2][7] ), .A2(n460), .ZN(n764) );
  OAI21_X1 U74 ( .B1(n477), .B2(n772), .A(n763), .ZN(n597) );
  NAND2_X1 U75 ( .A1(\mem[2][8] ), .A2(n460), .ZN(n763) );
  OAI21_X1 U76 ( .B1(n476), .B2(n772), .A(n762), .ZN(n596) );
  NAND2_X1 U77 ( .A1(\mem[2][9] ), .A2(n460), .ZN(n762) );
  OAI21_X1 U78 ( .B1(n475), .B2(n772), .A(n761), .ZN(n595) );
  NAND2_X1 U79 ( .A1(\mem[2][10] ), .A2(n460), .ZN(n761) );
  OAI21_X1 U80 ( .B1(n474), .B2(n772), .A(n760), .ZN(n594) );
  NAND2_X1 U81 ( .A1(\mem[2][11] ), .A2(n460), .ZN(n760) );
  OAI21_X1 U82 ( .B1(n473), .B2(n772), .A(n759), .ZN(n593) );
  NAND2_X1 U83 ( .A1(\mem[2][12] ), .A2(n772), .ZN(n759) );
  OAI21_X1 U84 ( .B1(n472), .B2(n772), .A(n758), .ZN(n592) );
  NAND2_X1 U85 ( .A1(\mem[2][13] ), .A2(n772), .ZN(n758) );
  OAI21_X1 U86 ( .B1(n471), .B2(n772), .A(n757), .ZN(n591) );
  NAND2_X1 U87 ( .A1(\mem[2][14] ), .A2(n772), .ZN(n757) );
  OAI21_X1 U88 ( .B1(n470), .B2(n772), .A(n756), .ZN(n590) );
  NAND2_X1 U89 ( .A1(\mem[2][15] ), .A2(n460), .ZN(n756) );
  OAI21_X1 U90 ( .B1(n469), .B2(n772), .A(n755), .ZN(n589) );
  NAND2_X1 U91 ( .A1(\mem[2][16] ), .A2(n772), .ZN(n755) );
  OAI21_X1 U92 ( .B1(n468), .B2(n772), .A(n754), .ZN(n588) );
  NAND2_X1 U93 ( .A1(\mem[2][17] ), .A2(n772), .ZN(n754) );
  OAI21_X1 U94 ( .B1(n467), .B2(n772), .A(n753), .ZN(n587) );
  NAND2_X1 U95 ( .A1(\mem[2][18] ), .A2(n772), .ZN(n753) );
  OAI21_X1 U96 ( .B1(n466), .B2(n772), .A(n752), .ZN(n586) );
  NAND2_X1 U97 ( .A1(\mem[2][19] ), .A2(n460), .ZN(n752) );
  OAI21_X1 U98 ( .B1(n485), .B2(n459), .A(n750), .ZN(n585) );
  NAND2_X1 U99 ( .A1(\mem[3][0] ), .A2(n459), .ZN(n750) );
  OAI21_X1 U100 ( .B1(n484), .B2(n459), .A(n749), .ZN(n584) );
  NAND2_X1 U101 ( .A1(\mem[3][1] ), .A2(n459), .ZN(n749) );
  OAI21_X1 U102 ( .B1(n483), .B2(n459), .A(n748), .ZN(n583) );
  NAND2_X1 U103 ( .A1(\mem[3][2] ), .A2(n751), .ZN(n748) );
  OAI21_X1 U104 ( .B1(n482), .B2(n751), .A(n747), .ZN(n582) );
  NAND2_X1 U105 ( .A1(\mem[3][3] ), .A2(n459), .ZN(n747) );
  OAI21_X1 U106 ( .B1(n481), .B2(n751), .A(n746), .ZN(n581) );
  NAND2_X1 U107 ( .A1(\mem[3][4] ), .A2(n459), .ZN(n746) );
  OAI21_X1 U108 ( .B1(n480), .B2(n751), .A(n745), .ZN(n580) );
  NAND2_X1 U109 ( .A1(\mem[3][5] ), .A2(n751), .ZN(n745) );
  OAI21_X1 U110 ( .B1(n479), .B2(n751), .A(n744), .ZN(n579) );
  NAND2_X1 U111 ( .A1(\mem[3][6] ), .A2(n751), .ZN(n744) );
  OAI21_X1 U112 ( .B1(n478), .B2(n751), .A(n743), .ZN(n578) );
  NAND2_X1 U113 ( .A1(\mem[3][7] ), .A2(n751), .ZN(n743) );
  OAI21_X1 U114 ( .B1(n477), .B2(n751), .A(n742), .ZN(n577) );
  NAND2_X1 U115 ( .A1(\mem[3][8] ), .A2(n751), .ZN(n742) );
  OAI21_X1 U116 ( .B1(n476), .B2(n459), .A(n741), .ZN(n576) );
  NAND2_X1 U117 ( .A1(\mem[3][9] ), .A2(n751), .ZN(n741) );
  OAI21_X1 U118 ( .B1(n475), .B2(n751), .A(n740), .ZN(n575) );
  NAND2_X1 U119 ( .A1(\mem[3][10] ), .A2(n751), .ZN(n740) );
  OAI21_X1 U120 ( .B1(n474), .B2(n751), .A(n739), .ZN(n574) );
  NAND2_X1 U121 ( .A1(\mem[3][11] ), .A2(n751), .ZN(n739) );
  OAI21_X1 U122 ( .B1(n473), .B2(n459), .A(n738), .ZN(n573) );
  NAND2_X1 U123 ( .A1(\mem[3][12] ), .A2(n459), .ZN(n738) );
  OAI21_X1 U124 ( .B1(n472), .B2(n459), .A(n737), .ZN(n572) );
  NAND2_X1 U125 ( .A1(\mem[3][13] ), .A2(n459), .ZN(n737) );
  OAI21_X1 U126 ( .B1(n471), .B2(n459), .A(n736), .ZN(n571) );
  NAND2_X1 U127 ( .A1(\mem[3][14] ), .A2(n459), .ZN(n736) );
  OAI21_X1 U128 ( .B1(n470), .B2(n751), .A(n735), .ZN(n570) );
  NAND2_X1 U129 ( .A1(\mem[3][15] ), .A2(n459), .ZN(n735) );
  OAI21_X1 U130 ( .B1(n469), .B2(n751), .A(n734), .ZN(n569) );
  NAND2_X1 U131 ( .A1(\mem[3][16] ), .A2(n459), .ZN(n734) );
  OAI21_X1 U132 ( .B1(n468), .B2(n751), .A(n733), .ZN(n568) );
  NAND2_X1 U133 ( .A1(\mem[3][17] ), .A2(n459), .ZN(n733) );
  OAI21_X1 U134 ( .B1(n467), .B2(n459), .A(n732), .ZN(n567) );
  NAND2_X1 U135 ( .A1(\mem[3][18] ), .A2(n459), .ZN(n732) );
  OAI21_X1 U136 ( .B1(n466), .B2(n459), .A(n731), .ZN(n566) );
  NAND2_X1 U137 ( .A1(\mem[3][19] ), .A2(n459), .ZN(n731) );
  OAI21_X1 U138 ( .B1(n485), .B2(n730), .A(n729), .ZN(n565) );
  NAND2_X1 U139 ( .A1(\mem[4][0] ), .A2(n458), .ZN(n729) );
  OAI21_X1 U140 ( .B1(n484), .B2(n730), .A(n728), .ZN(n564) );
  NAND2_X1 U141 ( .A1(\mem[4][1] ), .A2(n458), .ZN(n728) );
  OAI21_X1 U142 ( .B1(n483), .B2(n730), .A(n727), .ZN(n563) );
  NAND2_X1 U143 ( .A1(\mem[4][2] ), .A2(n458), .ZN(n727) );
  OAI21_X1 U144 ( .B1(n482), .B2(n730), .A(n726), .ZN(n562) );
  NAND2_X1 U145 ( .A1(\mem[4][3] ), .A2(n458), .ZN(n726) );
  OAI21_X1 U146 ( .B1(n481), .B2(n458), .A(n725), .ZN(n561) );
  NAND2_X1 U147 ( .A1(\mem[4][4] ), .A2(n458), .ZN(n725) );
  OAI21_X1 U148 ( .B1(n480), .B2(n730), .A(n724), .ZN(n560) );
  NAND2_X1 U149 ( .A1(\mem[4][5] ), .A2(n458), .ZN(n724) );
  OAI21_X1 U150 ( .B1(n479), .B2(n730), .A(n723), .ZN(n559) );
  NAND2_X1 U151 ( .A1(\mem[4][6] ), .A2(n458), .ZN(n723) );
  OAI21_X1 U152 ( .B1(n478), .B2(n730), .A(n722), .ZN(n558) );
  NAND2_X1 U153 ( .A1(\mem[4][7] ), .A2(n458), .ZN(n722) );
  OAI21_X1 U154 ( .B1(n477), .B2(n730), .A(n721), .ZN(n557) );
  NAND2_X1 U155 ( .A1(\mem[4][8] ), .A2(n458), .ZN(n721) );
  OAI21_X1 U156 ( .B1(n476), .B2(n730), .A(n720), .ZN(n556) );
  NAND2_X1 U157 ( .A1(\mem[4][9] ), .A2(n458), .ZN(n720) );
  OAI21_X1 U158 ( .B1(n475), .B2(n730), .A(n719), .ZN(n555) );
  NAND2_X1 U159 ( .A1(\mem[4][10] ), .A2(n458), .ZN(n719) );
  OAI21_X1 U160 ( .B1(n474), .B2(n730), .A(n718), .ZN(n554) );
  NAND2_X1 U161 ( .A1(\mem[4][11] ), .A2(n458), .ZN(n718) );
  OAI21_X1 U162 ( .B1(n473), .B2(n730), .A(n717), .ZN(n553) );
  NAND2_X1 U163 ( .A1(\mem[4][12] ), .A2(n730), .ZN(n717) );
  OAI21_X1 U164 ( .B1(n472), .B2(n458), .A(n716), .ZN(n552) );
  NAND2_X1 U165 ( .A1(\mem[4][13] ), .A2(n730), .ZN(n716) );
  OAI21_X1 U166 ( .B1(n471), .B2(n458), .A(n715), .ZN(n551) );
  NAND2_X1 U167 ( .A1(\mem[4][14] ), .A2(n730), .ZN(n715) );
  OAI21_X1 U168 ( .B1(n470), .B2(n730), .A(n714), .ZN(n550) );
  NAND2_X1 U169 ( .A1(\mem[4][15] ), .A2(n730), .ZN(n714) );
  OAI21_X1 U170 ( .B1(n469), .B2(n730), .A(n713), .ZN(n549) );
  NAND2_X1 U171 ( .A1(\mem[4][16] ), .A2(n730), .ZN(n713) );
  OAI21_X1 U172 ( .B1(n468), .B2(n730), .A(n712), .ZN(n548) );
  NAND2_X1 U173 ( .A1(\mem[4][17] ), .A2(n730), .ZN(n712) );
  OAI21_X1 U174 ( .B1(n467), .B2(n730), .A(n711), .ZN(n547) );
  NAND2_X1 U175 ( .A1(\mem[4][18] ), .A2(n730), .ZN(n711) );
  OAI21_X1 U176 ( .B1(n466), .B2(n730), .A(n710), .ZN(n546) );
  NAND2_X1 U177 ( .A1(\mem[4][19] ), .A2(n458), .ZN(n710) );
  OAI21_X1 U178 ( .B1(n485), .B2(n708), .A(n707), .ZN(n545) );
  NAND2_X1 U179 ( .A1(\mem[5][0] ), .A2(n457), .ZN(n707) );
  OAI21_X1 U180 ( .B1(n484), .B2(n708), .A(n706), .ZN(n544) );
  NAND2_X1 U181 ( .A1(\mem[5][1] ), .A2(n457), .ZN(n706) );
  OAI21_X1 U182 ( .B1(n483), .B2(n708), .A(n705), .ZN(n543) );
  NAND2_X1 U183 ( .A1(\mem[5][2] ), .A2(n457), .ZN(n705) );
  OAI21_X1 U184 ( .B1(n482), .B2(n708), .A(n704), .ZN(n542) );
  NAND2_X1 U185 ( .A1(\mem[5][3] ), .A2(n457), .ZN(n704) );
  OAI21_X1 U186 ( .B1(n481), .B2(n457), .A(n703), .ZN(n541) );
  NAND2_X1 U187 ( .A1(\mem[5][4] ), .A2(n457), .ZN(n703) );
  OAI21_X1 U188 ( .B1(n480), .B2(n708), .A(n702), .ZN(n540) );
  NAND2_X1 U189 ( .A1(\mem[5][5] ), .A2(n457), .ZN(n702) );
  OAI21_X1 U190 ( .B1(n479), .B2(n708), .A(n701), .ZN(n539) );
  NAND2_X1 U191 ( .A1(\mem[5][6] ), .A2(n457), .ZN(n701) );
  OAI21_X1 U192 ( .B1(n478), .B2(n708), .A(n700), .ZN(n538) );
  NAND2_X1 U193 ( .A1(\mem[5][7] ), .A2(n457), .ZN(n700) );
  OAI21_X1 U194 ( .B1(n477), .B2(n708), .A(n699), .ZN(n537) );
  NAND2_X1 U195 ( .A1(\mem[5][8] ), .A2(n457), .ZN(n699) );
  OAI21_X1 U196 ( .B1(n476), .B2(n708), .A(n698), .ZN(n536) );
  NAND2_X1 U197 ( .A1(\mem[5][9] ), .A2(n457), .ZN(n698) );
  OAI21_X1 U198 ( .B1(n475), .B2(n708), .A(n697), .ZN(n535) );
  NAND2_X1 U199 ( .A1(\mem[5][10] ), .A2(n457), .ZN(n697) );
  OAI21_X1 U200 ( .B1(n474), .B2(n708), .A(n696), .ZN(n534) );
  NAND2_X1 U201 ( .A1(\mem[5][11] ), .A2(n457), .ZN(n696) );
  OAI21_X1 U202 ( .B1(n473), .B2(n708), .A(n695), .ZN(n533) );
  NAND2_X1 U203 ( .A1(\mem[5][12] ), .A2(n708), .ZN(n695) );
  OAI21_X1 U204 ( .B1(n472), .B2(n457), .A(n694), .ZN(n532) );
  NAND2_X1 U205 ( .A1(\mem[5][13] ), .A2(n708), .ZN(n694) );
  OAI21_X1 U206 ( .B1(n471), .B2(n457), .A(n693), .ZN(n531) );
  NAND2_X1 U207 ( .A1(\mem[5][14] ), .A2(n708), .ZN(n693) );
  OAI21_X1 U208 ( .B1(n470), .B2(n708), .A(n692), .ZN(n530) );
  NAND2_X1 U209 ( .A1(\mem[5][15] ), .A2(n708), .ZN(n692) );
  OAI21_X1 U210 ( .B1(n469), .B2(n708), .A(n691), .ZN(n529) );
  NAND2_X1 U211 ( .A1(\mem[5][16] ), .A2(n708), .ZN(n691) );
  OAI21_X1 U212 ( .B1(n468), .B2(n708), .A(n690), .ZN(n528) );
  NAND2_X1 U213 ( .A1(\mem[5][17] ), .A2(n708), .ZN(n690) );
  OAI21_X1 U214 ( .B1(n467), .B2(n708), .A(n689), .ZN(n527) );
  NAND2_X1 U215 ( .A1(\mem[5][18] ), .A2(n708), .ZN(n689) );
  OAI21_X1 U216 ( .B1(n466), .B2(n708), .A(n688), .ZN(n526) );
  NAND2_X1 U217 ( .A1(\mem[5][19] ), .A2(n457), .ZN(n688) );
  OAI21_X1 U218 ( .B1(n485), .B2(n687), .A(n686), .ZN(n525) );
  NAND2_X1 U219 ( .A1(\mem[6][0] ), .A2(n456), .ZN(n686) );
  OAI21_X1 U220 ( .B1(n484), .B2(n687), .A(n685), .ZN(n524) );
  NAND2_X1 U221 ( .A1(\mem[6][1] ), .A2(n456), .ZN(n685) );
  OAI21_X1 U222 ( .B1(n483), .B2(n687), .A(n684), .ZN(n523) );
  NAND2_X1 U223 ( .A1(\mem[6][2] ), .A2(n456), .ZN(n684) );
  OAI21_X1 U224 ( .B1(n482), .B2(n687), .A(n683), .ZN(n522) );
  NAND2_X1 U225 ( .A1(\mem[6][3] ), .A2(n456), .ZN(n683) );
  OAI21_X1 U226 ( .B1(n481), .B2(n456), .A(n682), .ZN(n521) );
  NAND2_X1 U227 ( .A1(\mem[6][4] ), .A2(n456), .ZN(n682) );
  OAI21_X1 U228 ( .B1(n480), .B2(n687), .A(n681), .ZN(n520) );
  NAND2_X1 U229 ( .A1(\mem[6][5] ), .A2(n456), .ZN(n681) );
  OAI21_X1 U230 ( .B1(n479), .B2(n687), .A(n680), .ZN(n519) );
  NAND2_X1 U231 ( .A1(\mem[6][6] ), .A2(n456), .ZN(n680) );
  OAI21_X1 U232 ( .B1(n478), .B2(n687), .A(n679), .ZN(n518) );
  NAND2_X1 U233 ( .A1(\mem[6][7] ), .A2(n456), .ZN(n679) );
  OAI21_X1 U234 ( .B1(n477), .B2(n687), .A(n678), .ZN(n517) );
  NAND2_X1 U235 ( .A1(\mem[6][8] ), .A2(n456), .ZN(n678) );
  OAI21_X1 U236 ( .B1(n476), .B2(n687), .A(n677), .ZN(n516) );
  NAND2_X1 U237 ( .A1(\mem[6][9] ), .A2(n456), .ZN(n677) );
  OAI21_X1 U238 ( .B1(n475), .B2(n687), .A(n676), .ZN(n515) );
  NAND2_X1 U239 ( .A1(\mem[6][10] ), .A2(n456), .ZN(n676) );
  OAI21_X1 U240 ( .B1(n474), .B2(n687), .A(n675), .ZN(n514) );
  NAND2_X1 U241 ( .A1(\mem[6][11] ), .A2(n456), .ZN(n675) );
  OAI21_X1 U242 ( .B1(n473), .B2(n687), .A(n674), .ZN(n513) );
  NAND2_X1 U243 ( .A1(\mem[6][12] ), .A2(n687), .ZN(n674) );
  OAI21_X1 U244 ( .B1(n472), .B2(n456), .A(n673), .ZN(n512) );
  NAND2_X1 U245 ( .A1(\mem[6][13] ), .A2(n687), .ZN(n673) );
  OAI21_X1 U246 ( .B1(n471), .B2(n456), .A(n672), .ZN(n511) );
  NAND2_X1 U247 ( .A1(\mem[6][14] ), .A2(n687), .ZN(n672) );
  OAI21_X1 U248 ( .B1(n470), .B2(n687), .A(n671), .ZN(n510) );
  NAND2_X1 U249 ( .A1(\mem[6][15] ), .A2(n687), .ZN(n671) );
  OAI21_X1 U250 ( .B1(n469), .B2(n687), .A(n670), .ZN(n509) );
  NAND2_X1 U251 ( .A1(\mem[6][16] ), .A2(n687), .ZN(n670) );
  OAI21_X1 U252 ( .B1(n468), .B2(n687), .A(n669), .ZN(n508) );
  NAND2_X1 U253 ( .A1(\mem[6][17] ), .A2(n687), .ZN(n669) );
  OAI21_X1 U254 ( .B1(n467), .B2(n687), .A(n668), .ZN(n507) );
  NAND2_X1 U255 ( .A1(\mem[6][18] ), .A2(n687), .ZN(n668) );
  OAI21_X1 U256 ( .B1(n466), .B2(n687), .A(n667), .ZN(n506) );
  NAND2_X1 U257 ( .A1(\mem[6][19] ), .A2(n456), .ZN(n667) );
  OAI21_X1 U258 ( .B1(n485), .B2(n666), .A(n665), .ZN(n505) );
  NAND2_X1 U259 ( .A1(\mem[7][0] ), .A2(n666), .ZN(n665) );
  OAI21_X1 U260 ( .B1(n484), .B2(n455), .A(n664), .ZN(n504) );
  NAND2_X1 U261 ( .A1(\mem[7][1] ), .A2(n666), .ZN(n664) );
  OAI21_X1 U262 ( .B1(n483), .B2(n455), .A(n663), .ZN(n503) );
  NAND2_X1 U263 ( .A1(\mem[7][2] ), .A2(n666), .ZN(n663) );
  OAI21_X1 U264 ( .B1(n482), .B2(n455), .A(n662), .ZN(n502) );
  NAND2_X1 U265 ( .A1(\mem[7][3] ), .A2(n666), .ZN(n662) );
  OAI21_X1 U266 ( .B1(n481), .B2(n455), .A(n661), .ZN(n501) );
  NAND2_X1 U267 ( .A1(\mem[7][4] ), .A2(n666), .ZN(n661) );
  OAI21_X1 U268 ( .B1(n480), .B2(n455), .A(n660), .ZN(n500) );
  NAND2_X1 U269 ( .A1(\mem[7][5] ), .A2(n666), .ZN(n660) );
  OAI21_X1 U270 ( .B1(n479), .B2(n455), .A(n659), .ZN(n499) );
  NAND2_X1 U271 ( .A1(\mem[7][6] ), .A2(n666), .ZN(n659) );
  OAI21_X1 U272 ( .B1(n478), .B2(n455), .A(n658), .ZN(n498) );
  NAND2_X1 U273 ( .A1(\mem[7][7] ), .A2(n666), .ZN(n658) );
  OAI21_X1 U274 ( .B1(n477), .B2(n455), .A(n657), .ZN(n497) );
  NAND2_X1 U275 ( .A1(\mem[7][8] ), .A2(n666), .ZN(n657) );
  OAI21_X1 U276 ( .B1(n476), .B2(n666), .A(n656), .ZN(n496) );
  NAND2_X1 U277 ( .A1(\mem[7][9] ), .A2(n666), .ZN(n656) );
  OAI21_X1 U278 ( .B1(n475), .B2(n455), .A(n655), .ZN(n495) );
  NAND2_X1 U279 ( .A1(\mem[7][10] ), .A2(n666), .ZN(n655) );
  OAI21_X1 U280 ( .B1(n474), .B2(n455), .A(n654), .ZN(n494) );
  NAND2_X1 U281 ( .A1(\mem[7][11] ), .A2(n666), .ZN(n654) );
  OAI21_X1 U282 ( .B1(n473), .B2(n666), .A(n653), .ZN(n493) );
  NAND2_X1 U283 ( .A1(\mem[7][12] ), .A2(n666), .ZN(n653) );
  OAI21_X1 U284 ( .B1(n472), .B2(n455), .A(n652), .ZN(n492) );
  NAND2_X1 U285 ( .A1(\mem[7][13] ), .A2(n666), .ZN(n652) );
  OAI21_X1 U286 ( .B1(n471), .B2(n666), .A(n651), .ZN(n491) );
  NAND2_X1 U287 ( .A1(\mem[7][14] ), .A2(n666), .ZN(n651) );
  OAI21_X1 U288 ( .B1(n470), .B2(n455), .A(n650), .ZN(n490) );
  NAND2_X1 U289 ( .A1(\mem[7][15] ), .A2(n666), .ZN(n650) );
  OAI21_X1 U290 ( .B1(n469), .B2(n455), .A(n649), .ZN(n489) );
  NAND2_X1 U291 ( .A1(\mem[7][16] ), .A2(n666), .ZN(n649) );
  OAI21_X1 U292 ( .B1(n468), .B2(n455), .A(n648), .ZN(n488) );
  NAND2_X1 U293 ( .A1(\mem[7][17] ), .A2(n666), .ZN(n648) );
  OAI21_X1 U294 ( .B1(n467), .B2(n455), .A(n647), .ZN(n487) );
  NAND2_X1 U295 ( .A1(\mem[7][18] ), .A2(n666), .ZN(n647) );
  OAI21_X1 U296 ( .B1(n466), .B2(n455), .A(n646), .ZN(n486) );
  NAND2_X1 U297 ( .A1(\mem[7][19] ), .A2(n666), .ZN(n646) );
  OAI21_X1 U298 ( .B1(n815), .B2(n483), .A(n812), .ZN(n643) );
  NAND2_X1 U299 ( .A1(\mem[0][2] ), .A2(n462), .ZN(n812) );
  OAI21_X1 U300 ( .B1(n815), .B2(n482), .A(n811), .ZN(n642) );
  NAND2_X1 U301 ( .A1(\mem[0][3] ), .A2(n462), .ZN(n811) );
  OAI21_X1 U302 ( .B1(n815), .B2(n481), .A(n810), .ZN(n641) );
  NAND2_X1 U303 ( .A1(\mem[0][4] ), .A2(n462), .ZN(n810) );
  OAI21_X1 U304 ( .B1(n815), .B2(n480), .A(n809), .ZN(n640) );
  NAND2_X1 U305 ( .A1(\mem[0][5] ), .A2(n462), .ZN(n809) );
  OAI21_X1 U306 ( .B1(n815), .B2(n479), .A(n808), .ZN(n639) );
  NAND2_X1 U307 ( .A1(\mem[0][6] ), .A2(n462), .ZN(n808) );
  OAI21_X1 U308 ( .B1(n815), .B2(n478), .A(n807), .ZN(n638) );
  NAND2_X1 U309 ( .A1(\mem[0][7] ), .A2(n462), .ZN(n807) );
  OAI21_X1 U310 ( .B1(n815), .B2(n477), .A(n806), .ZN(n637) );
  NAND2_X1 U311 ( .A1(\mem[0][8] ), .A2(n462), .ZN(n806) );
  OAI21_X1 U312 ( .B1(n815), .B2(n476), .A(n805), .ZN(n636) );
  NAND2_X1 U313 ( .A1(\mem[0][9] ), .A2(n462), .ZN(n805) );
  OAI21_X1 U314 ( .B1(n815), .B2(n475), .A(n804), .ZN(n635) );
  NAND2_X1 U315 ( .A1(\mem[0][10] ), .A2(n462), .ZN(n804) );
  OAI21_X1 U316 ( .B1(n815), .B2(n474), .A(n803), .ZN(n634) );
  NAND2_X1 U317 ( .A1(\mem[0][11] ), .A2(n462), .ZN(n803) );
  OAI21_X1 U318 ( .B1(n815), .B2(n473), .A(n802), .ZN(n633) );
  NAND2_X1 U319 ( .A1(\mem[0][12] ), .A2(n815), .ZN(n802) );
  OAI21_X1 U320 ( .B1(n815), .B2(n472), .A(n801), .ZN(n632) );
  NAND2_X1 U321 ( .A1(\mem[0][13] ), .A2(n815), .ZN(n801) );
  OAI21_X1 U322 ( .B1(n462), .B2(n471), .A(n800), .ZN(n631) );
  NAND2_X1 U323 ( .A1(\mem[0][14] ), .A2(n815), .ZN(n800) );
  OAI21_X1 U324 ( .B1(n815), .B2(n470), .A(n799), .ZN(n630) );
  NAND2_X1 U325 ( .A1(\mem[0][15] ), .A2(n462), .ZN(n799) );
  OAI21_X1 U326 ( .B1(n815), .B2(n469), .A(n798), .ZN(n629) );
  NAND2_X1 U327 ( .A1(\mem[0][16] ), .A2(n815), .ZN(n798) );
  OAI21_X1 U328 ( .B1(n815), .B2(n468), .A(n797), .ZN(n628) );
  NAND2_X1 U329 ( .A1(\mem[0][17] ), .A2(n815), .ZN(n797) );
  OAI21_X1 U330 ( .B1(n815), .B2(n467), .A(n796), .ZN(n627) );
  NAND2_X1 U331 ( .A1(\mem[0][18] ), .A2(n815), .ZN(n796) );
  OAI21_X1 U332 ( .B1(n462), .B2(n485), .A(n814), .ZN(n645) );
  NAND2_X1 U333 ( .A1(\mem[0][0] ), .A2(n462), .ZN(n814) );
  OAI21_X1 U334 ( .B1(n815), .B2(n484), .A(n813), .ZN(n644) );
  NAND2_X1 U335 ( .A1(\mem[0][1] ), .A2(n462), .ZN(n813) );
  OAI21_X1 U336 ( .B1(n815), .B2(n466), .A(n795), .ZN(n626) );
  NAND2_X1 U337 ( .A1(\mem[0][19] ), .A2(n462), .ZN(n795) );
  INV_X1 U338 ( .A(N10), .ZN(n463) );
  INV_X1 U339 ( .A(N11), .ZN(n464) );
  INV_X1 U340 ( .A(data_in[0]), .ZN(n485) );
  INV_X1 U341 ( .A(data_in[1]), .ZN(n484) );
  INV_X1 U342 ( .A(data_in[2]), .ZN(n483) );
  INV_X1 U343 ( .A(data_in[3]), .ZN(n482) );
  INV_X1 U344 ( .A(data_in[4]), .ZN(n481) );
  INV_X1 U345 ( .A(data_in[5]), .ZN(n480) );
  INV_X1 U346 ( .A(data_in[6]), .ZN(n479) );
  INV_X1 U347 ( .A(data_in[7]), .ZN(n478) );
  INV_X1 U356 ( .A(data_in[8]), .ZN(n477) );
  INV_X1 U357 ( .A(data_in[9]), .ZN(n476) );
  INV_X1 U358 ( .A(data_in[10]), .ZN(n475) );
  INV_X1 U359 ( .A(data_in[11]), .ZN(n474) );
  INV_X1 U360 ( .A(data_in[12]), .ZN(n473) );
  INV_X1 U361 ( .A(data_in[13]), .ZN(n472) );
  INV_X1 U362 ( .A(data_in[14]), .ZN(n471) );
  INV_X1 U363 ( .A(data_in[15]), .ZN(n470) );
  INV_X1 U364 ( .A(data_in[16]), .ZN(n469) );
  INV_X1 U365 ( .A(data_in[17]), .ZN(n468) );
  INV_X1 U366 ( .A(data_in[18]), .ZN(n467) );
  INV_X1 U367 ( .A(data_in[19]), .ZN(n466) );
  MUX2_X1 U368 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(N10), .Z(n1) );
  MUX2_X1 U369 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(N10), .Z(n2) );
  MUX2_X1 U370 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U371 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n452), .Z(n4) );
  MUX2_X1 U372 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n453), .Z(n5) );
  MUX2_X1 U373 ( .A(n5), .B(n4), .S(n451), .Z(n6) );
  MUX2_X1 U374 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n452), .Z(n7) );
  MUX2_X1 U375 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n454), .Z(n8) );
  MUX2_X1 U376 ( .A(n8), .B(n7), .S(N11), .Z(n9) );
  MUX2_X1 U377 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n453), .Z(n10) );
  MUX2_X1 U378 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(N10), .Z(n11) );
  MUX2_X1 U379 ( .A(n11), .B(n10), .S(n451), .Z(n12) );
  MUX2_X1 U380 ( .A(n12), .B(n9), .S(N12), .Z(N31) );
  MUX2_X1 U381 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n454), .Z(n13) );
  MUX2_X1 U382 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(N10), .Z(n14) );
  MUX2_X1 U383 ( .A(n14), .B(n13), .S(n451), .Z(n15) );
  MUX2_X1 U384 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n453), .Z(n16) );
  MUX2_X1 U385 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n453), .Z(n17) );
  MUX2_X1 U386 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U387 ( .A(n18), .B(n15), .S(N12), .Z(N30) );
  MUX2_X1 U388 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n454), .Z(n19) );
  MUX2_X1 U389 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n454), .Z(n20) );
  MUX2_X1 U390 ( .A(n20), .B(n19), .S(N11), .Z(n21) );
  MUX2_X1 U391 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n453), .Z(n22) );
  MUX2_X1 U392 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n452), .Z(n23) );
  MUX2_X1 U393 ( .A(n23), .B(n22), .S(N11), .Z(n354) );
  MUX2_X1 U394 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n452), .Z(n355) );
  MUX2_X1 U395 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n452), .Z(n356) );
  MUX2_X1 U396 ( .A(n356), .B(n355), .S(n451), .Z(n357) );
  MUX2_X1 U397 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n454), .Z(n358) );
  MUX2_X1 U398 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n452), .Z(n359) );
  MUX2_X1 U399 ( .A(n359), .B(n358), .S(N11), .Z(n360) );
  MUX2_X1 U400 ( .A(n360), .B(n357), .S(N12), .Z(N28) );
  MUX2_X1 U401 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n452), .Z(n361) );
  MUX2_X1 U402 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n452), .Z(n362) );
  MUX2_X1 U403 ( .A(n362), .B(n361), .S(N11), .Z(n363) );
  MUX2_X1 U404 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n452), .Z(n364) );
  MUX2_X1 U405 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n452), .Z(n365) );
  MUX2_X1 U406 ( .A(n365), .B(n364), .S(N11), .Z(n366) );
  MUX2_X1 U407 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n452), .Z(n367) );
  MUX2_X1 U408 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n452), .Z(n368) );
  MUX2_X1 U409 ( .A(n368), .B(n367), .S(n451), .Z(n369) );
  MUX2_X1 U410 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n452), .Z(n370) );
  MUX2_X1 U411 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n452), .Z(n371) );
  MUX2_X1 U412 ( .A(n371), .B(n370), .S(N11), .Z(n372) );
  MUX2_X1 U413 ( .A(n372), .B(n369), .S(N12), .Z(N26) );
  MUX2_X1 U414 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n452), .Z(n373) );
  MUX2_X1 U415 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n452), .Z(n374) );
  MUX2_X1 U416 ( .A(n374), .B(n373), .S(N11), .Z(n375) );
  MUX2_X1 U417 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n452), .Z(n376) );
  MUX2_X1 U418 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n452), .Z(n377) );
  MUX2_X1 U419 ( .A(n377), .B(n376), .S(N11), .Z(n378) );
  MUX2_X1 U420 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n453), .Z(n379) );
  MUX2_X1 U421 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n453), .Z(n380) );
  MUX2_X1 U422 ( .A(n380), .B(n379), .S(n451), .Z(n381) );
  MUX2_X1 U423 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n453), .Z(n382) );
  MUX2_X1 U424 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n453), .Z(n383) );
  MUX2_X1 U425 ( .A(n383), .B(n382), .S(n451), .Z(n384) );
  MUX2_X1 U426 ( .A(n384), .B(n381), .S(N12), .Z(N24) );
  MUX2_X1 U427 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n453), .Z(n385) );
  MUX2_X1 U428 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n453), .Z(n386) );
  MUX2_X1 U429 ( .A(n386), .B(n385), .S(n451), .Z(n387) );
  MUX2_X1 U430 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n453), .Z(n388) );
  MUX2_X1 U431 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n453), .Z(n389) );
  MUX2_X1 U432 ( .A(n389), .B(n388), .S(n451), .Z(n390) );
  MUX2_X1 U433 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n453), .Z(n391) );
  MUX2_X1 U434 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n453), .Z(n392) );
  MUX2_X1 U435 ( .A(n392), .B(n391), .S(n451), .Z(n393) );
  MUX2_X1 U436 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n453), .Z(n394) );
  MUX2_X1 U437 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n453), .Z(n395) );
  MUX2_X1 U438 ( .A(n395), .B(n394), .S(n451), .Z(n396) );
  MUX2_X1 U439 ( .A(n396), .B(n393), .S(N12), .Z(N22) );
  MUX2_X1 U440 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n454), .Z(n397) );
  MUX2_X1 U441 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n454), .Z(n398) );
  MUX2_X1 U442 ( .A(n398), .B(n397), .S(n451), .Z(n399) );
  MUX2_X1 U443 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n454), .Z(n400) );
  MUX2_X1 U444 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n454), .Z(n401) );
  MUX2_X1 U445 ( .A(n401), .B(n400), .S(n451), .Z(n402) );
  MUX2_X1 U446 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n454), .Z(n403) );
  MUX2_X1 U447 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n454), .Z(n404) );
  MUX2_X1 U448 ( .A(n404), .B(n403), .S(n451), .Z(n405) );
  MUX2_X1 U449 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n454), .Z(n406) );
  MUX2_X1 U450 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n454), .Z(n407) );
  MUX2_X1 U451 ( .A(n407), .B(n406), .S(n451), .Z(n408) );
  MUX2_X1 U452 ( .A(n408), .B(n405), .S(N12), .Z(N20) );
  MUX2_X1 U453 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n454), .Z(n409) );
  MUX2_X1 U454 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n454), .Z(n410) );
  MUX2_X1 U455 ( .A(n410), .B(n409), .S(n451), .Z(n411) );
  MUX2_X1 U456 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n454), .Z(n412) );
  MUX2_X1 U457 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n454), .Z(n413) );
  MUX2_X1 U458 ( .A(n413), .B(n412), .S(n451), .Z(n414) );
  MUX2_X1 U459 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n453), .Z(n415) );
  MUX2_X1 U460 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n453), .Z(n416) );
  MUX2_X1 U461 ( .A(n416), .B(n415), .S(n451), .Z(n417) );
  MUX2_X1 U462 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n453), .Z(n418) );
  MUX2_X1 U463 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(N10), .Z(n419) );
  MUX2_X1 U464 ( .A(n419), .B(n418), .S(N11), .Z(n420) );
  MUX2_X1 U465 ( .A(n420), .B(n417), .S(N12), .Z(N18) );
  MUX2_X1 U466 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(N10), .Z(n421) );
  MUX2_X1 U467 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(N10), .Z(n422) );
  MUX2_X1 U468 ( .A(n422), .B(n421), .S(N11), .Z(n423) );
  MUX2_X1 U469 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(N10), .Z(n424) );
  MUX2_X1 U470 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(N10), .Z(n425) );
  MUX2_X1 U471 ( .A(n425), .B(n424), .S(n451), .Z(n426) );
  MUX2_X1 U472 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n454), .Z(n427) );
  MUX2_X1 U473 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n454), .Z(n428) );
  MUX2_X1 U474 ( .A(n428), .B(n427), .S(n451), .Z(n429) );
  MUX2_X1 U475 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n454), .Z(n430) );
  MUX2_X1 U476 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(N10), .Z(n431) );
  MUX2_X1 U477 ( .A(n431), .B(n430), .S(N11), .Z(n432) );
  MUX2_X1 U478 ( .A(n432), .B(n429), .S(N12), .Z(N16) );
  MUX2_X1 U479 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n452), .Z(n433) );
  MUX2_X1 U480 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n453), .Z(n434) );
  MUX2_X1 U481 ( .A(n434), .B(n433), .S(N11), .Z(n435) );
  MUX2_X1 U482 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(N10), .Z(n436) );
  MUX2_X1 U483 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n452), .Z(n437) );
  MUX2_X1 U484 ( .A(n437), .B(n436), .S(n451), .Z(n438) );
  MUX2_X1 U485 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n453), .Z(n439) );
  MUX2_X1 U486 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n454), .Z(n440) );
  MUX2_X1 U487 ( .A(n440), .B(n439), .S(n451), .Z(n441) );
  MUX2_X1 U488 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n452), .Z(n442) );
  MUX2_X1 U489 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n453), .Z(n443) );
  MUX2_X1 U490 ( .A(n443), .B(n442), .S(N11), .Z(n444) );
  MUX2_X1 U491 ( .A(n444), .B(n441), .S(N12), .Z(N14) );
  MUX2_X1 U492 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n454), .Z(n445) );
  MUX2_X1 U493 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n452), .Z(n446) );
  MUX2_X1 U494 ( .A(n446), .B(n445), .S(n451), .Z(n447) );
  MUX2_X1 U495 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n452), .Z(n448) );
  MUX2_X1 U496 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n454), .Z(n449) );
  MUX2_X1 U497 ( .A(n449), .B(n448), .S(N11), .Z(n450) );
  MUX2_X1 U498 ( .A(n450), .B(n447), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE3_5 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N13, N14, N16, N18, N20, N22, N24, N26, N28, N30, N31,
         N32, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[19]  ( .D(N13), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \data_out_reg[18]  ( .D(N14), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[16]  ( .D(N16), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N20), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N22), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[8]  ( .D(N24), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N26), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N28), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N30), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N32), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n486), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n487), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n488), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n489), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n490), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n491), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n492), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n493), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n494), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n495), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n496), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n497), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n498), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n499), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n500), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n501), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n502), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n503), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n504), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n505), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n506), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n507), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n508), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n509), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n510), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n511), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n512), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n513), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n514), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n515), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n516), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n517), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n518), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n519), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n520), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n521), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n522), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n523), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n524), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n525), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n526), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n527), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n528), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n529), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n530), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n531), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n532), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n533), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n534), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n535), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n536), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n537), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n538), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n539), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n540), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n541), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n542), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n543), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n544), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n545), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n546), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n547), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n548), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n549), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n550), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n551), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n552), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n553), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n554), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n555), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n556), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n557), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n558), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n559), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n560), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n561), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n562), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n563), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n564), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n565), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n566), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n567), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n568), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n569), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n570), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n571), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n572), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n573), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n574), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n575), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n576), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n577), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n578), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n579), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n580), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n581), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n582), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n583), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n584), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n585), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n586), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n587), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n588), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n589), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n590), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n591), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n592), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n593), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n594), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n595), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n596), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n597), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n598), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n599), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n600), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n601), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n602), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n603), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n604), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n605), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n606), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n607), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n608), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n609), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n610), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n611), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n612), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n613), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n614), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n615), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n616), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n617), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n618), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n619), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n620), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n621), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n622), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n623), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n624), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n625), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n626), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n627), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n628), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n629), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n630), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n631), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n632), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n633), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n634), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n635), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n636), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n637), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n638), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n639), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n640), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n641), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n642), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n643), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n644), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n645), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U348 ( .A1(n463), .A2(n464), .A3(n794), .ZN(n815) );
  NAND3_X1 U349 ( .A1(n794), .A2(n464), .A3(N10), .ZN(n793) );
  NAND3_X1 U350 ( .A1(n794), .A2(n463), .A3(N11), .ZN(n772) );
  NAND3_X1 U351 ( .A1(N10), .A2(n794), .A3(N11), .ZN(n751) );
  NAND3_X1 U352 ( .A1(n463), .A2(n464), .A3(n709), .ZN(n730) );
  NAND3_X1 U353 ( .A1(N10), .A2(n464), .A3(n709), .ZN(n708) );
  NAND3_X1 U354 ( .A1(N11), .A2(n463), .A3(n709), .ZN(n687) );
  NAND3_X1 U355 ( .A1(N11), .A2(N10), .A3(n709), .ZN(n666) );
  DFF_X1 \data_out_reg[1]  ( .D(N31), .CK(clk), .Q(data_out[1]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n402), .SI(n399), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n354), .SI(n21), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n414), .SI(n411), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n426), .SI(n423), .SE(N12), .CK(clk), .Q(
        data_out[15]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n366), .SI(n363), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[17]  ( .D(n438), .SI(n435), .SE(N12), .CK(clk), .Q(
        data_out[17]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n378), .SI(n375), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n390), .SI(n387), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  BUF_X1 U3 ( .A(n666), .Z(n455) );
  BUF_X1 U4 ( .A(n772), .Z(n460) );
  BUF_X1 U5 ( .A(n730), .Z(n458) );
  BUF_X1 U6 ( .A(n751), .Z(n459) );
  BUF_X1 U7 ( .A(n793), .Z(n461) );
  BUF_X1 U8 ( .A(n708), .Z(n457) );
  BUF_X1 U9 ( .A(n687), .Z(n456) );
  BUF_X1 U10 ( .A(n815), .Z(n462) );
  BUF_X1 U11 ( .A(N10), .Z(n454) );
  BUF_X1 U12 ( .A(N10), .Z(n453) );
  BUF_X1 U13 ( .A(N11), .Z(n451) );
  NOR2_X1 U14 ( .A1(n465), .A2(N12), .ZN(n794) );
  INV_X1 U15 ( .A(wr_en), .ZN(n465) );
  AND2_X1 U16 ( .A1(N12), .A2(wr_en), .ZN(n709) );
  OAI21_X1 U17 ( .B1(n485), .B2(n793), .A(n792), .ZN(n625) );
  NAND2_X1 U18 ( .A1(\mem[1][0] ), .A2(n461), .ZN(n792) );
  OAI21_X1 U19 ( .B1(n484), .B2(n793), .A(n791), .ZN(n624) );
  NAND2_X1 U20 ( .A1(\mem[1][1] ), .A2(n461), .ZN(n791) );
  OAI21_X1 U21 ( .B1(n483), .B2(n793), .A(n790), .ZN(n623) );
  NAND2_X1 U22 ( .A1(\mem[1][2] ), .A2(n461), .ZN(n790) );
  OAI21_X1 U23 ( .B1(n482), .B2(n793), .A(n789), .ZN(n622) );
  NAND2_X1 U24 ( .A1(\mem[1][3] ), .A2(n461), .ZN(n789) );
  OAI21_X1 U25 ( .B1(n481), .B2(n461), .A(n788), .ZN(n621) );
  NAND2_X1 U26 ( .A1(\mem[1][4] ), .A2(n461), .ZN(n788) );
  OAI21_X1 U27 ( .B1(n480), .B2(n461), .A(n787), .ZN(n620) );
  NAND2_X1 U28 ( .A1(\mem[1][5] ), .A2(n461), .ZN(n787) );
  OAI21_X1 U29 ( .B1(n479), .B2(n793), .A(n786), .ZN(n619) );
  NAND2_X1 U30 ( .A1(\mem[1][6] ), .A2(n461), .ZN(n786) );
  OAI21_X1 U31 ( .B1(n478), .B2(n793), .A(n785), .ZN(n618) );
  NAND2_X1 U32 ( .A1(\mem[1][7] ), .A2(n461), .ZN(n785) );
  OAI21_X1 U33 ( .B1(n477), .B2(n793), .A(n784), .ZN(n617) );
  NAND2_X1 U34 ( .A1(\mem[1][8] ), .A2(n461), .ZN(n784) );
  OAI21_X1 U35 ( .B1(n476), .B2(n793), .A(n783), .ZN(n616) );
  NAND2_X1 U36 ( .A1(\mem[1][9] ), .A2(n461), .ZN(n783) );
  OAI21_X1 U37 ( .B1(n475), .B2(n793), .A(n782), .ZN(n615) );
  NAND2_X1 U38 ( .A1(\mem[1][10] ), .A2(n461), .ZN(n782) );
  OAI21_X1 U39 ( .B1(n474), .B2(n793), .A(n781), .ZN(n614) );
  NAND2_X1 U40 ( .A1(\mem[1][11] ), .A2(n461), .ZN(n781) );
  OAI21_X1 U41 ( .B1(n473), .B2(n793), .A(n780), .ZN(n613) );
  NAND2_X1 U42 ( .A1(\mem[1][12] ), .A2(n793), .ZN(n780) );
  OAI21_X1 U43 ( .B1(n472), .B2(n793), .A(n779), .ZN(n612) );
  NAND2_X1 U44 ( .A1(\mem[1][13] ), .A2(n793), .ZN(n779) );
  OAI21_X1 U45 ( .B1(n471), .B2(n793), .A(n778), .ZN(n611) );
  NAND2_X1 U46 ( .A1(\mem[1][14] ), .A2(n793), .ZN(n778) );
  OAI21_X1 U47 ( .B1(n470), .B2(n793), .A(n777), .ZN(n610) );
  NAND2_X1 U48 ( .A1(\mem[1][15] ), .A2(n461), .ZN(n777) );
  OAI21_X1 U49 ( .B1(n469), .B2(n793), .A(n776), .ZN(n609) );
  NAND2_X1 U50 ( .A1(\mem[1][16] ), .A2(n793), .ZN(n776) );
  OAI21_X1 U51 ( .B1(n468), .B2(n793), .A(n775), .ZN(n608) );
  NAND2_X1 U52 ( .A1(\mem[1][17] ), .A2(n793), .ZN(n775) );
  OAI21_X1 U53 ( .B1(n467), .B2(n793), .A(n774), .ZN(n607) );
  NAND2_X1 U54 ( .A1(\mem[1][18] ), .A2(n793), .ZN(n774) );
  OAI21_X1 U55 ( .B1(n466), .B2(n793), .A(n773), .ZN(n606) );
  NAND2_X1 U56 ( .A1(\mem[1][19] ), .A2(n461), .ZN(n773) );
  OAI21_X1 U57 ( .B1(n485), .B2(n772), .A(n771), .ZN(n605) );
  NAND2_X1 U58 ( .A1(\mem[2][0] ), .A2(n772), .ZN(n771) );
  OAI21_X1 U59 ( .B1(n484), .B2(n772), .A(n770), .ZN(n604) );
  NAND2_X1 U60 ( .A1(\mem[2][1] ), .A2(n772), .ZN(n770) );
  OAI21_X1 U61 ( .B1(n483), .B2(n772), .A(n769), .ZN(n603) );
  NAND2_X1 U62 ( .A1(\mem[2][2] ), .A2(n772), .ZN(n769) );
  OAI21_X1 U63 ( .B1(n482), .B2(n460), .A(n768), .ZN(n602) );
  NAND2_X1 U64 ( .A1(\mem[2][3] ), .A2(n772), .ZN(n768) );
  OAI21_X1 U65 ( .B1(n481), .B2(n460), .A(n767), .ZN(n601) );
  NAND2_X1 U66 ( .A1(\mem[2][4] ), .A2(n772), .ZN(n767) );
  OAI21_X1 U67 ( .B1(n480), .B2(n460), .A(n766), .ZN(n600) );
  NAND2_X1 U68 ( .A1(\mem[2][5] ), .A2(n772), .ZN(n766) );
  OAI21_X1 U69 ( .B1(n479), .B2(n460), .A(n765), .ZN(n599) );
  NAND2_X1 U70 ( .A1(\mem[2][6] ), .A2(n772), .ZN(n765) );
  OAI21_X1 U71 ( .B1(n478), .B2(n460), .A(n764), .ZN(n598) );
  NAND2_X1 U72 ( .A1(\mem[2][7] ), .A2(n772), .ZN(n764) );
  OAI21_X1 U73 ( .B1(n477), .B2(n460), .A(n763), .ZN(n597) );
  NAND2_X1 U74 ( .A1(\mem[2][8] ), .A2(n772), .ZN(n763) );
  OAI21_X1 U75 ( .B1(n476), .B2(n460), .A(n762), .ZN(n596) );
  NAND2_X1 U76 ( .A1(\mem[2][9] ), .A2(n772), .ZN(n762) );
  OAI21_X1 U77 ( .B1(n475), .B2(n460), .A(n761), .ZN(n595) );
  NAND2_X1 U78 ( .A1(\mem[2][10] ), .A2(n772), .ZN(n761) );
  OAI21_X1 U79 ( .B1(n474), .B2(n460), .A(n760), .ZN(n594) );
  NAND2_X1 U80 ( .A1(\mem[2][11] ), .A2(n772), .ZN(n760) );
  OAI21_X1 U81 ( .B1(n473), .B2(n460), .A(n759), .ZN(n593) );
  NAND2_X1 U82 ( .A1(\mem[2][12] ), .A2(n772), .ZN(n759) );
  OAI21_X1 U83 ( .B1(n472), .B2(n460), .A(n758), .ZN(n592) );
  NAND2_X1 U84 ( .A1(\mem[2][13] ), .A2(n772), .ZN(n758) );
  OAI21_X1 U85 ( .B1(n471), .B2(n460), .A(n757), .ZN(n591) );
  NAND2_X1 U86 ( .A1(\mem[2][14] ), .A2(n772), .ZN(n757) );
  OAI21_X1 U87 ( .B1(n470), .B2(n460), .A(n756), .ZN(n590) );
  NAND2_X1 U88 ( .A1(\mem[2][15] ), .A2(n772), .ZN(n756) );
  OAI21_X1 U89 ( .B1(n469), .B2(n460), .A(n755), .ZN(n589) );
  NAND2_X1 U90 ( .A1(\mem[2][16] ), .A2(n772), .ZN(n755) );
  OAI21_X1 U91 ( .B1(n468), .B2(n460), .A(n754), .ZN(n588) );
  NAND2_X1 U92 ( .A1(\mem[2][17] ), .A2(n772), .ZN(n754) );
  OAI21_X1 U93 ( .B1(n467), .B2(n460), .A(n753), .ZN(n587) );
  NAND2_X1 U94 ( .A1(\mem[2][18] ), .A2(n772), .ZN(n753) );
  OAI21_X1 U95 ( .B1(n466), .B2(n772), .A(n752), .ZN(n586) );
  NAND2_X1 U96 ( .A1(\mem[2][19] ), .A2(n772), .ZN(n752) );
  OAI21_X1 U97 ( .B1(n485), .B2(n751), .A(n750), .ZN(n585) );
  NAND2_X1 U98 ( .A1(\mem[3][0] ), .A2(n459), .ZN(n750) );
  OAI21_X1 U99 ( .B1(n484), .B2(n751), .A(n749), .ZN(n584) );
  NAND2_X1 U100 ( .A1(\mem[3][1] ), .A2(n459), .ZN(n749) );
  OAI21_X1 U101 ( .B1(n483), .B2(n751), .A(n748), .ZN(n583) );
  NAND2_X1 U102 ( .A1(\mem[3][2] ), .A2(n459), .ZN(n748) );
  OAI21_X1 U103 ( .B1(n482), .B2(n751), .A(n747), .ZN(n582) );
  NAND2_X1 U104 ( .A1(\mem[3][3] ), .A2(n459), .ZN(n747) );
  OAI21_X1 U105 ( .B1(n481), .B2(n459), .A(n746), .ZN(n581) );
  NAND2_X1 U106 ( .A1(\mem[3][4] ), .A2(n459), .ZN(n746) );
  OAI21_X1 U107 ( .B1(n480), .B2(n459), .A(n745), .ZN(n580) );
  NAND2_X1 U108 ( .A1(\mem[3][5] ), .A2(n459), .ZN(n745) );
  OAI21_X1 U109 ( .B1(n479), .B2(n751), .A(n744), .ZN(n579) );
  NAND2_X1 U110 ( .A1(\mem[3][6] ), .A2(n459), .ZN(n744) );
  OAI21_X1 U111 ( .B1(n478), .B2(n751), .A(n743), .ZN(n578) );
  NAND2_X1 U112 ( .A1(\mem[3][7] ), .A2(n459), .ZN(n743) );
  OAI21_X1 U113 ( .B1(n477), .B2(n751), .A(n742), .ZN(n577) );
  NAND2_X1 U114 ( .A1(\mem[3][8] ), .A2(n459), .ZN(n742) );
  OAI21_X1 U115 ( .B1(n476), .B2(n751), .A(n741), .ZN(n576) );
  NAND2_X1 U116 ( .A1(\mem[3][9] ), .A2(n459), .ZN(n741) );
  OAI21_X1 U117 ( .B1(n475), .B2(n751), .A(n740), .ZN(n575) );
  NAND2_X1 U118 ( .A1(\mem[3][10] ), .A2(n459), .ZN(n740) );
  OAI21_X1 U119 ( .B1(n474), .B2(n751), .A(n739), .ZN(n574) );
  NAND2_X1 U120 ( .A1(\mem[3][11] ), .A2(n459), .ZN(n739) );
  OAI21_X1 U121 ( .B1(n473), .B2(n751), .A(n738), .ZN(n573) );
  NAND2_X1 U122 ( .A1(\mem[3][12] ), .A2(n751), .ZN(n738) );
  OAI21_X1 U123 ( .B1(n472), .B2(n751), .A(n737), .ZN(n572) );
  NAND2_X1 U124 ( .A1(\mem[3][13] ), .A2(n751), .ZN(n737) );
  OAI21_X1 U125 ( .B1(n471), .B2(n751), .A(n736), .ZN(n571) );
  NAND2_X1 U126 ( .A1(\mem[3][14] ), .A2(n751), .ZN(n736) );
  OAI21_X1 U127 ( .B1(n470), .B2(n751), .A(n735), .ZN(n570) );
  NAND2_X1 U128 ( .A1(\mem[3][15] ), .A2(n459), .ZN(n735) );
  OAI21_X1 U129 ( .B1(n469), .B2(n751), .A(n734), .ZN(n569) );
  NAND2_X1 U130 ( .A1(\mem[3][16] ), .A2(n751), .ZN(n734) );
  OAI21_X1 U131 ( .B1(n468), .B2(n751), .A(n733), .ZN(n568) );
  NAND2_X1 U132 ( .A1(\mem[3][17] ), .A2(n751), .ZN(n733) );
  OAI21_X1 U133 ( .B1(n467), .B2(n751), .A(n732), .ZN(n567) );
  NAND2_X1 U134 ( .A1(\mem[3][18] ), .A2(n751), .ZN(n732) );
  OAI21_X1 U135 ( .B1(n466), .B2(n751), .A(n731), .ZN(n566) );
  NAND2_X1 U136 ( .A1(\mem[3][19] ), .A2(n459), .ZN(n731) );
  OAI21_X1 U137 ( .B1(n485), .B2(n730), .A(n729), .ZN(n565) );
  NAND2_X1 U138 ( .A1(\mem[4][0] ), .A2(n730), .ZN(n729) );
  OAI21_X1 U139 ( .B1(n484), .B2(n458), .A(n728), .ZN(n564) );
  NAND2_X1 U140 ( .A1(\mem[4][1] ), .A2(n730), .ZN(n728) );
  OAI21_X1 U141 ( .B1(n483), .B2(n458), .A(n727), .ZN(n563) );
  NAND2_X1 U142 ( .A1(\mem[4][2] ), .A2(n730), .ZN(n727) );
  OAI21_X1 U143 ( .B1(n482), .B2(n458), .A(n726), .ZN(n562) );
  NAND2_X1 U144 ( .A1(\mem[4][3] ), .A2(n730), .ZN(n726) );
  OAI21_X1 U145 ( .B1(n481), .B2(n458), .A(n725), .ZN(n561) );
  NAND2_X1 U146 ( .A1(\mem[4][4] ), .A2(n730), .ZN(n725) );
  OAI21_X1 U147 ( .B1(n480), .B2(n458), .A(n724), .ZN(n560) );
  NAND2_X1 U148 ( .A1(\mem[4][5] ), .A2(n730), .ZN(n724) );
  OAI21_X1 U149 ( .B1(n479), .B2(n458), .A(n723), .ZN(n559) );
  NAND2_X1 U150 ( .A1(\mem[4][6] ), .A2(n730), .ZN(n723) );
  OAI21_X1 U151 ( .B1(n478), .B2(n458), .A(n722), .ZN(n558) );
  NAND2_X1 U152 ( .A1(\mem[4][7] ), .A2(n730), .ZN(n722) );
  OAI21_X1 U153 ( .B1(n477), .B2(n458), .A(n721), .ZN(n557) );
  NAND2_X1 U154 ( .A1(\mem[4][8] ), .A2(n730), .ZN(n721) );
  OAI21_X1 U155 ( .B1(n476), .B2(n730), .A(n720), .ZN(n556) );
  NAND2_X1 U156 ( .A1(\mem[4][9] ), .A2(n730), .ZN(n720) );
  OAI21_X1 U157 ( .B1(n475), .B2(n458), .A(n719), .ZN(n555) );
  NAND2_X1 U158 ( .A1(\mem[4][10] ), .A2(n730), .ZN(n719) );
  OAI21_X1 U159 ( .B1(n474), .B2(n458), .A(n718), .ZN(n554) );
  NAND2_X1 U160 ( .A1(\mem[4][11] ), .A2(n730), .ZN(n718) );
  OAI21_X1 U161 ( .B1(n473), .B2(n730), .A(n717), .ZN(n553) );
  NAND2_X1 U162 ( .A1(\mem[4][12] ), .A2(n730), .ZN(n717) );
  OAI21_X1 U163 ( .B1(n472), .B2(n458), .A(n716), .ZN(n552) );
  NAND2_X1 U164 ( .A1(\mem[4][13] ), .A2(n730), .ZN(n716) );
  OAI21_X1 U165 ( .B1(n471), .B2(n730), .A(n715), .ZN(n551) );
  NAND2_X1 U166 ( .A1(\mem[4][14] ), .A2(n730), .ZN(n715) );
  OAI21_X1 U167 ( .B1(n470), .B2(n458), .A(n714), .ZN(n550) );
  NAND2_X1 U168 ( .A1(\mem[4][15] ), .A2(n730), .ZN(n714) );
  OAI21_X1 U169 ( .B1(n469), .B2(n458), .A(n713), .ZN(n549) );
  NAND2_X1 U170 ( .A1(\mem[4][16] ), .A2(n730), .ZN(n713) );
  OAI21_X1 U171 ( .B1(n468), .B2(n458), .A(n712), .ZN(n548) );
  NAND2_X1 U172 ( .A1(\mem[4][17] ), .A2(n730), .ZN(n712) );
  OAI21_X1 U173 ( .B1(n467), .B2(n458), .A(n711), .ZN(n547) );
  NAND2_X1 U174 ( .A1(\mem[4][18] ), .A2(n730), .ZN(n711) );
  OAI21_X1 U175 ( .B1(n466), .B2(n458), .A(n710), .ZN(n546) );
  NAND2_X1 U176 ( .A1(\mem[4][19] ), .A2(n730), .ZN(n710) );
  OAI21_X1 U177 ( .B1(n485), .B2(n708), .A(n707), .ZN(n545) );
  NAND2_X1 U178 ( .A1(\mem[5][0] ), .A2(n457), .ZN(n707) );
  OAI21_X1 U179 ( .B1(n484), .B2(n708), .A(n706), .ZN(n544) );
  NAND2_X1 U180 ( .A1(\mem[5][1] ), .A2(n457), .ZN(n706) );
  OAI21_X1 U181 ( .B1(n483), .B2(n708), .A(n705), .ZN(n543) );
  NAND2_X1 U182 ( .A1(\mem[5][2] ), .A2(n457), .ZN(n705) );
  OAI21_X1 U183 ( .B1(n482), .B2(n708), .A(n704), .ZN(n542) );
  NAND2_X1 U184 ( .A1(\mem[5][3] ), .A2(n457), .ZN(n704) );
  OAI21_X1 U185 ( .B1(n481), .B2(n457), .A(n703), .ZN(n541) );
  NAND2_X1 U186 ( .A1(\mem[5][4] ), .A2(n457), .ZN(n703) );
  OAI21_X1 U187 ( .B1(n480), .B2(n708), .A(n702), .ZN(n540) );
  NAND2_X1 U188 ( .A1(\mem[5][5] ), .A2(n457), .ZN(n702) );
  OAI21_X1 U189 ( .B1(n479), .B2(n708), .A(n701), .ZN(n539) );
  NAND2_X1 U190 ( .A1(\mem[5][6] ), .A2(n457), .ZN(n701) );
  OAI21_X1 U191 ( .B1(n478), .B2(n708), .A(n700), .ZN(n538) );
  NAND2_X1 U192 ( .A1(\mem[5][7] ), .A2(n457), .ZN(n700) );
  OAI21_X1 U193 ( .B1(n477), .B2(n708), .A(n699), .ZN(n537) );
  NAND2_X1 U194 ( .A1(\mem[5][8] ), .A2(n457), .ZN(n699) );
  OAI21_X1 U195 ( .B1(n476), .B2(n708), .A(n698), .ZN(n536) );
  NAND2_X1 U196 ( .A1(\mem[5][9] ), .A2(n457), .ZN(n698) );
  OAI21_X1 U197 ( .B1(n475), .B2(n708), .A(n697), .ZN(n535) );
  NAND2_X1 U198 ( .A1(\mem[5][10] ), .A2(n457), .ZN(n697) );
  OAI21_X1 U199 ( .B1(n474), .B2(n708), .A(n696), .ZN(n534) );
  NAND2_X1 U200 ( .A1(\mem[5][11] ), .A2(n457), .ZN(n696) );
  OAI21_X1 U201 ( .B1(n473), .B2(n708), .A(n695), .ZN(n533) );
  NAND2_X1 U202 ( .A1(\mem[5][12] ), .A2(n708), .ZN(n695) );
  OAI21_X1 U203 ( .B1(n472), .B2(n457), .A(n694), .ZN(n532) );
  NAND2_X1 U204 ( .A1(\mem[5][13] ), .A2(n708), .ZN(n694) );
  OAI21_X1 U205 ( .B1(n471), .B2(n457), .A(n693), .ZN(n531) );
  NAND2_X1 U206 ( .A1(\mem[5][14] ), .A2(n708), .ZN(n693) );
  OAI21_X1 U207 ( .B1(n470), .B2(n708), .A(n692), .ZN(n530) );
  NAND2_X1 U208 ( .A1(\mem[5][15] ), .A2(n708), .ZN(n692) );
  OAI21_X1 U209 ( .B1(n469), .B2(n708), .A(n691), .ZN(n529) );
  NAND2_X1 U210 ( .A1(\mem[5][16] ), .A2(n708), .ZN(n691) );
  OAI21_X1 U211 ( .B1(n468), .B2(n708), .A(n690), .ZN(n528) );
  NAND2_X1 U212 ( .A1(\mem[5][17] ), .A2(n708), .ZN(n690) );
  OAI21_X1 U213 ( .B1(n467), .B2(n708), .A(n689), .ZN(n527) );
  NAND2_X1 U214 ( .A1(\mem[5][18] ), .A2(n708), .ZN(n689) );
  OAI21_X1 U215 ( .B1(n466), .B2(n708), .A(n688), .ZN(n526) );
  NAND2_X1 U216 ( .A1(\mem[5][19] ), .A2(n457), .ZN(n688) );
  OAI21_X1 U217 ( .B1(n485), .B2(n687), .A(n686), .ZN(n525) );
  NAND2_X1 U218 ( .A1(\mem[6][0] ), .A2(n456), .ZN(n686) );
  OAI21_X1 U219 ( .B1(n484), .B2(n687), .A(n685), .ZN(n524) );
  NAND2_X1 U220 ( .A1(\mem[6][1] ), .A2(n456), .ZN(n685) );
  OAI21_X1 U221 ( .B1(n483), .B2(n687), .A(n684), .ZN(n523) );
  NAND2_X1 U222 ( .A1(\mem[6][2] ), .A2(n456), .ZN(n684) );
  OAI21_X1 U223 ( .B1(n482), .B2(n687), .A(n683), .ZN(n522) );
  NAND2_X1 U224 ( .A1(\mem[6][3] ), .A2(n456), .ZN(n683) );
  OAI21_X1 U225 ( .B1(n481), .B2(n456), .A(n682), .ZN(n521) );
  NAND2_X1 U226 ( .A1(\mem[6][4] ), .A2(n456), .ZN(n682) );
  OAI21_X1 U227 ( .B1(n480), .B2(n687), .A(n681), .ZN(n520) );
  NAND2_X1 U228 ( .A1(\mem[6][5] ), .A2(n456), .ZN(n681) );
  OAI21_X1 U229 ( .B1(n479), .B2(n687), .A(n680), .ZN(n519) );
  NAND2_X1 U230 ( .A1(\mem[6][6] ), .A2(n456), .ZN(n680) );
  OAI21_X1 U231 ( .B1(n478), .B2(n687), .A(n679), .ZN(n518) );
  NAND2_X1 U232 ( .A1(\mem[6][7] ), .A2(n456), .ZN(n679) );
  OAI21_X1 U233 ( .B1(n477), .B2(n687), .A(n678), .ZN(n517) );
  NAND2_X1 U234 ( .A1(\mem[6][8] ), .A2(n456), .ZN(n678) );
  OAI21_X1 U235 ( .B1(n476), .B2(n687), .A(n677), .ZN(n516) );
  NAND2_X1 U236 ( .A1(\mem[6][9] ), .A2(n456), .ZN(n677) );
  OAI21_X1 U237 ( .B1(n475), .B2(n687), .A(n676), .ZN(n515) );
  NAND2_X1 U238 ( .A1(\mem[6][10] ), .A2(n456), .ZN(n676) );
  OAI21_X1 U239 ( .B1(n474), .B2(n687), .A(n675), .ZN(n514) );
  NAND2_X1 U240 ( .A1(\mem[6][11] ), .A2(n456), .ZN(n675) );
  OAI21_X1 U241 ( .B1(n473), .B2(n687), .A(n674), .ZN(n513) );
  NAND2_X1 U242 ( .A1(\mem[6][12] ), .A2(n687), .ZN(n674) );
  OAI21_X1 U243 ( .B1(n472), .B2(n456), .A(n673), .ZN(n512) );
  NAND2_X1 U244 ( .A1(\mem[6][13] ), .A2(n687), .ZN(n673) );
  OAI21_X1 U245 ( .B1(n471), .B2(n456), .A(n672), .ZN(n511) );
  NAND2_X1 U246 ( .A1(\mem[6][14] ), .A2(n687), .ZN(n672) );
  OAI21_X1 U247 ( .B1(n470), .B2(n687), .A(n671), .ZN(n510) );
  NAND2_X1 U248 ( .A1(\mem[6][15] ), .A2(n687), .ZN(n671) );
  OAI21_X1 U249 ( .B1(n469), .B2(n687), .A(n670), .ZN(n509) );
  NAND2_X1 U250 ( .A1(\mem[6][16] ), .A2(n687), .ZN(n670) );
  OAI21_X1 U251 ( .B1(n468), .B2(n687), .A(n669), .ZN(n508) );
  NAND2_X1 U252 ( .A1(\mem[6][17] ), .A2(n687), .ZN(n669) );
  OAI21_X1 U253 ( .B1(n467), .B2(n687), .A(n668), .ZN(n507) );
  NAND2_X1 U254 ( .A1(\mem[6][18] ), .A2(n687), .ZN(n668) );
  OAI21_X1 U255 ( .B1(n466), .B2(n687), .A(n667), .ZN(n506) );
  NAND2_X1 U256 ( .A1(\mem[6][19] ), .A2(n456), .ZN(n667) );
  OAI21_X1 U257 ( .B1(n485), .B2(n455), .A(n665), .ZN(n505) );
  NAND2_X1 U258 ( .A1(\mem[7][0] ), .A2(n455), .ZN(n665) );
  OAI21_X1 U259 ( .B1(n484), .B2(n455), .A(n664), .ZN(n504) );
  NAND2_X1 U260 ( .A1(\mem[7][1] ), .A2(n455), .ZN(n664) );
  OAI21_X1 U261 ( .B1(n483), .B2(n455), .A(n663), .ZN(n503) );
  NAND2_X1 U262 ( .A1(\mem[7][2] ), .A2(n666), .ZN(n663) );
  OAI21_X1 U263 ( .B1(n482), .B2(n666), .A(n662), .ZN(n502) );
  NAND2_X1 U264 ( .A1(\mem[7][3] ), .A2(n455), .ZN(n662) );
  OAI21_X1 U265 ( .B1(n481), .B2(n666), .A(n661), .ZN(n501) );
  NAND2_X1 U266 ( .A1(\mem[7][4] ), .A2(n666), .ZN(n661) );
  OAI21_X1 U267 ( .B1(n480), .B2(n666), .A(n660), .ZN(n500) );
  NAND2_X1 U268 ( .A1(\mem[7][5] ), .A2(n666), .ZN(n660) );
  OAI21_X1 U269 ( .B1(n479), .B2(n666), .A(n659), .ZN(n499) );
  NAND2_X1 U270 ( .A1(\mem[7][6] ), .A2(n666), .ZN(n659) );
  OAI21_X1 U271 ( .B1(n478), .B2(n666), .A(n658), .ZN(n498) );
  NAND2_X1 U272 ( .A1(\mem[7][7] ), .A2(n666), .ZN(n658) );
  OAI21_X1 U273 ( .B1(n477), .B2(n666), .A(n657), .ZN(n497) );
  NAND2_X1 U274 ( .A1(\mem[7][8] ), .A2(n666), .ZN(n657) );
  OAI21_X1 U275 ( .B1(n476), .B2(n455), .A(n656), .ZN(n496) );
  NAND2_X1 U276 ( .A1(\mem[7][9] ), .A2(n666), .ZN(n656) );
  OAI21_X1 U277 ( .B1(n475), .B2(n666), .A(n655), .ZN(n495) );
  NAND2_X1 U278 ( .A1(\mem[7][10] ), .A2(n666), .ZN(n655) );
  OAI21_X1 U279 ( .B1(n474), .B2(n666), .A(n654), .ZN(n494) );
  NAND2_X1 U280 ( .A1(\mem[7][11] ), .A2(n666), .ZN(n654) );
  OAI21_X1 U281 ( .B1(n473), .B2(n455), .A(n653), .ZN(n493) );
  NAND2_X1 U282 ( .A1(\mem[7][12] ), .A2(n455), .ZN(n653) );
  OAI21_X1 U283 ( .B1(n472), .B2(n455), .A(n652), .ZN(n492) );
  NAND2_X1 U284 ( .A1(\mem[7][13] ), .A2(n455), .ZN(n652) );
  OAI21_X1 U285 ( .B1(n471), .B2(n455), .A(n651), .ZN(n491) );
  NAND2_X1 U286 ( .A1(\mem[7][14] ), .A2(n455), .ZN(n651) );
  OAI21_X1 U287 ( .B1(n470), .B2(n666), .A(n650), .ZN(n490) );
  NAND2_X1 U288 ( .A1(\mem[7][15] ), .A2(n455), .ZN(n650) );
  OAI21_X1 U289 ( .B1(n469), .B2(n666), .A(n649), .ZN(n489) );
  NAND2_X1 U290 ( .A1(\mem[7][16] ), .A2(n455), .ZN(n649) );
  OAI21_X1 U291 ( .B1(n468), .B2(n666), .A(n648), .ZN(n488) );
  NAND2_X1 U292 ( .A1(\mem[7][17] ), .A2(n455), .ZN(n648) );
  OAI21_X1 U293 ( .B1(n467), .B2(n455), .A(n647), .ZN(n487) );
  NAND2_X1 U294 ( .A1(\mem[7][18] ), .A2(n455), .ZN(n647) );
  OAI21_X1 U295 ( .B1(n466), .B2(n455), .A(n646), .ZN(n486) );
  NAND2_X1 U296 ( .A1(\mem[7][19] ), .A2(n455), .ZN(n646) );
  OAI21_X1 U297 ( .B1(n815), .B2(n483), .A(n812), .ZN(n643) );
  NAND2_X1 U298 ( .A1(\mem[0][2] ), .A2(n815), .ZN(n812) );
  OAI21_X1 U299 ( .B1(n815), .B2(n482), .A(n811), .ZN(n642) );
  NAND2_X1 U300 ( .A1(\mem[0][3] ), .A2(n815), .ZN(n811) );
  OAI21_X1 U301 ( .B1(n815), .B2(n481), .A(n810), .ZN(n641) );
  NAND2_X1 U302 ( .A1(\mem[0][4] ), .A2(n815), .ZN(n810) );
  OAI21_X1 U303 ( .B1(n815), .B2(n480), .A(n809), .ZN(n640) );
  NAND2_X1 U304 ( .A1(\mem[0][5] ), .A2(n815), .ZN(n809) );
  OAI21_X1 U305 ( .B1(n815), .B2(n479), .A(n808), .ZN(n639) );
  NAND2_X1 U306 ( .A1(\mem[0][6] ), .A2(n815), .ZN(n808) );
  OAI21_X1 U307 ( .B1(n462), .B2(n478), .A(n807), .ZN(n638) );
  NAND2_X1 U308 ( .A1(\mem[0][7] ), .A2(n815), .ZN(n807) );
  OAI21_X1 U309 ( .B1(n462), .B2(n477), .A(n806), .ZN(n637) );
  NAND2_X1 U310 ( .A1(\mem[0][8] ), .A2(n815), .ZN(n806) );
  OAI21_X1 U311 ( .B1(n462), .B2(n476), .A(n805), .ZN(n636) );
  NAND2_X1 U312 ( .A1(\mem[0][9] ), .A2(n462), .ZN(n805) );
  OAI21_X1 U313 ( .B1(n462), .B2(n475), .A(n804), .ZN(n635) );
  NAND2_X1 U314 ( .A1(\mem[0][10] ), .A2(n815), .ZN(n804) );
  OAI21_X1 U315 ( .B1(n462), .B2(n474), .A(n803), .ZN(n634) );
  NAND2_X1 U316 ( .A1(\mem[0][11] ), .A2(n815), .ZN(n803) );
  OAI21_X1 U317 ( .B1(n815), .B2(n473), .A(n802), .ZN(n633) );
  NAND2_X1 U318 ( .A1(\mem[0][12] ), .A2(n462), .ZN(n802) );
  OAI21_X1 U319 ( .B1(n815), .B2(n472), .A(n801), .ZN(n632) );
  NAND2_X1 U320 ( .A1(\mem[0][13] ), .A2(n462), .ZN(n801) );
  OAI21_X1 U321 ( .B1(n462), .B2(n471), .A(n800), .ZN(n631) );
  NAND2_X1 U322 ( .A1(\mem[0][14] ), .A2(n462), .ZN(n800) );
  OAI21_X1 U323 ( .B1(n462), .B2(n470), .A(n799), .ZN(n630) );
  NAND2_X1 U324 ( .A1(\mem[0][15] ), .A2(n462), .ZN(n799) );
  OAI21_X1 U325 ( .B1(n815), .B2(n469), .A(n798), .ZN(n629) );
  NAND2_X1 U326 ( .A1(\mem[0][16] ), .A2(n462), .ZN(n798) );
  OAI21_X1 U327 ( .B1(n815), .B2(n468), .A(n797), .ZN(n628) );
  NAND2_X1 U328 ( .A1(\mem[0][17] ), .A2(n462), .ZN(n797) );
  OAI21_X1 U329 ( .B1(n815), .B2(n467), .A(n796), .ZN(n627) );
  NAND2_X1 U330 ( .A1(\mem[0][18] ), .A2(n462), .ZN(n796) );
  OAI21_X1 U331 ( .B1(n815), .B2(n485), .A(n814), .ZN(n645) );
  NAND2_X1 U332 ( .A1(\mem[0][0] ), .A2(n815), .ZN(n814) );
  OAI21_X1 U333 ( .B1(n815), .B2(n484), .A(n813), .ZN(n644) );
  NAND2_X1 U334 ( .A1(\mem[0][1] ), .A2(n815), .ZN(n813) );
  OAI21_X1 U335 ( .B1(n815), .B2(n466), .A(n795), .ZN(n626) );
  NAND2_X1 U336 ( .A1(\mem[0][19] ), .A2(n462), .ZN(n795) );
  INV_X1 U337 ( .A(N10), .ZN(n463) );
  INV_X1 U338 ( .A(N11), .ZN(n464) );
  INV_X1 U339 ( .A(data_in[0]), .ZN(n485) );
  INV_X1 U340 ( .A(data_in[1]), .ZN(n484) );
  INV_X1 U341 ( .A(data_in[2]), .ZN(n483) );
  INV_X1 U342 ( .A(data_in[3]), .ZN(n482) );
  INV_X1 U343 ( .A(data_in[4]), .ZN(n481) );
  INV_X1 U344 ( .A(data_in[5]), .ZN(n480) );
  INV_X1 U345 ( .A(data_in[6]), .ZN(n479) );
  INV_X1 U346 ( .A(data_in[7]), .ZN(n478) );
  INV_X1 U347 ( .A(data_in[8]), .ZN(n477) );
  INV_X1 U356 ( .A(data_in[9]), .ZN(n476) );
  INV_X1 U357 ( .A(data_in[10]), .ZN(n475) );
  INV_X1 U358 ( .A(data_in[11]), .ZN(n474) );
  INV_X1 U359 ( .A(data_in[12]), .ZN(n473) );
  INV_X1 U360 ( .A(data_in[13]), .ZN(n472) );
  INV_X1 U361 ( .A(data_in[14]), .ZN(n471) );
  INV_X1 U362 ( .A(data_in[15]), .ZN(n470) );
  INV_X1 U363 ( .A(data_in[16]), .ZN(n469) );
  INV_X1 U364 ( .A(data_in[17]), .ZN(n468) );
  INV_X1 U365 ( .A(data_in[18]), .ZN(n467) );
  INV_X1 U366 ( .A(data_in[19]), .ZN(n466) );
  MUX2_X1 U367 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n452), .Z(n1) );
  MUX2_X1 U368 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n452), .Z(n2) );
  MUX2_X1 U369 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U370 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n452), .Z(n4) );
  MUX2_X1 U371 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n452), .Z(n5) );
  MUX2_X1 U372 ( .A(n5), .B(n4), .S(N11), .Z(n6) );
  MUX2_X1 U373 ( .A(n6), .B(n3), .S(N12), .Z(N32) );
  MUX2_X1 U374 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n452), .Z(n7) );
  MUX2_X1 U375 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n452), .Z(n8) );
  MUX2_X1 U376 ( .A(n8), .B(n7), .S(N11), .Z(n9) );
  MUX2_X1 U377 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n452), .Z(n10) );
  MUX2_X1 U378 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n452), .Z(n11) );
  MUX2_X1 U379 ( .A(n11), .B(n10), .S(N11), .Z(n12) );
  MUX2_X1 U380 ( .A(n12), .B(n9), .S(N12), .Z(N31) );
  MUX2_X1 U381 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n453), .Z(n13) );
  MUX2_X1 U382 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n453), .Z(n14) );
  MUX2_X1 U383 ( .A(n14), .B(n13), .S(N11), .Z(n15) );
  MUX2_X1 U384 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n453), .Z(n16) );
  MUX2_X1 U385 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n453), .Z(n17) );
  MUX2_X1 U386 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U387 ( .A(n18), .B(n15), .S(N12), .Z(N30) );
  MUX2_X1 U388 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n453), .Z(n19) );
  MUX2_X1 U389 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n453), .Z(n20) );
  MUX2_X1 U390 ( .A(n20), .B(n19), .S(N11), .Z(n21) );
  MUX2_X1 U391 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n453), .Z(n22) );
  MUX2_X1 U392 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n453), .Z(n23) );
  MUX2_X1 U393 ( .A(n23), .B(n22), .S(N11), .Z(n354) );
  MUX2_X1 U394 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n453), .Z(n355) );
  MUX2_X1 U395 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n453), .Z(n356) );
  MUX2_X1 U396 ( .A(n356), .B(n355), .S(n451), .Z(n357) );
  MUX2_X1 U397 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n453), .Z(n358) );
  MUX2_X1 U398 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n453), .Z(n359) );
  MUX2_X1 U399 ( .A(n359), .B(n358), .S(N11), .Z(n360) );
  MUX2_X1 U400 ( .A(n360), .B(n357), .S(N12), .Z(N28) );
  MUX2_X1 U401 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n452), .Z(n361) );
  MUX2_X1 U402 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(N10), .Z(n362) );
  MUX2_X1 U403 ( .A(n362), .B(n361), .S(N11), .Z(n363) );
  MUX2_X1 U404 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n364) );
  MUX2_X1 U405 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(N10), .Z(n365) );
  MUX2_X1 U406 ( .A(n365), .B(n364), .S(N11), .Z(n366) );
  MUX2_X1 U407 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n454), .Z(n367) );
  MUX2_X1 U408 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n453), .Z(n368) );
  MUX2_X1 U409 ( .A(n368), .B(n367), .S(N11), .Z(n369) );
  MUX2_X1 U410 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n454), .Z(n370) );
  MUX2_X1 U411 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n452), .Z(n371) );
  MUX2_X1 U412 ( .A(n371), .B(n370), .S(N11), .Z(n372) );
  MUX2_X1 U413 ( .A(n372), .B(n369), .S(N12), .Z(N26) );
  MUX2_X1 U414 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n373) );
  MUX2_X1 U415 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n374) );
  MUX2_X1 U416 ( .A(n374), .B(n373), .S(N11), .Z(n375) );
  MUX2_X1 U417 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n376) );
  MUX2_X1 U418 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n377) );
  MUX2_X1 U419 ( .A(n377), .B(n376), .S(N11), .Z(n378) );
  MUX2_X1 U420 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n453), .Z(n379) );
  MUX2_X1 U421 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n454), .Z(n380) );
  MUX2_X1 U422 ( .A(n380), .B(n379), .S(n451), .Z(n381) );
  MUX2_X1 U423 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n453), .Z(n382) );
  MUX2_X1 U424 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n453), .Z(n383) );
  MUX2_X1 U425 ( .A(n383), .B(n382), .S(n451), .Z(n384) );
  MUX2_X1 U426 ( .A(n384), .B(n381), .S(N12), .Z(N24) );
  MUX2_X1 U427 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n453), .Z(n385) );
  MUX2_X1 U428 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(N10), .Z(n386) );
  MUX2_X1 U429 ( .A(n386), .B(n385), .S(n451), .Z(n387) );
  MUX2_X1 U430 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n454), .Z(n388) );
  MUX2_X1 U431 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n453), .Z(n389) );
  MUX2_X1 U432 ( .A(n389), .B(n388), .S(n451), .Z(n390) );
  MUX2_X1 U433 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n454), .Z(n391) );
  MUX2_X1 U434 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n452), .Z(n392) );
  MUX2_X1 U435 ( .A(n392), .B(n391), .S(n451), .Z(n393) );
  MUX2_X1 U436 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n452), .Z(n394) );
  MUX2_X1 U437 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n452), .Z(n395) );
  MUX2_X1 U438 ( .A(n395), .B(n394), .S(n451), .Z(n396) );
  MUX2_X1 U439 ( .A(n396), .B(n393), .S(N12), .Z(N22) );
  MUX2_X1 U440 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(N10), .Z(n397) );
  MUX2_X1 U441 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n453), .Z(n398) );
  MUX2_X1 U442 ( .A(n398), .B(n397), .S(n451), .Z(n399) );
  MUX2_X1 U443 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n452), .Z(n400) );
  MUX2_X1 U444 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n452), .Z(n401) );
  MUX2_X1 U445 ( .A(n401), .B(n400), .S(n451), .Z(n402) );
  MUX2_X1 U446 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n452), .Z(n403) );
  MUX2_X1 U447 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n453), .Z(n404) );
  MUX2_X1 U448 ( .A(n404), .B(n403), .S(n451), .Z(n405) );
  MUX2_X1 U449 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n452), .Z(n406) );
  MUX2_X1 U450 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n454), .Z(n407) );
  MUX2_X1 U451 ( .A(n407), .B(n406), .S(n451), .Z(n408) );
  MUX2_X1 U452 ( .A(n408), .B(n405), .S(N12), .Z(N20) );
  MUX2_X1 U453 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n452), .Z(n409) );
  MUX2_X1 U454 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n454), .Z(n410) );
  MUX2_X1 U455 ( .A(n410), .B(n409), .S(n451), .Z(n411) );
  MUX2_X1 U456 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(N10), .Z(n412) );
  MUX2_X1 U457 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n453), .Z(n413) );
  MUX2_X1 U458 ( .A(n413), .B(n412), .S(n451), .Z(n414) );
  MUX2_X1 U459 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n452), .Z(n415) );
  MUX2_X1 U460 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n454), .Z(n416) );
  MUX2_X1 U461 ( .A(n416), .B(n415), .S(n451), .Z(n417) );
  MUX2_X1 U462 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n452), .Z(n418) );
  MUX2_X1 U463 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n454), .Z(n419) );
  MUX2_X1 U464 ( .A(n419), .B(n418), .S(n451), .Z(n420) );
  MUX2_X1 U465 ( .A(n420), .B(n417), .S(N12), .Z(N18) );
  MUX2_X1 U466 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n452), .Z(n421) );
  MUX2_X1 U467 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n453), .Z(n422) );
  MUX2_X1 U468 ( .A(n422), .B(n421), .S(n451), .Z(n423) );
  MUX2_X1 U469 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n454), .Z(n424) );
  MUX2_X1 U470 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(N10), .Z(n425) );
  MUX2_X1 U471 ( .A(n425), .B(n424), .S(n451), .Z(n426) );
  MUX2_X1 U472 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n452), .Z(n427) );
  MUX2_X1 U473 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n453), .Z(n428) );
  MUX2_X1 U474 ( .A(n428), .B(n427), .S(N11), .Z(n429) );
  MUX2_X1 U475 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n454), .Z(n430) );
  MUX2_X1 U476 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n452), .Z(n431) );
  MUX2_X1 U477 ( .A(n431), .B(n430), .S(n451), .Z(n432) );
  MUX2_X1 U478 ( .A(n432), .B(n429), .S(N12), .Z(N16) );
  MUX2_X1 U479 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n454), .Z(n433) );
  MUX2_X1 U480 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n454), .Z(n434) );
  MUX2_X1 U481 ( .A(n434), .B(n433), .S(n451), .Z(n435) );
  MUX2_X1 U482 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n454), .Z(n436) );
  MUX2_X1 U483 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n454), .Z(n437) );
  MUX2_X1 U484 ( .A(n437), .B(n436), .S(n451), .Z(n438) );
  MUX2_X1 U485 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n454), .Z(n439) );
  MUX2_X1 U486 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n454), .Z(n440) );
  MUX2_X1 U487 ( .A(n440), .B(n439), .S(N11), .Z(n441) );
  MUX2_X1 U488 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n454), .Z(n442) );
  MUX2_X1 U489 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n454), .Z(n443) );
  MUX2_X1 U490 ( .A(n443), .B(n442), .S(n451), .Z(n444) );
  MUX2_X1 U491 ( .A(n444), .B(n441), .S(N12), .Z(N14) );
  MUX2_X1 U492 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n454), .Z(n445) );
  MUX2_X1 U493 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n454), .Z(n446) );
  MUX2_X1 U494 ( .A(n446), .B(n445), .S(n451), .Z(n447) );
  MUX2_X1 U495 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n454), .Z(n448) );
  MUX2_X1 U496 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n454), .Z(n449) );
  MUX2_X1 U497 ( .A(n449), .B(n448), .S(n451), .Z(n450) );
  MUX2_X1 U498 ( .A(n450), .B(n447), .S(N12), .Z(N13) );
  CLKBUF_X1 U499 ( .A(N10), .Z(n452) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE3_4 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N14, N18, N20, N26, N28, N30, N32, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[18]  ( .D(N14), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N20), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[6]  ( .D(N26), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N28), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N30), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N32), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n486), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n487), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n488), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n489), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n490), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n491), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n492), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n493), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n494), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n495), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n496), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n497), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n498), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n499), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n500), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n501), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n502), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n503), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n504), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n505), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n506), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n507), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n508), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n509), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n510), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n511), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n512), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n513), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n514), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n515), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n516), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n517), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n518), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n519), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n520), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n521), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n522), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n523), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n524), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n525), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n526), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n527), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n528), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n529), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n530), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n531), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n532), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n533), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n534), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n535), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n536), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n537), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n538), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n539), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n540), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n541), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n542), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n543), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n544), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n545), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n546), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n547), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n548), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n549), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n550), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n551), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n552), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n553), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n554), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n555), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n556), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n557), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n558), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n559), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n560), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n561), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n562), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n563), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n564), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n565), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n566), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n567), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n568), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n569), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n570), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n571), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n572), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n573), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n574), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n575), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n576), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n577), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n578), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n579), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n580), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n581), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n582), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n583), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n584), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n585), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n586), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n587), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n588), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n589), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n590), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n591), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n592), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n593), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n594), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n595), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n596), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n597), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n598), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n599), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n600), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n601), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n602), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n603), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n604), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n605), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n606), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n607), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n608), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n609), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n610), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n611), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n612), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n613), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n614), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n615), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n616), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n617), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n618), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n619), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n620), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n621), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n622), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n623), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n624), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n625), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n626), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n627), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n628), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n629), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n630), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n631), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n632), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n633), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n634), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n635), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n636), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n637), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n638), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n639), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n640), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n641), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n642), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n643), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n644), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n645), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U348 ( .A1(n463), .A2(n464), .A3(n794), .ZN(n815) );
  NAND3_X1 U349 ( .A1(n794), .A2(n464), .A3(N10), .ZN(n793) );
  NAND3_X1 U350 ( .A1(n794), .A2(n463), .A3(N11), .ZN(n772) );
  NAND3_X1 U351 ( .A1(N10), .A2(n794), .A3(N11), .ZN(n751) );
  NAND3_X1 U352 ( .A1(n463), .A2(n464), .A3(n709), .ZN(n730) );
  NAND3_X1 U353 ( .A1(N10), .A2(n464), .A3(n709), .ZN(n708) );
  NAND3_X1 U354 ( .A1(N11), .A2(n463), .A3(n709), .ZN(n687) );
  NAND3_X1 U355 ( .A1(N11), .A2(N10), .A3(n709), .ZN(n666) );
  SDFF_X1 \data_out_reg[1]  ( .D(n12), .SI(n9), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n354), .SI(n21), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n426), .SI(n423), .SE(N12), .CK(clk), .Q(
        data_out[15]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n378), .SI(n375), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n414), .SI(n411), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n366), .SI(n363), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[17]  ( .D(n438), .SI(n435), .SE(N12), .CK(clk), .Q(
        data_out[17]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n402), .SI(n399), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[19]  ( .D(n450), .SI(n447), .SE(N12), .CK(clk), .Q(
        data_out[19]) );
  SDFF_X1 \data_out_reg[16]  ( .D(n432), .SI(n429), .SE(N12), .CK(clk), .Q(
        data_out[16]) );
  SDFF_X1 \data_out_reg[10]  ( .D(n396), .SI(n393), .SE(N12), .CK(clk), .Q(
        data_out[10]) );
  SDFF_X1 \data_out_reg[8]  ( .D(n384), .SI(n381), .SE(N12), .CK(clk), .Q(
        data_out[8]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n390), .SI(n387), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  BUF_X1 U3 ( .A(n666), .Z(n455) );
  BUF_X1 U4 ( .A(n708), .Z(n457) );
  BUF_X1 U5 ( .A(n730), .Z(n458) );
  BUF_X1 U6 ( .A(n815), .Z(n462) );
  BUF_X1 U7 ( .A(n751), .Z(n459) );
  BUF_X1 U8 ( .A(n793), .Z(n461) );
  BUF_X1 U9 ( .A(n687), .Z(n456) );
  BUF_X1 U10 ( .A(n772), .Z(n460) );
  BUF_X1 U11 ( .A(N10), .Z(n452) );
  BUF_X1 U12 ( .A(N10), .Z(n453) );
  BUF_X1 U13 ( .A(N10), .Z(n454) );
  BUF_X1 U14 ( .A(N11), .Z(n451) );
  NOR2_X1 U15 ( .A1(n465), .A2(N12), .ZN(n794) );
  INV_X1 U16 ( .A(wr_en), .ZN(n465) );
  AND2_X1 U17 ( .A1(N12), .A2(wr_en), .ZN(n709) );
  OAI21_X1 U18 ( .B1(n485), .B2(n793), .A(n792), .ZN(n625) );
  NAND2_X1 U19 ( .A1(\mem[1][0] ), .A2(n461), .ZN(n792) );
  OAI21_X1 U20 ( .B1(n484), .B2(n793), .A(n791), .ZN(n624) );
  NAND2_X1 U21 ( .A1(\mem[1][1] ), .A2(n461), .ZN(n791) );
  OAI21_X1 U22 ( .B1(n483), .B2(n793), .A(n790), .ZN(n623) );
  NAND2_X1 U23 ( .A1(\mem[1][2] ), .A2(n461), .ZN(n790) );
  OAI21_X1 U24 ( .B1(n482), .B2(n793), .A(n789), .ZN(n622) );
  NAND2_X1 U25 ( .A1(\mem[1][3] ), .A2(n461), .ZN(n789) );
  OAI21_X1 U26 ( .B1(n481), .B2(n461), .A(n788), .ZN(n621) );
  NAND2_X1 U27 ( .A1(\mem[1][4] ), .A2(n461), .ZN(n788) );
  OAI21_X1 U28 ( .B1(n480), .B2(n461), .A(n787), .ZN(n620) );
  NAND2_X1 U29 ( .A1(\mem[1][5] ), .A2(n461), .ZN(n787) );
  OAI21_X1 U30 ( .B1(n479), .B2(n793), .A(n786), .ZN(n619) );
  NAND2_X1 U31 ( .A1(\mem[1][6] ), .A2(n461), .ZN(n786) );
  OAI21_X1 U32 ( .B1(n478), .B2(n793), .A(n785), .ZN(n618) );
  NAND2_X1 U33 ( .A1(\mem[1][7] ), .A2(n461), .ZN(n785) );
  OAI21_X1 U34 ( .B1(n477), .B2(n793), .A(n784), .ZN(n617) );
  NAND2_X1 U35 ( .A1(\mem[1][8] ), .A2(n461), .ZN(n784) );
  OAI21_X1 U36 ( .B1(n476), .B2(n793), .A(n783), .ZN(n616) );
  NAND2_X1 U37 ( .A1(\mem[1][9] ), .A2(n461), .ZN(n783) );
  OAI21_X1 U38 ( .B1(n475), .B2(n793), .A(n782), .ZN(n615) );
  NAND2_X1 U39 ( .A1(\mem[1][10] ), .A2(n461), .ZN(n782) );
  OAI21_X1 U40 ( .B1(n474), .B2(n793), .A(n781), .ZN(n614) );
  NAND2_X1 U41 ( .A1(\mem[1][11] ), .A2(n461), .ZN(n781) );
  OAI21_X1 U42 ( .B1(n473), .B2(n793), .A(n780), .ZN(n613) );
  NAND2_X1 U43 ( .A1(\mem[1][12] ), .A2(n793), .ZN(n780) );
  OAI21_X1 U44 ( .B1(n472), .B2(n793), .A(n779), .ZN(n612) );
  NAND2_X1 U45 ( .A1(\mem[1][13] ), .A2(n793), .ZN(n779) );
  OAI21_X1 U46 ( .B1(n471), .B2(n793), .A(n778), .ZN(n611) );
  NAND2_X1 U47 ( .A1(\mem[1][14] ), .A2(n793), .ZN(n778) );
  OAI21_X1 U48 ( .B1(n470), .B2(n793), .A(n777), .ZN(n610) );
  NAND2_X1 U49 ( .A1(\mem[1][15] ), .A2(n461), .ZN(n777) );
  OAI21_X1 U50 ( .B1(n469), .B2(n793), .A(n776), .ZN(n609) );
  NAND2_X1 U51 ( .A1(\mem[1][16] ), .A2(n793), .ZN(n776) );
  OAI21_X1 U52 ( .B1(n468), .B2(n793), .A(n775), .ZN(n608) );
  NAND2_X1 U53 ( .A1(\mem[1][17] ), .A2(n793), .ZN(n775) );
  OAI21_X1 U54 ( .B1(n467), .B2(n793), .A(n774), .ZN(n607) );
  NAND2_X1 U55 ( .A1(\mem[1][18] ), .A2(n793), .ZN(n774) );
  OAI21_X1 U56 ( .B1(n466), .B2(n793), .A(n773), .ZN(n606) );
  NAND2_X1 U57 ( .A1(\mem[1][19] ), .A2(n461), .ZN(n773) );
  OAI21_X1 U58 ( .B1(n485), .B2(n772), .A(n771), .ZN(n605) );
  NAND2_X1 U59 ( .A1(\mem[2][0] ), .A2(n772), .ZN(n771) );
  OAI21_X1 U60 ( .B1(n484), .B2(n772), .A(n770), .ZN(n604) );
  NAND2_X1 U61 ( .A1(\mem[2][1] ), .A2(n772), .ZN(n770) );
  OAI21_X1 U62 ( .B1(n483), .B2(n772), .A(n769), .ZN(n603) );
  NAND2_X1 U63 ( .A1(\mem[2][2] ), .A2(n772), .ZN(n769) );
  OAI21_X1 U64 ( .B1(n482), .B2(n460), .A(n768), .ZN(n602) );
  NAND2_X1 U65 ( .A1(\mem[2][3] ), .A2(n460), .ZN(n768) );
  OAI21_X1 U66 ( .B1(n481), .B2(n772), .A(n767), .ZN(n601) );
  NAND2_X1 U67 ( .A1(\mem[2][4] ), .A2(n460), .ZN(n767) );
  OAI21_X1 U68 ( .B1(n480), .B2(n772), .A(n766), .ZN(n600) );
  NAND2_X1 U69 ( .A1(\mem[2][5] ), .A2(n460), .ZN(n766) );
  OAI21_X1 U70 ( .B1(n479), .B2(n772), .A(n765), .ZN(n599) );
  NAND2_X1 U71 ( .A1(\mem[2][6] ), .A2(n772), .ZN(n765) );
  OAI21_X1 U72 ( .B1(n478), .B2(n772), .A(n764), .ZN(n598) );
  NAND2_X1 U73 ( .A1(\mem[2][7] ), .A2(n772), .ZN(n764) );
  OAI21_X1 U74 ( .B1(n477), .B2(n460), .A(n763), .ZN(n597) );
  NAND2_X1 U75 ( .A1(\mem[2][8] ), .A2(n772), .ZN(n763) );
  OAI21_X1 U76 ( .B1(n476), .B2(n772), .A(n762), .ZN(n596) );
  NAND2_X1 U77 ( .A1(\mem[2][9] ), .A2(n772), .ZN(n762) );
  OAI21_X1 U78 ( .B1(n475), .B2(n460), .A(n761), .ZN(n595) );
  NAND2_X1 U79 ( .A1(\mem[2][10] ), .A2(n772), .ZN(n761) );
  OAI21_X1 U80 ( .B1(n474), .B2(n460), .A(n760), .ZN(n594) );
  NAND2_X1 U81 ( .A1(\mem[2][11] ), .A2(n772), .ZN(n760) );
  OAI21_X1 U82 ( .B1(n473), .B2(n460), .A(n759), .ZN(n593) );
  NAND2_X1 U83 ( .A1(\mem[2][12] ), .A2(n460), .ZN(n759) );
  OAI21_X1 U84 ( .B1(n472), .B2(n772), .A(n758), .ZN(n592) );
  NAND2_X1 U85 ( .A1(\mem[2][13] ), .A2(n460), .ZN(n758) );
  OAI21_X1 U86 ( .B1(n471), .B2(n772), .A(n757), .ZN(n591) );
  NAND2_X1 U87 ( .A1(\mem[2][14] ), .A2(n460), .ZN(n757) );
  OAI21_X1 U88 ( .B1(n470), .B2(n772), .A(n756), .ZN(n590) );
  NAND2_X1 U89 ( .A1(\mem[2][15] ), .A2(n460), .ZN(n756) );
  OAI21_X1 U90 ( .B1(n469), .B2(n772), .A(n755), .ZN(n589) );
  NAND2_X1 U91 ( .A1(\mem[2][16] ), .A2(n460), .ZN(n755) );
  OAI21_X1 U92 ( .B1(n468), .B2(n772), .A(n754), .ZN(n588) );
  NAND2_X1 U93 ( .A1(\mem[2][17] ), .A2(n460), .ZN(n754) );
  OAI21_X1 U94 ( .B1(n467), .B2(n772), .A(n753), .ZN(n587) );
  NAND2_X1 U95 ( .A1(\mem[2][18] ), .A2(n460), .ZN(n753) );
  OAI21_X1 U96 ( .B1(n466), .B2(n772), .A(n752), .ZN(n586) );
  NAND2_X1 U97 ( .A1(\mem[2][19] ), .A2(n460), .ZN(n752) );
  OAI21_X1 U98 ( .B1(n485), .B2(n751), .A(n750), .ZN(n585) );
  NAND2_X1 U99 ( .A1(\mem[3][0] ), .A2(n459), .ZN(n750) );
  OAI21_X1 U100 ( .B1(n484), .B2(n751), .A(n749), .ZN(n584) );
  NAND2_X1 U101 ( .A1(\mem[3][1] ), .A2(n459), .ZN(n749) );
  OAI21_X1 U102 ( .B1(n483), .B2(n751), .A(n748), .ZN(n583) );
  NAND2_X1 U103 ( .A1(\mem[3][2] ), .A2(n459), .ZN(n748) );
  OAI21_X1 U104 ( .B1(n482), .B2(n751), .A(n747), .ZN(n582) );
  NAND2_X1 U105 ( .A1(\mem[3][3] ), .A2(n459), .ZN(n747) );
  OAI21_X1 U106 ( .B1(n481), .B2(n459), .A(n746), .ZN(n581) );
  NAND2_X1 U107 ( .A1(\mem[3][4] ), .A2(n459), .ZN(n746) );
  OAI21_X1 U108 ( .B1(n480), .B2(n459), .A(n745), .ZN(n580) );
  NAND2_X1 U109 ( .A1(\mem[3][5] ), .A2(n459), .ZN(n745) );
  OAI21_X1 U110 ( .B1(n479), .B2(n751), .A(n744), .ZN(n579) );
  NAND2_X1 U111 ( .A1(\mem[3][6] ), .A2(n459), .ZN(n744) );
  OAI21_X1 U112 ( .B1(n478), .B2(n751), .A(n743), .ZN(n578) );
  NAND2_X1 U113 ( .A1(\mem[3][7] ), .A2(n459), .ZN(n743) );
  OAI21_X1 U114 ( .B1(n477), .B2(n751), .A(n742), .ZN(n577) );
  NAND2_X1 U115 ( .A1(\mem[3][8] ), .A2(n459), .ZN(n742) );
  OAI21_X1 U116 ( .B1(n476), .B2(n751), .A(n741), .ZN(n576) );
  NAND2_X1 U117 ( .A1(\mem[3][9] ), .A2(n459), .ZN(n741) );
  OAI21_X1 U118 ( .B1(n475), .B2(n751), .A(n740), .ZN(n575) );
  NAND2_X1 U119 ( .A1(\mem[3][10] ), .A2(n459), .ZN(n740) );
  OAI21_X1 U120 ( .B1(n474), .B2(n751), .A(n739), .ZN(n574) );
  NAND2_X1 U121 ( .A1(\mem[3][11] ), .A2(n459), .ZN(n739) );
  OAI21_X1 U122 ( .B1(n473), .B2(n751), .A(n738), .ZN(n573) );
  NAND2_X1 U123 ( .A1(\mem[3][12] ), .A2(n751), .ZN(n738) );
  OAI21_X1 U124 ( .B1(n472), .B2(n751), .A(n737), .ZN(n572) );
  NAND2_X1 U125 ( .A1(\mem[3][13] ), .A2(n751), .ZN(n737) );
  OAI21_X1 U126 ( .B1(n471), .B2(n751), .A(n736), .ZN(n571) );
  NAND2_X1 U127 ( .A1(\mem[3][14] ), .A2(n751), .ZN(n736) );
  OAI21_X1 U128 ( .B1(n470), .B2(n751), .A(n735), .ZN(n570) );
  NAND2_X1 U129 ( .A1(\mem[3][15] ), .A2(n459), .ZN(n735) );
  OAI21_X1 U130 ( .B1(n469), .B2(n751), .A(n734), .ZN(n569) );
  NAND2_X1 U131 ( .A1(\mem[3][16] ), .A2(n751), .ZN(n734) );
  OAI21_X1 U132 ( .B1(n468), .B2(n751), .A(n733), .ZN(n568) );
  NAND2_X1 U133 ( .A1(\mem[3][17] ), .A2(n751), .ZN(n733) );
  OAI21_X1 U134 ( .B1(n467), .B2(n751), .A(n732), .ZN(n567) );
  NAND2_X1 U135 ( .A1(\mem[3][18] ), .A2(n751), .ZN(n732) );
  OAI21_X1 U136 ( .B1(n466), .B2(n751), .A(n731), .ZN(n566) );
  NAND2_X1 U137 ( .A1(\mem[3][19] ), .A2(n459), .ZN(n731) );
  OAI21_X1 U138 ( .B1(n485), .B2(n730), .A(n729), .ZN(n565) );
  NAND2_X1 U139 ( .A1(\mem[4][0] ), .A2(n730), .ZN(n729) );
  OAI21_X1 U140 ( .B1(n484), .B2(n458), .A(n728), .ZN(n564) );
  NAND2_X1 U141 ( .A1(\mem[4][1] ), .A2(n730), .ZN(n728) );
  OAI21_X1 U142 ( .B1(n483), .B2(n458), .A(n727), .ZN(n563) );
  NAND2_X1 U143 ( .A1(\mem[4][2] ), .A2(n730), .ZN(n727) );
  OAI21_X1 U144 ( .B1(n482), .B2(n458), .A(n726), .ZN(n562) );
  NAND2_X1 U145 ( .A1(\mem[4][3] ), .A2(n730), .ZN(n726) );
  OAI21_X1 U146 ( .B1(n481), .B2(n458), .A(n725), .ZN(n561) );
  NAND2_X1 U147 ( .A1(\mem[4][4] ), .A2(n730), .ZN(n725) );
  OAI21_X1 U148 ( .B1(n480), .B2(n458), .A(n724), .ZN(n560) );
  NAND2_X1 U149 ( .A1(\mem[4][5] ), .A2(n730), .ZN(n724) );
  OAI21_X1 U150 ( .B1(n479), .B2(n458), .A(n723), .ZN(n559) );
  NAND2_X1 U151 ( .A1(\mem[4][6] ), .A2(n730), .ZN(n723) );
  OAI21_X1 U152 ( .B1(n478), .B2(n458), .A(n722), .ZN(n558) );
  NAND2_X1 U153 ( .A1(\mem[4][7] ), .A2(n730), .ZN(n722) );
  OAI21_X1 U154 ( .B1(n477), .B2(n458), .A(n721), .ZN(n557) );
  NAND2_X1 U155 ( .A1(\mem[4][8] ), .A2(n730), .ZN(n721) );
  OAI21_X1 U156 ( .B1(n476), .B2(n730), .A(n720), .ZN(n556) );
  NAND2_X1 U157 ( .A1(\mem[4][9] ), .A2(n730), .ZN(n720) );
  OAI21_X1 U158 ( .B1(n475), .B2(n458), .A(n719), .ZN(n555) );
  NAND2_X1 U159 ( .A1(\mem[4][10] ), .A2(n730), .ZN(n719) );
  OAI21_X1 U160 ( .B1(n474), .B2(n458), .A(n718), .ZN(n554) );
  NAND2_X1 U161 ( .A1(\mem[4][11] ), .A2(n730), .ZN(n718) );
  OAI21_X1 U162 ( .B1(n473), .B2(n730), .A(n717), .ZN(n553) );
  NAND2_X1 U163 ( .A1(\mem[4][12] ), .A2(n730), .ZN(n717) );
  OAI21_X1 U164 ( .B1(n472), .B2(n458), .A(n716), .ZN(n552) );
  NAND2_X1 U165 ( .A1(\mem[4][13] ), .A2(n730), .ZN(n716) );
  OAI21_X1 U166 ( .B1(n471), .B2(n730), .A(n715), .ZN(n551) );
  NAND2_X1 U167 ( .A1(\mem[4][14] ), .A2(n730), .ZN(n715) );
  OAI21_X1 U168 ( .B1(n470), .B2(n458), .A(n714), .ZN(n550) );
  NAND2_X1 U169 ( .A1(\mem[4][15] ), .A2(n730), .ZN(n714) );
  OAI21_X1 U170 ( .B1(n469), .B2(n458), .A(n713), .ZN(n549) );
  NAND2_X1 U171 ( .A1(\mem[4][16] ), .A2(n730), .ZN(n713) );
  OAI21_X1 U172 ( .B1(n468), .B2(n458), .A(n712), .ZN(n548) );
  NAND2_X1 U173 ( .A1(\mem[4][17] ), .A2(n730), .ZN(n712) );
  OAI21_X1 U174 ( .B1(n467), .B2(n458), .A(n711), .ZN(n547) );
  NAND2_X1 U175 ( .A1(\mem[4][18] ), .A2(n730), .ZN(n711) );
  OAI21_X1 U176 ( .B1(n466), .B2(n458), .A(n710), .ZN(n546) );
  NAND2_X1 U177 ( .A1(\mem[4][19] ), .A2(n730), .ZN(n710) );
  OAI21_X1 U178 ( .B1(n485), .B2(n457), .A(n707), .ZN(n545) );
  NAND2_X1 U179 ( .A1(\mem[5][0] ), .A2(n457), .ZN(n707) );
  OAI21_X1 U180 ( .B1(n484), .B2(n457), .A(n706), .ZN(n544) );
  NAND2_X1 U181 ( .A1(\mem[5][1] ), .A2(n457), .ZN(n706) );
  OAI21_X1 U182 ( .B1(n483), .B2(n457), .A(n705), .ZN(n543) );
  NAND2_X1 U183 ( .A1(\mem[5][2] ), .A2(n708), .ZN(n705) );
  OAI21_X1 U184 ( .B1(n482), .B2(n708), .A(n704), .ZN(n542) );
  NAND2_X1 U185 ( .A1(\mem[5][3] ), .A2(n457), .ZN(n704) );
  OAI21_X1 U186 ( .B1(n481), .B2(n708), .A(n703), .ZN(n541) );
  NAND2_X1 U187 ( .A1(\mem[5][4] ), .A2(n708), .ZN(n703) );
  OAI21_X1 U188 ( .B1(n480), .B2(n708), .A(n702), .ZN(n540) );
  NAND2_X1 U189 ( .A1(\mem[5][5] ), .A2(n708), .ZN(n702) );
  OAI21_X1 U190 ( .B1(n479), .B2(n708), .A(n701), .ZN(n539) );
  NAND2_X1 U191 ( .A1(\mem[5][6] ), .A2(n708), .ZN(n701) );
  OAI21_X1 U192 ( .B1(n478), .B2(n708), .A(n700), .ZN(n538) );
  NAND2_X1 U193 ( .A1(\mem[5][7] ), .A2(n708), .ZN(n700) );
  OAI21_X1 U194 ( .B1(n477), .B2(n708), .A(n699), .ZN(n537) );
  NAND2_X1 U195 ( .A1(\mem[5][8] ), .A2(n708), .ZN(n699) );
  OAI21_X1 U196 ( .B1(n476), .B2(n457), .A(n698), .ZN(n536) );
  NAND2_X1 U197 ( .A1(\mem[5][9] ), .A2(n708), .ZN(n698) );
  OAI21_X1 U198 ( .B1(n475), .B2(n708), .A(n697), .ZN(n535) );
  NAND2_X1 U199 ( .A1(\mem[5][10] ), .A2(n708), .ZN(n697) );
  OAI21_X1 U200 ( .B1(n474), .B2(n708), .A(n696), .ZN(n534) );
  NAND2_X1 U201 ( .A1(\mem[5][11] ), .A2(n708), .ZN(n696) );
  OAI21_X1 U202 ( .B1(n473), .B2(n457), .A(n695), .ZN(n533) );
  NAND2_X1 U203 ( .A1(\mem[5][12] ), .A2(n457), .ZN(n695) );
  OAI21_X1 U204 ( .B1(n472), .B2(n457), .A(n694), .ZN(n532) );
  NAND2_X1 U205 ( .A1(\mem[5][13] ), .A2(n457), .ZN(n694) );
  OAI21_X1 U206 ( .B1(n471), .B2(n457), .A(n693), .ZN(n531) );
  NAND2_X1 U207 ( .A1(\mem[5][14] ), .A2(n457), .ZN(n693) );
  OAI21_X1 U208 ( .B1(n470), .B2(n708), .A(n692), .ZN(n530) );
  NAND2_X1 U209 ( .A1(\mem[5][15] ), .A2(n457), .ZN(n692) );
  OAI21_X1 U210 ( .B1(n469), .B2(n708), .A(n691), .ZN(n529) );
  NAND2_X1 U211 ( .A1(\mem[5][16] ), .A2(n457), .ZN(n691) );
  OAI21_X1 U212 ( .B1(n468), .B2(n708), .A(n690), .ZN(n528) );
  NAND2_X1 U213 ( .A1(\mem[5][17] ), .A2(n457), .ZN(n690) );
  OAI21_X1 U214 ( .B1(n467), .B2(n708), .A(n689), .ZN(n527) );
  NAND2_X1 U215 ( .A1(\mem[5][18] ), .A2(n457), .ZN(n689) );
  OAI21_X1 U216 ( .B1(n466), .B2(n457), .A(n688), .ZN(n526) );
  NAND2_X1 U217 ( .A1(\mem[5][19] ), .A2(n457), .ZN(n688) );
  OAI21_X1 U218 ( .B1(n485), .B2(n456), .A(n686), .ZN(n525) );
  NAND2_X1 U219 ( .A1(\mem[6][0] ), .A2(n687), .ZN(n686) );
  OAI21_X1 U220 ( .B1(n484), .B2(n456), .A(n685), .ZN(n524) );
  NAND2_X1 U221 ( .A1(\mem[6][1] ), .A2(n687), .ZN(n685) );
  OAI21_X1 U222 ( .B1(n483), .B2(n456), .A(n684), .ZN(n523) );
  NAND2_X1 U223 ( .A1(\mem[6][2] ), .A2(n687), .ZN(n684) );
  OAI21_X1 U224 ( .B1(n482), .B2(n687), .A(n683), .ZN(n522) );
  NAND2_X1 U225 ( .A1(\mem[6][3] ), .A2(n456), .ZN(n683) );
  OAI21_X1 U226 ( .B1(n481), .B2(n687), .A(n682), .ZN(n521) );
  NAND2_X1 U227 ( .A1(\mem[6][4] ), .A2(n456), .ZN(n682) );
  OAI21_X1 U228 ( .B1(n480), .B2(n687), .A(n681), .ZN(n520) );
  NAND2_X1 U229 ( .A1(\mem[6][5] ), .A2(n687), .ZN(n681) );
  OAI21_X1 U230 ( .B1(n479), .B2(n687), .A(n680), .ZN(n519) );
  NAND2_X1 U231 ( .A1(\mem[6][6] ), .A2(n687), .ZN(n680) );
  OAI21_X1 U232 ( .B1(n478), .B2(n687), .A(n679), .ZN(n518) );
  NAND2_X1 U233 ( .A1(\mem[6][7] ), .A2(n687), .ZN(n679) );
  OAI21_X1 U234 ( .B1(n477), .B2(n687), .A(n678), .ZN(n517) );
  NAND2_X1 U235 ( .A1(\mem[6][8] ), .A2(n687), .ZN(n678) );
  OAI21_X1 U236 ( .B1(n476), .B2(n456), .A(n677), .ZN(n516) );
  NAND2_X1 U237 ( .A1(\mem[6][9] ), .A2(n687), .ZN(n677) );
  OAI21_X1 U238 ( .B1(n475), .B2(n687), .A(n676), .ZN(n515) );
  NAND2_X1 U239 ( .A1(\mem[6][10] ), .A2(n687), .ZN(n676) );
  OAI21_X1 U240 ( .B1(n474), .B2(n687), .A(n675), .ZN(n514) );
  NAND2_X1 U241 ( .A1(\mem[6][11] ), .A2(n687), .ZN(n675) );
  OAI21_X1 U242 ( .B1(n473), .B2(n687), .A(n674), .ZN(n513) );
  NAND2_X1 U243 ( .A1(\mem[6][12] ), .A2(n456), .ZN(n674) );
  OAI21_X1 U244 ( .B1(n472), .B2(n456), .A(n673), .ZN(n512) );
  NAND2_X1 U245 ( .A1(\mem[6][13] ), .A2(n456), .ZN(n673) );
  OAI21_X1 U246 ( .B1(n471), .B2(n687), .A(n672), .ZN(n511) );
  NAND2_X1 U247 ( .A1(\mem[6][14] ), .A2(n456), .ZN(n672) );
  OAI21_X1 U248 ( .B1(n470), .B2(n687), .A(n671), .ZN(n510) );
  NAND2_X1 U249 ( .A1(\mem[6][15] ), .A2(n456), .ZN(n671) );
  OAI21_X1 U250 ( .B1(n469), .B2(n687), .A(n670), .ZN(n509) );
  NAND2_X1 U251 ( .A1(\mem[6][16] ), .A2(n456), .ZN(n670) );
  OAI21_X1 U252 ( .B1(n468), .B2(n687), .A(n669), .ZN(n508) );
  NAND2_X1 U253 ( .A1(\mem[6][17] ), .A2(n456), .ZN(n669) );
  OAI21_X1 U254 ( .B1(n467), .B2(n687), .A(n668), .ZN(n507) );
  NAND2_X1 U255 ( .A1(\mem[6][18] ), .A2(n456), .ZN(n668) );
  OAI21_X1 U256 ( .B1(n466), .B2(n456), .A(n667), .ZN(n506) );
  NAND2_X1 U257 ( .A1(\mem[6][19] ), .A2(n456), .ZN(n667) );
  OAI21_X1 U258 ( .B1(n485), .B2(n666), .A(n665), .ZN(n505) );
  NAND2_X1 U259 ( .A1(\mem[7][0] ), .A2(n455), .ZN(n665) );
  OAI21_X1 U260 ( .B1(n484), .B2(n455), .A(n664), .ZN(n504) );
  NAND2_X1 U261 ( .A1(\mem[7][1] ), .A2(n455), .ZN(n664) );
  OAI21_X1 U262 ( .B1(n483), .B2(n666), .A(n663), .ZN(n503) );
  NAND2_X1 U263 ( .A1(\mem[7][2] ), .A2(n455), .ZN(n663) );
  OAI21_X1 U264 ( .B1(n482), .B2(n666), .A(n662), .ZN(n502) );
  NAND2_X1 U265 ( .A1(\mem[7][3] ), .A2(n455), .ZN(n662) );
  OAI21_X1 U266 ( .B1(n481), .B2(n455), .A(n661), .ZN(n501) );
  NAND2_X1 U267 ( .A1(\mem[7][4] ), .A2(n455), .ZN(n661) );
  OAI21_X1 U268 ( .B1(n480), .B2(n666), .A(n660), .ZN(n500) );
  NAND2_X1 U269 ( .A1(\mem[7][5] ), .A2(n455), .ZN(n660) );
  OAI21_X1 U270 ( .B1(n479), .B2(n666), .A(n659), .ZN(n499) );
  NAND2_X1 U271 ( .A1(\mem[7][6] ), .A2(n455), .ZN(n659) );
  OAI21_X1 U272 ( .B1(n478), .B2(n666), .A(n658), .ZN(n498) );
  NAND2_X1 U273 ( .A1(\mem[7][7] ), .A2(n455), .ZN(n658) );
  OAI21_X1 U274 ( .B1(n477), .B2(n666), .A(n657), .ZN(n497) );
  NAND2_X1 U275 ( .A1(\mem[7][8] ), .A2(n455), .ZN(n657) );
  OAI21_X1 U276 ( .B1(n476), .B2(n666), .A(n656), .ZN(n496) );
  NAND2_X1 U277 ( .A1(\mem[7][9] ), .A2(n455), .ZN(n656) );
  OAI21_X1 U278 ( .B1(n475), .B2(n666), .A(n655), .ZN(n495) );
  NAND2_X1 U279 ( .A1(\mem[7][10] ), .A2(n455), .ZN(n655) );
  OAI21_X1 U280 ( .B1(n474), .B2(n666), .A(n654), .ZN(n494) );
  NAND2_X1 U281 ( .A1(\mem[7][11] ), .A2(n455), .ZN(n654) );
  OAI21_X1 U282 ( .B1(n473), .B2(n666), .A(n653), .ZN(n493) );
  NAND2_X1 U283 ( .A1(\mem[7][12] ), .A2(n666), .ZN(n653) );
  OAI21_X1 U284 ( .B1(n472), .B2(n666), .A(n652), .ZN(n492) );
  NAND2_X1 U285 ( .A1(\mem[7][13] ), .A2(n666), .ZN(n652) );
  OAI21_X1 U286 ( .B1(n471), .B2(n666), .A(n651), .ZN(n491) );
  NAND2_X1 U287 ( .A1(\mem[7][14] ), .A2(n666), .ZN(n651) );
  OAI21_X1 U288 ( .B1(n470), .B2(n666), .A(n650), .ZN(n490) );
  NAND2_X1 U289 ( .A1(\mem[7][15] ), .A2(n666), .ZN(n650) );
  OAI21_X1 U290 ( .B1(n469), .B2(n666), .A(n649), .ZN(n489) );
  NAND2_X1 U291 ( .A1(\mem[7][16] ), .A2(n666), .ZN(n649) );
  OAI21_X1 U292 ( .B1(n468), .B2(n666), .A(n648), .ZN(n488) );
  NAND2_X1 U293 ( .A1(\mem[7][17] ), .A2(n666), .ZN(n648) );
  OAI21_X1 U294 ( .B1(n467), .B2(n666), .A(n647), .ZN(n487) );
  NAND2_X1 U295 ( .A1(\mem[7][18] ), .A2(n666), .ZN(n647) );
  OAI21_X1 U296 ( .B1(n466), .B2(n455), .A(n646), .ZN(n486) );
  NAND2_X1 U297 ( .A1(\mem[7][19] ), .A2(n455), .ZN(n646) );
  OAI21_X1 U298 ( .B1(n815), .B2(n483), .A(n812), .ZN(n643) );
  NAND2_X1 U299 ( .A1(\mem[0][2] ), .A2(n462), .ZN(n812) );
  OAI21_X1 U300 ( .B1(n815), .B2(n482), .A(n811), .ZN(n642) );
  NAND2_X1 U301 ( .A1(\mem[0][3] ), .A2(n462), .ZN(n811) );
  OAI21_X1 U302 ( .B1(n815), .B2(n481), .A(n810), .ZN(n641) );
  NAND2_X1 U303 ( .A1(\mem[0][4] ), .A2(n462), .ZN(n810) );
  OAI21_X1 U304 ( .B1(n815), .B2(n480), .A(n809), .ZN(n640) );
  NAND2_X1 U305 ( .A1(\mem[0][5] ), .A2(n462), .ZN(n809) );
  OAI21_X1 U306 ( .B1(n815), .B2(n479), .A(n808), .ZN(n639) );
  NAND2_X1 U307 ( .A1(\mem[0][6] ), .A2(n462), .ZN(n808) );
  OAI21_X1 U308 ( .B1(n815), .B2(n478), .A(n807), .ZN(n638) );
  NAND2_X1 U309 ( .A1(\mem[0][7] ), .A2(n462), .ZN(n807) );
  OAI21_X1 U310 ( .B1(n815), .B2(n477), .A(n806), .ZN(n637) );
  NAND2_X1 U311 ( .A1(\mem[0][8] ), .A2(n462), .ZN(n806) );
  OAI21_X1 U312 ( .B1(n815), .B2(n476), .A(n805), .ZN(n636) );
  NAND2_X1 U313 ( .A1(\mem[0][9] ), .A2(n462), .ZN(n805) );
  OAI21_X1 U314 ( .B1(n815), .B2(n475), .A(n804), .ZN(n635) );
  NAND2_X1 U315 ( .A1(\mem[0][10] ), .A2(n462), .ZN(n804) );
  OAI21_X1 U316 ( .B1(n815), .B2(n474), .A(n803), .ZN(n634) );
  NAND2_X1 U317 ( .A1(\mem[0][11] ), .A2(n462), .ZN(n803) );
  OAI21_X1 U318 ( .B1(n815), .B2(n473), .A(n802), .ZN(n633) );
  NAND2_X1 U319 ( .A1(\mem[0][12] ), .A2(n815), .ZN(n802) );
  OAI21_X1 U320 ( .B1(n815), .B2(n472), .A(n801), .ZN(n632) );
  NAND2_X1 U321 ( .A1(\mem[0][13] ), .A2(n815), .ZN(n801) );
  OAI21_X1 U322 ( .B1(n462), .B2(n471), .A(n800), .ZN(n631) );
  NAND2_X1 U323 ( .A1(\mem[0][14] ), .A2(n815), .ZN(n800) );
  OAI21_X1 U324 ( .B1(n815), .B2(n470), .A(n799), .ZN(n630) );
  NAND2_X1 U325 ( .A1(\mem[0][15] ), .A2(n462), .ZN(n799) );
  OAI21_X1 U326 ( .B1(n815), .B2(n469), .A(n798), .ZN(n629) );
  NAND2_X1 U327 ( .A1(\mem[0][16] ), .A2(n815), .ZN(n798) );
  OAI21_X1 U328 ( .B1(n815), .B2(n468), .A(n797), .ZN(n628) );
  NAND2_X1 U329 ( .A1(\mem[0][17] ), .A2(n815), .ZN(n797) );
  OAI21_X1 U330 ( .B1(n815), .B2(n467), .A(n796), .ZN(n627) );
  NAND2_X1 U331 ( .A1(\mem[0][18] ), .A2(n815), .ZN(n796) );
  OAI21_X1 U332 ( .B1(n462), .B2(n485), .A(n814), .ZN(n645) );
  NAND2_X1 U333 ( .A1(\mem[0][0] ), .A2(n462), .ZN(n814) );
  OAI21_X1 U334 ( .B1(n815), .B2(n484), .A(n813), .ZN(n644) );
  NAND2_X1 U335 ( .A1(\mem[0][1] ), .A2(n462), .ZN(n813) );
  OAI21_X1 U336 ( .B1(n815), .B2(n466), .A(n795), .ZN(n626) );
  NAND2_X1 U337 ( .A1(\mem[0][19] ), .A2(n462), .ZN(n795) );
  INV_X1 U338 ( .A(N10), .ZN(n463) );
  INV_X1 U339 ( .A(N11), .ZN(n464) );
  INV_X1 U340 ( .A(data_in[0]), .ZN(n485) );
  INV_X1 U341 ( .A(data_in[1]), .ZN(n484) );
  INV_X1 U342 ( .A(data_in[2]), .ZN(n483) );
  INV_X1 U343 ( .A(data_in[3]), .ZN(n482) );
  INV_X1 U344 ( .A(data_in[4]), .ZN(n481) );
  INV_X1 U345 ( .A(data_in[5]), .ZN(n480) );
  INV_X1 U346 ( .A(data_in[6]), .ZN(n479) );
  INV_X1 U347 ( .A(data_in[7]), .ZN(n478) );
  INV_X1 U356 ( .A(data_in[8]), .ZN(n477) );
  INV_X1 U357 ( .A(data_in[9]), .ZN(n476) );
  INV_X1 U358 ( .A(data_in[10]), .ZN(n475) );
  INV_X1 U359 ( .A(data_in[11]), .ZN(n474) );
  INV_X1 U360 ( .A(data_in[12]), .ZN(n473) );
  INV_X1 U361 ( .A(data_in[13]), .ZN(n472) );
  INV_X1 U362 ( .A(data_in[14]), .ZN(n471) );
  INV_X1 U363 ( .A(data_in[15]), .ZN(n470) );
  INV_X1 U364 ( .A(data_in[16]), .ZN(n469) );
  INV_X1 U365 ( .A(data_in[17]), .ZN(n468) );
  INV_X1 U366 ( .A(data_in[18]), .ZN(n467) );
  INV_X1 U367 ( .A(data_in[19]), .ZN(n466) );
  MUX2_X1 U368 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n453), .Z(n1) );
  MUX2_X1 U369 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n452), .Z(n2) );
  MUX2_X1 U370 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U371 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n454), .Z(n4) );
  MUX2_X1 U372 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n454), .Z(n5) );
  MUX2_X1 U373 ( .A(n5), .B(n4), .S(N11), .Z(n6) );
  MUX2_X1 U374 ( .A(n6), .B(n3), .S(N12), .Z(N32) );
  MUX2_X1 U375 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n454), .Z(n7) );
  MUX2_X1 U376 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n453), .Z(n8) );
  MUX2_X1 U377 ( .A(n8), .B(n7), .S(N11), .Z(n9) );
  MUX2_X1 U378 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n454), .Z(n10) );
  MUX2_X1 U379 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n453), .Z(n11) );
  MUX2_X1 U380 ( .A(n11), .B(n10), .S(N11), .Z(n12) );
  MUX2_X1 U381 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n452), .Z(n13) );
  MUX2_X1 U382 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n453), .Z(n14) );
  MUX2_X1 U383 ( .A(n14), .B(n13), .S(N11), .Z(n15) );
  MUX2_X1 U384 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n452), .Z(n16) );
  MUX2_X1 U385 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n453), .Z(n17) );
  MUX2_X1 U386 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U387 ( .A(n18), .B(n15), .S(N12), .Z(N30) );
  MUX2_X1 U388 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(N10), .Z(n19) );
  MUX2_X1 U389 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n20) );
  MUX2_X1 U390 ( .A(n20), .B(n19), .S(N11), .Z(n21) );
  MUX2_X1 U391 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n22) );
  MUX2_X1 U392 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n23) );
  MUX2_X1 U393 ( .A(n23), .B(n22), .S(N11), .Z(n354) );
  MUX2_X1 U394 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n453), .Z(n355) );
  MUX2_X1 U395 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n452), .Z(n356) );
  MUX2_X1 U396 ( .A(n356), .B(n355), .S(n451), .Z(n357) );
  MUX2_X1 U397 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n454), .Z(n358) );
  MUX2_X1 U398 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n359) );
  MUX2_X1 U399 ( .A(n359), .B(n358), .S(N11), .Z(n360) );
  MUX2_X1 U400 ( .A(n360), .B(n357), .S(N12), .Z(N28) );
  MUX2_X1 U401 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n452), .Z(n361) );
  MUX2_X1 U402 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(N10), .Z(n362) );
  MUX2_X1 U403 ( .A(n362), .B(n361), .S(N11), .Z(n363) );
  MUX2_X1 U404 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n364) );
  MUX2_X1 U405 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(N10), .Z(n365) );
  MUX2_X1 U406 ( .A(n365), .B(n364), .S(N11), .Z(n366) );
  MUX2_X1 U407 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n453), .Z(n367) );
  MUX2_X1 U408 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n454), .Z(n368) );
  MUX2_X1 U409 ( .A(n368), .B(n367), .S(N11), .Z(n369) );
  MUX2_X1 U410 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n454), .Z(n370) );
  MUX2_X1 U411 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n454), .Z(n371) );
  MUX2_X1 U412 ( .A(n371), .B(n370), .S(N11), .Z(n372) );
  MUX2_X1 U413 ( .A(n372), .B(n369), .S(N12), .Z(N26) );
  MUX2_X1 U414 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n453), .Z(n373) );
  MUX2_X1 U415 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n452), .Z(n374) );
  MUX2_X1 U416 ( .A(n374), .B(n373), .S(N11), .Z(n375) );
  MUX2_X1 U417 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n454), .Z(n376) );
  MUX2_X1 U418 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n452), .Z(n377) );
  MUX2_X1 U419 ( .A(n377), .B(n376), .S(N11), .Z(n378) );
  MUX2_X1 U420 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(N10), .Z(n379) );
  MUX2_X1 U421 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n454), .Z(n380) );
  MUX2_X1 U422 ( .A(n380), .B(n379), .S(n451), .Z(n381) );
  MUX2_X1 U423 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n453), .Z(n382) );
  MUX2_X1 U424 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n454), .Z(n383) );
  MUX2_X1 U425 ( .A(n383), .B(n382), .S(n451), .Z(n384) );
  MUX2_X1 U426 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n453), .Z(n385) );
  MUX2_X1 U427 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(N10), .Z(n386) );
  MUX2_X1 U428 ( .A(n386), .B(n385), .S(n451), .Z(n387) );
  MUX2_X1 U429 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n453), .Z(n388) );
  MUX2_X1 U430 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(N10), .Z(n389) );
  MUX2_X1 U431 ( .A(n389), .B(n388), .S(n451), .Z(n390) );
  MUX2_X1 U432 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n452), .Z(n391) );
  MUX2_X1 U433 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n452), .Z(n392) );
  MUX2_X1 U434 ( .A(n392), .B(n391), .S(n451), .Z(n393) );
  MUX2_X1 U435 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n452), .Z(n394) );
  MUX2_X1 U436 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n452), .Z(n395) );
  MUX2_X1 U437 ( .A(n395), .B(n394), .S(n451), .Z(n396) );
  MUX2_X1 U438 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n452), .Z(n397) );
  MUX2_X1 U439 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n452), .Z(n398) );
  MUX2_X1 U440 ( .A(n398), .B(n397), .S(n451), .Z(n399) );
  MUX2_X1 U441 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n452), .Z(n400) );
  MUX2_X1 U442 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n452), .Z(n401) );
  MUX2_X1 U443 ( .A(n401), .B(n400), .S(n451), .Z(n402) );
  MUX2_X1 U444 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n452), .Z(n403) );
  MUX2_X1 U445 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n452), .Z(n404) );
  MUX2_X1 U446 ( .A(n404), .B(n403), .S(n451), .Z(n405) );
  MUX2_X1 U447 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n452), .Z(n406) );
  MUX2_X1 U448 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n452), .Z(n407) );
  MUX2_X1 U449 ( .A(n407), .B(n406), .S(n451), .Z(n408) );
  MUX2_X1 U450 ( .A(n408), .B(n405), .S(N12), .Z(N20) );
  MUX2_X1 U451 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n452), .Z(n409) );
  MUX2_X1 U452 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n452), .Z(n410) );
  MUX2_X1 U453 ( .A(n410), .B(n409), .S(n451), .Z(n411) );
  MUX2_X1 U454 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n452), .Z(n412) );
  MUX2_X1 U455 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n452), .Z(n413) );
  MUX2_X1 U456 ( .A(n413), .B(n412), .S(n451), .Z(n414) );
  MUX2_X1 U457 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n453), .Z(n415) );
  MUX2_X1 U458 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n453), .Z(n416) );
  MUX2_X1 U459 ( .A(n416), .B(n415), .S(n451), .Z(n417) );
  MUX2_X1 U460 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n453), .Z(n418) );
  MUX2_X1 U461 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n453), .Z(n419) );
  MUX2_X1 U462 ( .A(n419), .B(n418), .S(N11), .Z(n420) );
  MUX2_X1 U463 ( .A(n420), .B(n417), .S(N12), .Z(N18) );
  MUX2_X1 U464 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n453), .Z(n421) );
  MUX2_X1 U465 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n453), .Z(n422) );
  MUX2_X1 U466 ( .A(n422), .B(n421), .S(n451), .Z(n423) );
  MUX2_X1 U467 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n453), .Z(n424) );
  MUX2_X1 U468 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n453), .Z(n425) );
  MUX2_X1 U469 ( .A(n425), .B(n424), .S(n451), .Z(n426) );
  MUX2_X1 U470 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n453), .Z(n427) );
  MUX2_X1 U471 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n453), .Z(n428) );
  MUX2_X1 U472 ( .A(n428), .B(n427), .S(n451), .Z(n429) );
  MUX2_X1 U473 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n453), .Z(n430) );
  MUX2_X1 U474 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n453), .Z(n431) );
  MUX2_X1 U475 ( .A(n431), .B(n430), .S(n451), .Z(n432) );
  MUX2_X1 U476 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n454), .Z(n433) );
  MUX2_X1 U477 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n454), .Z(n434) );
  MUX2_X1 U478 ( .A(n434), .B(n433), .S(n451), .Z(n435) );
  MUX2_X1 U479 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n454), .Z(n436) );
  MUX2_X1 U480 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n454), .Z(n437) );
  MUX2_X1 U481 ( .A(n437), .B(n436), .S(n451), .Z(n438) );
  MUX2_X1 U482 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n454), .Z(n439) );
  MUX2_X1 U483 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n454), .Z(n440) );
  MUX2_X1 U484 ( .A(n440), .B(n439), .S(N11), .Z(n441) );
  MUX2_X1 U485 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n454), .Z(n442) );
  MUX2_X1 U486 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n454), .Z(n443) );
  MUX2_X1 U487 ( .A(n443), .B(n442), .S(n451), .Z(n444) );
  MUX2_X1 U488 ( .A(n444), .B(n441), .S(N12), .Z(N14) );
  MUX2_X1 U489 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n454), .Z(n445) );
  MUX2_X1 U490 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n454), .Z(n446) );
  MUX2_X1 U491 ( .A(n446), .B(n445), .S(n451), .Z(n447) );
  MUX2_X1 U492 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n454), .Z(n448) );
  MUX2_X1 U493 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n454), .Z(n449) );
  MUX2_X1 U494 ( .A(n449), .B(n448), .S(n451), .Z(n450) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE3_3 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N14, N16, N18, N20, N24, N26, N28, N30, N32, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[18]  ( .D(N14), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[16]  ( .D(N16), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N20), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[8]  ( .D(N24), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N26), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N28), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N30), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N32), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n486), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n487), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n488), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n489), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n490), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n491), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n492), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n493), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n494), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n495), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n496), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n497), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n498), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n499), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n500), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n501), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n502), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n503), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n504), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n505), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n506), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n507), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n508), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n509), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n510), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n511), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n512), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n513), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n514), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n515), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n516), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n517), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n518), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n519), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n520), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n521), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n522), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n523), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n524), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n525), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n526), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n527), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n528), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n529), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n530), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n531), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n532), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n533), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n534), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n535), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n536), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n537), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n538), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n539), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n540), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n541), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n542), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n543), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n544), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n545), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n546), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n547), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n548), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n549), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n550), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n551), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n552), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n553), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n554), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n555), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n556), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n557), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n558), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n559), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n560), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n561), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n562), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n563), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n564), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n565), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n566), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n567), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n568), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n569), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n570), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n571), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n572), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n573), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n574), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n575), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n576), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n577), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n578), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n579), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n580), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n581), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n582), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n583), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n584), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n585), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n586), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n587), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n588), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n589), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n590), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n591), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n592), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n593), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n594), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n595), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n596), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n597), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n598), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n599), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n600), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n601), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n602), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n603), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n604), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n605), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n606), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n607), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n608), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n609), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n610), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n611), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n612), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n613), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n614), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n615), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n616), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n617), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n618), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n619), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n620), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n621), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n622), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n623), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n624), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n625), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n626), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n627), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n628), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n629), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n630), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n631), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n632), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n633), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n634), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n635), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n636), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n637), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n638), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n639), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n640), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n641), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n642), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n643), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n644), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n645), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U348 ( .A1(n463), .A2(n464), .A3(n794), .ZN(n815) );
  NAND3_X1 U349 ( .A1(n794), .A2(n464), .A3(N10), .ZN(n793) );
  NAND3_X1 U350 ( .A1(n794), .A2(n463), .A3(N11), .ZN(n772) );
  NAND3_X1 U351 ( .A1(N10), .A2(n794), .A3(N11), .ZN(n751) );
  NAND3_X1 U352 ( .A1(n463), .A2(n464), .A3(n709), .ZN(n730) );
  NAND3_X1 U353 ( .A1(N10), .A2(n464), .A3(n709), .ZN(n708) );
  NAND3_X1 U354 ( .A1(N11), .A2(n463), .A3(n709), .ZN(n687) );
  NAND3_X1 U355 ( .A1(N11), .A2(N10), .A3(n709), .ZN(n666) );
  SDFF_X1 \data_out_reg[13]  ( .D(n414), .SI(n411), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n12), .SI(n9), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n402), .SI(n399), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[17]  ( .D(n438), .SI(n435), .SE(N12), .CK(clk), .Q(
        data_out[17]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n390), .SI(n387), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n366), .SI(n363), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n354), .SI(n21), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n378), .SI(n375), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n426), .SI(n423), .SE(N12), .CK(clk), .Q(
        data_out[15]) );
  SDFF_X1 \data_out_reg[19]  ( .D(n450), .SI(n447), .SE(N12), .CK(clk), .Q(
        data_out[19]) );
  SDFF_X1 \data_out_reg[10]  ( .D(n396), .SI(n393), .SE(N12), .CK(clk), .Q(
        data_out[10]) );
  BUF_X1 U3 ( .A(n772), .Z(n460) );
  BUF_X1 U4 ( .A(n730), .Z(n458) );
  BUF_X1 U5 ( .A(N11), .Z(n451) );
  BUF_X1 U6 ( .A(n815), .Z(n462) );
  BUF_X1 U7 ( .A(n751), .Z(n459) );
  BUF_X1 U8 ( .A(n793), .Z(n461) );
  BUF_X1 U9 ( .A(n666), .Z(n455) );
  BUF_X1 U10 ( .A(n708), .Z(n457) );
  BUF_X1 U11 ( .A(n687), .Z(n456) );
  BUF_X1 U12 ( .A(N10), .Z(n453) );
  BUF_X1 U13 ( .A(N10), .Z(n454) );
  NOR2_X1 U14 ( .A1(n465), .A2(N12), .ZN(n794) );
  INV_X1 U15 ( .A(wr_en), .ZN(n465) );
  AND2_X1 U16 ( .A1(N12), .A2(wr_en), .ZN(n709) );
  OAI21_X1 U17 ( .B1(n485), .B2(n793), .A(n792), .ZN(n625) );
  NAND2_X1 U18 ( .A1(\mem[1][0] ), .A2(n461), .ZN(n792) );
  OAI21_X1 U19 ( .B1(n484), .B2(n793), .A(n791), .ZN(n624) );
  NAND2_X1 U20 ( .A1(\mem[1][1] ), .A2(n461), .ZN(n791) );
  OAI21_X1 U21 ( .B1(n483), .B2(n793), .A(n790), .ZN(n623) );
  NAND2_X1 U22 ( .A1(\mem[1][2] ), .A2(n461), .ZN(n790) );
  OAI21_X1 U23 ( .B1(n482), .B2(n793), .A(n789), .ZN(n622) );
  NAND2_X1 U24 ( .A1(\mem[1][3] ), .A2(n461), .ZN(n789) );
  OAI21_X1 U25 ( .B1(n481), .B2(n461), .A(n788), .ZN(n621) );
  NAND2_X1 U26 ( .A1(\mem[1][4] ), .A2(n461), .ZN(n788) );
  OAI21_X1 U27 ( .B1(n480), .B2(n461), .A(n787), .ZN(n620) );
  NAND2_X1 U28 ( .A1(\mem[1][5] ), .A2(n461), .ZN(n787) );
  OAI21_X1 U29 ( .B1(n479), .B2(n793), .A(n786), .ZN(n619) );
  NAND2_X1 U30 ( .A1(\mem[1][6] ), .A2(n461), .ZN(n786) );
  OAI21_X1 U31 ( .B1(n478), .B2(n793), .A(n785), .ZN(n618) );
  NAND2_X1 U32 ( .A1(\mem[1][7] ), .A2(n461), .ZN(n785) );
  OAI21_X1 U33 ( .B1(n477), .B2(n793), .A(n784), .ZN(n617) );
  NAND2_X1 U34 ( .A1(\mem[1][8] ), .A2(n461), .ZN(n784) );
  OAI21_X1 U35 ( .B1(n476), .B2(n793), .A(n783), .ZN(n616) );
  NAND2_X1 U36 ( .A1(\mem[1][9] ), .A2(n461), .ZN(n783) );
  OAI21_X1 U37 ( .B1(n475), .B2(n793), .A(n782), .ZN(n615) );
  NAND2_X1 U38 ( .A1(\mem[1][10] ), .A2(n461), .ZN(n782) );
  OAI21_X1 U39 ( .B1(n474), .B2(n793), .A(n781), .ZN(n614) );
  NAND2_X1 U40 ( .A1(\mem[1][11] ), .A2(n461), .ZN(n781) );
  OAI21_X1 U41 ( .B1(n473), .B2(n793), .A(n780), .ZN(n613) );
  NAND2_X1 U42 ( .A1(\mem[1][12] ), .A2(n793), .ZN(n780) );
  OAI21_X1 U43 ( .B1(n472), .B2(n793), .A(n779), .ZN(n612) );
  NAND2_X1 U44 ( .A1(\mem[1][13] ), .A2(n793), .ZN(n779) );
  OAI21_X1 U45 ( .B1(n471), .B2(n793), .A(n778), .ZN(n611) );
  NAND2_X1 U46 ( .A1(\mem[1][14] ), .A2(n793), .ZN(n778) );
  OAI21_X1 U47 ( .B1(n470), .B2(n793), .A(n777), .ZN(n610) );
  NAND2_X1 U48 ( .A1(\mem[1][15] ), .A2(n461), .ZN(n777) );
  OAI21_X1 U49 ( .B1(n469), .B2(n793), .A(n776), .ZN(n609) );
  NAND2_X1 U50 ( .A1(\mem[1][16] ), .A2(n793), .ZN(n776) );
  OAI21_X1 U51 ( .B1(n468), .B2(n793), .A(n775), .ZN(n608) );
  NAND2_X1 U52 ( .A1(\mem[1][17] ), .A2(n793), .ZN(n775) );
  OAI21_X1 U53 ( .B1(n467), .B2(n793), .A(n774), .ZN(n607) );
  NAND2_X1 U54 ( .A1(\mem[1][18] ), .A2(n793), .ZN(n774) );
  OAI21_X1 U55 ( .B1(n466), .B2(n793), .A(n773), .ZN(n606) );
  NAND2_X1 U56 ( .A1(\mem[1][19] ), .A2(n461), .ZN(n773) );
  OAI21_X1 U57 ( .B1(n485), .B2(n772), .A(n771), .ZN(n605) );
  NAND2_X1 U58 ( .A1(\mem[2][0] ), .A2(n460), .ZN(n771) );
  OAI21_X1 U59 ( .B1(n484), .B2(n772), .A(n770), .ZN(n604) );
  NAND2_X1 U60 ( .A1(\mem[2][1] ), .A2(n460), .ZN(n770) );
  OAI21_X1 U61 ( .B1(n483), .B2(n772), .A(n769), .ZN(n603) );
  NAND2_X1 U62 ( .A1(\mem[2][2] ), .A2(n460), .ZN(n769) );
  OAI21_X1 U63 ( .B1(n482), .B2(n772), .A(n768), .ZN(n602) );
  NAND2_X1 U64 ( .A1(\mem[2][3] ), .A2(n460), .ZN(n768) );
  OAI21_X1 U65 ( .B1(n481), .B2(n460), .A(n767), .ZN(n601) );
  NAND2_X1 U66 ( .A1(\mem[2][4] ), .A2(n460), .ZN(n767) );
  OAI21_X1 U67 ( .B1(n480), .B2(n772), .A(n766), .ZN(n600) );
  NAND2_X1 U68 ( .A1(\mem[2][5] ), .A2(n460), .ZN(n766) );
  OAI21_X1 U69 ( .B1(n479), .B2(n460), .A(n765), .ZN(n599) );
  NAND2_X1 U70 ( .A1(\mem[2][6] ), .A2(n460), .ZN(n765) );
  OAI21_X1 U71 ( .B1(n478), .B2(n772), .A(n764), .ZN(n598) );
  NAND2_X1 U72 ( .A1(\mem[2][7] ), .A2(n460), .ZN(n764) );
  OAI21_X1 U73 ( .B1(n477), .B2(n772), .A(n763), .ZN(n597) );
  NAND2_X1 U74 ( .A1(\mem[2][8] ), .A2(n460), .ZN(n763) );
  OAI21_X1 U75 ( .B1(n476), .B2(n772), .A(n762), .ZN(n596) );
  NAND2_X1 U76 ( .A1(\mem[2][9] ), .A2(n460), .ZN(n762) );
  OAI21_X1 U77 ( .B1(n475), .B2(n772), .A(n761), .ZN(n595) );
  NAND2_X1 U78 ( .A1(\mem[2][10] ), .A2(n460), .ZN(n761) );
  OAI21_X1 U79 ( .B1(n474), .B2(n772), .A(n760), .ZN(n594) );
  NAND2_X1 U80 ( .A1(\mem[2][11] ), .A2(n460), .ZN(n760) );
  OAI21_X1 U81 ( .B1(n473), .B2(n772), .A(n759), .ZN(n593) );
  NAND2_X1 U82 ( .A1(\mem[2][12] ), .A2(n460), .ZN(n759) );
  OAI21_X1 U83 ( .B1(n472), .B2(n772), .A(n758), .ZN(n592) );
  NAND2_X1 U84 ( .A1(\mem[2][13] ), .A2(n772), .ZN(n758) );
  OAI21_X1 U85 ( .B1(n471), .B2(n772), .A(n757), .ZN(n591) );
  NAND2_X1 U86 ( .A1(\mem[2][14] ), .A2(n772), .ZN(n757) );
  OAI21_X1 U87 ( .B1(n470), .B2(n772), .A(n756), .ZN(n590) );
  NAND2_X1 U88 ( .A1(\mem[2][15] ), .A2(n772), .ZN(n756) );
  OAI21_X1 U89 ( .B1(n469), .B2(n772), .A(n755), .ZN(n589) );
  NAND2_X1 U90 ( .A1(\mem[2][16] ), .A2(n772), .ZN(n755) );
  OAI21_X1 U91 ( .B1(n468), .B2(n772), .A(n754), .ZN(n588) );
  NAND2_X1 U92 ( .A1(\mem[2][17] ), .A2(n772), .ZN(n754) );
  OAI21_X1 U93 ( .B1(n467), .B2(n772), .A(n753), .ZN(n587) );
  NAND2_X1 U94 ( .A1(\mem[2][18] ), .A2(n772), .ZN(n753) );
  OAI21_X1 U95 ( .B1(n466), .B2(n460), .A(n752), .ZN(n586) );
  NAND2_X1 U96 ( .A1(\mem[2][19] ), .A2(n460), .ZN(n752) );
  OAI21_X1 U97 ( .B1(n485), .B2(n751), .A(n750), .ZN(n585) );
  NAND2_X1 U98 ( .A1(\mem[3][0] ), .A2(n459), .ZN(n750) );
  OAI21_X1 U99 ( .B1(n484), .B2(n751), .A(n749), .ZN(n584) );
  NAND2_X1 U100 ( .A1(\mem[3][1] ), .A2(n459), .ZN(n749) );
  OAI21_X1 U101 ( .B1(n483), .B2(n751), .A(n748), .ZN(n583) );
  NAND2_X1 U102 ( .A1(\mem[3][2] ), .A2(n459), .ZN(n748) );
  OAI21_X1 U103 ( .B1(n482), .B2(n751), .A(n747), .ZN(n582) );
  NAND2_X1 U104 ( .A1(\mem[3][3] ), .A2(n459), .ZN(n747) );
  OAI21_X1 U105 ( .B1(n481), .B2(n459), .A(n746), .ZN(n581) );
  NAND2_X1 U106 ( .A1(\mem[3][4] ), .A2(n459), .ZN(n746) );
  OAI21_X1 U107 ( .B1(n480), .B2(n459), .A(n745), .ZN(n580) );
  NAND2_X1 U108 ( .A1(\mem[3][5] ), .A2(n459), .ZN(n745) );
  OAI21_X1 U109 ( .B1(n479), .B2(n751), .A(n744), .ZN(n579) );
  NAND2_X1 U110 ( .A1(\mem[3][6] ), .A2(n459), .ZN(n744) );
  OAI21_X1 U111 ( .B1(n478), .B2(n751), .A(n743), .ZN(n578) );
  NAND2_X1 U112 ( .A1(\mem[3][7] ), .A2(n459), .ZN(n743) );
  OAI21_X1 U113 ( .B1(n477), .B2(n751), .A(n742), .ZN(n577) );
  NAND2_X1 U114 ( .A1(\mem[3][8] ), .A2(n459), .ZN(n742) );
  OAI21_X1 U115 ( .B1(n476), .B2(n751), .A(n741), .ZN(n576) );
  NAND2_X1 U116 ( .A1(\mem[3][9] ), .A2(n459), .ZN(n741) );
  OAI21_X1 U117 ( .B1(n475), .B2(n751), .A(n740), .ZN(n575) );
  NAND2_X1 U118 ( .A1(\mem[3][10] ), .A2(n459), .ZN(n740) );
  OAI21_X1 U119 ( .B1(n474), .B2(n751), .A(n739), .ZN(n574) );
  NAND2_X1 U120 ( .A1(\mem[3][11] ), .A2(n459), .ZN(n739) );
  OAI21_X1 U121 ( .B1(n473), .B2(n751), .A(n738), .ZN(n573) );
  NAND2_X1 U122 ( .A1(\mem[3][12] ), .A2(n751), .ZN(n738) );
  OAI21_X1 U123 ( .B1(n472), .B2(n751), .A(n737), .ZN(n572) );
  NAND2_X1 U124 ( .A1(\mem[3][13] ), .A2(n751), .ZN(n737) );
  OAI21_X1 U125 ( .B1(n471), .B2(n751), .A(n736), .ZN(n571) );
  NAND2_X1 U126 ( .A1(\mem[3][14] ), .A2(n751), .ZN(n736) );
  OAI21_X1 U127 ( .B1(n470), .B2(n751), .A(n735), .ZN(n570) );
  NAND2_X1 U128 ( .A1(\mem[3][15] ), .A2(n459), .ZN(n735) );
  OAI21_X1 U129 ( .B1(n469), .B2(n751), .A(n734), .ZN(n569) );
  NAND2_X1 U130 ( .A1(\mem[3][16] ), .A2(n751), .ZN(n734) );
  OAI21_X1 U131 ( .B1(n468), .B2(n751), .A(n733), .ZN(n568) );
  NAND2_X1 U132 ( .A1(\mem[3][17] ), .A2(n751), .ZN(n733) );
  OAI21_X1 U133 ( .B1(n467), .B2(n751), .A(n732), .ZN(n567) );
  NAND2_X1 U134 ( .A1(\mem[3][18] ), .A2(n751), .ZN(n732) );
  OAI21_X1 U135 ( .B1(n466), .B2(n751), .A(n731), .ZN(n566) );
  NAND2_X1 U136 ( .A1(\mem[3][19] ), .A2(n459), .ZN(n731) );
  OAI21_X1 U137 ( .B1(n485), .B2(n458), .A(n729), .ZN(n565) );
  NAND2_X1 U138 ( .A1(\mem[4][0] ), .A2(n458), .ZN(n729) );
  OAI21_X1 U139 ( .B1(n484), .B2(n458), .A(n728), .ZN(n564) );
  NAND2_X1 U140 ( .A1(\mem[4][1] ), .A2(n458), .ZN(n728) );
  OAI21_X1 U141 ( .B1(n483), .B2(n458), .A(n727), .ZN(n563) );
  NAND2_X1 U142 ( .A1(\mem[4][2] ), .A2(n730), .ZN(n727) );
  OAI21_X1 U143 ( .B1(n482), .B2(n730), .A(n726), .ZN(n562) );
  NAND2_X1 U144 ( .A1(\mem[4][3] ), .A2(n458), .ZN(n726) );
  OAI21_X1 U145 ( .B1(n481), .B2(n730), .A(n725), .ZN(n561) );
  NAND2_X1 U146 ( .A1(\mem[4][4] ), .A2(n730), .ZN(n725) );
  OAI21_X1 U147 ( .B1(n480), .B2(n730), .A(n724), .ZN(n560) );
  NAND2_X1 U148 ( .A1(\mem[4][5] ), .A2(n730), .ZN(n724) );
  OAI21_X1 U149 ( .B1(n479), .B2(n730), .A(n723), .ZN(n559) );
  NAND2_X1 U150 ( .A1(\mem[4][6] ), .A2(n730), .ZN(n723) );
  OAI21_X1 U151 ( .B1(n478), .B2(n730), .A(n722), .ZN(n558) );
  NAND2_X1 U152 ( .A1(\mem[4][7] ), .A2(n730), .ZN(n722) );
  OAI21_X1 U153 ( .B1(n477), .B2(n730), .A(n721), .ZN(n557) );
  NAND2_X1 U154 ( .A1(\mem[4][8] ), .A2(n730), .ZN(n721) );
  OAI21_X1 U155 ( .B1(n476), .B2(n458), .A(n720), .ZN(n556) );
  NAND2_X1 U156 ( .A1(\mem[4][9] ), .A2(n730), .ZN(n720) );
  OAI21_X1 U157 ( .B1(n475), .B2(n730), .A(n719), .ZN(n555) );
  NAND2_X1 U158 ( .A1(\mem[4][10] ), .A2(n730), .ZN(n719) );
  OAI21_X1 U159 ( .B1(n474), .B2(n730), .A(n718), .ZN(n554) );
  NAND2_X1 U160 ( .A1(\mem[4][11] ), .A2(n730), .ZN(n718) );
  OAI21_X1 U161 ( .B1(n473), .B2(n458), .A(n717), .ZN(n553) );
  NAND2_X1 U162 ( .A1(\mem[4][12] ), .A2(n458), .ZN(n717) );
  OAI21_X1 U163 ( .B1(n472), .B2(n458), .A(n716), .ZN(n552) );
  NAND2_X1 U164 ( .A1(\mem[4][13] ), .A2(n458), .ZN(n716) );
  OAI21_X1 U165 ( .B1(n471), .B2(n458), .A(n715), .ZN(n551) );
  NAND2_X1 U166 ( .A1(\mem[4][14] ), .A2(n458), .ZN(n715) );
  OAI21_X1 U167 ( .B1(n470), .B2(n730), .A(n714), .ZN(n550) );
  NAND2_X1 U168 ( .A1(\mem[4][15] ), .A2(n458), .ZN(n714) );
  OAI21_X1 U169 ( .B1(n469), .B2(n730), .A(n713), .ZN(n549) );
  NAND2_X1 U170 ( .A1(\mem[4][16] ), .A2(n458), .ZN(n713) );
  OAI21_X1 U171 ( .B1(n468), .B2(n730), .A(n712), .ZN(n548) );
  NAND2_X1 U172 ( .A1(\mem[4][17] ), .A2(n458), .ZN(n712) );
  OAI21_X1 U173 ( .B1(n467), .B2(n458), .A(n711), .ZN(n547) );
  NAND2_X1 U174 ( .A1(\mem[4][18] ), .A2(n458), .ZN(n711) );
  OAI21_X1 U175 ( .B1(n466), .B2(n458), .A(n710), .ZN(n546) );
  NAND2_X1 U176 ( .A1(\mem[4][19] ), .A2(n458), .ZN(n710) );
  OAI21_X1 U177 ( .B1(n485), .B2(n708), .A(n707), .ZN(n545) );
  NAND2_X1 U178 ( .A1(\mem[5][0] ), .A2(n457), .ZN(n707) );
  OAI21_X1 U179 ( .B1(n484), .B2(n708), .A(n706), .ZN(n544) );
  NAND2_X1 U180 ( .A1(\mem[5][1] ), .A2(n457), .ZN(n706) );
  OAI21_X1 U181 ( .B1(n483), .B2(n708), .A(n705), .ZN(n543) );
  NAND2_X1 U182 ( .A1(\mem[5][2] ), .A2(n457), .ZN(n705) );
  OAI21_X1 U183 ( .B1(n482), .B2(n708), .A(n704), .ZN(n542) );
  NAND2_X1 U184 ( .A1(\mem[5][3] ), .A2(n457), .ZN(n704) );
  OAI21_X1 U185 ( .B1(n481), .B2(n457), .A(n703), .ZN(n541) );
  NAND2_X1 U186 ( .A1(\mem[5][4] ), .A2(n457), .ZN(n703) );
  OAI21_X1 U187 ( .B1(n480), .B2(n708), .A(n702), .ZN(n540) );
  NAND2_X1 U188 ( .A1(\mem[5][5] ), .A2(n457), .ZN(n702) );
  OAI21_X1 U189 ( .B1(n479), .B2(n708), .A(n701), .ZN(n539) );
  NAND2_X1 U190 ( .A1(\mem[5][6] ), .A2(n457), .ZN(n701) );
  OAI21_X1 U191 ( .B1(n478), .B2(n708), .A(n700), .ZN(n538) );
  NAND2_X1 U192 ( .A1(\mem[5][7] ), .A2(n457), .ZN(n700) );
  OAI21_X1 U193 ( .B1(n477), .B2(n708), .A(n699), .ZN(n537) );
  NAND2_X1 U194 ( .A1(\mem[5][8] ), .A2(n457), .ZN(n699) );
  OAI21_X1 U195 ( .B1(n476), .B2(n708), .A(n698), .ZN(n536) );
  NAND2_X1 U196 ( .A1(\mem[5][9] ), .A2(n457), .ZN(n698) );
  OAI21_X1 U197 ( .B1(n475), .B2(n708), .A(n697), .ZN(n535) );
  NAND2_X1 U198 ( .A1(\mem[5][10] ), .A2(n457), .ZN(n697) );
  OAI21_X1 U199 ( .B1(n474), .B2(n708), .A(n696), .ZN(n534) );
  NAND2_X1 U200 ( .A1(\mem[5][11] ), .A2(n457), .ZN(n696) );
  OAI21_X1 U201 ( .B1(n473), .B2(n708), .A(n695), .ZN(n533) );
  NAND2_X1 U202 ( .A1(\mem[5][12] ), .A2(n708), .ZN(n695) );
  OAI21_X1 U203 ( .B1(n472), .B2(n457), .A(n694), .ZN(n532) );
  NAND2_X1 U204 ( .A1(\mem[5][13] ), .A2(n708), .ZN(n694) );
  OAI21_X1 U205 ( .B1(n471), .B2(n457), .A(n693), .ZN(n531) );
  NAND2_X1 U206 ( .A1(\mem[5][14] ), .A2(n708), .ZN(n693) );
  OAI21_X1 U207 ( .B1(n470), .B2(n708), .A(n692), .ZN(n530) );
  NAND2_X1 U208 ( .A1(\mem[5][15] ), .A2(n708), .ZN(n692) );
  OAI21_X1 U209 ( .B1(n469), .B2(n708), .A(n691), .ZN(n529) );
  NAND2_X1 U210 ( .A1(\mem[5][16] ), .A2(n708), .ZN(n691) );
  OAI21_X1 U211 ( .B1(n468), .B2(n708), .A(n690), .ZN(n528) );
  NAND2_X1 U212 ( .A1(\mem[5][17] ), .A2(n708), .ZN(n690) );
  OAI21_X1 U213 ( .B1(n467), .B2(n708), .A(n689), .ZN(n527) );
  NAND2_X1 U214 ( .A1(\mem[5][18] ), .A2(n708), .ZN(n689) );
  OAI21_X1 U215 ( .B1(n466), .B2(n708), .A(n688), .ZN(n526) );
  NAND2_X1 U216 ( .A1(\mem[5][19] ), .A2(n457), .ZN(n688) );
  OAI21_X1 U217 ( .B1(n485), .B2(n687), .A(n686), .ZN(n525) );
  NAND2_X1 U218 ( .A1(\mem[6][0] ), .A2(n687), .ZN(n686) );
  OAI21_X1 U219 ( .B1(n484), .B2(n687), .A(n685), .ZN(n524) );
  NAND2_X1 U220 ( .A1(\mem[6][1] ), .A2(n687), .ZN(n685) );
  OAI21_X1 U221 ( .B1(n483), .B2(n687), .A(n684), .ZN(n523) );
  NAND2_X1 U222 ( .A1(\mem[6][2] ), .A2(n687), .ZN(n684) );
  OAI21_X1 U223 ( .B1(n482), .B2(n456), .A(n683), .ZN(n522) );
  NAND2_X1 U224 ( .A1(\mem[6][3] ), .A2(n456), .ZN(n683) );
  OAI21_X1 U225 ( .B1(n481), .B2(n687), .A(n682), .ZN(n521) );
  NAND2_X1 U226 ( .A1(\mem[6][4] ), .A2(n456), .ZN(n682) );
  OAI21_X1 U227 ( .B1(n480), .B2(n687), .A(n681), .ZN(n520) );
  NAND2_X1 U228 ( .A1(\mem[6][5] ), .A2(n687), .ZN(n681) );
  OAI21_X1 U229 ( .B1(n479), .B2(n687), .A(n680), .ZN(n519) );
  NAND2_X1 U230 ( .A1(\mem[6][6] ), .A2(n687), .ZN(n680) );
  OAI21_X1 U231 ( .B1(n478), .B2(n456), .A(n679), .ZN(n518) );
  NAND2_X1 U232 ( .A1(\mem[6][7] ), .A2(n687), .ZN(n679) );
  OAI21_X1 U233 ( .B1(n477), .B2(n456), .A(n678), .ZN(n517) );
  NAND2_X1 U234 ( .A1(\mem[6][8] ), .A2(n687), .ZN(n678) );
  OAI21_X1 U235 ( .B1(n476), .B2(n456), .A(n677), .ZN(n516) );
  NAND2_X1 U236 ( .A1(\mem[6][9] ), .A2(n687), .ZN(n677) );
  OAI21_X1 U237 ( .B1(n475), .B2(n456), .A(n676), .ZN(n515) );
  NAND2_X1 U238 ( .A1(\mem[6][10] ), .A2(n687), .ZN(n676) );
  OAI21_X1 U239 ( .B1(n474), .B2(n456), .A(n675), .ZN(n514) );
  NAND2_X1 U240 ( .A1(\mem[6][11] ), .A2(n687), .ZN(n675) );
  OAI21_X1 U241 ( .B1(n473), .B2(n687), .A(n674), .ZN(n513) );
  NAND2_X1 U242 ( .A1(\mem[6][12] ), .A2(n456), .ZN(n674) );
  OAI21_X1 U243 ( .B1(n472), .B2(n687), .A(n673), .ZN(n512) );
  NAND2_X1 U244 ( .A1(\mem[6][13] ), .A2(n456), .ZN(n673) );
  OAI21_X1 U245 ( .B1(n471), .B2(n687), .A(n672), .ZN(n511) );
  NAND2_X1 U246 ( .A1(\mem[6][14] ), .A2(n456), .ZN(n672) );
  OAI21_X1 U247 ( .B1(n470), .B2(n687), .A(n671), .ZN(n510) );
  NAND2_X1 U248 ( .A1(\mem[6][15] ), .A2(n456), .ZN(n671) );
  OAI21_X1 U249 ( .B1(n469), .B2(n687), .A(n670), .ZN(n509) );
  NAND2_X1 U250 ( .A1(\mem[6][16] ), .A2(n456), .ZN(n670) );
  OAI21_X1 U251 ( .B1(n468), .B2(n687), .A(n669), .ZN(n508) );
  NAND2_X1 U252 ( .A1(\mem[6][17] ), .A2(n456), .ZN(n669) );
  OAI21_X1 U253 ( .B1(n467), .B2(n687), .A(n668), .ZN(n507) );
  NAND2_X1 U254 ( .A1(\mem[6][18] ), .A2(n456), .ZN(n668) );
  OAI21_X1 U255 ( .B1(n466), .B2(n687), .A(n667), .ZN(n506) );
  NAND2_X1 U256 ( .A1(\mem[6][19] ), .A2(n456), .ZN(n667) );
  OAI21_X1 U257 ( .B1(n485), .B2(n666), .A(n665), .ZN(n505) );
  NAND2_X1 U258 ( .A1(\mem[7][0] ), .A2(n455), .ZN(n665) );
  OAI21_X1 U259 ( .B1(n484), .B2(n666), .A(n664), .ZN(n504) );
  NAND2_X1 U260 ( .A1(\mem[7][1] ), .A2(n455), .ZN(n664) );
  OAI21_X1 U261 ( .B1(n483), .B2(n666), .A(n663), .ZN(n503) );
  NAND2_X1 U262 ( .A1(\mem[7][2] ), .A2(n455), .ZN(n663) );
  OAI21_X1 U263 ( .B1(n482), .B2(n666), .A(n662), .ZN(n502) );
  NAND2_X1 U264 ( .A1(\mem[7][3] ), .A2(n455), .ZN(n662) );
  OAI21_X1 U265 ( .B1(n481), .B2(n455), .A(n661), .ZN(n501) );
  NAND2_X1 U266 ( .A1(\mem[7][4] ), .A2(n455), .ZN(n661) );
  OAI21_X1 U267 ( .B1(n480), .B2(n666), .A(n660), .ZN(n500) );
  NAND2_X1 U268 ( .A1(\mem[7][5] ), .A2(n455), .ZN(n660) );
  OAI21_X1 U269 ( .B1(n479), .B2(n666), .A(n659), .ZN(n499) );
  NAND2_X1 U270 ( .A1(\mem[7][6] ), .A2(n455), .ZN(n659) );
  OAI21_X1 U271 ( .B1(n478), .B2(n666), .A(n658), .ZN(n498) );
  NAND2_X1 U272 ( .A1(\mem[7][7] ), .A2(n455), .ZN(n658) );
  OAI21_X1 U273 ( .B1(n477), .B2(n666), .A(n657), .ZN(n497) );
  NAND2_X1 U274 ( .A1(\mem[7][8] ), .A2(n455), .ZN(n657) );
  OAI21_X1 U275 ( .B1(n476), .B2(n666), .A(n656), .ZN(n496) );
  NAND2_X1 U276 ( .A1(\mem[7][9] ), .A2(n455), .ZN(n656) );
  OAI21_X1 U277 ( .B1(n475), .B2(n666), .A(n655), .ZN(n495) );
  NAND2_X1 U278 ( .A1(\mem[7][10] ), .A2(n455), .ZN(n655) );
  OAI21_X1 U279 ( .B1(n474), .B2(n666), .A(n654), .ZN(n494) );
  NAND2_X1 U280 ( .A1(\mem[7][11] ), .A2(n455), .ZN(n654) );
  OAI21_X1 U281 ( .B1(n473), .B2(n666), .A(n653), .ZN(n493) );
  NAND2_X1 U282 ( .A1(\mem[7][12] ), .A2(n666), .ZN(n653) );
  OAI21_X1 U283 ( .B1(n472), .B2(n455), .A(n652), .ZN(n492) );
  NAND2_X1 U284 ( .A1(\mem[7][13] ), .A2(n666), .ZN(n652) );
  OAI21_X1 U285 ( .B1(n471), .B2(n455), .A(n651), .ZN(n491) );
  NAND2_X1 U286 ( .A1(\mem[7][14] ), .A2(n666), .ZN(n651) );
  OAI21_X1 U287 ( .B1(n470), .B2(n666), .A(n650), .ZN(n490) );
  NAND2_X1 U288 ( .A1(\mem[7][15] ), .A2(n666), .ZN(n650) );
  OAI21_X1 U289 ( .B1(n469), .B2(n666), .A(n649), .ZN(n489) );
  NAND2_X1 U290 ( .A1(\mem[7][16] ), .A2(n666), .ZN(n649) );
  OAI21_X1 U291 ( .B1(n468), .B2(n666), .A(n648), .ZN(n488) );
  NAND2_X1 U292 ( .A1(\mem[7][17] ), .A2(n666), .ZN(n648) );
  OAI21_X1 U293 ( .B1(n467), .B2(n666), .A(n647), .ZN(n487) );
  NAND2_X1 U294 ( .A1(\mem[7][18] ), .A2(n666), .ZN(n647) );
  OAI21_X1 U295 ( .B1(n466), .B2(n666), .A(n646), .ZN(n486) );
  NAND2_X1 U296 ( .A1(\mem[7][19] ), .A2(n455), .ZN(n646) );
  OAI21_X1 U297 ( .B1(n815), .B2(n483), .A(n812), .ZN(n643) );
  NAND2_X1 U298 ( .A1(\mem[0][2] ), .A2(n462), .ZN(n812) );
  OAI21_X1 U299 ( .B1(n815), .B2(n482), .A(n811), .ZN(n642) );
  NAND2_X1 U300 ( .A1(\mem[0][3] ), .A2(n462), .ZN(n811) );
  OAI21_X1 U301 ( .B1(n815), .B2(n481), .A(n810), .ZN(n641) );
  NAND2_X1 U302 ( .A1(\mem[0][4] ), .A2(n462), .ZN(n810) );
  OAI21_X1 U303 ( .B1(n815), .B2(n480), .A(n809), .ZN(n640) );
  NAND2_X1 U304 ( .A1(\mem[0][5] ), .A2(n462), .ZN(n809) );
  OAI21_X1 U305 ( .B1(n815), .B2(n479), .A(n808), .ZN(n639) );
  NAND2_X1 U306 ( .A1(\mem[0][6] ), .A2(n462), .ZN(n808) );
  OAI21_X1 U307 ( .B1(n815), .B2(n478), .A(n807), .ZN(n638) );
  NAND2_X1 U308 ( .A1(\mem[0][7] ), .A2(n462), .ZN(n807) );
  OAI21_X1 U309 ( .B1(n815), .B2(n477), .A(n806), .ZN(n637) );
  NAND2_X1 U310 ( .A1(\mem[0][8] ), .A2(n462), .ZN(n806) );
  OAI21_X1 U311 ( .B1(n815), .B2(n476), .A(n805), .ZN(n636) );
  NAND2_X1 U312 ( .A1(\mem[0][9] ), .A2(n462), .ZN(n805) );
  OAI21_X1 U313 ( .B1(n815), .B2(n475), .A(n804), .ZN(n635) );
  NAND2_X1 U314 ( .A1(\mem[0][10] ), .A2(n462), .ZN(n804) );
  OAI21_X1 U315 ( .B1(n815), .B2(n474), .A(n803), .ZN(n634) );
  NAND2_X1 U316 ( .A1(\mem[0][11] ), .A2(n462), .ZN(n803) );
  OAI21_X1 U317 ( .B1(n815), .B2(n473), .A(n802), .ZN(n633) );
  NAND2_X1 U318 ( .A1(\mem[0][12] ), .A2(n815), .ZN(n802) );
  OAI21_X1 U319 ( .B1(n815), .B2(n472), .A(n801), .ZN(n632) );
  NAND2_X1 U320 ( .A1(\mem[0][13] ), .A2(n815), .ZN(n801) );
  OAI21_X1 U321 ( .B1(n462), .B2(n471), .A(n800), .ZN(n631) );
  NAND2_X1 U322 ( .A1(\mem[0][14] ), .A2(n815), .ZN(n800) );
  OAI21_X1 U323 ( .B1(n815), .B2(n470), .A(n799), .ZN(n630) );
  NAND2_X1 U324 ( .A1(\mem[0][15] ), .A2(n462), .ZN(n799) );
  OAI21_X1 U325 ( .B1(n815), .B2(n469), .A(n798), .ZN(n629) );
  NAND2_X1 U326 ( .A1(\mem[0][16] ), .A2(n815), .ZN(n798) );
  OAI21_X1 U327 ( .B1(n815), .B2(n468), .A(n797), .ZN(n628) );
  NAND2_X1 U328 ( .A1(\mem[0][17] ), .A2(n815), .ZN(n797) );
  OAI21_X1 U329 ( .B1(n815), .B2(n467), .A(n796), .ZN(n627) );
  NAND2_X1 U330 ( .A1(\mem[0][18] ), .A2(n815), .ZN(n796) );
  OAI21_X1 U331 ( .B1(n462), .B2(n485), .A(n814), .ZN(n645) );
  NAND2_X1 U332 ( .A1(\mem[0][0] ), .A2(n462), .ZN(n814) );
  OAI21_X1 U333 ( .B1(n815), .B2(n484), .A(n813), .ZN(n644) );
  NAND2_X1 U334 ( .A1(\mem[0][1] ), .A2(n462), .ZN(n813) );
  OAI21_X1 U335 ( .B1(n815), .B2(n466), .A(n795), .ZN(n626) );
  NAND2_X1 U336 ( .A1(\mem[0][19] ), .A2(n462), .ZN(n795) );
  INV_X1 U337 ( .A(N10), .ZN(n463) );
  INV_X1 U338 ( .A(N11), .ZN(n464) );
  INV_X1 U339 ( .A(data_in[0]), .ZN(n485) );
  INV_X1 U340 ( .A(data_in[1]), .ZN(n484) );
  INV_X1 U341 ( .A(data_in[2]), .ZN(n483) );
  INV_X1 U342 ( .A(data_in[3]), .ZN(n482) );
  INV_X1 U343 ( .A(data_in[4]), .ZN(n481) );
  INV_X1 U344 ( .A(data_in[5]), .ZN(n480) );
  INV_X1 U345 ( .A(data_in[6]), .ZN(n479) );
  INV_X1 U346 ( .A(data_in[7]), .ZN(n478) );
  INV_X1 U347 ( .A(data_in[8]), .ZN(n477) );
  INV_X1 U356 ( .A(data_in[9]), .ZN(n476) );
  INV_X1 U357 ( .A(data_in[10]), .ZN(n475) );
  INV_X1 U358 ( .A(data_in[11]), .ZN(n474) );
  INV_X1 U359 ( .A(data_in[12]), .ZN(n473) );
  INV_X1 U360 ( .A(data_in[13]), .ZN(n472) );
  INV_X1 U361 ( .A(data_in[14]), .ZN(n471) );
  INV_X1 U362 ( .A(data_in[15]), .ZN(n470) );
  INV_X1 U363 ( .A(data_in[16]), .ZN(n469) );
  INV_X1 U364 ( .A(data_in[17]), .ZN(n468) );
  INV_X1 U365 ( .A(data_in[18]), .ZN(n467) );
  INV_X1 U366 ( .A(data_in[19]), .ZN(n466) );
  MUX2_X1 U367 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n452), .Z(n1) );
  MUX2_X1 U368 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n452), .Z(n2) );
  MUX2_X1 U369 ( .A(n2), .B(n1), .S(n451), .Z(n3) );
  MUX2_X1 U370 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n452), .Z(n4) );
  MUX2_X1 U371 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n452), .Z(n5) );
  MUX2_X1 U372 ( .A(n5), .B(n4), .S(n451), .Z(n6) );
  MUX2_X1 U373 ( .A(n6), .B(n3), .S(N12), .Z(N32) );
  MUX2_X1 U374 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n452), .Z(n7) );
  MUX2_X1 U375 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n452), .Z(n8) );
  MUX2_X1 U376 ( .A(n8), .B(n7), .S(n451), .Z(n9) );
  MUX2_X1 U377 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n452), .Z(n10) );
  MUX2_X1 U378 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n452), .Z(n11) );
  MUX2_X1 U379 ( .A(n11), .B(n10), .S(n451), .Z(n12) );
  MUX2_X1 U380 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n452), .Z(n13) );
  MUX2_X1 U381 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n454), .Z(n14) );
  MUX2_X1 U382 ( .A(n14), .B(n13), .S(N11), .Z(n15) );
  MUX2_X1 U383 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n452), .Z(n16) );
  MUX2_X1 U384 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n453), .Z(n17) );
  MUX2_X1 U385 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U386 ( .A(n18), .B(n15), .S(N12), .Z(N30) );
  MUX2_X1 U387 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n452), .Z(n19) );
  MUX2_X1 U388 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n453), .Z(n20) );
  MUX2_X1 U389 ( .A(n20), .B(n19), .S(N11), .Z(n21) );
  MUX2_X1 U390 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n454), .Z(n22) );
  MUX2_X1 U391 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n23) );
  MUX2_X1 U392 ( .A(n23), .B(n22), .S(N11), .Z(n354) );
  MUX2_X1 U393 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n452), .Z(n355) );
  MUX2_X1 U394 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n454), .Z(n356) );
  MUX2_X1 U395 ( .A(n356), .B(n355), .S(N11), .Z(n357) );
  MUX2_X1 U396 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n453), .Z(n358) );
  MUX2_X1 U397 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n453), .Z(n359) );
  MUX2_X1 U398 ( .A(n359), .B(n358), .S(N11), .Z(n360) );
  MUX2_X1 U399 ( .A(n360), .B(n357), .S(N12), .Z(N28) );
  MUX2_X1 U400 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n453), .Z(n361) );
  MUX2_X1 U401 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n453), .Z(n362) );
  MUX2_X1 U402 ( .A(n362), .B(n361), .S(N11), .Z(n363) );
  MUX2_X1 U403 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n453), .Z(n364) );
  MUX2_X1 U404 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n453), .Z(n365) );
  MUX2_X1 U405 ( .A(n365), .B(n364), .S(N11), .Z(n366) );
  MUX2_X1 U406 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n453), .Z(n367) );
  MUX2_X1 U407 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n453), .Z(n368) );
  MUX2_X1 U408 ( .A(n368), .B(n367), .S(N11), .Z(n369) );
  MUX2_X1 U409 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n453), .Z(n370) );
  MUX2_X1 U410 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n453), .Z(n371) );
  MUX2_X1 U411 ( .A(n371), .B(n370), .S(N11), .Z(n372) );
  MUX2_X1 U412 ( .A(n372), .B(n369), .S(N12), .Z(N26) );
  MUX2_X1 U413 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n453), .Z(n373) );
  MUX2_X1 U414 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n453), .Z(n374) );
  MUX2_X1 U415 ( .A(n374), .B(n373), .S(N11), .Z(n375) );
  MUX2_X1 U416 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n453), .Z(n376) );
  MUX2_X1 U417 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n453), .Z(n377) );
  MUX2_X1 U418 ( .A(n377), .B(n376), .S(N11), .Z(n378) );
  MUX2_X1 U419 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n454), .Z(n379) );
  MUX2_X1 U420 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n454), .Z(n380) );
  MUX2_X1 U421 ( .A(n380), .B(n379), .S(N11), .Z(n381) );
  MUX2_X1 U422 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n454), .Z(n382) );
  MUX2_X1 U423 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n454), .Z(n383) );
  MUX2_X1 U424 ( .A(n383), .B(n382), .S(N11), .Z(n384) );
  MUX2_X1 U425 ( .A(n384), .B(n381), .S(N12), .Z(N24) );
  MUX2_X1 U426 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n454), .Z(n385) );
  MUX2_X1 U427 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n454), .Z(n386) );
  MUX2_X1 U428 ( .A(n386), .B(n385), .S(N11), .Z(n387) );
  MUX2_X1 U429 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n454), .Z(n388) );
  MUX2_X1 U430 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n454), .Z(n389) );
  MUX2_X1 U431 ( .A(n389), .B(n388), .S(n451), .Z(n390) );
  MUX2_X1 U432 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n454), .Z(n391) );
  MUX2_X1 U433 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n454), .Z(n392) );
  MUX2_X1 U434 ( .A(n392), .B(n391), .S(n451), .Z(n393) );
  MUX2_X1 U435 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n454), .Z(n394) );
  MUX2_X1 U436 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n454), .Z(n395) );
  MUX2_X1 U437 ( .A(n395), .B(n394), .S(n451), .Z(n396) );
  MUX2_X1 U438 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n452), .Z(n397) );
  MUX2_X1 U439 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(N10), .Z(n398) );
  MUX2_X1 U440 ( .A(n398), .B(n397), .S(n451), .Z(n399) );
  MUX2_X1 U441 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(N10), .Z(n400) );
  MUX2_X1 U442 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(N10), .Z(n401) );
  MUX2_X1 U443 ( .A(n401), .B(n400), .S(n451), .Z(n402) );
  MUX2_X1 U444 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n454), .Z(n403) );
  MUX2_X1 U445 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n452), .Z(n404) );
  MUX2_X1 U446 ( .A(n404), .B(n403), .S(N11), .Z(n405) );
  MUX2_X1 U447 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n453), .Z(n406) );
  MUX2_X1 U448 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n452), .Z(n407) );
  MUX2_X1 U449 ( .A(n407), .B(n406), .S(N11), .Z(n408) );
  MUX2_X1 U450 ( .A(n408), .B(n405), .S(N12), .Z(N20) );
  MUX2_X1 U451 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(N10), .Z(n409) );
  MUX2_X1 U452 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(N10), .Z(n410) );
  MUX2_X1 U453 ( .A(n410), .B(n409), .S(n451), .Z(n411) );
  MUX2_X1 U454 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(N10), .Z(n412) );
  MUX2_X1 U455 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(N10), .Z(n413) );
  MUX2_X1 U456 ( .A(n413), .B(n412), .S(n451), .Z(n414) );
  MUX2_X1 U457 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n453), .Z(n415) );
  MUX2_X1 U458 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n454), .Z(n416) );
  MUX2_X1 U459 ( .A(n416), .B(n415), .S(n451), .Z(n417) );
  MUX2_X1 U460 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n452), .Z(n418) );
  MUX2_X1 U461 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n454), .Z(n419) );
  MUX2_X1 U462 ( .A(n419), .B(n418), .S(n451), .Z(n420) );
  MUX2_X1 U463 ( .A(n420), .B(n417), .S(N12), .Z(N18) );
  MUX2_X1 U464 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n452), .Z(n421) );
  MUX2_X1 U465 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n453), .Z(n422) );
  MUX2_X1 U466 ( .A(n422), .B(n421), .S(n451), .Z(n423) );
  MUX2_X1 U467 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(N10), .Z(n424) );
  MUX2_X1 U468 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n452), .Z(n425) );
  MUX2_X1 U469 ( .A(n425), .B(n424), .S(n451), .Z(n426) );
  MUX2_X1 U470 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n454), .Z(n427) );
  MUX2_X1 U471 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n453), .Z(n428) );
  MUX2_X1 U472 ( .A(n428), .B(n427), .S(n451), .Z(n429) );
  MUX2_X1 U473 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n453), .Z(n430) );
  MUX2_X1 U474 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n452), .Z(n431) );
  MUX2_X1 U475 ( .A(n431), .B(n430), .S(n451), .Z(n432) );
  MUX2_X1 U476 ( .A(n432), .B(n429), .S(N12), .Z(N16) );
  MUX2_X1 U477 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(N10), .Z(n433) );
  MUX2_X1 U478 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n454), .Z(n434) );
  MUX2_X1 U479 ( .A(n434), .B(n433), .S(n451), .Z(n435) );
  MUX2_X1 U480 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n454), .Z(n436) );
  MUX2_X1 U481 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n452), .Z(n437) );
  MUX2_X1 U482 ( .A(n437), .B(n436), .S(n451), .Z(n438) );
  MUX2_X1 U483 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n454), .Z(n439) );
  MUX2_X1 U484 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n452), .Z(n440) );
  MUX2_X1 U485 ( .A(n440), .B(n439), .S(n451), .Z(n441) );
  MUX2_X1 U486 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n452), .Z(n442) );
  MUX2_X1 U487 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n454), .Z(n443) );
  MUX2_X1 U488 ( .A(n443), .B(n442), .S(n451), .Z(n444) );
  MUX2_X1 U489 ( .A(n444), .B(n441), .S(N12), .Z(N14) );
  MUX2_X1 U490 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n452), .Z(n445) );
  MUX2_X1 U491 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n453), .Z(n446) );
  MUX2_X1 U492 ( .A(n446), .B(n445), .S(n451), .Z(n447) );
  MUX2_X1 U493 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(N10), .Z(n448) );
  MUX2_X1 U494 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n453), .Z(n449) );
  MUX2_X1 U495 ( .A(n449), .B(n448), .S(n451), .Z(n450) );
  CLKBUF_X1 U496 ( .A(N10), .Z(n452) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE3_2 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N13, N14, N15, N18, N22, N24, N28, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[19]  ( .D(N13), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \data_out_reg[18]  ( .D(N14), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[17]  ( .D(N15), .CK(clk), .Q(data_out[17]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[10]  ( .D(N22), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[8]  ( .D(N24), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[4]  ( .D(N28), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n487), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n488), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n489), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n490), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n491), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n492), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n493), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n494), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n495), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n496), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n497), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n498), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n499), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n500), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n501), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n502), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n503), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n504), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n505), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n506), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n507), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n508), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n509), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n510), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n511), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n512), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n513), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n514), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n515), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n516), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n517), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n518), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n519), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n520), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n521), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n522), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n523), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n524), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n525), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n526), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n527), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n528), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n529), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n530), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n531), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n532), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n533), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n534), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n535), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n536), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n537), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n538), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n539), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n540), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n541), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n542), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n543), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n544), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n545), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n546), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n547), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n548), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n549), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n550), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n551), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n552), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n553), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n554), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n555), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n556), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n557), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n558), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n559), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n560), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n561), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n562), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n563), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n564), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n565), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n566), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n567), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n568), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n569), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n570), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n571), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n572), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n573), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n574), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n575), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n576), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n577), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n578), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n579), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n580), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n581), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n582), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n583), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n584), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n585), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n586), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n587), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n588), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n589), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n590), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n591), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n592), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n593), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n594), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n595), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n596), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n597), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n598), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n599), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n600), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n601), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n602), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n603), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n604), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n605), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n606), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n607), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n608), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n609), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n610), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n611), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n612), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n613), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n614), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n615), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n616), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n617), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n618), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n619), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n620), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n621), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n622), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n623), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n624), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n625), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n626), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n627), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n628), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n629), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n630), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n631), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n632), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n633), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n634), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n635), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n636), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n637), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n638), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n639), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n640), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n641), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n642), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n643), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n644), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n645), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n646), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U348 ( .A1(n464), .A2(n465), .A3(n795), .ZN(n816) );
  NAND3_X1 U349 ( .A1(n795), .A2(n465), .A3(N10), .ZN(n794) );
  NAND3_X1 U350 ( .A1(n795), .A2(n464), .A3(N11), .ZN(n773) );
  NAND3_X1 U351 ( .A1(N10), .A2(n795), .A3(N11), .ZN(n752) );
  NAND3_X1 U352 ( .A1(n464), .A2(n465), .A3(n710), .ZN(n731) );
  NAND3_X1 U353 ( .A1(N10), .A2(n465), .A3(n710), .ZN(n709) );
  NAND3_X1 U354 ( .A1(N11), .A2(n464), .A3(n710), .ZN(n688) );
  NAND3_X1 U355 ( .A1(N11), .A2(N10), .A3(n710), .ZN(n667) );
  SDFF_X1 \data_out_reg[11]  ( .D(n402), .SI(n399), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n12), .SI(n9), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n390), .SI(n387), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n378), .SI(n375), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n414), .SI(n411), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n366), .SI(n363), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n6), .SI(n3), .SE(N12), .CK(clk), .Q(
        data_out[0]) );
  SDFF_X1 \data_out_reg[2]  ( .D(n18), .SI(n15), .SE(N12), .CK(clk), .Q(
        data_out[2]) );
  SDFF_X1 \data_out_reg[16]  ( .D(n432), .SI(n429), .SE(N12), .CK(clk), .Q(
        data_out[16]) );
  SDFF_X1 \data_out_reg[6]  ( .D(n372), .SI(n369), .SE(N12), .CK(clk), .Q(
        data_out[6]) );
  SDFF_X1 \data_out_reg[12]  ( .D(n408), .SI(n405), .SE(N12), .CK(clk), .Q(
        data_out[12]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n354), .SI(n21), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n426), .SI(n423), .SE(N12), .CK(clk), .Q(
        data_out[15]) );
  BUF_X1 U3 ( .A(n794), .Z(n462) );
  BUF_X1 U4 ( .A(n773), .Z(n461) );
  BUF_X1 U5 ( .A(n731), .Z(n459) );
  BUF_X1 U6 ( .A(n709), .Z(n458) );
  BUF_X1 U7 ( .A(n688), .Z(n457) );
  BUF_X1 U8 ( .A(n452), .Z(n451) );
  BUF_X1 U9 ( .A(n816), .Z(n463) );
  BUF_X1 U10 ( .A(n752), .Z(n460) );
  BUF_X1 U11 ( .A(n667), .Z(n456) );
  BUF_X1 U12 ( .A(N10), .Z(n453) );
  BUF_X1 U13 ( .A(N10), .Z(n454) );
  BUF_X1 U14 ( .A(N10), .Z(n455) );
  BUF_X1 U15 ( .A(N11), .Z(n452) );
  AND2_X1 U16 ( .A1(N12), .A2(wr_en), .ZN(n710) );
  OAI21_X1 U17 ( .B1(n486), .B2(n462), .A(n793), .ZN(n626) );
  NAND2_X1 U18 ( .A1(\mem[1][0] ), .A2(n462), .ZN(n793) );
  OAI21_X1 U19 ( .B1(n485), .B2(n462), .A(n792), .ZN(n625) );
  NAND2_X1 U20 ( .A1(\mem[1][1] ), .A2(n462), .ZN(n792) );
  OAI21_X1 U21 ( .B1(n484), .B2(n462), .A(n791), .ZN(n624) );
  NAND2_X1 U22 ( .A1(\mem[1][2] ), .A2(n794), .ZN(n791) );
  OAI21_X1 U23 ( .B1(n483), .B2(n794), .A(n790), .ZN(n623) );
  NAND2_X1 U24 ( .A1(\mem[1][3] ), .A2(n462), .ZN(n790) );
  OAI21_X1 U25 ( .B1(n482), .B2(n794), .A(n789), .ZN(n622) );
  NAND2_X1 U26 ( .A1(\mem[1][4] ), .A2(n462), .ZN(n789) );
  OAI21_X1 U27 ( .B1(n481), .B2(n794), .A(n788), .ZN(n621) );
  NAND2_X1 U28 ( .A1(\mem[1][5] ), .A2(n794), .ZN(n788) );
  OAI21_X1 U29 ( .B1(n480), .B2(n794), .A(n787), .ZN(n620) );
  NAND2_X1 U30 ( .A1(\mem[1][6] ), .A2(n794), .ZN(n787) );
  OAI21_X1 U31 ( .B1(n479), .B2(n794), .A(n786), .ZN(n619) );
  NAND2_X1 U32 ( .A1(\mem[1][7] ), .A2(n794), .ZN(n786) );
  OAI21_X1 U33 ( .B1(n478), .B2(n794), .A(n785), .ZN(n618) );
  NAND2_X1 U34 ( .A1(\mem[1][8] ), .A2(n794), .ZN(n785) );
  OAI21_X1 U35 ( .B1(n477), .B2(n462), .A(n784), .ZN(n617) );
  NAND2_X1 U36 ( .A1(\mem[1][9] ), .A2(n794), .ZN(n784) );
  OAI21_X1 U37 ( .B1(n476), .B2(n794), .A(n783), .ZN(n616) );
  NAND2_X1 U38 ( .A1(\mem[1][10] ), .A2(n794), .ZN(n783) );
  OAI21_X1 U39 ( .B1(n475), .B2(n794), .A(n782), .ZN(n615) );
  NAND2_X1 U40 ( .A1(\mem[1][11] ), .A2(n794), .ZN(n782) );
  OAI21_X1 U41 ( .B1(n474), .B2(n462), .A(n781), .ZN(n614) );
  NAND2_X1 U42 ( .A1(\mem[1][12] ), .A2(n462), .ZN(n781) );
  OAI21_X1 U43 ( .B1(n473), .B2(n462), .A(n780), .ZN(n613) );
  NAND2_X1 U44 ( .A1(\mem[1][13] ), .A2(n462), .ZN(n780) );
  OAI21_X1 U45 ( .B1(n472), .B2(n462), .A(n779), .ZN(n612) );
  NAND2_X1 U46 ( .A1(\mem[1][14] ), .A2(n462), .ZN(n779) );
  OAI21_X1 U47 ( .B1(n471), .B2(n794), .A(n778), .ZN(n611) );
  NAND2_X1 U48 ( .A1(\mem[1][15] ), .A2(n462), .ZN(n778) );
  OAI21_X1 U49 ( .B1(n470), .B2(n794), .A(n777), .ZN(n610) );
  NAND2_X1 U50 ( .A1(\mem[1][16] ), .A2(n462), .ZN(n777) );
  OAI21_X1 U51 ( .B1(n469), .B2(n794), .A(n776), .ZN(n609) );
  NAND2_X1 U52 ( .A1(\mem[1][17] ), .A2(n462), .ZN(n776) );
  OAI21_X1 U53 ( .B1(n468), .B2(n462), .A(n775), .ZN(n608) );
  NAND2_X1 U54 ( .A1(\mem[1][18] ), .A2(n462), .ZN(n775) );
  OAI21_X1 U55 ( .B1(n467), .B2(n462), .A(n774), .ZN(n607) );
  NAND2_X1 U56 ( .A1(\mem[1][19] ), .A2(n462), .ZN(n774) );
  OAI21_X1 U57 ( .B1(n486), .B2(n461), .A(n772), .ZN(n606) );
  NAND2_X1 U58 ( .A1(\mem[2][0] ), .A2(n461), .ZN(n772) );
  OAI21_X1 U59 ( .B1(n485), .B2(n461), .A(n771), .ZN(n605) );
  NAND2_X1 U60 ( .A1(\mem[2][1] ), .A2(n461), .ZN(n771) );
  OAI21_X1 U61 ( .B1(n484), .B2(n461), .A(n770), .ZN(n604) );
  NAND2_X1 U62 ( .A1(\mem[2][2] ), .A2(n773), .ZN(n770) );
  OAI21_X1 U63 ( .B1(n483), .B2(n773), .A(n769), .ZN(n603) );
  NAND2_X1 U64 ( .A1(\mem[2][3] ), .A2(n461), .ZN(n769) );
  OAI21_X1 U65 ( .B1(n482), .B2(n773), .A(n768), .ZN(n602) );
  NAND2_X1 U66 ( .A1(\mem[2][4] ), .A2(n461), .ZN(n768) );
  OAI21_X1 U67 ( .B1(n481), .B2(n773), .A(n767), .ZN(n601) );
  NAND2_X1 U68 ( .A1(\mem[2][5] ), .A2(n773), .ZN(n767) );
  OAI21_X1 U69 ( .B1(n480), .B2(n773), .A(n766), .ZN(n600) );
  NAND2_X1 U70 ( .A1(\mem[2][6] ), .A2(n773), .ZN(n766) );
  OAI21_X1 U71 ( .B1(n479), .B2(n773), .A(n765), .ZN(n599) );
  NAND2_X1 U72 ( .A1(\mem[2][7] ), .A2(n773), .ZN(n765) );
  OAI21_X1 U73 ( .B1(n478), .B2(n773), .A(n764), .ZN(n598) );
  NAND2_X1 U74 ( .A1(\mem[2][8] ), .A2(n773), .ZN(n764) );
  OAI21_X1 U75 ( .B1(n477), .B2(n461), .A(n763), .ZN(n597) );
  NAND2_X1 U76 ( .A1(\mem[2][9] ), .A2(n773), .ZN(n763) );
  OAI21_X1 U77 ( .B1(n476), .B2(n773), .A(n762), .ZN(n596) );
  NAND2_X1 U78 ( .A1(\mem[2][10] ), .A2(n773), .ZN(n762) );
  OAI21_X1 U79 ( .B1(n475), .B2(n773), .A(n761), .ZN(n595) );
  NAND2_X1 U80 ( .A1(\mem[2][11] ), .A2(n773), .ZN(n761) );
  OAI21_X1 U81 ( .B1(n474), .B2(n461), .A(n760), .ZN(n594) );
  NAND2_X1 U82 ( .A1(\mem[2][12] ), .A2(n461), .ZN(n760) );
  OAI21_X1 U83 ( .B1(n473), .B2(n461), .A(n759), .ZN(n593) );
  NAND2_X1 U84 ( .A1(\mem[2][13] ), .A2(n461), .ZN(n759) );
  OAI21_X1 U85 ( .B1(n472), .B2(n461), .A(n758), .ZN(n592) );
  NAND2_X1 U86 ( .A1(\mem[2][14] ), .A2(n461), .ZN(n758) );
  OAI21_X1 U87 ( .B1(n471), .B2(n773), .A(n757), .ZN(n591) );
  NAND2_X1 U88 ( .A1(\mem[2][15] ), .A2(n461), .ZN(n757) );
  OAI21_X1 U89 ( .B1(n470), .B2(n773), .A(n756), .ZN(n590) );
  NAND2_X1 U90 ( .A1(\mem[2][16] ), .A2(n461), .ZN(n756) );
  OAI21_X1 U91 ( .B1(n469), .B2(n773), .A(n755), .ZN(n589) );
  NAND2_X1 U92 ( .A1(\mem[2][17] ), .A2(n461), .ZN(n755) );
  OAI21_X1 U93 ( .B1(n468), .B2(n461), .A(n754), .ZN(n588) );
  NAND2_X1 U94 ( .A1(\mem[2][18] ), .A2(n461), .ZN(n754) );
  OAI21_X1 U95 ( .B1(n467), .B2(n461), .A(n753), .ZN(n587) );
  NAND2_X1 U96 ( .A1(\mem[2][19] ), .A2(n461), .ZN(n753) );
  OAI21_X1 U97 ( .B1(n486), .B2(n752), .A(n751), .ZN(n586) );
  NAND2_X1 U98 ( .A1(\mem[3][0] ), .A2(n460), .ZN(n751) );
  OAI21_X1 U99 ( .B1(n485), .B2(n752), .A(n750), .ZN(n585) );
  NAND2_X1 U100 ( .A1(\mem[3][1] ), .A2(n460), .ZN(n750) );
  OAI21_X1 U101 ( .B1(n484), .B2(n752), .A(n749), .ZN(n584) );
  NAND2_X1 U102 ( .A1(\mem[3][2] ), .A2(n460), .ZN(n749) );
  OAI21_X1 U103 ( .B1(n483), .B2(n752), .A(n748), .ZN(n583) );
  NAND2_X1 U104 ( .A1(\mem[3][3] ), .A2(n460), .ZN(n748) );
  OAI21_X1 U105 ( .B1(n482), .B2(n460), .A(n747), .ZN(n582) );
  NAND2_X1 U106 ( .A1(\mem[3][4] ), .A2(n460), .ZN(n747) );
  OAI21_X1 U107 ( .B1(n481), .B2(n460), .A(n746), .ZN(n581) );
  NAND2_X1 U108 ( .A1(\mem[3][5] ), .A2(n460), .ZN(n746) );
  OAI21_X1 U109 ( .B1(n480), .B2(n752), .A(n745), .ZN(n580) );
  NAND2_X1 U110 ( .A1(\mem[3][6] ), .A2(n460), .ZN(n745) );
  OAI21_X1 U111 ( .B1(n479), .B2(n752), .A(n744), .ZN(n579) );
  NAND2_X1 U112 ( .A1(\mem[3][7] ), .A2(n460), .ZN(n744) );
  OAI21_X1 U113 ( .B1(n478), .B2(n752), .A(n743), .ZN(n578) );
  NAND2_X1 U114 ( .A1(\mem[3][8] ), .A2(n460), .ZN(n743) );
  OAI21_X1 U115 ( .B1(n477), .B2(n752), .A(n742), .ZN(n577) );
  NAND2_X1 U116 ( .A1(\mem[3][9] ), .A2(n460), .ZN(n742) );
  OAI21_X1 U117 ( .B1(n476), .B2(n752), .A(n741), .ZN(n576) );
  NAND2_X1 U118 ( .A1(\mem[3][10] ), .A2(n460), .ZN(n741) );
  OAI21_X1 U119 ( .B1(n475), .B2(n752), .A(n740), .ZN(n575) );
  NAND2_X1 U120 ( .A1(\mem[3][11] ), .A2(n460), .ZN(n740) );
  OAI21_X1 U121 ( .B1(n474), .B2(n752), .A(n739), .ZN(n574) );
  NAND2_X1 U122 ( .A1(\mem[3][12] ), .A2(n752), .ZN(n739) );
  OAI21_X1 U123 ( .B1(n473), .B2(n752), .A(n738), .ZN(n573) );
  NAND2_X1 U124 ( .A1(\mem[3][13] ), .A2(n752), .ZN(n738) );
  OAI21_X1 U125 ( .B1(n472), .B2(n752), .A(n737), .ZN(n572) );
  NAND2_X1 U126 ( .A1(\mem[3][14] ), .A2(n752), .ZN(n737) );
  OAI21_X1 U127 ( .B1(n471), .B2(n752), .A(n736), .ZN(n571) );
  NAND2_X1 U128 ( .A1(\mem[3][15] ), .A2(n460), .ZN(n736) );
  OAI21_X1 U129 ( .B1(n470), .B2(n752), .A(n735), .ZN(n570) );
  NAND2_X1 U130 ( .A1(\mem[3][16] ), .A2(n752), .ZN(n735) );
  OAI21_X1 U131 ( .B1(n469), .B2(n752), .A(n734), .ZN(n569) );
  NAND2_X1 U132 ( .A1(\mem[3][17] ), .A2(n752), .ZN(n734) );
  OAI21_X1 U133 ( .B1(n468), .B2(n752), .A(n733), .ZN(n568) );
  NAND2_X1 U134 ( .A1(\mem[3][18] ), .A2(n752), .ZN(n733) );
  OAI21_X1 U135 ( .B1(n467), .B2(n752), .A(n732), .ZN(n567) );
  NAND2_X1 U136 ( .A1(\mem[3][19] ), .A2(n460), .ZN(n732) );
  OAI21_X1 U137 ( .B1(n486), .B2(n731), .A(n730), .ZN(n566) );
  NAND2_X1 U138 ( .A1(\mem[4][0] ), .A2(n731), .ZN(n730) );
  OAI21_X1 U139 ( .B1(n485), .B2(n459), .A(n729), .ZN(n565) );
  NAND2_X1 U140 ( .A1(\mem[4][1] ), .A2(n731), .ZN(n729) );
  OAI21_X1 U141 ( .B1(n484), .B2(n459), .A(n728), .ZN(n564) );
  NAND2_X1 U142 ( .A1(\mem[4][2] ), .A2(n731), .ZN(n728) );
  OAI21_X1 U143 ( .B1(n483), .B2(n459), .A(n727), .ZN(n563) );
  NAND2_X1 U144 ( .A1(\mem[4][3] ), .A2(n731), .ZN(n727) );
  OAI21_X1 U145 ( .B1(n482), .B2(n459), .A(n726), .ZN(n562) );
  NAND2_X1 U146 ( .A1(\mem[4][4] ), .A2(n731), .ZN(n726) );
  OAI21_X1 U147 ( .B1(n481), .B2(n459), .A(n725), .ZN(n561) );
  NAND2_X1 U148 ( .A1(\mem[4][5] ), .A2(n731), .ZN(n725) );
  OAI21_X1 U149 ( .B1(n480), .B2(n459), .A(n724), .ZN(n560) );
  NAND2_X1 U150 ( .A1(\mem[4][6] ), .A2(n731), .ZN(n724) );
  OAI21_X1 U151 ( .B1(n479), .B2(n459), .A(n723), .ZN(n559) );
  NAND2_X1 U152 ( .A1(\mem[4][7] ), .A2(n731), .ZN(n723) );
  OAI21_X1 U153 ( .B1(n478), .B2(n459), .A(n722), .ZN(n558) );
  NAND2_X1 U154 ( .A1(\mem[4][8] ), .A2(n731), .ZN(n722) );
  OAI21_X1 U155 ( .B1(n477), .B2(n731), .A(n721), .ZN(n557) );
  NAND2_X1 U156 ( .A1(\mem[4][9] ), .A2(n731), .ZN(n721) );
  OAI21_X1 U157 ( .B1(n476), .B2(n459), .A(n720), .ZN(n556) );
  NAND2_X1 U158 ( .A1(\mem[4][10] ), .A2(n731), .ZN(n720) );
  OAI21_X1 U159 ( .B1(n475), .B2(n459), .A(n719), .ZN(n555) );
  NAND2_X1 U160 ( .A1(\mem[4][11] ), .A2(n731), .ZN(n719) );
  OAI21_X1 U161 ( .B1(n474), .B2(n731), .A(n718), .ZN(n554) );
  NAND2_X1 U162 ( .A1(\mem[4][12] ), .A2(n731), .ZN(n718) );
  OAI21_X1 U163 ( .B1(n473), .B2(n459), .A(n717), .ZN(n553) );
  NAND2_X1 U164 ( .A1(\mem[4][13] ), .A2(n731), .ZN(n717) );
  OAI21_X1 U165 ( .B1(n472), .B2(n731), .A(n716), .ZN(n552) );
  NAND2_X1 U166 ( .A1(\mem[4][14] ), .A2(n731), .ZN(n716) );
  OAI21_X1 U167 ( .B1(n471), .B2(n459), .A(n715), .ZN(n551) );
  NAND2_X1 U168 ( .A1(\mem[4][15] ), .A2(n731), .ZN(n715) );
  OAI21_X1 U169 ( .B1(n470), .B2(n459), .A(n714), .ZN(n550) );
  NAND2_X1 U170 ( .A1(\mem[4][16] ), .A2(n731), .ZN(n714) );
  OAI21_X1 U171 ( .B1(n469), .B2(n459), .A(n713), .ZN(n549) );
  NAND2_X1 U172 ( .A1(\mem[4][17] ), .A2(n731), .ZN(n713) );
  OAI21_X1 U173 ( .B1(n468), .B2(n459), .A(n712), .ZN(n548) );
  NAND2_X1 U174 ( .A1(\mem[4][18] ), .A2(n731), .ZN(n712) );
  OAI21_X1 U175 ( .B1(n467), .B2(n459), .A(n711), .ZN(n547) );
  NAND2_X1 U176 ( .A1(\mem[4][19] ), .A2(n731), .ZN(n711) );
  OAI21_X1 U177 ( .B1(n486), .B2(n709), .A(n708), .ZN(n546) );
  NAND2_X1 U178 ( .A1(\mem[5][0] ), .A2(n709), .ZN(n708) );
  OAI21_X1 U179 ( .B1(n485), .B2(n458), .A(n707), .ZN(n545) );
  NAND2_X1 U180 ( .A1(\mem[5][1] ), .A2(n709), .ZN(n707) );
  OAI21_X1 U181 ( .B1(n484), .B2(n458), .A(n706), .ZN(n544) );
  NAND2_X1 U182 ( .A1(\mem[5][2] ), .A2(n709), .ZN(n706) );
  OAI21_X1 U183 ( .B1(n483), .B2(n458), .A(n705), .ZN(n543) );
  NAND2_X1 U184 ( .A1(\mem[5][3] ), .A2(n709), .ZN(n705) );
  OAI21_X1 U185 ( .B1(n482), .B2(n458), .A(n704), .ZN(n542) );
  NAND2_X1 U186 ( .A1(\mem[5][4] ), .A2(n709), .ZN(n704) );
  OAI21_X1 U187 ( .B1(n481), .B2(n458), .A(n703), .ZN(n541) );
  NAND2_X1 U188 ( .A1(\mem[5][5] ), .A2(n709), .ZN(n703) );
  OAI21_X1 U189 ( .B1(n480), .B2(n458), .A(n702), .ZN(n540) );
  NAND2_X1 U190 ( .A1(\mem[5][6] ), .A2(n709), .ZN(n702) );
  OAI21_X1 U191 ( .B1(n479), .B2(n458), .A(n701), .ZN(n539) );
  NAND2_X1 U192 ( .A1(\mem[5][7] ), .A2(n709), .ZN(n701) );
  OAI21_X1 U193 ( .B1(n478), .B2(n458), .A(n700), .ZN(n538) );
  NAND2_X1 U194 ( .A1(\mem[5][8] ), .A2(n709), .ZN(n700) );
  OAI21_X1 U195 ( .B1(n477), .B2(n709), .A(n699), .ZN(n537) );
  NAND2_X1 U196 ( .A1(\mem[5][9] ), .A2(n709), .ZN(n699) );
  OAI21_X1 U197 ( .B1(n476), .B2(n458), .A(n698), .ZN(n536) );
  NAND2_X1 U198 ( .A1(\mem[5][10] ), .A2(n709), .ZN(n698) );
  OAI21_X1 U199 ( .B1(n475), .B2(n458), .A(n697), .ZN(n535) );
  NAND2_X1 U200 ( .A1(\mem[5][11] ), .A2(n709), .ZN(n697) );
  OAI21_X1 U201 ( .B1(n474), .B2(n709), .A(n696), .ZN(n534) );
  NAND2_X1 U202 ( .A1(\mem[5][12] ), .A2(n709), .ZN(n696) );
  OAI21_X1 U203 ( .B1(n473), .B2(n458), .A(n695), .ZN(n533) );
  NAND2_X1 U204 ( .A1(\mem[5][13] ), .A2(n709), .ZN(n695) );
  OAI21_X1 U205 ( .B1(n472), .B2(n709), .A(n694), .ZN(n532) );
  NAND2_X1 U206 ( .A1(\mem[5][14] ), .A2(n709), .ZN(n694) );
  OAI21_X1 U207 ( .B1(n471), .B2(n458), .A(n693), .ZN(n531) );
  NAND2_X1 U208 ( .A1(\mem[5][15] ), .A2(n709), .ZN(n693) );
  OAI21_X1 U209 ( .B1(n470), .B2(n458), .A(n692), .ZN(n530) );
  NAND2_X1 U210 ( .A1(\mem[5][16] ), .A2(n709), .ZN(n692) );
  OAI21_X1 U211 ( .B1(n469), .B2(n458), .A(n691), .ZN(n529) );
  NAND2_X1 U212 ( .A1(\mem[5][17] ), .A2(n709), .ZN(n691) );
  OAI21_X1 U213 ( .B1(n468), .B2(n458), .A(n690), .ZN(n528) );
  NAND2_X1 U214 ( .A1(\mem[5][18] ), .A2(n709), .ZN(n690) );
  OAI21_X1 U215 ( .B1(n467), .B2(n458), .A(n689), .ZN(n527) );
  NAND2_X1 U216 ( .A1(\mem[5][19] ), .A2(n709), .ZN(n689) );
  OAI21_X1 U217 ( .B1(n486), .B2(n688), .A(n687), .ZN(n526) );
  NAND2_X1 U218 ( .A1(\mem[6][0] ), .A2(n688), .ZN(n687) );
  OAI21_X1 U219 ( .B1(n485), .B2(n457), .A(n686), .ZN(n525) );
  NAND2_X1 U220 ( .A1(\mem[6][1] ), .A2(n688), .ZN(n686) );
  OAI21_X1 U221 ( .B1(n484), .B2(n457), .A(n685), .ZN(n524) );
  NAND2_X1 U222 ( .A1(\mem[6][2] ), .A2(n688), .ZN(n685) );
  OAI21_X1 U223 ( .B1(n483), .B2(n457), .A(n684), .ZN(n523) );
  NAND2_X1 U224 ( .A1(\mem[6][3] ), .A2(n688), .ZN(n684) );
  OAI21_X1 U225 ( .B1(n482), .B2(n457), .A(n683), .ZN(n522) );
  NAND2_X1 U226 ( .A1(\mem[6][4] ), .A2(n688), .ZN(n683) );
  OAI21_X1 U227 ( .B1(n481), .B2(n457), .A(n682), .ZN(n521) );
  NAND2_X1 U228 ( .A1(\mem[6][5] ), .A2(n688), .ZN(n682) );
  OAI21_X1 U229 ( .B1(n480), .B2(n457), .A(n681), .ZN(n520) );
  NAND2_X1 U230 ( .A1(\mem[6][6] ), .A2(n688), .ZN(n681) );
  OAI21_X1 U231 ( .B1(n479), .B2(n457), .A(n680), .ZN(n519) );
  NAND2_X1 U232 ( .A1(\mem[6][7] ), .A2(n688), .ZN(n680) );
  OAI21_X1 U233 ( .B1(n478), .B2(n457), .A(n679), .ZN(n518) );
  NAND2_X1 U234 ( .A1(\mem[6][8] ), .A2(n688), .ZN(n679) );
  OAI21_X1 U235 ( .B1(n477), .B2(n688), .A(n678), .ZN(n517) );
  NAND2_X1 U236 ( .A1(\mem[6][9] ), .A2(n688), .ZN(n678) );
  OAI21_X1 U237 ( .B1(n476), .B2(n457), .A(n677), .ZN(n516) );
  NAND2_X1 U238 ( .A1(\mem[6][10] ), .A2(n688), .ZN(n677) );
  OAI21_X1 U239 ( .B1(n475), .B2(n457), .A(n676), .ZN(n515) );
  NAND2_X1 U240 ( .A1(\mem[6][11] ), .A2(n688), .ZN(n676) );
  OAI21_X1 U241 ( .B1(n474), .B2(n688), .A(n675), .ZN(n514) );
  NAND2_X1 U242 ( .A1(\mem[6][12] ), .A2(n688), .ZN(n675) );
  OAI21_X1 U243 ( .B1(n473), .B2(n457), .A(n674), .ZN(n513) );
  NAND2_X1 U244 ( .A1(\mem[6][13] ), .A2(n688), .ZN(n674) );
  OAI21_X1 U245 ( .B1(n472), .B2(n688), .A(n673), .ZN(n512) );
  NAND2_X1 U246 ( .A1(\mem[6][14] ), .A2(n688), .ZN(n673) );
  OAI21_X1 U247 ( .B1(n471), .B2(n457), .A(n672), .ZN(n511) );
  NAND2_X1 U248 ( .A1(\mem[6][15] ), .A2(n688), .ZN(n672) );
  OAI21_X1 U249 ( .B1(n470), .B2(n457), .A(n671), .ZN(n510) );
  NAND2_X1 U250 ( .A1(\mem[6][16] ), .A2(n688), .ZN(n671) );
  OAI21_X1 U251 ( .B1(n469), .B2(n457), .A(n670), .ZN(n509) );
  NAND2_X1 U252 ( .A1(\mem[6][17] ), .A2(n688), .ZN(n670) );
  OAI21_X1 U253 ( .B1(n468), .B2(n457), .A(n669), .ZN(n508) );
  NAND2_X1 U254 ( .A1(\mem[6][18] ), .A2(n688), .ZN(n669) );
  OAI21_X1 U255 ( .B1(n467), .B2(n457), .A(n668), .ZN(n507) );
  NAND2_X1 U256 ( .A1(\mem[6][19] ), .A2(n688), .ZN(n668) );
  OAI21_X1 U257 ( .B1(n486), .B2(n667), .A(n666), .ZN(n506) );
  NAND2_X1 U258 ( .A1(\mem[7][0] ), .A2(n456), .ZN(n666) );
  OAI21_X1 U259 ( .B1(n485), .B2(n667), .A(n665), .ZN(n505) );
  NAND2_X1 U260 ( .A1(\mem[7][1] ), .A2(n456), .ZN(n665) );
  OAI21_X1 U261 ( .B1(n484), .B2(n667), .A(n664), .ZN(n504) );
  NAND2_X1 U262 ( .A1(\mem[7][2] ), .A2(n456), .ZN(n664) );
  OAI21_X1 U263 ( .B1(n483), .B2(n667), .A(n663), .ZN(n503) );
  NAND2_X1 U264 ( .A1(\mem[7][3] ), .A2(n456), .ZN(n663) );
  OAI21_X1 U265 ( .B1(n482), .B2(n456), .A(n662), .ZN(n502) );
  NAND2_X1 U266 ( .A1(\mem[7][4] ), .A2(n456), .ZN(n662) );
  OAI21_X1 U267 ( .B1(n481), .B2(n667), .A(n661), .ZN(n501) );
  NAND2_X1 U268 ( .A1(\mem[7][5] ), .A2(n456), .ZN(n661) );
  OAI21_X1 U269 ( .B1(n480), .B2(n667), .A(n660), .ZN(n500) );
  NAND2_X1 U270 ( .A1(\mem[7][6] ), .A2(n456), .ZN(n660) );
  OAI21_X1 U271 ( .B1(n479), .B2(n667), .A(n659), .ZN(n499) );
  NAND2_X1 U272 ( .A1(\mem[7][7] ), .A2(n456), .ZN(n659) );
  OAI21_X1 U273 ( .B1(n478), .B2(n667), .A(n658), .ZN(n498) );
  NAND2_X1 U274 ( .A1(\mem[7][8] ), .A2(n456), .ZN(n658) );
  OAI21_X1 U275 ( .B1(n477), .B2(n667), .A(n657), .ZN(n497) );
  NAND2_X1 U276 ( .A1(\mem[7][9] ), .A2(n456), .ZN(n657) );
  OAI21_X1 U277 ( .B1(n476), .B2(n667), .A(n656), .ZN(n496) );
  NAND2_X1 U278 ( .A1(\mem[7][10] ), .A2(n456), .ZN(n656) );
  OAI21_X1 U279 ( .B1(n475), .B2(n667), .A(n655), .ZN(n495) );
  NAND2_X1 U280 ( .A1(\mem[7][11] ), .A2(n456), .ZN(n655) );
  OAI21_X1 U281 ( .B1(n474), .B2(n667), .A(n654), .ZN(n494) );
  NAND2_X1 U282 ( .A1(\mem[7][12] ), .A2(n667), .ZN(n654) );
  OAI21_X1 U283 ( .B1(n473), .B2(n456), .A(n653), .ZN(n493) );
  NAND2_X1 U284 ( .A1(\mem[7][13] ), .A2(n667), .ZN(n653) );
  OAI21_X1 U285 ( .B1(n472), .B2(n456), .A(n652), .ZN(n492) );
  NAND2_X1 U286 ( .A1(\mem[7][14] ), .A2(n667), .ZN(n652) );
  OAI21_X1 U287 ( .B1(n471), .B2(n667), .A(n651), .ZN(n491) );
  NAND2_X1 U288 ( .A1(\mem[7][15] ), .A2(n667), .ZN(n651) );
  OAI21_X1 U289 ( .B1(n470), .B2(n667), .A(n650), .ZN(n490) );
  NAND2_X1 U290 ( .A1(\mem[7][16] ), .A2(n667), .ZN(n650) );
  OAI21_X1 U291 ( .B1(n469), .B2(n667), .A(n649), .ZN(n489) );
  NAND2_X1 U292 ( .A1(\mem[7][17] ), .A2(n667), .ZN(n649) );
  OAI21_X1 U293 ( .B1(n468), .B2(n667), .A(n648), .ZN(n488) );
  NAND2_X1 U294 ( .A1(\mem[7][18] ), .A2(n667), .ZN(n648) );
  OAI21_X1 U295 ( .B1(n467), .B2(n667), .A(n647), .ZN(n487) );
  NAND2_X1 U296 ( .A1(\mem[7][19] ), .A2(n456), .ZN(n647) );
  OAI21_X1 U297 ( .B1(n816), .B2(n484), .A(n813), .ZN(n644) );
  NAND2_X1 U298 ( .A1(\mem[0][2] ), .A2(n463), .ZN(n813) );
  OAI21_X1 U299 ( .B1(n816), .B2(n483), .A(n812), .ZN(n643) );
  NAND2_X1 U300 ( .A1(\mem[0][3] ), .A2(n463), .ZN(n812) );
  OAI21_X1 U301 ( .B1(n816), .B2(n482), .A(n811), .ZN(n642) );
  NAND2_X1 U302 ( .A1(\mem[0][4] ), .A2(n463), .ZN(n811) );
  OAI21_X1 U303 ( .B1(n816), .B2(n481), .A(n810), .ZN(n641) );
  NAND2_X1 U304 ( .A1(\mem[0][5] ), .A2(n463), .ZN(n810) );
  OAI21_X1 U305 ( .B1(n816), .B2(n480), .A(n809), .ZN(n640) );
  NAND2_X1 U306 ( .A1(\mem[0][6] ), .A2(n463), .ZN(n809) );
  OAI21_X1 U307 ( .B1(n816), .B2(n479), .A(n808), .ZN(n639) );
  NAND2_X1 U308 ( .A1(\mem[0][7] ), .A2(n463), .ZN(n808) );
  OAI21_X1 U309 ( .B1(n816), .B2(n478), .A(n807), .ZN(n638) );
  NAND2_X1 U310 ( .A1(\mem[0][8] ), .A2(n463), .ZN(n807) );
  OAI21_X1 U311 ( .B1(n816), .B2(n477), .A(n806), .ZN(n637) );
  NAND2_X1 U312 ( .A1(\mem[0][9] ), .A2(n463), .ZN(n806) );
  OAI21_X1 U313 ( .B1(n816), .B2(n476), .A(n805), .ZN(n636) );
  NAND2_X1 U314 ( .A1(\mem[0][10] ), .A2(n463), .ZN(n805) );
  OAI21_X1 U315 ( .B1(n816), .B2(n475), .A(n804), .ZN(n635) );
  NAND2_X1 U316 ( .A1(\mem[0][11] ), .A2(n463), .ZN(n804) );
  OAI21_X1 U317 ( .B1(n816), .B2(n474), .A(n803), .ZN(n634) );
  NAND2_X1 U318 ( .A1(\mem[0][12] ), .A2(n816), .ZN(n803) );
  OAI21_X1 U319 ( .B1(n816), .B2(n473), .A(n802), .ZN(n633) );
  NAND2_X1 U320 ( .A1(\mem[0][13] ), .A2(n816), .ZN(n802) );
  OAI21_X1 U321 ( .B1(n463), .B2(n472), .A(n801), .ZN(n632) );
  NAND2_X1 U322 ( .A1(\mem[0][14] ), .A2(n816), .ZN(n801) );
  OAI21_X1 U323 ( .B1(n816), .B2(n471), .A(n800), .ZN(n631) );
  NAND2_X1 U324 ( .A1(\mem[0][15] ), .A2(n463), .ZN(n800) );
  OAI21_X1 U325 ( .B1(n816), .B2(n470), .A(n799), .ZN(n630) );
  NAND2_X1 U326 ( .A1(\mem[0][16] ), .A2(n816), .ZN(n799) );
  OAI21_X1 U327 ( .B1(n816), .B2(n469), .A(n798), .ZN(n629) );
  NAND2_X1 U328 ( .A1(\mem[0][17] ), .A2(n816), .ZN(n798) );
  OAI21_X1 U329 ( .B1(n816), .B2(n468), .A(n797), .ZN(n628) );
  NAND2_X1 U330 ( .A1(\mem[0][18] ), .A2(n816), .ZN(n797) );
  OAI21_X1 U331 ( .B1(n463), .B2(n486), .A(n815), .ZN(n646) );
  NAND2_X1 U332 ( .A1(\mem[0][0] ), .A2(n463), .ZN(n815) );
  OAI21_X1 U333 ( .B1(n816), .B2(n485), .A(n814), .ZN(n645) );
  NAND2_X1 U334 ( .A1(\mem[0][1] ), .A2(n463), .ZN(n814) );
  OAI21_X1 U335 ( .B1(n816), .B2(n467), .A(n796), .ZN(n627) );
  NAND2_X1 U336 ( .A1(\mem[0][19] ), .A2(n463), .ZN(n796) );
  NOR2_X1 U337 ( .A1(n466), .A2(N12), .ZN(n795) );
  INV_X1 U338 ( .A(wr_en), .ZN(n466) );
  INV_X1 U339 ( .A(N10), .ZN(n464) );
  INV_X1 U340 ( .A(N11), .ZN(n465) );
  INV_X1 U341 ( .A(data_in[0]), .ZN(n486) );
  INV_X1 U342 ( .A(data_in[1]), .ZN(n485) );
  INV_X1 U343 ( .A(data_in[2]), .ZN(n484) );
  INV_X1 U344 ( .A(data_in[3]), .ZN(n483) );
  INV_X1 U345 ( .A(data_in[4]), .ZN(n482) );
  INV_X1 U346 ( .A(data_in[5]), .ZN(n481) );
  INV_X1 U347 ( .A(data_in[6]), .ZN(n480) );
  INV_X1 U356 ( .A(data_in[7]), .ZN(n479) );
  INV_X1 U357 ( .A(data_in[8]), .ZN(n478) );
  INV_X1 U358 ( .A(data_in[9]), .ZN(n477) );
  INV_X1 U359 ( .A(data_in[10]), .ZN(n476) );
  INV_X1 U360 ( .A(data_in[11]), .ZN(n475) );
  INV_X1 U361 ( .A(data_in[12]), .ZN(n474) );
  INV_X1 U362 ( .A(data_in[13]), .ZN(n473) );
  INV_X1 U363 ( .A(data_in[14]), .ZN(n472) );
  INV_X1 U364 ( .A(data_in[15]), .ZN(n471) );
  INV_X1 U365 ( .A(data_in[16]), .ZN(n470) );
  INV_X1 U366 ( .A(data_in[17]), .ZN(n469) );
  INV_X1 U367 ( .A(data_in[18]), .ZN(n468) );
  INV_X1 U368 ( .A(data_in[19]), .ZN(n467) );
  MUX2_X1 U369 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n455), .Z(n1) );
  MUX2_X1 U370 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n453), .Z(n2) );
  MUX2_X1 U371 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U372 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n454), .Z(n4) );
  MUX2_X1 U373 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n455), .Z(n5) );
  MUX2_X1 U374 ( .A(n5), .B(n4), .S(N11), .Z(n6) );
  MUX2_X1 U375 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n454), .Z(n7) );
  MUX2_X1 U376 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n455), .Z(n8) );
  MUX2_X1 U377 ( .A(n8), .B(n7), .S(N11), .Z(n9) );
  MUX2_X1 U378 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(N10), .Z(n10) );
  MUX2_X1 U379 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n454), .Z(n11) );
  MUX2_X1 U380 ( .A(n11), .B(n10), .S(n452), .Z(n12) );
  MUX2_X1 U381 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(N10), .Z(n13) );
  MUX2_X1 U382 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(N10), .Z(n14) );
  MUX2_X1 U383 ( .A(n14), .B(n13), .S(N11), .Z(n15) );
  MUX2_X1 U384 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(N10), .Z(n16) );
  MUX2_X1 U385 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(N10), .Z(n17) );
  MUX2_X1 U386 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U387 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(N10), .Z(n19) );
  MUX2_X1 U388 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n20) );
  MUX2_X1 U389 ( .A(n20), .B(n19), .S(N11), .Z(n21) );
  MUX2_X1 U390 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n22) );
  MUX2_X1 U391 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n23) );
  MUX2_X1 U392 ( .A(n23), .B(n22), .S(N11), .Z(n354) );
  MUX2_X1 U393 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n453), .Z(n355) );
  MUX2_X1 U394 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n454), .Z(n356) );
  MUX2_X1 U395 ( .A(n356), .B(n355), .S(N11), .Z(n357) );
  MUX2_X1 U396 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n455), .Z(n358) );
  MUX2_X1 U397 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n454), .Z(n359) );
  MUX2_X1 U398 ( .A(n359), .B(n358), .S(n452), .Z(n360) );
  MUX2_X1 U399 ( .A(n360), .B(n357), .S(N12), .Z(N28) );
  MUX2_X1 U400 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n455), .Z(n361) );
  MUX2_X1 U401 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n453), .Z(n362) );
  MUX2_X1 U402 ( .A(n362), .B(n361), .S(N11), .Z(n363) );
  MUX2_X1 U403 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n364) );
  MUX2_X1 U404 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n454), .Z(n365) );
  MUX2_X1 U405 ( .A(n365), .B(n364), .S(N11), .Z(n366) );
  MUX2_X1 U406 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n455), .Z(n367) );
  MUX2_X1 U407 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n455), .Z(n368) );
  MUX2_X1 U408 ( .A(n368), .B(n367), .S(N11), .Z(n369) );
  MUX2_X1 U409 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n453), .Z(n370) );
  MUX2_X1 U410 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n453), .Z(n371) );
  MUX2_X1 U411 ( .A(n371), .B(n370), .S(N11), .Z(n372) );
  MUX2_X1 U412 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n454), .Z(n373) );
  MUX2_X1 U413 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n454), .Z(n374) );
  MUX2_X1 U414 ( .A(n374), .B(n373), .S(N11), .Z(n375) );
  MUX2_X1 U415 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n455), .Z(n376) );
  MUX2_X1 U416 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n377) );
  MUX2_X1 U417 ( .A(n377), .B(n376), .S(N11), .Z(n378) );
  MUX2_X1 U418 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n455), .Z(n379) );
  MUX2_X1 U419 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n455), .Z(n380) );
  MUX2_X1 U420 ( .A(n380), .B(n379), .S(n451), .Z(n381) );
  MUX2_X1 U421 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n453), .Z(n382) );
  MUX2_X1 U422 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n455), .Z(n383) );
  MUX2_X1 U423 ( .A(n383), .B(n382), .S(n451), .Z(n384) );
  MUX2_X1 U424 ( .A(n384), .B(n381), .S(N12), .Z(N24) );
  MUX2_X1 U425 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n453), .Z(n385) );
  MUX2_X1 U426 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n453), .Z(n386) );
  MUX2_X1 U427 ( .A(n386), .B(n385), .S(n451), .Z(n387) );
  MUX2_X1 U428 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n453), .Z(n388) );
  MUX2_X1 U429 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n454), .Z(n389) );
  MUX2_X1 U430 ( .A(n389), .B(n388), .S(n451), .Z(n390) );
  MUX2_X1 U431 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n454), .Z(n391) );
  MUX2_X1 U432 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n453), .Z(n392) );
  MUX2_X1 U433 ( .A(n392), .B(n391), .S(n451), .Z(n393) );
  MUX2_X1 U434 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n454), .Z(n394) );
  MUX2_X1 U435 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n453), .Z(n395) );
  MUX2_X1 U436 ( .A(n395), .B(n394), .S(n451), .Z(n396) );
  MUX2_X1 U437 ( .A(n396), .B(n393), .S(N12), .Z(N22) );
  MUX2_X1 U438 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n453), .Z(n397) );
  MUX2_X1 U439 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n453), .Z(n398) );
  MUX2_X1 U440 ( .A(n398), .B(n397), .S(n451), .Z(n399) );
  MUX2_X1 U441 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n453), .Z(n400) );
  MUX2_X1 U442 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n453), .Z(n401) );
  MUX2_X1 U443 ( .A(n401), .B(n400), .S(n451), .Z(n402) );
  MUX2_X1 U444 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n453), .Z(n403) );
  MUX2_X1 U445 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n453), .Z(n404) );
  MUX2_X1 U446 ( .A(n404), .B(n403), .S(n451), .Z(n405) );
  MUX2_X1 U447 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n453), .Z(n406) );
  MUX2_X1 U448 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n453), .Z(n407) );
  MUX2_X1 U449 ( .A(n407), .B(n406), .S(n451), .Z(n408) );
  MUX2_X1 U450 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n453), .Z(n409) );
  MUX2_X1 U451 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n453), .Z(n410) );
  MUX2_X1 U452 ( .A(n410), .B(n409), .S(n451), .Z(n411) );
  MUX2_X1 U453 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n453), .Z(n412) );
  MUX2_X1 U454 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n453), .Z(n413) );
  MUX2_X1 U455 ( .A(n413), .B(n412), .S(n451), .Z(n414) );
  MUX2_X1 U456 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n454), .Z(n415) );
  MUX2_X1 U457 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n454), .Z(n416) );
  MUX2_X1 U458 ( .A(n416), .B(n415), .S(n452), .Z(n417) );
  MUX2_X1 U459 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n454), .Z(n418) );
  MUX2_X1 U460 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n454), .Z(n419) );
  MUX2_X1 U461 ( .A(n419), .B(n418), .S(n452), .Z(n420) );
  MUX2_X1 U462 ( .A(n420), .B(n417), .S(N12), .Z(N18) );
  MUX2_X1 U463 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n454), .Z(n421) );
  MUX2_X1 U464 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n454), .Z(n422) );
  MUX2_X1 U465 ( .A(n422), .B(n421), .S(n452), .Z(n423) );
  MUX2_X1 U466 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n454), .Z(n424) );
  MUX2_X1 U467 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n454), .Z(n425) );
  MUX2_X1 U468 ( .A(n425), .B(n424), .S(n452), .Z(n426) );
  MUX2_X1 U469 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n454), .Z(n427) );
  MUX2_X1 U470 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n454), .Z(n428) );
  MUX2_X1 U471 ( .A(n428), .B(n427), .S(n452), .Z(n429) );
  MUX2_X1 U472 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n454), .Z(n430) );
  MUX2_X1 U473 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n454), .Z(n431) );
  MUX2_X1 U474 ( .A(n431), .B(n430), .S(n452), .Z(n432) );
  MUX2_X1 U475 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n455), .Z(n433) );
  MUX2_X1 U476 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n455), .Z(n434) );
  MUX2_X1 U477 ( .A(n434), .B(n433), .S(N11), .Z(n435) );
  MUX2_X1 U478 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n455), .Z(n436) );
  MUX2_X1 U479 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n455), .Z(n437) );
  MUX2_X1 U480 ( .A(n437), .B(n436), .S(n452), .Z(n438) );
  MUX2_X1 U481 ( .A(n438), .B(n435), .S(N12), .Z(N15) );
  MUX2_X1 U482 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n455), .Z(n439) );
  MUX2_X1 U483 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n455), .Z(n440) );
  MUX2_X1 U484 ( .A(n440), .B(n439), .S(N11), .Z(n441) );
  MUX2_X1 U485 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n455), .Z(n442) );
  MUX2_X1 U486 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n455), .Z(n443) );
  MUX2_X1 U487 ( .A(n443), .B(n442), .S(n452), .Z(n444) );
  MUX2_X1 U488 ( .A(n444), .B(n441), .S(N12), .Z(N14) );
  MUX2_X1 U489 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n455), .Z(n445) );
  MUX2_X1 U490 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n455), .Z(n446) );
  MUX2_X1 U491 ( .A(n446), .B(n445), .S(n452), .Z(n447) );
  MUX2_X1 U492 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n455), .Z(n448) );
  MUX2_X1 U493 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n455), .Z(n449) );
  MUX2_X1 U494 ( .A(n449), .B(n448), .S(n452), .Z(n450) );
  MUX2_X1 U495 ( .A(n450), .B(n447), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH20_SIZE8_LOGSIZE3_1 ( clk, data_in, data_out, addr, wr_en
 );
  input [19:0] data_in;
  output [19:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N14, N16, N18, N22, N24, N26, N28, N30, N32, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[18]  ( .D(N14), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[16]  ( .D(N16), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[14]  ( .D(N18), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[10]  ( .D(N22), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[8]  ( .D(N24), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N26), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N28), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N30), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N32), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][19]  ( .D(n487), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n488), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n489), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n490), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n491), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n492), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n493), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n494), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n495), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n496), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n497), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n498), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n499), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n500), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n501), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n502), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n503), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n504), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n505), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n506), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n507), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n508), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n509), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n510), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n511), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n512), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n513), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n514), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n515), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n516), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n517), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n518), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n519), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n520), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n521), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n522), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n523), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n524), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n525), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n526), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n527), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n528), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n529), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n530), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n531), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n532), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n533), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n534), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n535), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n536), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n537), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n538), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n539), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n540), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n541), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n542), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n543), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n544), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n545), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n546), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n547), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n548), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n549), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n550), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n551), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n552), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n553), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n554), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n555), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n556), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n557), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n558), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n559), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n560), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n561), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n562), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n563), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n564), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n565), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n566), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n567), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n568), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n569), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n570), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n571), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n572), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n573), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n574), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n575), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n576), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n577), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n578), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n579), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n580), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n581), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n582), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n583), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n584), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n585), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n586), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n587), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n588), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n589), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n590), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n591), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n592), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n593), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n594), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n595), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n596), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n597), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n598), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n599), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n600), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n601), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n602), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n603), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n604), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n605), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n606), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n607), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n608), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n609), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n610), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n611), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n612), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n613), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n614), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n615), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n616), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n617), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n618), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n619), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n620), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n621), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n622), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n623), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n624), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n625), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n626), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n627), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n628), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n629), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n630), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n631), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n632), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n633), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n634), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n635), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n636), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n637), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n638), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n639), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n640), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n641), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n642), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n643), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n644), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n645), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n646), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U348 ( .A1(n464), .A2(n465), .A3(n795), .ZN(n816) );
  NAND3_X1 U349 ( .A1(n795), .A2(n465), .A3(N10), .ZN(n794) );
  NAND3_X1 U350 ( .A1(n795), .A2(n464), .A3(N11), .ZN(n773) );
  NAND3_X1 U351 ( .A1(N10), .A2(n795), .A3(N11), .ZN(n752) );
  NAND3_X1 U352 ( .A1(n464), .A2(n465), .A3(n710), .ZN(n731) );
  NAND3_X1 U353 ( .A1(N10), .A2(n465), .A3(n710), .ZN(n709) );
  NAND3_X1 U354 ( .A1(N11), .A2(n464), .A3(n710), .ZN(n688) );
  NAND3_X1 U355 ( .A1(N11), .A2(N10), .A3(n710), .ZN(n667) );
  SDFF_X1 \data_out_reg[9]  ( .D(n390), .SI(n387), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[17]  ( .D(n438), .SI(n435), .SE(N12), .CK(clk), .Q(
        data_out[17]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n12), .SI(n9), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n414), .SI(n411), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n378), .SI(n375), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n354), .SI(n21), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n366), .SI(n363), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n402), .SI(n399), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[19]  ( .D(n450), .SI(n447), .SE(N12), .CK(clk), .Q(
        data_out[19]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n426), .SI(n423), .SE(N12), .CK(clk), .Q(
        data_out[15]) );
  SDFF_X1 \data_out_reg[12]  ( .D(n408), .SI(n405), .SE(N12), .CK(clk), .Q(
        data_out[12]) );
  BUF_X1 U3 ( .A(n773), .Z(n461) );
  BUF_X1 U4 ( .A(n667), .Z(n456) );
  BUF_X1 U5 ( .A(n794), .Z(n462) );
  BUF_X1 U6 ( .A(n452), .Z(n451) );
  BUF_X1 U7 ( .A(n816), .Z(n463) );
  BUF_X1 U8 ( .A(n752), .Z(n460) );
  BUF_X1 U9 ( .A(n709), .Z(n458) );
  BUF_X1 U10 ( .A(n688), .Z(n457) );
  BUF_X1 U11 ( .A(n731), .Z(n459) );
  BUF_X1 U12 ( .A(N10), .Z(n453) );
  BUF_X1 U13 ( .A(N10), .Z(n454) );
  BUF_X1 U14 ( .A(N10), .Z(n455) );
  BUF_X1 U15 ( .A(N11), .Z(n452) );
  NOR2_X1 U16 ( .A1(n466), .A2(N12), .ZN(n795) );
  INV_X1 U17 ( .A(wr_en), .ZN(n466) );
  AND2_X1 U18 ( .A1(N12), .A2(wr_en), .ZN(n710) );
  OAI21_X1 U19 ( .B1(n486), .B2(n794), .A(n793), .ZN(n626) );
  NAND2_X1 U20 ( .A1(\mem[1][0] ), .A2(n794), .ZN(n793) );
  OAI21_X1 U21 ( .B1(n485), .B2(n794), .A(n792), .ZN(n625) );
  NAND2_X1 U22 ( .A1(\mem[1][1] ), .A2(n794), .ZN(n792) );
  OAI21_X1 U23 ( .B1(n484), .B2(n794), .A(n791), .ZN(n624) );
  NAND2_X1 U24 ( .A1(\mem[1][2] ), .A2(n794), .ZN(n791) );
  OAI21_X1 U25 ( .B1(n483), .B2(n462), .A(n790), .ZN(n623) );
  NAND2_X1 U26 ( .A1(\mem[1][3] ), .A2(n794), .ZN(n790) );
  OAI21_X1 U27 ( .B1(n482), .B2(n462), .A(n789), .ZN(n622) );
  NAND2_X1 U28 ( .A1(\mem[1][4] ), .A2(n794), .ZN(n789) );
  OAI21_X1 U29 ( .B1(n481), .B2(n462), .A(n788), .ZN(n621) );
  NAND2_X1 U30 ( .A1(\mem[1][5] ), .A2(n794), .ZN(n788) );
  OAI21_X1 U31 ( .B1(n480), .B2(n462), .A(n787), .ZN(n620) );
  NAND2_X1 U32 ( .A1(\mem[1][6] ), .A2(n794), .ZN(n787) );
  OAI21_X1 U33 ( .B1(n479), .B2(n462), .A(n786), .ZN(n619) );
  NAND2_X1 U34 ( .A1(\mem[1][7] ), .A2(n794), .ZN(n786) );
  OAI21_X1 U35 ( .B1(n478), .B2(n462), .A(n785), .ZN(n618) );
  NAND2_X1 U36 ( .A1(\mem[1][8] ), .A2(n794), .ZN(n785) );
  OAI21_X1 U37 ( .B1(n477), .B2(n462), .A(n784), .ZN(n617) );
  NAND2_X1 U38 ( .A1(\mem[1][9] ), .A2(n794), .ZN(n784) );
  OAI21_X1 U39 ( .B1(n476), .B2(n462), .A(n783), .ZN(n616) );
  NAND2_X1 U40 ( .A1(\mem[1][10] ), .A2(n794), .ZN(n783) );
  OAI21_X1 U41 ( .B1(n475), .B2(n462), .A(n782), .ZN(n615) );
  NAND2_X1 U42 ( .A1(\mem[1][11] ), .A2(n794), .ZN(n782) );
  OAI21_X1 U43 ( .B1(n474), .B2(n462), .A(n781), .ZN(n614) );
  NAND2_X1 U44 ( .A1(\mem[1][12] ), .A2(n794), .ZN(n781) );
  OAI21_X1 U45 ( .B1(n473), .B2(n462), .A(n780), .ZN(n613) );
  NAND2_X1 U46 ( .A1(\mem[1][13] ), .A2(n794), .ZN(n780) );
  OAI21_X1 U47 ( .B1(n472), .B2(n462), .A(n779), .ZN(n612) );
  NAND2_X1 U48 ( .A1(\mem[1][14] ), .A2(n794), .ZN(n779) );
  OAI21_X1 U49 ( .B1(n471), .B2(n462), .A(n778), .ZN(n611) );
  NAND2_X1 U50 ( .A1(\mem[1][15] ), .A2(n794), .ZN(n778) );
  OAI21_X1 U51 ( .B1(n470), .B2(n462), .A(n777), .ZN(n610) );
  NAND2_X1 U52 ( .A1(\mem[1][16] ), .A2(n794), .ZN(n777) );
  OAI21_X1 U53 ( .B1(n469), .B2(n462), .A(n776), .ZN(n609) );
  NAND2_X1 U54 ( .A1(\mem[1][17] ), .A2(n794), .ZN(n776) );
  OAI21_X1 U55 ( .B1(n468), .B2(n462), .A(n775), .ZN(n608) );
  NAND2_X1 U56 ( .A1(\mem[1][18] ), .A2(n794), .ZN(n775) );
  OAI21_X1 U57 ( .B1(n467), .B2(n794), .A(n774), .ZN(n607) );
  NAND2_X1 U58 ( .A1(\mem[1][19] ), .A2(n794), .ZN(n774) );
  OAI21_X1 U59 ( .B1(n486), .B2(n773), .A(n772), .ZN(n606) );
  NAND2_X1 U60 ( .A1(\mem[2][0] ), .A2(n461), .ZN(n772) );
  OAI21_X1 U61 ( .B1(n485), .B2(n773), .A(n771), .ZN(n605) );
  NAND2_X1 U62 ( .A1(\mem[2][1] ), .A2(n461), .ZN(n771) );
  OAI21_X1 U63 ( .B1(n484), .B2(n773), .A(n770), .ZN(n604) );
  NAND2_X1 U64 ( .A1(\mem[2][2] ), .A2(n461), .ZN(n770) );
  OAI21_X1 U65 ( .B1(n483), .B2(n773), .A(n769), .ZN(n603) );
  NAND2_X1 U66 ( .A1(\mem[2][3] ), .A2(n461), .ZN(n769) );
  OAI21_X1 U67 ( .B1(n482), .B2(n461), .A(n768), .ZN(n602) );
  NAND2_X1 U68 ( .A1(\mem[2][4] ), .A2(n461), .ZN(n768) );
  OAI21_X1 U69 ( .B1(n481), .B2(n773), .A(n767), .ZN(n601) );
  NAND2_X1 U70 ( .A1(\mem[2][5] ), .A2(n461), .ZN(n767) );
  OAI21_X1 U71 ( .B1(n480), .B2(n461), .A(n766), .ZN(n600) );
  NAND2_X1 U72 ( .A1(\mem[2][6] ), .A2(n461), .ZN(n766) );
  OAI21_X1 U73 ( .B1(n479), .B2(n773), .A(n765), .ZN(n599) );
  NAND2_X1 U74 ( .A1(\mem[2][7] ), .A2(n461), .ZN(n765) );
  OAI21_X1 U75 ( .B1(n478), .B2(n773), .A(n764), .ZN(n598) );
  NAND2_X1 U76 ( .A1(\mem[2][8] ), .A2(n461), .ZN(n764) );
  OAI21_X1 U77 ( .B1(n477), .B2(n773), .A(n763), .ZN(n597) );
  NAND2_X1 U78 ( .A1(\mem[2][9] ), .A2(n461), .ZN(n763) );
  OAI21_X1 U79 ( .B1(n476), .B2(n773), .A(n762), .ZN(n596) );
  NAND2_X1 U80 ( .A1(\mem[2][10] ), .A2(n461), .ZN(n762) );
  OAI21_X1 U81 ( .B1(n475), .B2(n773), .A(n761), .ZN(n595) );
  NAND2_X1 U82 ( .A1(\mem[2][11] ), .A2(n461), .ZN(n761) );
  OAI21_X1 U83 ( .B1(n474), .B2(n773), .A(n760), .ZN(n594) );
  NAND2_X1 U84 ( .A1(\mem[2][12] ), .A2(n461), .ZN(n760) );
  OAI21_X1 U85 ( .B1(n473), .B2(n773), .A(n759), .ZN(n593) );
  NAND2_X1 U86 ( .A1(\mem[2][13] ), .A2(n773), .ZN(n759) );
  OAI21_X1 U87 ( .B1(n472), .B2(n773), .A(n758), .ZN(n592) );
  NAND2_X1 U88 ( .A1(\mem[2][14] ), .A2(n773), .ZN(n758) );
  OAI21_X1 U89 ( .B1(n471), .B2(n773), .A(n757), .ZN(n591) );
  NAND2_X1 U90 ( .A1(\mem[2][15] ), .A2(n773), .ZN(n757) );
  OAI21_X1 U91 ( .B1(n470), .B2(n773), .A(n756), .ZN(n590) );
  NAND2_X1 U92 ( .A1(\mem[2][16] ), .A2(n773), .ZN(n756) );
  OAI21_X1 U93 ( .B1(n469), .B2(n773), .A(n755), .ZN(n589) );
  NAND2_X1 U94 ( .A1(\mem[2][17] ), .A2(n773), .ZN(n755) );
  OAI21_X1 U95 ( .B1(n468), .B2(n773), .A(n754), .ZN(n588) );
  NAND2_X1 U96 ( .A1(\mem[2][18] ), .A2(n773), .ZN(n754) );
  OAI21_X1 U97 ( .B1(n467), .B2(n461), .A(n753), .ZN(n587) );
  NAND2_X1 U98 ( .A1(\mem[2][19] ), .A2(n461), .ZN(n753) );
  OAI21_X1 U99 ( .B1(n486), .B2(n752), .A(n751), .ZN(n586) );
  NAND2_X1 U100 ( .A1(\mem[3][0] ), .A2(n460), .ZN(n751) );
  OAI21_X1 U101 ( .B1(n485), .B2(n752), .A(n750), .ZN(n585) );
  NAND2_X1 U102 ( .A1(\mem[3][1] ), .A2(n460), .ZN(n750) );
  OAI21_X1 U103 ( .B1(n484), .B2(n752), .A(n749), .ZN(n584) );
  NAND2_X1 U104 ( .A1(\mem[3][2] ), .A2(n460), .ZN(n749) );
  OAI21_X1 U105 ( .B1(n483), .B2(n752), .A(n748), .ZN(n583) );
  NAND2_X1 U106 ( .A1(\mem[3][3] ), .A2(n460), .ZN(n748) );
  OAI21_X1 U107 ( .B1(n482), .B2(n460), .A(n747), .ZN(n582) );
  NAND2_X1 U108 ( .A1(\mem[3][4] ), .A2(n460), .ZN(n747) );
  OAI21_X1 U109 ( .B1(n481), .B2(n460), .A(n746), .ZN(n581) );
  NAND2_X1 U110 ( .A1(\mem[3][5] ), .A2(n460), .ZN(n746) );
  OAI21_X1 U111 ( .B1(n480), .B2(n752), .A(n745), .ZN(n580) );
  NAND2_X1 U112 ( .A1(\mem[3][6] ), .A2(n460), .ZN(n745) );
  OAI21_X1 U113 ( .B1(n479), .B2(n752), .A(n744), .ZN(n579) );
  NAND2_X1 U114 ( .A1(\mem[3][7] ), .A2(n460), .ZN(n744) );
  OAI21_X1 U115 ( .B1(n478), .B2(n752), .A(n743), .ZN(n578) );
  NAND2_X1 U116 ( .A1(\mem[3][8] ), .A2(n460), .ZN(n743) );
  OAI21_X1 U117 ( .B1(n477), .B2(n752), .A(n742), .ZN(n577) );
  NAND2_X1 U118 ( .A1(\mem[3][9] ), .A2(n460), .ZN(n742) );
  OAI21_X1 U119 ( .B1(n476), .B2(n752), .A(n741), .ZN(n576) );
  NAND2_X1 U120 ( .A1(\mem[3][10] ), .A2(n460), .ZN(n741) );
  OAI21_X1 U121 ( .B1(n475), .B2(n752), .A(n740), .ZN(n575) );
  NAND2_X1 U122 ( .A1(\mem[3][11] ), .A2(n460), .ZN(n740) );
  OAI21_X1 U123 ( .B1(n474), .B2(n752), .A(n739), .ZN(n574) );
  NAND2_X1 U124 ( .A1(\mem[3][12] ), .A2(n752), .ZN(n739) );
  OAI21_X1 U125 ( .B1(n473), .B2(n752), .A(n738), .ZN(n573) );
  NAND2_X1 U126 ( .A1(\mem[3][13] ), .A2(n752), .ZN(n738) );
  OAI21_X1 U127 ( .B1(n472), .B2(n752), .A(n737), .ZN(n572) );
  NAND2_X1 U128 ( .A1(\mem[3][14] ), .A2(n752), .ZN(n737) );
  OAI21_X1 U129 ( .B1(n471), .B2(n752), .A(n736), .ZN(n571) );
  NAND2_X1 U130 ( .A1(\mem[3][15] ), .A2(n460), .ZN(n736) );
  OAI21_X1 U131 ( .B1(n470), .B2(n752), .A(n735), .ZN(n570) );
  NAND2_X1 U132 ( .A1(\mem[3][16] ), .A2(n752), .ZN(n735) );
  OAI21_X1 U133 ( .B1(n469), .B2(n752), .A(n734), .ZN(n569) );
  NAND2_X1 U134 ( .A1(\mem[3][17] ), .A2(n752), .ZN(n734) );
  OAI21_X1 U135 ( .B1(n468), .B2(n752), .A(n733), .ZN(n568) );
  NAND2_X1 U136 ( .A1(\mem[3][18] ), .A2(n752), .ZN(n733) );
  OAI21_X1 U137 ( .B1(n467), .B2(n752), .A(n732), .ZN(n567) );
  NAND2_X1 U138 ( .A1(\mem[3][19] ), .A2(n460), .ZN(n732) );
  OAI21_X1 U139 ( .B1(n486), .B2(n731), .A(n730), .ZN(n566) );
  NAND2_X1 U140 ( .A1(\mem[4][0] ), .A2(n731), .ZN(n730) );
  OAI21_X1 U141 ( .B1(n485), .B2(n731), .A(n729), .ZN(n565) );
  NAND2_X1 U142 ( .A1(\mem[4][1] ), .A2(n731), .ZN(n729) );
  OAI21_X1 U143 ( .B1(n484), .B2(n731), .A(n728), .ZN(n564) );
  NAND2_X1 U144 ( .A1(\mem[4][2] ), .A2(n731), .ZN(n728) );
  OAI21_X1 U145 ( .B1(n483), .B2(n459), .A(n727), .ZN(n563) );
  NAND2_X1 U146 ( .A1(\mem[4][3] ), .A2(n459), .ZN(n727) );
  OAI21_X1 U147 ( .B1(n482), .B2(n731), .A(n726), .ZN(n562) );
  NAND2_X1 U148 ( .A1(\mem[4][4] ), .A2(n459), .ZN(n726) );
  OAI21_X1 U149 ( .B1(n481), .B2(n731), .A(n725), .ZN(n561) );
  NAND2_X1 U150 ( .A1(\mem[4][5] ), .A2(n731), .ZN(n725) );
  OAI21_X1 U151 ( .B1(n480), .B2(n731), .A(n724), .ZN(n560) );
  NAND2_X1 U152 ( .A1(\mem[4][6] ), .A2(n731), .ZN(n724) );
  OAI21_X1 U153 ( .B1(n479), .B2(n459), .A(n723), .ZN(n559) );
  NAND2_X1 U154 ( .A1(\mem[4][7] ), .A2(n731), .ZN(n723) );
  OAI21_X1 U155 ( .B1(n478), .B2(n459), .A(n722), .ZN(n558) );
  NAND2_X1 U156 ( .A1(\mem[4][8] ), .A2(n731), .ZN(n722) );
  OAI21_X1 U157 ( .B1(n477), .B2(n459), .A(n721), .ZN(n557) );
  NAND2_X1 U158 ( .A1(\mem[4][9] ), .A2(n731), .ZN(n721) );
  OAI21_X1 U159 ( .B1(n476), .B2(n459), .A(n720), .ZN(n556) );
  NAND2_X1 U160 ( .A1(\mem[4][10] ), .A2(n731), .ZN(n720) );
  OAI21_X1 U161 ( .B1(n475), .B2(n459), .A(n719), .ZN(n555) );
  NAND2_X1 U162 ( .A1(\mem[4][11] ), .A2(n731), .ZN(n719) );
  OAI21_X1 U163 ( .B1(n474), .B2(n731), .A(n718), .ZN(n554) );
  NAND2_X1 U164 ( .A1(\mem[4][12] ), .A2(n459), .ZN(n718) );
  OAI21_X1 U165 ( .B1(n473), .B2(n731), .A(n717), .ZN(n553) );
  NAND2_X1 U166 ( .A1(\mem[4][13] ), .A2(n459), .ZN(n717) );
  OAI21_X1 U167 ( .B1(n472), .B2(n731), .A(n716), .ZN(n552) );
  NAND2_X1 U168 ( .A1(\mem[4][14] ), .A2(n459), .ZN(n716) );
  OAI21_X1 U169 ( .B1(n471), .B2(n731), .A(n715), .ZN(n551) );
  NAND2_X1 U170 ( .A1(\mem[4][15] ), .A2(n459), .ZN(n715) );
  OAI21_X1 U171 ( .B1(n470), .B2(n731), .A(n714), .ZN(n550) );
  NAND2_X1 U172 ( .A1(\mem[4][16] ), .A2(n459), .ZN(n714) );
  OAI21_X1 U173 ( .B1(n469), .B2(n731), .A(n713), .ZN(n549) );
  NAND2_X1 U174 ( .A1(\mem[4][17] ), .A2(n459), .ZN(n713) );
  OAI21_X1 U175 ( .B1(n468), .B2(n731), .A(n712), .ZN(n548) );
  NAND2_X1 U176 ( .A1(\mem[4][18] ), .A2(n459), .ZN(n712) );
  OAI21_X1 U177 ( .B1(n467), .B2(n731), .A(n711), .ZN(n547) );
  NAND2_X1 U178 ( .A1(\mem[4][19] ), .A2(n459), .ZN(n711) );
  OAI21_X1 U179 ( .B1(n486), .B2(n709), .A(n708), .ZN(n546) );
  NAND2_X1 U180 ( .A1(\mem[5][0] ), .A2(n458), .ZN(n708) );
  OAI21_X1 U181 ( .B1(n485), .B2(n709), .A(n707), .ZN(n545) );
  NAND2_X1 U182 ( .A1(\mem[5][1] ), .A2(n458), .ZN(n707) );
  OAI21_X1 U183 ( .B1(n484), .B2(n709), .A(n706), .ZN(n544) );
  NAND2_X1 U184 ( .A1(\mem[5][2] ), .A2(n458), .ZN(n706) );
  OAI21_X1 U185 ( .B1(n483), .B2(n709), .A(n705), .ZN(n543) );
  NAND2_X1 U186 ( .A1(\mem[5][3] ), .A2(n458), .ZN(n705) );
  OAI21_X1 U187 ( .B1(n482), .B2(n458), .A(n704), .ZN(n542) );
  NAND2_X1 U188 ( .A1(\mem[5][4] ), .A2(n458), .ZN(n704) );
  OAI21_X1 U189 ( .B1(n481), .B2(n709), .A(n703), .ZN(n541) );
  NAND2_X1 U190 ( .A1(\mem[5][5] ), .A2(n458), .ZN(n703) );
  OAI21_X1 U191 ( .B1(n480), .B2(n709), .A(n702), .ZN(n540) );
  NAND2_X1 U192 ( .A1(\mem[5][6] ), .A2(n458), .ZN(n702) );
  OAI21_X1 U193 ( .B1(n479), .B2(n709), .A(n701), .ZN(n539) );
  NAND2_X1 U194 ( .A1(\mem[5][7] ), .A2(n458), .ZN(n701) );
  OAI21_X1 U195 ( .B1(n478), .B2(n709), .A(n700), .ZN(n538) );
  NAND2_X1 U196 ( .A1(\mem[5][8] ), .A2(n458), .ZN(n700) );
  OAI21_X1 U197 ( .B1(n477), .B2(n709), .A(n699), .ZN(n537) );
  NAND2_X1 U198 ( .A1(\mem[5][9] ), .A2(n458), .ZN(n699) );
  OAI21_X1 U199 ( .B1(n476), .B2(n709), .A(n698), .ZN(n536) );
  NAND2_X1 U200 ( .A1(\mem[5][10] ), .A2(n458), .ZN(n698) );
  OAI21_X1 U201 ( .B1(n475), .B2(n709), .A(n697), .ZN(n535) );
  NAND2_X1 U202 ( .A1(\mem[5][11] ), .A2(n458), .ZN(n697) );
  OAI21_X1 U203 ( .B1(n474), .B2(n709), .A(n696), .ZN(n534) );
  NAND2_X1 U204 ( .A1(\mem[5][12] ), .A2(n709), .ZN(n696) );
  OAI21_X1 U205 ( .B1(n473), .B2(n458), .A(n695), .ZN(n533) );
  NAND2_X1 U206 ( .A1(\mem[5][13] ), .A2(n709), .ZN(n695) );
  OAI21_X1 U207 ( .B1(n472), .B2(n458), .A(n694), .ZN(n532) );
  NAND2_X1 U208 ( .A1(\mem[5][14] ), .A2(n709), .ZN(n694) );
  OAI21_X1 U209 ( .B1(n471), .B2(n709), .A(n693), .ZN(n531) );
  NAND2_X1 U210 ( .A1(\mem[5][15] ), .A2(n709), .ZN(n693) );
  OAI21_X1 U211 ( .B1(n470), .B2(n709), .A(n692), .ZN(n530) );
  NAND2_X1 U212 ( .A1(\mem[5][16] ), .A2(n709), .ZN(n692) );
  OAI21_X1 U213 ( .B1(n469), .B2(n709), .A(n691), .ZN(n529) );
  NAND2_X1 U214 ( .A1(\mem[5][17] ), .A2(n709), .ZN(n691) );
  OAI21_X1 U215 ( .B1(n468), .B2(n709), .A(n690), .ZN(n528) );
  NAND2_X1 U216 ( .A1(\mem[5][18] ), .A2(n709), .ZN(n690) );
  OAI21_X1 U217 ( .B1(n467), .B2(n709), .A(n689), .ZN(n527) );
  NAND2_X1 U218 ( .A1(\mem[5][19] ), .A2(n458), .ZN(n689) );
  OAI21_X1 U219 ( .B1(n486), .B2(n457), .A(n687), .ZN(n526) );
  NAND2_X1 U220 ( .A1(\mem[6][0] ), .A2(n688), .ZN(n687) );
  OAI21_X1 U221 ( .B1(n485), .B2(n457), .A(n686), .ZN(n525) );
  NAND2_X1 U222 ( .A1(\mem[6][1] ), .A2(n688), .ZN(n686) );
  OAI21_X1 U223 ( .B1(n484), .B2(n457), .A(n685), .ZN(n524) );
  NAND2_X1 U224 ( .A1(\mem[6][2] ), .A2(n688), .ZN(n685) );
  OAI21_X1 U225 ( .B1(n483), .B2(n688), .A(n684), .ZN(n523) );
  NAND2_X1 U226 ( .A1(\mem[6][3] ), .A2(n457), .ZN(n684) );
  OAI21_X1 U227 ( .B1(n482), .B2(n688), .A(n683), .ZN(n522) );
  NAND2_X1 U228 ( .A1(\mem[6][4] ), .A2(n457), .ZN(n683) );
  OAI21_X1 U229 ( .B1(n481), .B2(n688), .A(n682), .ZN(n521) );
  NAND2_X1 U230 ( .A1(\mem[6][5] ), .A2(n688), .ZN(n682) );
  OAI21_X1 U231 ( .B1(n480), .B2(n688), .A(n681), .ZN(n520) );
  NAND2_X1 U232 ( .A1(\mem[6][6] ), .A2(n688), .ZN(n681) );
  OAI21_X1 U233 ( .B1(n479), .B2(n688), .A(n680), .ZN(n519) );
  NAND2_X1 U234 ( .A1(\mem[6][7] ), .A2(n688), .ZN(n680) );
  OAI21_X1 U235 ( .B1(n478), .B2(n688), .A(n679), .ZN(n518) );
  NAND2_X1 U236 ( .A1(\mem[6][8] ), .A2(n688), .ZN(n679) );
  OAI21_X1 U237 ( .B1(n477), .B2(n457), .A(n678), .ZN(n517) );
  NAND2_X1 U238 ( .A1(\mem[6][9] ), .A2(n688), .ZN(n678) );
  OAI21_X1 U239 ( .B1(n476), .B2(n688), .A(n677), .ZN(n516) );
  NAND2_X1 U240 ( .A1(\mem[6][10] ), .A2(n688), .ZN(n677) );
  OAI21_X1 U241 ( .B1(n475), .B2(n688), .A(n676), .ZN(n515) );
  NAND2_X1 U242 ( .A1(\mem[6][11] ), .A2(n688), .ZN(n676) );
  OAI21_X1 U243 ( .B1(n474), .B2(n688), .A(n675), .ZN(n514) );
  NAND2_X1 U244 ( .A1(\mem[6][12] ), .A2(n457), .ZN(n675) );
  OAI21_X1 U245 ( .B1(n473), .B2(n457), .A(n674), .ZN(n513) );
  NAND2_X1 U246 ( .A1(\mem[6][13] ), .A2(n457), .ZN(n674) );
  OAI21_X1 U247 ( .B1(n472), .B2(n688), .A(n673), .ZN(n512) );
  NAND2_X1 U248 ( .A1(\mem[6][14] ), .A2(n457), .ZN(n673) );
  OAI21_X1 U249 ( .B1(n471), .B2(n688), .A(n672), .ZN(n511) );
  NAND2_X1 U250 ( .A1(\mem[6][15] ), .A2(n457), .ZN(n672) );
  OAI21_X1 U251 ( .B1(n470), .B2(n688), .A(n671), .ZN(n510) );
  NAND2_X1 U252 ( .A1(\mem[6][16] ), .A2(n457), .ZN(n671) );
  OAI21_X1 U253 ( .B1(n469), .B2(n688), .A(n670), .ZN(n509) );
  NAND2_X1 U254 ( .A1(\mem[6][17] ), .A2(n457), .ZN(n670) );
  OAI21_X1 U255 ( .B1(n468), .B2(n688), .A(n669), .ZN(n508) );
  NAND2_X1 U256 ( .A1(\mem[6][18] ), .A2(n457), .ZN(n669) );
  OAI21_X1 U257 ( .B1(n467), .B2(n457), .A(n668), .ZN(n507) );
  NAND2_X1 U258 ( .A1(\mem[6][19] ), .A2(n457), .ZN(n668) );
  OAI21_X1 U259 ( .B1(n486), .B2(n667), .A(n666), .ZN(n506) );
  NAND2_X1 U260 ( .A1(\mem[7][0] ), .A2(n456), .ZN(n666) );
  OAI21_X1 U261 ( .B1(n485), .B2(n456), .A(n665), .ZN(n505) );
  NAND2_X1 U262 ( .A1(\mem[7][1] ), .A2(n456), .ZN(n665) );
  OAI21_X1 U263 ( .B1(n484), .B2(n667), .A(n664), .ZN(n504) );
  NAND2_X1 U264 ( .A1(\mem[7][2] ), .A2(n456), .ZN(n664) );
  OAI21_X1 U265 ( .B1(n483), .B2(n667), .A(n663), .ZN(n503) );
  NAND2_X1 U266 ( .A1(\mem[7][3] ), .A2(n456), .ZN(n663) );
  OAI21_X1 U267 ( .B1(n482), .B2(n456), .A(n662), .ZN(n502) );
  NAND2_X1 U268 ( .A1(\mem[7][4] ), .A2(n456), .ZN(n662) );
  OAI21_X1 U269 ( .B1(n481), .B2(n667), .A(n661), .ZN(n501) );
  NAND2_X1 U270 ( .A1(\mem[7][5] ), .A2(n456), .ZN(n661) );
  OAI21_X1 U271 ( .B1(n480), .B2(n667), .A(n660), .ZN(n500) );
  NAND2_X1 U272 ( .A1(\mem[7][6] ), .A2(n456), .ZN(n660) );
  OAI21_X1 U273 ( .B1(n479), .B2(n667), .A(n659), .ZN(n499) );
  NAND2_X1 U274 ( .A1(\mem[7][7] ), .A2(n456), .ZN(n659) );
  OAI21_X1 U275 ( .B1(n478), .B2(n667), .A(n658), .ZN(n498) );
  NAND2_X1 U276 ( .A1(\mem[7][8] ), .A2(n456), .ZN(n658) );
  OAI21_X1 U277 ( .B1(n477), .B2(n667), .A(n657), .ZN(n497) );
  NAND2_X1 U278 ( .A1(\mem[7][9] ), .A2(n456), .ZN(n657) );
  OAI21_X1 U279 ( .B1(n476), .B2(n667), .A(n656), .ZN(n496) );
  NAND2_X1 U280 ( .A1(\mem[7][10] ), .A2(n456), .ZN(n656) );
  OAI21_X1 U281 ( .B1(n475), .B2(n667), .A(n655), .ZN(n495) );
  NAND2_X1 U282 ( .A1(\mem[7][11] ), .A2(n456), .ZN(n655) );
  OAI21_X1 U283 ( .B1(n474), .B2(n667), .A(n654), .ZN(n494) );
  NAND2_X1 U284 ( .A1(\mem[7][12] ), .A2(n667), .ZN(n654) );
  OAI21_X1 U285 ( .B1(n473), .B2(n667), .A(n653), .ZN(n493) );
  NAND2_X1 U286 ( .A1(\mem[7][13] ), .A2(n667), .ZN(n653) );
  OAI21_X1 U287 ( .B1(n472), .B2(n667), .A(n652), .ZN(n492) );
  NAND2_X1 U288 ( .A1(\mem[7][14] ), .A2(n667), .ZN(n652) );
  OAI21_X1 U289 ( .B1(n471), .B2(n667), .A(n651), .ZN(n491) );
  NAND2_X1 U290 ( .A1(\mem[7][15] ), .A2(n667), .ZN(n651) );
  OAI21_X1 U291 ( .B1(n470), .B2(n667), .A(n650), .ZN(n490) );
  NAND2_X1 U292 ( .A1(\mem[7][16] ), .A2(n667), .ZN(n650) );
  OAI21_X1 U293 ( .B1(n469), .B2(n667), .A(n649), .ZN(n489) );
  NAND2_X1 U294 ( .A1(\mem[7][17] ), .A2(n667), .ZN(n649) );
  OAI21_X1 U295 ( .B1(n468), .B2(n667), .A(n648), .ZN(n488) );
  NAND2_X1 U296 ( .A1(\mem[7][18] ), .A2(n667), .ZN(n648) );
  OAI21_X1 U297 ( .B1(n467), .B2(n456), .A(n647), .ZN(n487) );
  NAND2_X1 U298 ( .A1(\mem[7][19] ), .A2(n456), .ZN(n647) );
  OAI21_X1 U299 ( .B1(n816), .B2(n484), .A(n813), .ZN(n644) );
  NAND2_X1 U300 ( .A1(\mem[0][2] ), .A2(n463), .ZN(n813) );
  OAI21_X1 U301 ( .B1(n816), .B2(n483), .A(n812), .ZN(n643) );
  NAND2_X1 U302 ( .A1(\mem[0][3] ), .A2(n463), .ZN(n812) );
  OAI21_X1 U303 ( .B1(n816), .B2(n482), .A(n811), .ZN(n642) );
  NAND2_X1 U304 ( .A1(\mem[0][4] ), .A2(n463), .ZN(n811) );
  OAI21_X1 U305 ( .B1(n816), .B2(n481), .A(n810), .ZN(n641) );
  NAND2_X1 U306 ( .A1(\mem[0][5] ), .A2(n463), .ZN(n810) );
  OAI21_X1 U307 ( .B1(n816), .B2(n480), .A(n809), .ZN(n640) );
  NAND2_X1 U308 ( .A1(\mem[0][6] ), .A2(n463), .ZN(n809) );
  OAI21_X1 U309 ( .B1(n816), .B2(n479), .A(n808), .ZN(n639) );
  NAND2_X1 U310 ( .A1(\mem[0][7] ), .A2(n463), .ZN(n808) );
  OAI21_X1 U311 ( .B1(n816), .B2(n478), .A(n807), .ZN(n638) );
  NAND2_X1 U312 ( .A1(\mem[0][8] ), .A2(n463), .ZN(n807) );
  OAI21_X1 U313 ( .B1(n816), .B2(n477), .A(n806), .ZN(n637) );
  NAND2_X1 U314 ( .A1(\mem[0][9] ), .A2(n463), .ZN(n806) );
  OAI21_X1 U315 ( .B1(n816), .B2(n476), .A(n805), .ZN(n636) );
  NAND2_X1 U316 ( .A1(\mem[0][10] ), .A2(n463), .ZN(n805) );
  OAI21_X1 U317 ( .B1(n816), .B2(n475), .A(n804), .ZN(n635) );
  NAND2_X1 U318 ( .A1(\mem[0][11] ), .A2(n463), .ZN(n804) );
  OAI21_X1 U319 ( .B1(n816), .B2(n474), .A(n803), .ZN(n634) );
  NAND2_X1 U320 ( .A1(\mem[0][12] ), .A2(n816), .ZN(n803) );
  OAI21_X1 U321 ( .B1(n816), .B2(n473), .A(n802), .ZN(n633) );
  NAND2_X1 U322 ( .A1(\mem[0][13] ), .A2(n816), .ZN(n802) );
  OAI21_X1 U323 ( .B1(n463), .B2(n472), .A(n801), .ZN(n632) );
  NAND2_X1 U324 ( .A1(\mem[0][14] ), .A2(n816), .ZN(n801) );
  OAI21_X1 U325 ( .B1(n816), .B2(n471), .A(n800), .ZN(n631) );
  NAND2_X1 U326 ( .A1(\mem[0][15] ), .A2(n463), .ZN(n800) );
  OAI21_X1 U327 ( .B1(n816), .B2(n470), .A(n799), .ZN(n630) );
  NAND2_X1 U328 ( .A1(\mem[0][16] ), .A2(n816), .ZN(n799) );
  OAI21_X1 U329 ( .B1(n816), .B2(n469), .A(n798), .ZN(n629) );
  NAND2_X1 U330 ( .A1(\mem[0][17] ), .A2(n816), .ZN(n798) );
  OAI21_X1 U331 ( .B1(n816), .B2(n468), .A(n797), .ZN(n628) );
  NAND2_X1 U332 ( .A1(\mem[0][18] ), .A2(n816), .ZN(n797) );
  OAI21_X1 U333 ( .B1(n463), .B2(n486), .A(n815), .ZN(n646) );
  NAND2_X1 U334 ( .A1(\mem[0][0] ), .A2(n463), .ZN(n815) );
  OAI21_X1 U335 ( .B1(n816), .B2(n485), .A(n814), .ZN(n645) );
  NAND2_X1 U336 ( .A1(\mem[0][1] ), .A2(n463), .ZN(n814) );
  OAI21_X1 U337 ( .B1(n816), .B2(n467), .A(n796), .ZN(n627) );
  NAND2_X1 U338 ( .A1(\mem[0][19] ), .A2(n463), .ZN(n796) );
  INV_X1 U339 ( .A(N10), .ZN(n464) );
  INV_X1 U340 ( .A(N11), .ZN(n465) );
  INV_X1 U341 ( .A(data_in[0]), .ZN(n486) );
  INV_X1 U342 ( .A(data_in[1]), .ZN(n485) );
  INV_X1 U343 ( .A(data_in[2]), .ZN(n484) );
  INV_X1 U344 ( .A(data_in[3]), .ZN(n483) );
  INV_X1 U345 ( .A(data_in[4]), .ZN(n482) );
  INV_X1 U346 ( .A(data_in[5]), .ZN(n481) );
  INV_X1 U347 ( .A(data_in[6]), .ZN(n480) );
  INV_X1 U356 ( .A(data_in[7]), .ZN(n479) );
  INV_X1 U357 ( .A(data_in[8]), .ZN(n478) );
  INV_X1 U358 ( .A(data_in[9]), .ZN(n477) );
  INV_X1 U359 ( .A(data_in[10]), .ZN(n476) );
  INV_X1 U360 ( .A(data_in[11]), .ZN(n475) );
  INV_X1 U361 ( .A(data_in[12]), .ZN(n474) );
  INV_X1 U362 ( .A(data_in[13]), .ZN(n473) );
  INV_X1 U363 ( .A(data_in[14]), .ZN(n472) );
  INV_X1 U364 ( .A(data_in[15]), .ZN(n471) );
  INV_X1 U365 ( .A(data_in[16]), .ZN(n470) );
  INV_X1 U366 ( .A(data_in[17]), .ZN(n469) );
  INV_X1 U367 ( .A(data_in[18]), .ZN(n468) );
  INV_X1 U368 ( .A(data_in[19]), .ZN(n467) );
  MUX2_X1 U369 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n455), .Z(n1) );
  MUX2_X1 U370 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n453), .Z(n2) );
  MUX2_X1 U371 ( .A(n2), .B(n1), .S(n452), .Z(n3) );
  MUX2_X1 U372 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(N10), .Z(n4) );
  MUX2_X1 U373 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n454), .Z(n5) );
  MUX2_X1 U374 ( .A(n5), .B(n4), .S(N11), .Z(n6) );
  MUX2_X1 U375 ( .A(n6), .B(n3), .S(N12), .Z(N32) );
  MUX2_X1 U376 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(N10), .Z(n7) );
  MUX2_X1 U377 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n453), .Z(n8) );
  MUX2_X1 U378 ( .A(n8), .B(n7), .S(N11), .Z(n9) );
  MUX2_X1 U379 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n455), .Z(n10) );
  MUX2_X1 U380 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n453), .Z(n11) );
  MUX2_X1 U381 ( .A(n11), .B(n10), .S(N11), .Z(n12) );
  MUX2_X1 U382 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n454), .Z(n13) );
  MUX2_X1 U383 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(N10), .Z(n14) );
  MUX2_X1 U384 ( .A(n14), .B(n13), .S(n451), .Z(n15) );
  MUX2_X1 U385 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n453), .Z(n16) );
  MUX2_X1 U386 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n455), .Z(n17) );
  MUX2_X1 U387 ( .A(n17), .B(n16), .S(n451), .Z(n18) );
  MUX2_X1 U388 ( .A(n18), .B(n15), .S(N12), .Z(N30) );
  MUX2_X1 U389 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n454), .Z(n19) );
  MUX2_X1 U390 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n20) );
  MUX2_X1 U391 ( .A(n20), .B(n19), .S(n451), .Z(n21) );
  MUX2_X1 U392 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n454), .Z(n22) );
  MUX2_X1 U393 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n455), .Z(n23) );
  MUX2_X1 U394 ( .A(n23), .B(n22), .S(n451), .Z(n354) );
  MUX2_X1 U395 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n454), .Z(n355) );
  MUX2_X1 U396 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n453), .Z(n356) );
  MUX2_X1 U397 ( .A(n356), .B(n355), .S(n451), .Z(n357) );
  MUX2_X1 U398 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n454), .Z(n358) );
  MUX2_X1 U399 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n453), .Z(n359) );
  MUX2_X1 U400 ( .A(n359), .B(n358), .S(n451), .Z(n360) );
  MUX2_X1 U401 ( .A(n360), .B(n357), .S(N12), .Z(N28) );
  MUX2_X1 U402 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n453), .Z(n361) );
  MUX2_X1 U403 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n453), .Z(n362) );
  MUX2_X1 U404 ( .A(n362), .B(n361), .S(n451), .Z(n363) );
  MUX2_X1 U405 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n453), .Z(n364) );
  MUX2_X1 U406 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n453), .Z(n365) );
  MUX2_X1 U407 ( .A(n365), .B(n364), .S(n451), .Z(n366) );
  MUX2_X1 U408 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n453), .Z(n367) );
  MUX2_X1 U409 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n453), .Z(n368) );
  MUX2_X1 U410 ( .A(n368), .B(n367), .S(n451), .Z(n369) );
  MUX2_X1 U411 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n453), .Z(n370) );
  MUX2_X1 U412 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n453), .Z(n371) );
  MUX2_X1 U413 ( .A(n371), .B(n370), .S(n451), .Z(n372) );
  MUX2_X1 U414 ( .A(n372), .B(n369), .S(N12), .Z(N26) );
  MUX2_X1 U415 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n453), .Z(n373) );
  MUX2_X1 U416 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n453), .Z(n374) );
  MUX2_X1 U417 ( .A(n374), .B(n373), .S(n451), .Z(n375) );
  MUX2_X1 U418 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n453), .Z(n376) );
  MUX2_X1 U419 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n453), .Z(n377) );
  MUX2_X1 U420 ( .A(n377), .B(n376), .S(n451), .Z(n378) );
  MUX2_X1 U421 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n454), .Z(n379) );
  MUX2_X1 U422 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n454), .Z(n380) );
  MUX2_X1 U423 ( .A(n380), .B(n379), .S(n452), .Z(n381) );
  MUX2_X1 U424 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n454), .Z(n382) );
  MUX2_X1 U425 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n454), .Z(n383) );
  MUX2_X1 U426 ( .A(n383), .B(n382), .S(n452), .Z(n384) );
  MUX2_X1 U427 ( .A(n384), .B(n381), .S(N12), .Z(N24) );
  MUX2_X1 U428 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n454), .Z(n385) );
  MUX2_X1 U429 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n454), .Z(n386) );
  MUX2_X1 U430 ( .A(n386), .B(n385), .S(n452), .Z(n387) );
  MUX2_X1 U431 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n454), .Z(n388) );
  MUX2_X1 U432 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n454), .Z(n389) );
  MUX2_X1 U433 ( .A(n389), .B(n388), .S(n452), .Z(n390) );
  MUX2_X1 U434 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n454), .Z(n391) );
  MUX2_X1 U435 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n454), .Z(n392) );
  MUX2_X1 U436 ( .A(n392), .B(n391), .S(n452), .Z(n393) );
  MUX2_X1 U437 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n454), .Z(n394) );
  MUX2_X1 U438 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n454), .Z(n395) );
  MUX2_X1 U439 ( .A(n395), .B(n394), .S(n452), .Z(n396) );
  MUX2_X1 U440 ( .A(n396), .B(n393), .S(N12), .Z(N22) );
  MUX2_X1 U441 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n455), .Z(n397) );
  MUX2_X1 U442 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n455), .Z(n398) );
  MUX2_X1 U443 ( .A(n398), .B(n397), .S(n452), .Z(n399) );
  MUX2_X1 U444 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n455), .Z(n400) );
  MUX2_X1 U445 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n455), .Z(n401) );
  MUX2_X1 U446 ( .A(n401), .B(n400), .S(n452), .Z(n402) );
  MUX2_X1 U447 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n455), .Z(n403) );
  MUX2_X1 U448 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n455), .Z(n404) );
  MUX2_X1 U449 ( .A(n404), .B(n403), .S(n452), .Z(n405) );
  MUX2_X1 U450 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n455), .Z(n406) );
  MUX2_X1 U451 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n455), .Z(n407) );
  MUX2_X1 U452 ( .A(n407), .B(n406), .S(n452), .Z(n408) );
  MUX2_X1 U453 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n455), .Z(n409) );
  MUX2_X1 U454 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n455), .Z(n410) );
  MUX2_X1 U455 ( .A(n410), .B(n409), .S(n452), .Z(n411) );
  MUX2_X1 U456 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n455), .Z(n412) );
  MUX2_X1 U457 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n455), .Z(n413) );
  MUX2_X1 U458 ( .A(n413), .B(n412), .S(n452), .Z(n414) );
  MUX2_X1 U459 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n454), .Z(n415) );
  MUX2_X1 U460 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n453), .Z(n416) );
  MUX2_X1 U461 ( .A(n416), .B(n415), .S(n452), .Z(n417) );
  MUX2_X1 U462 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n455), .Z(n418) );
  MUX2_X1 U463 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n453), .Z(n419) );
  MUX2_X1 U464 ( .A(n419), .B(n418), .S(n452), .Z(n420) );
  MUX2_X1 U465 ( .A(n420), .B(n417), .S(N12), .Z(N18) );
  MUX2_X1 U466 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(N10), .Z(n421) );
  MUX2_X1 U467 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(N10), .Z(n422) );
  MUX2_X1 U468 ( .A(n422), .B(n421), .S(N11), .Z(n423) );
  MUX2_X1 U469 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(N10), .Z(n424) );
  MUX2_X1 U470 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(N10), .Z(n425) );
  MUX2_X1 U471 ( .A(n425), .B(n424), .S(n452), .Z(n426) );
  MUX2_X1 U472 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(n453), .Z(n427) );
  MUX2_X1 U473 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n455), .Z(n428) );
  MUX2_X1 U474 ( .A(n428), .B(n427), .S(n452), .Z(n429) );
  MUX2_X1 U475 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n454), .Z(n430) );
  MUX2_X1 U476 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n455), .Z(n431) );
  MUX2_X1 U477 ( .A(n431), .B(n430), .S(n452), .Z(n432) );
  MUX2_X1 U478 ( .A(n432), .B(n429), .S(N12), .Z(N16) );
  MUX2_X1 U479 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(N10), .Z(n433) );
  MUX2_X1 U480 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n454), .Z(n434) );
  MUX2_X1 U481 ( .A(n434), .B(n433), .S(N11), .Z(n435) );
  MUX2_X1 U482 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n455), .Z(n436) );
  MUX2_X1 U483 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(N10), .Z(n437) );
  MUX2_X1 U484 ( .A(n437), .B(n436), .S(n452), .Z(n438) );
  MUX2_X1 U485 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n454), .Z(n439) );
  MUX2_X1 U486 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n453), .Z(n440) );
  MUX2_X1 U487 ( .A(n440), .B(n439), .S(n452), .Z(n441) );
  MUX2_X1 U488 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n455), .Z(n442) );
  MUX2_X1 U489 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n454), .Z(n443) );
  MUX2_X1 U490 ( .A(n443), .B(n442), .S(n451), .Z(n444) );
  MUX2_X1 U491 ( .A(n444), .B(n441), .S(N12), .Z(N14) );
  MUX2_X1 U492 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n455), .Z(n445) );
  MUX2_X1 U493 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(N10), .Z(n446) );
  MUX2_X1 U494 ( .A(n446), .B(n445), .S(n452), .Z(n447) );
  MUX2_X1 U495 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n453), .Z(n448) );
  MUX2_X1 U496 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n455), .Z(n449) );
  MUX2_X1 U497 ( .A(n449), .B(n448), .S(n452), .Z(n450) );
endmodule


module memory_WIDTH40_SIZE8_LOGSIZE3 ( clk, data_in, data_out, addr, wr_en );
  input [39:0] data_in;
  output [39:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][39] , \mem[7][38] , \mem[7][37] , \mem[7][36] ,
         \mem[7][35] , \mem[7][34] , \mem[7][33] , \mem[7][32] , \mem[7][31] ,
         \mem[7][30] , \mem[7][29] , \mem[7][28] , \mem[7][27] , \mem[7][26] ,
         \mem[7][25] , \mem[7][24] , \mem[7][23] , \mem[7][22] , \mem[7][21] ,
         \mem[7][20] , \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] ,
         \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] ,
         \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] ,
         \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] ,
         \mem[7][0] , \mem[6][39] , \mem[6][38] , \mem[6][37] , \mem[6][36] ,
         \mem[6][35] , \mem[6][34] , \mem[6][33] , \mem[6][32] , \mem[6][31] ,
         \mem[6][30] , \mem[6][29] , \mem[6][28] , \mem[6][27] , \mem[6][26] ,
         \mem[6][25] , \mem[6][24] , \mem[6][23] , \mem[6][22] , \mem[6][21] ,
         \mem[6][20] , \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] ,
         \mem[6][15] , \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] ,
         \mem[6][10] , \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] ,
         \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] ,
         \mem[6][0] , \mem[5][39] , \mem[5][38] , \mem[5][37] , \mem[5][36] ,
         \mem[5][35] , \mem[5][34] , \mem[5][33] , \mem[5][32] , \mem[5][31] ,
         \mem[5][30] , \mem[5][29] , \mem[5][28] , \mem[5][27] , \mem[5][26] ,
         \mem[5][25] , \mem[5][24] , \mem[5][23] , \mem[5][22] , \mem[5][21] ,
         \mem[5][20] , \mem[5][19] , \mem[5][18] , \mem[5][17] , \mem[5][16] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][39] , \mem[4][38] , \mem[4][37] , \mem[4][36] ,
         \mem[4][35] , \mem[4][34] , \mem[4][33] , \mem[4][32] , \mem[4][31] ,
         \mem[4][30] , \mem[4][29] , \mem[4][28] , \mem[4][27] , \mem[4][26] ,
         \mem[4][25] , \mem[4][24] , \mem[4][23] , \mem[4][22] , \mem[4][21] ,
         \mem[4][20] , \mem[4][19] , \mem[4][18] , \mem[4][17] , \mem[4][16] ,
         \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] ,
         \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][39] , \mem[3][38] , \mem[3][37] , \mem[3][36] ,
         \mem[3][35] , \mem[3][34] , \mem[3][33] , \mem[3][32] , \mem[3][31] ,
         \mem[3][30] , \mem[3][29] , \mem[3][28] , \mem[3][27] , \mem[3][26] ,
         \mem[3][25] , \mem[3][24] , \mem[3][23] , \mem[3][22] , \mem[3][21] ,
         \mem[3][20] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][39] , \mem[2][38] , \mem[2][37] , \mem[2][36] ,
         \mem[2][35] , \mem[2][34] , \mem[2][33] , \mem[2][32] , \mem[2][31] ,
         \mem[2][30] , \mem[2][29] , \mem[2][28] , \mem[2][27] , \mem[2][26] ,
         \mem[2][25] , \mem[2][24] , \mem[2][23] , \mem[2][22] , \mem[2][21] ,
         \mem[2][20] , \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] ,
         \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] ,
         \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] ,
         \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] ,
         \mem[2][0] , \mem[1][39] , \mem[1][38] , \mem[1][37] , \mem[1][36] ,
         \mem[1][35] , \mem[1][34] , \mem[1][33] , \mem[1][32] , \mem[1][31] ,
         \mem[1][30] , \mem[1][29] , \mem[1][28] , \mem[1][27] , \mem[1][26] ,
         \mem[1][25] , \mem[1][24] , \mem[1][23] , \mem[1][22] , \mem[1][21] ,
         \mem[1][20] , \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] ,
         \mem[1][15] , \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] ,
         \mem[1][10] , \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] ,
         \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] ,
         \mem[1][0] , \mem[0][39] , \mem[0][38] , \mem[0][37] , \mem[0][36] ,
         \mem[0][35] , \mem[0][34] , \mem[0][33] , \mem[0][32] , \mem[0][31] ,
         \mem[0][30] , \mem[0][29] , \mem[0][28] , \mem[0][27] , \mem[0][26] ,
         \mem[0][25] , \mem[0][24] , \mem[0][23] , \mem[0][22] , \mem[0][21] ,
         \mem[0][20] , \mem[0][19] , \mem[0][18] , \mem[0][17] , \mem[0][16] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51,
         N52, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[39]  ( .D(N13), .CK(clk), .Q(data_out[39]) );
  DFF_X1 \data_out_reg[38]  ( .D(N14), .CK(clk), .Q(data_out[38]) );
  DFF_X1 \data_out_reg[37]  ( .D(N15), .CK(clk), .Q(data_out[37]) );
  DFF_X1 \data_out_reg[36]  ( .D(N16), .CK(clk), .Q(data_out[36]) );
  DFF_X1 \data_out_reg[35]  ( .D(N17), .CK(clk), .Q(data_out[35]) );
  DFF_X1 \data_out_reg[34]  ( .D(N18), .CK(clk), .Q(data_out[34]) );
  DFF_X1 \data_out_reg[33]  ( .D(N19), .CK(clk), .Q(data_out[33]) );
  DFF_X1 \data_out_reg[32]  ( .D(N20), .CK(clk), .Q(data_out[32]) );
  DFF_X1 \data_out_reg[31]  ( .D(N21), .CK(clk), .Q(data_out[31]) );
  DFF_X1 \data_out_reg[30]  ( .D(N22), .CK(clk), .Q(data_out[30]) );
  DFF_X1 \data_out_reg[29]  ( .D(N23), .CK(clk), .Q(data_out[29]) );
  DFF_X1 \data_out_reg[28]  ( .D(N24), .CK(clk), .Q(data_out[28]) );
  DFF_X1 \data_out_reg[27]  ( .D(N25), .CK(clk), .Q(data_out[27]) );
  DFF_X1 \data_out_reg[26]  ( .D(N26), .CK(clk), .Q(data_out[26]) );
  DFF_X1 \data_out_reg[25]  ( .D(N27), .CK(clk), .Q(data_out[25]) );
  DFF_X1 \data_out_reg[24]  ( .D(N28), .CK(clk), .Q(data_out[24]) );
  DFF_X1 \data_out_reg[23]  ( .D(N29), .CK(clk), .Q(data_out[23]) );
  DFF_X1 \data_out_reg[22]  ( .D(N30), .CK(clk), .Q(data_out[22]) );
  DFF_X1 \data_out_reg[21]  ( .D(N31), .CK(clk), .Q(data_out[21]) );
  DFF_X1 \data_out_reg[20]  ( .D(N32), .CK(clk), .Q(data_out[20]) );
  DFF_X1 \data_out_reg[19]  ( .D(N33), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \data_out_reg[18]  ( .D(N34), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[17]  ( .D(N35), .CK(clk), .Q(data_out[17]) );
  DFF_X1 \data_out_reg[16]  ( .D(N36), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[15]  ( .D(N37), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N38), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(N39), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(N40), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(N41), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N42), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N43), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N44), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N45), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N46), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N47), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N48), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N49), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N50), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N51), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N52), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][39]  ( .D(n693), .CK(clk), .Q(\mem[7][39] ) );
  DFF_X1 \mem_reg[7][38]  ( .D(n692), .CK(clk), .Q(\mem[7][38] ) );
  DFF_X1 \mem_reg[7][37]  ( .D(n691), .CK(clk), .Q(\mem[7][37] ) );
  DFF_X1 \mem_reg[7][36]  ( .D(n690), .CK(clk), .Q(\mem[7][36] ) );
  DFF_X1 \mem_reg[7][35]  ( .D(n689), .CK(clk), .Q(\mem[7][35] ) );
  DFF_X1 \mem_reg[7][34]  ( .D(n688), .CK(clk), .Q(\mem[7][34] ) );
  DFF_X1 \mem_reg[7][33]  ( .D(n687), .CK(clk), .Q(\mem[7][33] ) );
  DFF_X1 \mem_reg[7][32]  ( .D(n686), .CK(clk), .Q(\mem[7][32] ) );
  DFF_X1 \mem_reg[7][31]  ( .D(n685), .CK(clk), .Q(\mem[7][31] ) );
  DFF_X1 \mem_reg[7][30]  ( .D(n684), .CK(clk), .Q(\mem[7][30] ) );
  DFF_X1 \mem_reg[7][29]  ( .D(n683), .CK(clk), .Q(\mem[7][29] ) );
  DFF_X1 \mem_reg[7][28]  ( .D(n682), .CK(clk), .Q(\mem[7][28] ) );
  DFF_X1 \mem_reg[7][27]  ( .D(n681), .CK(clk), .Q(\mem[7][27] ) );
  DFF_X1 \mem_reg[7][26]  ( .D(n680), .CK(clk), .Q(\mem[7][26] ) );
  DFF_X1 \mem_reg[7][25]  ( .D(n679), .CK(clk), .Q(\mem[7][25] ) );
  DFF_X1 \mem_reg[7][24]  ( .D(n678), .CK(clk), .Q(\mem[7][24] ) );
  DFF_X1 \mem_reg[7][23]  ( .D(n677), .CK(clk), .Q(\mem[7][23] ) );
  DFF_X1 \mem_reg[7][22]  ( .D(n676), .CK(clk), .Q(\mem[7][22] ) );
  DFF_X1 \mem_reg[7][21]  ( .D(n675), .CK(clk), .Q(\mem[7][21] ) );
  DFF_X1 \mem_reg[7][20]  ( .D(n674), .CK(clk), .Q(\mem[7][20] ) );
  DFF_X1 \mem_reg[7][19]  ( .D(n673), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n672), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n671), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n670), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n669), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n668), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n667), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n666), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n665), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n664), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n663), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n662), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n661), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n660), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n659), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n658), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n657), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n656), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n655), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n654), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][39]  ( .D(n653), .CK(clk), .Q(\mem[6][39] ) );
  DFF_X1 \mem_reg[6][38]  ( .D(n652), .CK(clk), .Q(\mem[6][38] ) );
  DFF_X1 \mem_reg[6][37]  ( .D(n651), .CK(clk), .Q(\mem[6][37] ) );
  DFF_X1 \mem_reg[6][36]  ( .D(n650), .CK(clk), .Q(\mem[6][36] ) );
  DFF_X1 \mem_reg[6][35]  ( .D(n649), .CK(clk), .Q(\mem[6][35] ) );
  DFF_X1 \mem_reg[6][34]  ( .D(n648), .CK(clk), .Q(\mem[6][34] ) );
  DFF_X1 \mem_reg[6][33]  ( .D(n647), .CK(clk), .Q(\mem[6][33] ) );
  DFF_X1 \mem_reg[6][32]  ( .D(n646), .CK(clk), .Q(\mem[6][32] ) );
  DFF_X1 \mem_reg[6][31]  ( .D(n645), .CK(clk), .Q(\mem[6][31] ) );
  DFF_X1 \mem_reg[6][30]  ( .D(n644), .CK(clk), .Q(\mem[6][30] ) );
  DFF_X1 \mem_reg[6][29]  ( .D(n643), .CK(clk), .Q(\mem[6][29] ) );
  DFF_X1 \mem_reg[6][28]  ( .D(n642), .CK(clk), .Q(\mem[6][28] ) );
  DFF_X1 \mem_reg[6][27]  ( .D(n641), .CK(clk), .Q(\mem[6][27] ) );
  DFF_X1 \mem_reg[6][26]  ( .D(n640), .CK(clk), .Q(\mem[6][26] ) );
  DFF_X1 \mem_reg[6][25]  ( .D(n639), .CK(clk), .Q(\mem[6][25] ) );
  DFF_X1 \mem_reg[6][24]  ( .D(n638), .CK(clk), .Q(\mem[6][24] ) );
  DFF_X1 \mem_reg[6][23]  ( .D(n637), .CK(clk), .Q(\mem[6][23] ) );
  DFF_X1 \mem_reg[6][22]  ( .D(n636), .CK(clk), .Q(\mem[6][22] ) );
  DFF_X1 \mem_reg[6][21]  ( .D(n635), .CK(clk), .Q(\mem[6][21] ) );
  DFF_X1 \mem_reg[6][20]  ( .D(n634), .CK(clk), .Q(\mem[6][20] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n633), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n632), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n631), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n630), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n629), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n628), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n627), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n626), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n625), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n624), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n623), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n622), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n621), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n620), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n619), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n618), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n617), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n616), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n615), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n614), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][39]  ( .D(n613), .CK(clk), .Q(\mem[5][39] ) );
  DFF_X1 \mem_reg[5][38]  ( .D(n612), .CK(clk), .Q(\mem[5][38] ) );
  DFF_X1 \mem_reg[5][37]  ( .D(n611), .CK(clk), .Q(\mem[5][37] ) );
  DFF_X1 \mem_reg[5][36]  ( .D(n610), .CK(clk), .Q(\mem[5][36] ) );
  DFF_X1 \mem_reg[5][35]  ( .D(n609), .CK(clk), .Q(\mem[5][35] ) );
  DFF_X1 \mem_reg[5][34]  ( .D(n608), .CK(clk), .Q(\mem[5][34] ) );
  DFF_X1 \mem_reg[5][33]  ( .D(n607), .CK(clk), .Q(\mem[5][33] ) );
  DFF_X1 \mem_reg[5][32]  ( .D(n606), .CK(clk), .Q(\mem[5][32] ) );
  DFF_X1 \mem_reg[5][31]  ( .D(n605), .CK(clk), .Q(\mem[5][31] ) );
  DFF_X1 \mem_reg[5][30]  ( .D(n604), .CK(clk), .Q(\mem[5][30] ) );
  DFF_X1 \mem_reg[5][29]  ( .D(n603), .CK(clk), .Q(\mem[5][29] ) );
  DFF_X1 \mem_reg[5][28]  ( .D(n602), .CK(clk), .Q(\mem[5][28] ) );
  DFF_X1 \mem_reg[5][27]  ( .D(n601), .CK(clk), .Q(\mem[5][27] ) );
  DFF_X1 \mem_reg[5][26]  ( .D(n600), .CK(clk), .Q(\mem[5][26] ) );
  DFF_X1 \mem_reg[5][25]  ( .D(n599), .CK(clk), .Q(\mem[5][25] ) );
  DFF_X1 \mem_reg[5][24]  ( .D(n598), .CK(clk), .Q(\mem[5][24] ) );
  DFF_X1 \mem_reg[5][23]  ( .D(n597), .CK(clk), .Q(\mem[5][23] ) );
  DFF_X1 \mem_reg[5][22]  ( .D(n596), .CK(clk), .Q(\mem[5][22] ) );
  DFF_X1 \mem_reg[5][21]  ( .D(n595), .CK(clk), .Q(\mem[5][21] ) );
  DFF_X1 \mem_reg[5][20]  ( .D(n594), .CK(clk), .Q(\mem[5][20] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n593), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n592), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n591), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n590), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n589), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n588), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n587), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n586), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n585), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n584), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n583), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n582), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n581), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n580), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n579), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n578), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n577), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n576), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n575), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n574), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][39]  ( .D(n573), .CK(clk), .Q(\mem[4][39] ) );
  DFF_X1 \mem_reg[4][38]  ( .D(n572), .CK(clk), .Q(\mem[4][38] ) );
  DFF_X1 \mem_reg[4][37]  ( .D(n571), .CK(clk), .Q(\mem[4][37] ) );
  DFF_X1 \mem_reg[4][36]  ( .D(n570), .CK(clk), .Q(\mem[4][36] ) );
  DFF_X1 \mem_reg[4][35]  ( .D(n569), .CK(clk), .Q(\mem[4][35] ) );
  DFF_X1 \mem_reg[4][34]  ( .D(n568), .CK(clk), .Q(\mem[4][34] ) );
  DFF_X1 \mem_reg[4][33]  ( .D(n567), .CK(clk), .Q(\mem[4][33] ) );
  DFF_X1 \mem_reg[4][32]  ( .D(n566), .CK(clk), .Q(\mem[4][32] ) );
  DFF_X1 \mem_reg[4][31]  ( .D(n565), .CK(clk), .Q(\mem[4][31] ) );
  DFF_X1 \mem_reg[4][30]  ( .D(n564), .CK(clk), .Q(\mem[4][30] ) );
  DFF_X1 \mem_reg[4][29]  ( .D(n563), .CK(clk), .Q(\mem[4][29] ) );
  DFF_X1 \mem_reg[4][28]  ( .D(n562), .CK(clk), .Q(\mem[4][28] ) );
  DFF_X1 \mem_reg[4][27]  ( .D(n561), .CK(clk), .Q(\mem[4][27] ) );
  DFF_X1 \mem_reg[4][26]  ( .D(n560), .CK(clk), .Q(\mem[4][26] ) );
  DFF_X1 \mem_reg[4][25]  ( .D(n559), .CK(clk), .Q(\mem[4][25] ) );
  DFF_X1 \mem_reg[4][24]  ( .D(n558), .CK(clk), .Q(\mem[4][24] ) );
  DFF_X1 \mem_reg[4][23]  ( .D(n557), .CK(clk), .Q(\mem[4][23] ) );
  DFF_X1 \mem_reg[4][22]  ( .D(n556), .CK(clk), .Q(\mem[4][22] ) );
  DFF_X1 \mem_reg[4][21]  ( .D(n555), .CK(clk), .Q(\mem[4][21] ) );
  DFF_X1 \mem_reg[4][20]  ( .D(n554), .CK(clk), .Q(\mem[4][20] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n553), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n552), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n551), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n550), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n549), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n548), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n547), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n546), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n545), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n544), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n543), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n542), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n541), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n540), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n539), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n538), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n537), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n536), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n535), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n534), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][39]  ( .D(n533), .CK(clk), .Q(\mem[3][39] ) );
  DFF_X1 \mem_reg[3][38]  ( .D(n532), .CK(clk), .Q(\mem[3][38] ) );
  DFF_X1 \mem_reg[3][37]  ( .D(n531), .CK(clk), .Q(\mem[3][37] ) );
  DFF_X1 \mem_reg[3][36]  ( .D(n530), .CK(clk), .Q(\mem[3][36] ) );
  DFF_X1 \mem_reg[3][35]  ( .D(n529), .CK(clk), .Q(\mem[3][35] ) );
  DFF_X1 \mem_reg[3][34]  ( .D(n528), .CK(clk), .Q(\mem[3][34] ) );
  DFF_X1 \mem_reg[3][33]  ( .D(n527), .CK(clk), .Q(\mem[3][33] ) );
  DFF_X1 \mem_reg[3][32]  ( .D(n526), .CK(clk), .Q(\mem[3][32] ) );
  DFF_X1 \mem_reg[3][31]  ( .D(n525), .CK(clk), .Q(\mem[3][31] ) );
  DFF_X1 \mem_reg[3][30]  ( .D(n524), .CK(clk), .Q(\mem[3][30] ) );
  DFF_X1 \mem_reg[3][29]  ( .D(n523), .CK(clk), .Q(\mem[3][29] ) );
  DFF_X1 \mem_reg[3][28]  ( .D(n522), .CK(clk), .Q(\mem[3][28] ) );
  DFF_X1 \mem_reg[3][27]  ( .D(n521), .CK(clk), .Q(\mem[3][27] ) );
  DFF_X1 \mem_reg[3][26]  ( .D(n520), .CK(clk), .Q(\mem[3][26] ) );
  DFF_X1 \mem_reg[3][25]  ( .D(n519), .CK(clk), .Q(\mem[3][25] ) );
  DFF_X1 \mem_reg[3][24]  ( .D(n518), .CK(clk), .Q(\mem[3][24] ) );
  DFF_X1 \mem_reg[3][23]  ( .D(n517), .CK(clk), .Q(\mem[3][23] ) );
  DFF_X1 \mem_reg[3][22]  ( .D(n516), .CK(clk), .Q(\mem[3][22] ) );
  DFF_X1 \mem_reg[3][21]  ( .D(n515), .CK(clk), .Q(\mem[3][21] ) );
  DFF_X1 \mem_reg[3][20]  ( .D(n514), .CK(clk), .Q(\mem[3][20] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n513), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n512), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n511), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n510), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n509), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n508), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n507), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n506), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n505), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n504), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n503), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n502), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n501), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n500), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n499), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n498), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n497), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n496), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n495), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n494), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][39]  ( .D(n493), .CK(clk), .Q(\mem[2][39] ) );
  DFF_X1 \mem_reg[2][38]  ( .D(n492), .CK(clk), .Q(\mem[2][38] ) );
  DFF_X1 \mem_reg[2][37]  ( .D(n491), .CK(clk), .Q(\mem[2][37] ) );
  DFF_X1 \mem_reg[2][36]  ( .D(n490), .CK(clk), .Q(\mem[2][36] ) );
  DFF_X1 \mem_reg[2][35]  ( .D(n489), .CK(clk), .Q(\mem[2][35] ) );
  DFF_X1 \mem_reg[2][34]  ( .D(n488), .CK(clk), .Q(\mem[2][34] ) );
  DFF_X1 \mem_reg[2][33]  ( .D(n487), .CK(clk), .Q(\mem[2][33] ) );
  DFF_X1 \mem_reg[2][32]  ( .D(n486), .CK(clk), .Q(\mem[2][32] ) );
  DFF_X1 \mem_reg[2][31]  ( .D(n485), .CK(clk), .Q(\mem[2][31] ) );
  DFF_X1 \mem_reg[2][30]  ( .D(n484), .CK(clk), .Q(\mem[2][30] ) );
  DFF_X1 \mem_reg[2][29]  ( .D(n483), .CK(clk), .Q(\mem[2][29] ) );
  DFF_X1 \mem_reg[2][28]  ( .D(n482), .CK(clk), .Q(\mem[2][28] ) );
  DFF_X1 \mem_reg[2][27]  ( .D(n481), .CK(clk), .Q(\mem[2][27] ) );
  DFF_X1 \mem_reg[2][26]  ( .D(n480), .CK(clk), .Q(\mem[2][26] ) );
  DFF_X1 \mem_reg[2][25]  ( .D(n479), .CK(clk), .Q(\mem[2][25] ) );
  DFF_X1 \mem_reg[2][24]  ( .D(n478), .CK(clk), .Q(\mem[2][24] ) );
  DFF_X1 \mem_reg[2][23]  ( .D(n477), .CK(clk), .Q(\mem[2][23] ) );
  DFF_X1 \mem_reg[2][22]  ( .D(n476), .CK(clk), .Q(\mem[2][22] ) );
  DFF_X1 \mem_reg[2][21]  ( .D(n475), .CK(clk), .Q(\mem[2][21] ) );
  DFF_X1 \mem_reg[2][20]  ( .D(n474), .CK(clk), .Q(\mem[2][20] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n473), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n472), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n471), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n470), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n469), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n468), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n467), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n466), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n465), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n464), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n463), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n462), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n461), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n460), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n459), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n458), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n457), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n456), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n455), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n454), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][39]  ( .D(n453), .CK(clk), .Q(\mem[1][39] ) );
  DFF_X1 \mem_reg[1][38]  ( .D(n452), .CK(clk), .Q(\mem[1][38] ) );
  DFF_X1 \mem_reg[1][37]  ( .D(n451), .CK(clk), .Q(\mem[1][37] ) );
  DFF_X1 \mem_reg[1][36]  ( .D(n450), .CK(clk), .Q(\mem[1][36] ) );
  DFF_X1 \mem_reg[1][35]  ( .D(n449), .CK(clk), .Q(\mem[1][35] ) );
  DFF_X1 \mem_reg[1][34]  ( .D(n448), .CK(clk), .Q(\mem[1][34] ) );
  DFF_X1 \mem_reg[1][33]  ( .D(n447), .CK(clk), .Q(\mem[1][33] ) );
  DFF_X1 \mem_reg[1][32]  ( .D(n446), .CK(clk), .Q(\mem[1][32] ) );
  DFF_X1 \mem_reg[1][31]  ( .D(n445), .CK(clk), .Q(\mem[1][31] ) );
  DFF_X1 \mem_reg[1][30]  ( .D(n444), .CK(clk), .Q(\mem[1][30] ) );
  DFF_X1 \mem_reg[1][29]  ( .D(n443), .CK(clk), .Q(\mem[1][29] ) );
  DFF_X1 \mem_reg[1][28]  ( .D(n442), .CK(clk), .Q(\mem[1][28] ) );
  DFF_X1 \mem_reg[1][27]  ( .D(n441), .CK(clk), .Q(\mem[1][27] ) );
  DFF_X1 \mem_reg[1][26]  ( .D(n440), .CK(clk), .Q(\mem[1][26] ) );
  DFF_X1 \mem_reg[1][25]  ( .D(n439), .CK(clk), .Q(\mem[1][25] ) );
  DFF_X1 \mem_reg[1][24]  ( .D(n438), .CK(clk), .Q(\mem[1][24] ) );
  DFF_X1 \mem_reg[1][23]  ( .D(n437), .CK(clk), .Q(\mem[1][23] ) );
  DFF_X1 \mem_reg[1][22]  ( .D(n436), .CK(clk), .Q(\mem[1][22] ) );
  DFF_X1 \mem_reg[1][21]  ( .D(n435), .CK(clk), .Q(\mem[1][21] ) );
  DFF_X1 \mem_reg[1][20]  ( .D(n434), .CK(clk), .Q(\mem[1][20] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n433), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n432), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n431), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n430), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n429), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n428), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n427), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n426), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n425), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n424), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n423), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n422), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n421), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n420), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n419), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n418), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n417), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n416), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n415), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n414), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][39]  ( .D(n413), .CK(clk), .Q(\mem[0][39] ) );
  DFF_X1 \mem_reg[0][38]  ( .D(n412), .CK(clk), .Q(\mem[0][38] ) );
  DFF_X1 \mem_reg[0][37]  ( .D(n411), .CK(clk), .Q(\mem[0][37] ) );
  DFF_X1 \mem_reg[0][36]  ( .D(n410), .CK(clk), .Q(\mem[0][36] ) );
  DFF_X1 \mem_reg[0][35]  ( .D(n409), .CK(clk), .Q(\mem[0][35] ) );
  DFF_X1 \mem_reg[0][34]  ( .D(n408), .CK(clk), .Q(\mem[0][34] ) );
  DFF_X1 \mem_reg[0][33]  ( .D(n407), .CK(clk), .Q(\mem[0][33] ) );
  DFF_X1 \mem_reg[0][32]  ( .D(n406), .CK(clk), .Q(\mem[0][32] ) );
  DFF_X1 \mem_reg[0][31]  ( .D(n405), .CK(clk), .Q(\mem[0][31] ) );
  DFF_X1 \mem_reg[0][30]  ( .D(n404), .CK(clk), .Q(\mem[0][30] ) );
  DFF_X1 \mem_reg[0][29]  ( .D(n403), .CK(clk), .Q(\mem[0][29] ) );
  DFF_X1 \mem_reg[0][28]  ( .D(n402), .CK(clk), .Q(\mem[0][28] ) );
  DFF_X1 \mem_reg[0][27]  ( .D(n401), .CK(clk), .Q(\mem[0][27] ) );
  DFF_X1 \mem_reg[0][26]  ( .D(n400), .CK(clk), .Q(\mem[0][26] ) );
  DFF_X1 \mem_reg[0][25]  ( .D(n399), .CK(clk), .Q(\mem[0][25] ) );
  DFF_X1 \mem_reg[0][24]  ( .D(n398), .CK(clk), .Q(\mem[0][24] ) );
  DFF_X1 \mem_reg[0][23]  ( .D(n397), .CK(clk), .Q(\mem[0][23] ) );
  DFF_X1 \mem_reg[0][22]  ( .D(n396), .CK(clk), .Q(\mem[0][22] ) );
  DFF_X1 \mem_reg[0][21]  ( .D(n395), .CK(clk), .Q(\mem[0][21] ) );
  DFF_X1 \mem_reg[0][20]  ( .D(n394), .CK(clk), .Q(\mem[0][20] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n393), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n392), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n391), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n390), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n389), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n388), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n387), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n386), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n385), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n384), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n383), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n382), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n381), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n380), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n379), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n378), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n377), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n376), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n375), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n374), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U688 ( .A1(n926), .A2(n927), .A3(n85), .ZN(n44) );
  NAND3_X1 U689 ( .A1(n85), .A2(n927), .A3(N10), .ZN(n86) );
  NAND3_X1 U690 ( .A1(n85), .A2(n926), .A3(N11), .ZN(n127) );
  NAND3_X1 U691 ( .A1(N10), .A2(n85), .A3(N11), .ZN(n168) );
  NAND3_X1 U692 ( .A1(n926), .A2(n927), .A3(n250), .ZN(n209) );
  NAND3_X1 U693 ( .A1(N10), .A2(n927), .A3(n250), .ZN(n251) );
  NAND3_X1 U694 ( .A1(N11), .A2(n926), .A3(n250), .ZN(n292) );
  NAND3_X1 U695 ( .A1(N11), .A2(N10), .A3(n250), .ZN(n333) );
  BUF_X1 U3 ( .A(n901), .Z(n898) );
  BUF_X1 U4 ( .A(n901), .Z(n899) );
  BUF_X1 U5 ( .A(n901), .Z(n897) );
  BUF_X1 U6 ( .A(n900), .Z(n896) );
  BUF_X1 U7 ( .A(N10), .Z(n901) );
  BUF_X1 U8 ( .A(N10), .Z(n900) );
  BUF_X1 U9 ( .A(N11), .Z(n892) );
  BUF_X1 U10 ( .A(N11), .Z(n893) );
  BUF_X1 U11 ( .A(N11), .Z(n894) );
  BUF_X1 U12 ( .A(n44), .Z(n925) );
  BUF_X1 U13 ( .A(n44), .Z(n924) );
  BUF_X1 U14 ( .A(n44), .Z(n923) );
  BUF_X1 U15 ( .A(n86), .Z(n922) );
  BUF_X1 U16 ( .A(n86), .Z(n921) );
  BUF_X1 U17 ( .A(n86), .Z(n920) );
  BUF_X1 U18 ( .A(n168), .Z(n915) );
  BUF_X1 U19 ( .A(n168), .Z(n914) );
  BUF_X1 U20 ( .A(n209), .Z(n913) );
  BUF_X1 U21 ( .A(n209), .Z(n912) );
  BUF_X1 U22 ( .A(n209), .Z(n911) );
  BUF_X1 U23 ( .A(n251), .Z(n910) );
  BUF_X1 U24 ( .A(n251), .Z(n909) );
  BUF_X1 U25 ( .A(n251), .Z(n908) );
  BUF_X1 U26 ( .A(n292), .Z(n907) );
  BUF_X1 U27 ( .A(n292), .Z(n906) );
  BUF_X1 U28 ( .A(n292), .Z(n905) );
  BUF_X1 U29 ( .A(n333), .Z(n902) );
  BUF_X1 U30 ( .A(n168), .Z(n916) );
  BUF_X1 U31 ( .A(n127), .Z(n917) );
  BUF_X1 U32 ( .A(n127), .Z(n918) );
  BUF_X1 U33 ( .A(n333), .Z(n903) );
  INV_X1 U34 ( .A(N10), .ZN(n926) );
  INV_X1 U35 ( .A(N11), .ZN(n927) );
  BUF_X1 U36 ( .A(N12), .Z(n891) );
  NOR2_X1 U37 ( .A1(n928), .A2(N12), .ZN(n85) );
  INV_X1 U38 ( .A(wr_en), .ZN(n928) );
  AND2_X1 U39 ( .A1(N12), .A2(wr_en), .ZN(n250) );
  OAI21_X1 U40 ( .B1(n937), .B2(n906), .A(n324), .ZN(n645) );
  NAND2_X1 U41 ( .A1(\mem[6][31] ), .A2(n906), .ZN(n324) );
  OAI21_X1 U42 ( .B1(n936), .B2(n907), .A(n325), .ZN(n646) );
  NAND2_X1 U43 ( .A1(\mem[6][32] ), .A2(n905), .ZN(n325) );
  OAI21_X1 U44 ( .B1(n935), .B2(n906), .A(n326), .ZN(n647) );
  NAND2_X1 U45 ( .A1(\mem[6][33] ), .A2(n905), .ZN(n326) );
  OAI21_X1 U46 ( .B1(n934), .B2(n905), .A(n327), .ZN(n648) );
  NAND2_X1 U47 ( .A1(\mem[6][34] ), .A2(n905), .ZN(n327) );
  OAI21_X1 U48 ( .B1(n933), .B2(n292), .A(n328), .ZN(n649) );
  NAND2_X1 U49 ( .A1(\mem[6][35] ), .A2(n905), .ZN(n328) );
  OAI21_X1 U50 ( .B1(n932), .B2(n292), .A(n329), .ZN(n650) );
  NAND2_X1 U51 ( .A1(\mem[6][36] ), .A2(n905), .ZN(n329) );
  OAI21_X1 U52 ( .B1(n931), .B2(n292), .A(n330), .ZN(n651) );
  NAND2_X1 U53 ( .A1(\mem[6][37] ), .A2(n905), .ZN(n330) );
  OAI21_X1 U54 ( .B1(n930), .B2(n292), .A(n331), .ZN(n652) );
  NAND2_X1 U55 ( .A1(\mem[6][38] ), .A2(n905), .ZN(n331) );
  OAI21_X1 U56 ( .B1(n937), .B2(n904), .A(n365), .ZN(n685) );
  NAND2_X1 U57 ( .A1(\mem[7][31] ), .A2(n902), .ZN(n365) );
  OAI21_X1 U58 ( .B1(n936), .B2(n904), .A(n366), .ZN(n686) );
  NAND2_X1 U59 ( .A1(\mem[7][32] ), .A2(n333), .ZN(n366) );
  OAI21_X1 U60 ( .B1(n935), .B2(n904), .A(n367), .ZN(n687) );
  NAND2_X1 U61 ( .A1(\mem[7][33] ), .A2(n333), .ZN(n367) );
  OAI21_X1 U62 ( .B1(n934), .B2(n904), .A(n368), .ZN(n688) );
  NAND2_X1 U63 ( .A1(\mem[7][34] ), .A2(n333), .ZN(n368) );
  OAI21_X1 U64 ( .B1(n933), .B2(n904), .A(n369), .ZN(n689) );
  NAND2_X1 U65 ( .A1(\mem[7][35] ), .A2(n333), .ZN(n369) );
  OAI21_X1 U66 ( .B1(n932), .B2(n904), .A(n370), .ZN(n690) );
  NAND2_X1 U67 ( .A1(\mem[7][36] ), .A2(n333), .ZN(n370) );
  OAI21_X1 U68 ( .B1(n931), .B2(n904), .A(n371), .ZN(n691) );
  NAND2_X1 U69 ( .A1(\mem[7][37] ), .A2(n333), .ZN(n371) );
  OAI21_X1 U70 ( .B1(n930), .B2(n904), .A(n372), .ZN(n692) );
  NAND2_X1 U71 ( .A1(\mem[7][38] ), .A2(n333), .ZN(n372) );
  OAI21_X1 U72 ( .B1(n937), .B2(n86), .A(n118), .ZN(n445) );
  NAND2_X1 U73 ( .A1(\mem[1][31] ), .A2(n921), .ZN(n118) );
  OAI21_X1 U74 ( .B1(n936), .B2(n86), .A(n119), .ZN(n446) );
  NAND2_X1 U75 ( .A1(\mem[1][32] ), .A2(n920), .ZN(n119) );
  OAI21_X1 U76 ( .B1(n935), .B2(n86), .A(n120), .ZN(n447) );
  NAND2_X1 U77 ( .A1(\mem[1][33] ), .A2(n920), .ZN(n120) );
  OAI21_X1 U78 ( .B1(n934), .B2(n86), .A(n121), .ZN(n448) );
  NAND2_X1 U79 ( .A1(\mem[1][34] ), .A2(n920), .ZN(n121) );
  OAI21_X1 U80 ( .B1(n933), .B2(n86), .A(n122), .ZN(n449) );
  NAND2_X1 U81 ( .A1(\mem[1][35] ), .A2(n920), .ZN(n122) );
  OAI21_X1 U82 ( .B1(n932), .B2(n86), .A(n123), .ZN(n450) );
  NAND2_X1 U83 ( .A1(\mem[1][36] ), .A2(n920), .ZN(n123) );
  OAI21_X1 U84 ( .B1(n931), .B2(n921), .A(n124), .ZN(n451) );
  NAND2_X1 U85 ( .A1(\mem[1][37] ), .A2(n920), .ZN(n124) );
  OAI21_X1 U86 ( .B1(n930), .B2(n86), .A(n125), .ZN(n452) );
  NAND2_X1 U87 ( .A1(\mem[1][38] ), .A2(n920), .ZN(n125) );
  OAI21_X1 U88 ( .B1(n937), .B2(n919), .A(n159), .ZN(n485) );
  NAND2_X1 U89 ( .A1(\mem[2][31] ), .A2(n127), .ZN(n159) );
  OAI21_X1 U90 ( .B1(n936), .B2(n919), .A(n160), .ZN(n486) );
  NAND2_X1 U91 ( .A1(\mem[2][32] ), .A2(n127), .ZN(n160) );
  OAI21_X1 U92 ( .B1(n935), .B2(n919), .A(n161), .ZN(n487) );
  NAND2_X1 U93 ( .A1(\mem[2][33] ), .A2(n127), .ZN(n161) );
  OAI21_X1 U94 ( .B1(n934), .B2(n919), .A(n162), .ZN(n488) );
  NAND2_X1 U95 ( .A1(\mem[2][34] ), .A2(n127), .ZN(n162) );
  OAI21_X1 U96 ( .B1(n933), .B2(n919), .A(n163), .ZN(n489) );
  NAND2_X1 U97 ( .A1(\mem[2][35] ), .A2(n127), .ZN(n163) );
  OAI21_X1 U98 ( .B1(n932), .B2(n919), .A(n164), .ZN(n490) );
  NAND2_X1 U99 ( .A1(\mem[2][36] ), .A2(n127), .ZN(n164) );
  OAI21_X1 U100 ( .B1(n931), .B2(n919), .A(n165), .ZN(n491) );
  NAND2_X1 U101 ( .A1(\mem[2][37] ), .A2(n127), .ZN(n165) );
  OAI21_X1 U102 ( .B1(n930), .B2(n919), .A(n166), .ZN(n492) );
  NAND2_X1 U103 ( .A1(\mem[2][38] ), .A2(n127), .ZN(n166) );
  OAI21_X1 U104 ( .B1(n937), .B2(n915), .A(n200), .ZN(n525) );
  NAND2_X1 U105 ( .A1(\mem[3][31] ), .A2(n915), .ZN(n200) );
  OAI21_X1 U106 ( .B1(n936), .B2(n916), .A(n201), .ZN(n526) );
  NAND2_X1 U107 ( .A1(\mem[3][32] ), .A2(n914), .ZN(n201) );
  OAI21_X1 U108 ( .B1(n935), .B2(n916), .A(n202), .ZN(n527) );
  NAND2_X1 U109 ( .A1(\mem[3][33] ), .A2(n914), .ZN(n202) );
  OAI21_X1 U110 ( .B1(n934), .B2(n915), .A(n203), .ZN(n528) );
  NAND2_X1 U111 ( .A1(\mem[3][34] ), .A2(n914), .ZN(n203) );
  OAI21_X1 U112 ( .B1(n933), .B2(n914), .A(n204), .ZN(n529) );
  NAND2_X1 U113 ( .A1(\mem[3][35] ), .A2(n914), .ZN(n204) );
  OAI21_X1 U114 ( .B1(n932), .B2(n914), .A(n205), .ZN(n530) );
  NAND2_X1 U115 ( .A1(\mem[3][36] ), .A2(n914), .ZN(n205) );
  OAI21_X1 U116 ( .B1(n931), .B2(n915), .A(n206), .ZN(n531) );
  NAND2_X1 U117 ( .A1(\mem[3][37] ), .A2(n914), .ZN(n206) );
  OAI21_X1 U118 ( .B1(n930), .B2(n916), .A(n207), .ZN(n532) );
  NAND2_X1 U119 ( .A1(\mem[3][38] ), .A2(n914), .ZN(n207) );
  OAI21_X1 U120 ( .B1(n937), .B2(n209), .A(n241), .ZN(n565) );
  NAND2_X1 U121 ( .A1(\mem[4][31] ), .A2(n912), .ZN(n241) );
  OAI21_X1 U122 ( .B1(n936), .B2(n209), .A(n242), .ZN(n566) );
  NAND2_X1 U123 ( .A1(\mem[4][32] ), .A2(n911), .ZN(n242) );
  OAI21_X1 U124 ( .B1(n935), .B2(n209), .A(n243), .ZN(n567) );
  NAND2_X1 U125 ( .A1(\mem[4][33] ), .A2(n911), .ZN(n243) );
  OAI21_X1 U126 ( .B1(n934), .B2(n209), .A(n244), .ZN(n568) );
  NAND2_X1 U127 ( .A1(\mem[4][34] ), .A2(n911), .ZN(n244) );
  OAI21_X1 U128 ( .B1(n933), .B2(n209), .A(n245), .ZN(n569) );
  NAND2_X1 U129 ( .A1(\mem[4][35] ), .A2(n911), .ZN(n245) );
  OAI21_X1 U130 ( .B1(n932), .B2(n209), .A(n246), .ZN(n570) );
  NAND2_X1 U131 ( .A1(\mem[4][36] ), .A2(n911), .ZN(n246) );
  OAI21_X1 U132 ( .B1(n931), .B2(n912), .A(n247), .ZN(n571) );
  NAND2_X1 U133 ( .A1(\mem[4][37] ), .A2(n911), .ZN(n247) );
  OAI21_X1 U134 ( .B1(n930), .B2(n209), .A(n248), .ZN(n572) );
  NAND2_X1 U135 ( .A1(\mem[4][38] ), .A2(n911), .ZN(n248) );
  OAI21_X1 U136 ( .B1(n937), .B2(n909), .A(n283), .ZN(n605) );
  NAND2_X1 U137 ( .A1(\mem[5][31] ), .A2(n909), .ZN(n283) );
  OAI21_X1 U138 ( .B1(n936), .B2(n910), .A(n284), .ZN(n606) );
  NAND2_X1 U139 ( .A1(\mem[5][32] ), .A2(n908), .ZN(n284) );
  OAI21_X1 U140 ( .B1(n935), .B2(n909), .A(n285), .ZN(n607) );
  NAND2_X1 U141 ( .A1(\mem[5][33] ), .A2(n908), .ZN(n285) );
  OAI21_X1 U142 ( .B1(n934), .B2(n908), .A(n286), .ZN(n608) );
  NAND2_X1 U143 ( .A1(\mem[5][34] ), .A2(n908), .ZN(n286) );
  OAI21_X1 U144 ( .B1(n933), .B2(n251), .A(n287), .ZN(n609) );
  NAND2_X1 U145 ( .A1(\mem[5][35] ), .A2(n908), .ZN(n287) );
  OAI21_X1 U146 ( .B1(n932), .B2(n251), .A(n288), .ZN(n610) );
  NAND2_X1 U147 ( .A1(\mem[5][36] ), .A2(n908), .ZN(n288) );
  OAI21_X1 U148 ( .B1(n931), .B2(n251), .A(n289), .ZN(n611) );
  NAND2_X1 U149 ( .A1(\mem[5][37] ), .A2(n908), .ZN(n289) );
  OAI21_X1 U150 ( .B1(n930), .B2(n251), .A(n290), .ZN(n612) );
  NAND2_X1 U151 ( .A1(\mem[5][38] ), .A2(n908), .ZN(n290) );
  OAI21_X1 U152 ( .B1(n925), .B2(n934), .A(n79), .ZN(n408) );
  NAND2_X1 U153 ( .A1(\mem[0][34] ), .A2(n924), .ZN(n79) );
  OAI21_X1 U154 ( .B1(n924), .B2(n933), .A(n80), .ZN(n409) );
  NAND2_X1 U155 ( .A1(\mem[0][35] ), .A2(n925), .ZN(n80) );
  OAI21_X1 U156 ( .B1(n923), .B2(n932), .A(n81), .ZN(n410) );
  NAND2_X1 U157 ( .A1(\mem[0][36] ), .A2(n923), .ZN(n81) );
  OAI21_X1 U158 ( .B1(n923), .B2(n931), .A(n82), .ZN(n411) );
  NAND2_X1 U159 ( .A1(\mem[0][37] ), .A2(n44), .ZN(n82) );
  OAI21_X1 U160 ( .B1(n44), .B2(n930), .A(n83), .ZN(n412) );
  NAND2_X1 U161 ( .A1(\mem[0][38] ), .A2(n925), .ZN(n83) );
  OAI21_X1 U162 ( .B1(n925), .B2(n967), .A(n46), .ZN(n375) );
  NAND2_X1 U163 ( .A1(\mem[0][1] ), .A2(n925), .ZN(n46) );
  OAI21_X1 U164 ( .B1(n925), .B2(n966), .A(n47), .ZN(n376) );
  NAND2_X1 U165 ( .A1(\mem[0][2] ), .A2(n923), .ZN(n47) );
  OAI21_X1 U166 ( .B1(n925), .B2(n965), .A(n48), .ZN(n377) );
  NAND2_X1 U167 ( .A1(\mem[0][3] ), .A2(n924), .ZN(n48) );
  OAI21_X1 U168 ( .B1(n925), .B2(n964), .A(n49), .ZN(n378) );
  NAND2_X1 U169 ( .A1(\mem[0][4] ), .A2(n923), .ZN(n49) );
  OAI21_X1 U170 ( .B1(n925), .B2(n963), .A(n50), .ZN(n379) );
  NAND2_X1 U171 ( .A1(\mem[0][5] ), .A2(n923), .ZN(n50) );
  OAI21_X1 U172 ( .B1(n925), .B2(n962), .A(n51), .ZN(n380) );
  NAND2_X1 U173 ( .A1(\mem[0][6] ), .A2(n923), .ZN(n51) );
  OAI21_X1 U174 ( .B1(n925), .B2(n960), .A(n53), .ZN(n382) );
  NAND2_X1 U175 ( .A1(\mem[0][8] ), .A2(n924), .ZN(n53) );
  OAI21_X1 U176 ( .B1(n925), .B2(n959), .A(n54), .ZN(n383) );
  NAND2_X1 U177 ( .A1(\mem[0][9] ), .A2(n924), .ZN(n54) );
  OAI21_X1 U178 ( .B1(n925), .B2(n929), .A(n84), .ZN(n413) );
  NAND2_X1 U179 ( .A1(\mem[0][39] ), .A2(n925), .ZN(n84) );
  OAI21_X1 U180 ( .B1(n967), .B2(n920), .A(n88), .ZN(n415) );
  NAND2_X1 U181 ( .A1(\mem[1][1] ), .A2(n920), .ZN(n88) );
  OAI21_X1 U182 ( .B1(n966), .B2(n921), .A(n89), .ZN(n416) );
  NAND2_X1 U183 ( .A1(\mem[1][2] ), .A2(n920), .ZN(n89) );
  OAI21_X1 U184 ( .B1(n965), .B2(n922), .A(n90), .ZN(n417) );
  NAND2_X1 U185 ( .A1(\mem[1][3] ), .A2(n920), .ZN(n90) );
  OAI21_X1 U186 ( .B1(n964), .B2(n920), .A(n91), .ZN(n418) );
  NAND2_X1 U187 ( .A1(\mem[1][4] ), .A2(n921), .ZN(n91) );
  OAI21_X1 U188 ( .B1(n963), .B2(n921), .A(n92), .ZN(n419) );
  NAND2_X1 U189 ( .A1(\mem[1][5] ), .A2(n921), .ZN(n92) );
  OAI21_X1 U190 ( .B1(n962), .B2(n922), .A(n93), .ZN(n420) );
  NAND2_X1 U191 ( .A1(\mem[1][6] ), .A2(n921), .ZN(n93) );
  OAI21_X1 U192 ( .B1(n960), .B2(n920), .A(n95), .ZN(n422) );
  NAND2_X1 U193 ( .A1(\mem[1][8] ), .A2(n922), .ZN(n95) );
  OAI21_X1 U194 ( .B1(n929), .B2(n921), .A(n126), .ZN(n453) );
  NAND2_X1 U195 ( .A1(\mem[1][39] ), .A2(n920), .ZN(n126) );
  OAI21_X1 U196 ( .B1(n967), .B2(n919), .A(n129), .ZN(n455) );
  NAND2_X1 U197 ( .A1(\mem[2][1] ), .A2(n919), .ZN(n129) );
  OAI21_X1 U198 ( .B1(n966), .B2(n919), .A(n130), .ZN(n456) );
  NAND2_X1 U199 ( .A1(\mem[2][2] ), .A2(n917), .ZN(n130) );
  OAI21_X1 U200 ( .B1(n965), .B2(n919), .A(n131), .ZN(n457) );
  NAND2_X1 U201 ( .A1(\mem[2][3] ), .A2(n917), .ZN(n131) );
  OAI21_X1 U202 ( .B1(n964), .B2(n919), .A(n132), .ZN(n458) );
  NAND2_X1 U203 ( .A1(\mem[2][4] ), .A2(n918), .ZN(n132) );
  OAI21_X1 U204 ( .B1(n963), .B2(n919), .A(n133), .ZN(n459) );
  NAND2_X1 U205 ( .A1(\mem[2][5] ), .A2(n917), .ZN(n133) );
  OAI21_X1 U206 ( .B1(n962), .B2(n917), .A(n134), .ZN(n460) );
  NAND2_X1 U207 ( .A1(\mem[2][6] ), .A2(n918), .ZN(n134) );
  OAI21_X1 U208 ( .B1(n960), .B2(n918), .A(n136), .ZN(n462) );
  NAND2_X1 U209 ( .A1(\mem[2][8] ), .A2(n918), .ZN(n136) );
  OAI21_X1 U210 ( .B1(n929), .B2(n127), .A(n167), .ZN(n493) );
  NAND2_X1 U211 ( .A1(\mem[2][39] ), .A2(n917), .ZN(n167) );
  OAI21_X1 U212 ( .B1(n967), .B2(n916), .A(n170), .ZN(n495) );
  NAND2_X1 U213 ( .A1(\mem[3][1] ), .A2(n914), .ZN(n170) );
  OAI21_X1 U214 ( .B1(n966), .B2(n916), .A(n171), .ZN(n496) );
  NAND2_X1 U215 ( .A1(\mem[3][2] ), .A2(n914), .ZN(n171) );
  OAI21_X1 U216 ( .B1(n965), .B2(n916), .A(n172), .ZN(n497) );
  NAND2_X1 U217 ( .A1(\mem[3][3] ), .A2(n914), .ZN(n172) );
  OAI21_X1 U218 ( .B1(n964), .B2(n916), .A(n173), .ZN(n498) );
  NAND2_X1 U219 ( .A1(\mem[3][4] ), .A2(n915), .ZN(n173) );
  OAI21_X1 U220 ( .B1(n963), .B2(n916), .A(n174), .ZN(n499) );
  NAND2_X1 U221 ( .A1(\mem[3][5] ), .A2(n915), .ZN(n174) );
  OAI21_X1 U222 ( .B1(n962), .B2(n916), .A(n175), .ZN(n500) );
  NAND2_X1 U223 ( .A1(\mem[3][6] ), .A2(n915), .ZN(n175) );
  OAI21_X1 U224 ( .B1(n960), .B2(n916), .A(n177), .ZN(n502) );
  NAND2_X1 U225 ( .A1(\mem[3][8] ), .A2(n914), .ZN(n177) );
  OAI21_X1 U226 ( .B1(n929), .B2(n916), .A(n208), .ZN(n533) );
  NAND2_X1 U227 ( .A1(\mem[3][39] ), .A2(n914), .ZN(n208) );
  OAI21_X1 U228 ( .B1(n967), .B2(n911), .A(n211), .ZN(n535) );
  NAND2_X1 U229 ( .A1(\mem[4][1] ), .A2(n911), .ZN(n211) );
  OAI21_X1 U230 ( .B1(n966), .B2(n912), .A(n212), .ZN(n536) );
  NAND2_X1 U231 ( .A1(\mem[4][2] ), .A2(n911), .ZN(n212) );
  OAI21_X1 U232 ( .B1(n965), .B2(n913), .A(n213), .ZN(n537) );
  NAND2_X1 U233 ( .A1(\mem[4][3] ), .A2(n911), .ZN(n213) );
  OAI21_X1 U234 ( .B1(n964), .B2(n911), .A(n214), .ZN(n538) );
  NAND2_X1 U235 ( .A1(\mem[4][4] ), .A2(n912), .ZN(n214) );
  OAI21_X1 U236 ( .B1(n963), .B2(n912), .A(n215), .ZN(n539) );
  NAND2_X1 U237 ( .A1(\mem[4][5] ), .A2(n912), .ZN(n215) );
  OAI21_X1 U238 ( .B1(n962), .B2(n913), .A(n216), .ZN(n540) );
  NAND2_X1 U239 ( .A1(\mem[4][6] ), .A2(n912), .ZN(n216) );
  OAI21_X1 U240 ( .B1(n960), .B2(n911), .A(n218), .ZN(n542) );
  NAND2_X1 U241 ( .A1(\mem[4][8] ), .A2(n913), .ZN(n218) );
  OAI21_X1 U242 ( .B1(n929), .B2(n912), .A(n249), .ZN(n573) );
  NAND2_X1 U243 ( .A1(\mem[4][39] ), .A2(n911), .ZN(n249) );
  OAI21_X1 U244 ( .B1(n967), .B2(n908), .A(n253), .ZN(n575) );
  NAND2_X1 U245 ( .A1(\mem[5][1] ), .A2(n908), .ZN(n253) );
  OAI21_X1 U246 ( .B1(n966), .B2(n909), .A(n254), .ZN(n576) );
  NAND2_X1 U247 ( .A1(\mem[5][2] ), .A2(n908), .ZN(n254) );
  OAI21_X1 U248 ( .B1(n965), .B2(n910), .A(n255), .ZN(n577) );
  NAND2_X1 U249 ( .A1(\mem[5][3] ), .A2(n908), .ZN(n255) );
  OAI21_X1 U250 ( .B1(n964), .B2(n908), .A(n256), .ZN(n578) );
  NAND2_X1 U251 ( .A1(\mem[5][4] ), .A2(n909), .ZN(n256) );
  OAI21_X1 U252 ( .B1(n963), .B2(n909), .A(n257), .ZN(n579) );
  NAND2_X1 U253 ( .A1(\mem[5][5] ), .A2(n909), .ZN(n257) );
  OAI21_X1 U254 ( .B1(n962), .B2(n910), .A(n258), .ZN(n580) );
  NAND2_X1 U255 ( .A1(\mem[5][6] ), .A2(n909), .ZN(n258) );
  OAI21_X1 U256 ( .B1(n960), .B2(n908), .A(n260), .ZN(n582) );
  NAND2_X1 U257 ( .A1(\mem[5][8] ), .A2(n910), .ZN(n260) );
  OAI21_X1 U258 ( .B1(n929), .B2(n909), .A(n291), .ZN(n613) );
  NAND2_X1 U259 ( .A1(\mem[5][39] ), .A2(n908), .ZN(n291) );
  OAI21_X1 U260 ( .B1(n967), .B2(n905), .A(n294), .ZN(n615) );
  NAND2_X1 U261 ( .A1(\mem[6][1] ), .A2(n905), .ZN(n294) );
  OAI21_X1 U262 ( .B1(n966), .B2(n906), .A(n295), .ZN(n616) );
  NAND2_X1 U263 ( .A1(\mem[6][2] ), .A2(n905), .ZN(n295) );
  OAI21_X1 U264 ( .B1(n965), .B2(n907), .A(n296), .ZN(n617) );
  NAND2_X1 U265 ( .A1(\mem[6][3] ), .A2(n905), .ZN(n296) );
  OAI21_X1 U266 ( .B1(n964), .B2(n905), .A(n297), .ZN(n618) );
  NAND2_X1 U267 ( .A1(\mem[6][4] ), .A2(n906), .ZN(n297) );
  OAI21_X1 U268 ( .B1(n963), .B2(n906), .A(n298), .ZN(n619) );
  NAND2_X1 U269 ( .A1(\mem[6][5] ), .A2(n906), .ZN(n298) );
  OAI21_X1 U270 ( .B1(n962), .B2(n907), .A(n299), .ZN(n620) );
  NAND2_X1 U271 ( .A1(\mem[6][6] ), .A2(n906), .ZN(n299) );
  OAI21_X1 U272 ( .B1(n960), .B2(n905), .A(n301), .ZN(n622) );
  NAND2_X1 U273 ( .A1(\mem[6][8] ), .A2(n907), .ZN(n301) );
  OAI21_X1 U274 ( .B1(n929), .B2(n906), .A(n332), .ZN(n653) );
  NAND2_X1 U275 ( .A1(\mem[6][39] ), .A2(n905), .ZN(n332) );
  OAI21_X1 U276 ( .B1(n967), .B2(n903), .A(n335), .ZN(n655) );
  NAND2_X1 U277 ( .A1(\mem[7][1] ), .A2(n333), .ZN(n335) );
  OAI21_X1 U278 ( .B1(n966), .B2(n902), .A(n336), .ZN(n656) );
  NAND2_X1 U279 ( .A1(\mem[7][2] ), .A2(n333), .ZN(n336) );
  OAI21_X1 U280 ( .B1(n965), .B2(n333), .A(n337), .ZN(n657) );
  NAND2_X1 U281 ( .A1(\mem[7][3] ), .A2(n902), .ZN(n337) );
  OAI21_X1 U282 ( .B1(n964), .B2(n333), .A(n338), .ZN(n658) );
  NAND2_X1 U283 ( .A1(\mem[7][4] ), .A2(n333), .ZN(n338) );
  OAI21_X1 U284 ( .B1(n963), .B2(n333), .A(n339), .ZN(n659) );
  NAND2_X1 U285 ( .A1(\mem[7][5] ), .A2(n333), .ZN(n339) );
  OAI21_X1 U286 ( .B1(n962), .B2(n333), .A(n340), .ZN(n660) );
  NAND2_X1 U287 ( .A1(\mem[7][6] ), .A2(n333), .ZN(n340) );
  OAI21_X1 U288 ( .B1(n960), .B2(n333), .A(n342), .ZN(n662) );
  NAND2_X1 U289 ( .A1(\mem[7][8] ), .A2(n902), .ZN(n342) );
  OAI21_X1 U290 ( .B1(n929), .B2(n333), .A(n373), .ZN(n693) );
  NAND2_X1 U291 ( .A1(\mem[7][39] ), .A2(n333), .ZN(n373) );
  OAI21_X1 U292 ( .B1(n968), .B2(n921), .A(n87), .ZN(n414) );
  NAND2_X1 U293 ( .A1(\mem[1][0] ), .A2(n920), .ZN(n87) );
  OAI21_X1 U294 ( .B1(n961), .B2(n922), .A(n94), .ZN(n421) );
  NAND2_X1 U295 ( .A1(\mem[1][7] ), .A2(n922), .ZN(n94) );
  OAI21_X1 U296 ( .B1(n959), .B2(n921), .A(n96), .ZN(n423) );
  NAND2_X1 U297 ( .A1(\mem[1][9] ), .A2(n922), .ZN(n96) );
  OAI21_X1 U298 ( .B1(n958), .B2(n920), .A(n97), .ZN(n424) );
  NAND2_X1 U299 ( .A1(\mem[1][10] ), .A2(n922), .ZN(n97) );
  OAI21_X1 U300 ( .B1(n957), .B2(n86), .A(n98), .ZN(n425) );
  NAND2_X1 U301 ( .A1(\mem[1][11] ), .A2(n920), .ZN(n98) );
  OAI21_X1 U302 ( .B1(n956), .B2(n86), .A(n99), .ZN(n426) );
  NAND2_X1 U303 ( .A1(\mem[1][12] ), .A2(n922), .ZN(n99) );
  OAI21_X1 U304 ( .B1(n955), .B2(n86), .A(n100), .ZN(n427) );
  NAND2_X1 U305 ( .A1(\mem[1][13] ), .A2(n921), .ZN(n100) );
  OAI21_X1 U306 ( .B1(n954), .B2(n86), .A(n101), .ZN(n428) );
  NAND2_X1 U307 ( .A1(\mem[1][14] ), .A2(n920), .ZN(n101) );
  OAI21_X1 U308 ( .B1(n953), .B2(n86), .A(n102), .ZN(n429) );
  NAND2_X1 U309 ( .A1(\mem[1][15] ), .A2(n922), .ZN(n102) );
  OAI21_X1 U310 ( .B1(n952), .B2(n86), .A(n103), .ZN(n430) );
  NAND2_X1 U311 ( .A1(\mem[1][16] ), .A2(n922), .ZN(n103) );
  OAI21_X1 U312 ( .B1(n951), .B2(n86), .A(n104), .ZN(n431) );
  NAND2_X1 U313 ( .A1(\mem[1][17] ), .A2(n922), .ZN(n104) );
  OAI21_X1 U314 ( .B1(n950), .B2(n86), .A(n105), .ZN(n432) );
  NAND2_X1 U315 ( .A1(\mem[1][18] ), .A2(n922), .ZN(n105) );
  OAI21_X1 U316 ( .B1(n968), .B2(n917), .A(n128), .ZN(n454) );
  NAND2_X1 U317 ( .A1(\mem[2][0] ), .A2(n918), .ZN(n128) );
  OAI21_X1 U318 ( .B1(n961), .B2(n917), .A(n135), .ZN(n461) );
  NAND2_X1 U319 ( .A1(\mem[2][7] ), .A2(n127), .ZN(n135) );
  OAI21_X1 U320 ( .B1(n959), .B2(n917), .A(n137), .ZN(n463) );
  NAND2_X1 U321 ( .A1(\mem[2][9] ), .A2(n127), .ZN(n137) );
  OAI21_X1 U322 ( .B1(n958), .B2(n917), .A(n138), .ZN(n464) );
  NAND2_X1 U323 ( .A1(\mem[2][10] ), .A2(n127), .ZN(n138) );
  OAI21_X1 U324 ( .B1(n957), .B2(n917), .A(n139), .ZN(n465) );
  NAND2_X1 U325 ( .A1(\mem[2][11] ), .A2(n917), .ZN(n139) );
  OAI21_X1 U326 ( .B1(n956), .B2(n917), .A(n140), .ZN(n466) );
  NAND2_X1 U327 ( .A1(\mem[2][12] ), .A2(n918), .ZN(n140) );
  OAI21_X1 U328 ( .B1(n955), .B2(n917), .A(n141), .ZN(n467) );
  NAND2_X1 U329 ( .A1(\mem[2][13] ), .A2(n127), .ZN(n141) );
  OAI21_X1 U330 ( .B1(n954), .B2(n917), .A(n142), .ZN(n468) );
  NAND2_X1 U331 ( .A1(\mem[2][14] ), .A2(n127), .ZN(n142) );
  OAI21_X1 U332 ( .B1(n953), .B2(n917), .A(n143), .ZN(n469) );
  NAND2_X1 U333 ( .A1(\mem[2][15] ), .A2(n918), .ZN(n143) );
  OAI21_X1 U334 ( .B1(n952), .B2(n917), .A(n144), .ZN(n470) );
  NAND2_X1 U335 ( .A1(\mem[2][16] ), .A2(n127), .ZN(n144) );
  OAI21_X1 U336 ( .B1(n951), .B2(n917), .A(n145), .ZN(n471) );
  NAND2_X1 U337 ( .A1(\mem[2][17] ), .A2(n918), .ZN(n145) );
  OAI21_X1 U338 ( .B1(n950), .B2(n917), .A(n146), .ZN(n472) );
  NAND2_X1 U339 ( .A1(\mem[2][18] ), .A2(n917), .ZN(n146) );
  OAI21_X1 U340 ( .B1(n968), .B2(n916), .A(n169), .ZN(n494) );
  NAND2_X1 U341 ( .A1(\mem[3][0] ), .A2(n914), .ZN(n169) );
  OAI21_X1 U342 ( .B1(n961), .B2(n914), .A(n176), .ZN(n501) );
  NAND2_X1 U343 ( .A1(\mem[3][7] ), .A2(n914), .ZN(n176) );
  OAI21_X1 U344 ( .B1(n959), .B2(n915), .A(n178), .ZN(n503) );
  NAND2_X1 U345 ( .A1(\mem[3][9] ), .A2(n916), .ZN(n178) );
  OAI21_X1 U346 ( .B1(n958), .B2(n168), .A(n179), .ZN(n504) );
  NAND2_X1 U347 ( .A1(\mem[3][10] ), .A2(n915), .ZN(n179) );
  OAI21_X1 U348 ( .B1(n957), .B2(n168), .A(n180), .ZN(n505) );
  NAND2_X1 U349 ( .A1(\mem[3][11] ), .A2(n916), .ZN(n180) );
  OAI21_X1 U350 ( .B1(n956), .B2(n168), .A(n181), .ZN(n506) );
  NAND2_X1 U351 ( .A1(\mem[3][12] ), .A2(n916), .ZN(n181) );
  OAI21_X1 U352 ( .B1(n955), .B2(n168), .A(n182), .ZN(n507) );
  NAND2_X1 U353 ( .A1(\mem[3][13] ), .A2(n915), .ZN(n182) );
  OAI21_X1 U354 ( .B1(n954), .B2(n168), .A(n183), .ZN(n508) );
  NAND2_X1 U355 ( .A1(\mem[3][14] ), .A2(n916), .ZN(n183) );
  OAI21_X1 U356 ( .B1(n953), .B2(n168), .A(n184), .ZN(n509) );
  NAND2_X1 U357 ( .A1(\mem[3][15] ), .A2(n916), .ZN(n184) );
  OAI21_X1 U358 ( .B1(n952), .B2(n168), .A(n185), .ZN(n510) );
  NAND2_X1 U359 ( .A1(\mem[3][16] ), .A2(n914), .ZN(n185) );
  OAI21_X1 U360 ( .B1(n951), .B2(n168), .A(n186), .ZN(n511) );
  NAND2_X1 U361 ( .A1(\mem[3][17] ), .A2(n168), .ZN(n186) );
  OAI21_X1 U362 ( .B1(n950), .B2(n168), .A(n187), .ZN(n512) );
  NAND2_X1 U363 ( .A1(\mem[3][18] ), .A2(n168), .ZN(n187) );
  OAI21_X1 U364 ( .B1(n968), .B2(n913), .A(n210), .ZN(n534) );
  NAND2_X1 U365 ( .A1(\mem[4][0] ), .A2(n911), .ZN(n210) );
  OAI21_X1 U366 ( .B1(n961), .B2(n912), .A(n217), .ZN(n541) );
  NAND2_X1 U367 ( .A1(\mem[4][7] ), .A2(n913), .ZN(n217) );
  OAI21_X1 U368 ( .B1(n959), .B2(n911), .A(n219), .ZN(n543) );
  NAND2_X1 U369 ( .A1(\mem[4][9] ), .A2(n913), .ZN(n219) );
  OAI21_X1 U370 ( .B1(n958), .B2(n209), .A(n220), .ZN(n544) );
  NAND2_X1 U371 ( .A1(\mem[4][10] ), .A2(n913), .ZN(n220) );
  OAI21_X1 U372 ( .B1(n957), .B2(n209), .A(n221), .ZN(n545) );
  NAND2_X1 U373 ( .A1(\mem[4][11] ), .A2(n913), .ZN(n221) );
  OAI21_X1 U374 ( .B1(n956), .B2(n209), .A(n222), .ZN(n546) );
  NAND2_X1 U375 ( .A1(\mem[4][12] ), .A2(n911), .ZN(n222) );
  OAI21_X1 U376 ( .B1(n955), .B2(n209), .A(n223), .ZN(n547) );
  NAND2_X1 U377 ( .A1(\mem[4][13] ), .A2(n912), .ZN(n223) );
  OAI21_X1 U378 ( .B1(n954), .B2(n209), .A(n224), .ZN(n548) );
  NAND2_X1 U379 ( .A1(\mem[4][14] ), .A2(n913), .ZN(n224) );
  OAI21_X1 U380 ( .B1(n953), .B2(n209), .A(n225), .ZN(n549) );
  NAND2_X1 U381 ( .A1(\mem[4][15] ), .A2(n911), .ZN(n225) );
  OAI21_X1 U382 ( .B1(n952), .B2(n209), .A(n226), .ZN(n550) );
  NAND2_X1 U383 ( .A1(\mem[4][16] ), .A2(n913), .ZN(n226) );
  OAI21_X1 U384 ( .B1(n951), .B2(n209), .A(n227), .ZN(n551) );
  NAND2_X1 U385 ( .A1(\mem[4][17] ), .A2(n913), .ZN(n227) );
  OAI21_X1 U386 ( .B1(n950), .B2(n209), .A(n228), .ZN(n552) );
  NAND2_X1 U387 ( .A1(\mem[4][18] ), .A2(n913), .ZN(n228) );
  OAI21_X1 U388 ( .B1(n968), .B2(n251), .A(n252), .ZN(n574) );
  NAND2_X1 U389 ( .A1(\mem[5][0] ), .A2(n908), .ZN(n252) );
  OAI21_X1 U390 ( .B1(n961), .B2(n251), .A(n259), .ZN(n581) );
  NAND2_X1 U391 ( .A1(\mem[5][7] ), .A2(n910), .ZN(n259) );
  OAI21_X1 U392 ( .B1(n959), .B2(n251), .A(n261), .ZN(n583) );
  NAND2_X1 U393 ( .A1(\mem[5][9] ), .A2(n910), .ZN(n261) );
  OAI21_X1 U394 ( .B1(n958), .B2(n251), .A(n262), .ZN(n584) );
  NAND2_X1 U395 ( .A1(\mem[5][10] ), .A2(n910), .ZN(n262) );
  OAI21_X1 U396 ( .B1(n957), .B2(n251), .A(n263), .ZN(n585) );
  NAND2_X1 U397 ( .A1(\mem[5][11] ), .A2(n910), .ZN(n263) );
  OAI21_X1 U398 ( .B1(n956), .B2(n251), .A(n264), .ZN(n586) );
  NAND2_X1 U399 ( .A1(\mem[5][12] ), .A2(n908), .ZN(n264) );
  OAI21_X1 U400 ( .B1(n955), .B2(n251), .A(n265), .ZN(n587) );
  NAND2_X1 U401 ( .A1(\mem[5][13] ), .A2(n909), .ZN(n265) );
  OAI21_X1 U402 ( .B1(n954), .B2(n251), .A(n266), .ZN(n588) );
  NAND2_X1 U403 ( .A1(\mem[5][14] ), .A2(n910), .ZN(n266) );
  OAI21_X1 U404 ( .B1(n953), .B2(n251), .A(n267), .ZN(n589) );
  NAND2_X1 U405 ( .A1(\mem[5][15] ), .A2(n908), .ZN(n267) );
  OAI21_X1 U406 ( .B1(n952), .B2(n251), .A(n268), .ZN(n590) );
  NAND2_X1 U407 ( .A1(\mem[5][16] ), .A2(n910), .ZN(n268) );
  OAI21_X1 U408 ( .B1(n951), .B2(n251), .A(n269), .ZN(n591) );
  NAND2_X1 U409 ( .A1(\mem[5][17] ), .A2(n910), .ZN(n269) );
  OAI21_X1 U410 ( .B1(n950), .B2(n251), .A(n270), .ZN(n592) );
  NAND2_X1 U411 ( .A1(\mem[5][18] ), .A2(n910), .ZN(n270) );
  OAI21_X1 U412 ( .B1(n968), .B2(n292), .A(n293), .ZN(n614) );
  NAND2_X1 U413 ( .A1(\mem[6][0] ), .A2(n905), .ZN(n293) );
  OAI21_X1 U414 ( .B1(n961), .B2(n292), .A(n300), .ZN(n621) );
  NAND2_X1 U415 ( .A1(\mem[6][7] ), .A2(n907), .ZN(n300) );
  OAI21_X1 U416 ( .B1(n959), .B2(n292), .A(n302), .ZN(n623) );
  NAND2_X1 U417 ( .A1(\mem[6][9] ), .A2(n907), .ZN(n302) );
  OAI21_X1 U418 ( .B1(n958), .B2(n292), .A(n303), .ZN(n624) );
  NAND2_X1 U419 ( .A1(\mem[6][10] ), .A2(n907), .ZN(n303) );
  OAI21_X1 U420 ( .B1(n957), .B2(n292), .A(n304), .ZN(n625) );
  NAND2_X1 U421 ( .A1(\mem[6][11] ), .A2(n907), .ZN(n304) );
  OAI21_X1 U422 ( .B1(n956), .B2(n292), .A(n305), .ZN(n626) );
  NAND2_X1 U423 ( .A1(\mem[6][12] ), .A2(n905), .ZN(n305) );
  OAI21_X1 U424 ( .B1(n955), .B2(n292), .A(n306), .ZN(n627) );
  NAND2_X1 U425 ( .A1(\mem[6][13] ), .A2(n906), .ZN(n306) );
  OAI21_X1 U426 ( .B1(n954), .B2(n292), .A(n307), .ZN(n628) );
  NAND2_X1 U427 ( .A1(\mem[6][14] ), .A2(n907), .ZN(n307) );
  OAI21_X1 U428 ( .B1(n953), .B2(n292), .A(n308), .ZN(n629) );
  NAND2_X1 U429 ( .A1(\mem[6][15] ), .A2(n905), .ZN(n308) );
  OAI21_X1 U430 ( .B1(n952), .B2(n292), .A(n309), .ZN(n630) );
  NAND2_X1 U431 ( .A1(\mem[6][16] ), .A2(n907), .ZN(n309) );
  OAI21_X1 U432 ( .B1(n951), .B2(n292), .A(n310), .ZN(n631) );
  NAND2_X1 U433 ( .A1(\mem[6][17] ), .A2(n907), .ZN(n310) );
  OAI21_X1 U434 ( .B1(n950), .B2(n292), .A(n311), .ZN(n632) );
  NAND2_X1 U435 ( .A1(\mem[6][18] ), .A2(n907), .ZN(n311) );
  OAI21_X1 U436 ( .B1(n968), .B2(n903), .A(n334), .ZN(n654) );
  NAND2_X1 U437 ( .A1(\mem[7][0] ), .A2(n333), .ZN(n334) );
  OAI21_X1 U438 ( .B1(n961), .B2(n903), .A(n341), .ZN(n661) );
  NAND2_X1 U439 ( .A1(\mem[7][7] ), .A2(n902), .ZN(n341) );
  OAI21_X1 U440 ( .B1(n959), .B2(n903), .A(n343), .ZN(n663) );
  NAND2_X1 U441 ( .A1(\mem[7][9] ), .A2(n902), .ZN(n343) );
  OAI21_X1 U442 ( .B1(n958), .B2(n903), .A(n344), .ZN(n664) );
  NAND2_X1 U443 ( .A1(\mem[7][10] ), .A2(n902), .ZN(n344) );
  OAI21_X1 U444 ( .B1(n957), .B2(n904), .A(n345), .ZN(n665) );
  NAND2_X1 U445 ( .A1(\mem[7][11] ), .A2(n333), .ZN(n345) );
  OAI21_X1 U446 ( .B1(n956), .B2(n903), .A(n346), .ZN(n666) );
  NAND2_X1 U447 ( .A1(\mem[7][12] ), .A2(n902), .ZN(n346) );
  OAI21_X1 U448 ( .B1(n955), .B2(n904), .A(n347), .ZN(n667) );
  NAND2_X1 U449 ( .A1(\mem[7][13] ), .A2(n333), .ZN(n347) );
  OAI21_X1 U450 ( .B1(n954), .B2(n903), .A(n348), .ZN(n668) );
  NAND2_X1 U451 ( .A1(\mem[7][14] ), .A2(n902), .ZN(n348) );
  OAI21_X1 U452 ( .B1(n953), .B2(n904), .A(n349), .ZN(n669) );
  NAND2_X1 U453 ( .A1(\mem[7][15] ), .A2(n902), .ZN(n349) );
  OAI21_X1 U454 ( .B1(n952), .B2(n903), .A(n350), .ZN(n670) );
  NAND2_X1 U455 ( .A1(\mem[7][16] ), .A2(n902), .ZN(n350) );
  OAI21_X1 U456 ( .B1(n951), .B2(n903), .A(n351), .ZN(n671) );
  NAND2_X1 U457 ( .A1(\mem[7][17] ), .A2(n902), .ZN(n351) );
  OAI21_X1 U458 ( .B1(n950), .B2(n904), .A(n352), .ZN(n672) );
  NAND2_X1 U459 ( .A1(\mem[7][18] ), .A2(n902), .ZN(n352) );
  OAI21_X1 U460 ( .B1(n44), .B2(n968), .A(n45), .ZN(n374) );
  NAND2_X1 U461 ( .A1(\mem[0][0] ), .A2(n924), .ZN(n45) );
  OAI21_X1 U462 ( .B1(n44), .B2(n961), .A(n52), .ZN(n381) );
  NAND2_X1 U463 ( .A1(\mem[0][7] ), .A2(n924), .ZN(n52) );
  OAI21_X1 U464 ( .B1(n44), .B2(n958), .A(n55), .ZN(n384) );
  NAND2_X1 U465 ( .A1(\mem[0][10] ), .A2(n924), .ZN(n55) );
  OAI21_X1 U466 ( .B1(n44), .B2(n957), .A(n56), .ZN(n385) );
  NAND2_X1 U467 ( .A1(\mem[0][11] ), .A2(n925), .ZN(n56) );
  OAI21_X1 U468 ( .B1(n44), .B2(n956), .A(n57), .ZN(n386) );
  NAND2_X1 U469 ( .A1(\mem[0][12] ), .A2(n925), .ZN(n57) );
  OAI21_X1 U470 ( .B1(n44), .B2(n955), .A(n58), .ZN(n387) );
  NAND2_X1 U471 ( .A1(\mem[0][13] ), .A2(n923), .ZN(n58) );
  OAI21_X1 U472 ( .B1(n44), .B2(n954), .A(n59), .ZN(n388) );
  NAND2_X1 U473 ( .A1(\mem[0][14] ), .A2(n925), .ZN(n59) );
  OAI21_X1 U474 ( .B1(n44), .B2(n953), .A(n60), .ZN(n389) );
  NAND2_X1 U475 ( .A1(\mem[0][15] ), .A2(n925), .ZN(n60) );
  OAI21_X1 U476 ( .B1(n44), .B2(n952), .A(n61), .ZN(n390) );
  NAND2_X1 U477 ( .A1(\mem[0][16] ), .A2(n924), .ZN(n61) );
  OAI21_X1 U478 ( .B1(n44), .B2(n951), .A(n62), .ZN(n391) );
  NAND2_X1 U479 ( .A1(\mem[0][17] ), .A2(n924), .ZN(n62) );
  OAI21_X1 U480 ( .B1(n44), .B2(n950), .A(n63), .ZN(n392) );
  NAND2_X1 U481 ( .A1(\mem[0][18] ), .A2(n924), .ZN(n63) );
  OAI21_X1 U482 ( .B1(n44), .B2(n949), .A(n64), .ZN(n393) );
  NAND2_X1 U483 ( .A1(\mem[0][19] ), .A2(n924), .ZN(n64) );
  OAI21_X1 U484 ( .B1(n44), .B2(n948), .A(n65), .ZN(n394) );
  NAND2_X1 U485 ( .A1(\mem[0][20] ), .A2(n924), .ZN(n65) );
  OAI21_X1 U486 ( .B1(n949), .B2(n86), .A(n106), .ZN(n433) );
  NAND2_X1 U487 ( .A1(\mem[1][19] ), .A2(n922), .ZN(n106) );
  OAI21_X1 U488 ( .B1(n948), .B2(n86), .A(n107), .ZN(n434) );
  NAND2_X1 U489 ( .A1(\mem[1][20] ), .A2(n922), .ZN(n107) );
  OAI21_X1 U490 ( .B1(n947), .B2(n86), .A(n108), .ZN(n435) );
  NAND2_X1 U491 ( .A1(\mem[1][21] ), .A2(n922), .ZN(n108) );
  OAI21_X1 U492 ( .B1(n949), .B2(n918), .A(n147), .ZN(n473) );
  NAND2_X1 U493 ( .A1(\mem[2][19] ), .A2(n919), .ZN(n147) );
  OAI21_X1 U494 ( .B1(n948), .B2(n918), .A(n148), .ZN(n474) );
  NAND2_X1 U495 ( .A1(\mem[2][20] ), .A2(n918), .ZN(n148) );
  OAI21_X1 U496 ( .B1(n947), .B2(n918), .A(n149), .ZN(n475) );
  NAND2_X1 U497 ( .A1(\mem[2][21] ), .A2(n917), .ZN(n149) );
  OAI21_X1 U498 ( .B1(n949), .B2(n168), .A(n188), .ZN(n513) );
  NAND2_X1 U499 ( .A1(\mem[3][19] ), .A2(n168), .ZN(n188) );
  OAI21_X1 U500 ( .B1(n948), .B2(n168), .A(n189), .ZN(n514) );
  NAND2_X1 U501 ( .A1(\mem[3][20] ), .A2(n168), .ZN(n189) );
  OAI21_X1 U502 ( .B1(n947), .B2(n168), .A(n190), .ZN(n515) );
  NAND2_X1 U503 ( .A1(\mem[3][21] ), .A2(n168), .ZN(n190) );
  OAI21_X1 U504 ( .B1(n949), .B2(n209), .A(n229), .ZN(n553) );
  NAND2_X1 U505 ( .A1(\mem[4][19] ), .A2(n913), .ZN(n229) );
  OAI21_X1 U506 ( .B1(n948), .B2(n209), .A(n230), .ZN(n554) );
  NAND2_X1 U507 ( .A1(\mem[4][20] ), .A2(n913), .ZN(n230) );
  OAI21_X1 U508 ( .B1(n947), .B2(n209), .A(n231), .ZN(n555) );
  NAND2_X1 U509 ( .A1(\mem[4][21] ), .A2(n913), .ZN(n231) );
  OAI21_X1 U510 ( .B1(n949), .B2(n910), .A(n271), .ZN(n593) );
  NAND2_X1 U511 ( .A1(\mem[5][19] ), .A2(n910), .ZN(n271) );
  OAI21_X1 U512 ( .B1(n948), .B2(n909), .A(n272), .ZN(n594) );
  NAND2_X1 U513 ( .A1(\mem[5][20] ), .A2(n910), .ZN(n272) );
  OAI21_X1 U514 ( .B1(n947), .B2(n908), .A(n273), .ZN(n595) );
  NAND2_X1 U515 ( .A1(\mem[5][21] ), .A2(n910), .ZN(n273) );
  OAI21_X1 U516 ( .B1(n949), .B2(n907), .A(n312), .ZN(n633) );
  NAND2_X1 U517 ( .A1(\mem[6][19] ), .A2(n907), .ZN(n312) );
  OAI21_X1 U518 ( .B1(n948), .B2(n906), .A(n313), .ZN(n634) );
  NAND2_X1 U519 ( .A1(\mem[6][20] ), .A2(n907), .ZN(n313) );
  OAI21_X1 U520 ( .B1(n947), .B2(n905), .A(n314), .ZN(n635) );
  NAND2_X1 U521 ( .A1(\mem[6][21] ), .A2(n907), .ZN(n314) );
  OAI21_X1 U522 ( .B1(n949), .B2(n903), .A(n353), .ZN(n673) );
  NAND2_X1 U523 ( .A1(\mem[7][19] ), .A2(n902), .ZN(n353) );
  OAI21_X1 U524 ( .B1(n948), .B2(n903), .A(n354), .ZN(n674) );
  NAND2_X1 U525 ( .A1(\mem[7][20] ), .A2(n902), .ZN(n354) );
  OAI21_X1 U526 ( .B1(n947), .B2(n903), .A(n355), .ZN(n675) );
  NAND2_X1 U527 ( .A1(\mem[7][21] ), .A2(n902), .ZN(n355) );
  OAI21_X1 U528 ( .B1(n946), .B2(n86), .A(n109), .ZN(n436) );
  NAND2_X1 U529 ( .A1(\mem[1][22] ), .A2(n922), .ZN(n109) );
  OAI21_X1 U530 ( .B1(n945), .B2(n922), .A(n110), .ZN(n437) );
  NAND2_X1 U531 ( .A1(\mem[1][23] ), .A2(n922), .ZN(n110) );
  OAI21_X1 U532 ( .B1(n944), .B2(n922), .A(n111), .ZN(n438) );
  NAND2_X1 U533 ( .A1(\mem[1][24] ), .A2(n921), .ZN(n111) );
  OAI21_X1 U534 ( .B1(n943), .B2(n921), .A(n112), .ZN(n439) );
  NAND2_X1 U535 ( .A1(\mem[1][25] ), .A2(n921), .ZN(n112) );
  OAI21_X1 U536 ( .B1(n942), .B2(n920), .A(n113), .ZN(n440) );
  NAND2_X1 U537 ( .A1(\mem[1][26] ), .A2(n921), .ZN(n113) );
  OAI21_X1 U538 ( .B1(n941), .B2(n86), .A(n114), .ZN(n441) );
  NAND2_X1 U539 ( .A1(\mem[1][27] ), .A2(n921), .ZN(n114) );
  OAI21_X1 U540 ( .B1(n940), .B2(n86), .A(n115), .ZN(n442) );
  NAND2_X1 U541 ( .A1(\mem[1][28] ), .A2(n921), .ZN(n115) );
  OAI21_X1 U542 ( .B1(n939), .B2(n86), .A(n116), .ZN(n443) );
  NAND2_X1 U543 ( .A1(\mem[1][29] ), .A2(n921), .ZN(n116) );
  OAI21_X1 U544 ( .B1(n938), .B2(n86), .A(n117), .ZN(n444) );
  NAND2_X1 U545 ( .A1(\mem[1][30] ), .A2(n921), .ZN(n117) );
  OAI21_X1 U546 ( .B1(n946), .B2(n918), .A(n150), .ZN(n476) );
  NAND2_X1 U547 ( .A1(\mem[2][22] ), .A2(n918), .ZN(n150) );
  OAI21_X1 U548 ( .B1(n945), .B2(n918), .A(n151), .ZN(n477) );
  NAND2_X1 U549 ( .A1(\mem[2][23] ), .A2(n917), .ZN(n151) );
  OAI21_X1 U550 ( .B1(n944), .B2(n918), .A(n152), .ZN(n478) );
  NAND2_X1 U551 ( .A1(\mem[2][24] ), .A2(n127), .ZN(n152) );
  OAI21_X1 U552 ( .B1(n943), .B2(n918), .A(n153), .ZN(n479) );
  NAND2_X1 U553 ( .A1(\mem[2][25] ), .A2(n127), .ZN(n153) );
  OAI21_X1 U554 ( .B1(n942), .B2(n918), .A(n154), .ZN(n480) );
  NAND2_X1 U555 ( .A1(\mem[2][26] ), .A2(n127), .ZN(n154) );
  OAI21_X1 U556 ( .B1(n941), .B2(n918), .A(n155), .ZN(n481) );
  NAND2_X1 U557 ( .A1(\mem[2][27] ), .A2(n127), .ZN(n155) );
  OAI21_X1 U558 ( .B1(n940), .B2(n918), .A(n156), .ZN(n482) );
  NAND2_X1 U559 ( .A1(\mem[2][28] ), .A2(n127), .ZN(n156) );
  OAI21_X1 U560 ( .B1(n939), .B2(n918), .A(n157), .ZN(n483) );
  NAND2_X1 U561 ( .A1(\mem[2][29] ), .A2(n127), .ZN(n157) );
  OAI21_X1 U562 ( .B1(n938), .B2(n918), .A(n158), .ZN(n484) );
  NAND2_X1 U563 ( .A1(\mem[2][30] ), .A2(n127), .ZN(n158) );
  OAI21_X1 U564 ( .B1(n946), .B2(n168), .A(n191), .ZN(n516) );
  NAND2_X1 U565 ( .A1(\mem[3][22] ), .A2(n168), .ZN(n191) );
  OAI21_X1 U566 ( .B1(n945), .B2(n168), .A(n192), .ZN(n517) );
  NAND2_X1 U567 ( .A1(\mem[3][23] ), .A2(n168), .ZN(n192) );
  OAI21_X1 U568 ( .B1(n944), .B2(n916), .A(n193), .ZN(n518) );
  NAND2_X1 U569 ( .A1(\mem[3][24] ), .A2(n915), .ZN(n193) );
  OAI21_X1 U570 ( .B1(n943), .B2(n915), .A(n194), .ZN(n519) );
  NAND2_X1 U571 ( .A1(\mem[3][25] ), .A2(n915), .ZN(n194) );
  OAI21_X1 U572 ( .B1(n942), .B2(n914), .A(n195), .ZN(n520) );
  NAND2_X1 U573 ( .A1(\mem[3][26] ), .A2(n915), .ZN(n195) );
  OAI21_X1 U574 ( .B1(n941), .B2(n168), .A(n196), .ZN(n521) );
  NAND2_X1 U575 ( .A1(\mem[3][27] ), .A2(n915), .ZN(n196) );
  OAI21_X1 U576 ( .B1(n940), .B2(n916), .A(n197), .ZN(n522) );
  NAND2_X1 U577 ( .A1(\mem[3][28] ), .A2(n915), .ZN(n197) );
  OAI21_X1 U578 ( .B1(n939), .B2(n915), .A(n198), .ZN(n523) );
  NAND2_X1 U579 ( .A1(\mem[3][29] ), .A2(n915), .ZN(n198) );
  OAI21_X1 U580 ( .B1(n938), .B2(n168), .A(n199), .ZN(n524) );
  NAND2_X1 U581 ( .A1(\mem[3][30] ), .A2(n915), .ZN(n199) );
  OAI21_X1 U582 ( .B1(n946), .B2(n913), .A(n232), .ZN(n556) );
  NAND2_X1 U583 ( .A1(\mem[4][22] ), .A2(n913), .ZN(n232) );
  OAI21_X1 U584 ( .B1(n945), .B2(n913), .A(n233), .ZN(n557) );
  NAND2_X1 U585 ( .A1(\mem[4][23] ), .A2(n913), .ZN(n233) );
  OAI21_X1 U586 ( .B1(n944), .B2(n912), .A(n234), .ZN(n558) );
  NAND2_X1 U587 ( .A1(\mem[4][24] ), .A2(n912), .ZN(n234) );
  OAI21_X1 U588 ( .B1(n943), .B2(n911), .A(n235), .ZN(n559) );
  NAND2_X1 U589 ( .A1(\mem[4][25] ), .A2(n912), .ZN(n235) );
  OAI21_X1 U590 ( .B1(n942), .B2(n209), .A(n236), .ZN(n560) );
  NAND2_X1 U591 ( .A1(\mem[4][26] ), .A2(n912), .ZN(n236) );
  OAI21_X1 U592 ( .B1(n941), .B2(n912), .A(n237), .ZN(n561) );
  NAND2_X1 U593 ( .A1(\mem[4][27] ), .A2(n912), .ZN(n237) );
  OAI21_X1 U594 ( .B1(n940), .B2(n209), .A(n238), .ZN(n562) );
  NAND2_X1 U595 ( .A1(\mem[4][28] ), .A2(n912), .ZN(n238) );
  OAI21_X1 U596 ( .B1(n939), .B2(n209), .A(n239), .ZN(n563) );
  NAND2_X1 U597 ( .A1(\mem[4][29] ), .A2(n912), .ZN(n239) );
  OAI21_X1 U598 ( .B1(n938), .B2(n209), .A(n240), .ZN(n564) );
  NAND2_X1 U599 ( .A1(\mem[4][30] ), .A2(n912), .ZN(n240) );
  OAI21_X1 U600 ( .B1(n946), .B2(n910), .A(n274), .ZN(n596) );
  NAND2_X1 U601 ( .A1(\mem[5][22] ), .A2(n910), .ZN(n274) );
  OAI21_X1 U602 ( .B1(n945), .B2(n909), .A(n275), .ZN(n597) );
  NAND2_X1 U603 ( .A1(\mem[5][23] ), .A2(n910), .ZN(n275) );
  OAI21_X1 U604 ( .B1(n944), .B2(n251), .A(n276), .ZN(n598) );
  NAND2_X1 U605 ( .A1(\mem[5][24] ), .A2(n909), .ZN(n276) );
  OAI21_X1 U606 ( .B1(n943), .B2(n251), .A(n277), .ZN(n599) );
  NAND2_X1 U607 ( .A1(\mem[5][25] ), .A2(n909), .ZN(n277) );
  OAI21_X1 U608 ( .B1(n942), .B2(n251), .A(n278), .ZN(n600) );
  NAND2_X1 U609 ( .A1(\mem[5][26] ), .A2(n909), .ZN(n278) );
  OAI21_X1 U610 ( .B1(n941), .B2(n251), .A(n279), .ZN(n601) );
  NAND2_X1 U611 ( .A1(\mem[5][27] ), .A2(n909), .ZN(n279) );
  OAI21_X1 U612 ( .B1(n940), .B2(n251), .A(n280), .ZN(n602) );
  NAND2_X1 U613 ( .A1(\mem[5][28] ), .A2(n909), .ZN(n280) );
  OAI21_X1 U614 ( .B1(n939), .B2(n251), .A(n281), .ZN(n603) );
  NAND2_X1 U615 ( .A1(\mem[5][29] ), .A2(n909), .ZN(n281) );
  OAI21_X1 U616 ( .B1(n938), .B2(n251), .A(n282), .ZN(n604) );
  NAND2_X1 U617 ( .A1(\mem[5][30] ), .A2(n909), .ZN(n282) );
  OAI21_X1 U618 ( .B1(n946), .B2(n907), .A(n315), .ZN(n636) );
  NAND2_X1 U619 ( .A1(\mem[6][22] ), .A2(n907), .ZN(n315) );
  OAI21_X1 U620 ( .B1(n945), .B2(n906), .A(n316), .ZN(n637) );
  NAND2_X1 U621 ( .A1(\mem[6][23] ), .A2(n907), .ZN(n316) );
  OAI21_X1 U622 ( .B1(n944), .B2(n292), .A(n317), .ZN(n638) );
  NAND2_X1 U623 ( .A1(\mem[6][24] ), .A2(n906), .ZN(n317) );
  OAI21_X1 U624 ( .B1(n943), .B2(n292), .A(n318), .ZN(n639) );
  NAND2_X1 U625 ( .A1(\mem[6][25] ), .A2(n906), .ZN(n318) );
  OAI21_X1 U626 ( .B1(n942), .B2(n292), .A(n319), .ZN(n640) );
  NAND2_X1 U627 ( .A1(\mem[6][26] ), .A2(n906), .ZN(n319) );
  OAI21_X1 U628 ( .B1(n941), .B2(n292), .A(n320), .ZN(n641) );
  NAND2_X1 U629 ( .A1(\mem[6][27] ), .A2(n906), .ZN(n320) );
  OAI21_X1 U630 ( .B1(n940), .B2(n292), .A(n321), .ZN(n642) );
  NAND2_X1 U631 ( .A1(\mem[6][28] ), .A2(n906), .ZN(n321) );
  OAI21_X1 U632 ( .B1(n939), .B2(n292), .A(n322), .ZN(n643) );
  NAND2_X1 U633 ( .A1(\mem[6][29] ), .A2(n906), .ZN(n322) );
  OAI21_X1 U634 ( .B1(n938), .B2(n292), .A(n323), .ZN(n644) );
  NAND2_X1 U635 ( .A1(\mem[6][30] ), .A2(n906), .ZN(n323) );
  OAI21_X1 U636 ( .B1(n946), .B2(n903), .A(n356), .ZN(n676) );
  NAND2_X1 U637 ( .A1(\mem[7][22] ), .A2(n902), .ZN(n356) );
  OAI21_X1 U638 ( .B1(n945), .B2(n903), .A(n357), .ZN(n677) );
  NAND2_X1 U639 ( .A1(\mem[7][23] ), .A2(n902), .ZN(n357) );
  OAI21_X1 U640 ( .B1(n944), .B2(n903), .A(n358), .ZN(n678) );
  NAND2_X1 U641 ( .A1(\mem[7][24] ), .A2(n904), .ZN(n358) );
  OAI21_X1 U642 ( .B1(n943), .B2(n903), .A(n359), .ZN(n679) );
  NAND2_X1 U643 ( .A1(\mem[7][25] ), .A2(n902), .ZN(n359) );
  OAI21_X1 U644 ( .B1(n942), .B2(n903), .A(n360), .ZN(n680) );
  NAND2_X1 U645 ( .A1(\mem[7][26] ), .A2(n904), .ZN(n360) );
  OAI21_X1 U646 ( .B1(n941), .B2(n903), .A(n361), .ZN(n681) );
  NAND2_X1 U647 ( .A1(\mem[7][27] ), .A2(n902), .ZN(n361) );
  OAI21_X1 U648 ( .B1(n940), .B2(n903), .A(n362), .ZN(n682) );
  NAND2_X1 U649 ( .A1(\mem[7][28] ), .A2(n902), .ZN(n362) );
  OAI21_X1 U650 ( .B1(n939), .B2(n903), .A(n363), .ZN(n683) );
  NAND2_X1 U651 ( .A1(\mem[7][29] ), .A2(n903), .ZN(n363) );
  OAI21_X1 U652 ( .B1(n938), .B2(n903), .A(n364), .ZN(n684) );
  NAND2_X1 U653 ( .A1(\mem[7][30] ), .A2(n904), .ZN(n364) );
  OAI21_X1 U654 ( .B1(n44), .B2(n947), .A(n66), .ZN(n395) );
  NAND2_X1 U655 ( .A1(\mem[0][21] ), .A2(n924), .ZN(n66) );
  OAI21_X1 U656 ( .B1(n44), .B2(n946), .A(n67), .ZN(n396) );
  NAND2_X1 U657 ( .A1(\mem[0][22] ), .A2(n924), .ZN(n67) );
  OAI21_X1 U658 ( .B1(n924), .B2(n945), .A(n68), .ZN(n397) );
  NAND2_X1 U659 ( .A1(\mem[0][23] ), .A2(n924), .ZN(n68) );
  OAI21_X1 U660 ( .B1(n923), .B2(n944), .A(n69), .ZN(n398) );
  NAND2_X1 U661 ( .A1(\mem[0][24] ), .A2(n923), .ZN(n69) );
  OAI21_X1 U662 ( .B1(n924), .B2(n943), .A(n70), .ZN(n399) );
  NAND2_X1 U663 ( .A1(\mem[0][25] ), .A2(n923), .ZN(n70) );
  OAI21_X1 U664 ( .B1(n44), .B2(n942), .A(n71), .ZN(n400) );
  NAND2_X1 U665 ( .A1(\mem[0][26] ), .A2(n923), .ZN(n71) );
  OAI21_X1 U666 ( .B1(n924), .B2(n941), .A(n72), .ZN(n401) );
  NAND2_X1 U667 ( .A1(\mem[0][27] ), .A2(n923), .ZN(n72) );
  OAI21_X1 U668 ( .B1(n923), .B2(n940), .A(n73), .ZN(n402) );
  NAND2_X1 U669 ( .A1(\mem[0][28] ), .A2(n923), .ZN(n73) );
  OAI21_X1 U670 ( .B1(n925), .B2(n939), .A(n74), .ZN(n403) );
  NAND2_X1 U671 ( .A1(\mem[0][29] ), .A2(n923), .ZN(n74) );
  OAI21_X1 U672 ( .B1(n925), .B2(n938), .A(n75), .ZN(n404) );
  NAND2_X1 U673 ( .A1(\mem[0][30] ), .A2(n923), .ZN(n75) );
  OAI21_X1 U674 ( .B1(n44), .B2(n937), .A(n76), .ZN(n405) );
  NAND2_X1 U675 ( .A1(\mem[0][31] ), .A2(n923), .ZN(n76) );
  OAI21_X1 U676 ( .B1(n44), .B2(n936), .A(n77), .ZN(n406) );
  NAND2_X1 U677 ( .A1(\mem[0][32] ), .A2(n923), .ZN(n77) );
  OAI21_X1 U678 ( .B1(n44), .B2(n935), .A(n78), .ZN(n407) );
  NAND2_X1 U679 ( .A1(\mem[0][33] ), .A2(n44), .ZN(n78) );
  INV_X1 U680 ( .A(data_in[0]), .ZN(n968) );
  INV_X1 U681 ( .A(data_in[1]), .ZN(n967) );
  INV_X1 U682 ( .A(data_in[2]), .ZN(n966) );
  INV_X1 U683 ( .A(data_in[3]), .ZN(n965) );
  INV_X1 U684 ( .A(data_in[4]), .ZN(n964) );
  INV_X1 U685 ( .A(data_in[5]), .ZN(n963) );
  INV_X1 U686 ( .A(data_in[6]), .ZN(n962) );
  INV_X1 U687 ( .A(data_in[7]), .ZN(n961) );
  INV_X1 U696 ( .A(data_in[8]), .ZN(n960) );
  INV_X1 U697 ( .A(data_in[9]), .ZN(n959) );
  INV_X1 U698 ( .A(data_in[10]), .ZN(n958) );
  INV_X1 U699 ( .A(data_in[11]), .ZN(n957) );
  INV_X1 U700 ( .A(data_in[12]), .ZN(n956) );
  INV_X1 U701 ( .A(data_in[13]), .ZN(n955) );
  INV_X1 U702 ( .A(data_in[14]), .ZN(n954) );
  INV_X1 U703 ( .A(data_in[15]), .ZN(n953) );
  INV_X1 U704 ( .A(data_in[16]), .ZN(n952) );
  INV_X1 U705 ( .A(data_in[17]), .ZN(n951) );
  INV_X1 U706 ( .A(data_in[18]), .ZN(n950) );
  INV_X1 U707 ( .A(data_in[19]), .ZN(n949) );
  INV_X1 U708 ( .A(data_in[20]), .ZN(n948) );
  INV_X1 U709 ( .A(data_in[21]), .ZN(n947) );
  INV_X1 U710 ( .A(data_in[22]), .ZN(n946) );
  INV_X1 U711 ( .A(data_in[23]), .ZN(n945) );
  INV_X1 U712 ( .A(data_in[24]), .ZN(n944) );
  INV_X1 U713 ( .A(data_in[25]), .ZN(n943) );
  INV_X1 U714 ( .A(data_in[26]), .ZN(n942) );
  INV_X1 U715 ( .A(data_in[27]), .ZN(n941) );
  INV_X1 U716 ( .A(data_in[28]), .ZN(n940) );
  INV_X1 U717 ( .A(data_in[29]), .ZN(n939) );
  INV_X1 U718 ( .A(data_in[30]), .ZN(n938) );
  INV_X1 U719 ( .A(data_in[31]), .ZN(n937) );
  INV_X1 U720 ( .A(data_in[32]), .ZN(n936) );
  INV_X1 U721 ( .A(data_in[33]), .ZN(n935) );
  INV_X1 U722 ( .A(data_in[34]), .ZN(n934) );
  INV_X1 U723 ( .A(data_in[35]), .ZN(n933) );
  INV_X1 U724 ( .A(data_in[36]), .ZN(n932) );
  INV_X1 U725 ( .A(data_in[37]), .ZN(n931) );
  INV_X1 U726 ( .A(data_in[38]), .ZN(n930) );
  INV_X1 U727 ( .A(data_in[39]), .ZN(n929) );
  MUX2_X1 U728 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n895), .Z(n1) );
  MUX2_X1 U729 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n895), .Z(n2) );
  MUX2_X1 U730 ( .A(n2), .B(n1), .S(n892), .Z(n3) );
  MUX2_X1 U731 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n895), .Z(n4) );
  MUX2_X1 U732 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n895), .Z(n5) );
  MUX2_X1 U733 ( .A(n5), .B(n4), .S(n894), .Z(n6) );
  MUX2_X1 U734 ( .A(n6), .B(n3), .S(n891), .Z(N52) );
  MUX2_X1 U735 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n896), .Z(n7) );
  MUX2_X1 U736 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n896), .Z(n8) );
  MUX2_X1 U737 ( .A(n8), .B(n7), .S(n893), .Z(n9) );
  MUX2_X1 U738 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n896), .Z(n10) );
  MUX2_X1 U739 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n896), .Z(n11) );
  MUX2_X1 U740 ( .A(n11), .B(n10), .S(n892), .Z(n12) );
  MUX2_X1 U741 ( .A(n12), .B(n9), .S(n891), .Z(N51) );
  MUX2_X1 U742 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n896), .Z(n13) );
  MUX2_X1 U743 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n896), .Z(n14) );
  MUX2_X1 U744 ( .A(n14), .B(n13), .S(n894), .Z(n15) );
  MUX2_X1 U745 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n896), .Z(n16) );
  MUX2_X1 U746 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n896), .Z(n17) );
  MUX2_X1 U747 ( .A(n17), .B(n16), .S(n892), .Z(n18) );
  MUX2_X1 U748 ( .A(n18), .B(n15), .S(n891), .Z(N50) );
  MUX2_X1 U749 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n896), .Z(n19) );
  MUX2_X1 U750 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n896), .Z(n20) );
  MUX2_X1 U751 ( .A(n20), .B(n19), .S(n894), .Z(n21) );
  MUX2_X1 U752 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n896), .Z(n22) );
  MUX2_X1 U753 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n896), .Z(n23) );
  MUX2_X1 U754 ( .A(n23), .B(n22), .S(n893), .Z(n24) );
  MUX2_X1 U755 ( .A(n24), .B(n21), .S(n891), .Z(N49) );
  MUX2_X1 U756 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(N10), .Z(n25) );
  MUX2_X1 U757 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n901), .Z(n26) );
  MUX2_X1 U758 ( .A(n26), .B(n25), .S(n894), .Z(n27) );
  MUX2_X1 U759 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n901), .Z(n28) );
  MUX2_X1 U760 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n900), .Z(n29) );
  MUX2_X1 U761 ( .A(n29), .B(n28), .S(N11), .Z(n30) );
  MUX2_X1 U762 ( .A(n30), .B(n27), .S(n891), .Z(N48) );
  MUX2_X1 U763 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n901), .Z(n31) );
  MUX2_X1 U764 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n901), .Z(n32) );
  MUX2_X1 U765 ( .A(n32), .B(n31), .S(n892), .Z(n33) );
  MUX2_X1 U766 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n901), .Z(n34) );
  MUX2_X1 U767 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n900), .Z(n35) );
  MUX2_X1 U768 ( .A(n35), .B(n34), .S(N11), .Z(n36) );
  MUX2_X1 U769 ( .A(n36), .B(n33), .S(n891), .Z(N47) );
  MUX2_X1 U770 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n896), .Z(n37) );
  MUX2_X1 U771 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n900), .Z(n38) );
  MUX2_X1 U772 ( .A(n38), .B(n37), .S(n893), .Z(n39) );
  MUX2_X1 U773 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n901), .Z(n40) );
  MUX2_X1 U774 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n901), .Z(n41) );
  MUX2_X1 U775 ( .A(n41), .B(n40), .S(N11), .Z(n42) );
  MUX2_X1 U776 ( .A(n42), .B(n39), .S(n891), .Z(N46) );
  MUX2_X1 U777 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n895), .Z(n43) );
  MUX2_X1 U778 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n895), .Z(n694) );
  MUX2_X1 U779 ( .A(n694), .B(n43), .S(n894), .Z(n695) );
  MUX2_X1 U780 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n895), .Z(n696) );
  MUX2_X1 U781 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n900), .Z(n697) );
  MUX2_X1 U782 ( .A(n697), .B(n696), .S(N11), .Z(n698) );
  MUX2_X1 U783 ( .A(n698), .B(n695), .S(n891), .Z(N45) );
  MUX2_X1 U784 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n895), .Z(n699) );
  MUX2_X1 U785 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n895), .Z(n700) );
  MUX2_X1 U786 ( .A(n700), .B(n699), .S(n892), .Z(n701) );
  MUX2_X1 U787 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n895), .Z(n702) );
  MUX2_X1 U788 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n900), .Z(n703) );
  MUX2_X1 U789 ( .A(n703), .B(n702), .S(N11), .Z(n704) );
  MUX2_X1 U790 ( .A(n704), .B(n701), .S(n891), .Z(N44) );
  MUX2_X1 U791 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n895), .Z(n705) );
  MUX2_X1 U792 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n895), .Z(n706) );
  MUX2_X1 U793 ( .A(n706), .B(n705), .S(n893), .Z(n707) );
  MUX2_X1 U794 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n900), .Z(n708) );
  MUX2_X1 U795 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n898), .Z(n709) );
  MUX2_X1 U796 ( .A(n709), .B(n708), .S(N11), .Z(n710) );
  MUX2_X1 U797 ( .A(n710), .B(n707), .S(n891), .Z(N43) );
  MUX2_X1 U798 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n897), .Z(n711) );
  MUX2_X1 U799 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n897), .Z(n712) );
  MUX2_X1 U800 ( .A(n712), .B(n711), .S(n892), .Z(n713) );
  MUX2_X1 U801 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n897), .Z(n714) );
  MUX2_X1 U802 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n897), .Z(n715) );
  MUX2_X1 U803 ( .A(n715), .B(n714), .S(n892), .Z(n716) );
  MUX2_X1 U804 ( .A(n716), .B(n713), .S(n891), .Z(N42) );
  MUX2_X1 U805 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n897), .Z(n717) );
  MUX2_X1 U806 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n897), .Z(n718) );
  MUX2_X1 U807 ( .A(n718), .B(n717), .S(n893), .Z(n719) );
  MUX2_X1 U808 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n897), .Z(n720) );
  MUX2_X1 U809 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n897), .Z(n721) );
  MUX2_X1 U810 ( .A(n721), .B(n720), .S(n894), .Z(n722) );
  MUX2_X1 U811 ( .A(n722), .B(n719), .S(n891), .Z(N41) );
  MUX2_X1 U812 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n897), .Z(n723) );
  MUX2_X1 U813 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n897), .Z(n724) );
  MUX2_X1 U814 ( .A(n724), .B(n723), .S(n892), .Z(n725) );
  MUX2_X1 U815 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n897), .Z(n726) );
  MUX2_X1 U816 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n897), .Z(n727) );
  MUX2_X1 U817 ( .A(n727), .B(n726), .S(N11), .Z(n728) );
  MUX2_X1 U818 ( .A(n728), .B(n725), .S(n891), .Z(N40) );
  MUX2_X1 U819 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n896), .Z(n729) );
  MUX2_X1 U820 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n900), .Z(n730) );
  MUX2_X1 U821 ( .A(n730), .B(n729), .S(n894), .Z(n731) );
  MUX2_X1 U822 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n901), .Z(n732) );
  MUX2_X1 U823 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(N10), .Z(n733) );
  MUX2_X1 U824 ( .A(n733), .B(n732), .S(n892), .Z(n734) );
  MUX2_X1 U825 ( .A(n734), .B(n731), .S(n891), .Z(N39) );
  MUX2_X1 U826 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n901), .Z(n735) );
  MUX2_X1 U827 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n901), .Z(n736) );
  MUX2_X1 U828 ( .A(n736), .B(n735), .S(n893), .Z(n737) );
  MUX2_X1 U829 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n895), .Z(n738) );
  MUX2_X1 U830 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(N10), .Z(n739) );
  MUX2_X1 U831 ( .A(n739), .B(n738), .S(n893), .Z(n740) );
  MUX2_X1 U832 ( .A(n740), .B(n737), .S(n891), .Z(N38) );
  MUX2_X1 U833 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(N10), .Z(n741) );
  MUX2_X1 U834 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n901), .Z(n742) );
  MUX2_X1 U835 ( .A(n742), .B(n741), .S(n892), .Z(n743) );
  MUX2_X1 U836 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(N10), .Z(n744) );
  MUX2_X1 U837 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(N10), .Z(n745) );
  MUX2_X1 U838 ( .A(n745), .B(n744), .S(N11), .Z(n746) );
  MUX2_X1 U839 ( .A(n746), .B(n743), .S(n891), .Z(N37) );
  MUX2_X1 U840 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(N10), .Z(n747) );
  MUX2_X1 U841 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n900), .Z(n748) );
  MUX2_X1 U842 ( .A(n748), .B(n747), .S(n893), .Z(n749) );
  MUX2_X1 U843 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n901), .Z(n750) );
  MUX2_X1 U844 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n901), .Z(n751) );
  MUX2_X1 U845 ( .A(n751), .B(n750), .S(n894), .Z(n752) );
  MUX2_X1 U846 ( .A(n752), .B(n749), .S(n891), .Z(N36) );
  MUX2_X1 U847 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n896), .Z(n753) );
  MUX2_X1 U848 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n901), .Z(n754) );
  MUX2_X1 U849 ( .A(n754), .B(n753), .S(n894), .Z(n755) );
  MUX2_X1 U850 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n900), .Z(n756) );
  MUX2_X1 U851 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n900), .Z(n757) );
  MUX2_X1 U852 ( .A(n757), .B(n756), .S(N11), .Z(n758) );
  MUX2_X1 U853 ( .A(n758), .B(n755), .S(N12), .Z(N35) );
  MUX2_X1 U854 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n900), .Z(n759) );
  MUX2_X1 U855 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n900), .Z(n760) );
  MUX2_X1 U856 ( .A(n760), .B(n759), .S(n894), .Z(n761) );
  MUX2_X1 U857 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(N10), .Z(n762) );
  MUX2_X1 U858 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n900), .Z(n763) );
  MUX2_X1 U859 ( .A(n763), .B(n762), .S(n893), .Z(n764) );
  MUX2_X1 U860 ( .A(n764), .B(n761), .S(N12), .Z(N34) );
  MUX2_X1 U861 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(N10), .Z(n765) );
  MUX2_X1 U862 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n901), .Z(n766) );
  MUX2_X1 U863 ( .A(n766), .B(n765), .S(n893), .Z(n767) );
  MUX2_X1 U864 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n900), .Z(n768) );
  MUX2_X1 U865 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n900), .Z(n769) );
  MUX2_X1 U866 ( .A(n769), .B(n768), .S(n894), .Z(n770) );
  MUX2_X1 U867 ( .A(n770), .B(n767), .S(N12), .Z(N33) );
  MUX2_X1 U868 ( .A(\mem[6][20] ), .B(\mem[7][20] ), .S(N10), .Z(n771) );
  MUX2_X1 U869 ( .A(\mem[4][20] ), .B(\mem[5][20] ), .S(n900), .Z(n772) );
  MUX2_X1 U870 ( .A(n772), .B(n771), .S(n892), .Z(n773) );
  MUX2_X1 U871 ( .A(\mem[2][20] ), .B(\mem[3][20] ), .S(n900), .Z(n774) );
  MUX2_X1 U872 ( .A(\mem[0][20] ), .B(\mem[1][20] ), .S(n901), .Z(n775) );
  MUX2_X1 U873 ( .A(n775), .B(n774), .S(N11), .Z(n776) );
  MUX2_X1 U874 ( .A(n776), .B(n773), .S(N12), .Z(N32) );
  MUX2_X1 U875 ( .A(\mem[6][21] ), .B(\mem[7][21] ), .S(n900), .Z(n777) );
  MUX2_X1 U876 ( .A(\mem[4][21] ), .B(\mem[5][21] ), .S(n900), .Z(n778) );
  MUX2_X1 U877 ( .A(n778), .B(n777), .S(n893), .Z(n779) );
  MUX2_X1 U878 ( .A(\mem[2][21] ), .B(\mem[3][21] ), .S(n901), .Z(n780) );
  MUX2_X1 U879 ( .A(\mem[0][21] ), .B(\mem[1][21] ), .S(n901), .Z(n781) );
  MUX2_X1 U880 ( .A(n781), .B(n780), .S(N11), .Z(n782) );
  MUX2_X1 U881 ( .A(n782), .B(n779), .S(N12), .Z(N31) );
  MUX2_X1 U882 ( .A(\mem[6][22] ), .B(\mem[7][22] ), .S(n896), .Z(n783) );
  MUX2_X1 U883 ( .A(\mem[4][22] ), .B(\mem[5][22] ), .S(n897), .Z(n784) );
  MUX2_X1 U884 ( .A(n784), .B(n783), .S(n892), .Z(n785) );
  MUX2_X1 U885 ( .A(\mem[2][22] ), .B(\mem[3][22] ), .S(n898), .Z(n786) );
  MUX2_X1 U886 ( .A(\mem[0][22] ), .B(\mem[1][22] ), .S(n896), .Z(n787) );
  MUX2_X1 U887 ( .A(n787), .B(n786), .S(n892), .Z(n788) );
  MUX2_X1 U888 ( .A(n788), .B(n785), .S(N12), .Z(N30) );
  MUX2_X1 U889 ( .A(\mem[6][23] ), .B(\mem[7][23] ), .S(n897), .Z(n789) );
  MUX2_X1 U890 ( .A(\mem[4][23] ), .B(\mem[5][23] ), .S(n898), .Z(n790) );
  MUX2_X1 U891 ( .A(n790), .B(n789), .S(n892), .Z(n791) );
  MUX2_X1 U892 ( .A(\mem[2][23] ), .B(\mem[3][23] ), .S(n899), .Z(n792) );
  MUX2_X1 U893 ( .A(\mem[0][23] ), .B(\mem[1][23] ), .S(n895), .Z(n793) );
  MUX2_X1 U894 ( .A(n793), .B(n792), .S(n892), .Z(n794) );
  MUX2_X1 U895 ( .A(n794), .B(n791), .S(N12), .Z(N29) );
  MUX2_X1 U896 ( .A(\mem[6][24] ), .B(\mem[7][24] ), .S(n897), .Z(n795) );
  MUX2_X1 U897 ( .A(\mem[4][24] ), .B(\mem[5][24] ), .S(n899), .Z(n796) );
  MUX2_X1 U898 ( .A(n796), .B(n795), .S(n892), .Z(n797) );
  MUX2_X1 U899 ( .A(\mem[2][24] ), .B(\mem[3][24] ), .S(n896), .Z(n798) );
  MUX2_X1 U900 ( .A(\mem[0][24] ), .B(\mem[1][24] ), .S(n897), .Z(n799) );
  MUX2_X1 U901 ( .A(n799), .B(n798), .S(n892), .Z(n800) );
  MUX2_X1 U902 ( .A(n800), .B(n797), .S(N12), .Z(N28) );
  MUX2_X1 U903 ( .A(\mem[6][25] ), .B(\mem[7][25] ), .S(n898), .Z(n801) );
  MUX2_X1 U904 ( .A(\mem[4][25] ), .B(\mem[5][25] ), .S(n896), .Z(n802) );
  MUX2_X1 U905 ( .A(n802), .B(n801), .S(n892), .Z(n803) );
  MUX2_X1 U906 ( .A(\mem[2][25] ), .B(\mem[3][25] ), .S(n898), .Z(n804) );
  MUX2_X1 U907 ( .A(\mem[0][25] ), .B(\mem[1][25] ), .S(n898), .Z(n805) );
  MUX2_X1 U908 ( .A(n805), .B(n804), .S(n892), .Z(n806) );
  MUX2_X1 U909 ( .A(n806), .B(n803), .S(N12), .Z(N27) );
  MUX2_X1 U910 ( .A(\mem[6][26] ), .B(\mem[7][26] ), .S(n901), .Z(n807) );
  MUX2_X1 U911 ( .A(\mem[4][26] ), .B(\mem[5][26] ), .S(n895), .Z(n808) );
  MUX2_X1 U912 ( .A(n808), .B(n807), .S(n892), .Z(n809) );
  MUX2_X1 U913 ( .A(\mem[2][26] ), .B(\mem[3][26] ), .S(n900), .Z(n810) );
  MUX2_X1 U914 ( .A(\mem[0][26] ), .B(\mem[1][26] ), .S(n897), .Z(n811) );
  MUX2_X1 U915 ( .A(n811), .B(n810), .S(n892), .Z(n812) );
  MUX2_X1 U916 ( .A(n812), .B(n809), .S(N12), .Z(N26) );
  MUX2_X1 U917 ( .A(\mem[6][27] ), .B(\mem[7][27] ), .S(n895), .Z(n813) );
  MUX2_X1 U918 ( .A(\mem[4][27] ), .B(\mem[5][27] ), .S(n900), .Z(n814) );
  MUX2_X1 U919 ( .A(n814), .B(n813), .S(n892), .Z(n815) );
  MUX2_X1 U920 ( .A(\mem[2][27] ), .B(\mem[3][27] ), .S(n897), .Z(n816) );
  MUX2_X1 U921 ( .A(\mem[0][27] ), .B(\mem[1][27] ), .S(n899), .Z(n817) );
  MUX2_X1 U922 ( .A(n817), .B(n816), .S(n892), .Z(n818) );
  MUX2_X1 U923 ( .A(n818), .B(n815), .S(N12), .Z(N25) );
  MUX2_X1 U924 ( .A(\mem[6][28] ), .B(\mem[7][28] ), .S(n897), .Z(n819) );
  MUX2_X1 U925 ( .A(\mem[4][28] ), .B(\mem[5][28] ), .S(n896), .Z(n820) );
  MUX2_X1 U926 ( .A(n820), .B(n819), .S(n893), .Z(n821) );
  MUX2_X1 U927 ( .A(\mem[2][28] ), .B(\mem[3][28] ), .S(n897), .Z(n822) );
  MUX2_X1 U928 ( .A(\mem[0][28] ), .B(\mem[1][28] ), .S(n899), .Z(n823) );
  MUX2_X1 U929 ( .A(n823), .B(n822), .S(n893), .Z(n824) );
  MUX2_X1 U930 ( .A(n824), .B(n821), .S(n891), .Z(N24) );
  MUX2_X1 U931 ( .A(\mem[6][29] ), .B(\mem[7][29] ), .S(n899), .Z(n825) );
  MUX2_X1 U932 ( .A(\mem[4][29] ), .B(\mem[5][29] ), .S(n900), .Z(n826) );
  MUX2_X1 U933 ( .A(n826), .B(n825), .S(n893), .Z(n827) );
  MUX2_X1 U934 ( .A(\mem[2][29] ), .B(\mem[3][29] ), .S(n899), .Z(n828) );
  MUX2_X1 U935 ( .A(\mem[0][29] ), .B(\mem[1][29] ), .S(n896), .Z(n829) );
  MUX2_X1 U936 ( .A(n829), .B(n828), .S(n893), .Z(n830) );
  MUX2_X1 U937 ( .A(n830), .B(n827), .S(n891), .Z(N23) );
  MUX2_X1 U938 ( .A(\mem[6][30] ), .B(\mem[7][30] ), .S(n898), .Z(n831) );
  MUX2_X1 U939 ( .A(\mem[4][30] ), .B(\mem[5][30] ), .S(n897), .Z(n832) );
  MUX2_X1 U940 ( .A(n832), .B(n831), .S(n893), .Z(n833) );
  MUX2_X1 U941 ( .A(\mem[2][30] ), .B(\mem[3][30] ), .S(n901), .Z(n834) );
  MUX2_X1 U942 ( .A(\mem[0][30] ), .B(\mem[1][30] ), .S(n898), .Z(n835) );
  MUX2_X1 U943 ( .A(n835), .B(n834), .S(n893), .Z(n836) );
  MUX2_X1 U944 ( .A(n836), .B(n833), .S(n891), .Z(N22) );
  MUX2_X1 U945 ( .A(\mem[6][31] ), .B(\mem[7][31] ), .S(n898), .Z(n837) );
  MUX2_X1 U946 ( .A(\mem[4][31] ), .B(\mem[5][31] ), .S(n898), .Z(n838) );
  MUX2_X1 U947 ( .A(n838), .B(n837), .S(n893), .Z(n839) );
  MUX2_X1 U948 ( .A(\mem[2][31] ), .B(\mem[3][31] ), .S(n898), .Z(n840) );
  MUX2_X1 U949 ( .A(\mem[0][31] ), .B(\mem[1][31] ), .S(n898), .Z(n841) );
  MUX2_X1 U950 ( .A(n841), .B(n840), .S(n893), .Z(n842) );
  MUX2_X1 U951 ( .A(n842), .B(n839), .S(n891), .Z(N21) );
  MUX2_X1 U952 ( .A(\mem[6][32] ), .B(\mem[7][32] ), .S(n898), .Z(n843) );
  MUX2_X1 U953 ( .A(\mem[4][32] ), .B(\mem[5][32] ), .S(n898), .Z(n844) );
  MUX2_X1 U954 ( .A(n844), .B(n843), .S(n893), .Z(n845) );
  MUX2_X1 U955 ( .A(\mem[2][32] ), .B(\mem[3][32] ), .S(n898), .Z(n846) );
  MUX2_X1 U956 ( .A(\mem[0][32] ), .B(\mem[1][32] ), .S(n898), .Z(n847) );
  MUX2_X1 U957 ( .A(n847), .B(n846), .S(n893), .Z(n848) );
  MUX2_X1 U958 ( .A(n848), .B(n845), .S(n891), .Z(N20) );
  MUX2_X1 U959 ( .A(\mem[6][33] ), .B(\mem[7][33] ), .S(n898), .Z(n849) );
  MUX2_X1 U960 ( .A(\mem[4][33] ), .B(\mem[5][33] ), .S(n898), .Z(n850) );
  MUX2_X1 U961 ( .A(n850), .B(n849), .S(n893), .Z(n851) );
  MUX2_X1 U962 ( .A(\mem[2][33] ), .B(\mem[3][33] ), .S(n898), .Z(n852) );
  MUX2_X1 U963 ( .A(\mem[0][33] ), .B(\mem[1][33] ), .S(n898), .Z(n853) );
  MUX2_X1 U964 ( .A(n853), .B(n852), .S(n893), .Z(n854) );
  MUX2_X1 U965 ( .A(n854), .B(n851), .S(n891), .Z(N19) );
  MUX2_X1 U966 ( .A(\mem[6][34] ), .B(\mem[7][34] ), .S(n899), .Z(n855) );
  MUX2_X1 U967 ( .A(\mem[4][34] ), .B(\mem[5][34] ), .S(n899), .Z(n856) );
  MUX2_X1 U968 ( .A(n856), .B(n855), .S(n894), .Z(n857) );
  MUX2_X1 U969 ( .A(\mem[2][34] ), .B(\mem[3][34] ), .S(n899), .Z(n858) );
  MUX2_X1 U970 ( .A(\mem[0][34] ), .B(\mem[1][34] ), .S(n899), .Z(n859) );
  MUX2_X1 U971 ( .A(n859), .B(n858), .S(n894), .Z(n860) );
  MUX2_X1 U972 ( .A(n860), .B(n857), .S(N12), .Z(N18) );
  MUX2_X1 U973 ( .A(\mem[6][35] ), .B(\mem[7][35] ), .S(n899), .Z(n861) );
  MUX2_X1 U974 ( .A(\mem[4][35] ), .B(\mem[5][35] ), .S(n899), .Z(n862) );
  MUX2_X1 U975 ( .A(n862), .B(n861), .S(n894), .Z(n863) );
  MUX2_X1 U976 ( .A(\mem[2][35] ), .B(\mem[3][35] ), .S(n899), .Z(n864) );
  MUX2_X1 U977 ( .A(\mem[0][35] ), .B(\mem[1][35] ), .S(n899), .Z(n865) );
  MUX2_X1 U978 ( .A(n865), .B(n864), .S(n894), .Z(n866) );
  MUX2_X1 U979 ( .A(n866), .B(n863), .S(N12), .Z(N17) );
  MUX2_X1 U980 ( .A(\mem[6][36] ), .B(\mem[7][36] ), .S(n899), .Z(n867) );
  MUX2_X1 U981 ( .A(\mem[4][36] ), .B(\mem[5][36] ), .S(n899), .Z(n868) );
  MUX2_X1 U982 ( .A(n868), .B(n867), .S(n894), .Z(n869) );
  MUX2_X1 U983 ( .A(\mem[2][36] ), .B(\mem[3][36] ), .S(n899), .Z(n870) );
  MUX2_X1 U984 ( .A(\mem[0][36] ), .B(\mem[1][36] ), .S(n899), .Z(n871) );
  MUX2_X1 U985 ( .A(n871), .B(n870), .S(n894), .Z(n872) );
  MUX2_X1 U986 ( .A(n872), .B(n869), .S(N12), .Z(N16) );
  MUX2_X1 U987 ( .A(\mem[6][37] ), .B(\mem[7][37] ), .S(n899), .Z(n873) );
  MUX2_X1 U988 ( .A(\mem[4][37] ), .B(\mem[5][37] ), .S(n898), .Z(n874) );
  MUX2_X1 U989 ( .A(n874), .B(n873), .S(n894), .Z(n875) );
  MUX2_X1 U990 ( .A(\mem[2][37] ), .B(\mem[3][37] ), .S(n899), .Z(n876) );
  MUX2_X1 U991 ( .A(\mem[0][37] ), .B(\mem[1][37] ), .S(n897), .Z(n877) );
  MUX2_X1 U992 ( .A(n877), .B(n876), .S(n894), .Z(n878) );
  MUX2_X1 U993 ( .A(n878), .B(n875), .S(N12), .Z(N15) );
  MUX2_X1 U994 ( .A(\mem[6][38] ), .B(\mem[7][38] ), .S(n901), .Z(n879) );
  MUX2_X1 U995 ( .A(\mem[4][38] ), .B(\mem[5][38] ), .S(n899), .Z(n880) );
  MUX2_X1 U996 ( .A(n880), .B(n879), .S(n894), .Z(n881) );
  MUX2_X1 U997 ( .A(\mem[2][38] ), .B(\mem[3][38] ), .S(n895), .Z(n882) );
  MUX2_X1 U998 ( .A(\mem[0][38] ), .B(\mem[1][38] ), .S(n898), .Z(n883) );
  MUX2_X1 U999 ( .A(n883), .B(n882), .S(n894), .Z(n884) );
  MUX2_X1 U1000 ( .A(n884), .B(n881), .S(N12), .Z(N14) );
  MUX2_X1 U1001 ( .A(\mem[6][39] ), .B(\mem[7][39] ), .S(n895), .Z(n885) );
  MUX2_X1 U1002 ( .A(\mem[4][39] ), .B(\mem[5][39] ), .S(n895), .Z(n886) );
  MUX2_X1 U1003 ( .A(n886), .B(n885), .S(n894), .Z(n887) );
  MUX2_X1 U1004 ( .A(\mem[2][39] ), .B(\mem[3][39] ), .S(n896), .Z(n888) );
  MUX2_X1 U1005 ( .A(\mem[0][39] ), .B(\mem[1][39] ), .S(n899), .Z(n889) );
  MUX2_X1 U1006 ( .A(n889), .B(n888), .S(n894), .Z(n890) );
  MUX2_X1 U1007 ( .A(n890), .B(n887), .S(N12), .Z(N13) );
  CLKBUF_X1 U1008 ( .A(n900), .Z(n895) );
  CLKBUF_X1 U1009 ( .A(n333), .Z(n904) );
  CLKBUF_X1 U1010 ( .A(n127), .Z(n919) );
endmodule


module datapath_DW_mult_tc_8 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n15, n16, n17, n18,
         n19, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34, n35,
         n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n51, n52,
         n53, n54, n55, n57, n58, n59, n60, n61, n63, n64, n65, n67, n68, n69,
         n82, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n105, n106, n107, n108, n109,
         n111, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n124, n126, n127, n128, n129, n130, n131, n134, n135, n136, n137,
         n139, n141, n142, n143, n144, n145, n146, n149, n150, n151, n152,
         n154, n156, n157, n158, n159, n160, n161, n165, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n190, n191, n192, n193,
         n195, n197, n198, n199, n200, n201, n202, n206, n208, n209, n210,
         n211, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n256, n257, n258, n259, n260, n261, n262, n263, n267, n268,
         n269, n270, n271, n273, n274, n275, n276, n277, n278, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n303, n304,
         n305, n306, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n329,
         n331, n332, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n344, n346, n347, n348, n349, n350, n351, n352, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n371, n373, n374, n376, n378, n379, n380, n382, n384,
         n385, n386, n387, n388, n390, n392, n393, n394, n395, n396, n398,
         n400, n401, n402, n403, n404, n405, n406, n407, n409, n418, n424,
         n427, n430, n434, n435, n436, n437, n441, n443, n445, n446, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n793, n794, n796, n797, n799, n800, n802, n803, n805,
         n806, n808, n809, n811, n812, n814, n815, n817, n818, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1484, n1485, n1486, n1487, n1488, n1489, n1490;
  assign product[39] = n105;

  FA_X1 U488 ( .A(n831), .B(n454), .CI(n850), .CO(n450), .S(n451) );
  FA_X1 U489 ( .A(n455), .B(n832), .CI(n458), .CO(n452), .S(n453) );
  FA_X1 U491 ( .A(n462), .B(n833), .CI(n459), .CO(n456), .S(n457) );
  FA_X1 U492 ( .A(n851), .B(n464), .CI(n870), .CO(n458), .S(n459) );
  FA_X1 U493 ( .A(n463), .B(n470), .CI(n468), .CO(n460), .S(n461) );
  FA_X1 U494 ( .A(n834), .B(n852), .CI(n465), .CO(n462), .S(n463) );
  FA_X1 U496 ( .A(n474), .B(n471), .CI(n469), .CO(n466), .S(n467) );
  FA_X1 U497 ( .A(n478), .B(n871), .CI(n476), .CO(n468), .S(n469) );
  FA_X1 U498 ( .A(n853), .B(n835), .CI(n890), .CO(n470), .S(n471) );
  FA_X1 U499 ( .A(n475), .B(n477), .CI(n482), .CO(n472), .S(n473) );
  FA_X1 U500 ( .A(n486), .B(n479), .CI(n484), .CO(n474), .S(n475) );
  FA_X1 U501 ( .A(n836), .B(n854), .CI(n872), .CO(n476), .S(n477) );
  FA_X1 U503 ( .A(n490), .B(n492), .CI(n483), .CO(n480), .S(n481) );
  FA_X1 U504 ( .A(n485), .B(n494), .CI(n487), .CO(n482), .S(n483) );
  FA_X1 U505 ( .A(n855), .B(n496), .CI(n873), .CO(n484), .S(n485) );
  FA_X1 U506 ( .A(n891), .B(n837), .CI(n910), .CO(n486), .S(n487) );
  FA_X1 U507 ( .A(n500), .B(n493), .CI(n491), .CO(n488), .S(n489) );
  FA_X1 U508 ( .A(n495), .B(n504), .CI(n502), .CO(n490), .S(n491) );
  FA_X1 U509 ( .A(n497), .B(n874), .CI(n506), .CO(n492), .S(n493) );
  FA_X1 U510 ( .A(n892), .B(n856), .CI(n838), .CO(n494), .S(n495) );
  FA_X1 U512 ( .A(n510), .B(n503), .CI(n501), .CO(n498), .S(n499) );
  FA_X1 U513 ( .A(n507), .B(n505), .CI(n512), .CO(n500), .S(n501) );
  FA_X1 U514 ( .A(n516), .B(n893), .CI(n514), .CO(n502), .S(n503) );
  FA_X1 U515 ( .A(n857), .B(n911), .CI(n875), .CO(n504), .S(n505) );
  FA_X1 U516 ( .A(n518), .B(n839), .CI(n930), .CO(n506), .S(n507) );
  FA_X1 U517 ( .A(n522), .B(n513), .CI(n511), .CO(n508), .S(n509) );
  FA_X1 U518 ( .A(n526), .B(n515), .CI(n524), .CO(n510), .S(n511) );
  FA_X1 U519 ( .A(n528), .B(n530), .CI(n517), .CO(n512), .S(n513) );
  FA_X1 U520 ( .A(n840), .B(n858), .CI(n519), .CO(n514), .S(n515) );
  FA_X1 U521 ( .A(n912), .B(n876), .CI(n894), .CO(n516), .S(n517) );
  FA_X1 U523 ( .A(n525), .B(n534), .CI(n523), .CO(n520), .S(n521) );
  FA_X1 U524 ( .A(n527), .B(n538), .CI(n536), .CO(n522), .S(n523) );
  FA_X1 U525 ( .A(n529), .B(n540), .CI(n531), .CO(n524), .S(n525) );
  FA_X1 U526 ( .A(n877), .B(n895), .CI(n542), .CO(n526), .S(n527) );
  FA_X1 U527 ( .A(n859), .B(n931), .CI(n913), .CO(n528), .S(n529) );
  FA_X1 U528 ( .A(n544), .B(n841), .CI(n950), .CO(n530), .S(n531) );
  FA_X1 U529 ( .A(n535), .B(n537), .CI(n548), .CO(n532), .S(n533) );
  FA_X1 U530 ( .A(n539), .B(n552), .CI(n550), .CO(n534), .S(n535) );
  FA_X1 U531 ( .A(n541), .B(n554), .CI(n543), .CO(n536), .S(n537) );
  FA_X1 U532 ( .A(n558), .B(n545), .CI(n556), .CO(n538), .S(n539) );
  FA_X1 U533 ( .A(n896), .B(n932), .CI(n914), .CO(n540), .S(n541) );
  FA_X1 U534 ( .A(n842), .B(n878), .CI(n860), .CO(n542), .S(n543) );
  FA_X1 U536 ( .A(n562), .B(n551), .CI(n549), .CO(n546), .S(n547) );
  FA_X1 U537 ( .A(n553), .B(n566), .CI(n564), .CO(n548), .S(n549) );
  FA_X1 U538 ( .A(n559), .B(n557), .CI(n568), .CO(n550), .S(n551) );
  FA_X1 U539 ( .A(n570), .B(n572), .CI(n555), .CO(n552), .S(n553) );
  FA_X1 U540 ( .A(n879), .B(n915), .CI(n897), .CO(n554), .S(n555) );
  FA_X1 U541 ( .A(n861), .B(n951), .CI(n933), .CO(n556), .S(n557) );
  FA_X1 U542 ( .A(n574), .B(n843), .CI(n970), .CO(n558), .S(n559) );
  FA_X1 U543 ( .A(n578), .B(n565), .CI(n563), .CO(n560), .S(n561) );
  FA_X1 U544 ( .A(n567), .B(n582), .CI(n580), .CO(n562), .S(n563) );
  FA_X1 U545 ( .A(n584), .B(n573), .CI(n569), .CO(n564), .S(n565) );
  FA_X1 U546 ( .A(n586), .B(n588), .CI(n571), .CO(n566), .S(n567) );
  FA_X1 U547 ( .A(n575), .B(n898), .CI(n590), .CO(n568), .S(n569) );
  FA_X1 U548 ( .A(n844), .B(n916), .CI(n862), .CO(n570), .S(n571) );
  FA_X1 U549 ( .A(n952), .B(n880), .CI(n934), .CO(n572), .S(n573) );
  FA_X1 U551 ( .A(n594), .B(n581), .CI(n579), .CO(n576), .S(n577) );
  FA_X1 U552 ( .A(n583), .B(n598), .CI(n596), .CO(n578), .S(n579) );
  FA_X1 U553 ( .A(n600), .B(n591), .CI(n585), .CO(n580), .S(n581) );
  FA_X1 U554 ( .A(n587), .B(n602), .CI(n589), .CO(n582), .S(n583) );
  FA_X1 U555 ( .A(n606), .B(n917), .CI(n604), .CO(n584), .S(n585) );
  FA_X1 U556 ( .A(n881), .B(n935), .CI(n899), .CO(n586), .S(n587) );
  FA_X1 U557 ( .A(n608), .B(n953), .CI(n863), .CO(n588), .S(n589) );
  FA_X1 U558 ( .A(n845), .B(n971), .CI(n990), .CO(n590), .S(n591) );
  FA_X1 U559 ( .A(n612), .B(n597), .CI(n595), .CO(n592), .S(n593) );
  FA_X1 U560 ( .A(n599), .B(n616), .CI(n614), .CO(n594), .S(n595) );
  FA_X1 U561 ( .A(n618), .B(n603), .CI(n601), .CO(n596), .S(n597) );
  FA_X1 U562 ( .A(n605), .B(n620), .CI(n607), .CO(n598), .S(n599) );
  FA_X1 U563 ( .A(n624), .B(n626), .CI(n622), .CO(n600), .S(n601) );
  FA_X1 U564 ( .A(n918), .B(n936), .CI(n609), .CO(n602), .S(n603) );
  FA_X1 U565 ( .A(n954), .B(n864), .CI(n882), .CO(n604), .S(n605) );
  FA_X1 U566 ( .A(n972), .B(n846), .CI(n900), .CO(n606), .S(n607) );
  FA_X1 U569 ( .A(n617), .B(n634), .CI(n632), .CO(n612), .S(n613) );
  FA_X1 U570 ( .A(n636), .B(n621), .CI(n619), .CO(n614), .S(n615) );
  FA_X1 U571 ( .A(n623), .B(n638), .CI(n625), .CO(n616), .S(n617) );
  FA_X1 U572 ( .A(n642), .B(n627), .CI(n640), .CO(n618), .S(n619) );
  FA_X1 U573 ( .A(n955), .B(n973), .CI(n644), .CO(n620), .S(n621) );
  FA_X1 U574 ( .A(n991), .B(n901), .CI(n883), .CO(n622), .S(n623) );
  FA_X1 U575 ( .A(n919), .B(n847), .CI(n1010), .CO(n624), .S(n625) );
  FA_X1 U578 ( .A(n648), .B(n633), .CI(n631), .CO(n628), .S(n629) );
  FA_X1 U579 ( .A(n650), .B(n637), .CI(n635), .CO(n630), .S(n631) );
  FA_X1 U580 ( .A(n654), .B(n643), .CI(n652), .CO(n632), .S(n633) );
  FA_X1 U581 ( .A(n639), .B(n656), .CI(n641), .CO(n634), .S(n635) );
  FA_X1 U582 ( .A(n660), .B(n645), .CI(n658), .CO(n636), .S(n637) );
  FA_X1 U583 ( .A(n920), .B(n992), .CI(n974), .CO(n638), .S(n639) );
  FA_X1 U584 ( .A(n1011), .B(n956), .CI(n902), .CO(n640), .S(n641) );
  FA_X1 U585 ( .A(n866), .B(n884), .CI(n938), .CO(n642), .S(n643) );
  HA_X1 U586 ( .A(n820), .B(n848), .CO(n644), .S(n645) );
  FA_X1 U587 ( .A(n664), .B(n651), .CI(n649), .CO(n646), .S(n647) );
  FA_X1 U588 ( .A(n653), .B(n655), .CI(n666), .CO(n648), .S(n649) );
  FA_X1 U589 ( .A(n670), .B(n659), .CI(n668), .CO(n650), .S(n651) );
  FA_X1 U590 ( .A(n661), .B(n672), .CI(n657), .CO(n652), .S(n653) );
  FA_X1 U591 ( .A(n676), .B(n957), .CI(n674), .CO(n654), .S(n655) );
  FA_X1 U592 ( .A(n921), .B(n975), .CI(n939), .CO(n656), .S(n657) );
  FA_X1 U593 ( .A(n867), .B(n993), .CI(n903), .CO(n658), .S(n659) );
  FA_X1 U594 ( .A(n849), .B(n885), .CI(n1012), .CO(n660), .S(n661) );
  FA_X1 U595 ( .A(n667), .B(n680), .CI(n665), .CO(n662), .S(n663) );
  FA_X1 U596 ( .A(n669), .B(n671), .CI(n682), .CO(n664), .S(n665) );
  FA_X1 U597 ( .A(n675), .B(n673), .CI(n684), .CO(n666), .S(n667) );
  FA_X1 U598 ( .A(n686), .B(n690), .CI(n688), .CO(n668), .S(n669) );
  FA_X1 U599 ( .A(n958), .B(n976), .CI(n677), .CO(n670), .S(n671) );
  FA_X1 U600 ( .A(n886), .B(n904), .CI(n922), .CO(n672), .S(n673) );
  FA_X1 U601 ( .A(n1013), .B(n940), .CI(n994), .CO(n674), .S(n675) );
  HA_X1 U602 ( .A(n821), .B(n868), .CO(n676), .S(n677) );
  FA_X1 U603 ( .A(n694), .B(n683), .CI(n681), .CO(n678), .S(n679) );
  FA_X1 U604 ( .A(n698), .B(n696), .CI(n685), .CO(n680), .S(n681) );
  FA_X1 U605 ( .A(n689), .B(n691), .CI(n687), .CO(n682), .S(n683) );
  FA_X1 U606 ( .A(n702), .B(n704), .CI(n700), .CO(n684), .S(n685) );
  FA_X1 U607 ( .A(n959), .B(n977), .CI(n941), .CO(n686), .S(n687) );
  FA_X1 U608 ( .A(n887), .B(n995), .CI(n923), .CO(n688), .S(n689) );
  FA_X1 U609 ( .A(n1014), .B(n869), .CI(n905), .CO(n690), .S(n691) );
  FA_X1 U610 ( .A(n697), .B(n708), .CI(n695), .CO(n692), .S(n693) );
  FA_X1 U611 ( .A(n710), .B(n703), .CI(n699), .CO(n694), .S(n695) );
  FA_X1 U613 ( .A(n716), .B(n996), .CI(n705), .CO(n698), .S(n699) );
  FA_X1 U614 ( .A(n1015), .B(n942), .CI(n978), .CO(n700), .S(n701) );
  HA_X1 U616 ( .A(n822), .B(n888), .CO(n704), .S(n705) );
  FA_X1 U617 ( .A(n711), .B(n720), .CI(n709), .CO(n706), .S(n707) );
  FA_X1 U618 ( .A(n713), .B(n715), .CI(n722), .CO(n708), .S(n709) );
  FA_X1 U619 ( .A(n724), .B(n726), .CI(n717), .CO(n710), .S(n711) );
  FA_X1 U620 ( .A(n961), .B(n979), .CI(n728), .CO(n712), .S(n713) );
  FA_X1 U621 ( .A(n907), .B(n997), .CI(n943), .CO(n714), .S(n715) );
  FA_X1 U622 ( .A(n1016), .B(n889), .CI(n925), .CO(n716), .S(n717) );
  FA_X1 U623 ( .A(n732), .B(n723), .CI(n721), .CO(n718), .S(n719) );
  FA_X1 U624 ( .A(n727), .B(n725), .CI(n734), .CO(n720), .S(n721) );
  FA_X1 U625 ( .A(n738), .B(n729), .CI(n736), .CO(n722), .S(n723) );
  FA_X1 U626 ( .A(n926), .B(n980), .CI(n944), .CO(n724), .S(n725) );
  FA_X1 U627 ( .A(n1017), .B(n962), .CI(n998), .CO(n726), .S(n727) );
  HA_X1 U628 ( .A(n908), .B(n823), .CO(n728), .S(n729) );
  FA_X1 U629 ( .A(n735), .B(n742), .CI(n733), .CO(n730), .S(n731) );
  FA_X1 U630 ( .A(n737), .B(n739), .CI(n744), .CO(n732), .S(n733) );
  FA_X1 U631 ( .A(n748), .B(n981), .CI(n746), .CO(n734), .S(n735) );
  FA_X1 U632 ( .A(n927), .B(n999), .CI(n963), .CO(n736), .S(n737) );
  FA_X1 U633 ( .A(n1018), .B(n909), .CI(n945), .CO(n738), .S(n739) );
  FA_X1 U634 ( .A(n752), .B(n745), .CI(n743), .CO(n740), .S(n741) );
  FA_X1 U635 ( .A(n754), .B(n756), .CI(n747), .CO(n742), .S(n743) );
  FA_X1 U636 ( .A(n964), .B(n1000), .CI(n749), .CO(n744), .S(n745) );
  FA_X1 U637 ( .A(n946), .B(n982), .CI(n1019), .CO(n746), .S(n747) );
  HA_X1 U638 ( .A(n824), .B(n928), .CO(n748), .S(n749) );
  FA_X1 U639 ( .A(n760), .B(n755), .CI(n753), .CO(n750), .S(n751) );
  FA_X1 U640 ( .A(n762), .B(n764), .CI(n757), .CO(n752), .S(n753) );
  FA_X1 U641 ( .A(n947), .B(n1001), .CI(n983), .CO(n754), .S(n755) );
  FA_X1 U642 ( .A(n965), .B(n929), .CI(n1020), .CO(n756), .S(n757) );
  FA_X1 U643 ( .A(n763), .B(n768), .CI(n761), .CO(n758), .S(n759) );
  FA_X1 U644 ( .A(n765), .B(n1021), .CI(n770), .CO(n760), .S(n761) );
  FA_X1 U645 ( .A(n966), .B(n984), .CI(n1002), .CO(n762), .S(n763) );
  HA_X1 U646 ( .A(n825), .B(n948), .CO(n764), .S(n765) );
  FA_X1 U647 ( .A(n771), .B(n774), .CI(n769), .CO(n766), .S(n767) );
  FA_X1 U648 ( .A(n967), .B(n1003), .CI(n776), .CO(n768), .S(n769) );
  FA_X1 U649 ( .A(n985), .B(n949), .CI(n1022), .CO(n770), .S(n771) );
  FA_X1 U650 ( .A(n780), .B(n777), .CI(n775), .CO(n772), .S(n773) );
  FA_X1 U651 ( .A(n986), .B(n1023), .CI(n1004), .CO(n774), .S(n775) );
  HA_X1 U652 ( .A(n826), .B(n968), .CO(n776), .S(n777) );
  FA_X1 U653 ( .A(n784), .B(n987), .CI(n781), .CO(n778), .S(n779) );
  FA_X1 U654 ( .A(n1024), .B(n969), .CI(n1005), .CO(n780), .S(n781) );
  FA_X1 U655 ( .A(n1006), .B(n1025), .CI(n785), .CO(n782), .S(n783) );
  HA_X1 U656 ( .A(n827), .B(n988), .CO(n784), .S(n785) );
  FA_X1 U657 ( .A(n1026), .B(n989), .CI(n1007), .CO(n786), .S(n787) );
  HA_X1 U658 ( .A(n1008), .B(n1027), .CO(n788), .S(n789) );
  CLKBUF_X3 U1180 ( .A(a[7]), .Z(n1383) );
  CLKBUF_X1 U1181 ( .A(a[7]), .Z(n19) );
  CLKBUF_X3 U1182 ( .A(n1277), .Z(n18) );
  AND2_X1 U1183 ( .A1(n521), .A2(n532), .ZN(n1384) );
  XNOR2_X1 U1184 ( .A(n298), .B(n1385), .ZN(product[22]) );
  AND2_X1 U1185 ( .A1(n1409), .A2(n297), .ZN(n1385) );
  CLKBUF_X3 U1186 ( .A(n291), .Z(n64) );
  CLKBUF_X1 U1187 ( .A(n64), .Z(n1386) );
  CLKBUF_X1 U1188 ( .A(n1123), .Z(n1443) );
  CLKBUF_X1 U1189 ( .A(n1284), .Z(n34) );
  CLKBUF_X2 U1190 ( .A(n1284), .Z(n33) );
  XNOR2_X1 U1191 ( .A(n1257), .B(n55), .ZN(n1387) );
  CLKBUF_X1 U1192 ( .A(n49), .Z(n1388) );
  CLKBUF_X3 U1193 ( .A(a[17]), .Z(n49) );
  CLKBUF_X3 U1194 ( .A(b[8]), .Z(n1251) );
  CLKBUF_X3 U1195 ( .A(b[13]), .Z(n1246) );
  CLKBUF_X1 U1196 ( .A(n1280), .Z(n58) );
  CLKBUF_X3 U1197 ( .A(b[10]), .Z(n1249) );
  CLKBUF_X3 U1198 ( .A(b[2]), .Z(n1257) );
  CLKBUF_X3 U1199 ( .A(b[4]), .Z(n1255) );
  AND2_X1 U1200 ( .A1(n509), .A2(n520), .ZN(n1389) );
  INV_X1 U1201 ( .A(n1389), .ZN(n256) );
  NAND2_X2 U1202 ( .A1(n282), .A2(n249), .ZN(n247) );
  CLKBUF_X1 U1203 ( .A(n1468), .Z(n1390) );
  CLKBUF_X1 U1204 ( .A(n283), .Z(n1391) );
  XOR2_X1 U1205 ( .A(n924), .B(n960), .Z(n1392) );
  XOR2_X1 U1206 ( .A(n906), .B(n1392), .Z(n703) );
  NAND2_X1 U1207 ( .A1(n906), .A2(n924), .ZN(n1393) );
  NAND2_X1 U1208 ( .A1(n906), .A2(n960), .ZN(n1394) );
  NAND2_X1 U1209 ( .A1(n924), .A2(n960), .ZN(n1395) );
  NAND3_X1 U1210 ( .A1(n1393), .A2(n1394), .A3(n1395), .ZN(n702) );
  CLKBUF_X3 U1211 ( .A(b[1]), .Z(n1258) );
  BUF_X1 U1212 ( .A(n1278), .Z(n12) );
  BUF_X1 U1213 ( .A(n1279), .Z(n6) );
  BUF_X1 U1214 ( .A(n61), .Z(n1489) );
  BUF_X2 U1215 ( .A(n1446), .Z(n1425) );
  BUF_X2 U1216 ( .A(b[14]), .Z(n1245) );
  CLKBUF_X3 U1217 ( .A(n43), .Z(n1487) );
  BUF_X2 U1218 ( .A(n61), .Z(n1442) );
  OAI22_X1 U1219 ( .A1(n60), .A2(n1031), .B1(n58), .B2(n1030), .ZN(n448) );
  BUF_X2 U1220 ( .A(n61), .Z(n1441) );
  NOR2_X1 U1221 ( .A1(n789), .A2(n828), .ZN(n402) );
  NOR2_X1 U1222 ( .A1(n481), .A2(n488), .ZN(n220) );
  BUF_X2 U1223 ( .A(n1274), .Z(n36) );
  CLKBUF_X3 U1224 ( .A(b[6]), .Z(n1253) );
  OR2_X1 U1225 ( .A1(n473), .A2(n480), .ZN(n1396) );
  OR2_X1 U1226 ( .A1(n759), .A2(n766), .ZN(n1397) );
  OR2_X1 U1227 ( .A1(n453), .A2(n456), .ZN(n1398) );
  OR2_X1 U1228 ( .A1(n467), .A2(n472), .ZN(n1399) );
  OR2_X1 U1229 ( .A1(n830), .A2(n448), .ZN(n1400) );
  OR2_X1 U1230 ( .A1(n452), .A2(n451), .ZN(n1401) );
  OR2_X1 U1231 ( .A1(n693), .A2(n706), .ZN(n1402) );
  OR2_X1 U1232 ( .A1(n450), .A2(n449), .ZN(n1403) );
  OR2_X1 U1233 ( .A1(n751), .A2(n758), .ZN(n1404) );
  OR2_X1 U1234 ( .A1(n457), .A2(n460), .ZN(n1405) );
  OR2_X1 U1235 ( .A1(n767), .A2(n772), .ZN(n1406) );
  OR2_X1 U1236 ( .A1(n779), .A2(n782), .ZN(n1407) );
  OR2_X1 U1237 ( .A1(n787), .A2(n788), .ZN(n1408) );
  OR2_X1 U1238 ( .A1(n1461), .A2(n592), .ZN(n1409) );
  OR2_X1 U1239 ( .A1(n1460), .A2(n628), .ZN(n1410) );
  NOR2_X1 U1240 ( .A1(n561), .A2(n576), .ZN(n289) );
  OR2_X1 U1241 ( .A1(n1029), .A2(n829), .ZN(n1411) );
  NOR2_X1 U1242 ( .A1(n489), .A2(n498), .ZN(n229) );
  NOR2_X1 U1243 ( .A1(n461), .A2(n466), .ZN(n179) );
  CLKBUF_X3 U1244 ( .A(b[9]), .Z(n1250) );
  CLKBUF_X3 U1245 ( .A(b[11]), .Z(n1248) );
  BUF_X2 U1246 ( .A(n1279), .Z(n1412) );
  INV_X1 U1247 ( .A(n1290), .ZN(n1413) );
  CLKBUF_X1 U1248 ( .A(n1250), .Z(n1414) );
  OAI22_X1 U1249 ( .A1(n42), .A2(n1094), .B1(n40), .B2(n1093), .ZN(n478) );
  XNOR2_X1 U1250 ( .A(n55), .B(n1258), .ZN(n1415) );
  CLKBUF_X1 U1251 ( .A(n1386), .Z(n1416) );
  NOR2_X1 U1252 ( .A1(n593), .A2(n610), .ZN(n1417) );
  BUF_X2 U1253 ( .A(n13), .Z(n1418) );
  BUF_X1 U1254 ( .A(n13), .Z(n1419) );
  BUF_X2 U1255 ( .A(n13), .Z(n1485) );
  BUF_X2 U1256 ( .A(a[5]), .Z(n13) );
  CLKBUF_X1 U1257 ( .A(n311), .Z(n1420) );
  CLKBUF_X1 U1258 ( .A(n1180), .Z(n1421) );
  CLKBUF_X1 U1259 ( .A(n1240), .Z(n1422) );
  XNOR2_X1 U1260 ( .A(n1487), .B(n1254), .ZN(n1423) );
  CLKBUF_X1 U1261 ( .A(n1446), .Z(n1424) );
  BUF_X1 U1262 ( .A(a[9]), .Z(n1446) );
  OR2_X1 U1263 ( .A1(n312), .A2(n317), .ZN(n1426) );
  XNOR2_X1 U1264 ( .A(n55), .B(n1256), .ZN(n1427) );
  BUF_X2 U1265 ( .A(n1270), .Z(n59) );
  BUF_X1 U1266 ( .A(n1271), .Z(n1428) );
  CLKBUF_X1 U1267 ( .A(n1240), .Z(n1429) );
  NOR2_X1 U1268 ( .A1(n593), .A2(n610), .ZN(n303) );
  NAND2_X1 U1269 ( .A1(n1266), .A2(n1286), .ZN(n1276) );
  BUF_X1 U1270 ( .A(n1464), .Z(n1452) );
  CLKBUF_X1 U1271 ( .A(n1184), .Z(n1430) );
  CLKBUF_X1 U1272 ( .A(n304), .Z(n1431) );
  OAI22_X1 U1273 ( .A1(n24), .A2(n1157), .B1(n22), .B2(n1156), .ZN(n544) );
  BUF_X1 U1274 ( .A(n1286), .Z(n22) );
  BUF_X2 U1275 ( .A(b[19]), .Z(n1240) );
  OR2_X1 U1276 ( .A1(n663), .A2(n678), .ZN(n1468) );
  OR2_X2 U1277 ( .A1(n509), .A2(n520), .ZN(n1432) );
  BUF_X1 U1278 ( .A(n320), .Z(n1476) );
  CLKBUF_X3 U1279 ( .A(b[18]), .Z(n1241) );
  XNOR2_X1 U1280 ( .A(n198), .B(n1433), .ZN(product[32]) );
  AND2_X1 U1281 ( .A1(n1399), .A2(n197), .ZN(n1433) );
  XOR2_X1 U1282 ( .A(n630), .B(n615), .Z(n1434) );
  XOR2_X1 U1283 ( .A(n613), .B(n1434), .Z(n611) );
  NAND2_X1 U1284 ( .A1(n613), .A2(n630), .ZN(n1435) );
  NAND2_X1 U1285 ( .A1(n613), .A2(n615), .ZN(n1436) );
  NAND2_X1 U1286 ( .A1(n630), .A2(n615), .ZN(n1437) );
  NAND3_X1 U1287 ( .A1(n1435), .A2(n1436), .A3(n1437), .ZN(n610) );
  BUF_X2 U1288 ( .A(n1280), .Z(n57) );
  CLKBUF_X1 U1289 ( .A(n1), .Z(n1438) );
  CLKBUF_X1 U1290 ( .A(n1278), .Z(n1439) );
  CLKBUF_X1 U1291 ( .A(n1278), .Z(n1440) );
  BUF_X1 U1292 ( .A(n1124), .Z(n1444) );
  BUF_X4 U1293 ( .A(a[19]), .Z(n55) );
  CLKBUF_X1 U1294 ( .A(n49), .Z(n1445) );
  CLKBUF_X1 U1295 ( .A(a[9]), .Z(n25) );
  XNOR2_X1 U1296 ( .A(n286), .B(n1447), .ZN(product[24]) );
  AND2_X1 U1297 ( .A1(n424), .A2(n285), .ZN(n1447) );
  CLKBUF_X3 U1298 ( .A(a[13]), .Z(n1448) );
  CLKBUF_X1 U1299 ( .A(a[13]), .Z(n37) );
  CLKBUF_X1 U1300 ( .A(n1257), .Z(n1449) );
  XNOR2_X1 U1301 ( .A(n1419), .B(n1242), .ZN(n1450) );
  BUF_X2 U1302 ( .A(n13), .Z(n1484) );
  XNOR2_X1 U1303 ( .A(n1240), .B(n1), .ZN(n1451) );
  BUF_X1 U1304 ( .A(n1464), .Z(n1453) );
  CLKBUF_X1 U1305 ( .A(n1464), .Z(n1454) );
  BUF_X1 U1306 ( .A(n248), .Z(n1464) );
  XNOR2_X1 U1307 ( .A(n244), .B(n1455), .ZN(product[28]) );
  AND2_X1 U1308 ( .A1(n240), .A2(n243), .ZN(n1455) );
  XNOR2_X1 U1309 ( .A(n257), .B(n1456), .ZN(product[27]) );
  AND2_X1 U1310 ( .A1(n1432), .A2(n256), .ZN(n1456) );
  XNOR2_X1 U1311 ( .A(n209), .B(n1457), .ZN(product[31]) );
  AND2_X1 U1312 ( .A1(n1396), .A2(n208), .ZN(n1457) );
  BUF_X1 U1313 ( .A(n248), .Z(n65) );
  XNOR2_X1 U1314 ( .A(n277), .B(n1458), .ZN(product[25]) );
  AND2_X1 U1315 ( .A1(n273), .A2(n276), .ZN(n1458) );
  NOR2_X2 U1316 ( .A1(n647), .A2(n662), .ZN(n323) );
  XNOR2_X1 U1317 ( .A(n231), .B(n1459), .ZN(product[29]) );
  AND2_X1 U1318 ( .A1(n227), .A2(n230), .ZN(n1459) );
  CLKBUF_X1 U1319 ( .A(n611), .Z(n1460) );
  CLKBUF_X1 U1320 ( .A(n577), .Z(n1461) );
  NOR2_X2 U1321 ( .A1(n707), .A2(n718), .ZN(n350) );
  CLKBUF_X1 U1322 ( .A(n31), .Z(n1462) );
  OAI21_X1 U1323 ( .B1(n368), .B2(n380), .A(n369), .ZN(n367) );
  NOR2_X1 U1324 ( .A1(n611), .A2(n628), .ZN(n1463) );
  NOR2_X1 U1325 ( .A1(n611), .A2(n628), .ZN(n312) );
  BUF_X2 U1326 ( .A(n1271), .Z(n53) );
  BUF_X1 U1327 ( .A(n1282), .Z(n46) );
  BUF_X1 U1328 ( .A(b[0]), .Z(n61) );
  NOR2_X1 U1329 ( .A1(n1417), .A2(n296), .ZN(n1465) );
  CLKBUF_X1 U1330 ( .A(n1453), .Z(n1466) );
  CLKBUF_X1 U1331 ( .A(n318), .Z(n1467) );
  NAND2_X1 U1332 ( .A1(n1265), .A2(n1285), .ZN(n1275) );
  BUF_X2 U1333 ( .A(n1285), .Z(n27) );
  BUF_X2 U1334 ( .A(n1285), .Z(n28) );
  CLKBUF_X3 U1335 ( .A(b[17]), .Z(n1242) );
  NOR2_X1 U1336 ( .A1(n533), .A2(n546), .ZN(n275) );
  CLKBUF_X3 U1337 ( .A(b[7]), .Z(n1252) );
  NOR2_X2 U1338 ( .A1(n547), .A2(n560), .ZN(n284) );
  NOR2_X1 U1339 ( .A1(n577), .A2(n592), .ZN(n1469) );
  CLKBUF_X1 U1340 ( .A(n1249), .Z(n1470) );
  NOR2_X1 U1341 ( .A1(n577), .A2(n592), .ZN(n296) );
  OR2_X1 U1342 ( .A1(n521), .A2(n532), .ZN(n1471) );
  BUF_X2 U1343 ( .A(n1274), .Z(n35) );
  BUF_X2 U1344 ( .A(n1282), .Z(n45) );
  BUF_X2 U1345 ( .A(n1272), .Z(n47) );
  BUF_X2 U1346 ( .A(n43), .Z(n1486) );
  CLKBUF_X3 U1347 ( .A(b[12]), .Z(n1247) );
  NAND2_X1 U1348 ( .A1(n1260), .A2(n1280), .ZN(n1270) );
  CLKBUF_X3 U1349 ( .A(b[5]), .Z(n1254) );
  XOR2_X1 U1350 ( .A(n701), .B(n714), .Z(n1472) );
  XOR2_X1 U1351 ( .A(n712), .B(n1472), .Z(n697) );
  NAND2_X1 U1352 ( .A1(n712), .A2(n701), .ZN(n1473) );
  NAND2_X1 U1353 ( .A1(n712), .A2(n714), .ZN(n1474) );
  NAND2_X1 U1354 ( .A1(n701), .A2(n714), .ZN(n1475) );
  NAND3_X1 U1355 ( .A1(n1473), .A2(n1474), .A3(n1475), .ZN(n696) );
  AOI21_X1 U1356 ( .B1(n1390), .B2(n336), .A(n329), .ZN(n1477) );
  CLKBUF_X3 U1357 ( .A(b[15]), .Z(n1244) );
  CLKBUF_X3 U1358 ( .A(b[16]), .Z(n1243) );
  OAI21_X1 U1359 ( .B1(n292), .B2(n320), .A(n293), .ZN(n291) );
  AOI21_X1 U1360 ( .B1(n340), .B2(n321), .A(n322), .ZN(n320) );
  BUF_X2 U1361 ( .A(n1276), .Z(n23) );
  BUF_X2 U1362 ( .A(n1286), .Z(n21) );
  NAND2_X1 U1363 ( .A1(n1267), .A2(n1287), .ZN(n1277) );
  BUF_X1 U1364 ( .A(n1287), .Z(n16) );
  BUF_X1 U1365 ( .A(n1287), .Z(n15) );
  XNOR2_X1 U1366 ( .A(a[4]), .B(a[3]), .ZN(n1287) );
  BUF_X2 U1367 ( .A(n1283), .Z(n40) );
  NAND2_X1 U1368 ( .A1(n1263), .A2(n1283), .ZN(n1273) );
  BUF_X2 U1369 ( .A(n1283), .Z(n39) );
  XNOR2_X1 U1370 ( .A(n268), .B(n1478), .ZN(product[26]) );
  AND2_X1 U1371 ( .A1(n262), .A2(n267), .ZN(n1478) );
  NOR2_X1 U1372 ( .A1(n251), .A2(n275), .ZN(n249) );
  AOI21_X1 U1373 ( .B1(n218), .B2(n241), .A(n219), .ZN(n217) );
  XNOR2_X1 U1374 ( .A(n222), .B(n1479), .ZN(product[30]) );
  AND2_X1 U1375 ( .A1(n418), .A2(n221), .ZN(n1479) );
  XNOR2_X1 U1376 ( .A(n181), .B(n1480), .ZN(product[33]) );
  AND2_X1 U1377 ( .A1(n177), .A2(n180), .ZN(n1480) );
  NOR2_X1 U1378 ( .A1(n629), .A2(n646), .ZN(n317) );
  NOR2_X1 U1379 ( .A1(n229), .A2(n220), .ZN(n218) );
  NAND2_X1 U1380 ( .A1(n533), .A2(n546), .ZN(n276) );
  XNOR2_X1 U1381 ( .A(n157), .B(n1481), .ZN(product[35]) );
  AND2_X1 U1382 ( .A1(n1398), .A2(n156), .ZN(n1481) );
  XNOR2_X1 U1383 ( .A(n168), .B(n1482), .ZN(product[34]) );
  AND2_X1 U1384 ( .A1(n1405), .A2(n167), .ZN(n1482) );
  NOR2_X1 U1385 ( .A1(n741), .A2(n750), .ZN(n364) );
  NOR2_X1 U1386 ( .A1(n499), .A2(n508), .ZN(n242) );
  NAND2_X1 U1387 ( .A1(n489), .A2(n498), .ZN(n230) );
  NAND2_X1 U1388 ( .A1(n461), .A2(n466), .ZN(n180) );
  NOR2_X1 U1389 ( .A1(n773), .A2(n778), .ZN(n386) );
  AND2_X1 U1390 ( .A1(n1411), .A2(n409), .ZN(product[1]) );
  BUF_X2 U1391 ( .A(n1281), .Z(n51) );
  BUF_X2 U1392 ( .A(n1270), .Z(n60) );
  BUF_X2 U1393 ( .A(n1273), .Z(n41) );
  BUF_X2 U1394 ( .A(n1277), .Z(n17) );
  NAND2_X1 U1395 ( .A1(n1261), .A2(n1281), .ZN(n1271) );
  NAND2_X1 U1396 ( .A1(n1262), .A2(n1282), .ZN(n1272) );
  INV_X1 U1397 ( .A(a[0]), .ZN(n1289) );
  NAND2_X1 U1398 ( .A1(n1284), .A2(n1264), .ZN(n1274) );
  NAND2_X1 U1399 ( .A1(n1269), .A2(n1289), .ZN(n1279) );
  NOR2_X1 U1400 ( .A1(n280), .A2(n260), .ZN(n258) );
  NOR2_X1 U1401 ( .A1(n280), .A2(n271), .ZN(n269) );
  NOR2_X1 U1402 ( .A1(n247), .A2(n184), .ZN(n182) );
  NOR2_X1 U1403 ( .A1(n247), .A2(n171), .ZN(n169) );
  NOR2_X1 U1404 ( .A1(n247), .A2(n216), .ZN(n210) );
  NOR2_X1 U1405 ( .A1(n247), .A2(n145), .ZN(n143) );
  NOR2_X1 U1406 ( .A1(n247), .A2(n130), .ZN(n128) );
  NOR2_X1 U1407 ( .A1(n247), .A2(n201), .ZN(n199) );
  NOR2_X1 U1408 ( .A1(n247), .A2(n117), .ZN(n115) );
  NOR2_X1 U1409 ( .A1(n247), .A2(n242), .ZN(n232) );
  NAND2_X1 U1410 ( .A1(n214), .A2(n134), .ZN(n130) );
  INV_X1 U1411 ( .A(n186), .ZN(n184) );
  INV_X1 U1412 ( .A(n173), .ZN(n171) );
  INV_X1 U1413 ( .A(n1426), .ZN(n306) );
  INV_X1 U1414 ( .A(n280), .ZN(n278) );
  INV_X1 U1415 ( .A(n247), .ZN(n245) );
  INV_X1 U1416 ( .A(n1476), .ZN(n319) );
  NOR2_X1 U1417 ( .A1(n216), .A2(n192), .ZN(n186) );
  NOR2_X1 U1418 ( .A1(n216), .A2(n175), .ZN(n173) );
  INV_X1 U1419 ( .A(n187), .ZN(n185) );
  INV_X1 U1420 ( .A(n282), .ZN(n280) );
  INV_X1 U1421 ( .A(n340), .ZN(n339) );
  NOR2_X1 U1422 ( .A1(n1426), .A2(n301), .ZN(n299) );
  INV_X1 U1423 ( .A(n1391), .ZN(n281) );
  INV_X1 U1424 ( .A(n216), .ZN(n214) );
  BUF_X2 U1425 ( .A(n291), .Z(n63) );
  NAND2_X1 U1426 ( .A1(n1471), .A2(n1432), .ZN(n251) );
  NAND2_X1 U1427 ( .A1(n273), .A2(n262), .ZN(n260) );
  OAI21_X1 U1428 ( .B1(n281), .B2(n260), .A(n261), .ZN(n259) );
  AOI21_X1 U1429 ( .B1(n274), .B2(n262), .A(n1384), .ZN(n261) );
  OAI21_X1 U1430 ( .B1(n281), .B2(n271), .A(n276), .ZN(n270) );
  INV_X1 U1431 ( .A(n1420), .ZN(n309) );
  INV_X1 U1432 ( .A(n273), .ZN(n271) );
  NOR2_X1 U1433 ( .A1(n247), .A2(n225), .ZN(n223) );
  NOR2_X1 U1434 ( .A1(n247), .A2(n160), .ZN(n158) );
  NAND2_X1 U1435 ( .A1(n186), .A2(n149), .ZN(n145) );
  NAND2_X1 U1436 ( .A1(n214), .A2(n1396), .ZN(n201) );
  INV_X1 U1437 ( .A(n192), .ZN(n190) );
  INV_X1 U1438 ( .A(n119), .ZN(n117) );
  NAND2_X1 U1439 ( .A1(n1468), .A2(n335), .ZN(n326) );
  INV_X1 U1440 ( .A(n263), .ZN(n262) );
  INV_X1 U1441 ( .A(n1471), .ZN(n263) );
  INV_X1 U1442 ( .A(n336), .ZN(n334) );
  INV_X1 U1443 ( .A(n1452), .ZN(n246) );
  NAND2_X1 U1444 ( .A1(n287), .A2(n290), .ZN(n82) );
  XOR2_X1 U1445 ( .A(n352), .B(n91), .Z(product[14]) );
  NAND2_X1 U1446 ( .A1(n434), .A2(n351), .ZN(n91) );
  AOI21_X1 U1447 ( .B1(n357), .B2(n435), .A(n354), .ZN(n352) );
  INV_X1 U1448 ( .A(n350), .ZN(n434) );
  XOR2_X1 U1449 ( .A(n339), .B(n89), .Z(product[16]) );
  NAND2_X1 U1450 ( .A1(n335), .A2(n338), .ZN(n89) );
  XOR2_X1 U1451 ( .A(n347), .B(n90), .Z(product[15]) );
  NAND2_X1 U1452 ( .A1(n1402), .A2(n346), .ZN(n90) );
  XNOR2_X1 U1453 ( .A(n325), .B(n87), .ZN(product[18]) );
  NAND2_X1 U1454 ( .A1(n430), .A2(n324), .ZN(n87) );
  INV_X1 U1455 ( .A(n323), .ZN(n430) );
  XNOR2_X1 U1456 ( .A(n332), .B(n88), .ZN(product[17]) );
  NAND2_X1 U1457 ( .A1(n1390), .A2(n331), .ZN(n88) );
  OAI21_X1 U1458 ( .B1(n339), .B2(n337), .A(n334), .ZN(n332) );
  NOR2_X1 U1459 ( .A1(n303), .A2(n296), .ZN(n294) );
  AOI21_X1 U1460 ( .B1(n299), .B2(n319), .A(n300), .ZN(n298) );
  OAI21_X1 U1461 ( .B1(n327), .B2(n323), .A(n324), .ZN(n322) );
  AOI21_X1 U1462 ( .B1(n1465), .B2(n311), .A(n295), .ZN(n293) );
  NAND2_X1 U1463 ( .A1(n294), .A2(n310), .ZN(n292) );
  OAI21_X1 U1464 ( .B1(n341), .B2(n358), .A(n342), .ZN(n340) );
  NAND2_X1 U1465 ( .A1(n348), .A2(n1402), .ZN(n341) );
  INV_X1 U1466 ( .A(n284), .ZN(n424) );
  XOR2_X1 U1467 ( .A(n314), .B(n85), .Z(product[20]) );
  NAND2_X1 U1468 ( .A1(n1410), .A2(n313), .ZN(n85) );
  AOI21_X1 U1469 ( .B1(n319), .B2(n315), .A(n316), .ZN(n314) );
  XOR2_X1 U1470 ( .A(n305), .B(n84), .Z(product[21]) );
  NAND2_X1 U1471 ( .A1(n427), .A2(n1431), .ZN(n84) );
  AOI21_X1 U1472 ( .B1(n319), .B2(n306), .A(n1420), .ZN(n305) );
  INV_X1 U1473 ( .A(n303), .ZN(n427) );
  OAI21_X1 U1474 ( .B1(n1463), .B2(n318), .A(n313), .ZN(n311) );
  OAI21_X1 U1475 ( .B1(n217), .B2(n192), .A(n193), .ZN(n187) );
  OAI21_X1 U1476 ( .B1(n284), .B2(n290), .A(n285), .ZN(n283) );
  AOI21_X1 U1477 ( .B1(n1468), .B2(n336), .A(n329), .ZN(n327) );
  INV_X1 U1478 ( .A(n331), .ZN(n329) );
  NOR2_X1 U1479 ( .A1(n216), .A2(n121), .ZN(n119) );
  NOR2_X1 U1480 ( .A1(n312), .A2(n317), .ZN(n310) );
  NAND2_X1 U1481 ( .A1(n218), .A2(n240), .ZN(n216) );
  AOI21_X1 U1482 ( .B1(n283), .B2(n249), .A(n250), .ZN(n248) );
  OAI21_X1 U1483 ( .B1(n251), .B2(n276), .A(n252), .ZN(n250) );
  AOI21_X1 U1484 ( .B1(n1432), .B2(n1384), .A(n1389), .ZN(n252) );
  XNOR2_X1 U1485 ( .A(n319), .B(n86), .ZN(product[19]) );
  NAND2_X1 U1486 ( .A1(n315), .A2(n1467), .ZN(n86) );
  AOI21_X1 U1487 ( .B1(n215), .B2(n1396), .A(n206), .ZN(n202) );
  INV_X1 U1488 ( .A(n174), .ZN(n172) );
  OAI21_X1 U1489 ( .B1(n309), .B2(n301), .A(n1431), .ZN(n300) );
  INV_X1 U1490 ( .A(n337), .ZN(n335) );
  INV_X1 U1491 ( .A(n217), .ZN(n215) );
  NOR2_X1 U1492 ( .A1(n192), .A2(n136), .ZN(n134) );
  INV_X1 U1493 ( .A(n275), .ZN(n273) );
  NAND2_X1 U1494 ( .A1(n190), .A2(n177), .ZN(n175) );
  NAND2_X1 U1495 ( .A1(n1396), .A2(n1399), .ZN(n192) );
  INV_X1 U1496 ( .A(n317), .ZN(n315) );
  INV_X1 U1497 ( .A(n276), .ZN(n274) );
  INV_X1 U1498 ( .A(n338), .ZN(n336) );
  NAND2_X1 U1499 ( .A1(n240), .A2(n227), .ZN(n225) );
  INV_X1 U1500 ( .A(n427), .ZN(n301) );
  INV_X1 U1501 ( .A(n193), .ZN(n191) );
  INV_X1 U1502 ( .A(n367), .ZN(n366) );
  NAND2_X1 U1503 ( .A1(n173), .A2(n1405), .ZN(n160) );
  INV_X1 U1504 ( .A(n1467), .ZN(n316) );
  INV_X1 U1505 ( .A(n290), .ZN(n288) );
  INV_X1 U1506 ( .A(n289), .ZN(n287) );
  INV_X1 U1507 ( .A(n346), .ZN(n344) );
  XOR2_X1 U1508 ( .A(n374), .B(n95), .Z(product[10]) );
  NAND2_X1 U1509 ( .A1(n1404), .A2(n373), .ZN(n95) );
  AOI21_X1 U1510 ( .B1(n379), .B2(n1397), .A(n376), .ZN(n374) );
  OAI21_X1 U1511 ( .B1(n230), .B2(n220), .A(n221), .ZN(n219) );
  XNOR2_X1 U1512 ( .A(n357), .B(n92), .ZN(product[13]) );
  NAND2_X1 U1513 ( .A1(n435), .A2(n356), .ZN(n92) );
  INV_X1 U1514 ( .A(n355), .ZN(n435) );
  XNOR2_X1 U1515 ( .A(n363), .B(n93), .ZN(product[12]) );
  NAND2_X1 U1516 ( .A1(n436), .A2(n362), .ZN(n93) );
  OAI21_X1 U1517 ( .B1(n366), .B2(n364), .A(n365), .ZN(n363) );
  XNOR2_X1 U1518 ( .A(n379), .B(n96), .ZN(product[9]) );
  NAND2_X1 U1519 ( .A1(n1397), .A2(n378), .ZN(n96) );
  NAND2_X1 U1520 ( .A1(n1404), .A2(n1397), .ZN(n368) );
  AOI21_X1 U1521 ( .B1(n1404), .B2(n376), .A(n371), .ZN(n369) );
  AOI21_X1 U1522 ( .B1(n1399), .B2(n206), .A(n195), .ZN(n193) );
  INV_X1 U1523 ( .A(n197), .ZN(n195) );
  INV_X1 U1524 ( .A(n220), .ZN(n418) );
  NOR2_X1 U1525 ( .A1(n350), .A2(n355), .ZN(n348) );
  AOI21_X1 U1526 ( .B1(n367), .B2(n359), .A(n360), .ZN(n358) );
  OAI21_X1 U1527 ( .B1(n217), .B2(n175), .A(n176), .ZN(n174) );
  AOI21_X1 U1528 ( .B1(n191), .B2(n177), .A(n178), .ZN(n176) );
  INV_X1 U1529 ( .A(n180), .ZN(n178) );
  NAND2_X1 U1530 ( .A1(n663), .A2(n678), .ZN(n331) );
  NAND2_X1 U1531 ( .A1(n149), .A2(n1401), .ZN(n136) );
  NAND2_X1 U1532 ( .A1(n693), .A2(n706), .ZN(n346) );
  NOR2_X1 U1533 ( .A1(n692), .A2(n679), .ZN(n337) );
  AOI21_X1 U1534 ( .B1(n174), .B2(n1405), .A(n165), .ZN(n161) );
  AOI21_X1 U1535 ( .B1(n187), .B2(n149), .A(n150), .ZN(n146) );
  AOI21_X1 U1536 ( .B1(n215), .B2(n134), .A(n135), .ZN(n131) );
  AOI21_X1 U1537 ( .B1(n241), .B2(n227), .A(n228), .ZN(n226) );
  INV_X1 U1538 ( .A(n230), .ZN(n228) );
  INV_X1 U1539 ( .A(n120), .ZN(n118) );
  NAND2_X1 U1540 ( .A1(n561), .A2(n576), .ZN(n290) );
  NAND2_X1 U1541 ( .A1(n629), .A2(n646), .ZN(n318) );
  NAND2_X1 U1542 ( .A1(n593), .A2(n610), .ZN(n304) );
  NOR2_X1 U1543 ( .A1(n179), .A2(n151), .ZN(n149) );
  INV_X1 U1544 ( .A(n380), .ZN(n379) );
  NAND2_X1 U1545 ( .A1(n679), .A2(n692), .ZN(n338) );
  NAND2_X1 U1546 ( .A1(n647), .A2(n662), .ZN(n324) );
  NAND2_X1 U1547 ( .A1(n547), .A2(n560), .ZN(n285) );
  NAND2_X1 U1548 ( .A1(n611), .A2(n628), .ZN(n313) );
  NAND2_X1 U1549 ( .A1(n521), .A2(n532), .ZN(n267) );
  INV_X1 U1550 ( .A(n229), .ZN(n227) );
  INV_X1 U1551 ( .A(n179), .ZN(n177) );
  NAND2_X1 U1552 ( .A1(n1405), .A2(n1398), .ZN(n151) );
  NAND2_X1 U1553 ( .A1(n707), .A2(n718), .ZN(n351) );
  INV_X1 U1554 ( .A(n378), .ZN(n376) );
  INV_X1 U1555 ( .A(n242), .ZN(n240) );
  NAND2_X1 U1556 ( .A1(n577), .A2(n592), .ZN(n297) );
  INV_X1 U1557 ( .A(n243), .ZN(n241) );
  INV_X1 U1558 ( .A(n208), .ZN(n206) );
  NOR2_X1 U1559 ( .A1(n247), .A2(n108), .ZN(n106) );
  NAND2_X1 U1560 ( .A1(n119), .A2(n1400), .ZN(n108) );
  XOR2_X1 U1561 ( .A(n366), .B(n94), .Z(product[11]) );
  NAND2_X1 U1562 ( .A1(n437), .A2(n365), .ZN(n94) );
  INV_X1 U1563 ( .A(n364), .ZN(n437) );
  INV_X1 U1564 ( .A(n356), .ZN(n354) );
  INV_X1 U1565 ( .A(n373), .ZN(n371) );
  XOR2_X1 U1566 ( .A(n114), .B(n67), .Z(product[38]) );
  NAND2_X1 U1567 ( .A1(n1400), .A2(n113), .ZN(n67) );
  NAND2_X1 U1568 ( .A1(n1403), .A2(n126), .ZN(n68) );
  NAND2_X1 U1569 ( .A1(n1401), .A2(n141), .ZN(n69) );
  OAI21_X1 U1570 ( .B1(n388), .B2(n386), .A(n387), .ZN(n385) );
  AOI21_X1 U1571 ( .B1(n1407), .B2(n393), .A(n390), .ZN(n388) );
  INV_X1 U1572 ( .A(n392), .ZN(n390) );
  OAI21_X1 U1573 ( .B1(n394), .B2(n396), .A(n395), .ZN(n393) );
  OAI21_X1 U1574 ( .B1(n151), .B2(n180), .A(n152), .ZN(n150) );
  AOI21_X1 U1575 ( .B1(n165), .B2(n1398), .A(n154), .ZN(n152) );
  INV_X1 U1576 ( .A(n156), .ZN(n154) );
  NOR2_X1 U1577 ( .A1(n719), .A2(n730), .ZN(n355) );
  OAI21_X1 U1578 ( .B1(n193), .B2(n136), .A(n137), .ZN(n135) );
  AOI21_X1 U1579 ( .B1(n150), .B2(n1401), .A(n139), .ZN(n137) );
  INV_X1 U1580 ( .A(n141), .ZN(n139) );
  OAI21_X1 U1581 ( .B1(n217), .B2(n121), .A(n122), .ZN(n120) );
  AOI21_X1 U1582 ( .B1(n135), .B2(n1403), .A(n124), .ZN(n122) );
  INV_X1 U1583 ( .A(n126), .ZN(n124) );
  XNOR2_X1 U1584 ( .A(n385), .B(n97), .ZN(product[8]) );
  NAND2_X1 U1585 ( .A1(n1406), .A2(n384), .ZN(n97) );
  NAND2_X1 U1586 ( .A1(n719), .A2(n730), .ZN(n356) );
  NAND2_X1 U1587 ( .A1(n741), .A2(n750), .ZN(n365) );
  AOI21_X1 U1588 ( .B1(n120), .B2(n1400), .A(n111), .ZN(n109) );
  INV_X1 U1589 ( .A(n113), .ZN(n111) );
  NAND2_X1 U1590 ( .A1(n473), .A2(n480), .ZN(n208) );
  NAND2_X1 U1591 ( .A1(n499), .A2(n508), .ZN(n243) );
  NAND2_X1 U1592 ( .A1(n467), .A2(n472), .ZN(n197) );
  NAND2_X1 U1593 ( .A1(n481), .A2(n488), .ZN(n221) );
  NAND2_X1 U1594 ( .A1(n751), .A2(n758), .ZN(n373) );
  NAND2_X1 U1595 ( .A1(n731), .A2(n740), .ZN(n362) );
  INV_X1 U1596 ( .A(n167), .ZN(n165) );
  NAND2_X1 U1597 ( .A1(n441), .A2(n387), .ZN(n98) );
  INV_X1 U1598 ( .A(n386), .ZN(n441) );
  NAND2_X1 U1599 ( .A1(n1407), .A2(n392), .ZN(n99) );
  AOI21_X1 U1600 ( .B1(n385), .B2(n1406), .A(n382), .ZN(n380) );
  INV_X1 U1601 ( .A(n384), .ZN(n382) );
  XOR2_X1 U1602 ( .A(n100), .B(n396), .Z(product[5]) );
  NAND2_X1 U1603 ( .A1(n443), .A2(n395), .ZN(n100) );
  INV_X1 U1604 ( .A(n394), .ZN(n443) );
  NOR2_X1 U1605 ( .A1(n1028), .A2(n1009), .ZN(n406) );
  XOR2_X1 U1606 ( .A(n102), .B(n404), .Z(product[3]) );
  NAND2_X1 U1607 ( .A1(n445), .A2(n403), .ZN(n102) );
  INV_X1 U1608 ( .A(n402), .ZN(n445) );
  OAI21_X1 U1609 ( .B1(n402), .B2(n404), .A(n403), .ZN(n401) );
  AOI21_X1 U1610 ( .B1(n1408), .B2(n401), .A(n398), .ZN(n396) );
  INV_X1 U1611 ( .A(n400), .ZN(n398) );
  NAND2_X1 U1612 ( .A1(n830), .A2(n448), .ZN(n113) );
  NOR2_X1 U1613 ( .A1(n783), .A2(n786), .ZN(n394) );
  INV_X1 U1614 ( .A(n448), .ZN(n449) );
  INV_X1 U1615 ( .A(n544), .ZN(n545) );
  INV_X1 U1616 ( .A(n478), .ZN(n479) );
  OR2_X1 U1617 ( .A1(n937), .A2(n865), .ZN(n626) );
  XNOR2_X1 U1618 ( .A(n937), .B(n865), .ZN(n627) );
  NAND2_X1 U1619 ( .A1(n453), .A2(n456), .ZN(n156) );
  NAND2_X1 U1620 ( .A1(n457), .A2(n460), .ZN(n167) );
  NAND2_X1 U1621 ( .A1(n779), .A2(n782), .ZN(n392) );
  NAND2_X1 U1622 ( .A1(n452), .A2(n451), .ZN(n141) );
  NAND2_X1 U1623 ( .A1(n450), .A2(n449), .ZN(n126) );
  NAND2_X1 U1624 ( .A1(n767), .A2(n772), .ZN(n384) );
  NAND2_X1 U1625 ( .A1(n783), .A2(n786), .ZN(n395) );
  NAND2_X1 U1626 ( .A1(n773), .A2(n778), .ZN(n387) );
  XOR2_X1 U1627 ( .A(n103), .B(n409), .Z(product[2]) );
  NAND2_X1 U1628 ( .A1(n446), .A2(n407), .ZN(n103) );
  INV_X1 U1629 ( .A(n406), .ZN(n446) );
  INV_X1 U1630 ( .A(n405), .ZN(n404) );
  OAI21_X1 U1631 ( .B1(n406), .B2(n409), .A(n407), .ZN(n405) );
  XNOR2_X1 U1632 ( .A(n101), .B(n401), .ZN(product[4]) );
  NAND2_X1 U1633 ( .A1(n1408), .A2(n400), .ZN(n101) );
  OAI22_X1 U1634 ( .A1(n30), .A2(n1136), .B1(n28), .B2(n1135), .ZN(n518) );
  OAI22_X1 U1635 ( .A1(n30), .A2(n1143), .B1(n28), .B2(n1142), .ZN(n937) );
  OAI22_X1 U1636 ( .A1(n18), .A2(n1178), .B1(n16), .B2(n1177), .ZN(n574) );
  OAI22_X1 U1637 ( .A1(n11), .A2(n1199), .B1(n10), .B2(n1198), .ZN(n608) );
  OAI22_X1 U1638 ( .A1(n48), .A2(n1073), .B1(n46), .B2(n1072), .ZN(n464) );
  OAI22_X1 U1639 ( .A1(n36), .A2(n1115), .B1(n34), .B2(n1114), .ZN(n496) );
  OAI22_X1 U1640 ( .A1(n1428), .A2(n1067), .B1(n51), .B2(n1066), .ZN(n865) );
  OAI22_X1 U1641 ( .A1(n54), .A2(n1065), .B1(n51), .B2(n1064), .ZN(n863) );
  OAI22_X1 U1642 ( .A1(n24), .A2(n1160), .B1(n22), .B2(n1159), .ZN(n953) );
  OAI22_X1 U1643 ( .A1(n53), .A2(n1068), .B1(n1067), .B2(n51), .ZN(n866) );
  OAI22_X1 U1644 ( .A1(n47), .A2(n1087), .B1(n45), .B2(n1086), .ZN(n884) );
  OAI22_X1 U1645 ( .A1(n30), .A2(n1144), .B1(n28), .B2(n1143), .ZN(n938) );
  OAI22_X1 U1646 ( .A1(n54), .A2(n1063), .B1(n51), .B2(n1062), .ZN(n861) );
  OAI22_X1 U1647 ( .A1(n24), .A2(n1158), .B1(n22), .B2(n1157), .ZN(n951) );
  OAI22_X1 U1648 ( .A1(n30), .A2(n1139), .B1(n28), .B2(n1138), .ZN(n933) );
  OAI22_X1 U1649 ( .A1(n60), .A2(n1034), .B1(n58), .B2(n1033), .ZN(n833) );
  OAI22_X1 U1650 ( .A1(n60), .A2(n1033), .B1(n58), .B2(n1032), .ZN(n832) );
  INV_X1 U1651 ( .A(n454), .ZN(n455) );
  OAI22_X1 U1652 ( .A1(n17), .A2(n1195), .B1(n15), .B2(n1194), .ZN(n987) );
  OAI22_X1 U1653 ( .A1(n1440), .A2(n1215), .B1(n9), .B2(n1214), .ZN(n1006) );
  OAI22_X1 U1654 ( .A1(n1412), .A2(n1234), .B1(n1233), .B2(n3), .ZN(n1025) );
  AND2_X1 U1655 ( .A1(n1490), .A2(n812), .ZN(n989) );
  OAI22_X1 U1656 ( .A1(n1440), .A2(n1216), .B1(n9), .B2(n1215), .ZN(n1007) );
  OAI22_X1 U1657 ( .A1(n5), .A2(n1235), .B1(n1234), .B2(n3), .ZN(n1026) );
  OAI22_X1 U1658 ( .A1(n47), .A2(n1091), .B1(n45), .B2(n1090), .ZN(n888) );
  OAI22_X1 U1659 ( .A1(n48), .A2(n1292), .B1(n1092), .B2(n46), .ZN(n822) );
  XNOR2_X1 U1660 ( .A(n1487), .B(n1490), .ZN(n1091) );
  OAI22_X1 U1661 ( .A1(n11), .A2(n1213), .B1(n9), .B2(n1212), .ZN(n1004) );
  OAI22_X1 U1662 ( .A1(n5), .A2(n1232), .B1(n1231), .B2(n3), .ZN(n1023) );
  OAI22_X1 U1663 ( .A1(n17), .A2(n1194), .B1(n15), .B2(n1193), .ZN(n986) );
  INV_X1 U1664 ( .A(n608), .ZN(n609) );
  OAI22_X1 U1665 ( .A1(n30), .A2(n1142), .B1(n28), .B2(n1141), .ZN(n936) );
  OAI22_X1 U1666 ( .A1(n36), .A2(n1443), .B1(n34), .B2(n1122), .ZN(n918) );
  INV_X1 U1667 ( .A(n793), .ZN(n850) );
  OAI22_X1 U1668 ( .A1(n60), .A2(n1032), .B1(n58), .B2(n1031), .ZN(n831) );
  AOI21_X1 U1669 ( .B1(n54), .B2(n52), .A(n1051), .ZN(n793) );
  OAI22_X1 U1670 ( .A1(n1166), .A2(n1276), .B1(n21), .B2(n1165), .ZN(n959) );
  OAI22_X1 U1671 ( .A1(n29), .A2(n1147), .B1(n27), .B2(n1146), .ZN(n941) );
  OAI22_X1 U1672 ( .A1(n1185), .A2(n18), .B1(n16), .B2(n1184), .ZN(n977) );
  OAI22_X1 U1673 ( .A1(n17), .A2(n1196), .B1(n15), .B2(n1195), .ZN(n988) );
  OAI22_X1 U1674 ( .A1(n18), .A2(n1297), .B1(n1197), .B2(n16), .ZN(n827) );
  XNOR2_X1 U1675 ( .A(n1485), .B(n1442), .ZN(n1196) );
  AOI21_X1 U1676 ( .B1(n42), .B2(n40), .A(n1093), .ZN(n799) );
  AOI21_X1 U1677 ( .B1(n6), .B2(n4), .A(n1219), .ZN(n817) );
  OAI22_X1 U1678 ( .A1(n54), .A2(n1053), .B1(n52), .B2(n1052), .ZN(n851) );
  INV_X1 U1679 ( .A(n796), .ZN(n870) );
  AOI21_X1 U1680 ( .B1(n48), .B2(n46), .A(n1072), .ZN(n796) );
  AOI21_X1 U1681 ( .B1(n12), .B2(n10), .A(n1198), .ZN(n814) );
  AOI21_X1 U1682 ( .B1(n36), .B2(n34), .A(n1114), .ZN(n802) );
  OAI22_X1 U1683 ( .A1(n53), .A2(n1291), .B1(n1071), .B2(n52), .ZN(n821) );
  OAI22_X1 U1684 ( .A1(n53), .A2(n1070), .B1(n51), .B2(n1069), .ZN(n868) );
  OR2_X1 U1685 ( .A1(n1489), .A2(n1291), .ZN(n1071) );
  NAND2_X1 U1686 ( .A1(n1029), .A2(n829), .ZN(n409) );
  AND2_X1 U1687 ( .A1(n1490), .A2(n818), .ZN(product[0]) );
  INV_X1 U1688 ( .A(n3), .ZN(n818) );
  OAI22_X1 U1689 ( .A1(n60), .A2(n1040), .B1(n57), .B2(n1039), .ZN(n839) );
  INV_X1 U1690 ( .A(n805), .ZN(n930) );
  AOI21_X1 U1691 ( .B1(n30), .B2(n28), .A(n1135), .ZN(n805) );
  OAI22_X1 U1692 ( .A1(n30), .A2(n1138), .B1(n28), .B2(n1137), .ZN(n932) );
  OAI22_X1 U1693 ( .A1(n36), .A2(n1119), .B1(n34), .B2(n1118), .ZN(n914) );
  OAI22_X1 U1694 ( .A1(n42), .A2(n1100), .B1(n40), .B2(n1099), .ZN(n896) );
  OAI22_X1 U1695 ( .A1(n1428), .A2(n1058), .B1(n52), .B2(n1057), .ZN(n856) );
  OAI22_X1 U1696 ( .A1(n60), .A2(n1039), .B1(n58), .B2(n1038), .ZN(n838) );
  OAI22_X1 U1697 ( .A1(n42), .A2(n1096), .B1(n40), .B2(n1095), .ZN(n892) );
  OAI22_X1 U1698 ( .A1(n53), .A2(n1061), .B1(n51), .B2(n1060), .ZN(n859) );
  OAI22_X1 U1699 ( .A1(n30), .A2(n1137), .B1(n28), .B2(n1136), .ZN(n931) );
  OAI22_X1 U1700 ( .A1(n35), .A2(n1118), .B1(n34), .B2(n1117), .ZN(n913) );
  OAI22_X1 U1701 ( .A1(n54), .A2(n1057), .B1(n52), .B2(n1056), .ZN(n855) );
  OAI22_X1 U1702 ( .A1(n48), .A2(n1076), .B1(n46), .B2(n1075), .ZN(n873) );
  OAI22_X1 U1703 ( .A1(n12), .A2(n1204), .B1(n10), .B2(n1203), .ZN(n995) );
  OAI22_X1 U1704 ( .A1(n35), .A2(n1128), .B1(n33), .B2(n1127), .ZN(n923) );
  OAI22_X1 U1705 ( .A1(n47), .A2(n1090), .B1(n45), .B2(n1089), .ZN(n887) );
  OAI22_X1 U1706 ( .A1(n1439), .A2(n1201), .B1(n10), .B2(n1200), .ZN(n992) );
  OAI22_X1 U1707 ( .A1(n18), .A2(n1182), .B1(n1181), .B2(n16), .ZN(n974) );
  OAI22_X1 U1708 ( .A1(n36), .A2(n1125), .B1(n33), .B2(n1444), .ZN(n920) );
  OAI22_X1 U1709 ( .A1(n48), .A2(n1080), .B1(n46), .B2(n1079), .ZN(n877) );
  OAI22_X1 U1710 ( .A1(n42), .A2(n1099), .B1(n40), .B2(n1098), .ZN(n895) );
  AND2_X1 U1711 ( .A1(n1441), .A2(n791), .ZN(n849) );
  OAI22_X1 U1712 ( .A1(n5), .A2(n1221), .B1(n1220), .B2(n4), .ZN(n1012) );
  OAI22_X1 U1713 ( .A1(n47), .A2(n1088), .B1(n1087), .B2(n45), .ZN(n885) );
  OAI22_X1 U1714 ( .A1(n30), .A2(n1141), .B1(n28), .B2(n1140), .ZN(n935) );
  OAI22_X1 U1715 ( .A1(n41), .A2(n1103), .B1(n39), .B2(n1102), .ZN(n899) );
  OAI22_X1 U1716 ( .A1(n47), .A2(n1084), .B1(n45), .B2(n1083), .ZN(n881) );
  OAI22_X1 U1717 ( .A1(n24), .A2(n1162), .B1(n22), .B2(n1161), .ZN(n955) );
  OAI22_X1 U1718 ( .A1(n18), .A2(n1181), .B1(n16), .B2(n1421), .ZN(n973) );
  OAI22_X1 U1719 ( .A1(n54), .A2(n1059), .B1(n52), .B2(n1058), .ZN(n857) );
  OAI22_X1 U1720 ( .A1(n48), .A2(n1078), .B1(n46), .B2(n1077), .ZN(n875) );
  OAI22_X1 U1721 ( .A1(n36), .A2(n1116), .B1(n34), .B2(n1115), .ZN(n911) );
  OAI22_X1 U1722 ( .A1(n24), .A2(n1165), .B1(n22), .B2(n1164), .ZN(n958) );
  OAI22_X1 U1723 ( .A1(n18), .A2(n1430), .B1(n1183), .B2(n16), .ZN(n976) );
  OAI22_X1 U1724 ( .A1(n1440), .A2(n1209), .B1(n9), .B2(n1208), .ZN(n1000) );
  OAI22_X1 U1725 ( .A1(n23), .A2(n1171), .B1(n21), .B2(n1170), .ZN(n964) );
  AND2_X1 U1726 ( .A1(n1442), .A2(n794), .ZN(n869) );
  OAI22_X1 U1727 ( .A1(n1223), .A2(n6), .B1(n1222), .B2(n4), .ZN(n1014) );
  OAI22_X1 U1728 ( .A1(n41), .A2(n1109), .B1(n39), .B2(n1108), .ZN(n905) );
  OAI22_X1 U1729 ( .A1(n1440), .A2(n1202), .B1(n10), .B2(n1201), .ZN(n993) );
  OAI22_X1 U1730 ( .A1(n54), .A2(n1069), .B1(n51), .B2(n1068), .ZN(n867) );
  OAI22_X1 U1731 ( .A1(n41), .A2(n1107), .B1(n39), .B2(n1106), .ZN(n903) );
  OAI22_X1 U1732 ( .A1(n30), .A2(n1140), .B1(n28), .B2(n1139), .ZN(n934) );
  OAI22_X1 U1733 ( .A1(n24), .A2(n1159), .B1(n22), .B2(n1158), .ZN(n952) );
  OAI22_X1 U1734 ( .A1(n47), .A2(n1083), .B1(n45), .B2(n1082), .ZN(n880) );
  INV_X1 U1735 ( .A(n1419), .ZN(n1297) );
  INV_X1 U1736 ( .A(n27), .ZN(n806) );
  INV_X1 U1737 ( .A(n21), .ZN(n809) );
  OAI22_X1 U1738 ( .A1(n11), .A2(n1211), .B1(n9), .B2(n1210), .ZN(n1002) );
  OAI22_X1 U1739 ( .A1(n23), .A2(n1173), .B1(n21), .B2(n1172), .ZN(n966) );
  OAI22_X1 U1740 ( .A1(n17), .A2(n1192), .B1(n15), .B2(n1191), .ZN(n984) );
  OAI22_X1 U1741 ( .A1(n29), .A2(n1150), .B1(n27), .B2(n1149), .ZN(n944) );
  OAI22_X1 U1742 ( .A1(n35), .A2(n1131), .B1(n33), .B2(n1130), .ZN(n926) );
  OAI22_X1 U1743 ( .A1(n17), .A2(n1188), .B1(n15), .B2(n1187), .ZN(n980) );
  OAI22_X1 U1744 ( .A1(n18), .A2(n1180), .B1(n16), .B2(n1179), .ZN(n972) );
  OAI22_X1 U1745 ( .A1(n41), .A2(n1104), .B1(n1103), .B2(n39), .ZN(n900) );
  OAI22_X1 U1746 ( .A1(n59), .A2(n1047), .B1(n57), .B2(n1046), .ZN(n846) );
  OAI22_X1 U1747 ( .A1(n1428), .A2(n1064), .B1(n51), .B2(n1063), .ZN(n862) );
  OAI22_X1 U1748 ( .A1(n36), .A2(n1121), .B1(n34), .B2(n1120), .ZN(n916) );
  OAI22_X1 U1749 ( .A1(n60), .A2(n1045), .B1(n57), .B2(n1044), .ZN(n844) );
  OAI22_X1 U1750 ( .A1(n36), .A2(n1122), .B1(n34), .B2(n1121), .ZN(n917) );
  OAI22_X1 U1751 ( .A1(n35), .A2(n1129), .B1(n33), .B2(n1128), .ZN(n924) );
  OAI22_X1 U1752 ( .A1(n23), .A2(n1167), .B1(n21), .B2(n1166), .ZN(n960) );
  OAI22_X1 U1753 ( .A1(n41), .A2(n1110), .B1(n1109), .B2(n39), .ZN(n906) );
  OAI22_X1 U1754 ( .A1(n42), .A2(n1098), .B1(n40), .B2(n1097), .ZN(n894) );
  OAI22_X1 U1755 ( .A1(n48), .A2(n1079), .B1(n46), .B2(n1078), .ZN(n876) );
  OAI22_X1 U1756 ( .A1(n36), .A2(n1117), .B1(n34), .B2(n1116), .ZN(n912) );
  OAI22_X1 U1757 ( .A1(n1439), .A2(n1210), .B1(n9), .B2(n1209), .ZN(n1001) );
  OAI22_X1 U1758 ( .A1(n17), .A2(n1191), .B1(n15), .B2(n1190), .ZN(n983) );
  OAI22_X1 U1759 ( .A1(n29), .A2(n1153), .B1(n27), .B2(n1152), .ZN(n947) );
  OAI22_X1 U1760 ( .A1(n24), .A2(n1164), .B1(n22), .B2(n1163), .ZN(n957) );
  AND2_X1 U1761 ( .A1(n1490), .A2(n800), .ZN(n909) );
  OAI22_X1 U1762 ( .A1(n1412), .A2(n1227), .B1(n1226), .B2(n4), .ZN(n1018) );
  OAI22_X1 U1763 ( .A1(n29), .A2(n1151), .B1(n27), .B2(n1150), .ZN(n945) );
  OAI22_X1 U1764 ( .A1(n60), .A2(n1044), .B1(n57), .B2(n1043), .ZN(n843) );
  INV_X1 U1765 ( .A(n811), .ZN(n970) );
  AOI21_X1 U1766 ( .B1(n18), .B2(n16), .A(n1177), .ZN(n811) );
  OAI22_X1 U1767 ( .A1(n23), .A2(n1168), .B1(n21), .B2(n1167), .ZN(n961) );
  OAI22_X1 U1768 ( .A1(n17), .A2(n1187), .B1(n15), .B2(n1186), .ZN(n979) );
  OAI22_X1 U1769 ( .A1(n1439), .A2(n1212), .B1(n9), .B2(n1211), .ZN(n1003) );
  OAI22_X1 U1770 ( .A1(n23), .A2(n1174), .B1(n21), .B2(n1173), .ZN(n967) );
  OAI22_X1 U1771 ( .A1(n59), .A2(n1042), .B1(n57), .B2(n1041), .ZN(n841) );
  INV_X1 U1772 ( .A(n808), .ZN(n950) );
  AOI21_X1 U1773 ( .B1(n24), .B2(n22), .A(n1156), .ZN(n808) );
  OAI22_X1 U1774 ( .A1(n1412), .A2(n1224), .B1(n1223), .B2(n4), .ZN(n1015) );
  OAI22_X1 U1775 ( .A1(n29), .A2(n1148), .B1(n27), .B2(n1147), .ZN(n942) );
  OAI22_X1 U1776 ( .A1(n18), .A2(n1186), .B1(n16), .B2(n1185), .ZN(n978) );
  OAI22_X1 U1777 ( .A1(n5), .A2(n1230), .B1(n1229), .B2(n3), .ZN(n1021) );
  OAI22_X1 U1778 ( .A1(n42), .A2(n1102), .B1(n40), .B2(n1101), .ZN(n898) );
  INV_X1 U1779 ( .A(n574), .ZN(n575) );
  OAI22_X1 U1780 ( .A1(n11), .A2(n1205), .B1(n10), .B2(n1204), .ZN(n996) );
  OAI22_X1 U1781 ( .A1(n42), .A2(n1101), .B1(n40), .B2(n1100), .ZN(n897) );
  OAI22_X1 U1782 ( .A1(n47), .A2(n1082), .B1(n45), .B2(n1081), .ZN(n879) );
  OAI22_X1 U1783 ( .A1(n36), .A2(n1120), .B1(n34), .B2(n1119), .ZN(n915) );
  OAI22_X1 U1784 ( .A1(n1428), .A2(n1062), .B1(n51), .B2(n1061), .ZN(n860) );
  OAI22_X1 U1785 ( .A1(n48), .A2(n1081), .B1(n46), .B2(n1080), .ZN(n878) );
  OAI22_X1 U1786 ( .A1(n60), .A2(n1043), .B1(n57), .B2(n1042), .ZN(n842) );
  AND2_X1 U1787 ( .A1(n1441), .A2(n797), .ZN(n889) );
  OAI22_X1 U1788 ( .A1(n6), .A2(n1225), .B1(n1224), .B2(n4), .ZN(n1016) );
  OAI22_X1 U1789 ( .A1(n35), .A2(n1130), .B1(n33), .B2(n1129), .ZN(n925) );
  AND2_X1 U1790 ( .A1(n1442), .A2(n803), .ZN(n929) );
  OAI22_X1 U1791 ( .A1(n1412), .A2(n1229), .B1(n1228), .B2(n3), .ZN(n1020) );
  OAI22_X1 U1792 ( .A1(n23), .A2(n1172), .B1(n21), .B2(n1171), .ZN(n965) );
  OAI22_X1 U1793 ( .A1(n29), .A2(n1145), .B1(n27), .B2(n1144), .ZN(n939) );
  OAI22_X1 U1794 ( .A1(n35), .A2(n1126), .B1(n33), .B2(n1125), .ZN(n921) );
  OAI22_X1 U1795 ( .A1(n18), .A2(n1183), .B1(n1182), .B2(n16), .ZN(n975) );
  AND2_X1 U1796 ( .A1(n1442), .A2(n809), .ZN(n969) );
  OAI22_X1 U1797 ( .A1(n1440), .A2(n1214), .B1(n9), .B2(n1213), .ZN(n1005) );
  OAI22_X1 U1798 ( .A1(n1412), .A2(n1233), .B1(n1232), .B2(n3), .ZN(n1024) );
  OAI22_X1 U1799 ( .A1(n1439), .A2(n1206), .B1(n10), .B2(n1205), .ZN(n997) );
  OAI22_X1 U1800 ( .A1(n29), .A2(n1149), .B1(n27), .B2(n1148), .ZN(n943) );
  OAI22_X1 U1801 ( .A1(n41), .A2(n1111), .B1(n39), .B2(n1110), .ZN(n907) );
  OAI22_X1 U1802 ( .A1(n48), .A2(n1077), .B1(n46), .B2(n1076), .ZN(n874) );
  INV_X1 U1803 ( .A(n496), .ZN(n497) );
  OAI22_X1 U1804 ( .A1(n36), .A2(n1127), .B1(n33), .B2(n1126), .ZN(n922) );
  OAI22_X1 U1805 ( .A1(n47), .A2(n1089), .B1(n45), .B2(n1088), .ZN(n886) );
  OAI22_X1 U1806 ( .A1(n41), .A2(n1108), .B1(n39), .B2(n1107), .ZN(n904) );
  OAI22_X1 U1807 ( .A1(n11), .A2(n1207), .B1(n10), .B2(n1206), .ZN(n998) );
  OAI22_X1 U1808 ( .A1(n1412), .A2(n1226), .B1(n1225), .B2(n4), .ZN(n1017) );
  OAI22_X1 U1809 ( .A1(n23), .A2(n1169), .B1(n21), .B2(n1168), .ZN(n962) );
  OAI22_X1 U1810 ( .A1(n1439), .A2(n1208), .B1(n9), .B2(n1207), .ZN(n999) );
  OAI22_X1 U1811 ( .A1(n23), .A2(n1170), .B1(n21), .B2(n1169), .ZN(n963) );
  OAI22_X1 U1812 ( .A1(n36), .A2(n1132), .B1(n33), .B2(n1131), .ZN(n927) );
  OAI22_X1 U1813 ( .A1(n48), .A2(n1074), .B1(n46), .B2(n1073), .ZN(n871) );
  INV_X1 U1814 ( .A(n814), .ZN(n990) );
  OAI22_X1 U1815 ( .A1(n18), .A2(n1450), .B1(n1178), .B2(n16), .ZN(n971) );
  OAI22_X1 U1816 ( .A1(n59), .A2(n1427), .B1(n57), .B2(n1045), .ZN(n845) );
  AND2_X1 U1817 ( .A1(n1442), .A2(n806), .ZN(n949) );
  OAI22_X1 U1818 ( .A1(n1412), .A2(n1231), .B1(n1230), .B2(n3), .ZN(n1022) );
  OAI22_X1 U1819 ( .A1(n17), .A2(n1193), .B1(n15), .B2(n1192), .ZN(n985) );
  OAI22_X1 U1820 ( .A1(n42), .A2(n1097), .B1(n40), .B2(n1096), .ZN(n893) );
  OAI22_X1 U1821 ( .A1(n1428), .A2(n1060), .B1(n52), .B2(n1059), .ZN(n858) );
  OAI22_X1 U1822 ( .A1(n60), .A2(n1041), .B1(n57), .B2(n1040), .ZN(n840) );
  INV_X1 U1823 ( .A(n518), .ZN(n519) );
  OAI22_X1 U1824 ( .A1(n1428), .A2(n1056), .B1(n52), .B2(n1055), .ZN(n854) );
  OAI22_X1 U1825 ( .A1(n48), .A2(n1075), .B1(n46), .B2(n1074), .ZN(n872) );
  OAI22_X1 U1826 ( .A1(n60), .A2(n1037), .B1(n58), .B2(n1036), .ZN(n836) );
  OAI22_X1 U1827 ( .A1(n12), .A2(n1200), .B1(n10), .B2(n1199), .ZN(n991) );
  OAI22_X1 U1828 ( .A1(n47), .A2(n1423), .B1(n45), .B2(n1085), .ZN(n883) );
  OAI22_X1 U1829 ( .A1(n41), .A2(n1105), .B1(n39), .B2(n1104), .ZN(n901) );
  OAI22_X1 U1830 ( .A1(n1440), .A2(n1203), .B1(n10), .B2(n1202), .ZN(n994) );
  OAI22_X1 U1831 ( .A1(n5), .A2(n1222), .B1(n1221), .B2(n4), .ZN(n1013) );
  OAI22_X1 U1832 ( .A1(n29), .A2(n1146), .B1(n27), .B2(n1145), .ZN(n940) );
  OAI22_X1 U1833 ( .A1(n17), .A2(n1189), .B1(n15), .B2(n1188), .ZN(n981) );
  OAI22_X1 U1834 ( .A1(n5), .A2(n1220), .B1(n1451), .B2(n4), .ZN(n1011) );
  OAI22_X1 U1835 ( .A1(n41), .A2(n1106), .B1(n39), .B2(n1105), .ZN(n902) );
  OAI22_X1 U1836 ( .A1(n24), .A2(n1163), .B1(n22), .B2(n1162), .ZN(n956) );
  OAI22_X1 U1837 ( .A1(n1412), .A2(n1228), .B1(n1227), .B2(n4), .ZN(n1019) );
  OAI22_X1 U1838 ( .A1(n29), .A2(n1152), .B1(n27), .B2(n1151), .ZN(n946) );
  OAI22_X1 U1839 ( .A1(n17), .A2(n1190), .B1(n15), .B2(n1189), .ZN(n982) );
  OAI22_X1 U1840 ( .A1(n53), .A2(n1066), .B1(n51), .B2(n1065), .ZN(n864) );
  OAI22_X1 U1841 ( .A1(n47), .A2(n1085), .B1(n45), .B2(n1084), .ZN(n882) );
  OAI22_X1 U1842 ( .A1(n24), .A2(n1161), .B1(n22), .B2(n1160), .ZN(n954) );
  INV_X1 U1843 ( .A(n1486), .ZN(n1292) );
  NAND2_X1 U1844 ( .A1(n787), .A2(n788), .ZN(n400) );
  OAI22_X1 U1845 ( .A1(n42), .A2(n1293), .B1(n1113), .B2(n40), .ZN(n823) );
  OAI22_X1 U1846 ( .A1(n1112), .A2(n41), .B1(n39), .B2(n1111), .ZN(n908) );
  OR2_X1 U1847 ( .A1(n1489), .A2(n1293), .ZN(n1113) );
  AND2_X1 U1848 ( .A1(n1490), .A2(n815), .ZN(n1009) );
  INV_X1 U1849 ( .A(n9), .ZN(n815) );
  INV_X1 U1850 ( .A(n790), .ZN(n830) );
  AOI21_X1 U1851 ( .B1(n60), .B2(n58), .A(n1030), .ZN(n790) );
  OAI22_X1 U1852 ( .A1(n1428), .A2(n1054), .B1(n52), .B2(n1053), .ZN(n852) );
  OAI22_X1 U1853 ( .A1(n60), .A2(n1035), .B1(n58), .B2(n1034), .ZN(n834) );
  INV_X1 U1854 ( .A(n464), .ZN(n465) );
  OR2_X1 U1855 ( .A1(n1490), .A2(n1296), .ZN(n1176) );
  OR2_X1 U1856 ( .A1(n1490), .A2(n1290), .ZN(n1050) );
  OR2_X1 U1857 ( .A1(n1442), .A2(n1297), .ZN(n1197) );
  OR2_X1 U1858 ( .A1(n1490), .A2(n1295), .ZN(n1155) );
  OR2_X1 U1859 ( .A1(n1489), .A2(n1292), .ZN(n1092) );
  OR2_X1 U1860 ( .A1(n1442), .A2(n1294), .ZN(n1134) );
  OAI22_X1 U1861 ( .A1(n54), .A2(n1055), .B1(n52), .B2(n1054), .ZN(n853) );
  OAI22_X1 U1862 ( .A1(n60), .A2(n1036), .B1(n58), .B2(n1035), .ZN(n835) );
  INV_X1 U1863 ( .A(n799), .ZN(n890) );
  OAI22_X1 U1864 ( .A1(n1124), .A2(n35), .B1(n1123), .B2(n33), .ZN(n919) );
  OAI22_X1 U1865 ( .A1(n1048), .A2(n59), .B1(n1387), .B2(n57), .ZN(n847) );
  INV_X1 U1866 ( .A(n817), .ZN(n1010) );
  OAI22_X1 U1867 ( .A1(n42), .A2(n1095), .B1(n40), .B2(n1094), .ZN(n891) );
  OAI22_X1 U1868 ( .A1(n60), .A2(n1038), .B1(n58), .B2(n1037), .ZN(n837) );
  INV_X1 U1869 ( .A(n802), .ZN(n910) );
  INV_X1 U1870 ( .A(n45), .ZN(n797) );
  INV_X1 U1871 ( .A(n39), .ZN(n800) );
  INV_X1 U1872 ( .A(n51), .ZN(n794) );
  INV_X1 U1873 ( .A(n57), .ZN(n791) );
  INV_X1 U1874 ( .A(n15), .ZN(n812) );
  INV_X1 U1875 ( .A(n33), .ZN(n803) );
  XNOR2_X1 U1876 ( .A(n1485), .B(n1255), .ZN(n1192) );
  XNOR2_X1 U1877 ( .A(n1418), .B(n1254), .ZN(n1191) );
  XNOR2_X1 U1878 ( .A(n1484), .B(n1449), .ZN(n1194) );
  XNOR2_X1 U1879 ( .A(n1419), .B(n1252), .ZN(n1189) );
  XNOR2_X1 U1880 ( .A(n1488), .B(n1242), .ZN(n1074) );
  OAI22_X1 U1881 ( .A1(n5), .A2(n1299), .B1(n1239), .B2(n4), .ZN(n829) );
  INV_X1 U1882 ( .A(n1), .ZN(n1299) );
  OAI22_X1 U1883 ( .A1(n11), .A2(n1298), .B1(n1218), .B2(n10), .ZN(n828) );
  OR2_X1 U1884 ( .A1(n1441), .A2(n1298), .ZN(n1218) );
  INV_X1 U1885 ( .A(n7), .ZN(n1298) );
  OAI22_X1 U1886 ( .A1(n1412), .A2(n1238), .B1(n1237), .B2(n3), .ZN(n1029) );
  OAI22_X1 U1887 ( .A1(n29), .A2(n1154), .B1(n27), .B2(n1153), .ZN(n948) );
  OAI22_X1 U1888 ( .A1(n30), .A2(n1295), .B1(n1155), .B2(n28), .ZN(n825) );
  XNOR2_X1 U1889 ( .A(n1425), .B(n1441), .ZN(n1154) );
  XNOR2_X1 U1890 ( .A(n1487), .B(n1252), .ZN(n1084) );
  XNOR2_X1 U1891 ( .A(n1256), .B(n1486), .ZN(n1088) );
  XNOR2_X1 U1892 ( .A(n1487), .B(n1253), .ZN(n1085) );
  XNOR2_X1 U1893 ( .A(n1486), .B(n1255), .ZN(n1087) );
  XNOR2_X1 U1894 ( .A(n1487), .B(n1422), .ZN(n1072) );
  OAI22_X1 U1895 ( .A1(n1439), .A2(n1217), .B1(n9), .B2(n1216), .ZN(n1008) );
  OAI22_X1 U1896 ( .A1(n1412), .A2(n1236), .B1(n1235), .B2(n3), .ZN(n1027) );
  XNOR2_X1 U1897 ( .A(n7), .B(n1490), .ZN(n1217) );
  XNOR2_X1 U1898 ( .A(n1242), .B(n1484), .ZN(n1179) );
  XNOR2_X1 U1899 ( .A(n1484), .B(n1243), .ZN(n1180) );
  XNOR2_X1 U1900 ( .A(n1484), .B(n1241), .ZN(n1178) );
  XNOR2_X1 U1901 ( .A(n1240), .B(n1484), .ZN(n1177) );
  XNOR2_X1 U1902 ( .A(n1425), .B(n1258), .ZN(n1153) );
  XNOR2_X1 U1903 ( .A(n7), .B(n1253), .ZN(n1211) );
  XNOR2_X1 U1904 ( .A(n7), .B(n1254), .ZN(n1212) );
  XNOR2_X1 U1905 ( .A(n1425), .B(n1244), .ZN(n1139) );
  XNOR2_X1 U1906 ( .A(n1425), .B(n1243), .ZN(n1138) );
  XNOR2_X1 U1907 ( .A(n1425), .B(n1245), .ZN(n1140) );
  XNOR2_X1 U1908 ( .A(n25), .B(n1242), .ZN(n1137) );
  XNOR2_X1 U1909 ( .A(n1425), .B(n1246), .ZN(n1141) );
  XNOR2_X1 U1910 ( .A(n1425), .B(n1247), .ZN(n1142) );
  XNOR2_X1 U1911 ( .A(n7), .B(n1246), .ZN(n1204) );
  XNOR2_X1 U1912 ( .A(n7), .B(n1247), .ZN(n1205) );
  XNOR2_X1 U1913 ( .A(n7), .B(n1255), .ZN(n1213) );
  XNOR2_X1 U1914 ( .A(n7), .B(n1252), .ZN(n1210) );
  XNOR2_X1 U1915 ( .A(n25), .B(n1241), .ZN(n1136) );
  XNOR2_X1 U1916 ( .A(n25), .B(n1248), .ZN(n1143) );
  XNOR2_X1 U1917 ( .A(n25), .B(n1252), .ZN(n1147) );
  XNOR2_X1 U1918 ( .A(n7), .B(n1241), .ZN(n1199) );
  XNOR2_X1 U1919 ( .A(n1424), .B(n1253), .ZN(n1148) );
  XNOR2_X1 U1920 ( .A(n7), .B(n1245), .ZN(n1203) );
  XNOR2_X1 U1921 ( .A(n25), .B(n1251), .ZN(n1146) );
  XNOR2_X1 U1922 ( .A(n7), .B(n1248), .ZN(n1206) );
  XNOR2_X1 U1923 ( .A(n1425), .B(n1254), .ZN(n1149) );
  XNOR2_X1 U1924 ( .A(n7), .B(n1244), .ZN(n1202) );
  XNOR2_X1 U1925 ( .A(n7), .B(n1251), .ZN(n1209) );
  XNOR2_X1 U1926 ( .A(n1425), .B(n1257), .ZN(n1152) );
  XNOR2_X1 U1927 ( .A(n7), .B(n1242), .ZN(n1200) );
  XNOR2_X1 U1928 ( .A(n7), .B(n1256), .ZN(n1214) );
  XNOR2_X1 U1929 ( .A(n1425), .B(n1250), .ZN(n1145) );
  XNOR2_X1 U1930 ( .A(n25), .B(n1255), .ZN(n1150) );
  XNOR2_X1 U1931 ( .A(n7), .B(n1249), .ZN(n1207) );
  XNOR2_X1 U1932 ( .A(n7), .B(n1243), .ZN(n1201) );
  XNOR2_X1 U1933 ( .A(n1250), .B(n7), .ZN(n1208) );
  XNOR2_X1 U1934 ( .A(n1424), .B(n1256), .ZN(n1151) );
  XNOR2_X1 U1935 ( .A(n7), .B(n1257), .ZN(n1215) );
  XNOR2_X1 U1936 ( .A(n25), .B(n1249), .ZN(n1144) );
  XNOR2_X1 U1937 ( .A(n7), .B(n1258), .ZN(n1216) );
  XNOR2_X1 U1938 ( .A(n55), .B(n1256), .ZN(n1046) );
  XNOR2_X1 U1939 ( .A(n1257), .B(n55), .ZN(n1047) );
  XNOR2_X1 U1940 ( .A(n19), .B(n1241), .ZN(n1157) );
  XNOR2_X1 U1941 ( .A(n31), .B(n1246), .ZN(n1120) );
  XNOR2_X1 U1942 ( .A(n55), .B(n1254), .ZN(n1044) );
  XNOR2_X1 U1943 ( .A(n1383), .B(n1257), .ZN(n1173) );
  XNOR2_X1 U1944 ( .A(n31), .B(n1245), .ZN(n1119) );
  XNOR2_X1 U1945 ( .A(n55), .B(n1253), .ZN(n1043) );
  XNOR2_X1 U1946 ( .A(n1383), .B(n1243), .ZN(n1159) );
  XNOR2_X1 U1947 ( .A(n1383), .B(n1258), .ZN(n1174) );
  XNOR2_X1 U1948 ( .A(n55), .B(n1244), .ZN(n1034) );
  XNOR2_X1 U1949 ( .A(n1383), .B(n1242), .ZN(n1158) );
  XNOR2_X1 U1950 ( .A(n55), .B(n1255), .ZN(n1045) );
  XNOR2_X1 U1951 ( .A(n31), .B(n1244), .ZN(n1118) );
  XNOR2_X1 U1952 ( .A(n55), .B(n1252), .ZN(n1042) );
  XNOR2_X1 U1953 ( .A(n55), .B(n1245), .ZN(n1035) );
  XNOR2_X1 U1954 ( .A(n55), .B(n1243), .ZN(n1033) );
  XNOR2_X1 U1955 ( .A(n19), .B(n1244), .ZN(n1160) );
  XNOR2_X1 U1956 ( .A(n55), .B(n1246), .ZN(n1036) );
  XNOR2_X1 U1957 ( .A(n31), .B(n1247), .ZN(n1121) );
  XNOR2_X1 U1958 ( .A(n55), .B(n1251), .ZN(n1041) );
  XNOR2_X1 U1959 ( .A(n1462), .B(n1241), .ZN(n1115) );
  XNOR2_X1 U1960 ( .A(n31), .B(n1249), .ZN(n1123) );
  XNOR2_X1 U1961 ( .A(n55), .B(n1248), .ZN(n1038) );
  XNOR2_X1 U1962 ( .A(n31), .B(n1243), .ZN(n1117) );
  XNOR2_X1 U1963 ( .A(n55), .B(n1414), .ZN(n1040) );
  XNOR2_X1 U1964 ( .A(n55), .B(n1247), .ZN(n1037) );
  XNOR2_X1 U1965 ( .A(n31), .B(n1242), .ZN(n1116) );
  XNOR2_X1 U1966 ( .A(n55), .B(n1470), .ZN(n1039) );
  XNOR2_X1 U1967 ( .A(n19), .B(n1249), .ZN(n1165) );
  XNOR2_X1 U1968 ( .A(n1383), .B(n1251), .ZN(n1167) );
  XNOR2_X1 U1969 ( .A(n1383), .B(n1256), .ZN(n1172) );
  XNOR2_X1 U1970 ( .A(n1250), .B(n19), .ZN(n1166) );
  XNOR2_X1 U1971 ( .A(n31), .B(n1254), .ZN(n1128) );
  XNOR2_X1 U1972 ( .A(n31), .B(n1248), .ZN(n1122) );
  XNOR2_X1 U1973 ( .A(n55), .B(n1242), .ZN(n1032) );
  XNOR2_X1 U1974 ( .A(n31), .B(n1253), .ZN(n1127) );
  XNOR2_X1 U1975 ( .A(n31), .B(n1255), .ZN(n1129) );
  XNOR2_X1 U1976 ( .A(n1383), .B(n1248), .ZN(n1164) );
  XNOR2_X1 U1977 ( .A(n1383), .B(n1252), .ZN(n1168) );
  XNOR2_X1 U1978 ( .A(n31), .B(n1256), .ZN(n1130) );
  XNOR2_X1 U1979 ( .A(n31), .B(n1250), .ZN(n1124) );
  XNOR2_X1 U1980 ( .A(n55), .B(n1258), .ZN(n1048) );
  XNOR2_X1 U1981 ( .A(n31), .B(n1252), .ZN(n1126) );
  XNOR2_X1 U1982 ( .A(n1383), .B(n1247), .ZN(n1163) );
  XNOR2_X1 U1983 ( .A(n31), .B(n1257), .ZN(n1131) );
  XNOR2_X1 U1984 ( .A(n1383), .B(n1253), .ZN(n1169) );
  XNOR2_X1 U1985 ( .A(n1383), .B(n1246), .ZN(n1162) );
  XNOR2_X1 U1986 ( .A(n1383), .B(n1254), .ZN(n1170) );
  XNOR2_X1 U1987 ( .A(n19), .B(n1245), .ZN(n1161) );
  XNOR2_X1 U1988 ( .A(n31), .B(n1258), .ZN(n1132) );
  XNOR2_X1 U1989 ( .A(n31), .B(n1251), .ZN(n1125) );
  XNOR2_X1 U1990 ( .A(n19), .B(n1255), .ZN(n1171) );
  XNOR2_X1 U1991 ( .A(n55), .B(n1241), .ZN(n1031) );
  XNOR2_X1 U1992 ( .A(n1487), .B(n1250), .ZN(n1082) );
  XNOR2_X1 U1993 ( .A(n1488), .B(n1249), .ZN(n1081) );
  XNOR2_X1 U1994 ( .A(n1487), .B(n1251), .ZN(n1083) );
  XNOR2_X1 U1995 ( .A(n1488), .B(n1241), .ZN(n1073) );
  XNOR2_X1 U1996 ( .A(n1487), .B(n1244), .ZN(n1076) );
  XNOR2_X1 U1997 ( .A(n1488), .B(n1248), .ZN(n1080) );
  XNOR2_X1 U1998 ( .A(n1487), .B(n1245), .ZN(n1077) );
  XNOR2_X1 U1999 ( .A(n1487), .B(n1247), .ZN(n1079) );
  XNOR2_X1 U2000 ( .A(n1487), .B(n1246), .ZN(n1078) );
  XNOR2_X1 U2001 ( .A(n1488), .B(n1243), .ZN(n1075) );
  XNOR2_X1 U2002 ( .A(n1486), .B(n1258), .ZN(n1090) );
  XNOR2_X1 U2003 ( .A(n1257), .B(n1486), .ZN(n1089) );
  XNOR2_X1 U2004 ( .A(n1487), .B(n1254), .ZN(n1086) );
  XNOR2_X1 U2005 ( .A(n1418), .B(n1256), .ZN(n1193) );
  XNOR2_X1 U2006 ( .A(n1484), .B(n1247), .ZN(n1184) );
  XNOR2_X1 U2007 ( .A(n1418), .B(n1249), .ZN(n1186) );
  XNOR2_X1 U2008 ( .A(n1418), .B(n1248), .ZN(n1185) );
  XNOR2_X1 U2009 ( .A(n1485), .B(n1246), .ZN(n1183) );
  XNOR2_X1 U2010 ( .A(n1419), .B(n1250), .ZN(n1187) );
  XNOR2_X1 U2011 ( .A(n1418), .B(n1251), .ZN(n1188) );
  XNOR2_X1 U2012 ( .A(n1419), .B(n1258), .ZN(n1195) );
  XNOR2_X1 U2013 ( .A(n1485), .B(n1253), .ZN(n1190) );
  XNOR2_X1 U2014 ( .A(n1485), .B(n1244), .ZN(n1181) );
  XNOR2_X1 U2015 ( .A(n1485), .B(n1245), .ZN(n1182) );
  XNOR2_X1 U2016 ( .A(n1240), .B(n1424), .ZN(n1135) );
  XNOR2_X1 U2017 ( .A(n7), .B(n1240), .ZN(n1198) );
  XNOR2_X1 U2018 ( .A(n19), .B(n1240), .ZN(n1156) );
  XNOR2_X1 U2019 ( .A(n1462), .B(n1240), .ZN(n1114) );
  XNOR2_X1 U2020 ( .A(n1413), .B(n1429), .ZN(n1030) );
  BUF_X1 U2021 ( .A(n1288), .Z(n9) );
  BUF_X1 U2022 ( .A(n1288), .Z(n10) );
  BUF_X1 U2023 ( .A(n1281), .Z(n52) );
  BUF_X1 U2024 ( .A(n1271), .Z(n54) );
  BUF_X1 U2025 ( .A(n61), .Z(n1490) );
  BUF_X1 U2026 ( .A(n1279), .Z(n5) );
  OAI22_X1 U2027 ( .A1(n36), .A2(n1133), .B1(n33), .B2(n1132), .ZN(n928) );
  OAI22_X1 U2028 ( .A1(n36), .A2(n1294), .B1(n1134), .B2(n34), .ZN(n824) );
  XNOR2_X1 U2029 ( .A(n31), .B(n1441), .ZN(n1133) );
  OAI22_X1 U2030 ( .A1(n23), .A2(n1175), .B1(n21), .B2(n1174), .ZN(n968) );
  OAI22_X1 U2031 ( .A1(n24), .A2(n1296), .B1(n1176), .B2(n22), .ZN(n826) );
  XNOR2_X1 U2032 ( .A(n1383), .B(n1441), .ZN(n1175) );
  OAI22_X1 U2033 ( .A1(n59), .A2(n1049), .B1(n57), .B2(n1415), .ZN(n848) );
  OAI22_X1 U2034 ( .A1(n59), .A2(n1290), .B1(n1050), .B2(n58), .ZN(n820) );
  XNOR2_X1 U2035 ( .A(n55), .B(n1442), .ZN(n1049) );
  INV_X1 U2036 ( .A(n37), .ZN(n1293) );
  BUF_X2 U2037 ( .A(n1275), .Z(n30) );
  BUF_X2 U2038 ( .A(n1276), .Z(n24) );
  BUF_X2 U2039 ( .A(n1275), .Z(n29) );
  INV_X1 U2040 ( .A(n1425), .ZN(n1295) );
  INV_X1 U2041 ( .A(n1383), .ZN(n1296) );
  INV_X1 U2042 ( .A(n31), .ZN(n1294) );
  INV_X1 U2043 ( .A(n55), .ZN(n1290) );
  BUF_X1 U2044 ( .A(n1289), .Z(n3) );
  BUF_X1 U2045 ( .A(n1289), .Z(n4) );
  BUF_X2 U2046 ( .A(n1273), .Z(n42) );
  BUF_X1 U2047 ( .A(n1272), .Z(n48) );
  INV_X1 U2048 ( .A(n49), .ZN(n1291) );
  XNOR2_X1 U2049 ( .A(a[9]), .B(a[10]), .ZN(n1284) );
  XNOR2_X1 U2050 ( .A(a[16]), .B(a[15]), .ZN(n1281) );
  XNOR2_X1 U2051 ( .A(a[18]), .B(a[17]), .ZN(n1280) );
  BUF_X4 U2052 ( .A(a[3]), .Z(n7) );
  BUF_X4 U2053 ( .A(a[11]), .Z(n31) );
  XNOR2_X1 U2054 ( .A(a[2]), .B(a[1]), .ZN(n1288) );
  CLKBUF_X3 U2055 ( .A(b[3]), .Z(n1256) );
  BUF_X4 U2056 ( .A(a[1]), .Z(n1) );
  BUF_X1 U2057 ( .A(a[15]), .Z(n43) );
  OAI21_X1 U2058 ( .B1(n1469), .B2(n304), .A(n297), .ZN(n295) );
  XOR2_X1 U2059 ( .A(n142), .B(n69), .Z(product[36]) );
  CLKBUF_X1 U2060 ( .A(n43), .Z(n1488) );
  OAI22_X1 U2061 ( .A1(n1428), .A2(n1052), .B1(n52), .B2(n1051), .ZN(n454) );
  XNOR2_X1 U2062 ( .A(n1448), .B(n1243), .ZN(n1096) );
  XNOR2_X1 U2063 ( .A(n1240), .B(n1448), .ZN(n1093) );
  XNOR2_X1 U2064 ( .A(n1448), .B(n1249), .ZN(n1102) );
  XNOR2_X1 U2065 ( .A(n1448), .B(n1253), .ZN(n1106) );
  XNOR2_X1 U2066 ( .A(n1448), .B(n1242), .ZN(n1095) );
  XNOR2_X1 U2067 ( .A(n1448), .B(n1241), .ZN(n1094) );
  XNOR2_X1 U2068 ( .A(n1448), .B(n1254), .ZN(n1107) );
  XNOR2_X1 U2069 ( .A(n1448), .B(n1245), .ZN(n1098) );
  XNOR2_X1 U2070 ( .A(n1448), .B(n1244), .ZN(n1097) );
  XNOR2_X1 U2071 ( .A(n1448), .B(n1248), .ZN(n1101) );
  XNOR2_X1 U2072 ( .A(n1448), .B(n1252), .ZN(n1105) );
  XNOR2_X1 U2073 ( .A(n1448), .B(n1257), .ZN(n1110) );
  XNOR2_X1 U2074 ( .A(n37), .B(n1256), .ZN(n1109) );
  XNOR2_X1 U2075 ( .A(n37), .B(n1255), .ZN(n1108) );
  XNOR2_X1 U2076 ( .A(n1448), .B(n1247), .ZN(n1100) );
  XNOR2_X1 U2077 ( .A(n1448), .B(n1489), .ZN(n1112) );
  XNOR2_X1 U2078 ( .A(n1448), .B(n1246), .ZN(n1099) );
  XNOR2_X1 U2079 ( .A(n37), .B(n1258), .ZN(n1111) );
  XNOR2_X1 U2080 ( .A(n37), .B(n1251), .ZN(n1104) );
  XNOR2_X1 U2081 ( .A(n1250), .B(n37), .ZN(n1103) );
  XNOR2_X1 U2082 ( .A(a[13]), .B(a[14]), .ZN(n1282) );
  XNOR2_X1 U2083 ( .A(n1445), .B(n1243), .ZN(n1054) );
  XNOR2_X1 U2084 ( .A(n1445), .B(n1247), .ZN(n1058) );
  XNOR2_X1 U2085 ( .A(n1445), .B(n1242), .ZN(n1053) );
  XNOR2_X1 U2086 ( .A(n1388), .B(n1246), .ZN(n1057) );
  XNOR2_X1 U2087 ( .A(n49), .B(n1489), .ZN(n1070) );
  XNOR2_X1 U2088 ( .A(n49), .B(n1253), .ZN(n1064) );
  XNOR2_X1 U2089 ( .A(n1388), .B(n1245), .ZN(n1056) );
  XNOR2_X1 U2090 ( .A(n1445), .B(n1244), .ZN(n1055) );
  XNOR2_X1 U2091 ( .A(n49), .B(n1258), .ZN(n1069) );
  XNOR2_X1 U2092 ( .A(n49), .B(n1252), .ZN(n1063) );
  XNOR2_X1 U2093 ( .A(n1388), .B(n1248), .ZN(n1059) );
  XNOR2_X1 U2094 ( .A(n1257), .B(n49), .ZN(n1068) );
  XNOR2_X1 U2095 ( .A(n49), .B(n1256), .ZN(n1067) );
  XNOR2_X1 U2096 ( .A(n49), .B(n1251), .ZN(n1062) );
  XNOR2_X1 U2097 ( .A(n49), .B(n1250), .ZN(n1061) );
  XNOR2_X1 U2098 ( .A(n49), .B(n1249), .ZN(n1060) );
  XNOR2_X1 U2099 ( .A(n49), .B(n1255), .ZN(n1066) );
  XNOR2_X1 U2100 ( .A(n49), .B(n1254), .ZN(n1065) );
  XNOR2_X1 U2101 ( .A(n1445), .B(n1241), .ZN(n1052) );
  XNOR2_X1 U2102 ( .A(n1445), .B(n1429), .ZN(n1051) );
  NAND2_X1 U2103 ( .A1(n1268), .A2(n1288), .ZN(n1278) );
  CLKBUF_X1 U2104 ( .A(n1278), .Z(n11) );
  OAI21_X1 U2105 ( .B1(n339), .B2(n326), .A(n1477), .ZN(n325) );
  NOR2_X1 U2106 ( .A1(n323), .A2(n326), .ZN(n321) );
  NAND2_X1 U2107 ( .A1(n1028), .A2(n1009), .ZN(n407) );
  XOR2_X1 U2108 ( .A(n388), .B(n98), .Z(product[7]) );
  XOR2_X1 U2109 ( .A(n127), .B(n68), .Z(product[37]) );
  OAI22_X1 U2110 ( .A1(n1412), .A2(n1237), .B1(n1236), .B2(n3), .ZN(n1028) );
  XOR2_X1 U2111 ( .A(a[10]), .B(a[11]), .Z(n1264) );
  XNOR2_X1 U2112 ( .A(a[12]), .B(a[11]), .ZN(n1283) );
  XNOR2_X1 U2113 ( .A(n99), .B(n393), .ZN(product[6]) );
  XNOR2_X1 U2114 ( .A(n1), .B(n1248), .ZN(n1227) );
  XNOR2_X1 U2115 ( .A(n1438), .B(n1251), .ZN(n1230) );
  XNOR2_X1 U2116 ( .A(n1438), .B(n1252), .ZN(n1231) );
  XNOR2_X1 U2117 ( .A(n1), .B(n1247), .ZN(n1226) );
  XNOR2_X1 U2118 ( .A(n1), .B(n1246), .ZN(n1225) );
  XNOR2_X1 U2119 ( .A(n1), .B(n1242), .ZN(n1221) );
  XNOR2_X1 U2120 ( .A(n1), .B(n1241), .ZN(n1220) );
  XNOR2_X1 U2121 ( .A(n1), .B(n1245), .ZN(n1224) );
  XNOR2_X1 U2122 ( .A(n1), .B(n1250), .ZN(n1229) );
  XNOR2_X1 U2123 ( .A(n1), .B(n1249), .ZN(n1228) );
  XNOR2_X1 U2124 ( .A(n1), .B(n1243), .ZN(n1222) );
  XNOR2_X1 U2125 ( .A(n1), .B(n1244), .ZN(n1223) );
  XNOR2_X1 U2126 ( .A(n1), .B(n1253), .ZN(n1232) );
  XNOR2_X1 U2127 ( .A(n1), .B(n1254), .ZN(n1233) );
  XNOR2_X1 U2128 ( .A(n1240), .B(n1), .ZN(n1219) );
  XNOR2_X1 U2129 ( .A(n1), .B(n1255), .ZN(n1234) );
  XNOR2_X1 U2130 ( .A(n1), .B(n1256), .ZN(n1235) );
  XNOR2_X1 U2131 ( .A(n1438), .B(n1441), .ZN(n1238) );
  XNOR2_X1 U2132 ( .A(n1), .B(n1258), .ZN(n1237) );
  XNOR2_X1 U2133 ( .A(n1438), .B(n1257), .ZN(n1236) );
  OAI21_X1 U2134 ( .B1(n1466), .B2(n108), .A(n109), .ZN(n107) );
  OAI21_X1 U2135 ( .B1(n1466), .B2(n117), .A(n118), .ZN(n116) );
  OAI21_X1 U2136 ( .B1(n225), .B2(n65), .A(n226), .ZN(n224) );
  OAI21_X1 U2137 ( .B1(n65), .B2(n242), .A(n243), .ZN(n233) );
  OAI21_X1 U2138 ( .B1(n65), .B2(n216), .A(n217), .ZN(n211) );
  OAI21_X1 U2139 ( .B1(n1453), .B2(n160), .A(n161), .ZN(n159) );
  OAI21_X1 U2140 ( .B1(n1454), .B2(n184), .A(n185), .ZN(n183) );
  OAI21_X1 U2141 ( .B1(n1454), .B2(n145), .A(n146), .ZN(n144) );
  OAI21_X1 U2142 ( .B1(n1453), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U2143 ( .B1(n1454), .B2(n171), .A(n172), .ZN(n170) );
  OAI21_X1 U2144 ( .B1(n1453), .B2(n201), .A(n202), .ZN(n200) );
  XNOR2_X1 U2145 ( .A(a[8]), .B(a[7]), .ZN(n1285) );
  XOR2_X1 U2146 ( .A(a[6]), .B(a[7]), .Z(n1266) );
  XOR2_X1 U2147 ( .A(a[18]), .B(a[19]), .Z(n1260) );
  OAI21_X1 U2148 ( .B1(n361), .B2(n365), .A(n362), .ZN(n360) );
  NOR2_X1 U2149 ( .A1(n361), .A2(n364), .ZN(n359) );
  INV_X1 U2150 ( .A(n361), .ZN(n436) );
  NOR2_X1 U2151 ( .A1(n731), .A2(n740), .ZN(n361) );
  XNOR2_X1 U2152 ( .A(n64), .B(n82), .ZN(product[23]) );
  AOI21_X1 U2153 ( .B1(n63), .B2(n232), .A(n233), .ZN(n231) );
  AOI21_X1 U2154 ( .B1(n64), .B2(n245), .A(n246), .ZN(n244) );
  AOI21_X1 U2155 ( .B1(n64), .B2(n223), .A(n224), .ZN(n222) );
  AOI21_X1 U2156 ( .B1(n63), .B2(n269), .A(n270), .ZN(n268) );
  AOI21_X1 U2157 ( .B1(n63), .B2(n287), .A(n288), .ZN(n286) );
  AOI21_X1 U2158 ( .B1(n357), .B2(n348), .A(n349), .ZN(n347) );
  AOI21_X1 U2159 ( .B1(n349), .B2(n1402), .A(n344), .ZN(n342) );
  XOR2_X1 U2160 ( .A(a[16]), .B(a[17]), .Z(n1261) );
  AOI21_X1 U2161 ( .B1(n1416), .B2(n106), .A(n107), .ZN(n105) );
  AOI21_X1 U2162 ( .B1(n1416), .B2(n115), .A(n116), .ZN(n114) );
  AOI21_X1 U2163 ( .B1(n1386), .B2(n128), .A(n129), .ZN(n127) );
  AOI21_X1 U2164 ( .B1(n63), .B2(n210), .A(n211), .ZN(n209) );
  AOI21_X1 U2165 ( .B1(n64), .B2(n158), .A(n159), .ZN(n157) );
  AOI21_X1 U2166 ( .B1(n64), .B2(n182), .A(n183), .ZN(n181) );
  AOI21_X1 U2167 ( .B1(n64), .B2(n169), .A(n170), .ZN(n168) );
  AOI21_X1 U2168 ( .B1(n1386), .B2(n143), .A(n144), .ZN(n142) );
  AOI21_X1 U2169 ( .B1(n1386), .B2(n199), .A(n200), .ZN(n198) );
  NAND2_X1 U2170 ( .A1(n134), .A2(n1403), .ZN(n121) );
  AOI21_X1 U2171 ( .B1(n63), .B2(n258), .A(n259), .ZN(n257) );
  NAND2_X1 U2172 ( .A1(n759), .A2(n766), .ZN(n378) );
  XOR2_X1 U2173 ( .A(a[9]), .B(a[8]), .Z(n1265) );
  XOR2_X1 U2174 ( .A(a[2]), .B(a[3]), .Z(n1268) );
  XOR2_X1 U2175 ( .A(a[14]), .B(a[15]), .Z(n1262) );
  OAI21_X1 U2176 ( .B1(n350), .B2(n356), .A(n351), .ZN(n349) );
  XOR2_X1 U2177 ( .A(a[12]), .B(a[13]), .Z(n1263) );
  NAND2_X1 U2178 ( .A1(n789), .A2(n828), .ZN(n403) );
  XOR2_X1 U2179 ( .A(a[4]), .B(a[5]), .Z(n1267) );
  XNOR2_X1 U2180 ( .A(a[6]), .B(a[5]), .ZN(n1286) );
  NOR2_X1 U2181 ( .A1(n289), .A2(n284), .ZN(n282) );
  INV_X1 U2182 ( .A(n358), .ZN(n357) );
  XOR2_X1 U2183 ( .A(a[0]), .B(a[1]), .Z(n1269) );
  AOI21_X1 U2184 ( .B1(n63), .B2(n278), .A(n1391), .ZN(n277) );
  OR2_X1 U2185 ( .A1(n1490), .A2(n1299), .ZN(n1239) );
endmodule


module datapath_DW_mult_tc_9 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n3, n4, n6, n7, n9, n10, n11, n12, n13, n15, n16, n18, n21, n22,
         n23, n24, n25, n27, n28, n29, n30, n31, n33, n34, n35, n36, n37, n39,
         n40, n41, n42, n43, n45, n46, n47, n48, n49, n51, n52, n53, n54, n55,
         n57, n58, n59, n60, n61, n63, n64, n65, n67, n68, n69, n70, n71, n72,
         n73, n82, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n105, n106, n107, n108, n109,
         n111, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n124, n126, n127, n128, n129, n130, n131, n134, n135, n136, n137,
         n139, n141, n142, n143, n144, n145, n146, n149, n150, n151, n152,
         n154, n156, n157, n158, n159, n160, n161, n165, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n190, n191, n192, n193,
         n195, n197, n198, n199, n200, n201, n202, n206, n208, n209, n210,
         n211, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n254, n256, n257, n258, n259, n260, n261, n262, n263, n265,
         n267, n268, n269, n270, n271, n273, n274, n275, n276, n277, n278,
         n280, n281, n282, n283, n284, n285, n286, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n303,
         n304, n305, n306, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n331, n332, n333, n334, n339, n340, n341, n342, n344, n346, n347,
         n348, n349, n350, n351, n352, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n371,
         n373, n374, n376, n378, n379, n380, n382, n384, n385, n386, n387,
         n388, n390, n392, n393, n394, n395, n396, n398, n400, n401, n402,
         n403, n404, n405, n406, n407, n409, n418, n424, n425, n428, n430,
         n435, n436, n437, n441, n443, n445, n446, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n793,
         n794, n796, n797, n799, n800, n802, n803, n805, n806, n808, n809,
         n811, n812, n814, n815, n817, n818, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1509, n1510, n1511;
  assign product[39] = n105;

  FA_X1 U488 ( .A(n831), .B(n454), .CI(n850), .CO(n450), .S(n451) );
  FA_X1 U489 ( .A(n455), .B(n832), .CI(n458), .CO(n452), .S(n453) );
  FA_X1 U491 ( .A(n462), .B(n833), .CI(n459), .CO(n456), .S(n457) );
  FA_X1 U492 ( .A(n851), .B(n464), .CI(n870), .CO(n458), .S(n459) );
  FA_X1 U493 ( .A(n463), .B(n470), .CI(n468), .CO(n460), .S(n461) );
  FA_X1 U494 ( .A(n834), .B(n852), .CI(n465), .CO(n462), .S(n463) );
  FA_X1 U496 ( .A(n474), .B(n471), .CI(n469), .CO(n466), .S(n467) );
  FA_X1 U497 ( .A(n478), .B(n871), .CI(n476), .CO(n468), .S(n469) );
  FA_X1 U498 ( .A(n853), .B(n835), .CI(n890), .CO(n470), .S(n471) );
  FA_X1 U499 ( .A(n475), .B(n477), .CI(n482), .CO(n472), .S(n473) );
  FA_X1 U500 ( .A(n486), .B(n479), .CI(n484), .CO(n474), .S(n475) );
  FA_X1 U501 ( .A(n836), .B(n854), .CI(n872), .CO(n476), .S(n477) );
  FA_X1 U503 ( .A(n490), .B(n492), .CI(n483), .CO(n480), .S(n481) );
  FA_X1 U504 ( .A(n485), .B(n494), .CI(n487), .CO(n482), .S(n483) );
  FA_X1 U505 ( .A(n855), .B(n496), .CI(n873), .CO(n484), .S(n485) );
  FA_X1 U506 ( .A(n891), .B(n837), .CI(n910), .CO(n486), .S(n487) );
  FA_X1 U507 ( .A(n500), .B(n493), .CI(n491), .CO(n488), .S(n489) );
  FA_X1 U508 ( .A(n495), .B(n504), .CI(n502), .CO(n490), .S(n491) );
  FA_X1 U509 ( .A(n497), .B(n874), .CI(n506), .CO(n492), .S(n493) );
  FA_X1 U510 ( .A(n892), .B(n856), .CI(n838), .CO(n494), .S(n495) );
  FA_X1 U512 ( .A(n510), .B(n503), .CI(n501), .CO(n498), .S(n499) );
  FA_X1 U513 ( .A(n507), .B(n505), .CI(n512), .CO(n500), .S(n501) );
  FA_X1 U514 ( .A(n516), .B(n893), .CI(n514), .CO(n502), .S(n503) );
  FA_X1 U515 ( .A(n857), .B(n911), .CI(n875), .CO(n504), .S(n505) );
  FA_X1 U516 ( .A(n518), .B(n839), .CI(n930), .CO(n506), .S(n507) );
  FA_X1 U517 ( .A(n522), .B(n513), .CI(n511), .CO(n508), .S(n509) );
  FA_X1 U518 ( .A(n526), .B(n515), .CI(n524), .CO(n510), .S(n511) );
  FA_X1 U519 ( .A(n528), .B(n530), .CI(n517), .CO(n512), .S(n513) );
  FA_X1 U520 ( .A(n840), .B(n858), .CI(n519), .CO(n514), .S(n515) );
  FA_X1 U521 ( .A(n912), .B(n876), .CI(n894), .CO(n516), .S(n517) );
  FA_X1 U523 ( .A(n534), .B(n525), .CI(n523), .CO(n520), .S(n521) );
  FA_X1 U524 ( .A(n527), .B(n538), .CI(n536), .CO(n522), .S(n523) );
  FA_X1 U525 ( .A(n529), .B(n540), .CI(n531), .CO(n524), .S(n525) );
  FA_X1 U526 ( .A(n877), .B(n895), .CI(n542), .CO(n526), .S(n527) );
  FA_X1 U527 ( .A(n859), .B(n931), .CI(n913), .CO(n528), .S(n529) );
  FA_X1 U528 ( .A(n950), .B(n841), .CI(n544), .CO(n530), .S(n531) );
  FA_X1 U529 ( .A(n548), .B(n537), .CI(n535), .CO(n532), .S(n533) );
  FA_X1 U531 ( .A(n541), .B(n554), .CI(n543), .CO(n536), .S(n537) );
  FA_X1 U532 ( .A(n558), .B(n545), .CI(n556), .CO(n538), .S(n539) );
  FA_X1 U533 ( .A(n896), .B(n932), .CI(n914), .CO(n540), .S(n541) );
  FA_X1 U534 ( .A(n842), .B(n878), .CI(n860), .CO(n542), .S(n543) );
  FA_X1 U536 ( .A(n562), .B(n551), .CI(n549), .CO(n546), .S(n547) );
  FA_X1 U538 ( .A(n559), .B(n557), .CI(n568), .CO(n550), .S(n551) );
  FA_X1 U539 ( .A(n570), .B(n572), .CI(n555), .CO(n552), .S(n553) );
  FA_X1 U540 ( .A(n879), .B(n915), .CI(n897), .CO(n554), .S(n555) );
  FA_X1 U541 ( .A(n861), .B(n951), .CI(n933), .CO(n556), .S(n557) );
  FA_X1 U542 ( .A(n574), .B(n843), .CI(n970), .CO(n558), .S(n559) );
  FA_X1 U543 ( .A(n578), .B(n565), .CI(n563), .CO(n560), .S(n561) );
  FA_X1 U544 ( .A(n567), .B(n582), .CI(n580), .CO(n562), .S(n563) );
  FA_X1 U545 ( .A(n584), .B(n573), .CI(n569), .CO(n564), .S(n565) );
  FA_X1 U546 ( .A(n586), .B(n588), .CI(n571), .CO(n566), .S(n567) );
  FA_X1 U547 ( .A(n575), .B(n898), .CI(n590), .CO(n568), .S(n569) );
  FA_X1 U548 ( .A(n844), .B(n916), .CI(n862), .CO(n570), .S(n571) );
  FA_X1 U549 ( .A(n952), .B(n880), .CI(n934), .CO(n572), .S(n573) );
  FA_X1 U551 ( .A(n594), .B(n581), .CI(n579), .CO(n576), .S(n577) );
  FA_X1 U552 ( .A(n583), .B(n598), .CI(n596), .CO(n578), .S(n579) );
  FA_X1 U553 ( .A(n600), .B(n591), .CI(n585), .CO(n580), .S(n581) );
  FA_X1 U554 ( .A(n587), .B(n602), .CI(n589), .CO(n582), .S(n583) );
  FA_X1 U555 ( .A(n606), .B(n917), .CI(n604), .CO(n584), .S(n585) );
  FA_X1 U556 ( .A(n881), .B(n935), .CI(n899), .CO(n586), .S(n587) );
  FA_X1 U557 ( .A(n608), .B(n953), .CI(n863), .CO(n588), .S(n589) );
  FA_X1 U558 ( .A(n845), .B(n971), .CI(n990), .CO(n590), .S(n591) );
  FA_X1 U559 ( .A(n612), .B(n597), .CI(n595), .CO(n592), .S(n593) );
  FA_X1 U560 ( .A(n599), .B(n616), .CI(n614), .CO(n594), .S(n595) );
  FA_X1 U561 ( .A(n618), .B(n603), .CI(n601), .CO(n596), .S(n597) );
  FA_X1 U562 ( .A(n605), .B(n620), .CI(n607), .CO(n598), .S(n599) );
  FA_X1 U563 ( .A(n626), .B(n624), .CI(n622), .CO(n600), .S(n601) );
  FA_X1 U564 ( .A(n918), .B(n936), .CI(n609), .CO(n602), .S(n603) );
  FA_X1 U565 ( .A(n864), .B(n954), .CI(n882), .CO(n604), .S(n605) );
  FA_X1 U568 ( .A(n630), .B(n615), .CI(n613), .CO(n610), .S(n611) );
  FA_X1 U569 ( .A(n617), .B(n634), .CI(n632), .CO(n612), .S(n613) );
  FA_X1 U570 ( .A(n636), .B(n621), .CI(n619), .CO(n614), .S(n615) );
  FA_X1 U571 ( .A(n623), .B(n638), .CI(n625), .CO(n616), .S(n617) );
  FA_X1 U572 ( .A(n642), .B(n627), .CI(n640), .CO(n618), .S(n619) );
  FA_X1 U573 ( .A(n955), .B(n973), .CI(n644), .CO(n620), .S(n621) );
  FA_X1 U574 ( .A(n883), .B(n901), .CI(n991), .CO(n622), .S(n623) );
  FA_X1 U575 ( .A(n919), .B(n847), .CI(n1010), .CO(n624), .S(n625) );
  FA_X1 U579 ( .A(n650), .B(n637), .CI(n635), .CO(n630), .S(n631) );
  FA_X1 U580 ( .A(n654), .B(n643), .CI(n652), .CO(n632), .S(n633) );
  FA_X1 U581 ( .A(n639), .B(n656), .CI(n641), .CO(n634), .S(n635) );
  FA_X1 U582 ( .A(n660), .B(n645), .CI(n658), .CO(n636), .S(n637) );
  FA_X1 U583 ( .A(n920), .B(n992), .CI(n974), .CO(n638), .S(n639) );
  FA_X1 U584 ( .A(n956), .B(n902), .CI(n1011), .CO(n640), .S(n641) );
  HA_X1 U586 ( .A(n848), .B(n820), .CO(n644), .S(n645) );
  FA_X1 U588 ( .A(n653), .B(n655), .CI(n666), .CO(n648), .S(n649) );
  FA_X1 U589 ( .A(n670), .B(n659), .CI(n668), .CO(n650), .S(n651) );
  FA_X1 U590 ( .A(n661), .B(n672), .CI(n657), .CO(n652), .S(n653) );
  FA_X1 U591 ( .A(n676), .B(n957), .CI(n674), .CO(n654), .S(n655) );
  FA_X1 U592 ( .A(n975), .B(n921), .CI(n939), .CO(n656), .S(n657) );
  FA_X1 U593 ( .A(n867), .B(n993), .CI(n903), .CO(n658), .S(n659) );
  FA_X1 U594 ( .A(n849), .B(n1012), .CI(n885), .CO(n660), .S(n661) );
  FA_X1 U595 ( .A(n667), .B(n680), .CI(n665), .CO(n662), .S(n663) );
  FA_X1 U596 ( .A(n682), .B(n671), .CI(n669), .CO(n664), .S(n665) );
  FA_X1 U597 ( .A(n675), .B(n673), .CI(n684), .CO(n666), .S(n667) );
  FA_X1 U598 ( .A(n686), .B(n690), .CI(n688), .CO(n668), .S(n669) );
  FA_X1 U599 ( .A(n958), .B(n976), .CI(n677), .CO(n670), .S(n671) );
  FA_X1 U600 ( .A(n886), .B(n904), .CI(n922), .CO(n672), .S(n673) );
  FA_X1 U601 ( .A(n1013), .B(n940), .CI(n994), .CO(n674), .S(n675) );
  HA_X1 U602 ( .A(n821), .B(n868), .CO(n676), .S(n677) );
  FA_X1 U603 ( .A(n694), .B(n683), .CI(n681), .CO(n678), .S(n679) );
  FA_X1 U604 ( .A(n685), .B(n698), .CI(n696), .CO(n680), .S(n681) );
  FA_X1 U605 ( .A(n689), .B(n691), .CI(n687), .CO(n682), .S(n683) );
  FA_X1 U606 ( .A(n702), .B(n704), .CI(n700), .CO(n684), .S(n685) );
  FA_X1 U607 ( .A(n977), .B(n959), .CI(n941), .CO(n686), .S(n687) );
  FA_X1 U608 ( .A(n887), .B(n995), .CI(n923), .CO(n688), .S(n689) );
  FA_X1 U609 ( .A(n869), .B(n1014), .CI(n905), .CO(n690), .S(n691) );
  FA_X1 U610 ( .A(n697), .B(n708), .CI(n695), .CO(n692), .S(n693) );
  FA_X1 U611 ( .A(n710), .B(n703), .CI(n699), .CO(n694), .S(n695) );
  FA_X1 U612 ( .A(n701), .B(n714), .CI(n712), .CO(n696), .S(n697) );
  FA_X1 U613 ( .A(n705), .B(n996), .CI(n716), .CO(n698), .S(n699) );
  FA_X1 U614 ( .A(n1015), .B(n942), .CI(n978), .CO(n700), .S(n701) );
  FA_X1 U615 ( .A(n924), .B(n906), .CI(n960), .CO(n702), .S(n703) );
  HA_X1 U616 ( .A(n822), .B(n888), .CO(n704), .S(n705) );
  FA_X1 U617 ( .A(n711), .B(n720), .CI(n709), .CO(n706), .S(n707) );
  FA_X1 U618 ( .A(n713), .B(n715), .CI(n722), .CO(n708), .S(n709) );
  FA_X1 U619 ( .A(n724), .B(n726), .CI(n717), .CO(n710), .S(n711) );
  FA_X1 U620 ( .A(n961), .B(n979), .CI(n728), .CO(n712), .S(n713) );
  FA_X1 U621 ( .A(n907), .B(n997), .CI(n943), .CO(n714), .S(n715) );
  FA_X1 U622 ( .A(n889), .B(n1016), .CI(n925), .CO(n716), .S(n717) );
  FA_X1 U623 ( .A(n732), .B(n723), .CI(n721), .CO(n718), .S(n719) );
  FA_X1 U624 ( .A(n727), .B(n725), .CI(n734), .CO(n720), .S(n721) );
  FA_X1 U625 ( .A(n738), .B(n729), .CI(n736), .CO(n722), .S(n723) );
  FA_X1 U626 ( .A(n926), .B(n980), .CI(n944), .CO(n724), .S(n725) );
  FA_X1 U627 ( .A(n1017), .B(n962), .CI(n998), .CO(n726), .S(n727) );
  HA_X1 U628 ( .A(n823), .B(n908), .CO(n728), .S(n729) );
  FA_X1 U629 ( .A(n735), .B(n742), .CI(n733), .CO(n730), .S(n731) );
  FA_X1 U630 ( .A(n737), .B(n739), .CI(n744), .CO(n732), .S(n733) );
  FA_X1 U631 ( .A(n748), .B(n981), .CI(n746), .CO(n734), .S(n735) );
  FA_X1 U632 ( .A(n927), .B(n999), .CI(n963), .CO(n736), .S(n737) );
  FA_X1 U633 ( .A(n945), .B(n909), .CI(n1018), .CO(n738), .S(n739) );
  FA_X1 U634 ( .A(n752), .B(n745), .CI(n743), .CO(n740), .S(n741) );
  FA_X1 U635 ( .A(n754), .B(n756), .CI(n747), .CO(n742), .S(n743) );
  FA_X1 U636 ( .A(n964), .B(n1000), .CI(n749), .CO(n744), .S(n745) );
  FA_X1 U637 ( .A(n946), .B(n982), .CI(n1019), .CO(n746), .S(n747) );
  HA_X1 U638 ( .A(n824), .B(n928), .CO(n748), .S(n749) );
  FA_X1 U639 ( .A(n760), .B(n755), .CI(n753), .CO(n750), .S(n751) );
  FA_X1 U640 ( .A(n762), .B(n764), .CI(n757), .CO(n752), .S(n753) );
  FA_X1 U641 ( .A(n947), .B(n1001), .CI(n983), .CO(n754), .S(n755) );
  FA_X1 U642 ( .A(n965), .B(n929), .CI(n1020), .CO(n756), .S(n757) );
  FA_X1 U643 ( .A(n763), .B(n768), .CI(n761), .CO(n758), .S(n759) );
  FA_X1 U644 ( .A(n765), .B(n1021), .CI(n770), .CO(n760), .S(n761) );
  FA_X1 U645 ( .A(n966), .B(n984), .CI(n1002), .CO(n762), .S(n763) );
  HA_X1 U646 ( .A(n825), .B(n948), .CO(n764), .S(n765) );
  FA_X1 U647 ( .A(n771), .B(n774), .CI(n769), .CO(n766), .S(n767) );
  FA_X1 U648 ( .A(n967), .B(n1003), .CI(n776), .CO(n768), .S(n769) );
  FA_X1 U649 ( .A(n985), .B(n949), .CI(n1022), .CO(n770), .S(n771) );
  FA_X1 U650 ( .A(n780), .B(n777), .CI(n775), .CO(n772), .S(n773) );
  FA_X1 U651 ( .A(n986), .B(n1023), .CI(n1004), .CO(n774), .S(n775) );
  HA_X1 U652 ( .A(n826), .B(n968), .CO(n776), .S(n777) );
  FA_X1 U653 ( .A(n784), .B(n987), .CI(n781), .CO(n778), .S(n779) );
  FA_X1 U654 ( .A(n1024), .B(n969), .CI(n1005), .CO(n780), .S(n781) );
  FA_X1 U655 ( .A(n1006), .B(n1025), .CI(n785), .CO(n782), .S(n783) );
  HA_X1 U656 ( .A(n827), .B(n988), .CO(n784), .S(n785) );
  FA_X1 U657 ( .A(n1026), .B(n989), .CI(n1007), .CO(n786), .S(n787) );
  HA_X1 U658 ( .A(n1008), .B(n1027), .CO(n788), .S(n789) );
  INV_X1 U1180 ( .A(n800), .ZN(n1383) );
  CLKBUF_X1 U1181 ( .A(n312), .Z(n1384) );
  CLKBUF_X3 U1182 ( .A(b[11]), .Z(n1248) );
  CLKBUF_X3 U1183 ( .A(b[7]), .Z(n1252) );
  CLKBUF_X1 U1184 ( .A(n64), .Z(n1385) );
  CLKBUF_X3 U1185 ( .A(b[12]), .Z(n1247) );
  CLKBUF_X3 U1186 ( .A(b[17]), .Z(n1242) );
  CLKBUF_X3 U1187 ( .A(b[3]), .Z(n1256) );
  CLKBUF_X3 U1188 ( .A(b[10]), .Z(n1249) );
  CLKBUF_X3 U1189 ( .A(b[2]), .Z(n1257) );
  CLKBUF_X3 U1190 ( .A(b[4]), .Z(n1255) );
  BUF_X1 U1191 ( .A(n1272), .Z(n47) );
  BUF_X2 U1192 ( .A(b[13]), .Z(n1246) );
  BUF_X2 U1193 ( .A(b[6]), .Z(n1253) );
  BUF_X1 U1194 ( .A(n1272), .Z(n48) );
  BUF_X2 U1195 ( .A(a[19]), .Z(n1450) );
  BUF_X2 U1196 ( .A(n61), .Z(n1506) );
  OR2_X1 U1197 ( .A1(n663), .A2(n678), .ZN(n1503) );
  BUF_X2 U1198 ( .A(n61), .Z(n1507) );
  NOR2_X1 U1199 ( .A1(n547), .A2(n560), .ZN(n284) );
  BUF_X2 U1200 ( .A(n61), .Z(n1511) );
  BUF_X2 U1201 ( .A(a[7]), .Z(n1510) );
  NAND2_X2 U1202 ( .A1(n282), .A2(n249), .ZN(n247) );
  NOR2_X1 U1203 ( .A1(n296), .A2(n303), .ZN(n1386) );
  BUF_X2 U1204 ( .A(n1272), .Z(n1387) );
  CLKBUF_X2 U1205 ( .A(n1282), .Z(n46) );
  BUF_X1 U1206 ( .A(n1284), .Z(n34) );
  CLKBUF_X1 U1207 ( .A(a[0]), .Z(n1388) );
  CLKBUF_X1 U1208 ( .A(n1251), .Z(n1389) );
  NOR2_X2 U1209 ( .A1(n251), .A2(n275), .ZN(n249) );
  CLKBUF_X3 U1210 ( .A(b[1]), .Z(n1258) );
  CLKBUF_X1 U1211 ( .A(n1246), .Z(n1390) );
  XNOR2_X1 U1212 ( .A(n1391), .B(n900), .ZN(n607) );
  XNOR2_X1 U1213 ( .A(n972), .B(n846), .ZN(n1391) );
  BUF_X2 U1214 ( .A(n1274), .Z(n35) );
  AND2_X1 U1215 ( .A1(n663), .A2(n678), .ZN(n1456) );
  BUF_X1 U1216 ( .A(n1277), .Z(n18) );
  BUF_X2 U1217 ( .A(b[8]), .Z(n1251) );
  OAI22_X1 U1218 ( .A1(n1068), .A2(n53), .B1(n1466), .B2(n51), .ZN(n866) );
  BUF_X2 U1219 ( .A(n1273), .Z(n41) );
  BUF_X2 U1220 ( .A(b[15]), .Z(n1244) );
  NOR2_X1 U1221 ( .A1(n789), .A2(n828), .ZN(n402) );
  OAI22_X1 U1222 ( .A1(n1429), .A2(n1031), .B1(n58), .B2(n1030), .ZN(n448) );
  BUF_X2 U1223 ( .A(n291), .Z(n64) );
  INV_X1 U1224 ( .A(n1456), .ZN(n331) );
  XNOR2_X1 U1225 ( .A(n1424), .B(n1244), .ZN(n1392) );
  CLKBUF_X1 U1226 ( .A(n1257), .Z(n1393) );
  BUF_X1 U1227 ( .A(n1285), .Z(n27) );
  BUF_X1 U1228 ( .A(n1285), .Z(n28) );
  BUF_X1 U1229 ( .A(n320), .Z(n1470) );
  XNOR2_X1 U1230 ( .A(n564), .B(n1394), .ZN(n549) );
  XNOR2_X1 U1231 ( .A(n553), .B(n566), .ZN(n1394) );
  OAI22_X1 U1232 ( .A1(n29), .A2(n1144), .B1(n1143), .B2(n28), .ZN(n938) );
  BUF_X2 U1233 ( .A(n1275), .Z(n29) );
  XOR2_X1 U1234 ( .A(n648), .B(n633), .Z(n1395) );
  XOR2_X1 U1235 ( .A(n631), .B(n1395), .Z(n629) );
  NAND2_X1 U1236 ( .A1(n631), .A2(n648), .ZN(n1396) );
  NAND2_X1 U1237 ( .A1(n631), .A2(n633), .ZN(n1397) );
  NAND2_X1 U1238 ( .A1(n648), .A2(n633), .ZN(n1398) );
  NAND3_X1 U1239 ( .A1(n1396), .A2(n1397), .A3(n1398), .ZN(n628) );
  XOR2_X1 U1240 ( .A(n664), .B(n651), .Z(n1399) );
  XOR2_X1 U1241 ( .A(n649), .B(n1399), .Z(n647) );
  NAND2_X1 U1242 ( .A1(n649), .A2(n664), .ZN(n1400) );
  NAND2_X1 U1243 ( .A1(n649), .A2(n651), .ZN(n1401) );
  NAND2_X1 U1244 ( .A1(n664), .A2(n651), .ZN(n1402) );
  NAND3_X1 U1245 ( .A1(n1400), .A2(n1401), .A3(n1402), .ZN(n646) );
  OR2_X1 U1246 ( .A1(n473), .A2(n480), .ZN(n1403) );
  OR2_X1 U1247 ( .A1(n453), .A2(n456), .ZN(n1404) );
  OR2_X1 U1248 ( .A1(n467), .A2(n472), .ZN(n1405) );
  OR2_X1 U1249 ( .A1(n830), .A2(n448), .ZN(n1406) );
  OR2_X1 U1250 ( .A1(n679), .A2(n692), .ZN(n1407) );
  OR2_X1 U1251 ( .A1(n452), .A2(n451), .ZN(n1408) );
  OR2_X1 U1252 ( .A1(n693), .A2(n706), .ZN(n1409) );
  OR2_X1 U1253 ( .A1(n759), .A2(n766), .ZN(n1410) );
  OR2_X1 U1254 ( .A1(n450), .A2(n449), .ZN(n1411) );
  OR2_X1 U1255 ( .A1(n457), .A2(n460), .ZN(n1412) );
  OR2_X1 U1256 ( .A1(n767), .A2(n772), .ZN(n1413) );
  OR2_X1 U1257 ( .A1(n779), .A2(n782), .ZN(n1414) );
  OR2_X1 U1258 ( .A1(n787), .A2(n788), .ZN(n1415) );
  OR2_X1 U1259 ( .A1(n707), .A2(n718), .ZN(n1416) );
  OR2_X1 U1260 ( .A1(n1029), .A2(n829), .ZN(n1417) );
  OR2_X1 U1261 ( .A1(n1480), .A2(n592), .ZN(n1418) );
  AND2_X1 U1262 ( .A1(n679), .A2(n692), .ZN(n1425) );
  OAI21_X1 U1263 ( .B1(n284), .B2(n290), .A(n285), .ZN(n1419) );
  XNOR2_X1 U1264 ( .A(n1424), .B(n1242), .ZN(n1420) );
  CLKBUF_X1 U1265 ( .A(n1282), .Z(n45) );
  CLKBUF_X1 U1266 ( .A(n1288), .Z(n9) );
  BUF_X2 U1267 ( .A(b[16]), .Z(n1243) );
  BUF_X1 U1268 ( .A(n1279), .Z(n6) );
  CLKBUF_X1 U1269 ( .A(n1240), .Z(n1421) );
  XNOR2_X1 U1270 ( .A(n1), .B(n1240), .ZN(n1422) );
  BUF_X2 U1271 ( .A(a[1]), .Z(n1) );
  XNOR2_X1 U1272 ( .A(n1), .B(n1241), .ZN(n1423) );
  BUF_X2 U1273 ( .A(a[1]), .Z(n1424) );
  BUF_X1 U1274 ( .A(b[0]), .Z(n61) );
  OR2_X1 U1275 ( .A1(n1384), .A2(n317), .ZN(n1426) );
  INV_X1 U1276 ( .A(n41), .ZN(n1427) );
  INV_X1 U1277 ( .A(n1427), .ZN(n1428) );
  BUF_X2 U1278 ( .A(n1277), .Z(n1462) );
  BUF_X1 U1279 ( .A(n1270), .Z(n1429) );
  BUF_X2 U1280 ( .A(n1270), .Z(n1430) );
  CLKBUF_X1 U1281 ( .A(n1270), .Z(n59) );
  CLKBUF_X1 U1282 ( .A(n1503), .Z(n1431) );
  CLKBUF_X1 U1283 ( .A(n313), .Z(n1432) );
  BUF_X2 U1284 ( .A(a[11]), .Z(n31) );
  BUF_X1 U1285 ( .A(a[11]), .Z(n1465) );
  XOR2_X1 U1286 ( .A(n866), .B(n938), .Z(n1433) );
  XOR2_X1 U1287 ( .A(n884), .B(n1433), .Z(n643) );
  NAND2_X1 U1288 ( .A1(n884), .A2(n866), .ZN(n1434) );
  NAND2_X1 U1289 ( .A1(n884), .A2(n938), .ZN(n1435) );
  NAND2_X1 U1290 ( .A1(n866), .A2(n938), .ZN(n1436) );
  NAND3_X1 U1291 ( .A1(n1434), .A2(n1435), .A3(n1436), .ZN(n642) );
  BUF_X2 U1292 ( .A(b[19]), .Z(n1240) );
  CLKBUF_X1 U1293 ( .A(n593), .Z(n1437) );
  BUF_X2 U1294 ( .A(b[18]), .Z(n1241) );
  CLKBUF_X1 U1295 ( .A(n64), .Z(n1438) );
  CLKBUF_X1 U1296 ( .A(n1384), .Z(n1439) );
  BUF_X1 U1297 ( .A(n1273), .Z(n42) );
  BUF_X2 U1298 ( .A(b[14]), .Z(n1245) );
  CLKBUF_X1 U1299 ( .A(n1283), .Z(n40) );
  CLKBUF_X3 U1300 ( .A(a[19]), .Z(n55) );
  OR2_X1 U1301 ( .A1(n1437), .A2(n610), .ZN(n1440) );
  XNOR2_X1 U1302 ( .A(n298), .B(n1441), .ZN(product[22]) );
  AND2_X1 U1303 ( .A1(n1418), .A2(n1447), .ZN(n1441) );
  BUF_X2 U1304 ( .A(n1274), .Z(n1442) );
  XNOR2_X1 U1305 ( .A(n1250), .B(n31), .ZN(n1443) );
  CLKBUF_X1 U1306 ( .A(n340), .Z(n1444) );
  CLKBUF_X1 U1307 ( .A(n304), .Z(n1445) );
  AOI21_X2 U1308 ( .B1(n1419), .B2(n249), .A(n250), .ZN(n1446) );
  AOI21_X1 U1309 ( .B1(n283), .B2(n249), .A(n250), .ZN(n248) );
  CLKBUF_X1 U1310 ( .A(n297), .Z(n1447) );
  BUF_X2 U1311 ( .A(n1279), .Z(n1448) );
  CLKBUF_X1 U1312 ( .A(n1279), .Z(n1449) );
  XNOR2_X1 U1313 ( .A(n1465), .B(n1249), .ZN(n1451) );
  BUF_X1 U1314 ( .A(n1465), .Z(n1499) );
  XNOR2_X1 U1315 ( .A(n43), .B(n1254), .ZN(n1452) );
  XNOR2_X1 U1316 ( .A(n1450), .B(n1258), .ZN(n1453) );
  XNOR2_X1 U1317 ( .A(n49), .B(n1257), .ZN(n1454) );
  XNOR2_X1 U1318 ( .A(n1257), .B(n1450), .ZN(n1455) );
  XNOR2_X1 U1319 ( .A(n43), .B(n1255), .ZN(n1457) );
  CLKBUF_X1 U1320 ( .A(n311), .Z(n1458) );
  CLKBUF_X1 U1321 ( .A(n248), .Z(n65) );
  XNOR2_X1 U1322 ( .A(n1250), .B(n31), .ZN(n1459) );
  NOR2_X1 U1323 ( .A1(n647), .A2(n662), .ZN(n1460) );
  NOR2_X1 U1324 ( .A1(n647), .A2(n662), .ZN(n323) );
  XNOR2_X1 U1325 ( .A(n49), .B(n1256), .ZN(n1461) );
  BUF_X1 U1326 ( .A(n1277), .Z(n1463) );
  XNOR2_X1 U1327 ( .A(n305), .B(n1464), .ZN(product[21]) );
  AND2_X1 U1328 ( .A1(n1440), .A2(n1445), .ZN(n1464) );
  CLKBUF_X2 U1329 ( .A(n1284), .Z(n33) );
  XNOR2_X1 U1330 ( .A(n49), .B(n1256), .ZN(n1466) );
  BUF_X1 U1331 ( .A(n1274), .Z(n36) );
  CLKBUF_X1 U1332 ( .A(n43), .Z(n1467) );
  CLKBUF_X1 U1333 ( .A(n49), .Z(n1468) );
  BUF_X1 U1334 ( .A(n574), .Z(n1469) );
  BUF_X2 U1335 ( .A(n1281), .Z(n52) );
  BUF_X2 U1336 ( .A(n1281), .Z(n51) );
  CLKBUF_X1 U1337 ( .A(n39), .Z(n1471) );
  BUF_X2 U1338 ( .A(n39), .Z(n1472) );
  CLKBUF_X1 U1339 ( .A(n39), .Z(n1473) );
  NAND2_X1 U1340 ( .A1(n564), .A2(n553), .ZN(n1474) );
  NAND2_X1 U1341 ( .A1(n564), .A2(n566), .ZN(n1475) );
  NAND2_X1 U1342 ( .A1(n553), .A2(n566), .ZN(n1476) );
  NAND3_X1 U1343 ( .A1(n1474), .A2(n1475), .A3(n1476), .ZN(n548) );
  OR2_X2 U1344 ( .A1(n509), .A2(n520), .ZN(n1477) );
  XNOR2_X1 U1345 ( .A(n244), .B(n1478), .ZN(product[28]) );
  AND2_X1 U1346 ( .A1(n240), .A2(n243), .ZN(n1478) );
  NOR2_X1 U1347 ( .A1(n707), .A2(n718), .ZN(n1479) );
  NOR2_X1 U1348 ( .A1(n707), .A2(n718), .ZN(n350) );
  CLKBUF_X1 U1349 ( .A(n577), .Z(n1480) );
  XOR2_X1 U1350 ( .A(n539), .B(n552), .Z(n1481) );
  XOR2_X1 U1351 ( .A(n550), .B(n1481), .Z(n535) );
  NAND2_X1 U1352 ( .A1(n550), .A2(n539), .ZN(n1482) );
  NAND2_X1 U1353 ( .A1(n550), .A2(n552), .ZN(n1483) );
  NAND2_X1 U1354 ( .A1(n539), .A2(n552), .ZN(n1484) );
  NAND3_X1 U1355 ( .A1(n1482), .A2(n1483), .A3(n1484), .ZN(n534) );
  CLKBUF_X1 U1356 ( .A(n1421), .Z(n1485) );
  NOR2_X1 U1357 ( .A1(n593), .A2(n610), .ZN(n303) );
  NOR2_X1 U1358 ( .A1(n611), .A2(n628), .ZN(n1486) );
  NOR2_X1 U1359 ( .A1(n611), .A2(n628), .ZN(n312) );
  BUF_X2 U1360 ( .A(n1275), .Z(n30) );
  NOR2_X1 U1361 ( .A1(n577), .A2(n592), .ZN(n1487) );
  NOR2_X1 U1362 ( .A1(n577), .A2(n592), .ZN(n296) );
  XNOR2_X1 U1363 ( .A(n277), .B(n1488), .ZN(product[25]) );
  AND2_X1 U1364 ( .A1(n273), .A2(n276), .ZN(n1488) );
  XNOR2_X1 U1365 ( .A(n257), .B(n1489), .ZN(product[27]) );
  AND2_X1 U1366 ( .A1(n1477), .A2(n256), .ZN(n1489) );
  XNOR2_X1 U1367 ( .A(n286), .B(n1490), .ZN(product[24]) );
  AND2_X1 U1368 ( .A1(n424), .A2(n285), .ZN(n1490) );
  BUF_X2 U1369 ( .A(n1280), .Z(n57) );
  AOI21_X1 U1370 ( .B1(n1431), .B2(n1425), .A(n1456), .ZN(n1491) );
  OR2_X1 U1371 ( .A1(n521), .A2(n532), .ZN(n1492) );
  XNOR2_X1 U1372 ( .A(n268), .B(n1493), .ZN(product[26]) );
  AND2_X1 U1373 ( .A1(n262), .A2(n267), .ZN(n1493) );
  CLKBUF_X1 U1374 ( .A(n1257), .Z(n1494) );
  BUF_X2 U1375 ( .A(n1271), .Z(n53) );
  OR2_X2 U1376 ( .A1(n751), .A2(n758), .ZN(n1495) );
  NAND2_X1 U1377 ( .A1(n900), .A2(n972), .ZN(n1496) );
  NAND2_X1 U1378 ( .A1(n900), .A2(n846), .ZN(n1497) );
  NAND2_X1 U1379 ( .A1(n972), .A2(n846), .ZN(n1498) );
  NAND3_X1 U1380 ( .A1(n1496), .A2(n1497), .A3(n1498), .ZN(n606) );
  CLKBUF_X2 U1381 ( .A(n1287), .Z(n16) );
  CLKBUF_X1 U1382 ( .A(n1258), .Z(n1500) );
  NOR2_X2 U1383 ( .A1(n731), .A2(n740), .ZN(n361) );
  BUF_X2 U1384 ( .A(n1286), .Z(n21) );
  BUF_X2 U1385 ( .A(n1278), .Z(n12) );
  XNOR2_X1 U1386 ( .A(n222), .B(n1501), .ZN(product[30]) );
  AND2_X1 U1387 ( .A1(n418), .A2(n221), .ZN(n1501) );
  BUF_X1 U1388 ( .A(n1286), .Z(n22) );
  BUF_X2 U1389 ( .A(n1276), .Z(n24) );
  NAND2_X1 U1390 ( .A1(n1266), .A2(n1286), .ZN(n1276) );
  BUF_X4 U1391 ( .A(a[17]), .Z(n49) );
  BUF_X4 U1392 ( .A(a[9]), .Z(n25) );
  BUF_X4 U1393 ( .A(a[3]), .Z(n7) );
  OAI22_X1 U1394 ( .A1(n1428), .A2(n1094), .B1(n1383), .B2(n1093), .ZN(n478)
         );
  BUF_X4 U1395 ( .A(a[15]), .Z(n43) );
  NAND2_X1 U1396 ( .A1(n1267), .A2(n1287), .ZN(n1277) );
  CLKBUF_X3 U1397 ( .A(b[5]), .Z(n1254) );
  CLKBUF_X1 U1398 ( .A(n65), .Z(n1502) );
  BUF_X4 U1399 ( .A(a[5]), .Z(n13) );
  BUF_X4 U1400 ( .A(a[13]), .Z(n37) );
  BUF_X2 U1401 ( .A(n291), .Z(n63) );
  BUF_X2 U1402 ( .A(n1276), .Z(n23) );
  XNOR2_X1 U1403 ( .A(n209), .B(n1504), .ZN(product[31]) );
  AND2_X1 U1404 ( .A1(n1403), .A2(n208), .ZN(n1504) );
  XNOR2_X1 U1405 ( .A(n231), .B(n1505), .ZN(product[29]) );
  AND2_X1 U1406 ( .A1(n227), .A2(n230), .ZN(n1505) );
  CLKBUF_X3 U1407 ( .A(b[9]), .Z(n1250) );
  NOR2_X1 U1408 ( .A1(n533), .A2(n546), .ZN(n275) );
  NOR2_X1 U1409 ( .A1(n461), .A2(n466), .ZN(n179) );
  NOR2_X1 U1410 ( .A1(n489), .A2(n498), .ZN(n229) );
  NOR2_X1 U1411 ( .A1(n741), .A2(n750), .ZN(n364) );
  NOR2_X1 U1412 ( .A1(n481), .A2(n488), .ZN(n220) );
  NOR2_X1 U1413 ( .A1(n499), .A2(n508), .ZN(n242) );
  NOR2_X1 U1414 ( .A1(n773), .A2(n778), .ZN(n386) );
  AND2_X1 U1415 ( .A1(n1417), .A2(n409), .ZN(product[1]) );
  BUF_X1 U1416 ( .A(n1280), .Z(n58) );
  BUF_X1 U1417 ( .A(n1270), .Z(n60) );
  BUF_X1 U1418 ( .A(n1283), .Z(n39) );
  NAND2_X1 U1419 ( .A1(n1262), .A2(n1282), .ZN(n1272) );
  NAND2_X1 U1420 ( .A1(n1264), .A2(n1284), .ZN(n1274) );
  INV_X1 U1421 ( .A(n1388), .ZN(n1289) );
  NOR2_X1 U1422 ( .A1(n280), .A2(n271), .ZN(n269) );
  NOR2_X1 U1423 ( .A1(n280), .A2(n260), .ZN(n258) );
  NOR2_X1 U1424 ( .A1(n247), .A2(n117), .ZN(n115) );
  NOR2_X1 U1425 ( .A1(n247), .A2(n130), .ZN(n128) );
  NOR2_X1 U1426 ( .A1(n247), .A2(n145), .ZN(n143) );
  NOR2_X1 U1427 ( .A1(n247), .A2(n201), .ZN(n199) );
  NOR2_X1 U1428 ( .A1(n247), .A2(n242), .ZN(n232) );
  NOR2_X1 U1429 ( .A1(n247), .A2(n171), .ZN(n169) );
  NOR2_X1 U1430 ( .A1(n247), .A2(n184), .ZN(n182) );
  NOR2_X1 U1431 ( .A1(n247), .A2(n216), .ZN(n210) );
  NAND2_X1 U1432 ( .A1(n214), .A2(n134), .ZN(n130) );
  INV_X1 U1433 ( .A(n186), .ZN(n184) );
  INV_X1 U1434 ( .A(n173), .ZN(n171) );
  INV_X1 U1435 ( .A(n1426), .ZN(n306) );
  INV_X1 U1436 ( .A(n280), .ZN(n278) );
  INV_X1 U1437 ( .A(n247), .ZN(n245) );
  INV_X1 U1438 ( .A(n1470), .ZN(n319) );
  INV_X1 U1439 ( .A(n282), .ZN(n280) );
  NOR2_X1 U1440 ( .A1(n216), .A2(n175), .ZN(n173) );
  NOR2_X1 U1441 ( .A1(n216), .A2(n192), .ZN(n186) );
  INV_X1 U1442 ( .A(n187), .ZN(n185) );
  INV_X1 U1443 ( .A(n1444), .ZN(n339) );
  NAND2_X1 U1444 ( .A1(n1503), .A2(n1407), .ZN(n326) );
  NOR2_X1 U1445 ( .A1(n1426), .A2(n301), .ZN(n299) );
  INV_X1 U1446 ( .A(n283), .ZN(n281) );
  INV_X1 U1447 ( .A(n216), .ZN(n214) );
  NAND2_X1 U1448 ( .A1(n1492), .A2(n1477), .ZN(n251) );
  NAND2_X1 U1449 ( .A1(n273), .A2(n262), .ZN(n260) );
  OAI21_X1 U1450 ( .B1(n281), .B2(n271), .A(n276), .ZN(n270) );
  OAI21_X1 U1451 ( .B1(n281), .B2(n260), .A(n261), .ZN(n259) );
  AOI21_X1 U1452 ( .B1(n274), .B2(n262), .A(n265), .ZN(n261) );
  INV_X1 U1453 ( .A(n1458), .ZN(n309) );
  INV_X1 U1454 ( .A(n273), .ZN(n271) );
  NOR2_X1 U1455 ( .A1(n247), .A2(n225), .ZN(n223) );
  NOR2_X1 U1456 ( .A1(n247), .A2(n160), .ZN(n158) );
  INV_X1 U1457 ( .A(n192), .ZN(n190) );
  INV_X1 U1458 ( .A(n263), .ZN(n262) );
  INV_X1 U1459 ( .A(n1492), .ZN(n263) );
  NAND2_X1 U1460 ( .A1(n214), .A2(n1403), .ZN(n201) );
  NAND2_X1 U1461 ( .A1(n186), .A2(n149), .ZN(n145) );
  INV_X1 U1462 ( .A(n119), .ZN(n117) );
  INV_X1 U1463 ( .A(n1407), .ZN(n333) );
  INV_X1 U1464 ( .A(n1425), .ZN(n334) );
  INV_X1 U1465 ( .A(n1446), .ZN(n246) );
  XOR2_X1 U1466 ( .A(n339), .B(n89), .Z(product[16]) );
  NAND2_X1 U1467 ( .A1(n1407), .A2(n334), .ZN(n89) );
  XOR2_X1 U1468 ( .A(n347), .B(n90), .Z(product[15]) );
  NAND2_X1 U1469 ( .A1(n1409), .A2(n346), .ZN(n90) );
  AOI21_X1 U1470 ( .B1(n357), .B2(n348), .A(n349), .ZN(n347) );
  XNOR2_X1 U1471 ( .A(n319), .B(n86), .ZN(product[19]) );
  NAND2_X1 U1472 ( .A1(n315), .A2(n318), .ZN(n86) );
  XNOR2_X1 U1473 ( .A(n325), .B(n87), .ZN(product[18]) );
  NAND2_X1 U1474 ( .A1(n430), .A2(n324), .ZN(n87) );
  INV_X1 U1475 ( .A(n1460), .ZN(n430) );
  XNOR2_X1 U1476 ( .A(n332), .B(n88), .ZN(product[17]) );
  NAND2_X1 U1477 ( .A1(n1431), .A2(n331), .ZN(n88) );
  OAI21_X1 U1478 ( .B1(n339), .B2(n333), .A(n334), .ZN(n332) );
  OAI21_X1 U1479 ( .B1(n1486), .B2(n318), .A(n313), .ZN(n311) );
  NOR2_X1 U1480 ( .A1(n312), .A2(n317), .ZN(n310) );
  NAND2_X1 U1481 ( .A1(n425), .A2(n290), .ZN(n82) );
  INV_X1 U1482 ( .A(n289), .ZN(n425) );
  XOR2_X1 U1483 ( .A(n314), .B(n85), .Z(product[20]) );
  NAND2_X1 U1484 ( .A1(n428), .A2(n1432), .ZN(n85) );
  AOI21_X1 U1485 ( .B1(n319), .B2(n315), .A(n316), .ZN(n314) );
  NAND2_X1 U1486 ( .A1(n294), .A2(n310), .ZN(n292) );
  AOI21_X1 U1487 ( .B1(n311), .B2(n1386), .A(n295), .ZN(n293) );
  NOR2_X1 U1488 ( .A1(n296), .A2(n303), .ZN(n294) );
  OAI21_X1 U1489 ( .B1(n341), .B2(n358), .A(n342), .ZN(n340) );
  NAND2_X1 U1490 ( .A1(n348), .A2(n1409), .ZN(n341) );
  AOI21_X1 U1491 ( .B1(n349), .B2(n1409), .A(n344), .ZN(n342) );
  AOI21_X1 U1492 ( .B1(n299), .B2(n319), .A(n300), .ZN(n298) );
  AOI21_X1 U1493 ( .B1(n319), .B2(n306), .A(n1458), .ZN(n305) );
  AOI21_X1 U1494 ( .B1(n340), .B2(n321), .A(n322), .ZN(n320) );
  NOR2_X1 U1495 ( .A1(n1460), .A2(n326), .ZN(n321) );
  OAI21_X1 U1496 ( .B1(n284), .B2(n290), .A(n285), .ZN(n283) );
  INV_X1 U1497 ( .A(n284), .ZN(n424) );
  INV_X1 U1498 ( .A(n358), .ZN(n357) );
  AOI21_X1 U1499 ( .B1(n1503), .B2(n1425), .A(n1456), .ZN(n327) );
  NOR2_X1 U1500 ( .A1(n192), .A2(n136), .ZN(n134) );
  NOR2_X1 U1501 ( .A1(n216), .A2(n121), .ZN(n119) );
  NAND2_X1 U1502 ( .A1(n218), .A2(n240), .ZN(n216) );
  AOI21_X1 U1503 ( .B1(n215), .B2(n1403), .A(n206), .ZN(n202) );
  INV_X1 U1504 ( .A(n174), .ZN(n172) );
  XOR2_X1 U1505 ( .A(n352), .B(n91), .Z(product[14]) );
  NAND2_X1 U1506 ( .A1(n1416), .A2(n351), .ZN(n91) );
  AOI21_X1 U1507 ( .B1(n357), .B2(n435), .A(n354), .ZN(n352) );
  OAI21_X1 U1508 ( .B1(n217), .B2(n192), .A(n193), .ZN(n187) );
  OAI21_X1 U1509 ( .B1(n251), .B2(n276), .A(n252), .ZN(n250) );
  AOI21_X1 U1510 ( .B1(n1477), .B2(n265), .A(n254), .ZN(n252) );
  OAI21_X1 U1511 ( .B1(n1487), .B2(n304), .A(n297), .ZN(n295) );
  OAI21_X1 U1512 ( .B1(n309), .B2(n301), .A(n1445), .ZN(n300) );
  INV_X1 U1513 ( .A(n367), .ZN(n366) );
  INV_X1 U1514 ( .A(n217), .ZN(n215) );
  INV_X1 U1515 ( .A(n275), .ZN(n273) );
  NAND2_X1 U1516 ( .A1(n190), .A2(n177), .ZN(n175) );
  NAND2_X1 U1517 ( .A1(n1403), .A2(n1405), .ZN(n192) );
  INV_X1 U1518 ( .A(n276), .ZN(n274) );
  INV_X1 U1519 ( .A(n267), .ZN(n265) );
  INV_X1 U1520 ( .A(n317), .ZN(n315) );
  NAND2_X1 U1521 ( .A1(n240), .A2(n227), .ZN(n225) );
  INV_X1 U1522 ( .A(n1440), .ZN(n301) );
  INV_X1 U1523 ( .A(n193), .ZN(n191) );
  NAND2_X1 U1524 ( .A1(n173), .A2(n1412), .ZN(n160) );
  INV_X1 U1525 ( .A(n380), .ZN(n379) );
  INV_X1 U1526 ( .A(n318), .ZN(n316) );
  INV_X1 U1527 ( .A(n346), .ZN(n344) );
  INV_X1 U1528 ( .A(n256), .ZN(n254) );
  INV_X1 U1529 ( .A(n290), .ZN(n288) );
  XOR2_X1 U1530 ( .A(n374), .B(n95), .Z(product[10]) );
  NAND2_X1 U1531 ( .A1(n1495), .A2(n373), .ZN(n95) );
  AOI21_X1 U1532 ( .B1(n379), .B2(n1410), .A(n376), .ZN(n374) );
  AOI21_X1 U1533 ( .B1(n218), .B2(n241), .A(n219), .ZN(n217) );
  OAI21_X1 U1534 ( .B1(n230), .B2(n220), .A(n221), .ZN(n219) );
  XNOR2_X1 U1535 ( .A(n385), .B(n97), .ZN(product[8]) );
  XNOR2_X1 U1536 ( .A(n363), .B(n93), .ZN(product[12]) );
  NAND2_X1 U1537 ( .A1(n436), .A2(n362), .ZN(n93) );
  OAI21_X1 U1538 ( .B1(n366), .B2(n364), .A(n365), .ZN(n363) );
  INV_X1 U1539 ( .A(n361), .ZN(n436) );
  XNOR2_X1 U1540 ( .A(n357), .B(n92), .ZN(product[13]) );
  NAND2_X1 U1541 ( .A1(n435), .A2(n356), .ZN(n92) );
  XNOR2_X1 U1542 ( .A(n379), .B(n96), .ZN(product[9]) );
  NAND2_X1 U1543 ( .A1(n1410), .A2(n378), .ZN(n96) );
  OAI21_X1 U1544 ( .B1(n1479), .B2(n356), .A(n351), .ZN(n349) );
  NOR2_X1 U1545 ( .A1(n350), .A2(n355), .ZN(n348) );
  AOI21_X1 U1546 ( .B1(n367), .B2(n359), .A(n360), .ZN(n358) );
  AOI21_X1 U1547 ( .B1(n385), .B2(n1413), .A(n382), .ZN(n380) );
  INV_X1 U1548 ( .A(n384), .ZN(n382) );
  AOI21_X1 U1549 ( .B1(n1405), .B2(n206), .A(n195), .ZN(n193) );
  INV_X1 U1550 ( .A(n197), .ZN(n195) );
  XOR2_X1 U1551 ( .A(n181), .B(n72), .Z(product[33]) );
  NAND2_X1 U1552 ( .A1(n177), .A2(n180), .ZN(n72) );
  OAI21_X1 U1553 ( .B1(n217), .B2(n175), .A(n176), .ZN(n174) );
  AOI21_X1 U1554 ( .B1(n191), .B2(n177), .A(n178), .ZN(n176) );
  INV_X1 U1555 ( .A(n180), .ZN(n178) );
  NAND2_X1 U1556 ( .A1(n629), .A2(n646), .ZN(n318) );
  NOR2_X1 U1557 ( .A1(n629), .A2(n646), .ZN(n317) );
  INV_X1 U1558 ( .A(n220), .ZN(n418) );
  XOR2_X1 U1559 ( .A(n198), .B(n73), .Z(product[32]) );
  NAND2_X1 U1560 ( .A1(n1405), .A2(n197), .ZN(n73) );
  NOR2_X1 U1561 ( .A1(n561), .A2(n576), .ZN(n289) );
  NOR2_X1 U1562 ( .A1(n229), .A2(n220), .ZN(n218) );
  NOR2_X1 U1563 ( .A1(n179), .A2(n151), .ZN(n149) );
  NAND2_X1 U1564 ( .A1(n521), .A2(n532), .ZN(n267) );
  NAND2_X1 U1565 ( .A1(n693), .A2(n706), .ZN(n346) );
  AOI21_X1 U1566 ( .B1(n187), .B2(n149), .A(n150), .ZN(n146) );
  AOI21_X1 U1567 ( .B1(n174), .B2(n1412), .A(n165), .ZN(n161) );
  AOI21_X1 U1568 ( .B1(n215), .B2(n134), .A(n135), .ZN(n131) );
  INV_X1 U1569 ( .A(n120), .ZN(n118) );
  AOI21_X1 U1570 ( .B1(n241), .B2(n227), .A(n228), .ZN(n226) );
  INV_X1 U1571 ( .A(n230), .ZN(n228) );
  NAND2_X1 U1572 ( .A1(n561), .A2(n576), .ZN(n290) );
  NAND2_X1 U1573 ( .A1(n533), .A2(n546), .ZN(n276) );
  NAND2_X1 U1574 ( .A1(n593), .A2(n610), .ZN(n304) );
  OAI21_X1 U1575 ( .B1(n368), .B2(n380), .A(n369), .ZN(n367) );
  NAND2_X1 U1576 ( .A1(n1495), .A2(n1410), .ZN(n368) );
  AOI21_X1 U1577 ( .B1(n1495), .B2(n376), .A(n371), .ZN(n369) );
  NAND2_X1 U1578 ( .A1(n547), .A2(n560), .ZN(n285) );
  NAND2_X1 U1579 ( .A1(n577), .A2(n592), .ZN(n297) );
  NAND2_X1 U1580 ( .A1(n509), .A2(n520), .ZN(n256) );
  INV_X1 U1581 ( .A(n179), .ZN(n177) );
  INV_X1 U1582 ( .A(n229), .ZN(n227) );
  NAND2_X1 U1583 ( .A1(n149), .A2(n1408), .ZN(n136) );
  NAND2_X1 U1584 ( .A1(n134), .A2(n1411), .ZN(n121) );
  NAND2_X1 U1585 ( .A1(n1412), .A2(n1404), .ZN(n151) );
  NAND2_X1 U1586 ( .A1(n647), .A2(n662), .ZN(n324) );
  INV_X1 U1587 ( .A(n378), .ZN(n376) );
  NAND2_X1 U1588 ( .A1(n611), .A2(n628), .ZN(n313) );
  INV_X1 U1589 ( .A(n242), .ZN(n240) );
  INV_X1 U1590 ( .A(n243), .ZN(n241) );
  INV_X1 U1591 ( .A(n208), .ZN(n206) );
  NOR2_X1 U1592 ( .A1(n247), .A2(n108), .ZN(n106) );
  NAND2_X1 U1593 ( .A1(n119), .A2(n1406), .ZN(n108) );
  INV_X1 U1594 ( .A(n373), .ZN(n371) );
  XOR2_X1 U1595 ( .A(n366), .B(n94), .Z(product[11]) );
  NAND2_X1 U1596 ( .A1(n437), .A2(n365), .ZN(n94) );
  INV_X1 U1597 ( .A(n364), .ZN(n437) );
  INV_X1 U1598 ( .A(n356), .ZN(n354) );
  NAND2_X1 U1599 ( .A1(n1414), .A2(n392), .ZN(n99) );
  XOR2_X1 U1600 ( .A(n114), .B(n67), .Z(product[38]) );
  NAND2_X1 U1601 ( .A1(n1406), .A2(n113), .ZN(n67) );
  XOR2_X1 U1602 ( .A(n100), .B(n396), .Z(product[5]) );
  NAND2_X1 U1603 ( .A1(n443), .A2(n395), .ZN(n100) );
  INV_X1 U1604 ( .A(n394), .ZN(n443) );
  INV_X1 U1605 ( .A(n392), .ZN(n390) );
  OAI21_X1 U1606 ( .B1(n388), .B2(n386), .A(n387), .ZN(n385) );
  XOR2_X1 U1607 ( .A(n127), .B(n68), .Z(product[37]) );
  NAND2_X1 U1608 ( .A1(n1411), .A2(n126), .ZN(n68) );
  XOR2_X1 U1609 ( .A(n168), .B(n71), .Z(product[34]) );
  NAND2_X1 U1610 ( .A1(n1412), .A2(n167), .ZN(n71) );
  XOR2_X1 U1611 ( .A(n157), .B(n70), .Z(product[35]) );
  NAND2_X1 U1612 ( .A1(n1404), .A2(n156), .ZN(n70) );
  XOR2_X1 U1613 ( .A(n142), .B(n69), .Z(product[36]) );
  NAND2_X1 U1614 ( .A1(n1408), .A2(n141), .ZN(n69) );
  OAI21_X1 U1615 ( .B1(n151), .B2(n180), .A(n152), .ZN(n150) );
  AOI21_X1 U1616 ( .B1(n165), .B2(n1404), .A(n154), .ZN(n152) );
  INV_X1 U1617 ( .A(n156), .ZN(n154) );
  OAI21_X1 U1618 ( .B1(n193), .B2(n136), .A(n137), .ZN(n135) );
  AOI21_X1 U1619 ( .B1(n150), .B2(n1408), .A(n139), .ZN(n137) );
  INV_X1 U1620 ( .A(n141), .ZN(n139) );
  OAI21_X1 U1621 ( .B1(n217), .B2(n121), .A(n122), .ZN(n120) );
  AOI21_X1 U1622 ( .B1(n135), .B2(n1411), .A(n124), .ZN(n122) );
  INV_X1 U1623 ( .A(n126), .ZN(n124) );
  NAND2_X1 U1624 ( .A1(n461), .A2(n466), .ZN(n180) );
  NAND2_X1 U1625 ( .A1(n489), .A2(n498), .ZN(n230) );
  NAND2_X1 U1626 ( .A1(n741), .A2(n750), .ZN(n365) );
  NAND2_X1 U1627 ( .A1(n719), .A2(n730), .ZN(n356) );
  AOI21_X1 U1628 ( .B1(n120), .B2(n1406), .A(n111), .ZN(n109) );
  INV_X1 U1629 ( .A(n113), .ZN(n111) );
  NAND2_X1 U1630 ( .A1(n499), .A2(n508), .ZN(n243) );
  NAND2_X1 U1631 ( .A1(n473), .A2(n480), .ZN(n208) );
  NAND2_X1 U1632 ( .A1(n467), .A2(n472), .ZN(n197) );
  NAND2_X1 U1633 ( .A1(n481), .A2(n488), .ZN(n221) );
  INV_X1 U1634 ( .A(n167), .ZN(n165) );
  NAND2_X1 U1635 ( .A1(n441), .A2(n387), .ZN(n98) );
  INV_X1 U1636 ( .A(n386), .ZN(n441) );
  NOR2_X1 U1637 ( .A1(n1028), .A2(n1009), .ZN(n406) );
  XOR2_X1 U1638 ( .A(n102), .B(n404), .Z(product[3]) );
  NAND2_X1 U1639 ( .A1(n445), .A2(n403), .ZN(n102) );
  INV_X1 U1640 ( .A(n402), .ZN(n445) );
  XOR2_X1 U1641 ( .A(n103), .B(n409), .Z(product[2]) );
  NAND2_X1 U1642 ( .A1(n446), .A2(n407), .ZN(n103) );
  INV_X1 U1643 ( .A(n406), .ZN(n446) );
  XNOR2_X1 U1644 ( .A(n101), .B(n401), .ZN(product[4]) );
  NAND2_X1 U1645 ( .A1(n1415), .A2(n400), .ZN(n101) );
  OAI21_X1 U1646 ( .B1(n402), .B2(n404), .A(n403), .ZN(n401) );
  NAND2_X1 U1647 ( .A1(n1028), .A2(n1009), .ZN(n407) );
  AOI21_X1 U1648 ( .B1(n1415), .B2(n401), .A(n398), .ZN(n396) );
  INV_X1 U1649 ( .A(n400), .ZN(n398) );
  NAND2_X1 U1650 ( .A1(n830), .A2(n448), .ZN(n113) );
  INV_X1 U1651 ( .A(n448), .ZN(n449) );
  NOR2_X1 U1652 ( .A1(n783), .A2(n786), .ZN(n394) );
  INV_X1 U1653 ( .A(n478), .ZN(n479) );
  INV_X1 U1654 ( .A(n544), .ZN(n545) );
  OR2_X1 U1655 ( .A1(n937), .A2(n865), .ZN(n626) );
  XNOR2_X1 U1656 ( .A(n937), .B(n865), .ZN(n627) );
  NAND2_X1 U1657 ( .A1(n457), .A2(n460), .ZN(n167) );
  NAND2_X1 U1658 ( .A1(n453), .A2(n456), .ZN(n156) );
  NAND2_X1 U1659 ( .A1(n452), .A2(n451), .ZN(n141) );
  NAND2_X1 U1660 ( .A1(n779), .A2(n782), .ZN(n392) );
  NAND2_X1 U1661 ( .A1(n450), .A2(n449), .ZN(n126) );
  NAND2_X1 U1662 ( .A1(n773), .A2(n778), .ZN(n387) );
  NAND2_X1 U1663 ( .A1(n783), .A2(n786), .ZN(n395) );
  INV_X1 U1664 ( .A(n405), .ZN(n404) );
  OAI21_X1 U1665 ( .B1(n406), .B2(n409), .A(n407), .ZN(n405) );
  OAI22_X1 U1666 ( .A1(n54), .A2(n1052), .B1(n52), .B2(n1051), .ZN(n454) );
  OAI22_X1 U1667 ( .A1(n24), .A2(n1157), .B1(n22), .B2(n1156), .ZN(n544) );
  OAI22_X1 U1668 ( .A1(n1463), .A2(n1178), .B1(n16), .B2(n1177), .ZN(n574) );
  OAI22_X1 U1669 ( .A1(n30), .A2(n1136), .B1(n28), .B2(n1135), .ZN(n518) );
  OAI22_X1 U1670 ( .A1(n12), .A2(n1199), .B1(n1198), .B2(n10), .ZN(n608) );
  OAI22_X1 U1671 ( .A1(n48), .A2(n1073), .B1(n46), .B2(n1072), .ZN(n464) );
  OAI22_X1 U1672 ( .A1(n1442), .A2(n1115), .B1(n34), .B2(n1114), .ZN(n496) );
  OAI22_X1 U1673 ( .A1(n53), .A2(n1461), .B1(n51), .B2(n1066), .ZN(n865) );
  OAI22_X1 U1674 ( .A1(n30), .A2(n1143), .B1(n28), .B2(n1142), .ZN(n937) );
  OAI22_X1 U1675 ( .A1(n53), .A2(n1065), .B1(n52), .B2(n1064), .ZN(n863) );
  OAI22_X1 U1676 ( .A1(n23), .A2(n1160), .B1(n22), .B2(n1159), .ZN(n953) );
  OAI22_X1 U1677 ( .A1(n30), .A2(n1139), .B1(n28), .B2(n1138), .ZN(n933) );
  OAI22_X1 U1678 ( .A1(n53), .A2(n1063), .B1(n52), .B2(n1062), .ZN(n861) );
  OAI22_X1 U1679 ( .A1(n23), .A2(n1158), .B1(n22), .B2(n1157), .ZN(n951) );
  OAI22_X1 U1680 ( .A1(n30), .A2(n1147), .B1(n27), .B2(n1146), .ZN(n941) );
  OAI22_X1 U1681 ( .A1(n24), .A2(n1166), .B1(n21), .B2(n1165), .ZN(n959) );
  OAI22_X1 U1682 ( .A1(n1462), .A2(n1185), .B1(n16), .B2(n1184), .ZN(n977) );
  OAI22_X1 U1683 ( .A1(n29), .A2(n1153), .B1(n27), .B2(n1152), .ZN(n947) );
  OAI22_X1 U1684 ( .A1(n11), .A2(n1210), .B1(n9), .B2(n1209), .ZN(n1001) );
  OAI22_X1 U1685 ( .A1(n1463), .A2(n1191), .B1(n15), .B2(n1190), .ZN(n983) );
  OAI22_X1 U1686 ( .A1(n29), .A2(n1148), .B1(n27), .B2(n1147), .ZN(n942) );
  OAI22_X1 U1687 ( .A1(n1448), .A2(n1224), .B1(n4), .B2(n1223), .ZN(n1015) );
  OAI22_X1 U1688 ( .A1(n1462), .A2(n1186), .B1(n16), .B2(n1185), .ZN(n978) );
  OAI22_X1 U1689 ( .A1(n23), .A2(n1175), .B1(n21), .B2(n1174), .ZN(n968) );
  OAI22_X1 U1690 ( .A1(n23), .A2(n1296), .B1(n1176), .B2(n22), .ZN(n826) );
  XNOR2_X1 U1691 ( .A(n1509), .B(n1511), .ZN(n1175) );
  OAI22_X1 U1692 ( .A1(n60), .A2(n1032), .B1(n58), .B2(n1031), .ZN(n831) );
  INV_X1 U1693 ( .A(n793), .ZN(n850) );
  AOI21_X1 U1694 ( .B1(n54), .B2(n52), .A(n1051), .ZN(n793) );
  OAI22_X1 U1695 ( .A1(n1430), .A2(n1034), .B1(n58), .B2(n1033), .ZN(n833) );
  OAI22_X1 U1696 ( .A1(n1430), .A2(n1033), .B1(n58), .B2(n1032), .ZN(n832) );
  INV_X1 U1697 ( .A(n454), .ZN(n455) );
  OAI22_X1 U1698 ( .A1(n11), .A2(n1215), .B1(n9), .B2(n1214), .ZN(n1006) );
  OAI22_X1 U1699 ( .A1(n1448), .A2(n1234), .B1(n1233), .B2(n3), .ZN(n1025) );
  OAI22_X1 U1700 ( .A1(n11), .A2(n1216), .B1(n9), .B2(n1215), .ZN(n1007) );
  AND2_X1 U1701 ( .A1(n1506), .A2(n812), .ZN(n989) );
  OAI22_X1 U1702 ( .A1(n1448), .A2(n1235), .B1(n1234), .B2(n3), .ZN(n1026) );
  OAI22_X1 U1703 ( .A1(n30), .A2(n1295), .B1(n1155), .B2(n28), .ZN(n825) );
  OAI22_X1 U1704 ( .A1(n29), .A2(n1154), .B1(n27), .B2(n1153), .ZN(n948) );
  OR2_X1 U1705 ( .A1(n1507), .A2(n1295), .ZN(n1155) );
  OAI22_X1 U1706 ( .A1(n30), .A2(n1142), .B1(n28), .B2(n1141), .ZN(n936) );
  INV_X1 U1707 ( .A(n608), .ZN(n609) );
  OAI22_X1 U1708 ( .A1(n36), .A2(n1451), .B1(n34), .B2(n1122), .ZN(n918) );
  OAI22_X1 U1709 ( .A1(n60), .A2(n1039), .B1(n58), .B2(n1038), .ZN(n838) );
  OAI22_X1 U1710 ( .A1(n1428), .A2(n1096), .B1(n1383), .B2(n1095), .ZN(n892)
         );
  OAI22_X1 U1711 ( .A1(n54), .A2(n1058), .B1(n52), .B2(n1057), .ZN(n856) );
  AND2_X1 U1712 ( .A1(n1507), .A2(n800), .ZN(n909) );
  OAI22_X1 U1713 ( .A1(n29), .A2(n1151), .B1(n27), .B2(n1150), .ZN(n945) );
  OAI22_X1 U1714 ( .A1(n1449), .A2(n1227), .B1(n1226), .B2(n4), .ZN(n1018) );
  OAI22_X1 U1715 ( .A1(n1430), .A2(n1037), .B1(n58), .B2(n1036), .ZN(n836) );
  OAI22_X1 U1716 ( .A1(n54), .A2(n1056), .B1(n52), .B2(n1055), .ZN(n854) );
  OAI22_X1 U1717 ( .A1(n1387), .A2(n1075), .B1(n46), .B2(n1074), .ZN(n872) );
  OAI22_X1 U1718 ( .A1(n41), .A2(n1105), .B1(n1473), .B2(n1104), .ZN(n901) );
  OAI22_X1 U1719 ( .A1(n12), .A2(n1200), .B1(n10), .B2(n1199), .ZN(n991) );
  OAI22_X1 U1720 ( .A1(n47), .A2(n1452), .B1(n45), .B2(n1085), .ZN(n883) );
  AOI21_X1 U1721 ( .B1(n6), .B2(n4), .A(n1219), .ZN(n817) );
  AOI21_X1 U1722 ( .B1(n1428), .B2(n1383), .A(n1093), .ZN(n799) );
  INV_X1 U1723 ( .A(n790), .ZN(n830) );
  AOI21_X1 U1724 ( .B1(n60), .B2(n58), .A(n1030), .ZN(n790) );
  AOI21_X1 U1725 ( .B1(n1442), .B2(n34), .A(n1114), .ZN(n802) );
  AOI21_X1 U1726 ( .B1(n12), .B2(n10), .A(n1198), .ZN(n814) );
  OAI22_X1 U1727 ( .A1(n1462), .A2(n1195), .B1(n15), .B2(n1194), .ZN(n987) );
  OAI22_X1 U1728 ( .A1(n18), .A2(n1297), .B1(n1197), .B2(n16), .ZN(n827) );
  OAI22_X1 U1729 ( .A1(n1462), .A2(n1196), .B1(n15), .B2(n1195), .ZN(n988) );
  OR2_X1 U1730 ( .A1(n1507), .A2(n1297), .ZN(n1197) );
  OAI22_X1 U1731 ( .A1(n53), .A2(n1070), .B1(n51), .B2(n1069), .ZN(n868) );
  NAND2_X1 U1732 ( .A1(n1029), .A2(n829), .ZN(n409) );
  OAI22_X1 U1733 ( .A1(n30), .A2(n1137), .B1(n27), .B2(n1136), .ZN(n931) );
  OAI22_X1 U1734 ( .A1(n53), .A2(n1061), .B1(n51), .B2(n1060), .ZN(n859) );
  OAI22_X1 U1735 ( .A1(n1442), .A2(n1118), .B1(n34), .B2(n1117), .ZN(n913) );
  OAI22_X1 U1736 ( .A1(n30), .A2(n1138), .B1(n28), .B2(n1137), .ZN(n932) );
  OAI22_X1 U1737 ( .A1(n42), .A2(n1100), .B1(n40), .B2(n1099), .ZN(n896) );
  OAI22_X1 U1738 ( .A1(n1442), .A2(n1119), .B1(n34), .B2(n1118), .ZN(n914) );
  OAI22_X1 U1739 ( .A1(n12), .A2(n1204), .B1(n1203), .B2(n10), .ZN(n995) );
  OAI22_X1 U1740 ( .A1(n35), .A2(n1128), .B1(n33), .B2(n1127), .ZN(n923) );
  OAI22_X1 U1741 ( .A1(n47), .A2(n1090), .B1(n1089), .B2(n45), .ZN(n887) );
  OAI22_X1 U1742 ( .A1(n29), .A2(n1146), .B1(n27), .B2(n1145), .ZN(n940) );
  OAI22_X1 U1743 ( .A1(n12), .A2(n1203), .B1(n10), .B2(n1202), .ZN(n994) );
  OAI22_X1 U1744 ( .A1(n1448), .A2(n1222), .B1(n1420), .B2(n4), .ZN(n1013) );
  OAI22_X1 U1745 ( .A1(n1428), .A2(n1099), .B1(n1383), .B2(n1098), .ZN(n895)
         );
  OAI22_X1 U1746 ( .A1(n1387), .A2(n1080), .B1(n46), .B2(n1079), .ZN(n877) );
  OAI22_X1 U1747 ( .A1(n54), .A2(n1057), .B1(n52), .B2(n1056), .ZN(n855) );
  OAI22_X1 U1748 ( .A1(n1387), .A2(n1076), .B1(n46), .B2(n1075), .ZN(n873) );
  OAI22_X1 U1749 ( .A1(n12), .A2(n1201), .B1(n10), .B2(n1200), .ZN(n992) );
  OAI22_X1 U1750 ( .A1(n1463), .A2(n1182), .B1(n16), .B2(n1181), .ZN(n974) );
  OAI22_X1 U1751 ( .A1(n1442), .A2(n1125), .B1(n33), .B2(n1443), .ZN(n920) );
  OAI22_X1 U1752 ( .A1(n41), .A2(n1108), .B1(n1472), .B2(n1107), .ZN(n904) );
  OAI22_X1 U1753 ( .A1(n36), .A2(n1127), .B1(n34), .B2(n1126), .ZN(n922) );
  OAI22_X1 U1754 ( .A1(n1387), .A2(n1089), .B1(n1088), .B2(n46), .ZN(n886) );
  OAI22_X1 U1755 ( .A1(n1387), .A2(n1077), .B1(n46), .B2(n1076), .ZN(n874) );
  INV_X1 U1756 ( .A(n496), .ZN(n497) );
  OAI22_X1 U1757 ( .A1(n54), .A2(n1059), .B1(n52), .B2(n1058), .ZN(n857) );
  OAI22_X1 U1758 ( .A1(n48), .A2(n1078), .B1(n46), .B2(n1077), .ZN(n875) );
  OAI22_X1 U1759 ( .A1(n36), .A2(n1116), .B1(n34), .B2(n1115), .ZN(n911) );
  INV_X1 U1760 ( .A(n15), .ZN(n812) );
  INV_X1 U1761 ( .A(n21), .ZN(n809) );
  OAI22_X1 U1762 ( .A1(n59), .A2(n1455), .B1(n57), .B2(n1046), .ZN(n846) );
  OAI22_X1 U1763 ( .A1(n42), .A2(n1104), .B1(n1103), .B2(n1472), .ZN(n900) );
  OAI22_X1 U1764 ( .A1(n1462), .A2(n1180), .B1(n16), .B2(n1179), .ZN(n972) );
  OAI22_X1 U1765 ( .A1(n36), .A2(n1122), .B1(n34), .B2(n1121), .ZN(n917) );
  OAI22_X1 U1766 ( .A1(n1448), .A2(n1230), .B1(n1229), .B2(n3), .ZN(n1021) );
  OAI22_X1 U1767 ( .A1(n23), .A2(n1164), .B1(n22), .B2(n1163), .ZN(n957) );
  OAI22_X1 U1768 ( .A1(n41), .A2(n1103), .B1(n1473), .B2(n1102), .ZN(n899) );
  OAI22_X1 U1769 ( .A1(n29), .A2(n1141), .B1(n28), .B2(n1140), .ZN(n935) );
  OAI22_X1 U1770 ( .A1(n48), .A2(n1084), .B1(n46), .B2(n1083), .ZN(n881) );
  OAI22_X1 U1771 ( .A1(n53), .A2(n1064), .B1(n52), .B2(n1063), .ZN(n862) );
  OAI22_X1 U1772 ( .A1(n60), .A2(n1045), .B1(n57), .B2(n1044), .ZN(n844) );
  OAI22_X1 U1773 ( .A1(n1442), .A2(n1121), .B1(n34), .B2(n1120), .ZN(n916) );
  OAI22_X1 U1774 ( .A1(n11), .A2(n1211), .B1(n9), .B2(n1210), .ZN(n1002) );
  OAI22_X1 U1775 ( .A1(n23), .A2(n1173), .B1(n21), .B2(n1172), .ZN(n966) );
  OAI22_X1 U1776 ( .A1(n1463), .A2(n1192), .B1(n15), .B2(n1191), .ZN(n984) );
  AND2_X1 U1777 ( .A1(n1511), .A2(n791), .ZN(n849) );
  OAI22_X1 U1778 ( .A1(n1221), .A2(n6), .B1(n1220), .B2(n4), .ZN(n1012) );
  OAI22_X1 U1779 ( .A1(n47), .A2(n1088), .B1(n1087), .B2(n45), .ZN(n885) );
  OAI22_X1 U1780 ( .A1(n23), .A2(n1165), .B1(n22), .B2(n1164), .ZN(n958) );
  OAI22_X1 U1781 ( .A1(n1462), .A2(n1184), .B1(n16), .B2(n1183), .ZN(n976) );
  OAI22_X1 U1782 ( .A1(n41), .A2(n1098), .B1(n40), .B2(n1097), .ZN(n894) );
  OAI22_X1 U1783 ( .A1(n36), .A2(n1117), .B1(n34), .B2(n1116), .ZN(n912) );
  OAI22_X1 U1784 ( .A1(n48), .A2(n1079), .B1(n46), .B2(n1078), .ZN(n876) );
  OAI22_X1 U1785 ( .A1(n1457), .A2(n47), .B1(n45), .B2(n1086), .ZN(n884) );
  OAI22_X1 U1786 ( .A1(n42), .A2(n1110), .B1(n1473), .B2(n1109), .ZN(n906) );
  OAI22_X1 U1787 ( .A1(n1129), .A2(n35), .B1(n33), .B2(n1128), .ZN(n924) );
  OAI22_X1 U1788 ( .A1(n23), .A2(n1167), .B1(n1166), .B2(n21), .ZN(n960) );
  OAI22_X1 U1789 ( .A1(n30), .A2(n1150), .B1(n27), .B2(n1149), .ZN(n944) );
  OAI22_X1 U1790 ( .A1(n1463), .A2(n1188), .B1(n15), .B2(n1187), .ZN(n980) );
  OAI22_X1 U1791 ( .A1(n1442), .A2(n1131), .B1(n33), .B2(n1130), .ZN(n926) );
  OAI22_X1 U1792 ( .A1(n1430), .A2(n1044), .B1(n57), .B2(n1043), .ZN(n843) );
  INV_X1 U1793 ( .A(n811), .ZN(n970) );
  AOI21_X1 U1794 ( .B1(n18), .B2(n16), .A(n1177), .ZN(n811) );
  OAI22_X1 U1795 ( .A1(n1048), .A2(n59), .B1(n1047), .B2(n57), .ZN(n847) );
  OAI22_X1 U1796 ( .A1(n35), .A2(n1459), .B1(n1123), .B2(n33), .ZN(n919) );
  INV_X1 U1797 ( .A(n817), .ZN(n1010) );
  OAI22_X1 U1798 ( .A1(n23), .A2(n1168), .B1(n21), .B2(n1167), .ZN(n961) );
  OAI22_X1 U1799 ( .A1(n1462), .A2(n1187), .B1(n15), .B2(n1186), .ZN(n979) );
  OAI22_X1 U1800 ( .A1(n11), .A2(n1212), .B1(n9), .B2(n1211), .ZN(n1003) );
  OAI22_X1 U1801 ( .A1(n23), .A2(n1174), .B1(n21), .B2(n1173), .ZN(n967) );
  OAI22_X1 U1802 ( .A1(n1429), .A2(n1042), .B1(n57), .B2(n1041), .ZN(n841) );
  INV_X1 U1803 ( .A(n808), .ZN(n950) );
  AOI21_X1 U1804 ( .B1(n24), .B2(n22), .A(n1156), .ZN(n808) );
  OAI22_X1 U1805 ( .A1(n11), .A2(n1213), .B1(n9), .B2(n1212), .ZN(n1004) );
  OAI22_X1 U1806 ( .A1(n1449), .A2(n1232), .B1(n1231), .B2(n3), .ZN(n1023) );
  OAI22_X1 U1807 ( .A1(n1462), .A2(n1194), .B1(n15), .B2(n1193), .ZN(n986) );
  OAI22_X1 U1808 ( .A1(n11), .A2(n1214), .B1(n9), .B2(n1213), .ZN(n1005) );
  AND2_X1 U1809 ( .A1(n1507), .A2(n809), .ZN(n969) );
  OAI22_X1 U1810 ( .A1(n1449), .A2(n1233), .B1(n1232), .B2(n3), .ZN(n1024) );
  OAI22_X1 U1811 ( .A1(n1428), .A2(n1102), .B1(n1383), .B2(n1101), .ZN(n898)
         );
  INV_X1 U1812 ( .A(n1469), .ZN(n575) );
  OAI22_X1 U1813 ( .A1(n12), .A2(n1205), .B1(n10), .B2(n1204), .ZN(n996) );
  OAI22_X1 U1814 ( .A1(n42), .A2(n1101), .B1(n40), .B2(n1100), .ZN(n897) );
  OAI22_X1 U1815 ( .A1(n1387), .A2(n1082), .B1(n46), .B2(n1081), .ZN(n879) );
  OAI22_X1 U1816 ( .A1(n1442), .A2(n1120), .B1(n34), .B2(n1119), .ZN(n915) );
  AND2_X1 U1817 ( .A1(n1506), .A2(n803), .ZN(n929) );
  OAI22_X1 U1818 ( .A1(n1448), .A2(n1229), .B1(n1228), .B2(n3), .ZN(n1020) );
  OAI22_X1 U1819 ( .A1(n24), .A2(n1172), .B1(n21), .B2(n1171), .ZN(n965) );
  OAI22_X1 U1820 ( .A1(n30), .A2(n1145), .B1(n27), .B2(n1144), .ZN(n939) );
  OAI22_X1 U1821 ( .A1(n18), .A2(n1183), .B1(n16), .B2(n1182), .ZN(n975) );
  OAI22_X1 U1822 ( .A1(n35), .A2(n1126), .B1(n33), .B2(n1125), .ZN(n921) );
  AND2_X1 U1823 ( .A1(n1506), .A2(n797), .ZN(n889) );
  OAI22_X1 U1824 ( .A1(n1448), .A2(n1225), .B1(n1224), .B2(n4), .ZN(n1016) );
  OAI22_X1 U1825 ( .A1(n35), .A2(n1130), .B1(n33), .B2(n1129), .ZN(n925) );
  OAI22_X1 U1826 ( .A1(n30), .A2(n1140), .B1(n28), .B2(n1139), .ZN(n934) );
  OAI22_X1 U1827 ( .A1(n23), .A2(n1159), .B1(n22), .B2(n1158), .ZN(n952) );
  OAI22_X1 U1828 ( .A1(n1387), .A2(n1083), .B1(n46), .B2(n1082), .ZN(n880) );
  OAI22_X1 U1829 ( .A1(n42), .A2(n1109), .B1(n1108), .B2(n1472), .ZN(n905) );
  AND2_X1 U1830 ( .A1(n1506), .A2(n794), .ZN(n869) );
  OAI22_X1 U1831 ( .A1(n6), .A2(n1392), .B1(n1222), .B2(n4), .ZN(n1014) );
  OAI22_X1 U1832 ( .A1(n12), .A2(n1207), .B1(n10), .B2(n1206), .ZN(n998) );
  OAI22_X1 U1833 ( .A1(n1448), .A2(n1226), .B1(n1225), .B2(n4), .ZN(n1017) );
  OAI22_X1 U1834 ( .A1(n24), .A2(n1169), .B1(n21), .B2(n1168), .ZN(n962) );
  OAI22_X1 U1835 ( .A1(n29), .A2(n1149), .B1(n27), .B2(n1148), .ZN(n943) );
  OAI22_X1 U1836 ( .A1(n41), .A2(n1111), .B1(n1473), .B2(n1110), .ZN(n907) );
  OAI22_X1 U1837 ( .A1(n12), .A2(n1206), .B1(n10), .B2(n1205), .ZN(n997) );
  OAI22_X1 U1838 ( .A1(n23), .A2(n1162), .B1(n22), .B2(n1161), .ZN(n955) );
  OAI22_X1 U1839 ( .A1(n1463), .A2(n1181), .B1(n16), .B2(n1180), .ZN(n973) );
  INV_X1 U1840 ( .A(n1510), .ZN(n1296) );
  OAI22_X1 U1841 ( .A1(n48), .A2(n1074), .B1(n46), .B2(n1073), .ZN(n871) );
  OAI22_X1 U1842 ( .A1(n11), .A2(n1208), .B1(n9), .B2(n1207), .ZN(n999) );
  OAI22_X1 U1843 ( .A1(n23), .A2(n1170), .B1(n21), .B2(n1169), .ZN(n963) );
  OAI22_X1 U1844 ( .A1(n1442), .A2(n1132), .B1(n33), .B2(n1131), .ZN(n927) );
  OAI22_X1 U1845 ( .A1(n1428), .A2(n1097), .B1(n1383), .B2(n1096), .ZN(n893)
         );
  OAI22_X1 U1846 ( .A1(n11), .A2(n1209), .B1(n9), .B2(n1208), .ZN(n1000) );
  OAI22_X1 U1847 ( .A1(n23), .A2(n1171), .B1(n21), .B2(n1170), .ZN(n964) );
  OAI22_X1 U1848 ( .A1(n1462), .A2(n1189), .B1(n15), .B2(n1188), .ZN(n981) );
  OAI22_X1 U1849 ( .A1(n1046), .A2(n1430), .B1(n1045), .B2(n57), .ZN(n845) );
  INV_X1 U1850 ( .A(n814), .ZN(n990) );
  OAI22_X1 U1851 ( .A1(n1179), .A2(n18), .B1(n1178), .B2(n16), .ZN(n971) );
  OAI22_X1 U1852 ( .A1(n53), .A2(n1062), .B1(n52), .B2(n1061), .ZN(n860) );
  OAI22_X1 U1853 ( .A1(n1430), .A2(n1043), .B1(n57), .B2(n1042), .ZN(n842) );
  OAI22_X1 U1854 ( .A1(n1387), .A2(n1081), .B1(n46), .B2(n1080), .ZN(n878) );
  OAI22_X1 U1855 ( .A1(n41), .A2(n1106), .B1(n1472), .B2(n1105), .ZN(n902) );
  OAI22_X1 U1856 ( .A1(n1449), .A2(n1423), .B1(n1422), .B2(n4), .ZN(n1011) );
  OAI22_X1 U1857 ( .A1(n24), .A2(n1163), .B1(n22), .B2(n1162), .ZN(n956) );
  OAI22_X1 U1858 ( .A1(n53), .A2(n1066), .B1(n51), .B2(n1065), .ZN(n864) );
  OAI22_X1 U1859 ( .A1(n48), .A2(n1085), .B1(n46), .B2(n1084), .ZN(n882) );
  OAI22_X1 U1860 ( .A1(n24), .A2(n1161), .B1(n22), .B2(n1160), .ZN(n954) );
  AND2_X1 U1861 ( .A1(n1511), .A2(n806), .ZN(n949) );
  OAI22_X1 U1862 ( .A1(n1448), .A2(n1231), .B1(n1230), .B2(n3), .ZN(n1022) );
  OAI22_X1 U1863 ( .A1(n1462), .A2(n1193), .B1(n15), .B2(n1192), .ZN(n985) );
  OAI22_X1 U1864 ( .A1(n41), .A2(n1107), .B1(n1472), .B2(n1106), .ZN(n903) );
  OAI22_X1 U1865 ( .A1(n53), .A2(n1069), .B1(n51), .B2(n1454), .ZN(n867) );
  OAI22_X1 U1866 ( .A1(n12), .A2(n1202), .B1(n10), .B2(n1201), .ZN(n993) );
  OAI22_X1 U1867 ( .A1(n29), .A2(n1152), .B1(n27), .B2(n1151), .ZN(n946) );
  OAI22_X1 U1868 ( .A1(n1449), .A2(n1228), .B1(n1227), .B2(n4), .ZN(n1019) );
  OAI22_X1 U1869 ( .A1(n18), .A2(n1190), .B1(n15), .B2(n1189), .ZN(n982) );
  NAND2_X1 U1870 ( .A1(n787), .A2(n788), .ZN(n400) );
  OAI22_X1 U1871 ( .A1(n48), .A2(n1292), .B1(n1092), .B2(n45), .ZN(n822) );
  OAI22_X1 U1872 ( .A1(n1387), .A2(n1091), .B1(n46), .B2(n1090), .ZN(n888) );
  OR2_X1 U1873 ( .A1(n1506), .A2(n1292), .ZN(n1092) );
  OAI22_X1 U1874 ( .A1(n1429), .A2(n1290), .B1(n1050), .B2(n58), .ZN(n820) );
  OAI22_X1 U1875 ( .A1(n60), .A2(n1049), .B1(n57), .B2(n1453), .ZN(n848) );
  OR2_X1 U1876 ( .A1(n1506), .A2(n1290), .ZN(n1050) );
  OAI22_X1 U1877 ( .A1(n41), .A2(n1293), .B1(n1113), .B2(n40), .ZN(n823) );
  OAI22_X1 U1878 ( .A1(n41), .A2(n1112), .B1(n1472), .B2(n1111), .ZN(n908) );
  OR2_X1 U1879 ( .A1(n1506), .A2(n1293), .ZN(n1113) );
  OAI22_X1 U1880 ( .A1(n1429), .A2(n1041), .B1(n57), .B2(n1040), .ZN(n840) );
  OAI22_X1 U1881 ( .A1(n54), .A2(n1060), .B1(n52), .B2(n1059), .ZN(n858) );
  INV_X1 U1882 ( .A(n518), .ZN(n519) );
  OAI22_X1 U1883 ( .A1(n60), .A2(n1035), .B1(n58), .B2(n1034), .ZN(n834) );
  OAI22_X1 U1884 ( .A1(n54), .A2(n1054), .B1(n52), .B2(n1053), .ZN(n852) );
  INV_X1 U1885 ( .A(n464), .ZN(n465) );
  INV_X1 U1886 ( .A(n27), .ZN(n806) );
  OR2_X1 U1887 ( .A1(n1507), .A2(n1296), .ZN(n1176) );
  OR2_X1 U1888 ( .A1(n1507), .A2(n1294), .ZN(n1134) );
  OAI22_X1 U1889 ( .A1(n1429), .A2(n1040), .B1(n57), .B2(n1039), .ZN(n839) );
  INV_X1 U1890 ( .A(n805), .ZN(n930) );
  AOI21_X1 U1891 ( .B1(n30), .B2(n28), .A(n1135), .ZN(n805) );
  OAI22_X1 U1892 ( .A1(n54), .A2(n1053), .B1(n52), .B2(n1052), .ZN(n851) );
  INV_X1 U1893 ( .A(n796), .ZN(n870) );
  AOI21_X1 U1894 ( .B1(n1387), .B2(n46), .A(n1072), .ZN(n796) );
  OAI22_X1 U1895 ( .A1(n54), .A2(n1055), .B1(n52), .B2(n1054), .ZN(n853) );
  OAI22_X1 U1896 ( .A1(n1429), .A2(n1036), .B1(n58), .B2(n1035), .ZN(n835) );
  INV_X1 U1897 ( .A(n799), .ZN(n890) );
  OAI22_X1 U1898 ( .A1(n41), .A2(n1095), .B1(n1383), .B2(n1094), .ZN(n891) );
  OAI22_X1 U1899 ( .A1(n1430), .A2(n1038), .B1(n58), .B2(n1037), .ZN(n837) );
  INV_X1 U1900 ( .A(n802), .ZN(n910) );
  INV_X1 U1901 ( .A(n57), .ZN(n791) );
  INV_X1 U1902 ( .A(n1471), .ZN(n800) );
  AND2_X1 U1903 ( .A1(n1506), .A2(n815), .ZN(n1009) );
  INV_X1 U1904 ( .A(n9), .ZN(n815) );
  INV_X1 U1905 ( .A(n33), .ZN(n803) );
  INV_X1 U1906 ( .A(n45), .ZN(n797) );
  INV_X1 U1907 ( .A(n51), .ZN(n794) );
  AND2_X1 U1908 ( .A1(n1511), .A2(n818), .ZN(product[0]) );
  INV_X1 U1909 ( .A(n3), .ZN(n818) );
  OR2_X1 U1910 ( .A1(n1507), .A2(n1298), .ZN(n1218) );
  INV_X1 U1911 ( .A(n7), .ZN(n1298) );
  OAI22_X1 U1912 ( .A1(n11), .A2(n1217), .B1(n9), .B2(n1216), .ZN(n1008) );
  OAI22_X1 U1913 ( .A1(n1448), .A2(n1236), .B1(n1235), .B2(n3), .ZN(n1027) );
  XNOR2_X1 U1914 ( .A(n7), .B(n1506), .ZN(n1217) );
  XNOR2_X1 U1915 ( .A(n1510), .B(n1253), .ZN(n1169) );
  XNOR2_X1 U1916 ( .A(n1509), .B(n1254), .ZN(n1170) );
  XNOR2_X1 U1917 ( .A(n1510), .B(n1248), .ZN(n1164) );
  OAI22_X1 U1918 ( .A1(n1448), .A2(n1299), .B1(n1239), .B2(n4), .ZN(n829) );
  OR2_X1 U1919 ( .A1(n1507), .A2(n1299), .ZN(n1239) );
  INV_X1 U1920 ( .A(n1424), .ZN(n1299) );
  OAI22_X1 U1921 ( .A1(n1449), .A2(n1238), .B1(n1237), .B2(n3), .ZN(n1029) );
  XNOR2_X1 U1922 ( .A(n1510), .B(n1255), .ZN(n1171) );
  XNOR2_X1 U1923 ( .A(n1510), .B(n1256), .ZN(n1172) );
  XNOR2_X1 U1924 ( .A(n1510), .B(n1244), .ZN(n1160) );
  XNOR2_X1 U1925 ( .A(n1510), .B(n1245), .ZN(n1161) );
  XNOR2_X1 U1926 ( .A(n7), .B(n1393), .ZN(n1215) );
  XNOR2_X1 U1927 ( .A(n7), .B(n1258), .ZN(n1216) );
  XNOR2_X1 U1928 ( .A(n7), .B(n1255), .ZN(n1213) );
  XNOR2_X1 U1929 ( .A(n7), .B(n1256), .ZN(n1214) );
  XNOR2_X1 U1930 ( .A(n7), .B(n1252), .ZN(n1210) );
  XNOR2_X1 U1931 ( .A(n7), .B(n1253), .ZN(n1211) );
  XNOR2_X1 U1932 ( .A(n31), .B(n1254), .ZN(n1128) );
  XNOR2_X1 U1933 ( .A(n1465), .B(n1249), .ZN(n1123) );
  XNOR2_X1 U1934 ( .A(n31), .B(n1255), .ZN(n1129) );
  XNOR2_X1 U1935 ( .A(n31), .B(n1245), .ZN(n1119) );
  XNOR2_X1 U1936 ( .A(n31), .B(n1246), .ZN(n1120) );
  XNOR2_X1 U1937 ( .A(n31), .B(n1243), .ZN(n1117) );
  XNOR2_X1 U1938 ( .A(n1465), .B(n1242), .ZN(n1116) );
  XNOR2_X1 U1939 ( .A(n1465), .B(n1244), .ZN(n1118) );
  XNOR2_X1 U1940 ( .A(n7), .B(n1241), .ZN(n1199) );
  XNOR2_X1 U1941 ( .A(n7), .B(n1242), .ZN(n1200) );
  XNOR2_X1 U1942 ( .A(n31), .B(n1247), .ZN(n1121) );
  XNOR2_X1 U1943 ( .A(n31), .B(n1251), .ZN(n1125) );
  XNOR2_X1 U1944 ( .A(n31), .B(n1252), .ZN(n1126) );
  XNOR2_X1 U1945 ( .A(n7), .B(n1243), .ZN(n1201) );
  XNOR2_X1 U1946 ( .A(n7), .B(n1244), .ZN(n1202) );
  XNOR2_X1 U1947 ( .A(n31), .B(n1256), .ZN(n1130) );
  XNOR2_X1 U1948 ( .A(n7), .B(n1245), .ZN(n1203) );
  XNOR2_X1 U1949 ( .A(n7), .B(n1246), .ZN(n1204) );
  XNOR2_X1 U1950 ( .A(n1499), .B(n1241), .ZN(n1115) );
  XNOR2_X1 U1951 ( .A(n1465), .B(n1257), .ZN(n1131) );
  XNOR2_X1 U1952 ( .A(n31), .B(n1253), .ZN(n1127) );
  XNOR2_X1 U1953 ( .A(n7), .B(n1249), .ZN(n1207) );
  XNOR2_X1 U1954 ( .A(n7), .B(n1250), .ZN(n1208) );
  XNOR2_X1 U1955 ( .A(n1465), .B(n1258), .ZN(n1132) );
  XNOR2_X1 U1956 ( .A(n1499), .B(n1248), .ZN(n1122) );
  XNOR2_X1 U1957 ( .A(n7), .B(n1247), .ZN(n1205) );
  XNOR2_X1 U1958 ( .A(n7), .B(n1248), .ZN(n1206) );
  XNOR2_X1 U1959 ( .A(n7), .B(n1254), .ZN(n1212) );
  XNOR2_X1 U1960 ( .A(n7), .B(n1389), .ZN(n1209) );
  XNOR2_X1 U1961 ( .A(n1510), .B(n1257), .ZN(n1173) );
  XNOR2_X1 U1962 ( .A(n1250), .B(n1510), .ZN(n1166) );
  XNOR2_X1 U1963 ( .A(n1510), .B(n1251), .ZN(n1167) );
  XNOR2_X1 U1964 ( .A(n1510), .B(n1241), .ZN(n1157) );
  XNOR2_X1 U1965 ( .A(n1509), .B(n1246), .ZN(n1162) );
  XNOR2_X1 U1966 ( .A(n1510), .B(n1247), .ZN(n1163) );
  XNOR2_X1 U1967 ( .A(n1510), .B(n1242), .ZN(n1158) );
  XNOR2_X1 U1968 ( .A(n1509), .B(n1243), .ZN(n1159) );
  XNOR2_X1 U1969 ( .A(n1510), .B(n1249), .ZN(n1165) );
  XNOR2_X1 U1970 ( .A(n1509), .B(n1252), .ZN(n1168) );
  XNOR2_X1 U1971 ( .A(n1509), .B(n1500), .ZN(n1174) );
  XNOR2_X1 U1972 ( .A(n7), .B(n1240), .ZN(n1198) );
  XNOR2_X1 U1973 ( .A(n1465), .B(n1421), .ZN(n1114) );
  XNOR2_X1 U1974 ( .A(n1510), .B(n1240), .ZN(n1156) );
  BUF_X1 U1975 ( .A(n1288), .Z(n10) );
  BUF_X1 U1976 ( .A(n1271), .Z(n54) );
  BUF_X1 U1977 ( .A(n1278), .Z(n11) );
  OAI22_X1 U1978 ( .A1(n1442), .A2(n1133), .B1(n33), .B2(n1132), .ZN(n928) );
  OAI22_X1 U1979 ( .A1(n36), .A2(n1294), .B1(n1134), .B2(n34), .ZN(n824) );
  XNOR2_X1 U1980 ( .A(n31), .B(n1507), .ZN(n1133) );
  INV_X1 U1981 ( .A(n31), .ZN(n1294) );
  BUF_X1 U1982 ( .A(n1289), .Z(n3) );
  BUF_X1 U1983 ( .A(n1289), .Z(n4) );
  INV_X1 U1984 ( .A(n25), .ZN(n1295) );
  INV_X1 U1985 ( .A(n43), .ZN(n1292) );
  INV_X1 U1986 ( .A(n37), .ZN(n1293) );
  INV_X1 U1987 ( .A(n13), .ZN(n1297) );
  INV_X1 U1988 ( .A(n55), .ZN(n1290) );
  XNOR2_X1 U1989 ( .A(a[10]), .B(a[9]), .ZN(n1284) );
  XNOR2_X1 U1990 ( .A(a[14]), .B(a[13]), .ZN(n1282) );
  XNOR2_X1 U1991 ( .A(a[1]), .B(a[2]), .ZN(n1288) );
  XNOR2_X1 U1992 ( .A(a[16]), .B(a[15]), .ZN(n1281) );
  NAND2_X1 U1993 ( .A1(n1269), .A2(n1289), .ZN(n1279) );
  NAND2_X1 U1994 ( .A1(n1268), .A2(n1288), .ZN(n1278) );
  NAND2_X1 U1995 ( .A1(n1265), .A2(n1285), .ZN(n1275) );
  XNOR2_X1 U1996 ( .A(n1468), .B(n1247), .ZN(n1058) );
  INV_X1 U1997 ( .A(n49), .ZN(n1291) );
  XNOR2_X1 U1998 ( .A(n49), .B(n1506), .ZN(n1070) );
  XNOR2_X1 U1999 ( .A(n49), .B(n1390), .ZN(n1057) );
  XNOR2_X1 U2000 ( .A(n49), .B(n1258), .ZN(n1069) );
  XNOR2_X1 U2001 ( .A(n49), .B(n1253), .ZN(n1064) );
  XNOR2_X1 U2002 ( .A(n1468), .B(n1243), .ZN(n1054) );
  XNOR2_X1 U2003 ( .A(n49), .B(n1252), .ZN(n1063) );
  XNOR2_X1 U2004 ( .A(n49), .B(n1248), .ZN(n1059) );
  XNOR2_X1 U2005 ( .A(n1468), .B(n1242), .ZN(n1053) );
  XNOR2_X1 U2006 ( .A(n49), .B(n1251), .ZN(n1062) );
  XNOR2_X1 U2007 ( .A(n49), .B(n1257), .ZN(n1068) );
  XNOR2_X1 U2008 ( .A(n49), .B(n1245), .ZN(n1056) );
  XNOR2_X1 U2009 ( .A(n1468), .B(n1244), .ZN(n1055) );
  XNOR2_X1 U2010 ( .A(n1250), .B(n49), .ZN(n1061) );
  XNOR2_X1 U2011 ( .A(n49), .B(n1249), .ZN(n1060) );
  XNOR2_X1 U2012 ( .A(n49), .B(n1255), .ZN(n1066) );
  XNOR2_X1 U2013 ( .A(n49), .B(n1254), .ZN(n1065) );
  XNOR2_X1 U2014 ( .A(n1468), .B(n1241), .ZN(n1052) );
  XNOR2_X1 U2015 ( .A(n1468), .B(n1485), .ZN(n1051) );
  INV_X1 U2016 ( .A(n355), .ZN(n435) );
  NOR2_X1 U2017 ( .A1(n719), .A2(n730), .ZN(n355) );
  CLKBUF_X1 U2018 ( .A(a[7]), .Z(n1509) );
  CLKBUF_X1 U2019 ( .A(n1287), .Z(n15) );
  INV_X1 U2020 ( .A(n1439), .ZN(n428) );
  OAI22_X1 U2021 ( .A1(n1448), .A2(n1237), .B1(n1236), .B2(n3), .ZN(n1028) );
  XNOR2_X1 U2022 ( .A(n1450), .B(n1485), .ZN(n1030) );
  XNOR2_X1 U2023 ( .A(n1450), .B(n1241), .ZN(n1031) );
  XNOR2_X1 U2024 ( .A(n1450), .B(n1243), .ZN(n1033) );
  XNOR2_X1 U2025 ( .A(n1450), .B(n1242), .ZN(n1032) );
  XNOR2_X1 U2026 ( .A(n1450), .B(n1249), .ZN(n1039) );
  XNOR2_X1 U2027 ( .A(n1450), .B(n1511), .ZN(n1049) );
  XNOR2_X1 U2028 ( .A(n1450), .B(n1245), .ZN(n1035) );
  XNOR2_X1 U2029 ( .A(n1450), .B(n1248), .ZN(n1038) );
  XNOR2_X1 U2030 ( .A(n1450), .B(n1244), .ZN(n1034) );
  XNOR2_X1 U2031 ( .A(n1250), .B(n1450), .ZN(n1040) );
  XNOR2_X1 U2032 ( .A(n55), .B(n1254), .ZN(n1044) );
  XNOR2_X1 U2033 ( .A(n55), .B(n1253), .ZN(n1043) );
  XNOR2_X1 U2034 ( .A(n1450), .B(n1247), .ZN(n1037) );
  XNOR2_X1 U2035 ( .A(n1450), .B(n1252), .ZN(n1042) );
  XNOR2_X1 U2036 ( .A(n1450), .B(n1390), .ZN(n1036) );
  XNOR2_X1 U2037 ( .A(n55), .B(n1258), .ZN(n1048) );
  XNOR2_X1 U2038 ( .A(n1450), .B(n1251), .ZN(n1041) );
  XNOR2_X1 U2039 ( .A(n55), .B(n1255), .ZN(n1045) );
  XNOR2_X1 U2040 ( .A(n1257), .B(n55), .ZN(n1047) );
  XNOR2_X1 U2041 ( .A(n1256), .B(n55), .ZN(n1046) );
  XNOR2_X1 U2042 ( .A(n1467), .B(n1245), .ZN(n1077) );
  XNOR2_X1 U2043 ( .A(n43), .B(n1507), .ZN(n1091) );
  XNOR2_X1 U2044 ( .A(n1467), .B(n1244), .ZN(n1076) );
  XNOR2_X1 U2045 ( .A(n43), .B(n1254), .ZN(n1086) );
  XNOR2_X1 U2046 ( .A(n1467), .B(n1243), .ZN(n1075) );
  XNOR2_X1 U2047 ( .A(n43), .B(n1251), .ZN(n1083) );
  XNOR2_X1 U2048 ( .A(n1467), .B(n1242), .ZN(n1074) );
  XNOR2_X1 U2049 ( .A(n43), .B(n1258), .ZN(n1090) );
  XNOR2_X1 U2050 ( .A(n43), .B(n1257), .ZN(n1089) );
  XNOR2_X1 U2051 ( .A(n43), .B(n1247), .ZN(n1079) );
  XNOR2_X1 U2052 ( .A(n1250), .B(n43), .ZN(n1082) );
  XNOR2_X1 U2053 ( .A(n43), .B(n1246), .ZN(n1078) );
  XNOR2_X1 U2054 ( .A(n43), .B(n1256), .ZN(n1088) );
  XNOR2_X1 U2055 ( .A(n43), .B(n1249), .ZN(n1081) );
  XNOR2_X1 U2056 ( .A(n43), .B(n1248), .ZN(n1080) );
  XNOR2_X1 U2057 ( .A(n43), .B(n1255), .ZN(n1087) );
  XNOR2_X1 U2058 ( .A(n1467), .B(n1241), .ZN(n1073) );
  XNOR2_X1 U2059 ( .A(n43), .B(n1253), .ZN(n1085) );
  XNOR2_X1 U2060 ( .A(n43), .B(n1252), .ZN(n1084) );
  XNOR2_X1 U2061 ( .A(n1467), .B(n1485), .ZN(n1072) );
  XOR2_X1 U2062 ( .A(n388), .B(n98), .Z(product[7]) );
  AOI21_X1 U2063 ( .B1(n1414), .B2(n393), .A(n390), .ZN(n388) );
  XNOR2_X1 U2064 ( .A(n13), .B(n1494), .ZN(n1194) );
  XNOR2_X1 U2065 ( .A(n13), .B(n1244), .ZN(n1181) );
  XNOR2_X1 U2066 ( .A(n13), .B(n1253), .ZN(n1190) );
  XNOR2_X1 U2067 ( .A(n13), .B(n1252), .ZN(n1189) );
  XNOR2_X1 U2068 ( .A(n13), .B(n1256), .ZN(n1193) );
  XNOR2_X1 U2069 ( .A(n13), .B(n1251), .ZN(n1188) );
  XNOR2_X1 U2070 ( .A(n13), .B(n1506), .ZN(n1196) );
  XNOR2_X1 U2071 ( .A(n13), .B(n1258), .ZN(n1195) );
  XNOR2_X1 U2072 ( .A(n1250), .B(n13), .ZN(n1187) );
  XNOR2_X1 U2073 ( .A(n13), .B(n1247), .ZN(n1184) );
  XNOR2_X1 U2074 ( .A(n13), .B(n1249), .ZN(n1186) );
  XNOR2_X1 U2075 ( .A(n13), .B(n1246), .ZN(n1183) );
  XNOR2_X1 U2076 ( .A(n13), .B(n1248), .ZN(n1185) );
  XNOR2_X1 U2077 ( .A(n13), .B(n1255), .ZN(n1192) );
  XNOR2_X1 U2078 ( .A(n13), .B(n1254), .ZN(n1191) );
  XNOR2_X1 U2079 ( .A(n13), .B(n1245), .ZN(n1182) );
  XNOR2_X1 U2080 ( .A(n13), .B(n1243), .ZN(n1180) );
  XNOR2_X1 U2081 ( .A(n13), .B(n1242), .ZN(n1179) );
  XNOR2_X1 U2082 ( .A(n13), .B(n1241), .ZN(n1178) );
  XNOR2_X1 U2083 ( .A(n13), .B(n1240), .ZN(n1177) );
  XNOR2_X1 U2084 ( .A(n37), .B(n1243), .ZN(n1096) );
  XNOR2_X1 U2085 ( .A(n37), .B(n1249), .ZN(n1102) );
  XNOR2_X1 U2086 ( .A(n37), .B(n1253), .ZN(n1106) );
  XNOR2_X1 U2087 ( .A(n37), .B(n1242), .ZN(n1095) );
  XNOR2_X1 U2088 ( .A(n37), .B(n1252), .ZN(n1105) );
  XNOR2_X1 U2089 ( .A(n37), .B(n1245), .ZN(n1098) );
  XNOR2_X1 U2090 ( .A(n37), .B(n1244), .ZN(n1097) );
  XNOR2_X1 U2091 ( .A(n37), .B(n1248), .ZN(n1101) );
  XNOR2_X1 U2092 ( .A(n37), .B(n1254), .ZN(n1107) );
  XNOR2_X1 U2093 ( .A(n37), .B(n1247), .ZN(n1100) );
  XNOR2_X1 U2094 ( .A(n37), .B(n1257), .ZN(n1110) );
  XNOR2_X1 U2095 ( .A(n37), .B(n1256), .ZN(n1109) );
  XNOR2_X1 U2096 ( .A(n37), .B(n1255), .ZN(n1108) );
  XNOR2_X1 U2097 ( .A(n37), .B(n1246), .ZN(n1099) );
  XNOR2_X1 U2098 ( .A(n37), .B(n1511), .ZN(n1112) );
  XNOR2_X1 U2099 ( .A(n37), .B(n1258), .ZN(n1111) );
  XNOR2_X1 U2100 ( .A(n37), .B(n1251), .ZN(n1104) );
  XNOR2_X1 U2101 ( .A(n37), .B(n1250), .ZN(n1103) );
  XNOR2_X1 U2102 ( .A(n37), .B(n1241), .ZN(n1094) );
  XNOR2_X1 U2103 ( .A(n37), .B(n1485), .ZN(n1093) );
  NAND2_X1 U2104 ( .A1(n751), .A2(n758), .ZN(n373) );
  XNOR2_X1 U2105 ( .A(n25), .B(n1246), .ZN(n1141) );
  XNOR2_X1 U2106 ( .A(n25), .B(n1245), .ZN(n1140) );
  XNOR2_X1 U2107 ( .A(n25), .B(n1255), .ZN(n1150) );
  XNOR2_X1 U2108 ( .A(n25), .B(n1244), .ZN(n1139) );
  XNOR2_X1 U2109 ( .A(n25), .B(n1254), .ZN(n1149) );
  XNOR2_X1 U2110 ( .A(n25), .B(n1511), .ZN(n1154) );
  XNOR2_X1 U2111 ( .A(n25), .B(n1257), .ZN(n1152) );
  XNOR2_X1 U2112 ( .A(n25), .B(n1256), .ZN(n1151) );
  XNOR2_X1 U2113 ( .A(n25), .B(n1247), .ZN(n1142) );
  XNOR2_X1 U2114 ( .A(n25), .B(n1248), .ZN(n1143) );
  XNOR2_X1 U2115 ( .A(n25), .B(n1250), .ZN(n1145) );
  XNOR2_X1 U2116 ( .A(n25), .B(n1258), .ZN(n1153) );
  XNOR2_X1 U2117 ( .A(n25), .B(n1243), .ZN(n1138) );
  XNOR2_X1 U2118 ( .A(n25), .B(n1253), .ZN(n1148) );
  XNOR2_X1 U2119 ( .A(n25), .B(n1249), .ZN(n1144) );
  XNOR2_X1 U2120 ( .A(n25), .B(n1242), .ZN(n1137) );
  XNOR2_X1 U2121 ( .A(n25), .B(n1252), .ZN(n1147) );
  XNOR2_X1 U2122 ( .A(n25), .B(n1251), .ZN(n1146) );
  XNOR2_X1 U2123 ( .A(n25), .B(n1241), .ZN(n1136) );
  XNOR2_X1 U2124 ( .A(n25), .B(n1240), .ZN(n1135) );
  OAI21_X1 U2125 ( .B1(n339), .B2(n326), .A(n1491), .ZN(n325) );
  OAI21_X1 U2126 ( .B1(n327), .B2(n323), .A(n324), .ZN(n322) );
  XNOR2_X1 U2127 ( .A(a[18]), .B(a[17]), .ZN(n1280) );
  OAI22_X1 U2128 ( .A1(n54), .A2(n1291), .B1(n1071), .B2(n51), .ZN(n821) );
  OR2_X1 U2129 ( .A1(n1511), .A2(n1291), .ZN(n1071) );
  OAI21_X1 U2130 ( .B1(n1502), .B2(n108), .A(n109), .ZN(n107) );
  OAI21_X1 U2131 ( .B1(n1502), .B2(n117), .A(n118), .ZN(n116) );
  OAI21_X1 U2132 ( .B1(n1446), .B2(n160), .A(n161), .ZN(n159) );
  OAI21_X1 U2133 ( .B1(n145), .B2(n65), .A(n146), .ZN(n144) );
  OAI21_X1 U2134 ( .B1(n248), .B2(n242), .A(n243), .ZN(n233) );
  OAI21_X1 U2135 ( .B1(n1446), .B2(n184), .A(n185), .ZN(n183) );
  OAI21_X1 U2136 ( .B1(n65), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U2137 ( .B1(n65), .B2(n171), .A(n172), .ZN(n170) );
  OAI21_X1 U2138 ( .B1(n1446), .B2(n201), .A(n202), .ZN(n200) );
  OAI21_X1 U2139 ( .B1(n248), .B2(n216), .A(n217), .ZN(n211) );
  OAI21_X1 U2140 ( .B1(n1446), .B2(n225), .A(n226), .ZN(n224) );
  OAI21_X1 U2141 ( .B1(n394), .B2(n396), .A(n395), .ZN(n393) );
  XNOR2_X1 U2142 ( .A(n99), .B(n393), .ZN(product[6]) );
  XNOR2_X1 U2143 ( .A(n1424), .B(n1248), .ZN(n1227) );
  XNOR2_X1 U2144 ( .A(n1), .B(n1389), .ZN(n1230) );
  XNOR2_X1 U2145 ( .A(n1424), .B(n1247), .ZN(n1226) );
  XNOR2_X1 U2146 ( .A(n1), .B(n1252), .ZN(n1231) );
  XNOR2_X1 U2147 ( .A(n1424), .B(n1246), .ZN(n1225) );
  XNOR2_X1 U2148 ( .A(n1), .B(n1245), .ZN(n1224) );
  XNOR2_X1 U2149 ( .A(n1424), .B(n1244), .ZN(n1223) );
  XNOR2_X1 U2150 ( .A(n1424), .B(n1242), .ZN(n1221) );
  XNOR2_X1 U2151 ( .A(n1), .B(n1243), .ZN(n1222) );
  XNOR2_X1 U2152 ( .A(n1), .B(n1241), .ZN(n1220) );
  XNOR2_X1 U2153 ( .A(n1250), .B(n1424), .ZN(n1229) );
  XNOR2_X1 U2154 ( .A(n1424), .B(n1249), .ZN(n1228) );
  XNOR2_X1 U2155 ( .A(n1424), .B(n1253), .ZN(n1232) );
  XNOR2_X1 U2156 ( .A(n1), .B(n1511), .ZN(n1238) );
  XNOR2_X1 U2157 ( .A(n1424), .B(n1254), .ZN(n1233) );
  XNOR2_X1 U2158 ( .A(n1), .B(n1240), .ZN(n1219) );
  XNOR2_X1 U2159 ( .A(n1424), .B(n1256), .ZN(n1235) );
  XNOR2_X1 U2160 ( .A(n1424), .B(n1255), .ZN(n1234) );
  XNOR2_X1 U2161 ( .A(n1424), .B(n1258), .ZN(n1237) );
  XNOR2_X1 U2162 ( .A(n1), .B(n1494), .ZN(n1236) );
  NAND2_X1 U2163 ( .A1(n1413), .A2(n384), .ZN(n97) );
  XNOR2_X1 U2164 ( .A(a[8]), .B(a[7]), .ZN(n1285) );
  XOR2_X1 U2165 ( .A(a[6]), .B(a[7]), .Z(n1266) );
  NAND2_X1 U2166 ( .A1(n767), .A2(n772), .ZN(n384) );
  NOR2_X1 U2167 ( .A1(n361), .A2(n364), .ZN(n359) );
  OAI21_X1 U2168 ( .B1(n361), .B2(n365), .A(n362), .ZN(n360) );
  NAND2_X1 U2169 ( .A1(n731), .A2(n740), .ZN(n362) );
  XNOR2_X1 U2170 ( .A(a[12]), .B(a[11]), .ZN(n1283) );
  XOR2_X1 U2171 ( .A(a[10]), .B(a[11]), .Z(n1264) );
  NAND2_X1 U2172 ( .A1(n1261), .A2(n1281), .ZN(n1271) );
  XOR2_X1 U2173 ( .A(a[18]), .B(a[19]), .Z(n1260) );
  NOR2_X1 U2174 ( .A1(n289), .A2(n284), .ZN(n282) );
  NAND2_X1 U2175 ( .A1(n1260), .A2(n1280), .ZN(n1270) );
  NAND2_X1 U2176 ( .A1(n1263), .A2(n1283), .ZN(n1273) );
  OAI21_X1 U2177 ( .B1(n320), .B2(n292), .A(n293), .ZN(n291) );
  XOR2_X1 U2178 ( .A(a[16]), .B(a[17]), .Z(n1261) );
  XOR2_X1 U2179 ( .A(a[14]), .B(a[15]), .Z(n1262) );
  AOI21_X1 U2180 ( .B1(n1438), .B2(n106), .A(n107), .ZN(n105) );
  AOI21_X1 U2181 ( .B1(n1438), .B2(n115), .A(n116), .ZN(n114) );
  AOI21_X1 U2182 ( .B1(n64), .B2(n182), .A(n183), .ZN(n181) );
  AOI21_X1 U2183 ( .B1(n1438), .B2(n143), .A(n144), .ZN(n142) );
  AOI21_X1 U2184 ( .B1(n1438), .B2(n128), .A(n129), .ZN(n127) );
  AOI21_X1 U2185 ( .B1(n64), .B2(n199), .A(n200), .ZN(n198) );
  AOI21_X1 U2186 ( .B1(n63), .B2(n210), .A(n211), .ZN(n209) );
  AOI21_X1 U2187 ( .B1(n1385), .B2(n169), .A(n170), .ZN(n168) );
  AOI21_X1 U2188 ( .B1(n64), .B2(n158), .A(n159), .ZN(n157) );
  NAND2_X1 U2189 ( .A1(n759), .A2(n766), .ZN(n378) );
  XOR2_X1 U2190 ( .A(a[8]), .B(a[9]), .Z(n1265) );
  NAND2_X1 U2191 ( .A1(n707), .A2(n718), .ZN(n351) );
  XOR2_X1 U2192 ( .A(a[13]), .B(a[12]), .Z(n1263) );
  XOR2_X1 U2193 ( .A(a[2]), .B(a[3]), .Z(n1268) );
  XNOR2_X1 U2194 ( .A(a[4]), .B(a[3]), .ZN(n1287) );
  OAI22_X1 U2195 ( .A1(n12), .A2(n1298), .B1(n1218), .B2(n10), .ZN(n828) );
  NAND2_X1 U2196 ( .A1(n789), .A2(n828), .ZN(n403) );
  AOI21_X1 U2197 ( .B1(n64), .B2(n245), .A(n246), .ZN(n244) );
  AOI21_X1 U2198 ( .B1(n63), .B2(n232), .A(n233), .ZN(n231) );
  AOI21_X1 U2199 ( .B1(n64), .B2(n223), .A(n224), .ZN(n222) );
  XNOR2_X1 U2200 ( .A(n64), .B(n82), .ZN(product[23]) );
  AOI21_X1 U2201 ( .B1(n63), .B2(n425), .A(n288), .ZN(n286) );
  AOI21_X1 U2202 ( .B1(n63), .B2(n269), .A(n270), .ZN(n268) );
  AOI21_X1 U2203 ( .B1(n63), .B2(n278), .A(n1419), .ZN(n277) );
  AOI21_X1 U2204 ( .B1(n63), .B2(n258), .A(n259), .ZN(n257) );
  XOR2_X1 U2205 ( .A(a[4]), .B(a[5]), .Z(n1267) );
  XNOR2_X1 U2206 ( .A(a[6]), .B(a[5]), .ZN(n1286) );
  XOR2_X1 U2207 ( .A(a[1]), .B(a[0]), .Z(n1269) );
endmodule


module datapath_DW_mult_tc_10 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n15, n16, n17, n18,
         n19, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34, n35,
         n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n51, n52,
         n53, n54, n55, n58, n59, n60, n61, n63, n64, n65, n67, n68, n69, n70,
         n71, n72, n73, n82, n83, n84, n85, n86, n87, n88, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n105, n106,
         n107, n108, n109, n111, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n124, n126, n127, n128, n129, n130, n131, n134,
         n135, n136, n137, n139, n141, n142, n143, n144, n145, n146, n149,
         n150, n151, n152, n154, n156, n157, n158, n159, n160, n161, n165,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n190,
         n191, n192, n193, n195, n197, n198, n199, n200, n201, n202, n206,
         n208, n209, n210, n211, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n254, n256, n257, n258, n259, n260, n261,
         n262, n263, n267, n268, n269, n270, n271, n273, n274, n275, n276,
         n277, n278, n280, n281, n282, n283, n284, n285, n286, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n302, n303, n304, n305, n306, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n332, n333, n334, n336, n338, n339, n340, n341, n342,
         n344, n346, n347, n348, n349, n350, n351, n352, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n371, n373, n374, n376, n378, n379, n380, n382, n384,
         n385, n386, n387, n388, n390, n392, n393, n394, n395, n396, n398,
         n400, n401, n402, n403, n404, n405, n406, n407, n409, n418, n424,
         n425, n426, n428, n430, n435, n436, n437, n441, n443, n445, n446,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n793, n794, n796, n797, n799, n800, n802, n803,
         n805, n806, n808, n809, n811, n812, n814, n815, n817, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1493,
         n1494;
  assign product[39] = n105;

  FA_X1 U488 ( .A(n831), .B(n454), .CI(n850), .CO(n450), .S(n451) );
  FA_X1 U489 ( .A(n455), .B(n832), .CI(n458), .CO(n452), .S(n453) );
  FA_X1 U491 ( .A(n462), .B(n833), .CI(n459), .CO(n456), .S(n457) );
  FA_X1 U492 ( .A(n851), .B(n464), .CI(n870), .CO(n458), .S(n459) );
  FA_X1 U493 ( .A(n463), .B(n470), .CI(n468), .CO(n460), .S(n461) );
  FA_X1 U494 ( .A(n834), .B(n852), .CI(n465), .CO(n462), .S(n463) );
  FA_X1 U496 ( .A(n474), .B(n471), .CI(n469), .CO(n466), .S(n467) );
  FA_X1 U497 ( .A(n478), .B(n871), .CI(n476), .CO(n468), .S(n469) );
  FA_X1 U498 ( .A(n853), .B(n835), .CI(n890), .CO(n470), .S(n471) );
  FA_X1 U499 ( .A(n475), .B(n477), .CI(n482), .CO(n472), .S(n473) );
  FA_X1 U500 ( .A(n486), .B(n479), .CI(n484), .CO(n474), .S(n475) );
  FA_X1 U501 ( .A(n836), .B(n854), .CI(n872), .CO(n476), .S(n477) );
  FA_X1 U503 ( .A(n490), .B(n492), .CI(n483), .CO(n480), .S(n481) );
  FA_X1 U504 ( .A(n485), .B(n494), .CI(n487), .CO(n482), .S(n483) );
  FA_X1 U505 ( .A(n855), .B(n496), .CI(n873), .CO(n484), .S(n485) );
  FA_X1 U506 ( .A(n891), .B(n837), .CI(n910), .CO(n486), .S(n487) );
  FA_X1 U507 ( .A(n500), .B(n493), .CI(n491), .CO(n488), .S(n489) );
  FA_X1 U508 ( .A(n495), .B(n504), .CI(n502), .CO(n490), .S(n491) );
  FA_X1 U509 ( .A(n497), .B(n874), .CI(n506), .CO(n492), .S(n493) );
  FA_X1 U510 ( .A(n892), .B(n856), .CI(n838), .CO(n494), .S(n495) );
  FA_X1 U512 ( .A(n510), .B(n503), .CI(n501), .CO(n498), .S(n499) );
  FA_X1 U513 ( .A(n507), .B(n505), .CI(n512), .CO(n500), .S(n501) );
  FA_X1 U514 ( .A(n516), .B(n893), .CI(n514), .CO(n502), .S(n503) );
  FA_X1 U515 ( .A(n857), .B(n911), .CI(n875), .CO(n504), .S(n505) );
  FA_X1 U516 ( .A(n518), .B(n839), .CI(n930), .CO(n506), .S(n507) );
  FA_X1 U517 ( .A(n522), .B(n513), .CI(n511), .CO(n508), .S(n509) );
  FA_X1 U518 ( .A(n526), .B(n515), .CI(n524), .CO(n510), .S(n511) );
  FA_X1 U519 ( .A(n528), .B(n530), .CI(n517), .CO(n512), .S(n513) );
  FA_X1 U520 ( .A(n840), .B(n858), .CI(n519), .CO(n514), .S(n515) );
  FA_X1 U521 ( .A(n912), .B(n876), .CI(n894), .CO(n516), .S(n517) );
  FA_X1 U523 ( .A(n525), .B(n534), .CI(n523), .CO(n520), .S(n521) );
  FA_X1 U524 ( .A(n527), .B(n538), .CI(n536), .CO(n522), .S(n523) );
  FA_X1 U525 ( .A(n529), .B(n540), .CI(n531), .CO(n524), .S(n525) );
  FA_X1 U526 ( .A(n877), .B(n895), .CI(n542), .CO(n526), .S(n527) );
  FA_X1 U527 ( .A(n913), .B(n859), .CI(n931), .CO(n528), .S(n529) );
  FA_X1 U528 ( .A(n544), .B(n841), .CI(n950), .CO(n530), .S(n531) );
  FA_X1 U529 ( .A(n548), .B(n537), .CI(n535), .CO(n532), .S(n533) );
  FA_X1 U530 ( .A(n539), .B(n552), .CI(n550), .CO(n534), .S(n535) );
  FA_X1 U531 ( .A(n541), .B(n554), .CI(n543), .CO(n536), .S(n537) );
  FA_X1 U532 ( .A(n558), .B(n545), .CI(n556), .CO(n538), .S(n539) );
  FA_X1 U533 ( .A(n896), .B(n932), .CI(n914), .CO(n540), .S(n541) );
  FA_X1 U534 ( .A(n842), .B(n878), .CI(n860), .CO(n542), .S(n543) );
  FA_X1 U536 ( .A(n562), .B(n551), .CI(n549), .CO(n546), .S(n547) );
  FA_X1 U537 ( .A(n553), .B(n566), .CI(n564), .CO(n548), .S(n549) );
  FA_X1 U538 ( .A(n559), .B(n557), .CI(n568), .CO(n550), .S(n551) );
  FA_X1 U539 ( .A(n570), .B(n572), .CI(n555), .CO(n552), .S(n553) );
  FA_X1 U540 ( .A(n879), .B(n915), .CI(n897), .CO(n554), .S(n555) );
  FA_X1 U541 ( .A(n861), .B(n951), .CI(n933), .CO(n556), .S(n557) );
  FA_X1 U542 ( .A(n574), .B(n843), .CI(n970), .CO(n558), .S(n559) );
  FA_X1 U543 ( .A(n578), .B(n565), .CI(n563), .CO(n560), .S(n561) );
  FA_X1 U544 ( .A(n567), .B(n582), .CI(n580), .CO(n562), .S(n563) );
  FA_X1 U545 ( .A(n584), .B(n573), .CI(n569), .CO(n564), .S(n565) );
  FA_X1 U546 ( .A(n586), .B(n588), .CI(n571), .CO(n566), .S(n567) );
  FA_X1 U547 ( .A(n575), .B(n898), .CI(n590), .CO(n568), .S(n569) );
  FA_X1 U548 ( .A(n844), .B(n916), .CI(n862), .CO(n570), .S(n571) );
  FA_X1 U549 ( .A(n952), .B(n880), .CI(n934), .CO(n572), .S(n573) );
  FA_X1 U553 ( .A(n600), .B(n591), .CI(n585), .CO(n580), .S(n581) );
  FA_X1 U554 ( .A(n587), .B(n602), .CI(n589), .CO(n582), .S(n583) );
  FA_X1 U555 ( .A(n606), .B(n917), .CI(n604), .CO(n584), .S(n585) );
  FA_X1 U556 ( .A(n881), .B(n935), .CI(n899), .CO(n586), .S(n587) );
  FA_X1 U557 ( .A(n608), .B(n953), .CI(n863), .CO(n588), .S(n589) );
  FA_X1 U558 ( .A(n845), .B(n971), .CI(n990), .CO(n590), .S(n591) );
  FA_X1 U559 ( .A(n612), .B(n597), .CI(n595), .CO(n592), .S(n593) );
  FA_X1 U560 ( .A(n599), .B(n616), .CI(n614), .CO(n594), .S(n595) );
  FA_X1 U561 ( .A(n618), .B(n603), .CI(n601), .CO(n596), .S(n597) );
  FA_X1 U562 ( .A(n605), .B(n620), .CI(n607), .CO(n598), .S(n599) );
  FA_X1 U563 ( .A(n626), .B(n624), .CI(n622), .CO(n600), .S(n601) );
  FA_X1 U564 ( .A(n918), .B(n936), .CI(n609), .CO(n602), .S(n603) );
  FA_X1 U565 ( .A(n882), .B(n864), .CI(n954), .CO(n604), .S(n605) );
  FA_X1 U569 ( .A(n617), .B(n634), .CI(n632), .CO(n612), .S(n613) );
  FA_X1 U570 ( .A(n636), .B(n621), .CI(n619), .CO(n614), .S(n615) );
  FA_X1 U571 ( .A(n623), .B(n638), .CI(n625), .CO(n616), .S(n617) );
  FA_X1 U572 ( .A(n627), .B(n642), .CI(n640), .CO(n618), .S(n619) );
  FA_X1 U573 ( .A(n955), .B(n973), .CI(n644), .CO(n620), .S(n621) );
  FA_X1 U574 ( .A(n991), .B(n901), .CI(n883), .CO(n622), .S(n623) );
  FA_X1 U575 ( .A(n919), .B(n847), .CI(n1010), .CO(n624), .S(n625) );
  FA_X1 U578 ( .A(n648), .B(n633), .CI(n631), .CO(n628), .S(n629) );
  FA_X1 U579 ( .A(n650), .B(n637), .CI(n635), .CO(n630), .S(n631) );
  FA_X1 U580 ( .A(n654), .B(n643), .CI(n652), .CO(n632), .S(n633) );
  FA_X1 U581 ( .A(n639), .B(n656), .CI(n641), .CO(n634), .S(n635) );
  FA_X1 U582 ( .A(n660), .B(n645), .CI(n658), .CO(n636), .S(n637) );
  FA_X1 U583 ( .A(n920), .B(n992), .CI(n974), .CO(n638), .S(n639) );
  FA_X1 U584 ( .A(n902), .B(n956), .CI(n1011), .CO(n640), .S(n641) );
  FA_X1 U585 ( .A(n866), .B(n884), .CI(n938), .CO(n642), .S(n643) );
  HA_X1 U586 ( .A(n820), .B(n848), .CO(n644), .S(n645) );
  FA_X1 U587 ( .A(n664), .B(n651), .CI(n649), .CO(n646), .S(n647) );
  FA_X1 U588 ( .A(n666), .B(n655), .CI(n653), .CO(n648), .S(n649) );
  FA_X1 U589 ( .A(n670), .B(n659), .CI(n668), .CO(n650), .S(n651) );
  FA_X1 U590 ( .A(n661), .B(n672), .CI(n657), .CO(n652), .S(n653) );
  FA_X1 U591 ( .A(n676), .B(n957), .CI(n674), .CO(n654), .S(n655) );
  FA_X1 U592 ( .A(n921), .B(n939), .CI(n975), .CO(n656), .S(n657) );
  FA_X1 U593 ( .A(n867), .B(n993), .CI(n903), .CO(n658), .S(n659) );
  FA_X1 U594 ( .A(n849), .B(n885), .CI(n1012), .CO(n660), .S(n661) );
  FA_X1 U595 ( .A(n667), .B(n680), .CI(n665), .CO(n662), .S(n663) );
  FA_X1 U596 ( .A(n669), .B(n671), .CI(n682), .CO(n664), .S(n665) );
  FA_X1 U598 ( .A(n686), .B(n690), .CI(n688), .CO(n668), .S(n669) );
  FA_X1 U599 ( .A(n958), .B(n976), .CI(n677), .CO(n670), .S(n671) );
  FA_X1 U600 ( .A(n886), .B(n904), .CI(n922), .CO(n672), .S(n673) );
  FA_X1 U601 ( .A(n1013), .B(n940), .CI(n994), .CO(n674), .S(n675) );
  HA_X1 U602 ( .A(n868), .B(n821), .CO(n676), .S(n677) );
  FA_X1 U603 ( .A(n694), .B(n683), .CI(n681), .CO(n678), .S(n679) );
  FA_X1 U604 ( .A(n685), .B(n698), .CI(n696), .CO(n680), .S(n681) );
  FA_X1 U605 ( .A(n689), .B(n691), .CI(n687), .CO(n682), .S(n683) );
  FA_X1 U606 ( .A(n702), .B(n704), .CI(n700), .CO(n684), .S(n685) );
  FA_X1 U607 ( .A(n941), .B(n959), .CI(n977), .CO(n686), .S(n687) );
  FA_X1 U608 ( .A(n887), .B(n923), .CI(n995), .CO(n688), .S(n689) );
  FA_X1 U609 ( .A(n869), .B(n905), .CI(n1014), .CO(n690), .S(n691) );
  FA_X1 U610 ( .A(n697), .B(n708), .CI(n695), .CO(n692), .S(n693) );
  FA_X1 U611 ( .A(n699), .B(n703), .CI(n710), .CO(n694), .S(n695) );
  FA_X1 U612 ( .A(n712), .B(n714), .CI(n701), .CO(n696), .S(n697) );
  FA_X1 U613 ( .A(n705), .B(n996), .CI(n716), .CO(n698), .S(n699) );
  FA_X1 U614 ( .A(n978), .B(n942), .CI(n1015), .CO(n700), .S(n701) );
  HA_X1 U616 ( .A(n822), .B(n888), .CO(n704), .S(n705) );
  FA_X1 U617 ( .A(n711), .B(n720), .CI(n709), .CO(n706), .S(n707) );
  FA_X1 U618 ( .A(n713), .B(n715), .CI(n722), .CO(n708), .S(n709) );
  FA_X1 U619 ( .A(n724), .B(n726), .CI(n717), .CO(n710), .S(n711) );
  FA_X1 U620 ( .A(n961), .B(n979), .CI(n728), .CO(n712), .S(n713) );
  FA_X1 U621 ( .A(n907), .B(n997), .CI(n943), .CO(n714), .S(n715) );
  FA_X1 U622 ( .A(n889), .B(n925), .CI(n1016), .CO(n716), .S(n717) );
  FA_X1 U623 ( .A(n732), .B(n723), .CI(n721), .CO(n718), .S(n719) );
  FA_X1 U624 ( .A(n727), .B(n725), .CI(n734), .CO(n720), .S(n721) );
  FA_X1 U625 ( .A(n738), .B(n729), .CI(n736), .CO(n722), .S(n723) );
  FA_X1 U626 ( .A(n926), .B(n980), .CI(n944), .CO(n724), .S(n725) );
  FA_X1 U627 ( .A(n1017), .B(n962), .CI(n998), .CO(n726), .S(n727) );
  HA_X1 U628 ( .A(n908), .B(n823), .CO(n728), .S(n729) );
  FA_X1 U629 ( .A(n735), .B(n742), .CI(n733), .CO(n730), .S(n731) );
  FA_X1 U630 ( .A(n737), .B(n739), .CI(n744), .CO(n732), .S(n733) );
  FA_X1 U631 ( .A(n748), .B(n981), .CI(n746), .CO(n734), .S(n735) );
  FA_X1 U632 ( .A(n927), .B(n999), .CI(n963), .CO(n736), .S(n737) );
  FA_X1 U633 ( .A(n945), .B(n909), .CI(n1018), .CO(n738), .S(n739) );
  FA_X1 U634 ( .A(n752), .B(n745), .CI(n743), .CO(n740), .S(n741) );
  FA_X1 U635 ( .A(n754), .B(n756), .CI(n747), .CO(n742), .S(n743) );
  FA_X1 U636 ( .A(n964), .B(n1000), .CI(n749), .CO(n744), .S(n745) );
  FA_X1 U637 ( .A(n946), .B(n982), .CI(n1019), .CO(n746), .S(n747) );
  HA_X1 U638 ( .A(n824), .B(n928), .CO(n748), .S(n749) );
  FA_X1 U639 ( .A(n760), .B(n755), .CI(n753), .CO(n750), .S(n751) );
  FA_X1 U640 ( .A(n762), .B(n764), .CI(n757), .CO(n752), .S(n753) );
  FA_X1 U641 ( .A(n947), .B(n1001), .CI(n983), .CO(n754), .S(n755) );
  FA_X1 U642 ( .A(n965), .B(n929), .CI(n1020), .CO(n756), .S(n757) );
  FA_X1 U643 ( .A(n763), .B(n768), .CI(n761), .CO(n758), .S(n759) );
  FA_X1 U644 ( .A(n765), .B(n1021), .CI(n770), .CO(n760), .S(n761) );
  FA_X1 U645 ( .A(n966), .B(n984), .CI(n1002), .CO(n762), .S(n763) );
  HA_X1 U646 ( .A(n825), .B(n948), .CO(n764), .S(n765) );
  FA_X1 U647 ( .A(n771), .B(n774), .CI(n769), .CO(n766), .S(n767) );
  FA_X1 U648 ( .A(n967), .B(n1003), .CI(n776), .CO(n768), .S(n769) );
  FA_X1 U649 ( .A(n1022), .B(n949), .CI(n985), .CO(n770), .S(n771) );
  FA_X1 U650 ( .A(n780), .B(n777), .CI(n775), .CO(n772), .S(n773) );
  FA_X1 U651 ( .A(n986), .B(n1023), .CI(n1004), .CO(n774), .S(n775) );
  HA_X1 U652 ( .A(n826), .B(n968), .CO(n776), .S(n777) );
  FA_X1 U653 ( .A(n784), .B(n987), .CI(n781), .CO(n778), .S(n779) );
  FA_X1 U654 ( .A(n1024), .B(n969), .CI(n1005), .CO(n780), .S(n781) );
  FA_X1 U655 ( .A(n1006), .B(n1025), .CI(n785), .CO(n782), .S(n783) );
  HA_X1 U656 ( .A(n827), .B(n988), .CO(n784), .S(n785) );
  FA_X1 U657 ( .A(n1026), .B(n989), .CI(n1007), .CO(n786), .S(n787) );
  HA_X1 U658 ( .A(n1008), .B(n1027), .CO(n788), .S(n789) );
  NOR2_X2 U1180 ( .A1(n251), .A2(n275), .ZN(n249) );
  CLKBUF_X2 U1181 ( .A(b[11]), .Z(n1248) );
  BUF_X1 U1182 ( .A(n1278), .Z(n1429) );
  AOI21_X1 U1183 ( .B1(n283), .B2(n249), .A(n250), .ZN(n1383) );
  BUF_X2 U1184 ( .A(b[13]), .Z(n1246) );
  BUF_X1 U1185 ( .A(n1), .Z(n1384) );
  BUF_X1 U1186 ( .A(n1146), .Z(n1385) );
  CLKBUF_X3 U1187 ( .A(b[15]), .Z(n1244) );
  CLKBUF_X2 U1188 ( .A(b[14]), .Z(n1245) );
  CLKBUF_X3 U1189 ( .A(b[16]), .Z(n1243) );
  CLKBUF_X3 U1190 ( .A(b[6]), .Z(n1253) );
  CLKBUF_X3 U1191 ( .A(b[2]), .Z(n1257) );
  CLKBUF_X3 U1192 ( .A(b[4]), .Z(n1255) );
  BUF_X2 U1193 ( .A(b[19]), .Z(n1240) );
  OR2_X1 U1194 ( .A1(n787), .A2(n788), .ZN(n1386) );
  NAND2_X2 U1195 ( .A1(n282), .A2(n249), .ZN(n247) );
  CLKBUF_X3 U1196 ( .A(b[18]), .Z(n1241) );
  BUF_X2 U1197 ( .A(a[17]), .Z(n49) );
  OR2_X1 U1198 ( .A1(n663), .A2(n678), .ZN(n1451) );
  AND2_X1 U1199 ( .A1(n521), .A2(n532), .ZN(n1466) );
  BUF_X2 U1200 ( .A(n1431), .Z(n51) );
  BUF_X1 U1201 ( .A(n1277), .Z(n18) );
  BUF_X1 U1202 ( .A(n1274), .Z(n36) );
  BUF_X1 U1203 ( .A(n1274), .Z(n35) );
  BUF_X1 U1204 ( .A(n1273), .Z(n42) );
  BUF_X2 U1205 ( .A(n1287), .Z(n16) );
  BUF_X2 U1206 ( .A(n1287), .Z(n15) );
  BUF_X2 U1207 ( .A(n1270), .Z(n1413) );
  OAI22_X1 U1208 ( .A1(n1413), .A2(n1031), .B1(n58), .B2(n1030), .ZN(n448) );
  NOR2_X1 U1209 ( .A1(n481), .A2(n488), .ZN(n220) );
  AOI21_X1 U1210 ( .B1(n1386), .B2(n401), .A(n398), .ZN(n396) );
  INV_X1 U1211 ( .A(n1466), .ZN(n267) );
  XNOR2_X1 U1212 ( .A(n325), .B(n87), .ZN(product[18]) );
  BUF_X2 U1213 ( .A(n1383), .Z(n65) );
  OR2_X1 U1214 ( .A1(n312), .A2(n317), .ZN(n1387) );
  INV_X1 U1215 ( .A(n282), .ZN(n280) );
  CLKBUF_X1 U1216 ( .A(n318), .Z(n1388) );
  OR2_X1 U1217 ( .A1(n473), .A2(n480), .ZN(n1389) );
  OR2_X1 U1218 ( .A1(n453), .A2(n456), .ZN(n1390) );
  OR2_X1 U1219 ( .A1(n759), .A2(n766), .ZN(n1391) );
  OR2_X1 U1220 ( .A1(n467), .A2(n472), .ZN(n1392) );
  OR2_X1 U1221 ( .A1(n830), .A2(n448), .ZN(n1393) );
  OR2_X1 U1222 ( .A1(n452), .A2(n451), .ZN(n1394) );
  OR2_X1 U1223 ( .A1(n450), .A2(n449), .ZN(n1395) );
  OR2_X1 U1224 ( .A1(n751), .A2(n758), .ZN(n1396) );
  OR2_X1 U1225 ( .A1(n679), .A2(n692), .ZN(n1397) );
  OR2_X1 U1226 ( .A1(n457), .A2(n460), .ZN(n1398) );
  OR2_X1 U1227 ( .A1(n767), .A2(n772), .ZN(n1399) );
  OR2_X1 U1228 ( .A1(n779), .A2(n782), .ZN(n1400) );
  BUF_X2 U1229 ( .A(n1280), .Z(n1484) );
  OR2_X1 U1230 ( .A1(n707), .A2(n718), .ZN(n1401) );
  NOR2_X1 U1231 ( .A1(n461), .A2(n466), .ZN(n179) );
  OR2_X1 U1232 ( .A1(n1029), .A2(n829), .ZN(n1402) );
  NOR2_X1 U1233 ( .A1(n489), .A2(n498), .ZN(n229) );
  NOR2_X1 U1234 ( .A1(n499), .A2(n508), .ZN(n242) );
  BUF_X1 U1235 ( .A(n248), .Z(n1410) );
  XOR2_X1 U1236 ( .A(n630), .B(n615), .Z(n1403) );
  XOR2_X1 U1237 ( .A(n613), .B(n1403), .Z(n611) );
  NAND2_X1 U1238 ( .A1(n613), .A2(n630), .ZN(n1404) );
  NAND2_X1 U1239 ( .A1(n613), .A2(n615), .ZN(n1405) );
  NAND2_X1 U1240 ( .A1(n630), .A2(n615), .ZN(n1406) );
  NAND3_X1 U1241 ( .A1(n1404), .A2(n1405), .A3(n1406), .ZN(n610) );
  XNOR2_X1 U1242 ( .A(n1407), .B(n579), .ZN(n577) );
  XNOR2_X1 U1243 ( .A(n594), .B(n581), .ZN(n1407) );
  CLKBUF_X1 U1244 ( .A(n340), .Z(n1408) );
  OAI22_X1 U1245 ( .A1(n24), .A2(n1157), .B1(n22), .B2(n1156), .ZN(n544) );
  NOR2_X1 U1246 ( .A1(n647), .A2(n662), .ZN(n1409) );
  NOR2_X1 U1247 ( .A1(n647), .A2(n662), .ZN(n323) );
  CLKBUF_X1 U1248 ( .A(n63), .Z(n1411) );
  BUF_X2 U1249 ( .A(n1282), .Z(n45) );
  CLKBUF_X1 U1250 ( .A(n1410), .Z(n1412) );
  CLKBUF_X1 U1251 ( .A(n1270), .Z(n59) );
  XOR2_X1 U1252 ( .A(n583), .B(n598), .Z(n1414) );
  XOR2_X1 U1253 ( .A(n1414), .B(n596), .Z(n579) );
  NAND2_X1 U1254 ( .A1(n583), .A2(n598), .ZN(n1415) );
  NAND2_X1 U1255 ( .A1(n583), .A2(n596), .ZN(n1416) );
  NAND2_X1 U1256 ( .A1(n598), .A2(n596), .ZN(n1417) );
  NAND3_X1 U1257 ( .A1(n1415), .A2(n1416), .A3(n1417), .ZN(n578) );
  NAND2_X1 U1258 ( .A1(n594), .A2(n581), .ZN(n1418) );
  NAND2_X1 U1259 ( .A1(n594), .A2(n579), .ZN(n1419) );
  NAND2_X1 U1260 ( .A1(n581), .A2(n579), .ZN(n1420) );
  NAND3_X1 U1261 ( .A1(n1418), .A2(n1419), .A3(n1420), .ZN(n576) );
  INV_X1 U1262 ( .A(n288), .ZN(n1421) );
  NOR2_X1 U1263 ( .A1(n533), .A2(n546), .ZN(n275) );
  BUF_X2 U1264 ( .A(n1277), .Z(n1437) );
  BUF_X2 U1265 ( .A(n291), .Z(n64) );
  BUF_X2 U1266 ( .A(n1273), .Z(n1422) );
  CLKBUF_X1 U1267 ( .A(n1273), .Z(n41) );
  INV_X1 U1268 ( .A(n55), .ZN(n1423) );
  INV_X2 U1269 ( .A(n1423), .ZN(n1424) );
  CLKBUF_X1 U1270 ( .A(b[0]), .Z(n61) );
  XNOR2_X1 U1271 ( .A(n55), .B(n1258), .ZN(n1425) );
  CLKBUF_X1 U1272 ( .A(n1283), .Z(n40) );
  XNOR2_X1 U1273 ( .A(n1257), .B(n55), .ZN(n1426) );
  CLKBUF_X1 U1274 ( .A(n317), .Z(n1427) );
  CLKBUF_X1 U1275 ( .A(n19), .Z(n1428) );
  CLKBUF_X1 U1276 ( .A(n1278), .Z(n12) );
  XNOR2_X1 U1277 ( .A(n13), .B(n1242), .ZN(n1430) );
  XNOR2_X1 U1278 ( .A(a[16]), .B(a[15]), .ZN(n1431) );
  BUF_X1 U1279 ( .A(n1274), .Z(n1432) );
  CLKBUF_X1 U1280 ( .A(n311), .Z(n1433) );
  CLKBUF_X1 U1281 ( .A(n1288), .Z(n9) );
  CLKBUF_X1 U1282 ( .A(n1240), .Z(n1434) );
  CLKBUF_X1 U1283 ( .A(n303), .Z(n1435) );
  CLKBUF_X1 U1284 ( .A(n49), .Z(n1436) );
  BUF_X1 U1285 ( .A(n61), .Z(n1438) );
  CLKBUF_X1 U1286 ( .A(n48), .Z(n1439) );
  CLKBUF_X1 U1287 ( .A(n13), .Z(n1440) );
  XNOR2_X1 U1288 ( .A(n1), .B(n1240), .ZN(n1441) );
  XNOR2_X1 U1289 ( .A(n244), .B(n1442), .ZN(product[28]) );
  AND2_X1 U1290 ( .A1(n240), .A2(n243), .ZN(n1442) );
  XNOR2_X1 U1291 ( .A(n268), .B(n1443), .ZN(product[26]) );
  AND2_X1 U1292 ( .A1(n262), .A2(n267), .ZN(n1443) );
  CLKBUF_X1 U1293 ( .A(n388), .Z(n1444) );
  XNOR2_X1 U1294 ( .A(n222), .B(n1445), .ZN(product[30]) );
  AND2_X1 U1295 ( .A1(n418), .A2(n221), .ZN(n1445) );
  CLKBUF_X1 U1296 ( .A(n313), .Z(n1446) );
  XNOR2_X1 U1297 ( .A(n231), .B(n1447), .ZN(product[29]) );
  AND2_X1 U1298 ( .A1(n227), .A2(n230), .ZN(n1447) );
  CLKBUF_X1 U1299 ( .A(n283), .Z(n1448) );
  XNOR2_X1 U1300 ( .A(n277), .B(n1449), .ZN(product[25]) );
  AND2_X1 U1301 ( .A1(n273), .A2(n276), .ZN(n1449) );
  XNOR2_X1 U1302 ( .A(n257), .B(n1450), .ZN(product[27]) );
  AND2_X1 U1303 ( .A1(n1482), .A2(n256), .ZN(n1450) );
  CLKBUF_X1 U1304 ( .A(n367), .Z(n1452) );
  NOR2_X1 U1305 ( .A1(n707), .A2(n718), .ZN(n1453) );
  NOR2_X1 U1306 ( .A1(n707), .A2(n718), .ZN(n350) );
  NAND2_X1 U1307 ( .A1(n561), .A2(n576), .ZN(n290) );
  NOR2_X1 U1308 ( .A1(n561), .A2(n576), .ZN(n289) );
  XNOR2_X1 U1309 ( .A(n43), .B(n1255), .ZN(n1454) );
  BUF_X2 U1310 ( .A(a[15]), .Z(n43) );
  BUF_X2 U1311 ( .A(n1276), .Z(n23) );
  CLKBUF_X3 U1312 ( .A(n1284), .Z(n33) );
  NOR2_X1 U1313 ( .A1(n593), .A2(n610), .ZN(n303) );
  AND2_X1 U1314 ( .A1(n663), .A2(n678), .ZN(n1455) );
  CLKBUF_X1 U1315 ( .A(n39), .Z(n1456) );
  CLKBUF_X2 U1316 ( .A(n39), .Z(n1457) );
  BUF_X1 U1317 ( .A(n39), .Z(n1458) );
  BUF_X1 U1318 ( .A(n1086), .Z(n1459) );
  CLKBUF_X3 U1319 ( .A(a[15]), .Z(n1460) );
  XOR2_X1 U1320 ( .A(n675), .B(n673), .Z(n1461) );
  XOR2_X1 U1321 ( .A(n684), .B(n1461), .Z(n667) );
  NAND2_X1 U1322 ( .A1(n684), .A2(n675), .ZN(n1462) );
  NAND2_X1 U1323 ( .A1(n684), .A2(n673), .ZN(n1463) );
  NAND2_X1 U1324 ( .A1(n675), .A2(n673), .ZN(n1464) );
  NAND3_X1 U1325 ( .A1(n1462), .A2(n1463), .A3(n1464), .ZN(n666) );
  CLKBUF_X1 U1326 ( .A(n1451), .Z(n1465) );
  INV_X1 U1327 ( .A(n1455), .ZN(n1467) );
  BUF_X1 U1328 ( .A(n304), .Z(n1468) );
  CLKBUF_X3 U1329 ( .A(b[3]), .Z(n1256) );
  CLKBUF_X3 U1330 ( .A(n61), .Z(n1494) );
  CLKBUF_X3 U1331 ( .A(b[17]), .Z(n1242) );
  NAND2_X1 U1332 ( .A1(n1261), .A2(n1281), .ZN(n1271) );
  OR2_X2 U1333 ( .A1(n693), .A2(n706), .ZN(n1469) );
  NOR2_X2 U1334 ( .A1(n731), .A2(n740), .ZN(n361) );
  CLKBUF_X1 U1335 ( .A(n336), .Z(n1470) );
  XOR2_X1 U1336 ( .A(n846), .B(n972), .Z(n1471) );
  XOR2_X1 U1337 ( .A(n900), .B(n1471), .Z(n607) );
  NAND2_X1 U1338 ( .A1(n900), .A2(n846), .ZN(n1472) );
  NAND2_X1 U1339 ( .A1(n900), .A2(n972), .ZN(n1473) );
  NAND2_X1 U1340 ( .A1(n846), .A2(n972), .ZN(n1474) );
  NAND3_X1 U1341 ( .A1(n1472), .A2(n1473), .A3(n1474), .ZN(n606) );
  CLKBUF_X1 U1342 ( .A(n1256), .Z(n1475) );
  BUF_X2 U1343 ( .A(n40), .Z(n1476) );
  NOR2_X2 U1344 ( .A1(n547), .A2(n560), .ZN(n284) );
  XOR2_X1 U1345 ( .A(n960), .B(n906), .Z(n1477) );
  XOR2_X1 U1346 ( .A(n924), .B(n1477), .Z(n703) );
  NAND2_X1 U1347 ( .A1(n924), .A2(n960), .ZN(n1478) );
  NAND2_X1 U1348 ( .A1(n924), .A2(n906), .ZN(n1479) );
  NAND2_X1 U1349 ( .A1(n960), .A2(n906), .ZN(n1480) );
  NAND3_X1 U1350 ( .A1(n1478), .A2(n1479), .A3(n1480), .ZN(n702) );
  BUF_X4 U1351 ( .A(a[5]), .Z(n13) );
  BUF_X1 U1352 ( .A(n1283), .Z(n39) );
  OAI22_X1 U1353 ( .A1(n1422), .A2(n1094), .B1(n1476), .B2(n1093), .ZN(n478)
         );
  NOR2_X1 U1354 ( .A1(n577), .A2(n592), .ZN(n1481) );
  NOR2_X1 U1355 ( .A1(n577), .A2(n592), .ZN(n296) );
  CLKBUF_X3 U1356 ( .A(b[10]), .Z(n1249) );
  CLKBUF_X3 U1357 ( .A(b[1]), .Z(n1258) );
  BUF_X4 U1358 ( .A(a[3]), .Z(n7) );
  CLKBUF_X3 U1359 ( .A(b[12]), .Z(n1247) );
  OR2_X2 U1360 ( .A1(n509), .A2(n520), .ZN(n1482) );
  BUF_X1 U1361 ( .A(n1288), .Z(n10) );
  CLKBUF_X3 U1362 ( .A(b[7]), .Z(n1252) );
  NAND2_X1 U1363 ( .A1(n1260), .A2(n1280), .ZN(n1270) );
  CLKBUF_X3 U1364 ( .A(n1286), .Z(n21) );
  CLKBUF_X3 U1365 ( .A(n1286), .Z(n22) );
  NAND2_X1 U1366 ( .A1(n1266), .A2(n1286), .ZN(n1276) );
  NOR2_X1 U1367 ( .A1(n611), .A2(n628), .ZN(n1483) );
  OR2_X1 U1368 ( .A1(n521), .A2(n532), .ZN(n1485) );
  XNOR2_X1 U1369 ( .A(a[1]), .B(a[2]), .ZN(n1288) );
  NAND2_X1 U1370 ( .A1(n1268), .A2(n1288), .ZN(n1278) );
  XNOR2_X1 U1371 ( .A(n209), .B(n1486), .ZN(product[31]) );
  AND2_X1 U1372 ( .A1(n1389), .A2(n208), .ZN(n1486) );
  BUF_X1 U1373 ( .A(n61), .Z(n1487) );
  BUF_X1 U1374 ( .A(n61), .Z(n1488) );
  AOI21_X1 U1375 ( .B1(n1465), .B2(n1470), .A(n1455), .ZN(n1489) );
  XNOR2_X1 U1376 ( .A(n339), .B(n1490), .ZN(product[16]) );
  AND2_X1 U1377 ( .A1(n1397), .A2(n338), .ZN(n1490) );
  XNOR2_X1 U1378 ( .A(n286), .B(n1491), .ZN(product[24]) );
  AND2_X1 U1379 ( .A1(n424), .A2(n285), .ZN(n1491) );
  NOR2_X1 U1380 ( .A1(n229), .A2(n220), .ZN(n218) );
  NOR2_X1 U1381 ( .A1(n179), .A2(n151), .ZN(n149) );
  NAND2_X1 U1382 ( .A1(n533), .A2(n546), .ZN(n276) );
  NAND2_X1 U1383 ( .A1(n593), .A2(n610), .ZN(n304) );
  INV_X1 U1384 ( .A(n242), .ZN(n240) );
  NOR2_X1 U1385 ( .A1(n741), .A2(n750), .ZN(n364) );
  NAND2_X1 U1386 ( .A1(n489), .A2(n498), .ZN(n230) );
  NAND2_X1 U1387 ( .A1(n751), .A2(n758), .ZN(n373) );
  NOR2_X1 U1388 ( .A1(n1028), .A2(n1009), .ZN(n406) );
  NOR2_X1 U1389 ( .A1(n783), .A2(n786), .ZN(n394) );
  NOR2_X1 U1390 ( .A1(n773), .A2(n778), .ZN(n386) );
  NAND2_X1 U1391 ( .A1(n779), .A2(n782), .ZN(n392) );
  NOR2_X1 U1392 ( .A1(n789), .A2(n828), .ZN(n402) );
  AND2_X1 U1393 ( .A1(n1402), .A2(n409), .ZN(product[1]) );
  BUF_X2 U1394 ( .A(n1279), .Z(n6) );
  BUF_X2 U1395 ( .A(n1272), .Z(n48) );
  BUF_X2 U1396 ( .A(n1275), .Z(n29) );
  BUF_X2 U1397 ( .A(n1272), .Z(n47) );
  BUF_X2 U1398 ( .A(n1270), .Z(n60) );
  NAND2_X1 U1399 ( .A1(n1267), .A2(n1287), .ZN(n1277) );
  INV_X1 U1400 ( .A(a[0]), .ZN(n1289) );
  NOR2_X1 U1401 ( .A1(n280), .A2(n271), .ZN(n269) );
  NOR2_X1 U1402 ( .A1(n280), .A2(n260), .ZN(n258) );
  NAND2_X1 U1403 ( .A1(n214), .A2(n134), .ZN(n130) );
  INV_X1 U1404 ( .A(n280), .ZN(n278) );
  INV_X1 U1405 ( .A(n173), .ZN(n171) );
  INV_X1 U1406 ( .A(n186), .ZN(n184) );
  INV_X1 U1407 ( .A(n1387), .ZN(n306) );
  NOR2_X1 U1408 ( .A1(n216), .A2(n192), .ZN(n186) );
  NOR2_X1 U1409 ( .A1(n216), .A2(n175), .ZN(n173) );
  OAI21_X1 U1410 ( .B1(n281), .B2(n260), .A(n261), .ZN(n259) );
  AOI21_X1 U1411 ( .B1(n274), .B2(n262), .A(n1466), .ZN(n261) );
  INV_X1 U1412 ( .A(n187), .ZN(n185) );
  INV_X1 U1413 ( .A(n1448), .ZN(n281) );
  INV_X1 U1414 ( .A(n216), .ZN(n214) );
  INV_X1 U1415 ( .A(n1433), .ZN(n309) );
  NAND2_X1 U1416 ( .A1(n1485), .A2(n1482), .ZN(n251) );
  NAND2_X1 U1417 ( .A1(n273), .A2(n262), .ZN(n260) );
  OAI21_X1 U1418 ( .B1(n281), .B2(n271), .A(n276), .ZN(n270) );
  INV_X1 U1419 ( .A(n273), .ZN(n271) );
  NAND2_X1 U1420 ( .A1(n1451), .A2(n1397), .ZN(n326) );
  NOR2_X1 U1421 ( .A1(n1387), .A2(n1435), .ZN(n299) );
  INV_X1 U1422 ( .A(n263), .ZN(n262) );
  INV_X1 U1423 ( .A(n1485), .ZN(n263) );
  INV_X1 U1424 ( .A(n192), .ZN(n190) );
  NAND2_X1 U1425 ( .A1(n186), .A2(n149), .ZN(n145) );
  INV_X1 U1426 ( .A(n1470), .ZN(n334) );
  INV_X1 U1427 ( .A(n119), .ZN(n117) );
  INV_X1 U1428 ( .A(n1397), .ZN(n333) );
  NAND2_X1 U1429 ( .A1(n214), .A2(n1389), .ZN(n201) );
  INV_X1 U1430 ( .A(n65), .ZN(n246) );
  XOR2_X1 U1431 ( .A(n347), .B(n90), .Z(product[15]) );
  NAND2_X1 U1432 ( .A1(n1469), .A2(n346), .ZN(n90) );
  NAND2_X1 U1433 ( .A1(n315), .A2(n1388), .ZN(n86) );
  XNOR2_X1 U1434 ( .A(n332), .B(n88), .ZN(product[17]) );
  NAND2_X1 U1435 ( .A1(n1465), .A2(n1467), .ZN(n88) );
  OAI21_X1 U1436 ( .B1(n339), .B2(n333), .A(n334), .ZN(n332) );
  XOR2_X1 U1437 ( .A(n352), .B(n91), .Z(product[14]) );
  NAND2_X1 U1438 ( .A1(n1401), .A2(n351), .ZN(n91) );
  AOI21_X1 U1439 ( .B1(n357), .B2(n435), .A(n354), .ZN(n352) );
  AOI21_X1 U1440 ( .B1(n1451), .B2(n336), .A(n1455), .ZN(n327) );
  NAND2_X1 U1441 ( .A1(n425), .A2(n1421), .ZN(n82) );
  INV_X1 U1442 ( .A(n289), .ZN(n425) );
  OAI21_X1 U1443 ( .B1(n284), .B2(n290), .A(n285), .ZN(n283) );
  OAI21_X1 U1444 ( .B1(n217), .B2(n192), .A(n193), .ZN(n187) );
  NAND2_X1 U1445 ( .A1(n428), .A2(n1446), .ZN(n85) );
  INV_X1 U1446 ( .A(n312), .ZN(n428) );
  INV_X1 U1447 ( .A(n284), .ZN(n424) );
  XOR2_X1 U1448 ( .A(n305), .B(n84), .Z(product[21]) );
  NAND2_X1 U1449 ( .A1(n302), .A2(n1468), .ZN(n84) );
  XOR2_X1 U1450 ( .A(n298), .B(n83), .Z(product[22]) );
  NAND2_X1 U1451 ( .A1(n426), .A2(n297), .ZN(n83) );
  NAND2_X1 U1452 ( .A1(n218), .A2(n240), .ZN(n216) );
  AOI21_X1 U1453 ( .B1(n215), .B2(n1389), .A(n206), .ZN(n202) );
  INV_X1 U1454 ( .A(n174), .ZN(n172) );
  AOI21_X1 U1455 ( .B1(n283), .B2(n249), .A(n250), .ZN(n248) );
  OAI21_X1 U1456 ( .B1(n251), .B2(n276), .A(n252), .ZN(n250) );
  AOI21_X1 U1457 ( .B1(n1482), .B2(n1466), .A(n254), .ZN(n252) );
  INV_X1 U1458 ( .A(n358), .ZN(n357) );
  NAND2_X1 U1459 ( .A1(n430), .A2(n324), .ZN(n87) );
  OAI21_X1 U1460 ( .B1(n339), .B2(n326), .A(n1489), .ZN(n325) );
  INV_X1 U1461 ( .A(n1409), .ZN(n430) );
  INV_X1 U1462 ( .A(n380), .ZN(n379) );
  NOR2_X1 U1463 ( .A1(n192), .A2(n136), .ZN(n134) );
  INV_X1 U1464 ( .A(n217), .ZN(n215) );
  NOR2_X1 U1465 ( .A1(n216), .A2(n121), .ZN(n119) );
  INV_X1 U1466 ( .A(n275), .ZN(n273) );
  NAND2_X1 U1467 ( .A1(n190), .A2(n177), .ZN(n175) );
  NAND2_X1 U1468 ( .A1(n1389), .A2(n1392), .ZN(n192) );
  OAI21_X1 U1469 ( .B1(n309), .B2(n1435), .A(n1468), .ZN(n300) );
  INV_X1 U1470 ( .A(n1452), .ZN(n366) );
  INV_X1 U1471 ( .A(n276), .ZN(n274) );
  INV_X1 U1472 ( .A(n1435), .ZN(n302) );
  INV_X1 U1473 ( .A(n193), .ZN(n191) );
  NAND2_X1 U1474 ( .A1(n240), .A2(n227), .ZN(n225) );
  NAND2_X1 U1475 ( .A1(n173), .A2(n1398), .ZN(n160) );
  INV_X1 U1476 ( .A(n256), .ZN(n254) );
  INV_X1 U1477 ( .A(n346), .ZN(n344) );
  INV_X1 U1478 ( .A(n290), .ZN(n288) );
  INV_X1 U1479 ( .A(n1388), .ZN(n316) );
  NAND2_X1 U1480 ( .A1(n1399), .A2(n384), .ZN(n97) );
  INV_X1 U1481 ( .A(n384), .ZN(n382) );
  XOR2_X1 U1482 ( .A(n366), .B(n94), .Z(product[11]) );
  NAND2_X1 U1483 ( .A1(n437), .A2(n365), .ZN(n94) );
  INV_X1 U1484 ( .A(n364), .ZN(n437) );
  AOI21_X2 U1485 ( .B1(n218), .B2(n241), .A(n219), .ZN(n217) );
  OAI21_X1 U1486 ( .B1(n230), .B2(n220), .A(n221), .ZN(n219) );
  XNOR2_X1 U1487 ( .A(n363), .B(n93), .ZN(product[12]) );
  NAND2_X1 U1488 ( .A1(n436), .A2(n362), .ZN(n93) );
  OAI21_X1 U1489 ( .B1(n366), .B2(n364), .A(n365), .ZN(n363) );
  INV_X1 U1490 ( .A(n361), .ZN(n436) );
  XNOR2_X1 U1491 ( .A(n379), .B(n96), .ZN(product[9]) );
  NAND2_X1 U1492 ( .A1(n1391), .A2(n378), .ZN(n96) );
  XNOR2_X1 U1493 ( .A(n357), .B(n92), .ZN(product[13]) );
  NAND2_X1 U1494 ( .A1(n435), .A2(n356), .ZN(n92) );
  INV_X1 U1495 ( .A(n355), .ZN(n435) );
  OAI21_X1 U1496 ( .B1(n368), .B2(n380), .A(n369), .ZN(n367) );
  AOI21_X1 U1497 ( .B1(n215), .B2(n134), .A(n135), .ZN(n131) );
  INV_X1 U1498 ( .A(n120), .ZN(n118) );
  AOI21_X1 U1499 ( .B1(n187), .B2(n149), .A(n150), .ZN(n146) );
  AOI21_X1 U1500 ( .B1(n174), .B2(n1398), .A(n165), .ZN(n161) );
  NAND2_X1 U1501 ( .A1(n177), .A2(n180), .ZN(n72) );
  NAND2_X1 U1502 ( .A1(n1392), .A2(n197), .ZN(n73) );
  INV_X1 U1503 ( .A(n220), .ZN(n418) );
  AOI21_X1 U1504 ( .B1(n1392), .B2(n206), .A(n195), .ZN(n193) );
  INV_X1 U1505 ( .A(n197), .ZN(n195) );
  OAI21_X1 U1506 ( .B1(n217), .B2(n175), .A(n176), .ZN(n174) );
  AOI21_X1 U1507 ( .B1(n191), .B2(n177), .A(n178), .ZN(n176) );
  INV_X1 U1508 ( .A(n180), .ZN(n178) );
  NOR2_X1 U1509 ( .A1(n629), .A2(n646), .ZN(n317) );
  NOR2_X1 U1510 ( .A1(n611), .A2(n628), .ZN(n312) );
  NAND2_X1 U1511 ( .A1(n134), .A2(n1395), .ZN(n121) );
  AOI21_X1 U1512 ( .B1(n367), .B2(n359), .A(n360), .ZN(n358) );
  NOR2_X1 U1513 ( .A1(n361), .A2(n364), .ZN(n359) );
  OAI21_X1 U1514 ( .B1(n361), .B2(n365), .A(n362), .ZN(n360) );
  AOI21_X1 U1515 ( .B1(n241), .B2(n227), .A(n228), .ZN(n226) );
  INV_X1 U1516 ( .A(n230), .ZN(n228) );
  XOR2_X1 U1517 ( .A(n374), .B(n95), .Z(product[10]) );
  NAND2_X1 U1518 ( .A1(n1396), .A2(n373), .ZN(n95) );
  AOI21_X1 U1519 ( .B1(n379), .B2(n1391), .A(n376), .ZN(n374) );
  NAND2_X1 U1520 ( .A1(n629), .A2(n646), .ZN(n318) );
  NAND2_X1 U1521 ( .A1(n509), .A2(n520), .ZN(n256) );
  NAND2_X1 U1522 ( .A1(n547), .A2(n560), .ZN(n285) );
  INV_X1 U1523 ( .A(n179), .ZN(n177) );
  INV_X1 U1524 ( .A(n229), .ZN(n227) );
  NAND2_X1 U1525 ( .A1(n1398), .A2(n1390), .ZN(n151) );
  NAND2_X1 U1526 ( .A1(n149), .A2(n1394), .ZN(n136) );
  NAND2_X1 U1527 ( .A1(n679), .A2(n692), .ZN(n338) );
  NAND2_X1 U1528 ( .A1(n647), .A2(n662), .ZN(n324) );
  NAND2_X1 U1529 ( .A1(n611), .A2(n628), .ZN(n313) );
  NAND2_X1 U1530 ( .A1(n577), .A2(n592), .ZN(n297) );
  INV_X1 U1531 ( .A(n243), .ZN(n241) );
  INV_X1 U1532 ( .A(n208), .ZN(n206) );
  AOI21_X1 U1533 ( .B1(n1411), .B2(n106), .A(n107), .ZN(n105) );
  INV_X1 U1534 ( .A(n378), .ZN(n376) );
  INV_X1 U1535 ( .A(n356), .ZN(n354) );
  INV_X1 U1536 ( .A(n373), .ZN(n371) );
  NAND2_X1 U1537 ( .A1(n443), .A2(n395), .ZN(n100) );
  INV_X1 U1538 ( .A(n394), .ZN(n443) );
  XOR2_X1 U1539 ( .A(n114), .B(n67), .Z(product[38]) );
  NAND2_X1 U1540 ( .A1(n1393), .A2(n113), .ZN(n67) );
  AOI21_X1 U1541 ( .B1(n63), .B2(n115), .A(n116), .ZN(n114) );
  INV_X1 U1542 ( .A(n392), .ZN(n390) );
  XOR2_X1 U1543 ( .A(n168), .B(n71), .Z(product[34]) );
  NAND2_X1 U1544 ( .A1(n1398), .A2(n167), .ZN(n71) );
  XOR2_X1 U1545 ( .A(n127), .B(n68), .Z(product[37]) );
  NAND2_X1 U1546 ( .A1(n1395), .A2(n126), .ZN(n68) );
  AOI21_X1 U1547 ( .B1(n63), .B2(n128), .A(n129), .ZN(n127) );
  XOR2_X1 U1548 ( .A(n142), .B(n69), .Z(product[36]) );
  NAND2_X1 U1549 ( .A1(n1394), .A2(n141), .ZN(n69) );
  AOI21_X1 U1550 ( .B1(n63), .B2(n143), .A(n144), .ZN(n142) );
  XOR2_X1 U1551 ( .A(n157), .B(n70), .Z(product[35]) );
  NAND2_X1 U1552 ( .A1(n1390), .A2(n156), .ZN(n70) );
  AOI21_X1 U1553 ( .B1(n63), .B2(n158), .A(n159), .ZN(n157) );
  NOR2_X1 U1554 ( .A1(n719), .A2(n730), .ZN(n355) );
  OAI21_X1 U1555 ( .B1(n193), .B2(n136), .A(n137), .ZN(n135) );
  AOI21_X1 U1556 ( .B1(n150), .B2(n1394), .A(n139), .ZN(n137) );
  INV_X1 U1557 ( .A(n141), .ZN(n139) );
  OAI21_X1 U1558 ( .B1(n217), .B2(n121), .A(n122), .ZN(n120) );
  AOI21_X1 U1559 ( .B1(n135), .B2(n1395), .A(n124), .ZN(n122) );
  INV_X1 U1560 ( .A(n126), .ZN(n124) );
  OAI21_X1 U1561 ( .B1(n151), .B2(n180), .A(n152), .ZN(n150) );
  AOI21_X1 U1562 ( .B1(n165), .B2(n1390), .A(n154), .ZN(n152) );
  INV_X1 U1563 ( .A(n156), .ZN(n154) );
  OAI21_X1 U1564 ( .B1(n388), .B2(n386), .A(n387), .ZN(n385) );
  NAND2_X1 U1565 ( .A1(n461), .A2(n466), .ZN(n180) );
  NAND2_X1 U1566 ( .A1(n741), .A2(n750), .ZN(n365) );
  NAND2_X1 U1567 ( .A1(n719), .A2(n730), .ZN(n356) );
  AOI21_X1 U1568 ( .B1(n120), .B2(n1393), .A(n111), .ZN(n109) );
  INV_X1 U1569 ( .A(n113), .ZN(n111) );
  NAND2_X1 U1570 ( .A1(n499), .A2(n508), .ZN(n243) );
  NAND2_X1 U1571 ( .A1(n473), .A2(n480), .ZN(n208) );
  NAND2_X1 U1572 ( .A1(n467), .A2(n472), .ZN(n197) );
  NAND2_X1 U1573 ( .A1(n481), .A2(n488), .ZN(n221) );
  NAND2_X1 U1574 ( .A1(n731), .A2(n740), .ZN(n362) );
  NAND2_X1 U1575 ( .A1(n759), .A2(n766), .ZN(n378) );
  NAND2_X1 U1576 ( .A1(n767), .A2(n772), .ZN(n384) );
  INV_X1 U1577 ( .A(n167), .ZN(n165) );
  NAND2_X1 U1578 ( .A1(n441), .A2(n387), .ZN(n98) );
  INV_X1 U1579 ( .A(n386), .ZN(n441) );
  NAND2_X1 U1580 ( .A1(n1400), .A2(n392), .ZN(n99) );
  XOR2_X1 U1581 ( .A(n102), .B(n404), .Z(product[3]) );
  NAND2_X1 U1582 ( .A1(n445), .A2(n403), .ZN(n102) );
  INV_X1 U1583 ( .A(n402), .ZN(n445) );
  XOR2_X1 U1584 ( .A(n103), .B(n409), .Z(product[2]) );
  NAND2_X1 U1585 ( .A1(n446), .A2(n407), .ZN(n103) );
  INV_X1 U1586 ( .A(n406), .ZN(n446) );
  XNOR2_X1 U1587 ( .A(n101), .B(n401), .ZN(product[4]) );
  NAND2_X1 U1588 ( .A1(n1386), .A2(n400), .ZN(n101) );
  OAI21_X1 U1589 ( .B1(n402), .B2(n404), .A(n403), .ZN(n401) );
  NAND2_X1 U1590 ( .A1(n830), .A2(n448), .ZN(n113) );
  INV_X1 U1591 ( .A(n448), .ZN(n449) );
  INV_X1 U1592 ( .A(n400), .ZN(n398) );
  NAND2_X1 U1593 ( .A1(n1028), .A2(n1009), .ZN(n407) );
  INV_X1 U1594 ( .A(n544), .ZN(n545) );
  INV_X1 U1595 ( .A(n478), .ZN(n479) );
  OR2_X1 U1596 ( .A1(n937), .A2(n865), .ZN(n626) );
  XNOR2_X1 U1597 ( .A(n937), .B(n865), .ZN(n627) );
  NAND2_X1 U1598 ( .A1(n457), .A2(n460), .ZN(n167) );
  NAND2_X1 U1599 ( .A1(n452), .A2(n451), .ZN(n141) );
  NAND2_X1 U1600 ( .A1(n450), .A2(n449), .ZN(n126) );
  NAND2_X1 U1601 ( .A1(n453), .A2(n456), .ZN(n156) );
  NAND2_X1 U1602 ( .A1(n773), .A2(n778), .ZN(n387) );
  NAND2_X1 U1603 ( .A1(n783), .A2(n786), .ZN(n395) );
  INV_X1 U1604 ( .A(n405), .ZN(n404) );
  OAI21_X1 U1605 ( .B1(n406), .B2(n409), .A(n407), .ZN(n405) );
  OAI22_X1 U1606 ( .A1(n54), .A2(n1052), .B1(n52), .B2(n1051), .ZN(n454) );
  OAI22_X1 U1607 ( .A1(n36), .A2(n1115), .B1(n34), .B2(n1114), .ZN(n496) );
  OAI22_X1 U1608 ( .A1(n5), .A2(n1237), .B1(n1236), .B2(n3), .ZN(n1028) );
  OAI22_X1 U1609 ( .A1(n11), .A2(n1199), .B1(n1198), .B2(n10), .ZN(n608) );
  OAI22_X1 U1610 ( .A1(n30), .A2(n1136), .B1(n28), .B2(n1135), .ZN(n518) );
  OAI22_X1 U1611 ( .A1(n1437), .A2(n1178), .B1(n16), .B2(n1177), .ZN(n574) );
  OAI22_X1 U1612 ( .A1(n1439), .A2(n1073), .B1(n46), .B2(n1072), .ZN(n464) );
  OAI22_X1 U1613 ( .A1(n53), .A2(n1067), .B1(n51), .B2(n1066), .ZN(n865) );
  OAI22_X1 U1614 ( .A1(n30), .A2(n1143), .B1(n28), .B2(n1142), .ZN(n937) );
  OAI22_X1 U1615 ( .A1(n60), .A2(n1032), .B1(n58), .B2(n1031), .ZN(n831) );
  INV_X1 U1616 ( .A(n793), .ZN(n850) );
  AOI21_X1 U1617 ( .B1(n54), .B2(n52), .A(n1051), .ZN(n793) );
  OAI22_X1 U1618 ( .A1(n5), .A2(n1234), .B1(n1233), .B2(n3), .ZN(n1025) );
  OAI22_X1 U1619 ( .A1(n1429), .A2(n1215), .B1(n9), .B2(n1214), .ZN(n1006) );
  OAI22_X1 U1620 ( .A1(n1413), .A2(n1034), .B1(n58), .B2(n1033), .ZN(n833) );
  OAI22_X1 U1621 ( .A1(n17), .A2(n1195), .B1(n15), .B2(n1194), .ZN(n987) );
  OAI22_X1 U1622 ( .A1(n30), .A2(n1295), .B1(n1155), .B2(n28), .ZN(n825) );
  OAI22_X1 U1623 ( .A1(n29), .A2(n1154), .B1(n27), .B2(n1153), .ZN(n948) );
  OR2_X1 U1624 ( .A1(n1438), .A2(n1295), .ZN(n1155) );
  OAI22_X1 U1625 ( .A1(n48), .A2(n1459), .B1(n45), .B2(n1085), .ZN(n883) );
  OAI22_X1 U1626 ( .A1(n1422), .A2(n1105), .B1(n1458), .B2(n1104), .ZN(n901)
         );
  OAI22_X1 U1627 ( .A1(n11), .A2(n1200), .B1(n10), .B2(n1199), .ZN(n991) );
  OAI22_X1 U1628 ( .A1(n30), .A2(n1140), .B1(n28), .B2(n1139), .ZN(n934) );
  OAI22_X1 U1629 ( .A1(n48), .A2(n1083), .B1(n45), .B2(n1082), .ZN(n880) );
  OAI22_X1 U1630 ( .A1(n24), .A2(n1159), .B1(n22), .B2(n1158), .ZN(n952) );
  OAI22_X1 U1631 ( .A1(n29), .A2(n1149), .B1(n27), .B2(n1148), .ZN(n943) );
  OAI22_X1 U1632 ( .A1(n1422), .A2(n1111), .B1(n1458), .B2(n1110), .ZN(n907)
         );
  OAI22_X1 U1633 ( .A1(n1429), .A2(n1206), .B1(n10), .B2(n1205), .ZN(n997) );
  OAI22_X1 U1634 ( .A1(n36), .A2(n1129), .B1(n33), .B2(n1128), .ZN(n924) );
  OAI22_X1 U1635 ( .A1(n1422), .A2(n1110), .B1(n1109), .B2(n1457), .ZN(n906)
         );
  OAI22_X1 U1636 ( .A1(n23), .A2(n1167), .B1(n1166), .B2(n21), .ZN(n960) );
  OAI22_X1 U1637 ( .A1(n53), .A2(n1065), .B1(n51), .B2(n1064), .ZN(n863) );
  OAI22_X1 U1638 ( .A1(n24), .A2(n1160), .B1(n22), .B2(n1159), .ZN(n953) );
  OAI22_X1 U1639 ( .A1(n24), .A2(n1296), .B1(n1176), .B2(n22), .ZN(n826) );
  OAI22_X1 U1640 ( .A1(n23), .A2(n1175), .B1(n21), .B2(n1174), .ZN(n968) );
  OR2_X1 U1641 ( .A1(n1488), .A2(n1296), .ZN(n1176) );
  OAI22_X1 U1642 ( .A1(n29), .A2(n1145), .B1(n27), .B2(n1144), .ZN(n939) );
  OAI22_X1 U1643 ( .A1(n35), .A2(n1126), .B1(n33), .B2(n1125), .ZN(n921) );
  OAI22_X1 U1644 ( .A1(n18), .A2(n1183), .B1(n16), .B2(n1182), .ZN(n975) );
  OAI22_X1 U1645 ( .A1(n29), .A2(n1153), .B1(n27), .B2(n1152), .ZN(n947) );
  OAI22_X1 U1646 ( .A1(n17), .A2(n1191), .B1(n15), .B2(n1190), .ZN(n983) );
  OAI22_X1 U1647 ( .A1(n1429), .A2(n1210), .B1(n9), .B2(n1209), .ZN(n1001) );
  AND2_X1 U1648 ( .A1(n1488), .A2(n794), .ZN(n869) );
  OAI22_X1 U1649 ( .A1(n42), .A2(n1109), .B1(n1108), .B2(n1458), .ZN(n905) );
  OAI22_X1 U1650 ( .A1(n6), .A2(n1223), .B1(n1222), .B2(n4), .ZN(n1014) );
  OAI22_X1 U1651 ( .A1(n29), .A2(n1148), .B1(n1147), .B2(n27), .ZN(n942) );
  OAI22_X1 U1652 ( .A1(n6), .A2(n1224), .B1(n1223), .B2(n4), .ZN(n1015) );
  OAI22_X1 U1653 ( .A1(n18), .A2(n1186), .B1(n16), .B2(n1185), .ZN(n978) );
  OAI22_X1 U1654 ( .A1(n36), .A2(n1125), .B1(n33), .B2(n1124), .ZN(n920) );
  OAI22_X1 U1655 ( .A1(n11), .A2(n1201), .B1(n10), .B2(n1200), .ZN(n992) );
  OAI22_X1 U1656 ( .A1(n1437), .A2(n1182), .B1(n16), .B2(n1181), .ZN(n974) );
  AND2_X1 U1657 ( .A1(n1488), .A2(n812), .ZN(n989) );
  OAI22_X1 U1658 ( .A1(n5), .A2(n1235), .B1(n1234), .B2(n3), .ZN(n1026) );
  OAI22_X1 U1659 ( .A1(n11), .A2(n1216), .B1(n9), .B2(n1215), .ZN(n1007) );
  AOI21_X1 U1660 ( .B1(n12), .B2(n10), .A(n1198), .ZN(n814) );
  AOI21_X1 U1661 ( .B1(n1432), .B2(n34), .A(n1114), .ZN(n802) );
  AOI21_X1 U1662 ( .B1(n6), .B2(n4), .A(n1219), .ZN(n817) );
  AOI21_X1 U1663 ( .B1(n41), .B2(n1476), .A(n1093), .ZN(n799) );
  OAI22_X1 U1664 ( .A1(n36), .A2(n1294), .B1(n1134), .B2(n34), .ZN(n824) );
  OAI22_X1 U1665 ( .A1(n36), .A2(n1133), .B1(n33), .B2(n1132), .ZN(n928) );
  OR2_X1 U1666 ( .A1(n1488), .A2(n1294), .ZN(n1134) );
  NAND2_X1 U1667 ( .A1(n1029), .A2(n829), .ZN(n409) );
  OAI22_X1 U1668 ( .A1(n60), .A2(n1033), .B1(n58), .B2(n1032), .ZN(n832) );
  INV_X1 U1669 ( .A(n454), .ZN(n455) );
  NAND2_X1 U1670 ( .A1(n789), .A2(n828), .ZN(n403) );
  AND2_X1 U1671 ( .A1(n1438), .A2(n815), .ZN(n1009) );
  INV_X1 U1672 ( .A(n9), .ZN(n815) );
  INV_X1 U1673 ( .A(n805), .ZN(n930) );
  OAI22_X1 U1674 ( .A1(n60), .A2(n1040), .B1(n1484), .B2(n1039), .ZN(n839) );
  AOI21_X1 U1675 ( .B1(n30), .B2(n28), .A(n1135), .ZN(n805) );
  OAI22_X1 U1676 ( .A1(n29), .A2(n1385), .B1(n27), .B2(n1145), .ZN(n940) );
  OAI22_X1 U1677 ( .A1(n6), .A2(n1222), .B1(n1221), .B2(n4), .ZN(n1013) );
  OAI22_X1 U1678 ( .A1(n1429), .A2(n1203), .B1(n10), .B2(n1202), .ZN(n994) );
  OAI22_X1 U1679 ( .A1(n1422), .A2(n1096), .B1(n1476), .B2(n1095), .ZN(n892)
         );
  OAI22_X1 U1680 ( .A1(n1413), .A2(n1039), .B1(n58), .B2(n1038), .ZN(n838) );
  OAI22_X1 U1681 ( .A1(n54), .A2(n1058), .B1(n52), .B2(n1057), .ZN(n856) );
  OAI22_X1 U1682 ( .A1(n48), .A2(n1076), .B1(n46), .B2(n1075), .ZN(n873) );
  OAI22_X1 U1683 ( .A1(n54), .A2(n1057), .B1(n52), .B2(n1056), .ZN(n855) );
  OAI22_X1 U1684 ( .A1(n1422), .A2(n1099), .B1(n1476), .B2(n1098), .ZN(n895)
         );
  OAI22_X1 U1685 ( .A1(n48), .A2(n1080), .B1(n46), .B2(n1079), .ZN(n877) );
  OAI22_X1 U1686 ( .A1(n1437), .A2(n1189), .B1(n15), .B2(n1188), .ZN(n981) );
  OAI22_X1 U1687 ( .A1(n47), .A2(n1088), .B1(n45), .B2(n1087), .ZN(n885) );
  AND2_X1 U1688 ( .A1(n1488), .A2(n791), .ZN(n849) );
  OAI22_X1 U1689 ( .A1(n6), .A2(n1221), .B1(n1220), .B2(n4), .ZN(n1012) );
  OAI22_X1 U1690 ( .A1(n35), .A2(n1128), .B1(n33), .B2(n1127), .ZN(n923) );
  OAI22_X1 U1691 ( .A1(n47), .A2(n1090), .B1(n1089), .B2(n45), .ZN(n887) );
  OAI22_X1 U1692 ( .A1(n12), .A2(n1204), .B1(n1203), .B2(n10), .ZN(n995) );
  OAI22_X1 U1693 ( .A1(n35), .A2(n1118), .B1(n34), .B2(n1117), .ZN(n913) );
  OAI22_X1 U1694 ( .A1(n30), .A2(n1137), .B1(n28), .B2(n1136), .ZN(n931) );
  OAI22_X1 U1695 ( .A1(n53), .A2(n1061), .B1(n51), .B2(n1060), .ZN(n859) );
  OAI22_X1 U1696 ( .A1(n1432), .A2(n1119), .B1(n34), .B2(n1118), .ZN(n914) );
  OAI22_X1 U1697 ( .A1(n30), .A2(n1138), .B1(n28), .B2(n1137), .ZN(n932) );
  OAI22_X1 U1698 ( .A1(n42), .A2(n1100), .B1(n1476), .B2(n1099), .ZN(n896) );
  OAI22_X1 U1699 ( .A1(n1432), .A2(n1132), .B1(n33), .B2(n1131), .ZN(n927) );
  OAI22_X1 U1700 ( .A1(n11), .A2(n1208), .B1(n9), .B2(n1207), .ZN(n999) );
  OAI22_X1 U1701 ( .A1(n23), .A2(n1170), .B1(n21), .B2(n1169), .ZN(n963) );
  INV_X1 U1702 ( .A(n799), .ZN(n890) );
  OAI22_X1 U1703 ( .A1(n54), .A2(n1055), .B1(n52), .B2(n1054), .ZN(n853) );
  OAI22_X1 U1704 ( .A1(n60), .A2(n1036), .B1(n58), .B2(n1035), .ZN(n835) );
  OAI22_X1 U1705 ( .A1(n1437), .A2(n1181), .B1(n16), .B2(n1180), .ZN(n973) );
  OAI22_X1 U1706 ( .A1(n24), .A2(n1162), .B1(n22), .B2(n1161), .ZN(n955) );
  OAI22_X1 U1707 ( .A1(n24), .A2(n1164), .B1(n22), .B2(n1163), .ZN(n957) );
  OAI22_X1 U1708 ( .A1(n24), .A2(n1165), .B1(n22), .B2(n1164), .ZN(n958) );
  OAI22_X1 U1709 ( .A1(n1437), .A2(n1184), .B1(n16), .B2(n1183), .ZN(n976) );
  OAI22_X1 U1710 ( .A1(n30), .A2(n1139), .B1(n28), .B2(n1138), .ZN(n933) );
  OAI22_X1 U1711 ( .A1(n24), .A2(n1158), .B1(n22), .B2(n1157), .ZN(n951) );
  OAI22_X1 U1712 ( .A1(n53), .A2(n1063), .B1(n51), .B2(n1062), .ZN(n861) );
  OAI22_X1 U1713 ( .A1(n1432), .A2(n1127), .B1(n33), .B2(n1126), .ZN(n922) );
  OAI22_X1 U1714 ( .A1(n41), .A2(n1108), .B1(n1457), .B2(n1107), .ZN(n904) );
  OAI22_X1 U1715 ( .A1(n48), .A2(n1089), .B1(n45), .B2(n1088), .ZN(n886) );
  AND2_X1 U1716 ( .A1(n1438), .A2(n800), .ZN(n909) );
  OAI22_X1 U1717 ( .A1(n29), .A2(n1151), .B1(n27), .B2(n1150), .ZN(n945) );
  OAI22_X1 U1718 ( .A1(n6), .A2(n1227), .B1(n1226), .B2(n4), .ZN(n1018) );
  OAI22_X1 U1719 ( .A1(n1432), .A2(n1121), .B1(n34), .B2(n1120), .ZN(n916) );
  OAI22_X1 U1720 ( .A1(n53), .A2(n1064), .B1(n51), .B2(n1063), .ZN(n862) );
  OAI22_X1 U1721 ( .A1(n60), .A2(n1045), .B1(n1484), .B2(n1044), .ZN(n844) );
  OAI22_X1 U1722 ( .A1(n11), .A2(n1211), .B1(n9), .B2(n1210), .ZN(n1002) );
  OAI22_X1 U1723 ( .A1(n17), .A2(n1192), .B1(n15), .B2(n1191), .ZN(n984) );
  OAI22_X1 U1724 ( .A1(n23), .A2(n1173), .B1(n21), .B2(n1172), .ZN(n966) );
  OAI22_X1 U1725 ( .A1(n1432), .A2(n1122), .B1(n34), .B2(n1121), .ZN(n917) );
  OAI22_X1 U1726 ( .A1(n29), .A2(n1150), .B1(n27), .B2(n1149), .ZN(n944) );
  OAI22_X1 U1727 ( .A1(n1432), .A2(n1131), .B1(n33), .B2(n1130), .ZN(n926) );
  OAI22_X1 U1728 ( .A1(n18), .A2(n1188), .B1(n15), .B2(n1187), .ZN(n980) );
  OAI22_X1 U1729 ( .A1(n1422), .A2(n1104), .B1(n1103), .B2(n1458), .ZN(n900)
         );
  OAI22_X1 U1730 ( .A1(n1437), .A2(n1180), .B1(n16), .B2(n1179), .ZN(n972) );
  OAI22_X1 U1731 ( .A1(n60), .A2(n1426), .B1(n1484), .B2(n1046), .ZN(n846) );
  OAI22_X1 U1732 ( .A1(n47), .A2(n1454), .B1(n45), .B2(n1086), .ZN(n884) );
  OAI22_X1 U1733 ( .A1(n30), .A2(n1144), .B1(n28), .B2(n1143), .ZN(n938) );
  OAI22_X1 U1734 ( .A1(n1068), .A2(n53), .B1(n1067), .B2(n51), .ZN(n866) );
  OAI22_X1 U1735 ( .A1(n1422), .A2(n1103), .B1(n1457), .B2(n1102), .ZN(n899)
         );
  OAI22_X1 U1736 ( .A1(n30), .A2(n1141), .B1(n28), .B2(n1140), .ZN(n935) );
  OAI22_X1 U1737 ( .A1(n48), .A2(n1084), .B1(n45), .B2(n1083), .ZN(n881) );
  OAI22_X1 U1738 ( .A1(n41), .A2(n1098), .B1(n1476), .B2(n1097), .ZN(n894) );
  OAI22_X1 U1739 ( .A1(n36), .A2(n1117), .B1(n34), .B2(n1116), .ZN(n912) );
  OAI22_X1 U1740 ( .A1(n48), .A2(n1079), .B1(n46), .B2(n1078), .ZN(n876) );
  OAI22_X1 U1741 ( .A1(n18), .A2(n1187), .B1(n15), .B2(n1186), .ZN(n979) );
  OAI22_X1 U1742 ( .A1(n23), .A2(n1168), .B1(n21), .B2(n1167), .ZN(n961) );
  OAI22_X1 U1743 ( .A1(n1124), .A2(n35), .B1(n1123), .B2(n33), .ZN(n919) );
  INV_X1 U1744 ( .A(n817), .ZN(n1010) );
  OAI22_X1 U1745 ( .A1(n1048), .A2(n1413), .B1(n1047), .B2(n1484), .ZN(n847)
         );
  OAI22_X1 U1746 ( .A1(n41), .A2(n1095), .B1(n1476), .B2(n1094), .ZN(n891) );
  INV_X1 U1747 ( .A(n802), .ZN(n910) );
  OAI22_X1 U1748 ( .A1(n60), .A2(n1038), .B1(n58), .B2(n1037), .ZN(n837) );
  INV_X1 U1749 ( .A(n464), .ZN(n465) );
  OAI22_X1 U1750 ( .A1(n1413), .A2(n1035), .B1(n58), .B2(n1034), .ZN(n834) );
  OAI22_X1 U1751 ( .A1(n54), .A2(n1054), .B1(n52), .B2(n1053), .ZN(n852) );
  INV_X1 U1752 ( .A(n796), .ZN(n870) );
  OAI22_X1 U1753 ( .A1(n54), .A2(n1053), .B1(n52), .B2(n1052), .ZN(n851) );
  AOI21_X1 U1754 ( .B1(n1439), .B2(n46), .A(n1072), .ZN(n796) );
  OAI22_X1 U1755 ( .A1(n11), .A2(n1212), .B1(n9), .B2(n1211), .ZN(n1003) );
  OAI22_X1 U1756 ( .A1(n23), .A2(n1174), .B1(n21), .B2(n1173), .ZN(n967) );
  OAI22_X1 U1757 ( .A1(n5), .A2(n1232), .B1(n1231), .B2(n3), .ZN(n1023) );
  OAI22_X1 U1758 ( .A1(n11), .A2(n1213), .B1(n9), .B2(n1212), .ZN(n1004) );
  OAI22_X1 U1759 ( .A1(n17), .A2(n1194), .B1(n15), .B2(n1193), .ZN(n986) );
  OAI22_X1 U1760 ( .A1(n48), .A2(n1081), .B1(n46), .B2(n1080), .ZN(n878) );
  OAI22_X1 U1761 ( .A1(n53), .A2(n1062), .B1(n51), .B2(n1061), .ZN(n860) );
  OAI22_X1 U1762 ( .A1(n60), .A2(n1043), .B1(n1484), .B2(n1042), .ZN(n842) );
  AND2_X1 U1763 ( .A1(n1487), .A2(n809), .ZN(n969) );
  OAI22_X1 U1764 ( .A1(n5), .A2(n1233), .B1(n1232), .B2(n3), .ZN(n1024) );
  OAI22_X1 U1765 ( .A1(n1429), .A2(n1214), .B1(n9), .B2(n1213), .ZN(n1005) );
  OAI22_X1 U1766 ( .A1(n1429), .A2(n1205), .B1(n10), .B2(n1204), .ZN(n996) );
  OAI22_X1 U1767 ( .A1(n5), .A2(n1230), .B1(n1229), .B2(n3), .ZN(n1021) );
  OAI22_X1 U1768 ( .A1(n1439), .A2(n1074), .B1(n46), .B2(n1073), .ZN(n871) );
  OAI22_X1 U1769 ( .A1(n29), .A2(n1147), .B1(n27), .B2(n1146), .ZN(n941) );
  OAI22_X1 U1770 ( .A1(n23), .A2(n1166), .B1(n21), .B2(n1165), .ZN(n959) );
  OAI22_X1 U1771 ( .A1(n18), .A2(n1185), .B1(n16), .B2(n1184), .ZN(n977) );
  OAI22_X1 U1772 ( .A1(n1422), .A2(n1101), .B1(n1476), .B2(n1100), .ZN(n897)
         );
  OAI22_X1 U1773 ( .A1(n48), .A2(n1082), .B1(n45), .B2(n1081), .ZN(n879) );
  OAI22_X1 U1774 ( .A1(n36), .A2(n1120), .B1(n34), .B2(n1119), .ZN(n915) );
  AND2_X1 U1775 ( .A1(n1438), .A2(n797), .ZN(n889) );
  OAI22_X1 U1776 ( .A1(n35), .A2(n1130), .B1(n33), .B2(n1129), .ZN(n925) );
  OAI22_X1 U1777 ( .A1(n6), .A2(n1225), .B1(n1224), .B2(n4), .ZN(n1016) );
  AND2_X1 U1778 ( .A1(n1487), .A2(n803), .ZN(n929) );
  OAI22_X1 U1779 ( .A1(n5), .A2(n1229), .B1(n1228), .B2(n3), .ZN(n1020) );
  OAI22_X1 U1780 ( .A1(n23), .A2(n1172), .B1(n21), .B2(n1171), .ZN(n965) );
  OAI22_X1 U1781 ( .A1(n29), .A2(n1152), .B1(n27), .B2(n1151), .ZN(n946) );
  OAI22_X1 U1782 ( .A1(n6), .A2(n1228), .B1(n1227), .B2(n4), .ZN(n1019) );
  OAI22_X1 U1783 ( .A1(n17), .A2(n1190), .B1(n15), .B2(n1189), .ZN(n982) );
  OAI22_X1 U1784 ( .A1(n6), .A2(n1226), .B1(n1225), .B2(n4), .ZN(n1017) );
  OAI22_X1 U1785 ( .A1(n1429), .A2(n1207), .B1(n10), .B2(n1206), .ZN(n998) );
  OAI22_X1 U1786 ( .A1(n23), .A2(n1169), .B1(n21), .B2(n1168), .ZN(n962) );
  OAI22_X1 U1787 ( .A1(n1439), .A2(n1077), .B1(n46), .B2(n1076), .ZN(n874) );
  INV_X1 U1788 ( .A(n496), .ZN(n497) );
  OAI22_X1 U1789 ( .A1(n1439), .A2(n1078), .B1(n46), .B2(n1077), .ZN(n875) );
  OAI22_X1 U1790 ( .A1(n36), .A2(n1116), .B1(n34), .B2(n1115), .ZN(n911) );
  OAI22_X1 U1791 ( .A1(n54), .A2(n1059), .B1(n52), .B2(n1058), .ZN(n857) );
  OAI22_X1 U1792 ( .A1(n59), .A2(n1042), .B1(n1484), .B2(n1041), .ZN(n841) );
  INV_X1 U1793 ( .A(n808), .ZN(n950) );
  AOI21_X1 U1794 ( .B1(n24), .B2(n22), .A(n1156), .ZN(n808) );
  OAI22_X1 U1795 ( .A1(n1422), .A2(n1102), .B1(n1476), .B2(n1101), .ZN(n898)
         );
  INV_X1 U1796 ( .A(n574), .ZN(n575) );
  AND2_X1 U1797 ( .A1(n1438), .A2(n806), .ZN(n949) );
  OAI22_X1 U1798 ( .A1(n5), .A2(n1231), .B1(n1230), .B2(n3), .ZN(n1022) );
  OAI22_X1 U1799 ( .A1(n18), .A2(n1193), .B1(n15), .B2(n1192), .ZN(n985) );
  OAI22_X1 U1800 ( .A1(n1437), .A2(n1430), .B1(n1178), .B2(n16), .ZN(n971) );
  OAI22_X1 U1801 ( .A1(n59), .A2(n1046), .B1(n1045), .B2(n1484), .ZN(n845) );
  INV_X1 U1802 ( .A(n814), .ZN(n990) );
  OAI22_X1 U1803 ( .A1(n47), .A2(n1085), .B1(n45), .B2(n1084), .ZN(n882) );
  OAI22_X1 U1804 ( .A1(n24), .A2(n1161), .B1(n22), .B2(n1160), .ZN(n954) );
  OAI22_X1 U1805 ( .A1(n53), .A2(n1066), .B1(n51), .B2(n1065), .ZN(n864) );
  OAI22_X1 U1806 ( .A1(n41), .A2(n1107), .B1(n1457), .B2(n1106), .ZN(n903) );
  OAI22_X1 U1807 ( .A1(n11), .A2(n1202), .B1(n10), .B2(n1201), .ZN(n993) );
  OAI22_X1 U1808 ( .A1(n53), .A2(n1069), .B1(n51), .B2(n1068), .ZN(n867) );
  OAI22_X1 U1809 ( .A1(n1422), .A2(n1097), .B1(n1476), .B2(n1096), .ZN(n893)
         );
  OAI22_X1 U1810 ( .A1(n1422), .A2(n1106), .B1(n1458), .B2(n1105), .ZN(n902)
         );
  OAI22_X1 U1811 ( .A1(n6), .A2(n1220), .B1(n1441), .B2(n4), .ZN(n1011) );
  OAI22_X1 U1812 ( .A1(n24), .A2(n1163), .B1(n22), .B2(n1162), .ZN(n956) );
  OAI22_X1 U1813 ( .A1(n1439), .A2(n1075), .B1(n46), .B2(n1074), .ZN(n872) );
  OAI22_X1 U1814 ( .A1(n1413), .A2(n1037), .B1(n58), .B2(n1036), .ZN(n836) );
  OAI22_X1 U1815 ( .A1(n54), .A2(n1056), .B1(n52), .B2(n1055), .ZN(n854) );
  INV_X1 U1816 ( .A(n518), .ZN(n519) );
  OAI22_X1 U1817 ( .A1(n54), .A2(n1060), .B1(n52), .B2(n1059), .ZN(n858) );
  OAI22_X1 U1818 ( .A1(n1413), .A2(n1041), .B1(n1484), .B2(n1040), .ZN(n840)
         );
  OAI22_X1 U1819 ( .A1(n1429), .A2(n1209), .B1(n9), .B2(n1208), .ZN(n1000) );
  OAI22_X1 U1820 ( .A1(n23), .A2(n1171), .B1(n21), .B2(n1170), .ZN(n964) );
  NAND2_X1 U1821 ( .A1(n787), .A2(n788), .ZN(n400) );
  OAI22_X1 U1822 ( .A1(n42), .A2(n1293), .B1(n1113), .B2(n1456), .ZN(n823) );
  OAI22_X1 U1823 ( .A1(n42), .A2(n1112), .B1(n1111), .B2(n1457), .ZN(n908) );
  OR2_X1 U1824 ( .A1(n1488), .A2(n1293), .ZN(n1113) );
  INV_X1 U1825 ( .A(n790), .ZN(n830) );
  AOI21_X1 U1826 ( .B1(n60), .B2(n58), .A(n1030), .ZN(n790) );
  OAI22_X1 U1827 ( .A1(n1432), .A2(n1123), .B1(n34), .B2(n1122), .ZN(n918) );
  OAI22_X1 U1828 ( .A1(n30), .A2(n1142), .B1(n28), .B2(n1141), .ZN(n936) );
  INV_X1 U1829 ( .A(n608), .ZN(n609) );
  INV_X1 U1830 ( .A(n27), .ZN(n806) );
  OR2_X1 U1831 ( .A1(n1488), .A2(n1423), .ZN(n1050) );
  OR2_X1 U1832 ( .A1(n1438), .A2(n1297), .ZN(n1197) );
  OR2_X1 U1833 ( .A1(n1438), .A2(n1292), .ZN(n1092) );
  OAI22_X1 U1834 ( .A1(n1413), .A2(n1044), .B1(n1484), .B2(n1043), .ZN(n843)
         );
  INV_X1 U1835 ( .A(n811), .ZN(n970) );
  AOI21_X1 U1836 ( .B1(n17), .B2(n16), .A(n1177), .ZN(n811) );
  INV_X1 U1837 ( .A(n15), .ZN(n812) );
  INV_X1 U1838 ( .A(n51), .ZN(n794) );
  INV_X1 U1839 ( .A(n1456), .ZN(n800) );
  INV_X1 U1840 ( .A(n33), .ZN(n803) );
  INV_X1 U1841 ( .A(n1484), .ZN(n791) );
  INV_X1 U1842 ( .A(n21), .ZN(n809) );
  INV_X1 U1843 ( .A(n45), .ZN(n797) );
  AND2_X1 U1844 ( .A1(n1488), .A2(a[0]), .ZN(product[0]) );
  OAI22_X1 U1845 ( .A1(n5), .A2(n1236), .B1(n1235), .B2(n3), .ZN(n1027) );
  OAI22_X1 U1846 ( .A1(n11), .A2(n1217), .B1(n9), .B2(n1216), .ZN(n1008) );
  XNOR2_X1 U1847 ( .A(n7), .B(n1487), .ZN(n1217) );
  OAI22_X1 U1848 ( .A1(n11), .A2(n1298), .B1(n1218), .B2(n10), .ZN(n828) );
  OR2_X1 U1849 ( .A1(n1487), .A2(n1298), .ZN(n1218) );
  INV_X1 U1850 ( .A(n7), .ZN(n1298) );
  OAI22_X1 U1851 ( .A1(n6), .A2(n1299), .B1(n1239), .B2(n4), .ZN(n829) );
  OR2_X1 U1852 ( .A1(n1438), .A2(n1299), .ZN(n1239) );
  INV_X1 U1853 ( .A(n1), .ZN(n1299) );
  OAI22_X1 U1854 ( .A1(n5), .A2(n1238), .B1(n1237), .B2(n3), .ZN(n1029) );
  OAI22_X1 U1855 ( .A1(n47), .A2(n1091), .B1(n45), .B2(n1090), .ZN(n888) );
  OAI22_X1 U1856 ( .A1(n48), .A2(n1292), .B1(n1092), .B2(n46), .ZN(n822) );
  XNOR2_X1 U1857 ( .A(n1460), .B(n1493), .ZN(n1091) );
  BUF_X1 U1858 ( .A(n61), .Z(n1493) );
  OAI22_X1 U1859 ( .A1(n53), .A2(n1070), .B1(n51), .B2(n1069), .ZN(n868) );
  XNOR2_X1 U1860 ( .A(n49), .B(n1487), .ZN(n1070) );
  OAI22_X1 U1861 ( .A1(n17), .A2(n1196), .B1(n15), .B2(n1195), .ZN(n988) );
  OAI22_X1 U1862 ( .A1(n17), .A2(n1297), .B1(n1197), .B2(n16), .ZN(n827) );
  XNOR2_X1 U1863 ( .A(n1440), .B(n1494), .ZN(n1196) );
  XNOR2_X1 U1864 ( .A(n13), .B(n1249), .ZN(n1186) );
  XNOR2_X1 U1865 ( .A(n13), .B(n1248), .ZN(n1185) );
  XNOR2_X1 U1866 ( .A(n1440), .B(n1475), .ZN(n1193) );
  XNOR2_X1 U1867 ( .A(n13), .B(n1250), .ZN(n1187) );
  XNOR2_X1 U1868 ( .A(n13), .B(n1255), .ZN(n1192) );
  XNOR2_X1 U1869 ( .A(n13), .B(n1243), .ZN(n1180) );
  XNOR2_X1 U1870 ( .A(n13), .B(n1251), .ZN(n1188) );
  XNOR2_X1 U1871 ( .A(n13), .B(n1241), .ZN(n1178) );
  XNOR2_X1 U1872 ( .A(n13), .B(n1254), .ZN(n1191) );
  XNOR2_X1 U1873 ( .A(n13), .B(n1244), .ZN(n1181) );
  XNOR2_X1 U1874 ( .A(n13), .B(n1245), .ZN(n1182) );
  XNOR2_X1 U1875 ( .A(n13), .B(n1247), .ZN(n1184) );
  XNOR2_X1 U1876 ( .A(n13), .B(n1252), .ZN(n1189) );
  XNOR2_X1 U1877 ( .A(n1440), .B(n1257), .ZN(n1194) );
  XNOR2_X1 U1878 ( .A(n13), .B(n1246), .ZN(n1183) );
  XNOR2_X1 U1879 ( .A(n13), .B(n1242), .ZN(n1179) );
  XNOR2_X1 U1880 ( .A(n13), .B(n1253), .ZN(n1190) );
  XNOR2_X1 U1881 ( .A(n13), .B(n1258), .ZN(n1195) );
  XNOR2_X1 U1882 ( .A(n7), .B(n1257), .ZN(n1215) );
  XNOR2_X1 U1883 ( .A(n7), .B(n1256), .ZN(n1214) );
  XNOR2_X1 U1884 ( .A(n49), .B(n1258), .ZN(n1069) );
  XNOR2_X1 U1885 ( .A(n7), .B(n1247), .ZN(n1205) );
  XNOR2_X1 U1886 ( .A(n7), .B(n1246), .ZN(n1204) );
  XNOR2_X1 U1887 ( .A(n43), .B(n1258), .ZN(n1090) );
  XNOR2_X1 U1888 ( .A(n7), .B(n1253), .ZN(n1211) );
  XNOR2_X1 U1889 ( .A(n55), .B(n1254), .ZN(n1044) );
  XNOR2_X1 U1890 ( .A(n7), .B(n1254), .ZN(n1212) );
  XNOR2_X1 U1891 ( .A(n55), .B(n1253), .ZN(n1043) );
  XNOR2_X1 U1892 ( .A(n43), .B(n1257), .ZN(n1089) );
  XNOR2_X1 U1893 ( .A(n7), .B(n1245), .ZN(n1203) );
  XNOR2_X1 U1894 ( .A(n49), .B(n1252), .ZN(n1063) );
  XNOR2_X1 U1895 ( .A(n1436), .B(n1241), .ZN(n1052) );
  XNOR2_X1 U1896 ( .A(n49), .B(n1255), .ZN(n1066) );
  XNOR2_X1 U1897 ( .A(n55), .B(n1252), .ZN(n1042) );
  XNOR2_X1 U1898 ( .A(n1460), .B(n1248), .ZN(n1080) );
  XNOR2_X1 U1899 ( .A(n49), .B(n1253), .ZN(n1064) );
  XNOR2_X1 U1900 ( .A(n49), .B(n1251), .ZN(n1062) );
  XNOR2_X1 U1901 ( .A(n49), .B(n1254), .ZN(n1065) );
  XNOR2_X1 U1902 ( .A(n7), .B(n1248), .ZN(n1206) );
  XNOR2_X1 U1903 ( .A(n1460), .B(n1250), .ZN(n1082) );
  XNOR2_X1 U1904 ( .A(n1424), .B(n1243), .ZN(n1033) );
  XNOR2_X1 U1905 ( .A(n1256), .B(n43), .ZN(n1088) );
  XNOR2_X1 U1906 ( .A(n49), .B(n1256), .ZN(n1067) );
  XNOR2_X1 U1907 ( .A(n7), .B(n1244), .ZN(n1202) );
  XNOR2_X1 U1908 ( .A(n1460), .B(n1244), .ZN(n1076) );
  XNOR2_X1 U1909 ( .A(n49), .B(n1250), .ZN(n1061) );
  XNOR2_X1 U1910 ( .A(n1251), .B(n55), .ZN(n1041) );
  XNOR2_X1 U1911 ( .A(n1424), .B(n1242), .ZN(n1032) );
  XNOR2_X1 U1912 ( .A(n7), .B(n1255), .ZN(n1213) );
  XNOR2_X1 U1913 ( .A(n1460), .B(n1251), .ZN(n1083) );
  XNOR2_X1 U1914 ( .A(n1460), .B(n1247), .ZN(n1079) );
  XNOR2_X1 U1915 ( .A(n1460), .B(n1249), .ZN(n1081) );
  XNOR2_X1 U1916 ( .A(n1257), .B(n55), .ZN(n1047) );
  XNOR2_X1 U1917 ( .A(n1460), .B(n1245), .ZN(n1077) );
  XNOR2_X1 U1918 ( .A(n49), .B(n1249), .ZN(n1060) );
  XNOR2_X1 U1919 ( .A(n7), .B(n1252), .ZN(n1210) );
  XNOR2_X1 U1920 ( .A(n1460), .B(n1252), .ZN(n1084) );
  XNOR2_X1 U1921 ( .A(n55), .B(n1258), .ZN(n1048) );
  XNOR2_X1 U1922 ( .A(n43), .B(n1255), .ZN(n1087) );
  XNOR2_X1 U1923 ( .A(n55), .B(n1255), .ZN(n1045) );
  XNOR2_X1 U1924 ( .A(n1460), .B(n1253), .ZN(n1085) );
  XNOR2_X1 U1925 ( .A(n7), .B(n1249), .ZN(n1207) );
  XNOR2_X1 U1926 ( .A(n1460), .B(n1242), .ZN(n1074) );
  XNOR2_X1 U1927 ( .A(n1424), .B(n1244), .ZN(n1034) );
  XNOR2_X1 U1928 ( .A(n1460), .B(n1241), .ZN(n1073) );
  XNOR2_X1 U1929 ( .A(n49), .B(n1257), .ZN(n1068) );
  XNOR2_X1 U1930 ( .A(n7), .B(n1241), .ZN(n1199) );
  XNOR2_X1 U1931 ( .A(n7), .B(n1242), .ZN(n1200) );
  XNOR2_X1 U1932 ( .A(n55), .B(n1248), .ZN(n1038) );
  XNOR2_X1 U1933 ( .A(n49), .B(n1246), .ZN(n1057) );
  XNOR2_X1 U1934 ( .A(n43), .B(n1254), .ZN(n1086) );
  XNOR2_X1 U1935 ( .A(n1424), .B(n1241), .ZN(n1031) );
  XNOR2_X1 U1936 ( .A(n49), .B(n1245), .ZN(n1056) );
  XNOR2_X1 U1937 ( .A(n55), .B(n1247), .ZN(n1037) );
  XNOR2_X1 U1938 ( .A(n7), .B(n1243), .ZN(n1201) );
  XNOR2_X1 U1939 ( .A(n1250), .B(n55), .ZN(n1040) );
  XNOR2_X1 U1940 ( .A(n1460), .B(n1243), .ZN(n1075) );
  XNOR2_X1 U1941 ( .A(n1436), .B(n1244), .ZN(n1055) );
  XNOR2_X1 U1942 ( .A(n1424), .B(n1246), .ZN(n1036) );
  XNOR2_X1 U1943 ( .A(n49), .B(n1248), .ZN(n1059) );
  XNOR2_X1 U1944 ( .A(n1436), .B(n1247), .ZN(n1058) );
  XNOR2_X1 U1945 ( .A(n1424), .B(n1249), .ZN(n1039) );
  XNOR2_X1 U1946 ( .A(n1436), .B(n1242), .ZN(n1053) );
  XNOR2_X1 U1947 ( .A(n1436), .B(n1243), .ZN(n1054) );
  XNOR2_X1 U1948 ( .A(n1424), .B(n1245), .ZN(n1035) );
  XNOR2_X1 U1949 ( .A(n1460), .B(n1246), .ZN(n1078) );
  XNOR2_X1 U1950 ( .A(n7), .B(n1250), .ZN(n1208) );
  XNOR2_X1 U1951 ( .A(n1256), .B(n55), .ZN(n1046) );
  XNOR2_X1 U1952 ( .A(n7), .B(n1251), .ZN(n1209) );
  XNOR2_X1 U1953 ( .A(n7), .B(n1258), .ZN(n1216) );
  XNOR2_X1 U1954 ( .A(n1240), .B(n13), .ZN(n1177) );
  XNOR2_X1 U1955 ( .A(n7), .B(n1240), .ZN(n1198) );
  XNOR2_X1 U1956 ( .A(n1460), .B(n1434), .ZN(n1072) );
  XNOR2_X1 U1957 ( .A(n1436), .B(n1434), .ZN(n1051) );
  XNOR2_X1 U1958 ( .A(n1424), .B(n1434), .ZN(n1030) );
  BUF_X2 U1959 ( .A(n1284), .Z(n34) );
  BUF_X2 U1960 ( .A(n1285), .Z(n28) );
  BUF_X1 U1961 ( .A(n1280), .Z(n58) );
  BUF_X1 U1962 ( .A(n1282), .Z(n46) );
  BUF_X2 U1963 ( .A(n1275), .Z(n30) );
  BUF_X2 U1964 ( .A(n1431), .Z(n52) );
  BUF_X1 U1965 ( .A(n1279), .Z(n5) );
  OAI22_X1 U1966 ( .A1(n1413), .A2(n1049), .B1(n1484), .B2(n1425), .ZN(n848)
         );
  OAI22_X1 U1967 ( .A1(n1413), .A2(n1423), .B1(n1050), .B2(n58), .ZN(n820) );
  XNOR2_X1 U1968 ( .A(n55), .B(n1494), .ZN(n1049) );
  INV_X1 U1969 ( .A(n25), .ZN(n1295) );
  INV_X1 U1970 ( .A(n31), .ZN(n1294) );
  BUF_X2 U1971 ( .A(n1271), .Z(n54) );
  BUF_X2 U1972 ( .A(n1271), .Z(n53) );
  INV_X1 U1973 ( .A(n13), .ZN(n1297) );
  INV_X1 U1974 ( .A(n43), .ZN(n1292) );
  BUF_X1 U1975 ( .A(n1289), .Z(n3) );
  BUF_X1 U1976 ( .A(n1289), .Z(n4) );
  INV_X1 U1977 ( .A(n49), .ZN(n1291) );
  BUF_X2 U1978 ( .A(n1276), .Z(n24) );
  INV_X1 U1979 ( .A(n37), .ZN(n1293) );
  INV_X1 U1980 ( .A(n19), .ZN(n1296) );
  BUF_X1 U1981 ( .A(n1277), .Z(n17) );
  BUF_X2 U1982 ( .A(n1278), .Z(n11) );
  XNOR2_X1 U1983 ( .A(a[6]), .B(a[5]), .ZN(n1286) );
  XNOR2_X1 U1984 ( .A(a[17]), .B(a[18]), .ZN(n1280) );
  BUF_X4 U1985 ( .A(a[19]), .Z(n55) );
  XNOR2_X1 U1986 ( .A(a[13]), .B(a[14]), .ZN(n1282) );
  CLKBUF_X3 U1987 ( .A(b[5]), .Z(n1254) );
  CLKBUF_X3 U1988 ( .A(b[8]), .Z(n1251) );
  CLKBUF_X3 U1989 ( .A(b[9]), .Z(n1250) );
  BUF_X4 U1990 ( .A(a[13]), .Z(n37) );
  BUF_X4 U1991 ( .A(a[7]), .Z(n19) );
  NAND2_X1 U1992 ( .A1(n1269), .A2(n1289), .ZN(n1279) );
  XNOR2_X1 U1993 ( .A(a[4]), .B(a[3]), .ZN(n1287) );
  AOI21_X1 U1994 ( .B1(n63), .B2(n182), .A(n183), .ZN(n181) );
  INV_X1 U1995 ( .A(n1481), .ZN(n426) );
  OAI21_X1 U1996 ( .B1(n296), .B2(n304), .A(n297), .ZN(n295) );
  AOI21_X1 U1997 ( .B1(n63), .B2(n169), .A(n170), .ZN(n168) );
  BUF_X2 U1998 ( .A(n291), .Z(n63) );
  NOR2_X1 U1999 ( .A1(n247), .A2(n117), .ZN(n115) );
  NOR2_X1 U2000 ( .A1(n247), .A2(n108), .ZN(n106) );
  NOR2_X1 U2001 ( .A1(n247), .A2(n160), .ZN(n158) );
  NOR2_X1 U2002 ( .A1(n247), .A2(n130), .ZN(n128) );
  NOR2_X1 U2003 ( .A1(n247), .A2(n145), .ZN(n143) );
  NOR2_X1 U2004 ( .A1(n247), .A2(n184), .ZN(n182) );
  NOR2_X1 U2005 ( .A1(n247), .A2(n225), .ZN(n223) );
  NOR2_X1 U2006 ( .A1(n247), .A2(n216), .ZN(n210) );
  INV_X1 U2007 ( .A(n247), .ZN(n245) );
  NOR2_X1 U2008 ( .A1(n247), .A2(n171), .ZN(n169) );
  NOR2_X1 U2009 ( .A1(n247), .A2(n242), .ZN(n232) );
  XNOR2_X1 U2010 ( .A(n1428), .B(n1248), .ZN(n1164) );
  XNOR2_X1 U2011 ( .A(n1428), .B(n1494), .ZN(n1175) );
  XNOR2_X1 U2012 ( .A(n19), .B(n1254), .ZN(n1170) );
  XNOR2_X1 U2013 ( .A(n19), .B(n1249), .ZN(n1165) );
  XNOR2_X1 U2014 ( .A(n19), .B(n1258), .ZN(n1174) );
  XNOR2_X1 U2015 ( .A(n19), .B(n1253), .ZN(n1169) );
  XNOR2_X1 U2016 ( .A(n1257), .B(n19), .ZN(n1173) );
  XNOR2_X1 U2017 ( .A(n19), .B(n1252), .ZN(n1168) );
  XNOR2_X1 U2018 ( .A(n19), .B(n1243), .ZN(n1159) );
  XNOR2_X1 U2019 ( .A(n19), .B(n1256), .ZN(n1172) );
  XNOR2_X1 U2020 ( .A(n19), .B(n1247), .ZN(n1163) );
  XNOR2_X1 U2021 ( .A(n19), .B(n1246), .ZN(n1162) );
  XNOR2_X1 U2022 ( .A(n19), .B(n1242), .ZN(n1158) );
  XNOR2_X1 U2023 ( .A(n19), .B(n1255), .ZN(n1171) );
  XNOR2_X1 U2024 ( .A(n19), .B(n1251), .ZN(n1167) );
  XNOR2_X1 U2025 ( .A(n19), .B(n1250), .ZN(n1166) );
  XNOR2_X1 U2026 ( .A(n19), .B(n1241), .ZN(n1157) );
  XNOR2_X1 U2027 ( .A(n19), .B(n1245), .ZN(n1161) );
  XNOR2_X1 U2028 ( .A(n19), .B(n1244), .ZN(n1160) );
  XNOR2_X1 U2029 ( .A(n19), .B(n1240), .ZN(n1156) );
  AOI21_X1 U2030 ( .B1(n349), .B2(n1469), .A(n344), .ZN(n342) );
  NAND2_X1 U2031 ( .A1(n693), .A2(n706), .ZN(n346) );
  XOR2_X1 U2032 ( .A(n314), .B(n85), .Z(product[20]) );
  INV_X1 U2033 ( .A(n338), .ZN(n336) );
  AOI21_X1 U2034 ( .B1(n64), .B2(n210), .A(n211), .ZN(n209) );
  CLKBUF_X3 U2035 ( .A(n1285), .Z(n27) );
  NAND2_X1 U2036 ( .A1(n1265), .A2(n1285), .ZN(n1275) );
  XNOR2_X1 U2037 ( .A(n385), .B(n97), .ZN(product[8]) );
  XOR2_X1 U2038 ( .A(n198), .B(n73), .Z(product[32]) );
  XNOR2_X1 U2039 ( .A(n25), .B(n1250), .ZN(n1145) );
  XNOR2_X1 U2040 ( .A(n25), .B(n1246), .ZN(n1141) );
  XNOR2_X1 U2041 ( .A(n25), .B(n1494), .ZN(n1154) );
  XNOR2_X1 U2042 ( .A(n25), .B(n1245), .ZN(n1140) );
  XNOR2_X1 U2043 ( .A(n25), .B(n1254), .ZN(n1149) );
  XNOR2_X1 U2044 ( .A(n25), .B(n1251), .ZN(n1146) );
  XNOR2_X1 U2045 ( .A(n25), .B(n1255), .ZN(n1150) );
  XNOR2_X1 U2046 ( .A(n25), .B(n1247), .ZN(n1142) );
  XNOR2_X1 U2047 ( .A(n25), .B(n1258), .ZN(n1153) );
  XNOR2_X1 U2048 ( .A(n25), .B(n1244), .ZN(n1139) );
  XNOR2_X1 U2049 ( .A(n25), .B(n1257), .ZN(n1152) );
  XNOR2_X1 U2050 ( .A(n25), .B(n1256), .ZN(n1151) );
  XNOR2_X1 U2051 ( .A(n25), .B(n1253), .ZN(n1148) );
  XNOR2_X1 U2052 ( .A(n25), .B(n1249), .ZN(n1144) );
  XNOR2_X1 U2053 ( .A(n25), .B(n1248), .ZN(n1143) );
  XNOR2_X1 U2054 ( .A(n25), .B(n1252), .ZN(n1147) );
  XNOR2_X1 U2055 ( .A(n25), .B(n1243), .ZN(n1138) );
  XNOR2_X1 U2056 ( .A(n25), .B(n1242), .ZN(n1137) );
  XNOR2_X1 U2057 ( .A(n25), .B(n1241), .ZN(n1136) );
  XNOR2_X1 U2058 ( .A(n25), .B(n1240), .ZN(n1135) );
  XNOR2_X1 U2059 ( .A(a[10]), .B(a[9]), .ZN(n1284) );
  BUF_X4 U2060 ( .A(a[9]), .Z(n25) );
  NAND2_X1 U2061 ( .A1(n119), .A2(n1393), .ZN(n108) );
  OAI22_X1 U2062 ( .A1(n54), .A2(n1291), .B1(n1071), .B2(n52), .ZN(n821) );
  OR2_X1 U2063 ( .A1(n1438), .A2(n1291), .ZN(n1071) );
  XOR2_X1 U2064 ( .A(n181), .B(n72), .Z(product[33]) );
  AOI21_X1 U2065 ( .B1(n357), .B2(n348), .A(n349), .ZN(n347) );
  NAND2_X1 U2066 ( .A1(n348), .A2(n1469), .ZN(n341) );
  XNOR2_X1 U2067 ( .A(n31), .B(n1248), .ZN(n1122) );
  XNOR2_X1 U2068 ( .A(n31), .B(n1252), .ZN(n1126) );
  XNOR2_X1 U2069 ( .A(n31), .B(n1251), .ZN(n1125) );
  XNOR2_X1 U2070 ( .A(n31), .B(n1247), .ZN(n1121) );
  XNOR2_X1 U2071 ( .A(n31), .B(n1494), .ZN(n1133) );
  XNOR2_X1 U2072 ( .A(n31), .B(n1257), .ZN(n1131) );
  XNOR2_X1 U2073 ( .A(n31), .B(n1254), .ZN(n1128) );
  XNOR2_X1 U2074 ( .A(n31), .B(n1258), .ZN(n1132) );
  XNOR2_X1 U2075 ( .A(n31), .B(n1246), .ZN(n1120) );
  XNOR2_X1 U2076 ( .A(n31), .B(n1245), .ZN(n1119) );
  XNOR2_X1 U2077 ( .A(n1250), .B(n31), .ZN(n1124) );
  XNOR2_X1 U2078 ( .A(n31), .B(n1249), .ZN(n1123) );
  XNOR2_X1 U2079 ( .A(n31), .B(n1256), .ZN(n1130) );
  XNOR2_X1 U2080 ( .A(n31), .B(n1253), .ZN(n1127) );
  XNOR2_X1 U2081 ( .A(n31), .B(n1244), .ZN(n1118) );
  XNOR2_X1 U2082 ( .A(n31), .B(n1243), .ZN(n1117) );
  XNOR2_X1 U2083 ( .A(n31), .B(n1242), .ZN(n1116) );
  XNOR2_X1 U2084 ( .A(n31), .B(n1255), .ZN(n1129) );
  XNOR2_X1 U2085 ( .A(n31), .B(n1241), .ZN(n1115) );
  XNOR2_X1 U2086 ( .A(n31), .B(n1240), .ZN(n1114) );
  BUF_X4 U2087 ( .A(a[11]), .Z(n31) );
  NOR2_X1 U2088 ( .A1(n303), .A2(n1481), .ZN(n294) );
  NOR2_X1 U2089 ( .A1(n312), .A2(n317), .ZN(n310) );
  NAND2_X1 U2090 ( .A1(n294), .A2(n310), .ZN(n292) );
  INV_X1 U2091 ( .A(n1427), .ZN(n315) );
  XNOR2_X1 U2092 ( .A(n37), .B(n1243), .ZN(n1096) );
  XNOR2_X1 U2093 ( .A(n37), .B(n1242), .ZN(n1095) );
  XNOR2_X1 U2094 ( .A(n37), .B(n1248), .ZN(n1101) );
  XNOR2_X1 U2095 ( .A(n37), .B(n1254), .ZN(n1107) );
  XNOR2_X1 U2096 ( .A(n37), .B(n1247), .ZN(n1100) );
  XNOR2_X1 U2097 ( .A(n37), .B(n1253), .ZN(n1106) );
  XNOR2_X1 U2098 ( .A(n37), .B(n1249), .ZN(n1102) );
  XNOR2_X1 U2099 ( .A(n37), .B(n1245), .ZN(n1098) );
  XNOR2_X1 U2100 ( .A(n37), .B(n1244), .ZN(n1097) );
  XNOR2_X1 U2101 ( .A(n37), .B(n1246), .ZN(n1099) );
  XNOR2_X1 U2102 ( .A(n37), .B(n1252), .ZN(n1105) );
  XNOR2_X1 U2103 ( .A(n37), .B(n1257), .ZN(n1110) );
  XNOR2_X1 U2104 ( .A(n37), .B(n1251), .ZN(n1104) );
  XNOR2_X1 U2105 ( .A(n37), .B(n1250), .ZN(n1103) );
  XNOR2_X1 U2106 ( .A(n37), .B(n1493), .ZN(n1112) );
  XNOR2_X1 U2107 ( .A(n37), .B(n1256), .ZN(n1109) );
  XNOR2_X1 U2108 ( .A(n37), .B(n1255), .ZN(n1108) );
  XNOR2_X1 U2109 ( .A(n37), .B(n1258), .ZN(n1111) );
  XNOR2_X1 U2110 ( .A(n37), .B(n1241), .ZN(n1094) );
  XNOR2_X1 U2111 ( .A(n37), .B(n1434), .ZN(n1093) );
  NAND2_X1 U2112 ( .A1(n1396), .A2(n1391), .ZN(n368) );
  AOI21_X1 U2113 ( .B1(n1396), .B2(n376), .A(n371), .ZN(n369) );
  AOI21_X1 U2114 ( .B1(n63), .B2(n245), .A(n246), .ZN(n244) );
  AOI21_X1 U2115 ( .B1(n63), .B2(n223), .A(n224), .ZN(n222) );
  XNOR2_X1 U2116 ( .A(n63), .B(n82), .ZN(product[23]) );
  AOI21_X1 U2117 ( .B1(n64), .B2(n232), .A(n233), .ZN(n231) );
  AOI21_X1 U2118 ( .B1(n64), .B2(n258), .A(n259), .ZN(n257) );
  AOI21_X1 U2119 ( .B1(n64), .B2(n278), .A(n1448), .ZN(n277) );
  AOI21_X1 U2120 ( .B1(n64), .B2(n425), .A(n288), .ZN(n286) );
  XOR2_X1 U2121 ( .A(n1444), .B(n98), .Z(product[7]) );
  NOR2_X1 U2122 ( .A1(n1409), .A2(n326), .ZN(n321) );
  AOI21_X1 U2123 ( .B1(n1400), .B2(n393), .A(n390), .ZN(n388) );
  OAI21_X1 U2124 ( .B1(n394), .B2(n396), .A(n395), .ZN(n393) );
  NAND2_X1 U2125 ( .A1(n1262), .A2(n1282), .ZN(n1272) );
  OAI21_X1 U2126 ( .B1(n1483), .B2(n318), .A(n313), .ZN(n311) );
  OAI21_X1 U2127 ( .B1(n1412), .B2(n108), .A(n109), .ZN(n107) );
  OAI21_X1 U2128 ( .B1(n1412), .B2(n117), .A(n118), .ZN(n116) );
  OAI21_X1 U2129 ( .B1(n1410), .B2(n201), .A(n202), .ZN(n200) );
  OAI21_X1 U2130 ( .B1(n1410), .B2(n171), .A(n172), .ZN(n170) );
  OAI21_X1 U2131 ( .B1(n65), .B2(n242), .A(n243), .ZN(n233) );
  OAI21_X1 U2132 ( .B1(n1410), .B2(n160), .A(n161), .ZN(n159) );
  OAI21_X1 U2133 ( .B1(n1410), .B2(n184), .A(n185), .ZN(n183) );
  OAI21_X1 U2134 ( .B1(n65), .B2(n216), .A(n217), .ZN(n211) );
  OAI21_X1 U2135 ( .B1(n65), .B2(n225), .A(n226), .ZN(n224) );
  OAI21_X1 U2136 ( .B1(n1410), .B2(n145), .A(n146), .ZN(n144) );
  OAI21_X1 U2137 ( .B1(n1410), .B2(n130), .A(n131), .ZN(n129) );
  XNOR2_X1 U2138 ( .A(n1), .B(n1248), .ZN(n1227) );
  XNOR2_X1 U2139 ( .A(n1), .B(n1251), .ZN(n1230) );
  XNOR2_X1 U2140 ( .A(n1), .B(n1252), .ZN(n1231) );
  XNOR2_X1 U2141 ( .A(n1), .B(n1247), .ZN(n1226) );
  XNOR2_X1 U2142 ( .A(n1), .B(n1246), .ZN(n1225) );
  XNOR2_X1 U2143 ( .A(n1), .B(n1243), .ZN(n1222) );
  XNOR2_X1 U2144 ( .A(n1), .B(n1242), .ZN(n1221) );
  XNOR2_X1 U2145 ( .A(n1), .B(n1241), .ZN(n1220) );
  XNOR2_X1 U2146 ( .A(n1), .B(n1245), .ZN(n1224) );
  XNOR2_X1 U2147 ( .A(n1), .B(n1244), .ZN(n1223) );
  XNOR2_X1 U2148 ( .A(n1), .B(n1253), .ZN(n1232) );
  XNOR2_X1 U2149 ( .A(n1), .B(n1254), .ZN(n1233) );
  XNOR2_X1 U2150 ( .A(n1), .B(n1255), .ZN(n1234) );
  XNOR2_X1 U2151 ( .A(n1250), .B(n1), .ZN(n1229) );
  XNOR2_X1 U2152 ( .A(n1), .B(n1249), .ZN(n1228) );
  XNOR2_X1 U2153 ( .A(n1384), .B(n1487), .ZN(n1238) );
  XNOR2_X1 U2154 ( .A(n1), .B(n1475), .ZN(n1235) );
  XNOR2_X1 U2155 ( .A(n1384), .B(n1258), .ZN(n1237) );
  XNOR2_X1 U2156 ( .A(n1), .B(n1240), .ZN(n1219) );
  XNOR2_X1 U2157 ( .A(n1384), .B(n1257), .ZN(n1236) );
  BUF_X4 U2158 ( .A(a[1]), .Z(n1) );
  AOI21_X1 U2159 ( .B1(n63), .B2(n199), .A(n200), .ZN(n198) );
  NOR2_X1 U2160 ( .A1(n247), .A2(n201), .ZN(n199) );
  AOI21_X1 U2161 ( .B1(n385), .B2(n1399), .A(n382), .ZN(n380) );
  AOI21_X1 U2162 ( .B1(n64), .B2(n269), .A(n270), .ZN(n268) );
  AOI21_X1 U2163 ( .B1(n311), .B2(n294), .A(n295), .ZN(n293) );
  XNOR2_X1 U2164 ( .A(a[8]), .B(a[7]), .ZN(n1285) );
  XOR2_X1 U2165 ( .A(a[6]), .B(a[7]), .Z(n1266) );
  XNOR2_X1 U2166 ( .A(n319), .B(n86), .ZN(product[19]) );
  AOI21_X1 U2167 ( .B1(n319), .B2(n306), .A(n1433), .ZN(n305) );
  AOI21_X1 U2168 ( .B1(n319), .B2(n315), .A(n316), .ZN(n314) );
  AOI21_X1 U2169 ( .B1(n299), .B2(n319), .A(n300), .ZN(n298) );
  XOR2_X1 U2170 ( .A(a[10]), .B(a[11]), .Z(n1264) );
  XNOR2_X1 U2171 ( .A(a[12]), .B(a[11]), .ZN(n1283) );
  NAND2_X1 U2172 ( .A1(n1264), .A2(n1284), .ZN(n1274) );
  XOR2_X1 U2173 ( .A(a[4]), .B(a[5]), .Z(n1267) );
  NAND2_X1 U2174 ( .A1(n1263), .A2(n1283), .ZN(n1273) );
  OAI21_X1 U2175 ( .B1(n292), .B2(n320), .A(n293), .ZN(n291) );
  INV_X1 U2176 ( .A(n320), .ZN(n319) );
  XOR2_X1 U2177 ( .A(a[16]), .B(a[17]), .Z(n1261) );
  NOR2_X1 U2178 ( .A1(n350), .A2(n355), .ZN(n348) );
  OAI21_X1 U2179 ( .B1(n1453), .B2(n356), .A(n351), .ZN(n349) );
  NAND2_X1 U2180 ( .A1(n707), .A2(n718), .ZN(n351) );
  XOR2_X1 U2181 ( .A(a[13]), .B(a[12]), .Z(n1263) );
  NOR2_X1 U2182 ( .A1(n289), .A2(n284), .ZN(n282) );
  XOR2_X1 U2183 ( .A(a[18]), .B(a[19]), .Z(n1260) );
  XOR2_X1 U2184 ( .A(a[8]), .B(a[9]), .Z(n1265) );
  XNOR2_X1 U2185 ( .A(n99), .B(n393), .ZN(product[6]) );
  XOR2_X1 U2186 ( .A(a[14]), .B(a[15]), .Z(n1262) );
  XNOR2_X1 U2187 ( .A(a[16]), .B(a[15]), .ZN(n1281) );
  XOR2_X1 U2188 ( .A(a[2]), .B(a[3]), .Z(n1268) );
  INV_X1 U2189 ( .A(n1408), .ZN(n339) );
  AOI21_X1 U2190 ( .B1(n340), .B2(n321), .A(n322), .ZN(n320) );
  OAI21_X1 U2191 ( .B1(n327), .B2(n323), .A(n324), .ZN(n322) );
  OAI21_X1 U2192 ( .B1(n341), .B2(n358), .A(n342), .ZN(n340) );
  XOR2_X1 U2193 ( .A(a[1]), .B(a[0]), .Z(n1269) );
  XOR2_X1 U2194 ( .A(n100), .B(n396), .Z(product[5]) );
endmodule


module datapath_DW_mult_tc_11 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n15, n16, n17, n18,
         n19, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34, n35,
         n36, n37, n40, n41, n42, n43, n45, n47, n48, n49, n51, n52, n54, n55,
         n57, n58, n59, n60, n61, n63, n64, n66, n67, n68, n69, n70, n71, n72,
         n73, n77, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n105, n106,
         n107, n108, n109, n111, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n124, n126, n127, n128, n129, n130, n131, n134,
         n135, n136, n137, n139, n141, n142, n143, n144, n145, n146, n149,
         n150, n151, n152, n154, n156, n157, n158, n159, n160, n161, n165,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n190,
         n191, n192, n193, n195, n197, n198, n199, n200, n201, n202, n206,
         n208, n209, n210, n211, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n254, n256, n257, n258, n259, n260, n261,
         n262, n263, n265, n267, n268, n269, n270, n273, n274, n275, n276,
         n277, n278, n280, n281, n282, n283, n284, n285, n286, n288, n289,
         n290, n291, n292, n293, n294, n295, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n309, n310, n311, n312, n313, n314,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n329, n331, n332, n333, n334, n339, n341, n342, n344, n346,
         n347, n348, n349, n350, n351, n352, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n371, n373, n374, n376, n378, n379, n380, n382, n384, n385, n386,
         n387, n388, n390, n392, n393, n394, n395, n396, n398, n400, n401,
         n402, n403, n404, n405, n406, n407, n409, n418, n424, n425, n426,
         n429, n435, n436, n437, n441, n443, n445, n446, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n793, n794, n796, n797, n799, n800, n802, n803, n805, n806, n808,
         n809, n811, n812, n814, n815, n817, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483;
  assign product[39] = n105;

  FA_X1 U488 ( .A(n831), .B(n454), .CI(n850), .CO(n450), .S(n451) );
  FA_X1 U489 ( .A(n455), .B(n832), .CI(n458), .CO(n452), .S(n453) );
  FA_X1 U491 ( .A(n462), .B(n833), .CI(n459), .CO(n456), .S(n457) );
  FA_X1 U492 ( .A(n851), .B(n464), .CI(n870), .CO(n458), .S(n459) );
  FA_X1 U493 ( .A(n463), .B(n470), .CI(n468), .CO(n460), .S(n461) );
  FA_X1 U494 ( .A(n834), .B(n852), .CI(n465), .CO(n462), .S(n463) );
  FA_X1 U496 ( .A(n474), .B(n471), .CI(n469), .CO(n466), .S(n467) );
  FA_X1 U497 ( .A(n478), .B(n871), .CI(n476), .CO(n468), .S(n469) );
  FA_X1 U498 ( .A(n853), .B(n835), .CI(n890), .CO(n470), .S(n471) );
  FA_X1 U499 ( .A(n475), .B(n477), .CI(n482), .CO(n472), .S(n473) );
  FA_X1 U500 ( .A(n486), .B(n479), .CI(n484), .CO(n474), .S(n475) );
  FA_X1 U501 ( .A(n836), .B(n854), .CI(n872), .CO(n476), .S(n477) );
  FA_X1 U503 ( .A(n490), .B(n492), .CI(n483), .CO(n480), .S(n481) );
  FA_X1 U504 ( .A(n485), .B(n494), .CI(n487), .CO(n482), .S(n483) );
  FA_X1 U505 ( .A(n855), .B(n496), .CI(n873), .CO(n484), .S(n485) );
  FA_X1 U506 ( .A(n891), .B(n837), .CI(n910), .CO(n486), .S(n487) );
  FA_X1 U507 ( .A(n500), .B(n493), .CI(n491), .CO(n488), .S(n489) );
  FA_X1 U508 ( .A(n495), .B(n504), .CI(n502), .CO(n490), .S(n491) );
  FA_X1 U509 ( .A(n497), .B(n874), .CI(n506), .CO(n492), .S(n493) );
  FA_X1 U510 ( .A(n892), .B(n856), .CI(n838), .CO(n494), .S(n495) );
  FA_X1 U512 ( .A(n510), .B(n503), .CI(n501), .CO(n498), .S(n499) );
  FA_X1 U513 ( .A(n507), .B(n505), .CI(n512), .CO(n500), .S(n501) );
  FA_X1 U514 ( .A(n516), .B(n893), .CI(n514), .CO(n502), .S(n503) );
  FA_X1 U515 ( .A(n857), .B(n911), .CI(n875), .CO(n504), .S(n505) );
  FA_X1 U516 ( .A(n518), .B(n839), .CI(n930), .CO(n506), .S(n507) );
  FA_X1 U517 ( .A(n522), .B(n513), .CI(n511), .CO(n508), .S(n509) );
  FA_X1 U518 ( .A(n526), .B(n515), .CI(n524), .CO(n510), .S(n511) );
  FA_X1 U519 ( .A(n528), .B(n530), .CI(n517), .CO(n512), .S(n513) );
  FA_X1 U520 ( .A(n840), .B(n858), .CI(n519), .CO(n514), .S(n515) );
  FA_X1 U521 ( .A(n912), .B(n876), .CI(n894), .CO(n516), .S(n517) );
  FA_X1 U523 ( .A(n534), .B(n525), .CI(n523), .CO(n520), .S(n521) );
  FA_X1 U524 ( .A(n527), .B(n538), .CI(n536), .CO(n522), .S(n523) );
  FA_X1 U525 ( .A(n529), .B(n540), .CI(n531), .CO(n524), .S(n525) );
  FA_X1 U526 ( .A(n877), .B(n895), .CI(n542), .CO(n526), .S(n527) );
  FA_X1 U527 ( .A(n859), .B(n931), .CI(n913), .CO(n528), .S(n529) );
  FA_X1 U528 ( .A(n544), .B(n841), .CI(n950), .CO(n530), .S(n531) );
  FA_X1 U529 ( .A(n548), .B(n537), .CI(n535), .CO(n532), .S(n533) );
  FA_X1 U530 ( .A(n539), .B(n552), .CI(n550), .CO(n534), .S(n535) );
  FA_X1 U531 ( .A(n541), .B(n554), .CI(n543), .CO(n536), .S(n537) );
  FA_X1 U532 ( .A(n558), .B(n545), .CI(n556), .CO(n538), .S(n539) );
  FA_X1 U533 ( .A(n896), .B(n932), .CI(n914), .CO(n540), .S(n541) );
  FA_X1 U534 ( .A(n842), .B(n878), .CI(n860), .CO(n542), .S(n543) );
  FA_X1 U536 ( .A(n562), .B(n551), .CI(n549), .CO(n546), .S(n547) );
  FA_X1 U537 ( .A(n553), .B(n566), .CI(n564), .CO(n548), .S(n549) );
  FA_X1 U538 ( .A(n559), .B(n557), .CI(n568), .CO(n550), .S(n551) );
  FA_X1 U539 ( .A(n570), .B(n572), .CI(n555), .CO(n552), .S(n553) );
  FA_X1 U540 ( .A(n879), .B(n915), .CI(n897), .CO(n554), .S(n555) );
  FA_X1 U541 ( .A(n861), .B(n951), .CI(n933), .CO(n556), .S(n557) );
  FA_X1 U542 ( .A(n574), .B(n843), .CI(n970), .CO(n558), .S(n559) );
  FA_X1 U543 ( .A(n578), .B(n565), .CI(n563), .CO(n560), .S(n561) );
  FA_X1 U544 ( .A(n567), .B(n582), .CI(n580), .CO(n562), .S(n563) );
  FA_X1 U545 ( .A(n584), .B(n573), .CI(n569), .CO(n564), .S(n565) );
  FA_X1 U546 ( .A(n586), .B(n588), .CI(n571), .CO(n566), .S(n567) );
  FA_X1 U547 ( .A(n575), .B(n898), .CI(n590), .CO(n568), .S(n569) );
  FA_X1 U548 ( .A(n844), .B(n916), .CI(n862), .CO(n570), .S(n571) );
  FA_X1 U549 ( .A(n952), .B(n880), .CI(n934), .CO(n572), .S(n573) );
  FA_X1 U552 ( .A(n583), .B(n598), .CI(n596), .CO(n578), .S(n579) );
  FA_X1 U553 ( .A(n600), .B(n591), .CI(n585), .CO(n580), .S(n581) );
  FA_X1 U554 ( .A(n587), .B(n602), .CI(n589), .CO(n582), .S(n583) );
  FA_X1 U555 ( .A(n606), .B(n917), .CI(n604), .CO(n584), .S(n585) );
  FA_X1 U556 ( .A(n881), .B(n935), .CI(n899), .CO(n586), .S(n587) );
  FA_X1 U557 ( .A(n608), .B(n953), .CI(n863), .CO(n588), .S(n589) );
  FA_X1 U558 ( .A(n971), .B(n845), .CI(n990), .CO(n590), .S(n591) );
  FA_X1 U559 ( .A(n612), .B(n597), .CI(n595), .CO(n592), .S(n593) );
  FA_X1 U560 ( .A(n599), .B(n616), .CI(n614), .CO(n594), .S(n595) );
  FA_X1 U561 ( .A(n618), .B(n603), .CI(n601), .CO(n596), .S(n597) );
  FA_X1 U562 ( .A(n605), .B(n620), .CI(n607), .CO(n598), .S(n599) );
  FA_X1 U563 ( .A(n624), .B(n626), .CI(n622), .CO(n600), .S(n601) );
  FA_X1 U564 ( .A(n918), .B(n936), .CI(n609), .CO(n602), .S(n603) );
  FA_X1 U565 ( .A(n954), .B(n864), .CI(n882), .CO(n604), .S(n605) );
  FA_X1 U566 ( .A(n900), .B(n846), .CI(n972), .CO(n606), .S(n607) );
  FA_X1 U568 ( .A(n630), .B(n615), .CI(n613), .CO(n610), .S(n611) );
  FA_X1 U569 ( .A(n617), .B(n634), .CI(n632), .CO(n612), .S(n613) );
  FA_X1 U570 ( .A(n636), .B(n621), .CI(n619), .CO(n614), .S(n615) );
  FA_X1 U571 ( .A(n623), .B(n638), .CI(n625), .CO(n616), .S(n617) );
  FA_X1 U572 ( .A(n627), .B(n642), .CI(n640), .CO(n618), .S(n619) );
  FA_X1 U573 ( .A(n955), .B(n973), .CI(n644), .CO(n620), .S(n621) );
  FA_X1 U574 ( .A(n991), .B(n901), .CI(n883), .CO(n622), .S(n623) );
  FA_X1 U575 ( .A(n847), .B(n919), .CI(n1010), .CO(n624), .S(n625) );
  FA_X1 U578 ( .A(n648), .B(n633), .CI(n631), .CO(n628), .S(n629) );
  FA_X1 U579 ( .A(n650), .B(n637), .CI(n635), .CO(n630), .S(n631) );
  FA_X1 U580 ( .A(n654), .B(n643), .CI(n652), .CO(n632), .S(n633) );
  FA_X1 U581 ( .A(n639), .B(n656), .CI(n641), .CO(n634), .S(n635) );
  FA_X1 U582 ( .A(n660), .B(n645), .CI(n658), .CO(n636), .S(n637) );
  FA_X1 U583 ( .A(n920), .B(n992), .CI(n974), .CO(n638), .S(n639) );
  FA_X1 U584 ( .A(n1011), .B(n956), .CI(n902), .CO(n640), .S(n641) );
  FA_X1 U585 ( .A(n866), .B(n884), .CI(n938), .CO(n642), .S(n643) );
  HA_X1 U586 ( .A(n820), .B(n848), .CO(n644), .S(n645) );
  FA_X1 U587 ( .A(n664), .B(n651), .CI(n649), .CO(n646), .S(n647) );
  FA_X1 U588 ( .A(n666), .B(n655), .CI(n653), .CO(n648), .S(n649) );
  FA_X1 U589 ( .A(n670), .B(n659), .CI(n668), .CO(n650), .S(n651) );
  FA_X1 U590 ( .A(n661), .B(n672), .CI(n657), .CO(n652), .S(n653) );
  FA_X1 U591 ( .A(n676), .B(n957), .CI(n674), .CO(n654), .S(n655) );
  FA_X1 U592 ( .A(n939), .B(n975), .CI(n921), .CO(n656), .S(n657) );
  FA_X1 U593 ( .A(n867), .B(n993), .CI(n903), .CO(n658), .S(n659) );
  FA_X1 U594 ( .A(n849), .B(n885), .CI(n1012), .CO(n660), .S(n661) );
  FA_X1 U595 ( .A(n667), .B(n680), .CI(n665), .CO(n662), .S(n663) );
  FA_X1 U596 ( .A(n682), .B(n671), .CI(n669), .CO(n664), .S(n665) );
  FA_X1 U597 ( .A(n675), .B(n673), .CI(n684), .CO(n666), .S(n667) );
  FA_X1 U598 ( .A(n686), .B(n688), .CI(n690), .CO(n668), .S(n669) );
  FA_X1 U599 ( .A(n958), .B(n976), .CI(n677), .CO(n670), .S(n671) );
  FA_X1 U600 ( .A(n886), .B(n904), .CI(n922), .CO(n672), .S(n673) );
  FA_X1 U601 ( .A(n1013), .B(n940), .CI(n994), .CO(n674), .S(n675) );
  HA_X1 U602 ( .A(n821), .B(n868), .CO(n676), .S(n677) );
  FA_X1 U604 ( .A(n696), .B(n698), .CI(n685), .CO(n680), .S(n681) );
  FA_X1 U606 ( .A(n702), .B(n704), .CI(n700), .CO(n684), .S(n685) );
  FA_X1 U607 ( .A(n959), .B(n977), .CI(n941), .CO(n686), .S(n687) );
  FA_X1 U608 ( .A(n923), .B(n887), .CI(n995), .CO(n688), .S(n689) );
  FA_X1 U609 ( .A(n869), .B(n905), .CI(n1014), .CO(n690), .S(n691) );
  FA_X1 U610 ( .A(n697), .B(n708), .CI(n695), .CO(n692), .S(n693) );
  FA_X1 U611 ( .A(n710), .B(n703), .CI(n699), .CO(n694), .S(n695) );
  FA_X1 U612 ( .A(n712), .B(n714), .CI(n701), .CO(n696), .S(n697) );
  FA_X1 U613 ( .A(n705), .B(n996), .CI(n716), .CO(n698), .S(n699) );
  FA_X1 U614 ( .A(n978), .B(n942), .CI(n1015), .CO(n700), .S(n701) );
  FA_X1 U615 ( .A(n960), .B(n906), .CI(n924), .CO(n702), .S(n703) );
  HA_X1 U616 ( .A(n822), .B(n888), .CO(n704), .S(n705) );
  FA_X1 U617 ( .A(n711), .B(n720), .CI(n709), .CO(n706), .S(n707) );
  FA_X1 U618 ( .A(n713), .B(n715), .CI(n722), .CO(n708), .S(n709) );
  FA_X1 U619 ( .A(n724), .B(n726), .CI(n717), .CO(n710), .S(n711) );
  FA_X1 U620 ( .A(n961), .B(n979), .CI(n728), .CO(n712), .S(n713) );
  FA_X1 U621 ( .A(n907), .B(n997), .CI(n943), .CO(n714), .S(n715) );
  FA_X1 U622 ( .A(n925), .B(n889), .CI(n1016), .CO(n716), .S(n717) );
  FA_X1 U623 ( .A(n732), .B(n723), .CI(n721), .CO(n718), .S(n719) );
  FA_X1 U624 ( .A(n727), .B(n725), .CI(n734), .CO(n720), .S(n721) );
  FA_X1 U625 ( .A(n738), .B(n729), .CI(n736), .CO(n722), .S(n723) );
  FA_X1 U626 ( .A(n926), .B(n980), .CI(n944), .CO(n724), .S(n725) );
  FA_X1 U627 ( .A(n1017), .B(n962), .CI(n998), .CO(n726), .S(n727) );
  HA_X1 U628 ( .A(n823), .B(n908), .CO(n728), .S(n729) );
  FA_X1 U629 ( .A(n735), .B(n742), .CI(n733), .CO(n730), .S(n731) );
  FA_X1 U630 ( .A(n737), .B(n739), .CI(n744), .CO(n732), .S(n733) );
  FA_X1 U631 ( .A(n748), .B(n981), .CI(n746), .CO(n734), .S(n735) );
  FA_X1 U632 ( .A(n927), .B(n999), .CI(n963), .CO(n736), .S(n737) );
  FA_X1 U633 ( .A(n945), .B(n909), .CI(n1018), .CO(n738), .S(n739) );
  FA_X1 U634 ( .A(n752), .B(n745), .CI(n743), .CO(n740), .S(n741) );
  FA_X1 U635 ( .A(n754), .B(n756), .CI(n747), .CO(n742), .S(n743) );
  FA_X1 U636 ( .A(n964), .B(n1000), .CI(n749), .CO(n744), .S(n745) );
  FA_X1 U637 ( .A(n946), .B(n982), .CI(n1019), .CO(n746), .S(n747) );
  HA_X1 U638 ( .A(n824), .B(n928), .CO(n748), .S(n749) );
  FA_X1 U639 ( .A(n760), .B(n755), .CI(n753), .CO(n750), .S(n751) );
  FA_X1 U640 ( .A(n762), .B(n764), .CI(n757), .CO(n752), .S(n753) );
  FA_X1 U641 ( .A(n947), .B(n1001), .CI(n983), .CO(n754), .S(n755) );
  FA_X1 U642 ( .A(n965), .B(n929), .CI(n1020), .CO(n756), .S(n757) );
  FA_X1 U643 ( .A(n763), .B(n768), .CI(n761), .CO(n758), .S(n759) );
  FA_X1 U644 ( .A(n765), .B(n1021), .CI(n770), .CO(n760), .S(n761) );
  FA_X1 U645 ( .A(n966), .B(n984), .CI(n1002), .CO(n762), .S(n763) );
  HA_X1 U646 ( .A(n825), .B(n948), .CO(n764), .S(n765) );
  FA_X1 U647 ( .A(n771), .B(n774), .CI(n769), .CO(n766), .S(n767) );
  FA_X1 U648 ( .A(n967), .B(n1003), .CI(n776), .CO(n768), .S(n769) );
  FA_X1 U649 ( .A(n985), .B(n949), .CI(n1022), .CO(n770), .S(n771) );
  FA_X1 U650 ( .A(n780), .B(n777), .CI(n775), .CO(n772), .S(n773) );
  FA_X1 U651 ( .A(n986), .B(n1023), .CI(n1004), .CO(n774), .S(n775) );
  HA_X1 U652 ( .A(n826), .B(n968), .CO(n776), .S(n777) );
  FA_X1 U653 ( .A(n784), .B(n987), .CI(n781), .CO(n778), .S(n779) );
  FA_X1 U654 ( .A(n1024), .B(n969), .CI(n1005), .CO(n780), .S(n781) );
  FA_X1 U655 ( .A(n1006), .B(n1025), .CI(n785), .CO(n782), .S(n783) );
  HA_X1 U656 ( .A(n827), .B(n988), .CO(n784), .S(n785) );
  FA_X1 U657 ( .A(n1026), .B(n989), .CI(n1007), .CO(n786), .S(n787) );
  HA_X1 U658 ( .A(n1008), .B(n1027), .CO(n788), .S(n789) );
  CLKBUF_X1 U1180 ( .A(n611), .Z(n1383) );
  CLKBUF_X1 U1181 ( .A(n1286), .Z(n21) );
  CLKBUF_X1 U1182 ( .A(n1277), .Z(n17) );
  CLKBUF_X3 U1183 ( .A(n1277), .Z(n18) );
  CLKBUF_X3 U1184 ( .A(n1276), .Z(n24) );
  INV_X1 U1185 ( .A(n1413), .ZN(n1384) );
  AOI21_X1 U1186 ( .B1(n283), .B2(n249), .A(n250), .ZN(n1432) );
  CLKBUF_X3 U1187 ( .A(n1270), .Z(n59) );
  CLKBUF_X1 U1188 ( .A(n1184), .Z(n1385) );
  CLKBUF_X1 U1189 ( .A(n1127), .Z(n1386) );
  CLKBUF_X1 U1190 ( .A(n1288), .Z(n9) );
  BUF_X1 U1191 ( .A(n1288), .Z(n10) );
  CLKBUF_X3 U1192 ( .A(b[4]), .Z(n1255) );
  CLKBUF_X2 U1193 ( .A(b[7]), .Z(n1252) );
  CLKBUF_X2 U1194 ( .A(b[16]), .Z(n1243) );
  BUF_X1 U1195 ( .A(n1462), .Z(n1387) );
  CLKBUF_X1 U1196 ( .A(n21), .Z(n1388) );
  BUF_X2 U1197 ( .A(n21), .Z(n1389) );
  BUF_X2 U1198 ( .A(n1282), .Z(n45) );
  CLKBUF_X3 U1199 ( .A(n1273), .Z(n41) );
  NOR2_X2 U1200 ( .A1(n577), .A2(n592), .ZN(n1466) );
  CLKBUF_X3 U1201 ( .A(n1276), .Z(n23) );
  CLKBUF_X1 U1202 ( .A(n1), .Z(n1390) );
  XOR2_X1 U1203 ( .A(n689), .B(n687), .Z(n1391) );
  XOR2_X1 U1204 ( .A(n691), .B(n1391), .Z(n683) );
  NAND2_X1 U1205 ( .A1(n691), .A2(n689), .ZN(n1392) );
  NAND2_X1 U1206 ( .A1(n691), .A2(n687), .ZN(n1393) );
  NAND2_X1 U1207 ( .A1(n689), .A2(n687), .ZN(n1394) );
  NAND3_X1 U1208 ( .A1(n1392), .A2(n1393), .A3(n1394), .ZN(n682) );
  CLKBUF_X3 U1209 ( .A(b[13]), .Z(n1246) );
  CLKBUF_X3 U1210 ( .A(b[6]), .Z(n1253) );
  OR2_X1 U1211 ( .A1(n692), .A2(n679), .ZN(n1460) );
  BUF_X1 U1212 ( .A(b[9]), .Z(n1477) );
  CLKBUF_X3 U1213 ( .A(b[18]), .Z(n1241) );
  CLKBUF_X3 U1214 ( .A(n49), .Z(n1480) );
  CLKBUF_X3 U1215 ( .A(b[1]), .Z(n1258) );
  BUF_X1 U1216 ( .A(n1279), .Z(n6) );
  BUF_X1 U1217 ( .A(a[17]), .Z(n49) );
  BUF_X2 U1218 ( .A(b[14]), .Z(n1245) );
  BUF_X2 U1219 ( .A(n61), .Z(n1450) );
  BUF_X2 U1220 ( .A(n61), .Z(n1449) );
  BUF_X2 U1221 ( .A(n248), .Z(n1453) );
  OR2_X1 U1222 ( .A1(n473), .A2(n480), .ZN(n1395) );
  OR2_X1 U1223 ( .A1(n759), .A2(n766), .ZN(n1396) );
  OR2_X1 U1224 ( .A1(n453), .A2(n456), .ZN(n1397) );
  OR2_X1 U1225 ( .A1(n467), .A2(n472), .ZN(n1398) );
  OR2_X1 U1226 ( .A1(n779), .A2(n782), .ZN(n1399) );
  OR2_X1 U1227 ( .A1(n830), .A2(n448), .ZN(n1400) );
  OR2_X1 U1228 ( .A1(n452), .A2(n451), .ZN(n1401) );
  OR2_X1 U1229 ( .A1(n693), .A2(n706), .ZN(n1402) );
  OR2_X1 U1230 ( .A1(n450), .A2(n449), .ZN(n1403) );
  OR2_X1 U1231 ( .A1(n751), .A2(n758), .ZN(n1404) );
  OR2_X1 U1232 ( .A1(n509), .A2(n520), .ZN(n1405) );
  AND2_X1 U1233 ( .A1(n1411), .A2(n409), .ZN(product[1]) );
  OR2_X1 U1234 ( .A1(n457), .A2(n460), .ZN(n1407) );
  OR2_X1 U1235 ( .A1(n767), .A2(n772), .ZN(n1408) );
  OR2_X1 U1236 ( .A1(n787), .A2(n788), .ZN(n1409) );
  AND2_X1 U1237 ( .A1(n679), .A2(n692), .ZN(n1410) );
  OR2_X1 U1238 ( .A1(n1029), .A2(n829), .ZN(n1411) );
  NOR2_X1 U1239 ( .A1(n593), .A2(n610), .ZN(n303) );
  OR2_X1 U1240 ( .A1(n707), .A2(n718), .ZN(n1412) );
  OR2_X1 U1241 ( .A1(n1383), .A2(n628), .ZN(n1413) );
  CLKBUF_X1 U1242 ( .A(n311), .Z(n1414) );
  OR2_X1 U1243 ( .A1(n1384), .A2(n317), .ZN(n1415) );
  CLKBUF_X1 U1244 ( .A(n19), .Z(n1416) );
  OAI22_X1 U1245 ( .A1(n60), .A2(n1031), .B1(n58), .B2(n1030), .ZN(n448) );
  CLKBUF_X1 U1246 ( .A(n63), .Z(n1417) );
  XNOR2_X1 U1247 ( .A(a[12]), .B(a[11]), .ZN(n1418) );
  BUF_X2 U1248 ( .A(n1418), .Z(n1422) );
  OAI21_X1 U1249 ( .B1(n284), .B2(n290), .A(n285), .ZN(n1419) );
  NOR2_X2 U1250 ( .A1(n547), .A2(n560), .ZN(n284) );
  OR2_X1 U1251 ( .A1(n521), .A2(n532), .ZN(n1420) );
  BUF_X2 U1252 ( .A(n1418), .Z(n1421) );
  BUF_X1 U1253 ( .A(n291), .Z(n1478) );
  BUF_X1 U1254 ( .A(n1283), .Z(n40) );
  BUF_X1 U1255 ( .A(n1272), .Z(n47) );
  NAND2_X2 U1256 ( .A1(n1261), .A2(n1281), .ZN(n1423) );
  XNOR2_X2 U1257 ( .A(a[16]), .B(a[15]), .ZN(n1281) );
  OR2_X2 U1258 ( .A1(n663), .A2(n678), .ZN(n1424) );
  XNOR2_X1 U1259 ( .A(n579), .B(n1425), .ZN(n577) );
  XNOR2_X1 U1260 ( .A(n594), .B(n581), .ZN(n1425) );
  BUF_X2 U1261 ( .A(n1270), .Z(n60) );
  NAND2_X1 U1262 ( .A1(n579), .A2(n594), .ZN(n1426) );
  NAND2_X1 U1263 ( .A1(n579), .A2(n581), .ZN(n1427) );
  NAND2_X1 U1264 ( .A1(n594), .A2(n581), .ZN(n1428) );
  NAND3_X1 U1265 ( .A1(n1426), .A2(n1427), .A3(n1428), .ZN(n576) );
  BUF_X2 U1266 ( .A(n1272), .Z(n48) );
  BUF_X2 U1267 ( .A(n1279), .Z(n1429) );
  NOR2_X1 U1268 ( .A1(n611), .A2(n628), .ZN(n1430) );
  NOR2_X1 U1269 ( .A1(n611), .A2(n628), .ZN(n312) );
  XNOR2_X1 U1270 ( .A(n7), .B(n1245), .ZN(n1431) );
  BUF_X1 U1271 ( .A(n61), .Z(n1482) );
  BUF_X1 U1272 ( .A(n1282), .Z(n1433) );
  CLKBUF_X3 U1273 ( .A(n1272), .Z(n1434) );
  CLKBUF_X3 U1274 ( .A(a[5]), .Z(n1435) );
  CLKBUF_X1 U1275 ( .A(a[5]), .Z(n13) );
  CLKBUF_X1 U1276 ( .A(b[0]), .Z(n61) );
  OR2_X1 U1277 ( .A1(n647), .A2(n662), .ZN(n1436) );
  INV_X1 U1278 ( .A(n1290), .ZN(n1437) );
  INV_X1 U1279 ( .A(n1480), .ZN(n1438) );
  INV_X1 U1280 ( .A(n1438), .ZN(n1439) );
  CLKBUF_X1 U1281 ( .A(n37), .Z(n1440) );
  XNOR2_X1 U1282 ( .A(n43), .B(n1255), .ZN(n1441) );
  CLKBUF_X1 U1283 ( .A(n322), .Z(n1442) );
  BUF_X2 U1284 ( .A(n1281), .Z(n52) );
  BUF_X2 U1285 ( .A(n1280), .Z(n57) );
  CLKBUF_X3 U1286 ( .A(a[11]), .Z(n1443) );
  CLKBUF_X1 U1287 ( .A(a[11]), .Z(n31) );
  CLKBUF_X1 U1288 ( .A(n43), .Z(n1444) );
  CLKBUF_X3 U1289 ( .A(n1273), .Z(n42) );
  BUF_X2 U1290 ( .A(n1281), .Z(n51) );
  BUF_X1 U1291 ( .A(n1278), .Z(n1445) );
  BUF_X1 U1292 ( .A(n1278), .Z(n1446) );
  BUF_X1 U1293 ( .A(n1275), .Z(n1447) );
  BUF_X1 U1294 ( .A(n1275), .Z(n1448) );
  XNOR2_X1 U1295 ( .A(n277), .B(n1451), .ZN(product[25]) );
  AND2_X1 U1296 ( .A1(n273), .A2(n276), .ZN(n1451) );
  NOR2_X1 U1297 ( .A1(n707), .A2(n718), .ZN(n350) );
  CLKBUF_X1 U1298 ( .A(n1), .Z(n1452) );
  CLKBUF_X3 U1299 ( .A(b[15]), .Z(n1244) );
  CLKBUF_X3 U1300 ( .A(b[12]), .Z(n1247) );
  XNOR2_X1 U1301 ( .A(n257), .B(n1454), .ZN(product[27]) );
  AND2_X1 U1302 ( .A1(n1405), .A2(n256), .ZN(n1454) );
  XNOR2_X1 U1303 ( .A(n268), .B(n1455), .ZN(product[26]) );
  AND2_X1 U1304 ( .A1(n262), .A2(n267), .ZN(n1455) );
  BUF_X2 U1305 ( .A(n1274), .Z(n35) );
  XOR2_X1 U1306 ( .A(n694), .B(n683), .Z(n1456) );
  XOR2_X1 U1307 ( .A(n681), .B(n1456), .Z(n679) );
  NAND2_X1 U1308 ( .A1(n681), .A2(n694), .ZN(n1457) );
  NAND2_X1 U1309 ( .A1(n681), .A2(n683), .ZN(n1458) );
  NAND2_X1 U1310 ( .A1(n694), .A2(n683), .ZN(n1459) );
  NAND3_X1 U1311 ( .A1(n1457), .A2(n1458), .A3(n1459), .ZN(n678) );
  CLKBUF_X3 U1312 ( .A(b[17]), .Z(n1242) );
  BUF_X4 U1313 ( .A(a[9]), .Z(n25) );
  BUF_X4 U1314 ( .A(a[13]), .Z(n37) );
  BUF_X4 U1315 ( .A(a[3]), .Z(n7) );
  CLKBUF_X1 U1316 ( .A(b[19]), .Z(n1469) );
  CLKBUF_X1 U1317 ( .A(b[19]), .Z(n1240) );
  CLKBUF_X1 U1318 ( .A(b[2]), .Z(n1472) );
  CLKBUF_X1 U1319 ( .A(b[2]), .Z(n1471) );
  CLKBUF_X1 U1320 ( .A(b[2]), .Z(n1257) );
  CLKBUF_X1 U1321 ( .A(n1453), .Z(n1461) );
  BUF_X4 U1322 ( .A(a[15]), .Z(n43) );
  CLKBUF_X1 U1323 ( .A(b[8]), .Z(n1473) );
  CLKBUF_X1 U1324 ( .A(b[8]), .Z(n1474) );
  CLKBUF_X1 U1325 ( .A(b[8]), .Z(n1251) );
  CLKBUF_X1 U1326 ( .A(b[19]), .Z(n1468) );
  CLKBUF_X3 U1327 ( .A(b[10]), .Z(n1249) );
  BUF_X4 U1328 ( .A(a[1]), .Z(n1) );
  BUF_X2 U1329 ( .A(n1271), .Z(n54) );
  OAI21_X1 U1330 ( .B1(n341), .B2(n358), .A(n342), .ZN(n1462) );
  BUF_X4 U1331 ( .A(n49), .Z(n1479) );
  XNOR2_X1 U1332 ( .A(n286), .B(n1463), .ZN(product[24]) );
  AND2_X1 U1333 ( .A1(n424), .A2(n285), .ZN(n1463) );
  BUF_X4 U1334 ( .A(a[7]), .Z(n19) );
  CLKBUF_X3 U1335 ( .A(b[11]), .Z(n1248) );
  CLKBUF_X3 U1336 ( .A(b[5]), .Z(n1254) );
  XNOR2_X1 U1337 ( .A(n222), .B(n1464), .ZN(product[30]) );
  AND2_X1 U1338 ( .A1(n418), .A2(n221), .ZN(n1464) );
  NOR2_X1 U1339 ( .A1(n303), .A2(n1466), .ZN(n1465) );
  CLKBUF_X1 U1340 ( .A(b[3]), .Z(n1256) );
  CLKBUF_X1 U1341 ( .A(b[3]), .Z(n1475) );
  CLKBUF_X1 U1342 ( .A(b[3]), .Z(n1476) );
  CLKBUF_X1 U1343 ( .A(b[9]), .Z(n1250) );
  XNOR2_X1 U1344 ( .A(n231), .B(n1467), .ZN(product[29]) );
  AND2_X1 U1345 ( .A1(n227), .A2(n230), .ZN(n1467) );
  XNOR2_X1 U1346 ( .A(n209), .B(n1470), .ZN(product[31]) );
  AND2_X1 U1347 ( .A1(n1395), .A2(n208), .ZN(n1470) );
  BUF_X1 U1348 ( .A(n61), .Z(n1483) );
  BUF_X2 U1349 ( .A(n247), .Z(n66) );
  CLKBUF_X3 U1350 ( .A(a[19]), .Z(n55) );
  NOR2_X1 U1351 ( .A1(n629), .A2(n646), .ZN(n317) );
  NOR2_X1 U1352 ( .A1(n533), .A2(n546), .ZN(n275) );
  NOR2_X1 U1353 ( .A1(n647), .A2(n662), .ZN(n323) );
  NOR2_X1 U1354 ( .A1(n461), .A2(n466), .ZN(n179) );
  NOR2_X1 U1355 ( .A1(n489), .A2(n498), .ZN(n229) );
  NOR2_X1 U1356 ( .A1(n731), .A2(n740), .ZN(n361) );
  NOR2_X1 U1357 ( .A1(n719), .A2(n730), .ZN(n355) );
  NOR2_X1 U1358 ( .A1(n481), .A2(n488), .ZN(n220) );
  NOR2_X1 U1359 ( .A1(n741), .A2(n750), .ZN(n364) );
  NOR2_X1 U1360 ( .A1(n499), .A2(n508), .ZN(n242) );
  NOR2_X1 U1361 ( .A1(n1028), .A2(n1009), .ZN(n406) );
  NOR2_X1 U1362 ( .A1(n783), .A2(n786), .ZN(n394) );
  NOR2_X1 U1363 ( .A1(n773), .A2(n778), .ZN(n386) );
  NOR2_X1 U1364 ( .A1(n789), .A2(n828), .ZN(n402) );
  BUF_X1 U1365 ( .A(n1287), .Z(n15) );
  NAND2_X1 U1366 ( .A1(n1265), .A2(n1285), .ZN(n1275) );
  NAND2_X1 U1367 ( .A1(n1266), .A2(n1286), .ZN(n1276) );
  NAND2_X1 U1368 ( .A1(n1260), .A2(n1280), .ZN(n1270) );
  NAND2_X1 U1369 ( .A1(n1263), .A2(n1283), .ZN(n1273) );
  NAND2_X1 U1370 ( .A1(n1262), .A2(n1282), .ZN(n1272) );
  NAND2_X1 U1371 ( .A1(n1264), .A2(n1284), .ZN(n1274) );
  INV_X1 U1372 ( .A(a[0]), .ZN(n1289) );
  BUF_X1 U1373 ( .A(n291), .Z(n63) );
  BUF_X1 U1374 ( .A(n291), .Z(n64) );
  NOR2_X1 U1375 ( .A1(n280), .A2(n275), .ZN(n269) );
  NOR2_X1 U1376 ( .A1(n280), .A2(n260), .ZN(n258) );
  NAND2_X1 U1377 ( .A1(n214), .A2(n134), .ZN(n130) );
  INV_X1 U1378 ( .A(n1415), .ZN(n306) );
  INV_X1 U1379 ( .A(n280), .ZN(n278) );
  INV_X1 U1380 ( .A(n173), .ZN(n171) );
  INV_X1 U1381 ( .A(n186), .ZN(n184) );
  INV_X1 U1382 ( .A(n66), .ZN(n245) );
  INV_X1 U1383 ( .A(n1481), .ZN(n319) );
  INV_X1 U1384 ( .A(n282), .ZN(n280) );
  INV_X1 U1385 ( .A(n1387), .ZN(n339) );
  NAND2_X1 U1386 ( .A1(n310), .A2(n294), .ZN(n292) );
  AOI21_X1 U1387 ( .B1(n311), .B2(n1465), .A(n295), .ZN(n293) );
  NOR2_X1 U1388 ( .A1(n216), .A2(n192), .ZN(n186) );
  NOR2_X1 U1389 ( .A1(n216), .A2(n175), .ZN(n173) );
  INV_X1 U1390 ( .A(n187), .ZN(n185) );
  NAND2_X1 U1391 ( .A1(n282), .A2(n249), .ZN(n247) );
  NOR2_X1 U1392 ( .A1(n1415), .A2(n301), .ZN(n299) );
  INV_X1 U1393 ( .A(n283), .ZN(n281) );
  INV_X1 U1394 ( .A(n216), .ZN(n214) );
  NAND2_X1 U1395 ( .A1(n1424), .A2(n1460), .ZN(n326) );
  NAND2_X1 U1396 ( .A1(n1420), .A2(n1405), .ZN(n251) );
  NAND2_X1 U1397 ( .A1(n273), .A2(n262), .ZN(n260) );
  OAI21_X1 U1398 ( .B1(n281), .B2(n275), .A(n276), .ZN(n270) );
  OAI21_X1 U1399 ( .B1(n281), .B2(n260), .A(n261), .ZN(n259) );
  AOI21_X1 U1400 ( .B1(n274), .B2(n262), .A(n265), .ZN(n261) );
  INV_X1 U1401 ( .A(n1414), .ZN(n309) );
  INV_X1 U1402 ( .A(n192), .ZN(n190) );
  INV_X1 U1403 ( .A(n263), .ZN(n262) );
  INV_X1 U1404 ( .A(n1420), .ZN(n263) );
  INV_X1 U1405 ( .A(n1460), .ZN(n333) );
  NAND2_X1 U1406 ( .A1(n186), .A2(n149), .ZN(n145) );
  NAND2_X1 U1407 ( .A1(n214), .A2(n1395), .ZN(n201) );
  INV_X1 U1408 ( .A(n1410), .ZN(n334) );
  INV_X1 U1409 ( .A(n119), .ZN(n117) );
  INV_X1 U1410 ( .A(n1432), .ZN(n246) );
  XOR2_X1 U1411 ( .A(n339), .B(n89), .Z(product[16]) );
  NAND2_X1 U1412 ( .A1(n1460), .A2(n334), .ZN(n89) );
  NOR2_X1 U1413 ( .A1(n303), .A2(n1466), .ZN(n294) );
  NAND2_X1 U1414 ( .A1(n425), .A2(n290), .ZN(n82) );
  INV_X1 U1415 ( .A(n289), .ZN(n425) );
  XNOR2_X1 U1416 ( .A(n325), .B(n87), .ZN(product[18]) );
  NAND2_X1 U1417 ( .A1(n1436), .A2(n324), .ZN(n87) );
  OAI21_X1 U1418 ( .B1(n339), .B2(n326), .A(n327), .ZN(n325) );
  XNOR2_X1 U1419 ( .A(n332), .B(n88), .ZN(product[17]) );
  NAND2_X1 U1420 ( .A1(n1424), .A2(n331), .ZN(n88) );
  OAI21_X1 U1421 ( .B1(n339), .B2(n333), .A(n334), .ZN(n332) );
  XOR2_X1 U1422 ( .A(n352), .B(n91), .Z(product[14]) );
  NAND2_X1 U1423 ( .A1(n1412), .A2(n351), .ZN(n91) );
  AOI21_X1 U1424 ( .B1(n357), .B2(n435), .A(n354), .ZN(n352) );
  NAND2_X1 U1425 ( .A1(n1402), .A2(n346), .ZN(n90) );
  AOI21_X1 U1426 ( .B1(n357), .B2(n348), .A(n349), .ZN(n347) );
  INV_X1 U1427 ( .A(n284), .ZN(n424) );
  AOI21_X1 U1428 ( .B1(n1424), .B2(n1410), .A(n329), .ZN(n327) );
  INV_X1 U1429 ( .A(n331), .ZN(n329) );
  XOR2_X1 U1430 ( .A(n298), .B(n83), .Z(product[22]) );
  NAND2_X1 U1431 ( .A1(n426), .A2(n297), .ZN(n83) );
  AOI21_X1 U1432 ( .B1(n299), .B2(n319), .A(n300), .ZN(n298) );
  INV_X1 U1433 ( .A(n1466), .ZN(n426) );
  XOR2_X1 U1434 ( .A(n305), .B(n84), .Z(product[21]) );
  NAND2_X1 U1435 ( .A1(n302), .A2(n304), .ZN(n84) );
  AOI21_X1 U1436 ( .B1(n319), .B2(n306), .A(n1414), .ZN(n305) );
  OAI21_X1 U1437 ( .B1(n284), .B2(n290), .A(n285), .ZN(n283) );
  OAI21_X1 U1438 ( .B1(n1430), .B2(n318), .A(n313), .ZN(n311) );
  OAI21_X1 U1439 ( .B1(n217), .B2(n192), .A(n193), .ZN(n187) );
  INV_X1 U1440 ( .A(n358), .ZN(n357) );
  XOR2_X1 U1441 ( .A(n314), .B(n85), .Z(product[20]) );
  NAND2_X1 U1442 ( .A1(n1413), .A2(n313), .ZN(n85) );
  AOI21_X1 U1443 ( .B1(n319), .B2(n429), .A(n316), .ZN(n314) );
  NOR2_X1 U1444 ( .A1(n312), .A2(n317), .ZN(n310) );
  NOR2_X1 U1445 ( .A1(n216), .A2(n121), .ZN(n119) );
  NAND2_X1 U1446 ( .A1(n218), .A2(n240), .ZN(n216) );
  AOI21_X1 U1447 ( .B1(n1419), .B2(n249), .A(n250), .ZN(n248) );
  OAI21_X1 U1448 ( .B1(n251), .B2(n276), .A(n252), .ZN(n250) );
  AOI21_X1 U1449 ( .B1(n1405), .B2(n265), .A(n254), .ZN(n252) );
  NOR2_X1 U1450 ( .A1(n251), .A2(n275), .ZN(n249) );
  AOI21_X1 U1451 ( .B1(n215), .B2(n1395), .A(n206), .ZN(n202) );
  INV_X1 U1452 ( .A(n174), .ZN(n172) );
  OAI21_X1 U1453 ( .B1(n1466), .B2(n304), .A(n297), .ZN(n295) );
  OAI21_X1 U1454 ( .B1(n309), .B2(n301), .A(n304), .ZN(n300) );
  NAND2_X1 U1455 ( .A1(n348), .A2(n1402), .ZN(n341) );
  AOI21_X1 U1456 ( .B1(n349), .B2(n1402), .A(n344), .ZN(n342) );
  INV_X1 U1457 ( .A(n302), .ZN(n301) );
  OAI21_X1 U1458 ( .B1(n327), .B2(n323), .A(n324), .ZN(n322) );
  NOR2_X1 U1459 ( .A1(n192), .A2(n136), .ZN(n134) );
  INV_X1 U1460 ( .A(n217), .ZN(n215) );
  INV_X1 U1461 ( .A(n275), .ZN(n273) );
  NAND2_X1 U1462 ( .A1(n190), .A2(n177), .ZN(n175) );
  NAND2_X1 U1463 ( .A1(n1395), .A2(n1398), .ZN(n192) );
  NOR2_X1 U1464 ( .A1(n323), .A2(n326), .ZN(n321) );
  INV_X1 U1465 ( .A(n276), .ZN(n274) );
  INV_X1 U1466 ( .A(n267), .ZN(n265) );
  INV_X1 U1467 ( .A(n193), .ZN(n191) );
  INV_X1 U1468 ( .A(n290), .ZN(n288) );
  XNOR2_X1 U1469 ( .A(n319), .B(n86), .ZN(product[19]) );
  NAND2_X1 U1470 ( .A1(n429), .A2(n318), .ZN(n86) );
  INV_X1 U1471 ( .A(n317), .ZN(n429) );
  NAND2_X1 U1472 ( .A1(n240), .A2(n227), .ZN(n225) );
  INV_X1 U1473 ( .A(n318), .ZN(n316) );
  NAND2_X1 U1474 ( .A1(n173), .A2(n1407), .ZN(n160) );
  INV_X1 U1475 ( .A(n346), .ZN(n344) );
  INV_X1 U1476 ( .A(n256), .ZN(n254) );
  INV_X1 U1477 ( .A(n220), .ZN(n418) );
  XOR2_X1 U1478 ( .A(n374), .B(n95), .Z(product[10]) );
  NAND2_X1 U1479 ( .A1(n1404), .A2(n373), .ZN(n95) );
  AOI21_X1 U1480 ( .B1(n379), .B2(n1396), .A(n376), .ZN(n374) );
  AOI21_X1 U1481 ( .B1(n218), .B2(n241), .A(n219), .ZN(n217) );
  OAI21_X1 U1482 ( .B1(n230), .B2(n220), .A(n221), .ZN(n219) );
  XNOR2_X1 U1483 ( .A(n379), .B(n96), .ZN(product[9]) );
  NAND2_X1 U1484 ( .A1(n1396), .A2(n378), .ZN(n96) );
  NOR2_X1 U1485 ( .A1(n350), .A2(n355), .ZN(n348) );
  NOR2_X1 U1486 ( .A1(n561), .A2(n576), .ZN(n289) );
  XOR2_X1 U1487 ( .A(n198), .B(n73), .Z(product[32]) );
  NAND2_X1 U1488 ( .A1(n1398), .A2(n197), .ZN(n73) );
  AOI21_X1 U1489 ( .B1(n1398), .B2(n206), .A(n195), .ZN(n193) );
  INV_X1 U1490 ( .A(n197), .ZN(n195) );
  NAND2_X1 U1491 ( .A1(n1404), .A2(n1396), .ZN(n368) );
  AOI21_X1 U1492 ( .B1(n1404), .B2(n376), .A(n371), .ZN(n369) );
  XOR2_X1 U1493 ( .A(n181), .B(n72), .Z(product[33]) );
  NAND2_X1 U1494 ( .A1(n177), .A2(n180), .ZN(n72) );
  OAI21_X1 U1495 ( .B1(n217), .B2(n175), .A(n176), .ZN(n174) );
  AOI21_X1 U1496 ( .B1(n191), .B2(n177), .A(n178), .ZN(n176) );
  INV_X1 U1497 ( .A(n180), .ZN(n178) );
  XOR2_X1 U1498 ( .A(n244), .B(n77), .Z(product[28]) );
  NAND2_X1 U1499 ( .A1(n240), .A2(n243), .ZN(n77) );
  NOR2_X1 U1500 ( .A1(n229), .A2(n220), .ZN(n218) );
  NOR2_X1 U1501 ( .A1(n179), .A2(n151), .ZN(n149) );
  NAND2_X1 U1502 ( .A1(n134), .A2(n1403), .ZN(n121) );
  AOI21_X1 U1503 ( .B1(n187), .B2(n149), .A(n150), .ZN(n146) );
  AOI21_X1 U1504 ( .B1(n174), .B2(n1407), .A(n165), .ZN(n161) );
  AOI21_X1 U1505 ( .B1(n215), .B2(n134), .A(n135), .ZN(n131) );
  AOI21_X1 U1506 ( .B1(n241), .B2(n227), .A(n228), .ZN(n226) );
  INV_X1 U1507 ( .A(n230), .ZN(n228) );
  INV_X1 U1508 ( .A(n120), .ZN(n118) );
  NAND2_X1 U1509 ( .A1(n629), .A2(n646), .ZN(n318) );
  NAND2_X1 U1510 ( .A1(n533), .A2(n546), .ZN(n276) );
  NAND2_X1 U1511 ( .A1(n593), .A2(n610), .ZN(n304) );
  INV_X1 U1512 ( .A(n380), .ZN(n379) );
  NAND2_X1 U1513 ( .A1(n521), .A2(n532), .ZN(n267) );
  NAND2_X1 U1514 ( .A1(n693), .A2(n706), .ZN(n346) );
  NAND2_X1 U1515 ( .A1(n509), .A2(n520), .ZN(n256) );
  NAND2_X1 U1516 ( .A1(n611), .A2(n628), .ZN(n313) );
  NAND2_X1 U1517 ( .A1(n647), .A2(n662), .ZN(n324) );
  NAND2_X1 U1518 ( .A1(n547), .A2(n560), .ZN(n285) );
  NAND2_X1 U1519 ( .A1(n577), .A2(n592), .ZN(n297) );
  NOR2_X1 U1520 ( .A1(n361), .A2(n364), .ZN(n359) );
  OAI21_X1 U1521 ( .B1(n361), .B2(n365), .A(n362), .ZN(n360) );
  INV_X1 U1522 ( .A(n179), .ZN(n177) );
  INV_X1 U1523 ( .A(n229), .ZN(n227) );
  NAND2_X1 U1524 ( .A1(n149), .A2(n1401), .ZN(n136) );
  NAND2_X1 U1525 ( .A1(n1407), .A2(n1397), .ZN(n151) );
  INV_X1 U1526 ( .A(n242), .ZN(n240) );
  INV_X1 U1527 ( .A(n243), .ZN(n241) );
  INV_X1 U1528 ( .A(n208), .ZN(n206) );
  INV_X1 U1529 ( .A(n378), .ZN(n376) );
  XOR2_X1 U1530 ( .A(n366), .B(n94), .Z(product[11]) );
  NAND2_X1 U1531 ( .A1(n437), .A2(n365), .ZN(n94) );
  INV_X1 U1532 ( .A(n364), .ZN(n437) );
  XNOR2_X1 U1533 ( .A(n357), .B(n92), .ZN(product[13]) );
  NAND2_X1 U1534 ( .A1(n435), .A2(n356), .ZN(n92) );
  INV_X1 U1535 ( .A(n355), .ZN(n435) );
  XNOR2_X1 U1536 ( .A(n363), .B(n93), .ZN(product[12]) );
  OAI21_X1 U1537 ( .B1(n366), .B2(n364), .A(n365), .ZN(n363) );
  NAND2_X1 U1538 ( .A1(n436), .A2(n362), .ZN(n93) );
  INV_X1 U1539 ( .A(n361), .ZN(n436) );
  NAND2_X1 U1540 ( .A1(n119), .A2(n1400), .ZN(n108) );
  INV_X1 U1541 ( .A(n356), .ZN(n354) );
  INV_X1 U1542 ( .A(n373), .ZN(n371) );
  NAND2_X1 U1543 ( .A1(n441), .A2(n387), .ZN(n98) );
  INV_X1 U1544 ( .A(n386), .ZN(n441) );
  NAND2_X1 U1545 ( .A1(n1403), .A2(n126), .ZN(n68) );
  XNOR2_X1 U1546 ( .A(n385), .B(n97), .ZN(product[8]) );
  NAND2_X1 U1547 ( .A1(n1408), .A2(n384), .ZN(n97) );
  XOR2_X1 U1548 ( .A(n157), .B(n70), .Z(product[35]) );
  NAND2_X1 U1549 ( .A1(n1397), .A2(n156), .ZN(n70) );
  OAI21_X1 U1550 ( .B1(n388), .B2(n386), .A(n387), .ZN(n385) );
  XOR2_X1 U1551 ( .A(n142), .B(n69), .Z(product[36]) );
  NAND2_X1 U1552 ( .A1(n1401), .A2(n141), .ZN(n69) );
  XOR2_X1 U1553 ( .A(n114), .B(n67), .Z(product[38]) );
  NAND2_X1 U1554 ( .A1(n1400), .A2(n113), .ZN(n67) );
  INV_X1 U1555 ( .A(n392), .ZN(n390) );
  XOR2_X1 U1556 ( .A(n168), .B(n71), .Z(product[34]) );
  NAND2_X1 U1557 ( .A1(n1407), .A2(n167), .ZN(n71) );
  OAI21_X1 U1558 ( .B1(n193), .B2(n136), .A(n137), .ZN(n135) );
  AOI21_X1 U1559 ( .B1(n150), .B2(n1401), .A(n139), .ZN(n137) );
  INV_X1 U1560 ( .A(n141), .ZN(n139) );
  OAI21_X1 U1561 ( .B1(n394), .B2(n396), .A(n395), .ZN(n393) );
  OAI21_X1 U1562 ( .B1(n217), .B2(n121), .A(n122), .ZN(n120) );
  AOI21_X1 U1563 ( .B1(n135), .B2(n1403), .A(n124), .ZN(n122) );
  INV_X1 U1564 ( .A(n126), .ZN(n124) );
  OAI21_X1 U1565 ( .B1(n151), .B2(n180), .A(n152), .ZN(n150) );
  AOI21_X1 U1566 ( .B1(n165), .B2(n1397), .A(n154), .ZN(n152) );
  INV_X1 U1567 ( .A(n156), .ZN(n154) );
  AOI21_X1 U1568 ( .B1(n385), .B2(n1408), .A(n382), .ZN(n380) );
  INV_X1 U1569 ( .A(n384), .ZN(n382) );
  NAND2_X1 U1570 ( .A1(n461), .A2(n466), .ZN(n180) );
  NAND2_X1 U1571 ( .A1(n741), .A2(n750), .ZN(n365) );
  NAND2_X1 U1572 ( .A1(n489), .A2(n498), .ZN(n230) );
  NAND2_X1 U1573 ( .A1(n719), .A2(n730), .ZN(n356) );
  AOI21_X1 U1574 ( .B1(n120), .B2(n1400), .A(n111), .ZN(n109) );
  INV_X1 U1575 ( .A(n113), .ZN(n111) );
  NAND2_X1 U1576 ( .A1(n499), .A2(n508), .ZN(n243) );
  NAND2_X1 U1577 ( .A1(n473), .A2(n480), .ZN(n208) );
  NAND2_X1 U1578 ( .A1(n467), .A2(n472), .ZN(n197) );
  NAND2_X1 U1579 ( .A1(n731), .A2(n740), .ZN(n362) );
  NAND2_X1 U1580 ( .A1(n481), .A2(n488), .ZN(n221) );
  NAND2_X1 U1581 ( .A1(n759), .A2(n766), .ZN(n378) );
  NAND2_X1 U1582 ( .A1(n751), .A2(n758), .ZN(n373) );
  INV_X1 U1583 ( .A(n167), .ZN(n165) );
  NAND2_X1 U1584 ( .A1(n443), .A2(n395), .ZN(n100) );
  INV_X1 U1585 ( .A(n394), .ZN(n443) );
  NAND2_X1 U1586 ( .A1(n1399), .A2(n392), .ZN(n99) );
  NAND2_X1 U1587 ( .A1(n446), .A2(n407), .ZN(n103) );
  INV_X1 U1588 ( .A(n406), .ZN(n446) );
  XOR2_X1 U1589 ( .A(n102), .B(n404), .Z(product[3]) );
  NAND2_X1 U1590 ( .A1(n445), .A2(n403), .ZN(n102) );
  INV_X1 U1591 ( .A(n402), .ZN(n445) );
  OAI21_X1 U1592 ( .B1(n402), .B2(n404), .A(n403), .ZN(n401) );
  NAND2_X1 U1593 ( .A1(n830), .A2(n448), .ZN(n113) );
  AOI21_X1 U1594 ( .B1(n1409), .B2(n401), .A(n398), .ZN(n396) );
  INV_X1 U1595 ( .A(n400), .ZN(n398) );
  INV_X1 U1596 ( .A(n448), .ZN(n449) );
  INV_X1 U1597 ( .A(n478), .ZN(n479) );
  INV_X1 U1598 ( .A(n544), .ZN(n545) );
  NAND2_X1 U1599 ( .A1(n1028), .A2(n1009), .ZN(n407) );
  XNOR2_X1 U1600 ( .A(n937), .B(n865), .ZN(n627) );
  OR2_X1 U1601 ( .A1(n937), .A2(n865), .ZN(n626) );
  NAND2_X1 U1602 ( .A1(n457), .A2(n460), .ZN(n167) );
  NAND2_X1 U1603 ( .A1(n767), .A2(n772), .ZN(n384) );
  NAND2_X1 U1604 ( .A1(n779), .A2(n782), .ZN(n392) );
  NAND2_X1 U1605 ( .A1(n453), .A2(n456), .ZN(n156) );
  NAND2_X1 U1606 ( .A1(n452), .A2(n451), .ZN(n141) );
  NAND2_X1 U1607 ( .A1(n450), .A2(n449), .ZN(n126) );
  NAND2_X1 U1608 ( .A1(n783), .A2(n786), .ZN(n395) );
  NAND2_X1 U1609 ( .A1(n773), .A2(n778), .ZN(n387) );
  INV_X1 U1610 ( .A(n405), .ZN(n404) );
  OAI21_X1 U1611 ( .B1(n406), .B2(n409), .A(n407), .ZN(n405) );
  XNOR2_X1 U1612 ( .A(n101), .B(n401), .ZN(product[4]) );
  NAND2_X1 U1613 ( .A1(n1409), .A2(n400), .ZN(n101) );
  OAI22_X1 U1614 ( .A1(n1429), .A2(n1237), .B1(n1236), .B2(n3), .ZN(n1028) );
  OAI22_X1 U1615 ( .A1(n42), .A2(n1094), .B1(n40), .B2(n1093), .ZN(n478) );
  OAI22_X1 U1616 ( .A1(n24), .A2(n1157), .B1(n22), .B2(n1156), .ZN(n544) );
  OAI22_X1 U1617 ( .A1(n29), .A2(n1136), .B1(n28), .B2(n1135), .ZN(n518) );
  OAI22_X1 U1618 ( .A1(n18), .A2(n1178), .B1(n16), .B2(n1177), .ZN(n574) );
  OAI22_X1 U1619 ( .A1(n1445), .A2(n1199), .B1(n10), .B2(n1198), .ZN(n608) );
  OAI22_X1 U1620 ( .A1(n36), .A2(n1115), .B1(n33), .B2(n1114), .ZN(n496) );
  OAI22_X1 U1621 ( .A1(n1434), .A2(n1073), .B1(n45), .B2(n1072), .ZN(n464) );
  OAI22_X1 U1622 ( .A1(n1423), .A2(n1067), .B1(n51), .B2(n1066), .ZN(n865) );
  OAI22_X1 U1623 ( .A1(n1448), .A2(n1143), .B1(n28), .B2(n1142), .ZN(n937) );
  INV_X1 U1624 ( .A(n793), .ZN(n850) );
  OAI22_X1 U1625 ( .A1(n60), .A2(n1032), .B1(n58), .B2(n1031), .ZN(n831) );
  AOI21_X1 U1626 ( .B1(n54), .B2(n52), .A(n1051), .ZN(n793) );
  OAI22_X1 U1627 ( .A1(n17), .A2(n1195), .B1(n15), .B2(n1194), .ZN(n987) );
  OAI22_X1 U1628 ( .A1(n60), .A2(n1034), .B1(n58), .B2(n1033), .ZN(n833) );
  OAI22_X1 U1629 ( .A1(n1445), .A2(n1215), .B1(n9), .B2(n1214), .ZN(n1006) );
  OAI22_X1 U1630 ( .A1(n1429), .A2(n1234), .B1(n1233), .B2(n3), .ZN(n1025) );
  AND2_X1 U1631 ( .A1(n1449), .A2(n812), .ZN(n989) );
  OAI22_X1 U1632 ( .A1(n1445), .A2(n1216), .B1(n9), .B2(n1215), .ZN(n1007) );
  OAI22_X1 U1633 ( .A1(n1429), .A2(n1235), .B1(n1234), .B2(n3), .ZN(n1026) );
  AND2_X1 U1634 ( .A1(n1449), .A2(n794), .ZN(n869) );
  OAI22_X1 U1635 ( .A1(n6), .A2(n1223), .B1(n1222), .B2(n4), .ZN(n1014) );
  OAI22_X1 U1636 ( .A1(n41), .A2(n1109), .B1(n1108), .B2(n1421), .ZN(n905) );
  OAI22_X1 U1637 ( .A1(n11), .A2(n1213), .B1(n9), .B2(n1212), .ZN(n1004) );
  OAI22_X1 U1638 ( .A1(n17), .A2(n1194), .B1(n15), .B2(n1193), .ZN(n986) );
  OAI22_X1 U1639 ( .A1(n5), .A2(n1232), .B1(n1231), .B2(n3), .ZN(n1023) );
  OAI22_X1 U1640 ( .A1(n1434), .A2(n1089), .B1(n45), .B2(n1088), .ZN(n886) );
  OAI22_X1 U1641 ( .A1(n35), .A2(n1386), .B1(n33), .B2(n1126), .ZN(n922) );
  OAI22_X1 U1642 ( .A1(n41), .A2(n1108), .B1(n1107), .B2(n1421), .ZN(n904) );
  OAI22_X1 U1643 ( .A1(n11), .A2(n1200), .B1(n10), .B2(n1199), .ZN(n991) );
  OAI22_X1 U1644 ( .A1(n48), .A2(n1086), .B1(n1433), .B2(n1085), .ZN(n883) );
  OAI22_X1 U1645 ( .A1(n41), .A2(n1105), .B1(n1104), .B2(n1422), .ZN(n901) );
  OAI22_X1 U1646 ( .A1(n42), .A2(n1293), .B1(n1113), .B2(n40), .ZN(n823) );
  OAI22_X1 U1647 ( .A1(n41), .A2(n1112), .B1(n1111), .B2(n1422), .ZN(n908) );
  OR2_X1 U1648 ( .A1(n1449), .A2(n1293), .ZN(n1113) );
  OAI22_X1 U1649 ( .A1(n1423), .A2(n1061), .B1(n51), .B2(n1060), .ZN(n859) );
  OAI22_X1 U1650 ( .A1(n36), .A2(n1118), .B1(n34), .B2(n1117), .ZN(n913) );
  OAI22_X1 U1651 ( .A1(n29), .A2(n1137), .B1(n28), .B2(n1136), .ZN(n931) );
  OAI22_X1 U1652 ( .A1(n1423), .A2(n1063), .B1(n51), .B2(n1062), .ZN(n861) );
  OAI22_X1 U1653 ( .A1(n30), .A2(n1139), .B1(n28), .B2(n1138), .ZN(n933) );
  OAI22_X1 U1654 ( .A1(n24), .A2(n1158), .B1(n22), .B2(n1157), .ZN(n951) );
  OAI22_X1 U1655 ( .A1(n1423), .A2(n1065), .B1(n51), .B2(n1064), .ZN(n863) );
  OAI22_X1 U1656 ( .A1(n24), .A2(n1160), .B1(n22), .B2(n1159), .ZN(n953) );
  INV_X1 U1657 ( .A(n608), .ZN(n609) );
  OAI22_X1 U1658 ( .A1(n36), .A2(n1123), .B1(n33), .B2(n1122), .ZN(n918) );
  OAI22_X1 U1659 ( .A1(n1448), .A2(n1142), .B1(n28), .B2(n1141), .ZN(n936) );
  OAI22_X1 U1660 ( .A1(n11), .A2(n1431), .B1(n10), .B2(n1202), .ZN(n994) );
  OAI22_X1 U1661 ( .A1(n1429), .A2(n1222), .B1(n1221), .B2(n4), .ZN(n1013) );
  OAI22_X1 U1662 ( .A1(n30), .A2(n1146), .B1(n27), .B2(n1145), .ZN(n940) );
  OAI22_X1 U1663 ( .A1(n18), .A2(n1179), .B1(n16), .B2(n1178), .ZN(n971) );
  INV_X1 U1664 ( .A(n814), .ZN(n990) );
  OAI22_X1 U1665 ( .A1(n59), .A2(n1046), .B1(n57), .B2(n1045), .ZN(n845) );
  OAI22_X1 U1666 ( .A1(n1434), .A2(n1079), .B1(n45), .B2(n1078), .ZN(n876) );
  OAI22_X1 U1667 ( .A1(n36), .A2(n1117), .B1(n33), .B2(n1116), .ZN(n912) );
  OAI22_X1 U1668 ( .A1(n42), .A2(n1098), .B1(n40), .B2(n1097), .ZN(n894) );
  AOI21_X1 U1669 ( .B1(n6), .B2(n4), .A(n1219), .ZN(n817) );
  AOI21_X1 U1670 ( .B1(n42), .B2(n40), .A(n1093), .ZN(n799) );
  AOI21_X1 U1671 ( .B1(n36), .B2(n33), .A(n1114), .ZN(n802) );
  AOI21_X1 U1672 ( .B1(n12), .B2(n10), .A(n1198), .ZN(n814) );
  OAI22_X1 U1673 ( .A1(n1423), .A2(n1070), .B1(n51), .B2(n1069), .ZN(n868) );
  XNOR2_X1 U1674 ( .A(n1480), .B(n1482), .ZN(n1070) );
  OAI22_X1 U1675 ( .A1(n60), .A2(n1033), .B1(n58), .B2(n1032), .ZN(n832) );
  INV_X1 U1676 ( .A(n454), .ZN(n455) );
  NAND2_X1 U1677 ( .A1(n789), .A2(n828), .ZN(n403) );
  XNOR2_X1 U1678 ( .A(n37), .B(n1482), .ZN(n1112) );
  AND2_X1 U1679 ( .A1(n1483), .A2(n815), .ZN(n1009) );
  INV_X1 U1680 ( .A(n9), .ZN(n815) );
  INV_X1 U1681 ( .A(n811), .ZN(n970) );
  OAI22_X1 U1682 ( .A1(n59), .A2(n1044), .B1(n57), .B2(n1043), .ZN(n843) );
  AOI21_X1 U1683 ( .B1(n18), .B2(n16), .A(n1177), .ZN(n811) );
  OAI22_X1 U1684 ( .A1(n36), .A2(n1119), .B1(n34), .B2(n1118), .ZN(n914) );
  OAI22_X1 U1685 ( .A1(n42), .A2(n1100), .B1(n40), .B2(n1099), .ZN(n896) );
  OAI22_X1 U1686 ( .A1(n1447), .A2(n1138), .B1(n28), .B2(n1137), .ZN(n932) );
  OAI22_X1 U1687 ( .A1(n54), .A2(n1057), .B1(n52), .B2(n1056), .ZN(n855) );
  OAI22_X1 U1688 ( .A1(n1434), .A2(n1076), .B1(n1433), .B2(n1075), .ZN(n873)
         );
  OAI22_X1 U1689 ( .A1(n54), .A2(n1058), .B1(n52), .B2(n1057), .ZN(n856) );
  OAI22_X1 U1690 ( .A1(n60), .A2(n1039), .B1(n58), .B2(n1038), .ZN(n838) );
  OAI22_X1 U1691 ( .A1(n42), .A2(n1096), .B1(n40), .B2(n1095), .ZN(n892) );
  OAI22_X1 U1692 ( .A1(n1446), .A2(n1208), .B1(n9), .B2(n1207), .ZN(n999) );
  OAI22_X1 U1693 ( .A1(n35), .A2(n1132), .B1(n33), .B2(n1131), .ZN(n927) );
  OAI22_X1 U1694 ( .A1(n23), .A2(n1170), .B1(n1389), .B2(n1169), .ZN(n963) );
  OAI22_X1 U1695 ( .A1(n11), .A2(n1207), .B1(n10), .B2(n1206), .ZN(n998) );
  OAI22_X1 U1696 ( .A1(n5), .A2(n1226), .B1(n1225), .B2(n4), .ZN(n1017) );
  OAI22_X1 U1697 ( .A1(n23), .A2(n1169), .B1(n1389), .B2(n1168), .ZN(n962) );
  OAI22_X1 U1698 ( .A1(n12), .A2(n1204), .B1(n10), .B2(n1203), .ZN(n995) );
  OAI22_X1 U1699 ( .A1(n1090), .A2(n47), .B1(n45), .B2(n1089), .ZN(n887) );
  OAI22_X1 U1700 ( .A1(n35), .A2(n1128), .B1(n34), .B2(n1127), .ZN(n923) );
  OAI22_X1 U1701 ( .A1(n18), .A2(n1182), .B1(n16), .B2(n1181), .ZN(n974) );
  OAI22_X1 U1702 ( .A1(n1446), .A2(n1201), .B1(n10), .B2(n1200), .ZN(n992) );
  OAI22_X1 U1703 ( .A1(n35), .A2(n1125), .B1(n33), .B2(n1124), .ZN(n920) );
  OAI22_X1 U1704 ( .A1(n1434), .A2(n1084), .B1(n1433), .B2(n1083), .ZN(n881)
         );
  OAI22_X1 U1705 ( .A1(n41), .A2(n1103), .B1(n1102), .B2(n1422), .ZN(n899) );
  OAI22_X1 U1706 ( .A1(n30), .A2(n1141), .B1(n28), .B2(n1140), .ZN(n935) );
  OAI22_X1 U1707 ( .A1(n48), .A2(n1080), .B1(n1433), .B2(n1079), .ZN(n877) );
  OAI22_X1 U1708 ( .A1(n42), .A2(n1099), .B1(n40), .B2(n1098), .ZN(n895) );
  AND2_X1 U1709 ( .A1(n1450), .A2(n791), .ZN(n849) );
  OAI22_X1 U1710 ( .A1(n6), .A2(n1221), .B1(n1220), .B2(n4), .ZN(n1012) );
  OAI22_X1 U1711 ( .A1(n47), .A2(n1088), .B1(n45), .B2(n1087), .ZN(n885) );
  OAI22_X1 U1712 ( .A1(n18), .A2(n1181), .B1(n15), .B2(n1180), .ZN(n973) );
  OAI22_X1 U1713 ( .A1(n24), .A2(n1162), .B1(n22), .B2(n1161), .ZN(n955) );
  OAI22_X1 U1714 ( .A1(n54), .A2(n1059), .B1(n52), .B2(n1058), .ZN(n857) );
  OAI22_X1 U1715 ( .A1(n48), .A2(n1078), .B1(n1433), .B2(n1077), .ZN(n875) );
  OAI22_X1 U1716 ( .A1(n36), .A2(n1116), .B1(n33), .B2(n1115), .ZN(n911) );
  OAI22_X1 U1717 ( .A1(n48), .A2(n1083), .B1(n1433), .B2(n1082), .ZN(n880) );
  OAI22_X1 U1718 ( .A1(n1447), .A2(n1140), .B1(n28), .B2(n1139), .ZN(n934) );
  OAI22_X1 U1719 ( .A1(n24), .A2(n1159), .B1(n22), .B2(n1158), .ZN(n952) );
  OAI22_X1 U1720 ( .A1(n17), .A2(n1188), .B1(n15), .B2(n1187), .ZN(n980) );
  OAI22_X1 U1721 ( .A1(n35), .A2(n1131), .B1(n33), .B2(n1130), .ZN(n926) );
  OAI22_X1 U1722 ( .A1(n1447), .A2(n1150), .B1(n27), .B2(n1149), .ZN(n944) );
  OAI22_X1 U1723 ( .A1(n48), .A2(n1077), .B1(n1433), .B2(n1076), .ZN(n874) );
  INV_X1 U1724 ( .A(n496), .ZN(n497) );
  OAI22_X1 U1725 ( .A1(n18), .A2(n1385), .B1(n15), .B2(n1183), .ZN(n976) );
  OAI22_X1 U1726 ( .A1(n24), .A2(n1165), .B1(n22), .B2(n1164), .ZN(n958) );
  AND2_X1 U1727 ( .A1(n1483), .A2(n800), .ZN(n909) );
  OAI22_X1 U1728 ( .A1(n5), .A2(n1227), .B1(n1226), .B2(n4), .ZN(n1018) );
  OAI22_X1 U1729 ( .A1(n29), .A2(n1151), .B1(n27), .B2(n1150), .ZN(n945) );
  OAI22_X1 U1730 ( .A1(n36), .A2(n1122), .B1(n33), .B2(n1121), .ZN(n917) );
  OAI22_X1 U1731 ( .A1(n24), .A2(n1164), .B1(n22), .B2(n1163), .ZN(n957) );
  OAI22_X1 U1732 ( .A1(n1423), .A2(n1064), .B1(n51), .B2(n1063), .ZN(n862) );
  OAI22_X1 U1733 ( .A1(n59), .A2(n1045), .B1(n57), .B2(n1044), .ZN(n844) );
  OAI22_X1 U1734 ( .A1(n36), .A2(n1121), .B1(n33), .B2(n1120), .ZN(n916) );
  OAI22_X1 U1735 ( .A1(n35), .A2(n1129), .B1(n34), .B2(n1128), .ZN(n924) );
  OAI22_X1 U1736 ( .A1(n41), .A2(n1110), .B1(n1422), .B2(n1109), .ZN(n906) );
  OAI22_X1 U1737 ( .A1(n23), .A2(n1167), .B1(n1388), .B2(n1166), .ZN(n960) );
  OAI22_X1 U1738 ( .A1(n18), .A2(n1185), .B1(n16), .B2(n1184), .ZN(n977) );
  OAI22_X1 U1739 ( .A1(n23), .A2(n1166), .B1(n1388), .B2(n1165), .ZN(n959) );
  OAI22_X1 U1740 ( .A1(n30), .A2(n1147), .B1(n27), .B2(n1146), .ZN(n941) );
  OAI22_X1 U1741 ( .A1(n48), .A2(n1441), .B1(n45), .B2(n1086), .ZN(n884) );
  OAI22_X1 U1742 ( .A1(n1423), .A2(n1068), .B1(n51), .B2(n1067), .ZN(n866) );
  OAI22_X1 U1743 ( .A1(n29), .A2(n1144), .B1(n28), .B2(n1143), .ZN(n938) );
  OAI22_X1 U1744 ( .A1(n18), .A2(n1180), .B1(n16), .B2(n1179), .ZN(n972) );
  OAI22_X1 U1745 ( .A1(n59), .A2(n1047), .B1(n57), .B2(n1046), .ZN(n846) );
  OAI22_X1 U1746 ( .A1(n41), .A2(n1104), .B1(n1422), .B2(n1103), .ZN(n900) );
  OAI22_X1 U1747 ( .A1(n17), .A2(n1191), .B1(n15), .B2(n1190), .ZN(n983) );
  OAI22_X1 U1748 ( .A1(n1446), .A2(n1210), .B1(n9), .B2(n1209), .ZN(n1001) );
  OAI22_X1 U1749 ( .A1(n1448), .A2(n1153), .B1(n27), .B2(n1152), .ZN(n947) );
  OAI22_X1 U1750 ( .A1(n1445), .A2(n1211), .B1(n9), .B2(n1210), .ZN(n1002) );
  OAI22_X1 U1751 ( .A1(n17), .A2(n1192), .B1(n15), .B2(n1191), .ZN(n984) );
  OAI22_X1 U1752 ( .A1(n23), .A2(n1173), .B1(n1389), .B2(n1172), .ZN(n966) );
  OAI22_X1 U1753 ( .A1(n17), .A2(n1187), .B1(n15), .B2(n1186), .ZN(n979) );
  OAI22_X1 U1754 ( .A1(n23), .A2(n1168), .B1(n1389), .B2(n1167), .ZN(n961) );
  INV_X1 U1755 ( .A(n817), .ZN(n1010) );
  OAI22_X1 U1756 ( .A1(n59), .A2(n1048), .B1(n57), .B2(n1047), .ZN(n847) );
  OAI22_X1 U1757 ( .A1(n35), .A2(n1124), .B1(n34), .B2(n1123), .ZN(n919) );
  OAI22_X1 U1758 ( .A1(n1446), .A2(n1212), .B1(n9), .B2(n1211), .ZN(n1003) );
  OAI22_X1 U1759 ( .A1(n23), .A2(n1174), .B1(n1389), .B2(n1173), .ZN(n967) );
  OAI22_X1 U1760 ( .A1(n18), .A2(n1186), .B1(n16), .B2(n1185), .ZN(n978) );
  OAI22_X1 U1761 ( .A1(n1429), .A2(n1224), .B1(n1223), .B2(n4), .ZN(n1015) );
  OAI22_X1 U1762 ( .A1(n1447), .A2(n1148), .B1(n27), .B2(n1147), .ZN(n942) );
  OAI22_X1 U1763 ( .A1(n18), .A2(n1183), .B1(n16), .B2(n1182), .ZN(n975) );
  OAI22_X1 U1764 ( .A1(n35), .A2(n1126), .B1(n34), .B2(n1125), .ZN(n921) );
  OAI22_X1 U1765 ( .A1(n1448), .A2(n1145), .B1(n27), .B2(n1144), .ZN(n939) );
  OAI22_X1 U1766 ( .A1(n11), .A2(n1214), .B1(n9), .B2(n1213), .ZN(n1005) );
  AND2_X1 U1767 ( .A1(n1449), .A2(n809), .ZN(n969) );
  OAI22_X1 U1768 ( .A1(n1429), .A2(n1233), .B1(n1232), .B2(n3), .ZN(n1024) );
  OAI22_X1 U1769 ( .A1(n1434), .A2(n1082), .B1(n45), .B2(n1081), .ZN(n879) );
  OAI22_X1 U1770 ( .A1(n42), .A2(n1101), .B1(n40), .B2(n1100), .ZN(n897) );
  OAI22_X1 U1771 ( .A1(n36), .A2(n1120), .B1(n33), .B2(n1119), .ZN(n915) );
  OAI22_X1 U1772 ( .A1(n1423), .A2(n1062), .B1(n51), .B2(n1061), .ZN(n860) );
  OAI22_X1 U1773 ( .A1(n1434), .A2(n1081), .B1(n1433), .B2(n1080), .ZN(n878)
         );
  OAI22_X1 U1774 ( .A1(n59), .A2(n1043), .B1(n57), .B2(n1042), .ZN(n842) );
  OAI22_X1 U1775 ( .A1(n1445), .A2(n1205), .B1(n10), .B2(n1204), .ZN(n996) );
  OAI22_X1 U1776 ( .A1(n5), .A2(n1230), .B1(n1229), .B2(n3), .ZN(n1021) );
  INV_X1 U1777 ( .A(n574), .ZN(n575) );
  OAI22_X1 U1778 ( .A1(n42), .A2(n1102), .B1(n40), .B2(n1101), .ZN(n898) );
  AND2_X1 U1779 ( .A1(n1450), .A2(n803), .ZN(n929) );
  OAI22_X1 U1780 ( .A1(n1429), .A2(n1229), .B1(n1228), .B2(n3), .ZN(n1020) );
  OAI22_X1 U1781 ( .A1(n23), .A2(n1172), .B1(n1389), .B2(n1171), .ZN(n965) );
  AND2_X1 U1782 ( .A1(n1449), .A2(n797), .ZN(n889) );
  OAI22_X1 U1783 ( .A1(n1429), .A2(n1225), .B1(n1224), .B2(n4), .ZN(n1016) );
  OAI22_X1 U1784 ( .A1(n35), .A2(n1130), .B1(n34), .B2(n1129), .ZN(n925) );
  OAI22_X1 U1785 ( .A1(n1445), .A2(n1206), .B1(n10), .B2(n1205), .ZN(n997) );
  OAI22_X1 U1786 ( .A1(n1447), .A2(n1149), .B1(n27), .B2(n1148), .ZN(n943) );
  OAI22_X1 U1787 ( .A1(n41), .A2(n1111), .B1(n1110), .B2(n1421), .ZN(n907) );
  NAND2_X1 U1788 ( .A1(n1029), .A2(n829), .ZN(n409) );
  OAI22_X1 U1789 ( .A1(n42), .A2(n1097), .B1(n40), .B2(n1096), .ZN(n893) );
  OAI22_X1 U1790 ( .A1(n1446), .A2(n1209), .B1(n9), .B2(n1208), .ZN(n1000) );
  OAI22_X1 U1791 ( .A1(n23), .A2(n1171), .B1(n1389), .B2(n1170), .ZN(n964) );
  OAI22_X1 U1792 ( .A1(n17), .A2(n1189), .B1(n15), .B2(n1188), .ZN(n981) );
  OAI22_X1 U1793 ( .A1(n1434), .A2(n1074), .B1(n1433), .B2(n1073), .ZN(n871)
         );
  OAI22_X1 U1794 ( .A1(n1446), .A2(n1202), .B1(n10), .B2(n1201), .ZN(n993) );
  OAI22_X1 U1795 ( .A1(n41), .A2(n1107), .B1(n1106), .B2(n1421), .ZN(n903) );
  OAI22_X1 U1796 ( .A1(n1423), .A2(n1069), .B1(n51), .B2(n1068), .ZN(n867) );
  OAI22_X1 U1797 ( .A1(n54), .A2(n1056), .B1(n52), .B2(n1055), .ZN(n854) );
  OAI22_X1 U1798 ( .A1(n1434), .A2(n1075), .B1(n1433), .B2(n1074), .ZN(n872)
         );
  OAI22_X1 U1799 ( .A1(n60), .A2(n1037), .B1(n58), .B2(n1036), .ZN(n836) );
  OAI22_X1 U1800 ( .A1(n17), .A2(n1190), .B1(n15), .B2(n1189), .ZN(n982) );
  OAI22_X1 U1801 ( .A1(n5), .A2(n1228), .B1(n1227), .B2(n4), .ZN(n1019) );
  OAI22_X1 U1802 ( .A1(n1448), .A2(n1152), .B1(n27), .B2(n1151), .ZN(n946) );
  OAI22_X1 U1803 ( .A1(n1434), .A2(n1085), .B1(n1433), .B2(n1084), .ZN(n882)
         );
  OAI22_X1 U1804 ( .A1(n1423), .A2(n1066), .B1(n51), .B2(n1065), .ZN(n864) );
  OAI22_X1 U1805 ( .A1(n24), .A2(n1161), .B1(n22), .B2(n1160), .ZN(n954) );
  AND2_X1 U1806 ( .A1(n1450), .A2(n806), .ZN(n949) );
  OAI22_X1 U1807 ( .A1(n17), .A2(n1193), .B1(n15), .B2(n1192), .ZN(n985) );
  OAI22_X1 U1808 ( .A1(n1429), .A2(n1231), .B1(n1230), .B2(n3), .ZN(n1022) );
  OAI22_X1 U1809 ( .A1(n1429), .A2(n1220), .B1(n1219), .B2(n4), .ZN(n1011) );
  OAI22_X1 U1810 ( .A1(n41), .A2(n1106), .B1(n1105), .B2(n1422), .ZN(n902) );
  OAI22_X1 U1811 ( .A1(n24), .A2(n1163), .B1(n22), .B2(n1162), .ZN(n956) );
  NAND2_X1 U1812 ( .A1(n787), .A2(n788), .ZN(n400) );
  INV_X1 U1813 ( .A(n790), .ZN(n830) );
  AOI21_X1 U1814 ( .B1(n60), .B2(n58), .A(n1030), .ZN(n790) );
  OAI22_X1 U1815 ( .A1(n54), .A2(n1060), .B1(n52), .B2(n1059), .ZN(n858) );
  OAI22_X1 U1816 ( .A1(n59), .A2(n1041), .B1(n57), .B2(n1040), .ZN(n840) );
  INV_X1 U1817 ( .A(n518), .ZN(n519) );
  OAI22_X1 U1818 ( .A1(n54), .A2(n1054), .B1(n52), .B2(n1053), .ZN(n852) );
  OAI22_X1 U1819 ( .A1(n60), .A2(n1035), .B1(n58), .B2(n1034), .ZN(n834) );
  INV_X1 U1820 ( .A(n464), .ZN(n465) );
  INV_X1 U1821 ( .A(n15), .ZN(n812) );
  OR2_X1 U1822 ( .A1(n1483), .A2(n1290), .ZN(n1050) );
  OR2_X1 U1823 ( .A1(n1450), .A2(n1297), .ZN(n1197) );
  OR2_X1 U1824 ( .A1(n1483), .A2(n1296), .ZN(n1176) );
  OR2_X1 U1825 ( .A1(n1450), .A2(n1294), .ZN(n1134) );
  OR2_X1 U1826 ( .A1(n1449), .A2(n1295), .ZN(n1155) );
  INV_X1 U1827 ( .A(n1480), .ZN(n1291) );
  OR2_X1 U1828 ( .A1(n1483), .A2(n1292), .ZN(n1092) );
  OAI22_X1 U1829 ( .A1(n54), .A2(n1055), .B1(n52), .B2(n1054), .ZN(n853) );
  OAI22_X1 U1830 ( .A1(n60), .A2(n1036), .B1(n58), .B2(n1035), .ZN(n835) );
  INV_X1 U1831 ( .A(n799), .ZN(n890) );
  OAI22_X1 U1832 ( .A1(n59), .A2(n1042), .B1(n57), .B2(n1041), .ZN(n841) );
  INV_X1 U1833 ( .A(n808), .ZN(n950) );
  AOI21_X1 U1834 ( .B1(n24), .B2(n22), .A(n1156), .ZN(n808) );
  OAI22_X1 U1835 ( .A1(n60), .A2(n1038), .B1(n58), .B2(n1037), .ZN(n837) );
  OAI22_X1 U1836 ( .A1(n42), .A2(n1095), .B1(n40), .B2(n1094), .ZN(n891) );
  INV_X1 U1837 ( .A(n802), .ZN(n910) );
  OAI22_X1 U1838 ( .A1(n59), .A2(n1040), .B1(n57), .B2(n1039), .ZN(n839) );
  INV_X1 U1839 ( .A(n805), .ZN(n930) );
  AOI21_X1 U1840 ( .B1(n29), .B2(n28), .A(n1135), .ZN(n805) );
  OAI22_X1 U1841 ( .A1(n54), .A2(n1053), .B1(n52), .B2(n1052), .ZN(n851) );
  INV_X1 U1842 ( .A(n796), .ZN(n870) );
  AOI21_X1 U1843 ( .B1(n48), .B2(n45), .A(n1072), .ZN(n796) );
  INV_X1 U1844 ( .A(n57), .ZN(n791) );
  INV_X1 U1845 ( .A(n1389), .ZN(n809) );
  INV_X1 U1846 ( .A(n1421), .ZN(n800) );
  INV_X1 U1847 ( .A(n27), .ZN(n806) );
  INV_X1 U1848 ( .A(n1281), .ZN(n794) );
  INV_X1 U1849 ( .A(n34), .ZN(n803) );
  INV_X1 U1850 ( .A(n45), .ZN(n797) );
  AND2_X1 U1851 ( .A1(n1483), .A2(a[0]), .ZN(product[0]) );
  OAI22_X1 U1852 ( .A1(n11), .A2(n1298), .B1(n1218), .B2(n10), .ZN(n828) );
  OR2_X1 U1853 ( .A1(n1483), .A2(n1298), .ZN(n1218) );
  INV_X1 U1854 ( .A(n7), .ZN(n1298) );
  OAI22_X1 U1855 ( .A1(n1429), .A2(n1299), .B1(n1239), .B2(n4), .ZN(n829) );
  OR2_X1 U1856 ( .A1(n1483), .A2(n1299), .ZN(n1239) );
  OAI22_X1 U1857 ( .A1(n5), .A2(n1238), .B1(n1237), .B2(n3), .ZN(n1029) );
  XNOR2_X1 U1858 ( .A(n1479), .B(n1254), .ZN(n1065) );
  XNOR2_X1 U1859 ( .A(n1479), .B(n1255), .ZN(n1066) );
  XNOR2_X1 U1860 ( .A(n1479), .B(n1249), .ZN(n1060) );
  XNOR2_X1 U1861 ( .A(n1479), .B(n1477), .ZN(n1061) );
  XNOR2_X1 U1862 ( .A(n1479), .B(n1244), .ZN(n1055) );
  XNOR2_X1 U1863 ( .A(n1479), .B(n1475), .ZN(n1067) );
  XNOR2_X1 U1864 ( .A(n1479), .B(n1245), .ZN(n1056) );
  XNOR2_X1 U1865 ( .A(n1479), .B(n1257), .ZN(n1068) );
  XNOR2_X1 U1866 ( .A(n1479), .B(n1474), .ZN(n1062) );
  OAI22_X1 U1867 ( .A1(n29), .A2(n1154), .B1(n27), .B2(n1153), .ZN(n948) );
  OAI22_X1 U1868 ( .A1(n30), .A2(n1295), .B1(n1155), .B2(n28), .ZN(n825) );
  XNOR2_X1 U1869 ( .A(n25), .B(n1449), .ZN(n1154) );
  OAI22_X1 U1870 ( .A1(n11), .A2(n1217), .B1(n9), .B2(n1216), .ZN(n1008) );
  OAI22_X1 U1871 ( .A1(n5), .A2(n1236), .B1(n1235), .B2(n3), .ZN(n1027) );
  XNOR2_X1 U1872 ( .A(n7), .B(n1449), .ZN(n1217) );
  XNOR2_X1 U1873 ( .A(n1479), .B(n1241), .ZN(n1052) );
  XNOR2_X1 U1874 ( .A(n1479), .B(n1240), .ZN(n1051) );
  XNOR2_X1 U1875 ( .A(n37), .B(n1250), .ZN(n1103) );
  XNOR2_X1 U1876 ( .A(n37), .B(n1251), .ZN(n1104) );
  XNOR2_X1 U1877 ( .A(n37), .B(n1244), .ZN(n1097) );
  XNOR2_X1 U1878 ( .A(n37), .B(n1258), .ZN(n1111) );
  XNOR2_X1 U1879 ( .A(n37), .B(n1246), .ZN(n1099) );
  XNOR2_X1 U1880 ( .A(n37), .B(n1247), .ZN(n1100) );
  XNOR2_X1 U1881 ( .A(n37), .B(n1255), .ZN(n1108) );
  XNOR2_X1 U1882 ( .A(n37), .B(n1476), .ZN(n1109) );
  XNOR2_X1 U1883 ( .A(n37), .B(n1254), .ZN(n1107) );
  XNOR2_X1 U1884 ( .A(n37), .B(n1472), .ZN(n1110) );
  XNOR2_X1 U1885 ( .A(n37), .B(n1252), .ZN(n1105) );
  XNOR2_X1 U1886 ( .A(n37), .B(n1248), .ZN(n1101) );
  XNOR2_X1 U1887 ( .A(n37), .B(n1245), .ZN(n1098) );
  XNOR2_X1 U1888 ( .A(n37), .B(n1253), .ZN(n1106) );
  XNOR2_X1 U1889 ( .A(n1440), .B(n1243), .ZN(n1096) );
  XNOR2_X1 U1890 ( .A(n1440), .B(n1241), .ZN(n1094) );
  XNOR2_X1 U1891 ( .A(n37), .B(n1249), .ZN(n1102) );
  XNOR2_X1 U1892 ( .A(n1440), .B(n1242), .ZN(n1095) );
  XNOR2_X1 U1893 ( .A(n1440), .B(n1240), .ZN(n1093) );
  OAI22_X1 U1894 ( .A1(n35), .A2(n1133), .B1(n33), .B2(n1132), .ZN(n928) );
  OAI22_X1 U1895 ( .A1(n36), .A2(n1294), .B1(n1134), .B2(n33), .ZN(n824) );
  XNOR2_X1 U1896 ( .A(n1443), .B(n1449), .ZN(n1133) );
  OAI22_X1 U1897 ( .A1(n17), .A2(n1196), .B1(n15), .B2(n1195), .ZN(n988) );
  OAI22_X1 U1898 ( .A1(n18), .A2(n1297), .B1(n1197), .B2(n15), .ZN(n827) );
  XNOR2_X1 U1899 ( .A(n1435), .B(n1450), .ZN(n1196) );
  XNOR2_X1 U1900 ( .A(n1480), .B(n1252), .ZN(n1063) );
  XNOR2_X1 U1901 ( .A(n1480), .B(n1258), .ZN(n1069) );
  XNOR2_X1 U1902 ( .A(n1480), .B(n1248), .ZN(n1059) );
  XNOR2_X1 U1903 ( .A(n1480), .B(n1253), .ZN(n1064) );
  XNOR2_X1 U1904 ( .A(n1439), .B(n1242), .ZN(n1053) );
  XNOR2_X1 U1905 ( .A(n1439), .B(n1243), .ZN(n1054) );
  XNOR2_X1 U1906 ( .A(n1439), .B(n1246), .ZN(n1057) );
  XNOR2_X1 U1907 ( .A(n1439), .B(n1247), .ZN(n1058) );
  XNOR2_X1 U1908 ( .A(n25), .B(n1241), .ZN(n1136) );
  XNOR2_X1 U1909 ( .A(n1255), .B(n43), .ZN(n1087) );
  XNOR2_X1 U1910 ( .A(n43), .B(n1475), .ZN(n1088) );
  XNOR2_X1 U1911 ( .A(n43), .B(n1252), .ZN(n1084) );
  XNOR2_X1 U1912 ( .A(n43), .B(n1253), .ZN(n1085) );
  XNOR2_X1 U1913 ( .A(n25), .B(n1248), .ZN(n1143) );
  XNOR2_X1 U1914 ( .A(n25), .B(n1251), .ZN(n1146) );
  XNOR2_X1 U1915 ( .A(n25), .B(n1242), .ZN(n1137) );
  XNOR2_X1 U1916 ( .A(n25), .B(n1249), .ZN(n1144) );
  XNOR2_X1 U1917 ( .A(n25), .B(n1252), .ZN(n1147) );
  XNOR2_X1 U1918 ( .A(n25), .B(n1243), .ZN(n1138) );
  XNOR2_X1 U1919 ( .A(n43), .B(n1249), .ZN(n1081) );
  XNOR2_X1 U1920 ( .A(n43), .B(n1477), .ZN(n1082) );
  XNOR2_X1 U1921 ( .A(n43), .B(n1248), .ZN(n1080) );
  XNOR2_X1 U1922 ( .A(n1444), .B(n1241), .ZN(n1073) );
  XNOR2_X1 U1923 ( .A(n25), .B(n1477), .ZN(n1145) );
  XNOR2_X1 U1924 ( .A(n43), .B(n1471), .ZN(n1089) );
  XNOR2_X1 U1925 ( .A(n43), .B(n1246), .ZN(n1078) );
  XNOR2_X1 U1926 ( .A(n25), .B(n1256), .ZN(n1151) );
  XNOR2_X1 U1927 ( .A(n43), .B(n1247), .ZN(n1079) );
  XNOR2_X1 U1928 ( .A(n25), .B(n1472), .ZN(n1152) );
  XNOR2_X1 U1929 ( .A(n1444), .B(n1242), .ZN(n1074) );
  XNOR2_X1 U1930 ( .A(n43), .B(n1254), .ZN(n1086) );
  XNOR2_X1 U1931 ( .A(n1444), .B(n1243), .ZN(n1075) );
  XNOR2_X1 U1932 ( .A(n43), .B(n1258), .ZN(n1090) );
  XNOR2_X1 U1933 ( .A(n25), .B(n1253), .ZN(n1148) );
  XNOR2_X1 U1934 ( .A(n43), .B(n1251), .ZN(n1083) );
  XNOR2_X1 U1935 ( .A(n25), .B(n1247), .ZN(n1142) );
  XNOR2_X1 U1936 ( .A(n25), .B(n1244), .ZN(n1139) );
  XNOR2_X1 U1937 ( .A(n25), .B(n1245), .ZN(n1140) );
  XNOR2_X1 U1938 ( .A(n25), .B(n1246), .ZN(n1141) );
  XNOR2_X1 U1939 ( .A(n25), .B(n1254), .ZN(n1149) );
  XNOR2_X1 U1940 ( .A(n1444), .B(n1244), .ZN(n1076) );
  XNOR2_X1 U1941 ( .A(n25), .B(n1255), .ZN(n1150) );
  XNOR2_X1 U1942 ( .A(n25), .B(n1258), .ZN(n1153) );
  XNOR2_X1 U1943 ( .A(n1444), .B(n1245), .ZN(n1077) );
  XNOR2_X1 U1944 ( .A(n55), .B(n1256), .ZN(n1046) );
  XNOR2_X1 U1945 ( .A(n55), .B(n1257), .ZN(n1047) );
  XNOR2_X1 U1946 ( .A(n55), .B(n1255), .ZN(n1045) );
  XNOR2_X1 U1947 ( .A(n13), .B(n1241), .ZN(n1178) );
  XNOR2_X1 U1948 ( .A(n13), .B(n1242), .ZN(n1179) );
  XNOR2_X1 U1949 ( .A(n1435), .B(n1243), .ZN(n1180) );
  XNOR2_X1 U1950 ( .A(n19), .B(n1244), .ZN(n1160) );
  XNOR2_X1 U1951 ( .A(n19), .B(n1245), .ZN(n1161) );
  XNOR2_X1 U1952 ( .A(n1443), .B(n1249), .ZN(n1123) );
  XNOR2_X1 U1953 ( .A(n1443), .B(n1477), .ZN(n1124) );
  XNOR2_X1 U1954 ( .A(n1435), .B(n1252), .ZN(n1189) );
  XNOR2_X1 U1955 ( .A(n55), .B(n1258), .ZN(n1048) );
  XNOR2_X1 U1956 ( .A(n7), .B(n1246), .ZN(n1204) );
  XNOR2_X1 U1957 ( .A(n31), .B(n1474), .ZN(n1125) );
  XNOR2_X1 U1958 ( .A(n31), .B(n1252), .ZN(n1126) );
  XNOR2_X1 U1959 ( .A(n13), .B(n1247), .ZN(n1184) );
  XNOR2_X1 U1960 ( .A(n1443), .B(n1245), .ZN(n1119) );
  XNOR2_X1 U1961 ( .A(n1437), .B(n1244), .ZN(n1034) );
  XNOR2_X1 U1962 ( .A(n1435), .B(n1248), .ZN(n1185) );
  XNOR2_X1 U1963 ( .A(n19), .B(n1241), .ZN(n1157) );
  XNOR2_X1 U1964 ( .A(n1443), .B(n1246), .ZN(n1120) );
  XNOR2_X1 U1965 ( .A(n13), .B(n1245), .ZN(n1182) );
  XNOR2_X1 U1966 ( .A(n1437), .B(n1246), .ZN(n1036) );
  XNOR2_X1 U1967 ( .A(n55), .B(n1247), .ZN(n1037) );
  XNOR2_X1 U1968 ( .A(n55), .B(n1253), .ZN(n1043) );
  XNOR2_X1 U1969 ( .A(n55), .B(n1254), .ZN(n1044) );
  XNOR2_X1 U1970 ( .A(n19), .B(n1250), .ZN(n1166) );
  XNOR2_X1 U1971 ( .A(n13), .B(n1246), .ZN(n1183) );
  XNOR2_X1 U1972 ( .A(n19), .B(n1473), .ZN(n1167) );
  XNOR2_X1 U1973 ( .A(n55), .B(n1252), .ZN(n1042) );
  XNOR2_X1 U1974 ( .A(n31), .B(n1243), .ZN(n1117) );
  XNOR2_X1 U1975 ( .A(n1443), .B(n1244), .ZN(n1118) );
  XNOR2_X1 U1976 ( .A(n1435), .B(n1253), .ZN(n1190) );
  XNOR2_X1 U1977 ( .A(n7), .B(n1258), .ZN(n1216) );
  XNOR2_X1 U1978 ( .A(n7), .B(n1247), .ZN(n1205) );
  XNOR2_X1 U1979 ( .A(n1443), .B(n1242), .ZN(n1116) );
  XNOR2_X1 U1980 ( .A(n7), .B(n1241), .ZN(n1199) );
  XNOR2_X1 U1981 ( .A(n7), .B(n1242), .ZN(n1200) );
  XNOR2_X1 U1982 ( .A(n19), .B(n1249), .ZN(n1165) );
  XNOR2_X1 U1983 ( .A(n7), .B(n1245), .ZN(n1203) );
  XNOR2_X1 U1984 ( .A(n19), .B(n1246), .ZN(n1162) );
  XNOR2_X1 U1985 ( .A(n55), .B(n1473), .ZN(n1041) );
  XNOR2_X1 U1986 ( .A(n19), .B(n1247), .ZN(n1163) );
  XNOR2_X1 U1987 ( .A(n31), .B(n1254), .ZN(n1128) );
  XNOR2_X1 U1988 ( .A(n31), .B(n1255), .ZN(n1129) );
  XNOR2_X1 U1989 ( .A(n19), .B(n1242), .ZN(n1158) );
  XNOR2_X1 U1990 ( .A(n7), .B(n1244), .ZN(n1202) );
  XNOR2_X1 U1991 ( .A(n31), .B(n1253), .ZN(n1127) );
  XNOR2_X1 U1992 ( .A(n7), .B(n1472), .ZN(n1215) );
  XNOR2_X1 U1993 ( .A(n55), .B(n1250), .ZN(n1040) );
  XNOR2_X1 U1994 ( .A(n7), .B(n1255), .ZN(n1213) );
  XNOR2_X1 U1995 ( .A(n1443), .B(n1247), .ZN(n1121) );
  XNOR2_X1 U1996 ( .A(n7), .B(n1475), .ZN(n1214) );
  XNOR2_X1 U1997 ( .A(n19), .B(n1243), .ZN(n1159) );
  XNOR2_X1 U1998 ( .A(n1443), .B(n1258), .ZN(n1132) );
  XNOR2_X1 U1999 ( .A(n1435), .B(n1249), .ZN(n1186) );
  XNOR2_X1 U2000 ( .A(n7), .B(n1248), .ZN(n1206) );
  XNOR2_X1 U2001 ( .A(n1435), .B(n1477), .ZN(n1187) );
  XNOR2_X1 U2002 ( .A(n19), .B(n1252), .ZN(n1168) );
  XNOR2_X1 U2003 ( .A(n7), .B(n1243), .ZN(n1201) );
  XNOR2_X1 U2004 ( .A(n1435), .B(n1473), .ZN(n1188) );
  XNOR2_X1 U2005 ( .A(n1443), .B(n1256), .ZN(n1130) );
  XNOR2_X1 U2006 ( .A(n19), .B(n1255), .ZN(n1171) );
  XNOR2_X1 U2007 ( .A(n1435), .B(n1258), .ZN(n1195) );
  XNOR2_X1 U2008 ( .A(n19), .B(n1476), .ZN(n1172) );
  XNOR2_X1 U2009 ( .A(n1443), .B(n1241), .ZN(n1115) );
  XNOR2_X1 U2010 ( .A(n19), .B(n1253), .ZN(n1169) );
  XNOR2_X1 U2011 ( .A(n55), .B(n1248), .ZN(n1038) );
  XNOR2_X1 U2012 ( .A(n1437), .B(n1245), .ZN(n1035) );
  XNOR2_X1 U2013 ( .A(n1443), .B(n1471), .ZN(n1131) );
  XNOR2_X1 U2014 ( .A(n1435), .B(n1254), .ZN(n1191) );
  XNOR2_X1 U2015 ( .A(n1435), .B(n1244), .ZN(n1181) );
  XNOR2_X1 U2016 ( .A(n1435), .B(n1255), .ZN(n1192) );
  XNOR2_X1 U2017 ( .A(n19), .B(n1257), .ZN(n1173) );
  XNOR2_X1 U2018 ( .A(n1443), .B(n1248), .ZN(n1122) );
  XNOR2_X1 U2019 ( .A(n7), .B(n1249), .ZN(n1207) );
  XNOR2_X1 U2020 ( .A(n7), .B(n1477), .ZN(n1208) );
  XNOR2_X1 U2021 ( .A(n7), .B(n1251), .ZN(n1209) );
  XNOR2_X1 U2022 ( .A(n1435), .B(n1256), .ZN(n1193) );
  XNOR2_X1 U2023 ( .A(n7), .B(n1252), .ZN(n1210) );
  XNOR2_X1 U2024 ( .A(n7), .B(n1253), .ZN(n1211) );
  XNOR2_X1 U2025 ( .A(n19), .B(n1254), .ZN(n1170) );
  XNOR2_X1 U2026 ( .A(n1435), .B(n1257), .ZN(n1194) );
  XNOR2_X1 U2027 ( .A(n1416), .B(n1248), .ZN(n1164) );
  XNOR2_X1 U2028 ( .A(n1416), .B(n1258), .ZN(n1174) );
  XNOR2_X1 U2029 ( .A(n1437), .B(n1249), .ZN(n1039) );
  XNOR2_X1 U2030 ( .A(n1437), .B(n1243), .ZN(n1033) );
  XNOR2_X1 U2031 ( .A(n7), .B(n1254), .ZN(n1212) );
  XNOR2_X1 U2032 ( .A(n1437), .B(n1242), .ZN(n1032) );
  XNOR2_X1 U2033 ( .A(n1437), .B(n1241), .ZN(n1031) );
  BUF_X1 U2034 ( .A(n1285), .Z(n27) );
  BUF_X1 U2035 ( .A(n1284), .Z(n33) );
  XNOR2_X1 U2036 ( .A(n25), .B(n1468), .ZN(n1135) );
  XNOR2_X1 U2037 ( .A(n1444), .B(n1468), .ZN(n1072) );
  XNOR2_X1 U2038 ( .A(n7), .B(n1469), .ZN(n1198) );
  XNOR2_X1 U2039 ( .A(n1435), .B(n1240), .ZN(n1177) );
  XNOR2_X1 U2040 ( .A(n19), .B(n1468), .ZN(n1156) );
  XNOR2_X1 U2041 ( .A(n1443), .B(n1469), .ZN(n1114) );
  XNOR2_X1 U2042 ( .A(n1437), .B(n1240), .ZN(n1030) );
  BUF_X1 U2043 ( .A(n1280), .Z(n58) );
  BUF_X1 U2044 ( .A(n1286), .Z(n22) );
  BUF_X1 U2045 ( .A(n1285), .Z(n28) );
  BUF_X1 U2046 ( .A(n1287), .Z(n16) );
  BUF_X1 U2047 ( .A(n1284), .Z(n34) );
  BUF_X1 U2048 ( .A(n1278), .Z(n12) );
  BUF_X1 U2049 ( .A(n1278), .Z(n11) );
  BUF_X1 U2050 ( .A(n1279), .Z(n5) );
  OAI22_X1 U2051 ( .A1(n1434), .A2(n1091), .B1(n1433), .B2(n1090), .ZN(n888)
         );
  XNOR2_X1 U2052 ( .A(n43), .B(n1449), .ZN(n1091) );
  INV_X1 U2053 ( .A(n37), .ZN(n1293) );
  OAI22_X1 U2054 ( .A1(n23), .A2(n1175), .B1(n1389), .B2(n1174), .ZN(n968) );
  OAI22_X1 U2055 ( .A1(n24), .A2(n1296), .B1(n1176), .B2(n22), .ZN(n826) );
  XNOR2_X1 U2056 ( .A(n1416), .B(n1450), .ZN(n1175) );
  OAI22_X1 U2057 ( .A1(n59), .A2(n1049), .B1(n57), .B2(n1048), .ZN(n848) );
  OAI22_X1 U2058 ( .A1(n60), .A2(n1290), .B1(n1050), .B2(n58), .ZN(n820) );
  XNOR2_X1 U2059 ( .A(n55), .B(n1450), .ZN(n1049) );
  INV_X1 U2060 ( .A(n25), .ZN(n1295) );
  INV_X1 U2061 ( .A(n1443), .ZN(n1294) );
  INV_X1 U2062 ( .A(n1435), .ZN(n1297) );
  INV_X1 U2063 ( .A(n1416), .ZN(n1296) );
  INV_X1 U2064 ( .A(n55), .ZN(n1290) );
  BUF_X1 U2065 ( .A(n1289), .Z(n3) );
  INV_X1 U2066 ( .A(n43), .ZN(n1292) );
  BUF_X1 U2067 ( .A(n1289), .Z(n4) );
  BUF_X1 U2068 ( .A(n1275), .Z(n30) );
  BUF_X1 U2069 ( .A(n1274), .Z(n36) );
  BUF_X1 U2070 ( .A(n1275), .Z(n29) );
  XNOR2_X1 U2071 ( .A(a[10]), .B(a[9]), .ZN(n1284) );
  XNOR2_X1 U2072 ( .A(a[13]), .B(a[14]), .ZN(n1282) );
  NAND2_X1 U2073 ( .A1(n1261), .A2(n1281), .ZN(n1271) );
  NAND2_X1 U2074 ( .A1(n1268), .A2(n1288), .ZN(n1278) );
  NAND2_X1 U2075 ( .A1(n1269), .A2(n1289), .ZN(n1279) );
  INV_X1 U2076 ( .A(n303), .ZN(n302) );
  XOR2_X1 U2077 ( .A(n347), .B(n90), .Z(product[15]) );
  XNOR2_X1 U2078 ( .A(n1452), .B(n1474), .ZN(n1230) );
  XNOR2_X1 U2079 ( .A(n1390), .B(n1252), .ZN(n1231) );
  XNOR2_X1 U2080 ( .A(n1), .B(n1247), .ZN(n1226) );
  XNOR2_X1 U2081 ( .A(n1390), .B(n1483), .ZN(n1238) );
  XNOR2_X1 U2082 ( .A(n1), .B(n1246), .ZN(n1225) );
  XNOR2_X1 U2083 ( .A(n1), .B(n1248), .ZN(n1227) );
  INV_X1 U2084 ( .A(n1), .ZN(n1299) );
  XNOR2_X1 U2085 ( .A(n1), .B(n1253), .ZN(n1232) );
  XNOR2_X1 U2086 ( .A(n1), .B(n1243), .ZN(n1222) );
  XNOR2_X1 U2087 ( .A(n1), .B(n1254), .ZN(n1233) );
  XNOR2_X1 U2088 ( .A(n1), .B(n1255), .ZN(n1234) );
  XNOR2_X1 U2089 ( .A(n1), .B(n1476), .ZN(n1235) );
  XNOR2_X1 U2090 ( .A(n1), .B(n1258), .ZN(n1237) );
  XNOR2_X1 U2091 ( .A(n1452), .B(n1471), .ZN(n1236) );
  XNOR2_X1 U2092 ( .A(n1), .B(n1250), .ZN(n1229) );
  XNOR2_X1 U2093 ( .A(n1), .B(n1242), .ZN(n1221) );
  XNOR2_X1 U2094 ( .A(n1), .B(n1244), .ZN(n1223) );
  XNOR2_X1 U2095 ( .A(n1), .B(n1249), .ZN(n1228) );
  XNOR2_X1 U2096 ( .A(n1), .B(n1245), .ZN(n1224) );
  XNOR2_X1 U2097 ( .A(n1), .B(n1241), .ZN(n1220) );
  XNOR2_X1 U2098 ( .A(n1), .B(n1469), .ZN(n1219) );
  OAI22_X1 U2099 ( .A1(n54), .A2(n1052), .B1(n52), .B2(n1051), .ZN(n454) );
  AOI21_X1 U2100 ( .B1(n321), .B2(n1387), .A(n1442), .ZN(n1481) );
  OAI21_X1 U2101 ( .B1(n1461), .B2(n108), .A(n109), .ZN(n107) );
  OAI21_X1 U2102 ( .B1(n1461), .B2(n117), .A(n118), .ZN(n116) );
  OAI21_X1 U2103 ( .B1(n1453), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U2104 ( .B1(n1453), .B2(n171), .A(n172), .ZN(n170) );
  OAI21_X1 U2105 ( .B1(n1453), .B2(n160), .A(n161), .ZN(n159) );
  OAI21_X1 U2106 ( .B1(n1453), .B2(n145), .A(n146), .ZN(n144) );
  OAI21_X1 U2107 ( .B1(n1453), .B2(n201), .A(n202), .ZN(n200) );
  OAI21_X1 U2108 ( .B1(n1453), .B2(n184), .A(n185), .ZN(n183) );
  OAI21_X1 U2109 ( .B1(n1432), .B2(n216), .A(n217), .ZN(n211) );
  OAI21_X1 U2110 ( .B1(n1432), .B2(n242), .A(n243), .ZN(n233) );
  OAI21_X1 U2111 ( .B1(n1432), .B2(n225), .A(n226), .ZN(n224) );
  NAND2_X1 U2112 ( .A1(n1267), .A2(n1287), .ZN(n1277) );
  XOR2_X1 U2113 ( .A(n103), .B(n409), .Z(product[2]) );
  XNOR2_X1 U2114 ( .A(a[18]), .B(a[17]), .ZN(n1280) );
  NAND2_X1 U2115 ( .A1(n663), .A2(n678), .ZN(n331) );
  OAI22_X1 U2116 ( .A1(n54), .A2(n1291), .B1(n1071), .B2(n52), .ZN(n821) );
  OR2_X1 U2117 ( .A1(n1483), .A2(n1291), .ZN(n1071) );
  OAI21_X1 U2118 ( .B1(n368), .B2(n380), .A(n369), .ZN(n367) );
  AOI21_X1 U2119 ( .B1(n367), .B2(n359), .A(n360), .ZN(n358) );
  INV_X1 U2120 ( .A(n367), .ZN(n366) );
  AOI21_X1 U2121 ( .B1(n321), .B2(n1462), .A(n322), .ZN(n320) );
  NOR2_X1 U2122 ( .A1(n66), .A2(n108), .ZN(n106) );
  NOR2_X1 U2123 ( .A1(n66), .A2(n117), .ZN(n115) );
  NOR2_X1 U2124 ( .A1(n66), .A2(n160), .ZN(n158) );
  NOR2_X1 U2125 ( .A1(n66), .A2(n130), .ZN(n128) );
  NOR2_X1 U2126 ( .A1(n66), .A2(n216), .ZN(n210) );
  NOR2_X1 U2127 ( .A1(n66), .A2(n201), .ZN(n199) );
  NOR2_X1 U2128 ( .A1(n66), .A2(n242), .ZN(n232) );
  NOR2_X1 U2129 ( .A1(n66), .A2(n145), .ZN(n143) );
  NOR2_X1 U2130 ( .A1(n66), .A2(n225), .ZN(n223) );
  NOR2_X1 U2131 ( .A1(n66), .A2(n184), .ZN(n182) );
  NOR2_X1 U2132 ( .A1(n66), .A2(n171), .ZN(n169) );
  NAND2_X1 U2133 ( .A1(n561), .A2(n576), .ZN(n290) );
  XNOR2_X1 U2134 ( .A(a[8]), .B(a[7]), .ZN(n1285) );
  XOR2_X1 U2135 ( .A(a[6]), .B(a[7]), .Z(n1266) );
  XNOR2_X1 U2136 ( .A(a[4]), .B(a[3]), .ZN(n1287) );
  XOR2_X1 U2137 ( .A(a[2]), .B(a[3]), .Z(n1268) );
  XOR2_X1 U2138 ( .A(a[4]), .B(a[5]), .Z(n1267) );
  XNOR2_X1 U2139 ( .A(a[6]), .B(a[5]), .ZN(n1286) );
  AOI21_X1 U2140 ( .B1(n1417), .B2(n106), .A(n107), .ZN(n105) );
  AOI21_X1 U2141 ( .B1(n1417), .B2(n115), .A(n116), .ZN(n114) );
  AOI21_X1 U2142 ( .B1(n64), .B2(n158), .A(n159), .ZN(n157) );
  AOI21_X1 U2143 ( .B1(n64), .B2(n128), .A(n129), .ZN(n127) );
  AOI21_X1 U2144 ( .B1(n1417), .B2(n143), .A(n144), .ZN(n142) );
  AOI21_X1 U2145 ( .B1(n64), .B2(n169), .A(n170), .ZN(n168) );
  AOI21_X1 U2146 ( .B1(n63), .B2(n199), .A(n200), .ZN(n198) );
  AOI21_X1 U2147 ( .B1(n1478), .B2(n210), .A(n211), .ZN(n209) );
  AOI21_X1 U2148 ( .B1(n64), .B2(n182), .A(n183), .ZN(n181) );
  XOR2_X1 U2149 ( .A(n127), .B(n68), .Z(product[37]) );
  XOR2_X1 U2150 ( .A(a[8]), .B(a[9]), .Z(n1265) );
  OAI21_X1 U2151 ( .B1(n320), .B2(n292), .A(n293), .ZN(n291) );
  XOR2_X1 U2152 ( .A(a[14]), .B(a[15]), .Z(n1262) );
  NOR2_X1 U2153 ( .A1(n289), .A2(n284), .ZN(n282) );
  XOR2_X1 U2154 ( .A(a[18]), .B(a[19]), .Z(n1260) );
  OAI22_X1 U2155 ( .A1(n1434), .A2(n1292), .B1(n1092), .B2(n1433), .ZN(n822)
         );
  OAI21_X1 U2156 ( .B1(n350), .B2(n356), .A(n351), .ZN(n349) );
  NAND2_X1 U2157 ( .A1(n707), .A2(n718), .ZN(n351) );
  XOR2_X1 U2158 ( .A(a[12]), .B(a[13]), .Z(n1263) );
  XOR2_X1 U2159 ( .A(a[16]), .B(a[17]), .Z(n1261) );
  AOI21_X1 U2160 ( .B1(n63), .B2(n223), .A(n224), .ZN(n222) );
  AOI21_X1 U2161 ( .B1(n64), .B2(n269), .A(n270), .ZN(n268) );
  AOI21_X1 U2162 ( .B1(n64), .B2(n232), .A(n233), .ZN(n231) );
  XNOR2_X1 U2163 ( .A(n63), .B(n82), .ZN(product[23]) );
  AOI21_X1 U2164 ( .B1(n1478), .B2(n245), .A(n246), .ZN(n244) );
  AOI21_X1 U2165 ( .B1(n1478), .B2(n258), .A(n259), .ZN(n257) );
  AOI21_X1 U2166 ( .B1(n1478), .B2(n425), .A(n288), .ZN(n286) );
  AOI21_X1 U2167 ( .B1(n1478), .B2(n278), .A(n1419), .ZN(n277) );
  XOR2_X1 U2168 ( .A(a[11]), .B(a[10]), .Z(n1264) );
  XNOR2_X1 U2169 ( .A(a[12]), .B(a[11]), .ZN(n1283) );
  XNOR2_X1 U2170 ( .A(a[1]), .B(a[2]), .ZN(n1288) );
  XOR2_X1 U2171 ( .A(a[1]), .B(a[0]), .Z(n1269) );
  XOR2_X1 U2172 ( .A(n388), .B(n98), .Z(product[7]) );
  XNOR2_X1 U2173 ( .A(n99), .B(n393), .ZN(product[6]) );
  AOI21_X1 U2174 ( .B1(n1399), .B2(n393), .A(n390), .ZN(n388) );
  XOR2_X1 U2175 ( .A(n100), .B(n396), .Z(product[5]) );
endmodule


module datapath_DW_mult_tc_12 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n4, n5, n6, n7, n9, n10, n11, n12, n13, n15, n16, n17, n18, n19,
         n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34, n35, n36, n37,
         n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n51, n52, n53, n54,
         n55, n58, n59, n60, n61, n63, n64, n65, n67, n68, n69, n70, n71, n72,
         n73, n82, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n105, n106, n107, n108, n109,
         n111, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n124, n126, n127, n128, n129, n130, n131, n134, n135, n136, n137,
         n139, n141, n142, n143, n144, n145, n146, n149, n150, n151, n152,
         n154, n156, n157, n158, n159, n160, n161, n165, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n190, n191, n192, n193,
         n195, n197, n198, n199, n200, n201, n202, n206, n208, n209, n210,
         n211, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n240, n241, n242, n243, n244, n245, n246, n248, n249, n250, n251,
         n252, n254, n256, n257, n258, n259, n260, n261, n262, n263, n267,
         n268, n269, n270, n271, n273, n274, n275, n276, n277, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n331, n332, n333, n334, n339, n340, n341, n342, n344, n346,
         n347, n348, n349, n350, n351, n352, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n371, n373, n374, n376, n378, n379, n380, n382, n384, n385, n386,
         n387, n388, n390, n392, n393, n394, n395, n396, n398, n400, n401,
         n402, n403, n404, n405, n406, n407, n409, n418, n424, n426, n428,
         n430, n434, n435, n436, n437, n441, n443, n445, n446, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n793, n794, n796, n797, n799, n800, n802, n803, n805, n806,
         n808, n809, n811, n812, n814, n815, n817, n818, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1489, n1490, n1491, n1492;
  assign product[39] = n105;

  FA_X1 U488 ( .A(n831), .B(n454), .CI(n850), .CO(n450), .S(n451) );
  FA_X1 U489 ( .A(n455), .B(n832), .CI(n458), .CO(n452), .S(n453) );
  FA_X1 U491 ( .A(n462), .B(n833), .CI(n459), .CO(n456), .S(n457) );
  FA_X1 U492 ( .A(n851), .B(n464), .CI(n870), .CO(n458), .S(n459) );
  FA_X1 U493 ( .A(n463), .B(n470), .CI(n468), .CO(n460), .S(n461) );
  FA_X1 U494 ( .A(n834), .B(n852), .CI(n465), .CO(n462), .S(n463) );
  FA_X1 U496 ( .A(n474), .B(n471), .CI(n469), .CO(n466), .S(n467) );
  FA_X1 U497 ( .A(n478), .B(n871), .CI(n476), .CO(n468), .S(n469) );
  FA_X1 U498 ( .A(n853), .B(n835), .CI(n890), .CO(n470), .S(n471) );
  FA_X1 U499 ( .A(n475), .B(n477), .CI(n482), .CO(n472), .S(n473) );
  FA_X1 U500 ( .A(n486), .B(n479), .CI(n484), .CO(n474), .S(n475) );
  FA_X1 U501 ( .A(n836), .B(n854), .CI(n872), .CO(n476), .S(n477) );
  FA_X1 U503 ( .A(n490), .B(n492), .CI(n483), .CO(n480), .S(n481) );
  FA_X1 U504 ( .A(n485), .B(n494), .CI(n487), .CO(n482), .S(n483) );
  FA_X1 U505 ( .A(n855), .B(n496), .CI(n873), .CO(n484), .S(n485) );
  FA_X1 U506 ( .A(n891), .B(n837), .CI(n910), .CO(n486), .S(n487) );
  FA_X1 U507 ( .A(n500), .B(n493), .CI(n491), .CO(n488), .S(n489) );
  FA_X1 U508 ( .A(n495), .B(n504), .CI(n502), .CO(n490), .S(n491) );
  FA_X1 U509 ( .A(n497), .B(n874), .CI(n506), .CO(n492), .S(n493) );
  FA_X1 U510 ( .A(n892), .B(n856), .CI(n838), .CO(n494), .S(n495) );
  FA_X1 U512 ( .A(n510), .B(n503), .CI(n501), .CO(n498), .S(n499) );
  FA_X1 U513 ( .A(n507), .B(n505), .CI(n512), .CO(n500), .S(n501) );
  FA_X1 U514 ( .A(n516), .B(n893), .CI(n514), .CO(n502), .S(n503) );
  FA_X1 U515 ( .A(n857), .B(n911), .CI(n875), .CO(n504), .S(n505) );
  FA_X1 U516 ( .A(n518), .B(n839), .CI(n930), .CO(n506), .S(n507) );
  FA_X1 U517 ( .A(n522), .B(n513), .CI(n511), .CO(n508), .S(n509) );
  FA_X1 U519 ( .A(n528), .B(n530), .CI(n517), .CO(n512), .S(n513) );
  FA_X1 U520 ( .A(n840), .B(n858), .CI(n519), .CO(n514), .S(n515) );
  FA_X1 U521 ( .A(n912), .B(n876), .CI(n894), .CO(n516), .S(n517) );
  FA_X1 U523 ( .A(n523), .B(n525), .CI(n534), .CO(n520), .S(n521) );
  FA_X1 U524 ( .A(n527), .B(n538), .CI(n536), .CO(n522), .S(n523) );
  FA_X1 U526 ( .A(n877), .B(n895), .CI(n542), .CO(n526), .S(n527) );
  FA_X1 U527 ( .A(n859), .B(n931), .CI(n913), .CO(n528), .S(n529) );
  FA_X1 U528 ( .A(n544), .B(n841), .CI(n950), .CO(n530), .S(n531) );
  FA_X1 U529 ( .A(n535), .B(n537), .CI(n548), .CO(n532), .S(n533) );
  FA_X1 U530 ( .A(n539), .B(n552), .CI(n550), .CO(n534), .S(n535) );
  FA_X1 U531 ( .A(n541), .B(n554), .CI(n543), .CO(n536), .S(n537) );
  FA_X1 U532 ( .A(n558), .B(n545), .CI(n556), .CO(n538), .S(n539) );
  FA_X1 U533 ( .A(n896), .B(n932), .CI(n914), .CO(n540), .S(n541) );
  FA_X1 U534 ( .A(n842), .B(n878), .CI(n860), .CO(n542), .S(n543) );
  FA_X1 U536 ( .A(n562), .B(n551), .CI(n549), .CO(n546), .S(n547) );
  FA_X1 U537 ( .A(n553), .B(n566), .CI(n564), .CO(n548), .S(n549) );
  FA_X1 U538 ( .A(n559), .B(n557), .CI(n568), .CO(n550), .S(n551) );
  FA_X1 U539 ( .A(n570), .B(n572), .CI(n555), .CO(n552), .S(n553) );
  FA_X1 U540 ( .A(n879), .B(n915), .CI(n897), .CO(n554), .S(n555) );
  FA_X1 U541 ( .A(n861), .B(n951), .CI(n933), .CO(n556), .S(n557) );
  FA_X1 U542 ( .A(n574), .B(n843), .CI(n970), .CO(n558), .S(n559) );
  FA_X1 U544 ( .A(n567), .B(n582), .CI(n580), .CO(n562), .S(n563) );
  FA_X1 U545 ( .A(n584), .B(n573), .CI(n569), .CO(n564), .S(n565) );
  FA_X1 U546 ( .A(n586), .B(n588), .CI(n571), .CO(n566), .S(n567) );
  FA_X1 U547 ( .A(n575), .B(n898), .CI(n590), .CO(n568), .S(n569) );
  FA_X1 U548 ( .A(n844), .B(n916), .CI(n862), .CO(n570), .S(n571) );
  FA_X1 U549 ( .A(n952), .B(n880), .CI(n934), .CO(n572), .S(n573) );
  FA_X1 U551 ( .A(n594), .B(n581), .CI(n579), .CO(n576), .S(n577) );
  FA_X1 U552 ( .A(n583), .B(n598), .CI(n596), .CO(n578), .S(n579) );
  FA_X1 U553 ( .A(n600), .B(n591), .CI(n585), .CO(n580), .S(n581) );
  FA_X1 U554 ( .A(n587), .B(n602), .CI(n589), .CO(n582), .S(n583) );
  FA_X1 U555 ( .A(n606), .B(n917), .CI(n604), .CO(n584), .S(n585) );
  FA_X1 U556 ( .A(n881), .B(n935), .CI(n899), .CO(n586), .S(n587) );
  FA_X1 U557 ( .A(n608), .B(n953), .CI(n863), .CO(n588), .S(n589) );
  FA_X1 U558 ( .A(n845), .B(n971), .CI(n990), .CO(n590), .S(n591) );
  FA_X1 U560 ( .A(n599), .B(n616), .CI(n614), .CO(n594), .S(n595) );
  FA_X1 U561 ( .A(n618), .B(n603), .CI(n601), .CO(n596), .S(n597) );
  FA_X1 U562 ( .A(n605), .B(n620), .CI(n607), .CO(n598), .S(n599) );
  FA_X1 U563 ( .A(n626), .B(n624), .CI(n622), .CO(n600), .S(n601) );
  FA_X1 U564 ( .A(n918), .B(n936), .CI(n609), .CO(n602), .S(n603) );
  FA_X1 U565 ( .A(n954), .B(n864), .CI(n882), .CO(n604), .S(n605) );
  FA_X1 U566 ( .A(n900), .B(n846), .CI(n972), .CO(n606), .S(n607) );
  FA_X1 U568 ( .A(n630), .B(n615), .CI(n613), .CO(n610), .S(n611) );
  FA_X1 U569 ( .A(n617), .B(n634), .CI(n632), .CO(n612), .S(n613) );
  FA_X1 U570 ( .A(n636), .B(n621), .CI(n619), .CO(n614), .S(n615) );
  FA_X1 U571 ( .A(n623), .B(n638), .CI(n625), .CO(n616), .S(n617) );
  FA_X1 U572 ( .A(n642), .B(n627), .CI(n640), .CO(n618), .S(n619) );
  FA_X1 U573 ( .A(n955), .B(n973), .CI(n644), .CO(n620), .S(n621) );
  FA_X1 U574 ( .A(n991), .B(n901), .CI(n883), .CO(n622), .S(n623) );
  FA_X1 U575 ( .A(n919), .B(n847), .CI(n1010), .CO(n624), .S(n625) );
  FA_X1 U578 ( .A(n648), .B(n633), .CI(n631), .CO(n628), .S(n629) );
  FA_X1 U579 ( .A(n650), .B(n637), .CI(n635), .CO(n630), .S(n631) );
  FA_X1 U580 ( .A(n654), .B(n643), .CI(n652), .CO(n632), .S(n633) );
  FA_X1 U581 ( .A(n639), .B(n656), .CI(n641), .CO(n634), .S(n635) );
  FA_X1 U582 ( .A(n660), .B(n645), .CI(n658), .CO(n636), .S(n637) );
  FA_X1 U583 ( .A(n920), .B(n992), .CI(n974), .CO(n638), .S(n639) );
  FA_X1 U584 ( .A(n1011), .B(n956), .CI(n902), .CO(n640), .S(n641) );
  FA_X1 U585 ( .A(n866), .B(n938), .CI(n884), .CO(n642), .S(n643) );
  HA_X1 U586 ( .A(n848), .B(n820), .CO(n644), .S(n645) );
  FA_X1 U588 ( .A(n666), .B(n655), .CI(n653), .CO(n648), .S(n649) );
  FA_X1 U589 ( .A(n670), .B(n659), .CI(n668), .CO(n650), .S(n651) );
  FA_X1 U590 ( .A(n661), .B(n672), .CI(n657), .CO(n652), .S(n653) );
  FA_X1 U591 ( .A(n676), .B(n957), .CI(n674), .CO(n654), .S(n655) );
  FA_X1 U592 ( .A(n921), .B(n975), .CI(n939), .CO(n656), .S(n657) );
  FA_X1 U593 ( .A(n867), .B(n993), .CI(n903), .CO(n658), .S(n659) );
  FA_X1 U594 ( .A(n1012), .B(n849), .CI(n885), .CO(n660), .S(n661) );
  FA_X1 U595 ( .A(n667), .B(n680), .CI(n665), .CO(n662), .S(n663) );
  FA_X1 U596 ( .A(n682), .B(n671), .CI(n669), .CO(n664), .S(n665) );
  FA_X1 U597 ( .A(n675), .B(n673), .CI(n684), .CO(n666), .S(n667) );
  FA_X1 U598 ( .A(n686), .B(n690), .CI(n688), .CO(n668), .S(n669) );
  FA_X1 U599 ( .A(n958), .B(n976), .CI(n677), .CO(n670), .S(n671) );
  FA_X1 U600 ( .A(n886), .B(n904), .CI(n922), .CO(n672), .S(n673) );
  FA_X1 U601 ( .A(n1013), .B(n940), .CI(n994), .CO(n674), .S(n675) );
  HA_X1 U602 ( .A(n821), .B(n868), .CO(n676), .S(n677) );
  FA_X1 U603 ( .A(n694), .B(n683), .CI(n681), .CO(n678), .S(n679) );
  FA_X1 U604 ( .A(n685), .B(n698), .CI(n696), .CO(n680), .S(n681) );
  FA_X1 U606 ( .A(n702), .B(n704), .CI(n700), .CO(n684), .S(n685) );
  FA_X1 U607 ( .A(n941), .B(n977), .CI(n959), .CO(n686), .S(n687) );
  FA_X1 U608 ( .A(n995), .B(n887), .CI(n923), .CO(n688), .S(n689) );
  FA_X1 U609 ( .A(n1014), .B(n869), .CI(n905), .CO(n690), .S(n691) );
  FA_X1 U610 ( .A(n697), .B(n708), .CI(n695), .CO(n692), .S(n693) );
  FA_X1 U611 ( .A(n710), .B(n703), .CI(n699), .CO(n694), .S(n695) );
  FA_X1 U612 ( .A(n701), .B(n714), .CI(n712), .CO(n696), .S(n697) );
  FA_X1 U613 ( .A(n716), .B(n996), .CI(n705), .CO(n698), .S(n699) );
  FA_X1 U614 ( .A(n1015), .B(n942), .CI(n978), .CO(n700), .S(n701) );
  FA_X1 U615 ( .A(n906), .B(n924), .CI(n960), .CO(n702), .S(n703) );
  HA_X1 U616 ( .A(n822), .B(n888), .CO(n704), .S(n705) );
  FA_X1 U617 ( .A(n711), .B(n720), .CI(n709), .CO(n706), .S(n707) );
  FA_X1 U618 ( .A(n713), .B(n715), .CI(n722), .CO(n708), .S(n709) );
  FA_X1 U619 ( .A(n724), .B(n726), .CI(n717), .CO(n710), .S(n711) );
  FA_X1 U620 ( .A(n961), .B(n979), .CI(n728), .CO(n712), .S(n713) );
  FA_X1 U621 ( .A(n907), .B(n997), .CI(n943), .CO(n714), .S(n715) );
  FA_X1 U622 ( .A(n925), .B(n889), .CI(n1016), .CO(n716), .S(n717) );
  FA_X1 U623 ( .A(n732), .B(n723), .CI(n721), .CO(n718), .S(n719) );
  FA_X1 U624 ( .A(n727), .B(n725), .CI(n734), .CO(n720), .S(n721) );
  FA_X1 U625 ( .A(n738), .B(n729), .CI(n736), .CO(n722), .S(n723) );
  FA_X1 U626 ( .A(n926), .B(n980), .CI(n944), .CO(n724), .S(n725) );
  FA_X1 U627 ( .A(n1017), .B(n962), .CI(n998), .CO(n726), .S(n727) );
  HA_X1 U628 ( .A(n908), .B(n823), .CO(n728), .S(n729) );
  FA_X1 U629 ( .A(n735), .B(n742), .CI(n733), .CO(n730), .S(n731) );
  FA_X1 U630 ( .A(n737), .B(n739), .CI(n744), .CO(n732), .S(n733) );
  FA_X1 U631 ( .A(n748), .B(n981), .CI(n746), .CO(n734), .S(n735) );
  FA_X1 U632 ( .A(n927), .B(n999), .CI(n963), .CO(n736), .S(n737) );
  FA_X1 U633 ( .A(n945), .B(n909), .CI(n1018), .CO(n738), .S(n739) );
  FA_X1 U634 ( .A(n752), .B(n745), .CI(n743), .CO(n740), .S(n741) );
  FA_X1 U635 ( .A(n754), .B(n756), .CI(n747), .CO(n742), .S(n743) );
  FA_X1 U636 ( .A(n964), .B(n1000), .CI(n749), .CO(n744), .S(n745) );
  FA_X1 U637 ( .A(n946), .B(n982), .CI(n1019), .CO(n746), .S(n747) );
  HA_X1 U638 ( .A(n824), .B(n928), .CO(n748), .S(n749) );
  FA_X1 U639 ( .A(n760), .B(n755), .CI(n753), .CO(n750), .S(n751) );
  FA_X1 U640 ( .A(n762), .B(n764), .CI(n757), .CO(n752), .S(n753) );
  FA_X1 U641 ( .A(n947), .B(n1001), .CI(n983), .CO(n754), .S(n755) );
  FA_X1 U642 ( .A(n965), .B(n929), .CI(n1020), .CO(n756), .S(n757) );
  FA_X1 U643 ( .A(n763), .B(n768), .CI(n761), .CO(n758), .S(n759) );
  FA_X1 U644 ( .A(n765), .B(n1021), .CI(n770), .CO(n760), .S(n761) );
  FA_X1 U645 ( .A(n966), .B(n984), .CI(n1002), .CO(n762), .S(n763) );
  HA_X1 U646 ( .A(n825), .B(n948), .CO(n764), .S(n765) );
  FA_X1 U647 ( .A(n771), .B(n774), .CI(n769), .CO(n766), .S(n767) );
  FA_X1 U648 ( .A(n967), .B(n1003), .CI(n776), .CO(n768), .S(n769) );
  FA_X1 U649 ( .A(n985), .B(n949), .CI(n1022), .CO(n770), .S(n771) );
  FA_X1 U650 ( .A(n780), .B(n777), .CI(n775), .CO(n772), .S(n773) );
  FA_X1 U651 ( .A(n986), .B(n1023), .CI(n1004), .CO(n774), .S(n775) );
  HA_X1 U652 ( .A(n826), .B(n968), .CO(n776), .S(n777) );
  FA_X1 U653 ( .A(n784), .B(n987), .CI(n781), .CO(n778), .S(n779) );
  FA_X1 U654 ( .A(n1024), .B(n969), .CI(n1005), .CO(n780), .S(n781) );
  FA_X1 U655 ( .A(n1006), .B(n1025), .CI(n785), .CO(n782), .S(n783) );
  HA_X1 U656 ( .A(n827), .B(n988), .CO(n784), .S(n785) );
  FA_X1 U657 ( .A(n1026), .B(n989), .CI(n1007), .CO(n786), .S(n787) );
  HA_X1 U658 ( .A(n1008), .B(n1027), .CO(n788), .S(n789) );
  CLKBUF_X3 U1180 ( .A(n1275), .Z(n29) );
  BUF_X1 U1181 ( .A(n1275), .Z(n30) );
  CLKBUF_X2 U1182 ( .A(n1283), .Z(n39) );
  BUF_X1 U1183 ( .A(n1283), .Z(n40) );
  CLKBUF_X3 U1184 ( .A(n1274), .Z(n36) );
  AOI21_X1 U1185 ( .B1(n283), .B2(n249), .A(n250), .ZN(n1383) );
  BUF_X4 U1186 ( .A(a[1]), .Z(n1384) );
  CLKBUF_X1 U1187 ( .A(a[1]), .Z(n1) );
  CLKBUF_X3 U1188 ( .A(b[17]), .Z(n1385) );
  CLKBUF_X3 U1189 ( .A(n1270), .Z(n59) );
  CLKBUF_X1 U1190 ( .A(n37), .Z(n1386) );
  CLKBUF_X3 U1191 ( .A(b[7]), .Z(n1252) );
  BUF_X1 U1192 ( .A(n1278), .Z(n1387) );
  CLKBUF_X3 U1193 ( .A(b[12]), .Z(n1247) );
  OR2_X2 U1194 ( .A1(n751), .A2(n758), .ZN(n1388) );
  CLKBUF_X1 U1195 ( .A(n358), .Z(n1389) );
  BUF_X1 U1196 ( .A(n1279), .Z(n1390) );
  BUF_X1 U1197 ( .A(n1279), .Z(n1391) );
  CLKBUF_X2 U1198 ( .A(n1282), .Z(n46) );
  CLKBUF_X3 U1199 ( .A(b[15]), .Z(n1244) );
  CLKBUF_X3 U1200 ( .A(b[14]), .Z(n1245) );
  CLKBUF_X3 U1201 ( .A(b[16]), .Z(n1243) );
  CLKBUF_X3 U1202 ( .A(b[17]), .Z(n1242) );
  CLKBUF_X3 U1203 ( .A(b[4]), .Z(n1255) );
  BUF_X2 U1204 ( .A(b[19]), .Z(n1240) );
  BUF_X2 U1205 ( .A(b[1]), .Z(n1258) );
  CLKBUF_X3 U1206 ( .A(b[13]), .Z(n1246) );
  CLKBUF_X1 U1207 ( .A(b[0]), .Z(n61) );
  XOR2_X1 U1208 ( .A(n691), .B(n687), .Z(n1392) );
  XOR2_X1 U1209 ( .A(n689), .B(n1392), .Z(n683) );
  NAND2_X2 U1210 ( .A1(n689), .A2(n691), .ZN(n1393) );
  NAND2_X1 U1211 ( .A1(n687), .A2(n689), .ZN(n1394) );
  NAND2_X1 U1212 ( .A1(n691), .A2(n687), .ZN(n1395) );
  NAND3_X1 U1213 ( .A1(n1393), .A2(n1394), .A3(n1395), .ZN(n682) );
  CLKBUF_X3 U1214 ( .A(b[11]), .Z(n1248) );
  CLKBUF_X3 U1215 ( .A(b[2]), .Z(n1257) );
  CLKBUF_X3 U1216 ( .A(b[6]), .Z(n1253) );
  AND2_X1 U1217 ( .A1(n521), .A2(n532), .ZN(n1474) );
  BUF_X1 U1218 ( .A(n61), .Z(n1491) );
  BUF_X1 U1219 ( .A(n43), .Z(n1484) );
  OAI22_X1 U1220 ( .A1(n60), .A2(n1031), .B1(n58), .B2(n1030), .ZN(n448) );
  INV_X1 U1221 ( .A(n1474), .ZN(n267) );
  XOR2_X1 U1222 ( .A(n664), .B(n651), .Z(n1396) );
  XOR2_X1 U1223 ( .A(n649), .B(n1396), .Z(n647) );
  NAND2_X1 U1224 ( .A1(n649), .A2(n664), .ZN(n1397) );
  NAND2_X1 U1225 ( .A1(n649), .A2(n651), .ZN(n1398) );
  NAND2_X1 U1226 ( .A1(n664), .A2(n651), .ZN(n1399) );
  NAND3_X1 U1227 ( .A1(n1397), .A2(n1398), .A3(n1399), .ZN(n646) );
  OR2_X1 U1228 ( .A1(n473), .A2(n480), .ZN(n1400) );
  OR2_X1 U1229 ( .A1(n453), .A2(n456), .ZN(n1401) );
  OR2_X1 U1230 ( .A1(n467), .A2(n472), .ZN(n1402) );
  OR2_X1 U1231 ( .A1(n830), .A2(n448), .ZN(n1403) );
  OR2_X1 U1232 ( .A1(n452), .A2(n451), .ZN(n1404) );
  OR2_X1 U1233 ( .A1(n759), .A2(n766), .ZN(n1405) );
  OR2_X1 U1234 ( .A1(n450), .A2(n449), .ZN(n1406) );
  OR2_X1 U1235 ( .A1(n457), .A2(n460), .ZN(n1407) );
  OR2_X1 U1236 ( .A1(n767), .A2(n772), .ZN(n1408) );
  OR2_X1 U1237 ( .A1(n779), .A2(n782), .ZN(n1409) );
  OR2_X1 U1238 ( .A1(n787), .A2(n788), .ZN(n1410) );
  NOR2_X1 U1239 ( .A1(n561), .A2(n576), .ZN(n289) );
  OR2_X1 U1240 ( .A1(n1029), .A2(n829), .ZN(n1411) );
  NOR2_X1 U1241 ( .A1(n499), .A2(n508), .ZN(n242) );
  BUF_X1 U1242 ( .A(n248), .Z(n65) );
  CLKBUF_X1 U1243 ( .A(n1250), .Z(n1412) );
  XNOR2_X1 U1244 ( .A(n19), .B(n1250), .ZN(n1413) );
  CLKBUF_X3 U1245 ( .A(b[9]), .Z(n1250) );
  BUF_X2 U1246 ( .A(n1383), .Z(n1414) );
  INV_X1 U1247 ( .A(n1298), .ZN(n1415) );
  INV_X1 U1248 ( .A(n1241), .ZN(n1416) );
  INV_X2 U1249 ( .A(n1416), .ZN(n1417) );
  BUF_X1 U1250 ( .A(b[18]), .Z(n1241) );
  XNOR2_X1 U1251 ( .A(n13), .B(n1242), .ZN(n1418) );
  BUF_X2 U1252 ( .A(n1280), .Z(n1481) );
  CLKBUF_X1 U1253 ( .A(n1240), .Z(n1419) );
  BUF_X2 U1254 ( .A(n61), .Z(n1420) );
  BUF_X2 U1255 ( .A(n61), .Z(n1492) );
  CLKBUF_X1 U1256 ( .A(n1250), .Z(n1421) );
  BUF_X1 U1257 ( .A(n1287), .Z(n16) );
  CLKBUF_X1 U1258 ( .A(n1287), .Z(n15) );
  NOR2_X1 U1259 ( .A1(n593), .A2(n610), .ZN(n303) );
  XNOR2_X1 U1260 ( .A(n7), .B(n1245), .ZN(n1422) );
  XNOR2_X1 U1261 ( .A(n298), .B(n1423), .ZN(product[22]) );
  AND2_X1 U1262 ( .A1(n426), .A2(n297), .ZN(n1423) );
  AND2_X1 U1263 ( .A1(n679), .A2(n692), .ZN(n1469) );
  XNOR2_X1 U1264 ( .A(n1384), .B(n1240), .ZN(n1424) );
  XNOR2_X1 U1265 ( .A(n563), .B(n1425), .ZN(n561) );
  XNOR2_X1 U1266 ( .A(n578), .B(n565), .ZN(n1425) );
  INV_X1 U1267 ( .A(n1468), .ZN(n331) );
  CLKBUF_X2 U1268 ( .A(n1284), .Z(n33) );
  BUF_X1 U1269 ( .A(n1284), .Z(n34) );
  BUF_X2 U1270 ( .A(n1273), .Z(n42) );
  AND2_X1 U1271 ( .A1(n663), .A2(n678), .ZN(n1468) );
  XOR2_X1 U1272 ( .A(n529), .B(n540), .Z(n1426) );
  XOR2_X1 U1273 ( .A(n1426), .B(n531), .Z(n525) );
  NAND2_X1 U1274 ( .A1(n529), .A2(n540), .ZN(n1427) );
  NAND2_X1 U1275 ( .A1(n529), .A2(n531), .ZN(n1428) );
  NAND2_X1 U1276 ( .A1(n540), .A2(n531), .ZN(n1429) );
  NAND3_X1 U1277 ( .A1(n1427), .A2(n1428), .A3(n1429), .ZN(n524) );
  XOR2_X1 U1278 ( .A(n526), .B(n515), .Z(n1430) );
  XOR2_X1 U1279 ( .A(n1430), .B(n524), .Z(n511) );
  NAND2_X1 U1280 ( .A1(n526), .A2(n515), .ZN(n1431) );
  NAND2_X1 U1281 ( .A1(n526), .A2(n524), .ZN(n1432) );
  NAND2_X1 U1282 ( .A1(n515), .A2(n524), .ZN(n1433) );
  NAND3_X1 U1283 ( .A1(n1431), .A2(n1432), .A3(n1433), .ZN(n510) );
  CLKBUF_X2 U1284 ( .A(a[9]), .Z(n1435) );
  BUF_X1 U1285 ( .A(n1123), .Z(n1434) );
  CLKBUF_X1 U1286 ( .A(a[9]), .Z(n25) );
  OAI22_X1 U1287 ( .A1(n24), .A2(n1157), .B1(n1156), .B2(n1443), .ZN(n1436) );
  XNOR2_X1 U1288 ( .A(n1490), .B(n1255), .ZN(n1437) );
  XNOR2_X1 U1289 ( .A(n55), .B(n1258), .ZN(n1438) );
  BUF_X4 U1290 ( .A(a[19]), .Z(n55) );
  BUF_X1 U1291 ( .A(n1124), .Z(n1439) );
  CLKBUF_X1 U1292 ( .A(n37), .Z(n1440) );
  XNOR2_X1 U1293 ( .A(n55), .B(n1257), .ZN(n1441) );
  CLKBUF_X1 U1294 ( .A(n1419), .Z(n1442) );
  BUF_X1 U1295 ( .A(n1286), .Z(n1443) );
  CLKBUF_X1 U1296 ( .A(n31), .Z(n1444) );
  CLKBUF_X1 U1297 ( .A(n311), .Z(n1445) );
  CLKBUF_X1 U1298 ( .A(n1478), .Z(n1446) );
  CLKBUF_X1 U1299 ( .A(n320), .Z(n1447) );
  CLKBUF_X1 U1300 ( .A(n64), .Z(n1448) );
  BUF_X1 U1301 ( .A(n1286), .Z(n22) );
  XNOR2_X1 U1302 ( .A(n268), .B(n1449), .ZN(product[26]) );
  AND2_X1 U1303 ( .A1(n262), .A2(n267), .ZN(n1449) );
  NAND2_X1 U1304 ( .A1(n563), .A2(n578), .ZN(n1450) );
  NAND2_X1 U1305 ( .A1(n563), .A2(n565), .ZN(n1451) );
  NAND2_X1 U1306 ( .A1(n578), .A2(n565), .ZN(n1452) );
  NAND3_X1 U1307 ( .A1(n1450), .A2(n1451), .A3(n1452), .ZN(n560) );
  XNOR2_X1 U1308 ( .A(n286), .B(n1453), .ZN(product[24]) );
  AND2_X1 U1309 ( .A1(n424), .A2(n285), .ZN(n1453) );
  CLKBUF_X1 U1310 ( .A(n282), .Z(n1454) );
  NAND2_X2 U1311 ( .A1(n282), .A2(n249), .ZN(n1455) );
  XNOR2_X1 U1312 ( .A(n277), .B(n1456), .ZN(product[25]) );
  AND2_X1 U1313 ( .A1(n273), .A2(n276), .ZN(n1456) );
  OR2_X2 U1314 ( .A1(n693), .A2(n706), .ZN(n1457) );
  CLKBUF_X1 U1315 ( .A(n1414), .Z(n1458) );
  XNOR2_X1 U1316 ( .A(n1256), .B(n1484), .ZN(n1459) );
  OR2_X1 U1317 ( .A1(n312), .A2(n317), .ZN(n1460) );
  XNOR2_X1 U1318 ( .A(n257), .B(n1461), .ZN(product[27]) );
  AND2_X1 U1319 ( .A1(n1471), .A2(n256), .ZN(n1461) );
  NOR2_X1 U1320 ( .A1(n533), .A2(n546), .ZN(n275) );
  XNOR2_X1 U1321 ( .A(n595), .B(n1462), .ZN(n593) );
  XNOR2_X1 U1322 ( .A(n612), .B(n597), .ZN(n1462) );
  NOR2_X2 U1323 ( .A1(n707), .A2(n718), .ZN(n350) );
  NOR2_X2 U1324 ( .A1(n731), .A2(n740), .ZN(n361) );
  NAND2_X1 U1325 ( .A1(n595), .A2(n612), .ZN(n1463) );
  NAND2_X1 U1326 ( .A1(n595), .A2(n597), .ZN(n1464) );
  NAND2_X1 U1327 ( .A1(n612), .A2(n597), .ZN(n1465) );
  NAND3_X1 U1328 ( .A1(n1463), .A2(n1464), .A3(n1465), .ZN(n592) );
  OR2_X2 U1329 ( .A1(n679), .A2(n692), .ZN(n1466) );
  CLKBUF_X1 U1330 ( .A(n313), .Z(n1467) );
  BUF_X2 U1331 ( .A(n1282), .Z(n45) );
  XNOR2_X1 U1332 ( .A(n231), .B(n1470), .ZN(product[29]) );
  AND2_X1 U1333 ( .A1(n227), .A2(n230), .ZN(n1470) );
  OR2_X2 U1334 ( .A1(n509), .A2(n520), .ZN(n1471) );
  INV_X1 U1335 ( .A(n316), .ZN(n1472) );
  XNOR2_X1 U1336 ( .A(n222), .B(n1473), .ZN(product[30]) );
  AND2_X1 U1337 ( .A1(n418), .A2(n221), .ZN(n1473) );
  BUF_X2 U1338 ( .A(n1276), .Z(n23) );
  CLKBUF_X1 U1339 ( .A(n1285), .Z(n27) );
  BUF_X1 U1340 ( .A(n1285), .Z(n28) );
  NOR2_X1 U1341 ( .A1(n647), .A2(n662), .ZN(n323) );
  BUF_X2 U1342 ( .A(n1271), .Z(n53) );
  NAND2_X1 U1343 ( .A1(n509), .A2(n520), .ZN(n256) );
  CLKBUF_X3 U1344 ( .A(b[10]), .Z(n1249) );
  NOR2_X1 U1345 ( .A1(n547), .A2(n560), .ZN(n1475) );
  NOR2_X1 U1346 ( .A1(n547), .A2(n560), .ZN(n284) );
  NOR2_X1 U1347 ( .A1(n611), .A2(n628), .ZN(n1476) );
  BUF_X2 U1348 ( .A(n1272), .Z(n1477) );
  NOR2_X1 U1349 ( .A1(n611), .A2(n628), .ZN(n312) );
  CLKBUF_X1 U1350 ( .A(n1272), .Z(n47) );
  NAND2_X1 U1351 ( .A1(n1264), .A2(n1284), .ZN(n1274) );
  NOR2_X1 U1352 ( .A1(n577), .A2(n592), .ZN(n1478) );
  NOR2_X1 U1353 ( .A1(n577), .A2(n592), .ZN(n296) );
  BUF_X2 U1354 ( .A(n1276), .Z(n24) );
  OR2_X2 U1355 ( .A1(n663), .A2(n678), .ZN(n1479) );
  OR2_X1 U1356 ( .A1(n521), .A2(n532), .ZN(n1480) );
  BUF_X2 U1357 ( .A(n1272), .Z(n48) );
  NOR2_X1 U1358 ( .A1(n629), .A2(n646), .ZN(n317) );
  CLKBUF_X3 U1359 ( .A(b[5]), .Z(n1254) );
  BUF_X2 U1360 ( .A(n1273), .Z(n41) );
  NAND2_X1 U1361 ( .A1(n1260), .A2(n1280), .ZN(n1270) );
  BUF_X1 U1362 ( .A(n1280), .Z(n58) );
  AOI21_X1 U1363 ( .B1(n1479), .B2(n1469), .A(n1468), .ZN(n1482) );
  BUF_X1 U1364 ( .A(n43), .Z(n1483) );
  XNOR2_X1 U1365 ( .A(n305), .B(n1485), .ZN(product[21]) );
  AND2_X1 U1366 ( .A1(n302), .A2(n304), .ZN(n1485) );
  OAI21_X1 U1367 ( .B1(n1476), .B2(n318), .A(n313), .ZN(n311) );
  NAND2_X1 U1368 ( .A1(n218), .A2(n240), .ZN(n216) );
  XNOR2_X1 U1369 ( .A(n209), .B(n1486), .ZN(product[31]) );
  AND2_X1 U1370 ( .A1(n1400), .A2(n208), .ZN(n1486) );
  XNOR2_X1 U1371 ( .A(n244), .B(n1487), .ZN(product[28]) );
  AND2_X1 U1372 ( .A1(n240), .A2(n243), .ZN(n1487) );
  NAND2_X1 U1373 ( .A1(n629), .A2(n646), .ZN(n318) );
  NAND2_X1 U1374 ( .A1(n533), .A2(n546), .ZN(n276) );
  NOR2_X1 U1375 ( .A1(n461), .A2(n466), .ZN(n179) );
  NOR2_X1 U1376 ( .A1(n719), .A2(n730), .ZN(n355) );
  NOR2_X1 U1377 ( .A1(n741), .A2(n750), .ZN(n364) );
  NOR2_X1 U1378 ( .A1(n481), .A2(n488), .ZN(n220) );
  NAND2_X1 U1379 ( .A1(n473), .A2(n480), .ZN(n208) );
  NOR2_X1 U1380 ( .A1(n1028), .A2(n1009), .ZN(n406) );
  NOR2_X1 U1381 ( .A1(n773), .A2(n778), .ZN(n386) );
  NOR2_X1 U1382 ( .A1(n789), .A2(n828), .ZN(n402) );
  AND2_X1 U1383 ( .A1(n1411), .A2(n409), .ZN(product[1]) );
  BUF_X2 U1384 ( .A(n1281), .Z(n51) );
  BUF_X2 U1385 ( .A(n1278), .Z(n12) );
  BUF_X1 U1386 ( .A(n1279), .Z(n5) );
  BUF_X2 U1387 ( .A(n1270), .Z(n60) );
  NAND2_X1 U1388 ( .A1(n1261), .A2(n1281), .ZN(n1271) );
  BUF_X1 U1389 ( .A(a[15]), .Z(n43) );
  NAND2_X1 U1390 ( .A1(n1262), .A2(n1282), .ZN(n1272) );
  NAND2_X1 U1391 ( .A1(n214), .A2(n134), .ZN(n130) );
  NOR2_X1 U1392 ( .A1(n280), .A2(n260), .ZN(n258) );
  NOR2_X1 U1393 ( .A1(n280), .A2(n271), .ZN(n269) );
  INV_X1 U1394 ( .A(n186), .ZN(n184) );
  INV_X1 U1395 ( .A(n173), .ZN(n171) );
  NOR2_X1 U1396 ( .A1(n1455), .A2(n216), .ZN(n210) );
  NOR2_X1 U1397 ( .A1(n1455), .A2(n242), .ZN(n232) );
  NOR2_X1 U1398 ( .A1(n1455), .A2(n145), .ZN(n143) );
  NOR2_X1 U1399 ( .A1(n1455), .A2(n117), .ZN(n115) );
  NOR2_X1 U1400 ( .A1(n1455), .A2(n130), .ZN(n128) );
  NOR2_X1 U1401 ( .A1(n1455), .A2(n201), .ZN(n199) );
  NOR2_X1 U1402 ( .A1(n1455), .A2(n171), .ZN(n169) );
  NOR2_X1 U1403 ( .A1(n1455), .A2(n184), .ZN(n182) );
  INV_X1 U1404 ( .A(n1460), .ZN(n306) );
  INV_X1 U1405 ( .A(n281), .ZN(n279) );
  INV_X1 U1406 ( .A(n1455), .ZN(n245) );
  INV_X1 U1407 ( .A(n1447), .ZN(n319) );
  INV_X1 U1408 ( .A(n283), .ZN(n281) );
  NOR2_X1 U1409 ( .A1(n216), .A2(n175), .ZN(n173) );
  NOR2_X1 U1410 ( .A1(n216), .A2(n192), .ZN(n186) );
  INV_X1 U1411 ( .A(n340), .ZN(n339) );
  INV_X1 U1412 ( .A(n216), .ZN(n214) );
  NOR2_X1 U1413 ( .A1(n1460), .A2(n301), .ZN(n299) );
  OAI21_X1 U1414 ( .B1(n65), .B2(n216), .A(n213), .ZN(n211) );
  INV_X1 U1415 ( .A(n215), .ZN(n213) );
  OAI21_X1 U1416 ( .B1(n65), .B2(n242), .A(n243), .ZN(n233) );
  OAI21_X1 U1417 ( .B1(n1414), .B2(n184), .A(n185), .ZN(n183) );
  INV_X1 U1418 ( .A(n187), .ZN(n185) );
  OAI21_X1 U1419 ( .B1(n281), .B2(n260), .A(n261), .ZN(n259) );
  AOI21_X1 U1420 ( .B1(n274), .B2(n262), .A(n1474), .ZN(n261) );
  OAI21_X1 U1421 ( .B1(n281), .B2(n271), .A(n276), .ZN(n270) );
  NAND2_X1 U1422 ( .A1(n273), .A2(n262), .ZN(n260) );
  NAND2_X1 U1423 ( .A1(n214), .A2(n1400), .ZN(n201) );
  NAND2_X1 U1424 ( .A1(n186), .A2(n149), .ZN(n145) );
  INV_X1 U1425 ( .A(n1445), .ZN(n309) );
  INV_X1 U1426 ( .A(n273), .ZN(n271) );
  NAND2_X1 U1427 ( .A1(n1479), .A2(n1466), .ZN(n326) );
  INV_X1 U1428 ( .A(n119), .ZN(n117) );
  NOR2_X1 U1429 ( .A1(n1455), .A2(n225), .ZN(n223) );
  NOR2_X1 U1430 ( .A1(n1455), .A2(n160), .ZN(n158) );
  INV_X1 U1431 ( .A(n192), .ZN(n190) );
  INV_X1 U1432 ( .A(n1414), .ZN(n246) );
  INV_X1 U1433 ( .A(n1466), .ZN(n333) );
  INV_X1 U1434 ( .A(n263), .ZN(n262) );
  INV_X1 U1435 ( .A(n1480), .ZN(n263) );
  INV_X1 U1436 ( .A(n1469), .ZN(n334) );
  NAND2_X1 U1437 ( .A1(n287), .A2(n290), .ZN(n82) );
  AOI21_X1 U1438 ( .B1(n299), .B2(n319), .A(n300), .ZN(n298) );
  AOI21_X1 U1439 ( .B1(n1471), .B2(n1474), .A(n254), .ZN(n252) );
  XOR2_X1 U1440 ( .A(n347), .B(n90), .Z(product[15]) );
  NAND2_X1 U1441 ( .A1(n1457), .A2(n346), .ZN(n90) );
  XOR2_X1 U1442 ( .A(n339), .B(n89), .Z(product[16]) );
  NAND2_X1 U1443 ( .A1(n1466), .A2(n334), .ZN(n89) );
  XNOR2_X1 U1444 ( .A(n332), .B(n88), .ZN(product[17]) );
  NAND2_X1 U1445 ( .A1(n1479), .A2(n331), .ZN(n88) );
  OAI21_X1 U1446 ( .B1(n339), .B2(n333), .A(n334), .ZN(n332) );
  NOR2_X1 U1447 ( .A1(n323), .A2(n326), .ZN(n321) );
  INV_X1 U1448 ( .A(n1475), .ZN(n424) );
  AOI21_X1 U1449 ( .B1(n311), .B2(n294), .A(n295), .ZN(n293) );
  NAND2_X1 U1450 ( .A1(n315), .A2(n1472), .ZN(n86) );
  XOR2_X1 U1451 ( .A(n314), .B(n85), .Z(product[20]) );
  NAND2_X1 U1452 ( .A1(n428), .A2(n1467), .ZN(n85) );
  AOI21_X1 U1453 ( .B1(n319), .B2(n315), .A(n316), .ZN(n314) );
  INV_X1 U1454 ( .A(n312), .ZN(n428) );
  INV_X1 U1455 ( .A(n217), .ZN(n215) );
  NOR2_X1 U1456 ( .A1(n216), .A2(n121), .ZN(n119) );
  XOR2_X1 U1457 ( .A(n352), .B(n91), .Z(product[14]) );
  NAND2_X1 U1458 ( .A1(n434), .A2(n351), .ZN(n91) );
  AOI21_X1 U1459 ( .B1(n357), .B2(n435), .A(n354), .ZN(n352) );
  INV_X1 U1460 ( .A(n350), .ZN(n434) );
  AOI21_X1 U1461 ( .B1(n319), .B2(n306), .A(n1445), .ZN(n305) );
  AOI21_X1 U1462 ( .B1(n1469), .B2(n1479), .A(n1468), .ZN(n327) );
  OAI21_X1 U1463 ( .B1(n309), .B2(n301), .A(n304), .ZN(n300) );
  INV_X1 U1464 ( .A(n1389), .ZN(n357) );
  NOR2_X1 U1465 ( .A1(n312), .A2(n317), .ZN(n310) );
  INV_X1 U1466 ( .A(n367), .ZN(n366) );
  NOR2_X1 U1467 ( .A1(n192), .A2(n136), .ZN(n134) );
  OAI21_X1 U1468 ( .B1(n1414), .B2(n201), .A(n202), .ZN(n200) );
  AOI21_X1 U1469 ( .B1(n215), .B2(n1400), .A(n206), .ZN(n202) );
  OAI21_X1 U1470 ( .B1(n1414), .B2(n171), .A(n172), .ZN(n170) );
  INV_X1 U1471 ( .A(n174), .ZN(n172) );
  NAND2_X1 U1472 ( .A1(n240), .A2(n227), .ZN(n225) );
  NAND2_X1 U1473 ( .A1(n1400), .A2(n1402), .ZN(n192) );
  NAND2_X1 U1474 ( .A1(n173), .A2(n1407), .ZN(n160) );
  INV_X1 U1475 ( .A(n275), .ZN(n273) );
  NAND2_X1 U1476 ( .A1(n190), .A2(n177), .ZN(n175) );
  INV_X1 U1477 ( .A(n317), .ZN(n315) );
  INV_X1 U1478 ( .A(n302), .ZN(n301) );
  INV_X1 U1479 ( .A(n276), .ZN(n274) );
  INV_X1 U1480 ( .A(n193), .ZN(n191) );
  XNOR2_X1 U1481 ( .A(n325), .B(n87), .ZN(product[18]) );
  NAND2_X1 U1482 ( .A1(n430), .A2(n324), .ZN(n87) );
  INV_X1 U1483 ( .A(n323), .ZN(n430) );
  INV_X1 U1484 ( .A(n256), .ZN(n254) );
  INV_X1 U1485 ( .A(n318), .ZN(n316) );
  INV_X1 U1486 ( .A(n290), .ZN(n288) );
  INV_X1 U1487 ( .A(n346), .ZN(n344) );
  XOR2_X1 U1488 ( .A(n374), .B(n95), .Z(product[10]) );
  NAND2_X1 U1489 ( .A1(n1388), .A2(n373), .ZN(n95) );
  AOI21_X1 U1490 ( .B1(n379), .B2(n1405), .A(n376), .ZN(n374) );
  XNOR2_X1 U1491 ( .A(n363), .B(n93), .ZN(product[12]) );
  NAND2_X1 U1492 ( .A1(n436), .A2(n362), .ZN(n93) );
  OAI21_X1 U1493 ( .B1(n366), .B2(n364), .A(n365), .ZN(n363) );
  XNOR2_X1 U1494 ( .A(n357), .B(n92), .ZN(product[13]) );
  NAND2_X1 U1495 ( .A1(n435), .A2(n356), .ZN(n92) );
  INV_X1 U1496 ( .A(n355), .ZN(n435) );
  XNOR2_X1 U1497 ( .A(n379), .B(n96), .ZN(product[9]) );
  NAND2_X1 U1498 ( .A1(n1405), .A2(n378), .ZN(n96) );
  OAI21_X1 U1499 ( .B1(n217), .B2(n175), .A(n176), .ZN(n174) );
  AOI21_X1 U1500 ( .B1(n191), .B2(n177), .A(n178), .ZN(n176) );
  INV_X1 U1501 ( .A(n180), .ZN(n178) );
  XOR2_X1 U1502 ( .A(n198), .B(n73), .Z(product[32]) );
  NAND2_X1 U1503 ( .A1(n1402), .A2(n197), .ZN(n73) );
  XOR2_X1 U1504 ( .A(n181), .B(n72), .Z(product[33]) );
  NAND2_X1 U1505 ( .A1(n177), .A2(n180), .ZN(n72) );
  AOI21_X1 U1506 ( .B1(n1402), .B2(n206), .A(n195), .ZN(n193) );
  INV_X1 U1507 ( .A(n197), .ZN(n195) );
  INV_X1 U1508 ( .A(n220), .ZN(n418) );
  AOI21_X1 U1509 ( .B1(n218), .B2(n241), .A(n219), .ZN(n217) );
  OAI21_X1 U1510 ( .B1(n230), .B2(n220), .A(n221), .ZN(n219) );
  OAI21_X1 U1511 ( .B1(n368), .B2(n380), .A(n369), .ZN(n367) );
  NAND2_X1 U1512 ( .A1(n1388), .A2(n1405), .ZN(n368) );
  AOI21_X1 U1513 ( .B1(n1388), .B2(n376), .A(n371), .ZN(n369) );
  AOI21_X1 U1514 ( .B1(n367), .B2(n359), .A(n360), .ZN(n358) );
  NOR2_X1 U1515 ( .A1(n179), .A2(n151), .ZN(n149) );
  OAI21_X1 U1516 ( .B1(n1414), .B2(n130), .A(n131), .ZN(n129) );
  AOI21_X1 U1517 ( .B1(n215), .B2(n134), .A(n135), .ZN(n131) );
  OAI21_X1 U1518 ( .B1(n1414), .B2(n160), .A(n161), .ZN(n159) );
  AOI21_X1 U1519 ( .B1(n174), .B2(n1407), .A(n165), .ZN(n161) );
  INV_X1 U1520 ( .A(n229), .ZN(n227) );
  NAND2_X1 U1521 ( .A1(n134), .A2(n1406), .ZN(n121) );
  INV_X1 U1522 ( .A(n380), .ZN(n379) );
  NAND2_X1 U1523 ( .A1(n611), .A2(n628), .ZN(n313) );
  NAND2_X1 U1524 ( .A1(n561), .A2(n576), .ZN(n290) );
  NAND2_X1 U1525 ( .A1(n593), .A2(n610), .ZN(n304) );
  OAI21_X1 U1526 ( .B1(n1458), .B2(n117), .A(n118), .ZN(n116) );
  INV_X1 U1527 ( .A(n120), .ZN(n118) );
  OAI21_X1 U1528 ( .B1(n65), .B2(n225), .A(n226), .ZN(n224) );
  AOI21_X1 U1529 ( .B1(n241), .B2(n227), .A(n228), .ZN(n226) );
  INV_X1 U1530 ( .A(n230), .ZN(n228) );
  OAI21_X1 U1531 ( .B1(n1414), .B2(n145), .A(n146), .ZN(n144) );
  AOI21_X1 U1532 ( .B1(n187), .B2(n149), .A(n150), .ZN(n146) );
  NAND2_X1 U1533 ( .A1(n693), .A2(n706), .ZN(n346) );
  INV_X1 U1534 ( .A(n179), .ZN(n177) );
  NAND2_X1 U1535 ( .A1(n119), .A2(n1403), .ZN(n108) );
  NAND2_X1 U1536 ( .A1(n149), .A2(n1404), .ZN(n136) );
  NAND2_X1 U1537 ( .A1(n547), .A2(n560), .ZN(n285) );
  NAND2_X1 U1538 ( .A1(n647), .A2(n662), .ZN(n324) );
  NAND2_X1 U1539 ( .A1(n707), .A2(n718), .ZN(n351) );
  NAND2_X1 U1540 ( .A1(n1407), .A2(n1401), .ZN(n151) );
  INV_X1 U1541 ( .A(n242), .ZN(n240) );
  NAND2_X1 U1542 ( .A1(n577), .A2(n592), .ZN(n297) );
  INV_X1 U1543 ( .A(n243), .ZN(n241) );
  INV_X1 U1544 ( .A(n208), .ZN(n206) );
  NOR2_X1 U1545 ( .A1(n1455), .A2(n108), .ZN(n106) );
  OAI21_X1 U1546 ( .B1(n1458), .B2(n108), .A(n109), .ZN(n107) );
  INV_X1 U1547 ( .A(n378), .ZN(n376) );
  XOR2_X1 U1548 ( .A(n366), .B(n94), .Z(product[11]) );
  NAND2_X1 U1549 ( .A1(n437), .A2(n365), .ZN(n94) );
  INV_X1 U1550 ( .A(n364), .ZN(n437) );
  INV_X1 U1551 ( .A(n356), .ZN(n354) );
  INV_X1 U1552 ( .A(n373), .ZN(n371) );
  NAND2_X1 U1553 ( .A1(n1408), .A2(n384), .ZN(n97) );
  AOI21_X1 U1554 ( .B1(n135), .B2(n1406), .A(n124), .ZN(n122) );
  INV_X1 U1555 ( .A(n126), .ZN(n124) );
  NAND2_X1 U1556 ( .A1(n1401), .A2(n156), .ZN(n70) );
  XOR2_X1 U1557 ( .A(n142), .B(n69), .Z(product[36]) );
  NAND2_X1 U1558 ( .A1(n1404), .A2(n141), .ZN(n69) );
  XOR2_X1 U1559 ( .A(n114), .B(n67), .Z(product[38]) );
  NAND2_X1 U1560 ( .A1(n1403), .A2(n113), .ZN(n67) );
  XOR2_X1 U1561 ( .A(n168), .B(n71), .Z(product[34]) );
  NAND2_X1 U1562 ( .A1(n1407), .A2(n167), .ZN(n71) );
  XOR2_X1 U1563 ( .A(n127), .B(n68), .Z(product[37]) );
  NAND2_X1 U1564 ( .A1(n1406), .A2(n126), .ZN(n68) );
  AOI21_X1 U1565 ( .B1(n385), .B2(n1408), .A(n382), .ZN(n380) );
  INV_X1 U1566 ( .A(n384), .ZN(n382) );
  AOI21_X1 U1567 ( .B1(n1409), .B2(n393), .A(n390), .ZN(n388) );
  INV_X1 U1568 ( .A(n392), .ZN(n390) );
  OAI21_X1 U1569 ( .B1(n394), .B2(n396), .A(n395), .ZN(n393) );
  OAI21_X1 U1570 ( .B1(n388), .B2(n386), .A(n387), .ZN(n385) );
  NOR2_X1 U1571 ( .A1(n489), .A2(n498), .ZN(n229) );
  OAI21_X1 U1572 ( .B1(n151), .B2(n180), .A(n152), .ZN(n150) );
  AOI21_X1 U1573 ( .B1(n165), .B2(n1401), .A(n154), .ZN(n152) );
  INV_X1 U1574 ( .A(n156), .ZN(n154) );
  OAI21_X1 U1575 ( .B1(n193), .B2(n136), .A(n137), .ZN(n135) );
  AOI21_X1 U1576 ( .B1(n150), .B2(n1404), .A(n139), .ZN(n137) );
  INV_X1 U1577 ( .A(n141), .ZN(n139) );
  AOI21_X1 U1578 ( .B1(n120), .B2(n1403), .A(n111), .ZN(n109) );
  INV_X1 U1579 ( .A(n113), .ZN(n111) );
  NAND2_X1 U1580 ( .A1(n461), .A2(n466), .ZN(n180) );
  NAND2_X1 U1581 ( .A1(n489), .A2(n498), .ZN(n230) );
  NAND2_X1 U1582 ( .A1(n719), .A2(n730), .ZN(n356) );
  NAND2_X1 U1583 ( .A1(n741), .A2(n750), .ZN(n365) );
  NAND2_X1 U1584 ( .A1(n751), .A2(n758), .ZN(n373) );
  NAND2_X1 U1585 ( .A1(n499), .A2(n508), .ZN(n243) );
  NAND2_X1 U1586 ( .A1(n467), .A2(n472), .ZN(n197) );
  NAND2_X1 U1587 ( .A1(n481), .A2(n488), .ZN(n221) );
  NAND2_X1 U1588 ( .A1(n759), .A2(n766), .ZN(n378) );
  NAND2_X1 U1589 ( .A1(n731), .A2(n740), .ZN(n362) );
  INV_X1 U1590 ( .A(n167), .ZN(n165) );
  NAND2_X1 U1591 ( .A1(n441), .A2(n387), .ZN(n98) );
  INV_X1 U1592 ( .A(n386), .ZN(n441) );
  NAND2_X1 U1593 ( .A1(n1409), .A2(n392), .ZN(n99) );
  XOR2_X1 U1594 ( .A(n100), .B(n396), .Z(product[5]) );
  NAND2_X1 U1595 ( .A1(n443), .A2(n395), .ZN(n100) );
  INV_X1 U1596 ( .A(n394), .ZN(n443) );
  XOR2_X1 U1597 ( .A(n102), .B(n404), .Z(product[3]) );
  NAND2_X1 U1598 ( .A1(n445), .A2(n403), .ZN(n102) );
  INV_X1 U1599 ( .A(n402), .ZN(n445) );
  XOR2_X1 U1600 ( .A(n103), .B(n409), .Z(product[2]) );
  NAND2_X1 U1601 ( .A1(n446), .A2(n407), .ZN(n103) );
  INV_X1 U1602 ( .A(n406), .ZN(n446) );
  XNOR2_X1 U1603 ( .A(n101), .B(n401), .ZN(product[4]) );
  NAND2_X1 U1604 ( .A1(n1410), .A2(n400), .ZN(n101) );
  OAI21_X1 U1605 ( .B1(n402), .B2(n404), .A(n403), .ZN(n401) );
  AOI21_X1 U1606 ( .B1(n1410), .B2(n401), .A(n398), .ZN(n396) );
  INV_X1 U1607 ( .A(n400), .ZN(n398) );
  NAND2_X1 U1608 ( .A1(n1028), .A2(n1009), .ZN(n407) );
  NAND2_X1 U1609 ( .A1(n830), .A2(n448), .ZN(n113) );
  NOR2_X1 U1610 ( .A1(n783), .A2(n786), .ZN(n394) );
  INV_X1 U1611 ( .A(n448), .ZN(n449) );
  INV_X1 U1612 ( .A(n1436), .ZN(n545) );
  INV_X1 U1613 ( .A(n478), .ZN(n479) );
  OR2_X1 U1614 ( .A1(n937), .A2(n865), .ZN(n626) );
  XNOR2_X1 U1615 ( .A(n937), .B(n865), .ZN(n627) );
  NAND2_X1 U1616 ( .A1(n779), .A2(n782), .ZN(n392) );
  NAND2_X1 U1617 ( .A1(n457), .A2(n460), .ZN(n167) );
  NAND2_X1 U1618 ( .A1(n453), .A2(n456), .ZN(n156) );
  NAND2_X1 U1619 ( .A1(n452), .A2(n451), .ZN(n141) );
  NAND2_X1 U1620 ( .A1(n450), .A2(n449), .ZN(n126) );
  NAND2_X1 U1621 ( .A1(n773), .A2(n778), .ZN(n387) );
  NAND2_X1 U1622 ( .A1(n783), .A2(n786), .ZN(n395) );
  INV_X1 U1623 ( .A(n405), .ZN(n404) );
  OAI21_X1 U1624 ( .B1(n406), .B2(n409), .A(n407), .ZN(n405) );
  OAI22_X1 U1625 ( .A1(n42), .A2(n1094), .B1(n40), .B2(n1093), .ZN(n478) );
  OAI22_X1 U1626 ( .A1(n30), .A2(n1136), .B1(n28), .B2(n1135), .ZN(n518) );
  OAI22_X1 U1627 ( .A1(n24), .A2(n1157), .B1(n1156), .B2(n22), .ZN(n544) );
  OAI22_X1 U1628 ( .A1(n18), .A2(n1178), .B1(n16), .B2(n1177), .ZN(n574) );
  OAI22_X1 U1629 ( .A1(n1387), .A2(n1199), .B1(n1198), .B2(n10), .ZN(n608) );
  OAI22_X1 U1630 ( .A1(n48), .A2(n1073), .B1(n46), .B2(n1072), .ZN(n464) );
  OAI22_X1 U1631 ( .A1(n36), .A2(n1115), .B1(n34), .B2(n1114), .ZN(n496) );
  OAI22_X1 U1632 ( .A1(n53), .A2(n1067), .B1(n51), .B2(n1066), .ZN(n865) );
  OAI22_X1 U1633 ( .A1(n30), .A2(n1143), .B1(n28), .B2(n1142), .ZN(n937) );
  INV_X1 U1634 ( .A(n793), .ZN(n850) );
  OAI22_X1 U1635 ( .A1(n60), .A2(n1032), .B1(n58), .B2(n1031), .ZN(n831) );
  AOI21_X1 U1636 ( .B1(n54), .B2(n52), .A(n1051), .ZN(n793) );
  OAI22_X1 U1637 ( .A1(n60), .A2(n1034), .B1(n58), .B2(n1033), .ZN(n833) );
  OAI22_X1 U1638 ( .A1(n60), .A2(n1033), .B1(n58), .B2(n1032), .ZN(n832) );
  INV_X1 U1639 ( .A(n454), .ZN(n455) );
  OAI22_X1 U1640 ( .A1(n1390), .A2(n1234), .B1(n1233), .B2(n4), .ZN(n1025) );
  OAI22_X1 U1641 ( .A1(n1387), .A2(n1215), .B1(n9), .B2(n1214), .ZN(n1006) );
  OAI22_X1 U1642 ( .A1(n17), .A2(n1195), .B1(n15), .B2(n1194), .ZN(n987) );
  AND2_X1 U1643 ( .A1(n1492), .A2(n812), .ZN(n989) );
  OAI22_X1 U1644 ( .A1(n11), .A2(n1216), .B1(n9), .B2(n1215), .ZN(n1007) );
  OAI22_X1 U1645 ( .A1(n1391), .A2(n1235), .B1(n1234), .B2(n4), .ZN(n1026) );
  OAI22_X1 U1646 ( .A1(n30), .A2(n1295), .B1(n1155), .B2(n28), .ZN(n825) );
  OAI22_X1 U1647 ( .A1(n29), .A2(n1154), .B1(n27), .B2(n1153), .ZN(n948) );
  OR2_X1 U1648 ( .A1(n1492), .A2(n1295), .ZN(n1155) );
  OAI22_X1 U1649 ( .A1(n1387), .A2(n1207), .B1(n10), .B2(n1206), .ZN(n998) );
  OAI22_X1 U1650 ( .A1(n5), .A2(n1226), .B1(n1225), .B2(n4), .ZN(n1017) );
  OAI22_X1 U1651 ( .A1(n23), .A2(n1169), .B1(n1443), .B2(n1168), .ZN(n962) );
  OAI22_X1 U1652 ( .A1(n1391), .A2(n1232), .B1(n1231), .B2(n4), .ZN(n1023) );
  OAI22_X1 U1653 ( .A1(n1387), .A2(n1213), .B1(n9), .B2(n1212), .ZN(n1004) );
  OAI22_X1 U1654 ( .A1(n17), .A2(n1194), .B1(n15), .B2(n1193), .ZN(n986) );
  OAI22_X1 U1655 ( .A1(n30), .A2(n1140), .B1(n28), .B2(n1139), .ZN(n934) );
  OAI22_X1 U1656 ( .A1(n24), .A2(n1159), .B1(n22), .B2(n1158), .ZN(n952) );
  OAI22_X1 U1657 ( .A1(n48), .A2(n1083), .B1(n45), .B2(n1082), .ZN(n880) );
  OAI22_X1 U1658 ( .A1(n53), .A2(n1062), .B1(n51), .B2(n1061), .ZN(n860) );
  OAI22_X1 U1659 ( .A1(n59), .A2(n1043), .B1(n1481), .B2(n1042), .ZN(n842) );
  OAI22_X1 U1660 ( .A1(n1477), .A2(n1081), .B1(n46), .B2(n1080), .ZN(n878) );
  OAI22_X1 U1661 ( .A1(n41), .A2(n1106), .B1(n39), .B2(n1105), .ZN(n902) );
  OAI22_X1 U1662 ( .A1(n5), .A2(n1220), .B1(n1424), .B2(n4), .ZN(n1011) );
  OAI22_X1 U1663 ( .A1(n24), .A2(n1163), .B1(n1443), .B2(n1162), .ZN(n956) );
  OAI22_X1 U1664 ( .A1(n24), .A2(n1160), .B1(n22), .B2(n1159), .ZN(n953) );
  OAI22_X1 U1665 ( .A1(n53), .A2(n1065), .B1(n51), .B2(n1064), .ZN(n863) );
  OAI22_X1 U1666 ( .A1(n41), .A2(n1105), .B1(n39), .B2(n1104), .ZN(n901) );
  OAI22_X1 U1667 ( .A1(n12), .A2(n1200), .B1(n10), .B2(n1199), .ZN(n991) );
  OAI22_X1 U1668 ( .A1(n48), .A2(n1086), .B1(n45), .B2(n1085), .ZN(n883) );
  OAI22_X1 U1669 ( .A1(n29), .A2(n1144), .B1(n28), .B2(n1143), .ZN(n938) );
  OAI22_X1 U1670 ( .A1(n53), .A2(n1068), .B1(n1067), .B2(n51), .ZN(n866) );
  OAI22_X1 U1671 ( .A1(n1477), .A2(n1437), .B1(n45), .B2(n1086), .ZN(n884) );
  AOI21_X1 U1672 ( .B1(n42), .B2(n40), .A(n1093), .ZN(n799) );
  AOI21_X1 U1673 ( .B1(n36), .B2(n34), .A(n1114), .ZN(n802) );
  AOI21_X1 U1674 ( .B1(n12), .B2(n10), .A(n1198), .ZN(n814) );
  OAI22_X1 U1675 ( .A1(n54), .A2(n1291), .B1(n1071), .B2(n52), .ZN(n821) );
  OAI22_X1 U1676 ( .A1(n53), .A2(n1070), .B1(n51), .B2(n1069), .ZN(n868) );
  OR2_X1 U1677 ( .A1(n1491), .A2(n1291), .ZN(n1071) );
  NAND2_X1 U1678 ( .A1(n1029), .A2(n829), .ZN(n409) );
  NAND2_X1 U1679 ( .A1(n789), .A2(n828), .ZN(n403) );
  XNOR2_X1 U1680 ( .A(n1483), .B(n1420), .ZN(n1091) );
  AND2_X1 U1681 ( .A1(n1492), .A2(n815), .ZN(n1009) );
  INV_X1 U1682 ( .A(n9), .ZN(n815) );
  AND2_X1 U1683 ( .A1(n1492), .A2(n818), .ZN(product[0]) );
  INV_X1 U1684 ( .A(n1289), .ZN(n818) );
  INV_X1 U1685 ( .A(n805), .ZN(n930) );
  OAI22_X1 U1686 ( .A1(n59), .A2(n1040), .B1(n1481), .B2(n1039), .ZN(n839) );
  AOI21_X1 U1687 ( .B1(n30), .B2(n28), .A(n1135), .ZN(n805) );
  OAI22_X1 U1688 ( .A1(n54), .A2(n1054), .B1(n52), .B2(n1053), .ZN(n852) );
  OAI22_X1 U1689 ( .A1(n60), .A2(n1035), .B1(n58), .B2(n1034), .ZN(n834) );
  INV_X1 U1690 ( .A(n464), .ZN(n465) );
  OAI22_X1 U1691 ( .A1(n30), .A2(n1138), .B1(n28), .B2(n1137), .ZN(n932) );
  OAI22_X1 U1692 ( .A1(n42), .A2(n1100), .B1(n40), .B2(n1099), .ZN(n896) );
  OAI22_X1 U1693 ( .A1(n35), .A2(n1119), .B1(n34), .B2(n1118), .ZN(n914) );
  OAI22_X1 U1694 ( .A1(n30), .A2(n1137), .B1(n28), .B2(n1136), .ZN(n931) );
  OAI22_X1 U1695 ( .A1(n53), .A2(n1061), .B1(n51), .B2(n1060), .ZN(n859) );
  OAI22_X1 U1696 ( .A1(n36), .A2(n1118), .B1(n34), .B2(n1117), .ZN(n913) );
  OAI22_X1 U1697 ( .A1(n54), .A2(n1057), .B1(n52), .B2(n1056), .ZN(n855) );
  OAI22_X1 U1698 ( .A1(n1477), .A2(n1076), .B1(n46), .B2(n1075), .ZN(n873) );
  OAI22_X1 U1699 ( .A1(n12), .A2(n1204), .B1(n10), .B2(n1203), .ZN(n995) );
  OAI22_X1 U1700 ( .A1(n35), .A2(n1128), .B1(n33), .B2(n1127), .ZN(n923) );
  OAI22_X1 U1701 ( .A1(n47), .A2(n1090), .B1(n1089), .B2(n45), .ZN(n887) );
  OAI22_X1 U1702 ( .A1(n42), .A2(n1099), .B1(n40), .B2(n1098), .ZN(n895) );
  OAI22_X1 U1703 ( .A1(n48), .A2(n1080), .B1(n46), .B2(n1079), .ZN(n877) );
  OAI22_X1 U1704 ( .A1(n18), .A2(n1182), .B1(n16), .B2(n1181), .ZN(n974) );
  OAI22_X1 U1705 ( .A1(n11), .A2(n1201), .B1(n10), .B2(n1200), .ZN(n992) );
  OAI22_X1 U1706 ( .A1(n36), .A2(n1125), .B1(n33), .B2(n1439), .ZN(n920) );
  OAI22_X1 U1707 ( .A1(n6), .A2(n1221), .B1(n1220), .B2(n4), .ZN(n1012) );
  AND2_X1 U1708 ( .A1(n1420), .A2(n791), .ZN(n849) );
  OAI22_X1 U1709 ( .A1(n47), .A2(n1459), .B1(n45), .B2(n1087), .ZN(n885) );
  OAI22_X1 U1710 ( .A1(n42), .A2(n1096), .B1(n40), .B2(n1095), .ZN(n892) );
  OAI22_X1 U1711 ( .A1(n54), .A2(n1058), .B1(n52), .B2(n1057), .ZN(n856) );
  OAI22_X1 U1712 ( .A1(n60), .A2(n1039), .B1(n58), .B2(n1038), .ZN(n838) );
  OAI22_X1 U1713 ( .A1(n24), .A2(n1162), .B1(n1443), .B2(n1161), .ZN(n955) );
  OAI22_X1 U1714 ( .A1(n18), .A2(n1181), .B1(n16), .B2(n1180), .ZN(n973) );
  OAI22_X1 U1715 ( .A1(n54), .A2(n1059), .B1(n52), .B2(n1058), .ZN(n857) );
  OAI22_X1 U1716 ( .A1(n48), .A2(n1078), .B1(n46), .B2(n1077), .ZN(n875) );
  OAI22_X1 U1717 ( .A1(n36), .A2(n1116), .B1(n34), .B2(n1115), .ZN(n911) );
  OAI22_X1 U1718 ( .A1(n1477), .A2(n1077), .B1(n46), .B2(n1076), .ZN(n874) );
  INV_X1 U1719 ( .A(n496), .ZN(n497) );
  OAI22_X1 U1720 ( .A1(n30), .A2(n1139), .B1(n28), .B2(n1138), .ZN(n933) );
  OAI22_X1 U1721 ( .A1(n24), .A2(n1158), .B1(n1443), .B2(n1157), .ZN(n951) );
  OAI22_X1 U1722 ( .A1(n53), .A2(n1063), .B1(n51), .B2(n1062), .ZN(n861) );
  OAI22_X1 U1723 ( .A1(n41), .A2(n1107), .B1(n39), .B2(n1106), .ZN(n903) );
  OAI22_X1 U1724 ( .A1(n11), .A2(n1202), .B1(n10), .B2(n1201), .ZN(n993) );
  OAI22_X1 U1725 ( .A1(n53), .A2(n1069), .B1(n51), .B2(n1068), .ZN(n867) );
  INV_X1 U1726 ( .A(n1481), .ZN(n791) );
  OAI22_X1 U1727 ( .A1(n18), .A2(n1180), .B1(n16), .B2(n1418), .ZN(n972) );
  OAI22_X1 U1728 ( .A1(n59), .A2(n1441), .B1(n1481), .B2(n1046), .ZN(n846) );
  OAI22_X1 U1729 ( .A1(n53), .A2(n1064), .B1(n51), .B2(n1063), .ZN(n862) );
  OAI22_X1 U1730 ( .A1(n59), .A2(n1045), .B1(n1481), .B2(n1044), .ZN(n844) );
  OAI22_X1 U1731 ( .A1(n36), .A2(n1121), .B1(n34), .B2(n1120), .ZN(n916) );
  OAI22_X1 U1732 ( .A1(n36), .A2(n1122), .B1(n34), .B2(n1121), .ZN(n917) );
  OAI22_X1 U1733 ( .A1(n41), .A2(n1103), .B1(n39), .B2(n1102), .ZN(n899) );
  OAI22_X1 U1734 ( .A1(n30), .A2(n1141), .B1(n28), .B2(n1140), .ZN(n935) );
  OAI22_X1 U1735 ( .A1(n1477), .A2(n1084), .B1(n45), .B2(n1083), .ZN(n881) );
  OAI22_X1 U1736 ( .A1(n24), .A2(n1164), .B1(n22), .B2(n1163), .ZN(n957) );
  OAI22_X1 U1737 ( .A1(n24), .A2(n1165), .B1(n22), .B2(n1164), .ZN(n958) );
  OAI22_X1 U1738 ( .A1(n18), .A2(n1184), .B1(n16), .B2(n1183), .ZN(n976) );
  OAI22_X1 U1739 ( .A1(n41), .A2(n1110), .B1(n39), .B2(n1109), .ZN(n906) );
  OAI22_X1 U1740 ( .A1(n1167), .A2(n23), .B1(n1166), .B2(n22), .ZN(n960) );
  OAI22_X1 U1741 ( .A1(n35), .A2(n1129), .B1(n33), .B2(n1128), .ZN(n924) );
  OAI22_X1 U1742 ( .A1(n29), .A2(n1150), .B1(n27), .B2(n1149), .ZN(n944) );
  OAI22_X1 U1743 ( .A1(n17), .A2(n1188), .B1(n15), .B2(n1187), .ZN(n980) );
  OAI22_X1 U1744 ( .A1(n36), .A2(n1131), .B1(n33), .B2(n1130), .ZN(n926) );
  OAI22_X1 U1745 ( .A1(n23), .A2(n1413), .B1(n22), .B2(n1165), .ZN(n959) );
  OAI22_X1 U1746 ( .A1(n29), .A2(n1147), .B1(n27), .B2(n1146), .ZN(n941) );
  OAI22_X1 U1747 ( .A1(n18), .A2(n1185), .B1(n1184), .B2(n16), .ZN(n977) );
  OAI22_X1 U1748 ( .A1(n1391), .A2(n1227), .B1(n1226), .B2(n4), .ZN(n1018) );
  AND2_X1 U1749 ( .A1(n1420), .A2(n800), .ZN(n909) );
  OAI22_X1 U1750 ( .A1(n1151), .A2(n29), .B1(n27), .B2(n1150), .ZN(n945) );
  OAI22_X1 U1751 ( .A1(n17), .A2(n1191), .B1(n15), .B2(n1190), .ZN(n983) );
  OAI22_X1 U1752 ( .A1(n29), .A2(n1153), .B1(n27), .B2(n1152), .ZN(n947) );
  OAI22_X1 U1753 ( .A1(n11), .A2(n1210), .B1(n9), .B2(n1209), .ZN(n1001) );
  OAI22_X1 U1754 ( .A1(n1387), .A2(n1211), .B1(n9), .B2(n1210), .ZN(n1002) );
  OAI22_X1 U1755 ( .A1(n23), .A2(n1173), .B1(n22), .B2(n1172), .ZN(n966) );
  OAI22_X1 U1756 ( .A1(n17), .A2(n1192), .B1(n15), .B2(n1191), .ZN(n984) );
  INV_X1 U1757 ( .A(n811), .ZN(n970) );
  OAI22_X1 U1758 ( .A1(n59), .A2(n1044), .B1(n1481), .B2(n1043), .ZN(n843) );
  AOI21_X1 U1759 ( .B1(n18), .B2(n16), .A(n1177), .ZN(n811) );
  OAI22_X1 U1760 ( .A1(n59), .A2(n1048), .B1(n1047), .B2(n1481), .ZN(n847) );
  OAI22_X1 U1761 ( .A1(n1124), .A2(n35), .B1(n1123), .B2(n33), .ZN(n919) );
  OAI22_X1 U1762 ( .A1(n23), .A2(n1168), .B1(n22), .B2(n1167), .ZN(n961) );
  OAI22_X1 U1763 ( .A1(n17), .A2(n1187), .B1(n15), .B2(n1186), .ZN(n979) );
  INV_X1 U1764 ( .A(n808), .ZN(n950) );
  OAI22_X1 U1765 ( .A1(n59), .A2(n1042), .B1(n1481), .B2(n1041), .ZN(n841) );
  AOI21_X1 U1766 ( .B1(n24), .B2(n1443), .A(n1156), .ZN(n808) );
  OAI22_X1 U1767 ( .A1(n23), .A2(n1174), .B1(n1443), .B2(n1173), .ZN(n967) );
  OAI22_X1 U1768 ( .A1(n1387), .A2(n1212), .B1(n9), .B2(n1211), .ZN(n1003) );
  AND2_X1 U1769 ( .A1(n1420), .A2(n809), .ZN(n969) );
  OAI22_X1 U1770 ( .A1(n1391), .A2(n1233), .B1(n1232), .B2(n4), .ZN(n1024) );
  OAI22_X1 U1771 ( .A1(n1387), .A2(n1214), .B1(n9), .B2(n1213), .ZN(n1005) );
  OAI22_X1 U1772 ( .A1(n42), .A2(n1102), .B1(n40), .B2(n1101), .ZN(n898) );
  INV_X1 U1773 ( .A(n574), .ZN(n575) );
  OAI22_X1 U1774 ( .A1(n5), .A2(n1230), .B1(n1229), .B2(n4), .ZN(n1021) );
  OAI22_X1 U1775 ( .A1(n42), .A2(n1101), .B1(n40), .B2(n1100), .ZN(n897) );
  OAI22_X1 U1776 ( .A1(n1477), .A2(n1082), .B1(n45), .B2(n1081), .ZN(n879) );
  OAI22_X1 U1777 ( .A1(n36), .A2(n1120), .B1(n34), .B2(n1119), .ZN(n915) );
  OAI22_X1 U1778 ( .A1(n42), .A2(n1098), .B1(n40), .B2(n1097), .ZN(n894) );
  OAI22_X1 U1779 ( .A1(n1477), .A2(n1079), .B1(n46), .B2(n1078), .ZN(n876) );
  OAI22_X1 U1780 ( .A1(n36), .A2(n1117), .B1(n34), .B2(n1116), .ZN(n912) );
  OAI22_X1 U1781 ( .A1(n29), .A2(n1145), .B1(n27), .B2(n1144), .ZN(n939) );
  OAI22_X1 U1782 ( .A1(n18), .A2(n1183), .B1(n16), .B2(n1182), .ZN(n975) );
  OAI22_X1 U1783 ( .A1(n35), .A2(n1126), .B1(n33), .B2(n1125), .ZN(n921) );
  OAI22_X1 U1784 ( .A1(n1390), .A2(n1225), .B1(n1224), .B2(n4), .ZN(n1016) );
  AND2_X1 U1785 ( .A1(n1420), .A2(n797), .ZN(n889) );
  OAI22_X1 U1786 ( .A1(n35), .A2(n1130), .B1(n33), .B2(n1129), .ZN(n925) );
  OAI22_X1 U1787 ( .A1(n1391), .A2(n1229), .B1(n1228), .B2(n4), .ZN(n1020) );
  OAI22_X1 U1788 ( .A1(n23), .A2(n1172), .B1(n1443), .B2(n1171), .ZN(n965) );
  AND2_X1 U1789 ( .A1(n1420), .A2(n803), .ZN(n929) );
  OAI22_X1 U1790 ( .A1(n41), .A2(n1108), .B1(n39), .B2(n1107), .ZN(n904) );
  OAI22_X1 U1791 ( .A1(n48), .A2(n1089), .B1(n45), .B2(n1459), .ZN(n886) );
  OAI22_X1 U1792 ( .A1(n36), .A2(n1127), .B1(n33), .B2(n1126), .ZN(n922) );
  OAI22_X1 U1793 ( .A1(n11), .A2(n1205), .B1(n10), .B2(n1204), .ZN(n996) );
  OAI22_X1 U1794 ( .A1(n6), .A2(n1223), .B1(n1222), .B2(n4), .ZN(n1014) );
  AND2_X1 U1795 ( .A1(n1492), .A2(n794), .ZN(n869) );
  OAI22_X1 U1796 ( .A1(n41), .A2(n1109), .B1(n39), .B2(n1108), .ZN(n905) );
  OAI22_X1 U1797 ( .A1(n29), .A2(n1149), .B1(n27), .B2(n1148), .ZN(n943) );
  OAI22_X1 U1798 ( .A1(n41), .A2(n1111), .B1(n39), .B2(n1110), .ZN(n907) );
  OAI22_X1 U1799 ( .A1(n1387), .A2(n1206), .B1(n10), .B2(n1205), .ZN(n997) );
  OAI22_X1 U1800 ( .A1(n30), .A2(n1142), .B1(n28), .B2(n1141), .ZN(n936) );
  INV_X1 U1801 ( .A(n608), .ZN(n609) );
  OAI22_X1 U1802 ( .A1(n36), .A2(n1434), .B1(n34), .B2(n1122), .ZN(n918) );
  OAI22_X1 U1803 ( .A1(n54), .A2(n1055), .B1(n52), .B2(n1054), .ZN(n853) );
  INV_X1 U1804 ( .A(n799), .ZN(n890) );
  OAI22_X1 U1805 ( .A1(n60), .A2(n1036), .B1(n58), .B2(n1035), .ZN(n835) );
  OAI22_X1 U1806 ( .A1(n18), .A2(n1179), .B1(n1178), .B2(n16), .ZN(n971) );
  INV_X1 U1807 ( .A(n814), .ZN(n990) );
  OAI22_X1 U1808 ( .A1(n1046), .A2(n59), .B1(n1481), .B2(n1045), .ZN(n845) );
  OAI22_X1 U1809 ( .A1(n54), .A2(n1060), .B1(n52), .B2(n1059), .ZN(n858) );
  INV_X1 U1810 ( .A(n518), .ZN(n519) );
  OAI22_X1 U1811 ( .A1(n59), .A2(n1041), .B1(n1481), .B2(n1040), .ZN(n840) );
  OAI22_X1 U1812 ( .A1(n54), .A2(n1056), .B1(n52), .B2(n1055), .ZN(n854) );
  OAI22_X1 U1813 ( .A1(n1477), .A2(n1075), .B1(n46), .B2(n1074), .ZN(n872) );
  OAI22_X1 U1814 ( .A1(n60), .A2(n1037), .B1(n58), .B2(n1036), .ZN(n836) );
  OAI22_X1 U1815 ( .A1(n23), .A2(n1171), .B1(n22), .B2(n1170), .ZN(n964) );
  OAI22_X1 U1816 ( .A1(n11), .A2(n1209), .B1(n9), .B2(n1208), .ZN(n1000) );
  OAI22_X1 U1817 ( .A1(n42), .A2(n1097), .B1(n40), .B2(n1096), .ZN(n893) );
  OAI22_X1 U1818 ( .A1(n17), .A2(n1189), .B1(n15), .B2(n1188), .ZN(n981) );
  OAI22_X1 U1819 ( .A1(n23), .A2(n1170), .B1(n1443), .B2(n1169), .ZN(n963) );
  OAI22_X1 U1820 ( .A1(n12), .A2(n1208), .B1(n9), .B2(n1207), .ZN(n999) );
  OAI22_X1 U1821 ( .A1(n36), .A2(n1132), .B1(n33), .B2(n1131), .ZN(n927) );
  OAI22_X1 U1822 ( .A1(n1387), .A2(n1422), .B1(n10), .B2(n1202), .ZN(n994) );
  OAI22_X1 U1823 ( .A1(n1390), .A2(n1222), .B1(n1221), .B2(n4), .ZN(n1013) );
  OAI22_X1 U1824 ( .A1(n29), .A2(n1146), .B1(n27), .B2(n1145), .ZN(n940) );
  OAI22_X1 U1825 ( .A1(n18), .A2(n1186), .B1(n16), .B2(n1185), .ZN(n978) );
  OAI22_X1 U1826 ( .A1(n1390), .A2(n1224), .B1(n1223), .B2(n4), .ZN(n1015) );
  OAI22_X1 U1827 ( .A1(n29), .A2(n1148), .B1(n27), .B2(n1147), .ZN(n942) );
  OAI22_X1 U1828 ( .A1(n1390), .A2(n1228), .B1(n1227), .B2(n4), .ZN(n1019) );
  OAI22_X1 U1829 ( .A1(n29), .A2(n1152), .B1(n27), .B2(n1151), .ZN(n946) );
  OAI22_X1 U1830 ( .A1(n17), .A2(n1190), .B1(n15), .B2(n1189), .ZN(n982) );
  OAI22_X1 U1831 ( .A1(n5), .A2(n1231), .B1(n1230), .B2(n4), .ZN(n1022) );
  AND2_X1 U1832 ( .A1(n1420), .A2(n806), .ZN(n949) );
  OAI22_X1 U1833 ( .A1(n17), .A2(n1193), .B1(n15), .B2(n1192), .ZN(n985) );
  OAI22_X1 U1834 ( .A1(n48), .A2(n1074), .B1(n46), .B2(n1073), .ZN(n871) );
  OAI22_X1 U1835 ( .A1(n24), .A2(n1161), .B1(n22), .B2(n1160), .ZN(n954) );
  OAI22_X1 U1836 ( .A1(n53), .A2(n1066), .B1(n51), .B2(n1065), .ZN(n864) );
  OAI22_X1 U1837 ( .A1(n48), .A2(n1085), .B1(n45), .B2(n1084), .ZN(n882) );
  NAND2_X1 U1838 ( .A1(n787), .A2(n788), .ZN(n400) );
  INV_X1 U1839 ( .A(n1490), .ZN(n1292) );
  OAI22_X1 U1840 ( .A1(n48), .A2(n1292), .B1(n1092), .B2(n46), .ZN(n822) );
  OAI22_X1 U1841 ( .A1(n48), .A2(n1091), .B1(n45), .B2(n1090), .ZN(n888) );
  OR2_X1 U1842 ( .A1(n1492), .A2(n1292), .ZN(n1092) );
  INV_X1 U1843 ( .A(n790), .ZN(n830) );
  AOI21_X1 U1844 ( .B1(n60), .B2(n58), .A(n1030), .ZN(n790) );
  OAI22_X1 U1845 ( .A1(n42), .A2(n1293), .B1(n1113), .B2(n40), .ZN(n823) );
  OAI22_X1 U1846 ( .A1(n1112), .A2(n41), .B1(n39), .B2(n1111), .ZN(n908) );
  OR2_X1 U1847 ( .A1(n1491), .A2(n1293), .ZN(n1113) );
  INV_X1 U1848 ( .A(n33), .ZN(n803) );
  INV_X1 U1849 ( .A(n22), .ZN(n809) );
  INV_X1 U1850 ( .A(n39), .ZN(n800) );
  OR2_X1 U1851 ( .A1(n1492), .A2(n1290), .ZN(n1050) );
  OR2_X1 U1852 ( .A1(n1420), .A2(n1296), .ZN(n1176) );
  OR2_X1 U1853 ( .A1(n1420), .A2(n1297), .ZN(n1197) );
  OR2_X1 U1854 ( .A1(n1492), .A2(n1294), .ZN(n1134) );
  OAI22_X1 U1855 ( .A1(n54), .A2(n1053), .B1(n52), .B2(n1052), .ZN(n851) );
  INV_X1 U1856 ( .A(n796), .ZN(n870) );
  AOI21_X1 U1857 ( .B1(n1477), .B2(n46), .A(n1072), .ZN(n796) );
  OAI22_X1 U1858 ( .A1(n42), .A2(n1095), .B1(n40), .B2(n1094), .ZN(n891) );
  OAI22_X1 U1859 ( .A1(n60), .A2(n1038), .B1(n58), .B2(n1037), .ZN(n837) );
  INV_X1 U1860 ( .A(n802), .ZN(n910) );
  INV_X1 U1861 ( .A(n45), .ZN(n797) );
  INV_X1 U1862 ( .A(n27), .ZN(n806) );
  INV_X1 U1863 ( .A(n15), .ZN(n812) );
  INV_X1 U1864 ( .A(n51), .ZN(n794) );
  OAI22_X1 U1865 ( .A1(n1391), .A2(n1236), .B1(n1235), .B2(n4), .ZN(n1027) );
  OAI22_X1 U1866 ( .A1(n11), .A2(n1217), .B1(n9), .B2(n1216), .ZN(n1008) );
  XNOR2_X1 U1867 ( .A(n1415), .B(n1492), .ZN(n1217) );
  BUF_X1 U1868 ( .A(n43), .Z(n1490) );
  OAI22_X1 U1869 ( .A1(n5), .A2(n1299), .B1(n1239), .B2(n4), .ZN(n829) );
  OR2_X1 U1870 ( .A1(n1420), .A2(n1299), .ZN(n1239) );
  INV_X1 U1871 ( .A(n1384), .ZN(n1299) );
  XNOR2_X1 U1872 ( .A(n1490), .B(n1245), .ZN(n1077) );
  XNOR2_X1 U1873 ( .A(n1483), .B(n1252), .ZN(n1084) );
  XNOR2_X1 U1874 ( .A(n1490), .B(n1255), .ZN(n1087) );
  XNOR2_X1 U1875 ( .A(n1484), .B(n1253), .ZN(n1085) );
  XNOR2_X1 U1876 ( .A(n1483), .B(n1442), .ZN(n1072) );
  BUF_X2 U1877 ( .A(n1277), .Z(n17) );
  OAI22_X1 U1878 ( .A1(n36), .A2(n1133), .B1(n33), .B2(n1132), .ZN(n928) );
  OAI22_X1 U1879 ( .A1(n36), .A2(n1294), .B1(n1134), .B2(n34), .ZN(n824) );
  XNOR2_X1 U1880 ( .A(n31), .B(n1491), .ZN(n1133) );
  OAI22_X1 U1881 ( .A1(n17), .A2(n1196), .B1(n15), .B2(n1195), .ZN(n988) );
  OAI22_X1 U1882 ( .A1(n18), .A2(n1297), .B1(n1197), .B2(n16), .ZN(n827) );
  XNOR2_X1 U1883 ( .A(n13), .B(n1492), .ZN(n1196) );
  XNOR2_X1 U1884 ( .A(n1483), .B(n1248), .ZN(n1080) );
  XNOR2_X1 U1885 ( .A(n1483), .B(n1412), .ZN(n1082) );
  XNOR2_X1 U1886 ( .A(n1483), .B(n1247), .ZN(n1079) );
  XNOR2_X1 U1887 ( .A(n1489), .B(n1249), .ZN(n1081) );
  XNOR2_X1 U1888 ( .A(n1484), .B(n1251), .ZN(n1083) );
  XNOR2_X1 U1889 ( .A(n1484), .B(n1244), .ZN(n1076) );
  XNOR2_X1 U1890 ( .A(n1483), .B(n1243), .ZN(n1075) );
  XNOR2_X1 U1891 ( .A(n1489), .B(n1246), .ZN(n1078) );
  XNOR2_X1 U1892 ( .A(n1489), .B(n1254), .ZN(n1086) );
  XNOR2_X1 U1893 ( .A(n1490), .B(n1257), .ZN(n1089) );
  XNOR2_X1 U1894 ( .A(n1490), .B(n1258), .ZN(n1090) );
  XNOR2_X1 U1895 ( .A(n1489), .B(n1242), .ZN(n1074) );
  XNOR2_X1 U1896 ( .A(n1484), .B(n1417), .ZN(n1073) );
  XNOR2_X1 U1897 ( .A(n55), .B(n1256), .ZN(n1046) );
  XNOR2_X1 U1898 ( .A(n55), .B(n1257), .ZN(n1047) );
  XNOR2_X1 U1899 ( .A(n13), .B(n1385), .ZN(n1179) );
  XNOR2_X1 U1900 ( .A(n13), .B(n1243), .ZN(n1180) );
  XNOR2_X1 U1901 ( .A(n19), .B(n1241), .ZN(n1157) );
  XNOR2_X1 U1902 ( .A(n31), .B(n1245), .ZN(n1119) );
  XNOR2_X1 U1903 ( .A(n55), .B(n1254), .ZN(n1044) );
  XNOR2_X1 U1904 ( .A(n55), .B(n1253), .ZN(n1043) );
  XNOR2_X1 U1905 ( .A(n31), .B(n1244), .ZN(n1118) );
  XNOR2_X1 U1906 ( .A(n31), .B(n1246), .ZN(n1120) );
  XNOR2_X1 U1907 ( .A(n55), .B(n1252), .ZN(n1042) );
  XNOR2_X1 U1908 ( .A(n19), .B(n1242), .ZN(n1158) );
  XNOR2_X1 U1909 ( .A(n55), .B(n1251), .ZN(n1041) );
  XNOR2_X1 U1910 ( .A(n13), .B(n1241), .ZN(n1178) );
  XNOR2_X1 U1911 ( .A(n55), .B(n1255), .ZN(n1045) );
  XNOR2_X1 U1912 ( .A(n19), .B(n1243), .ZN(n1159) );
  XNOR2_X1 U1913 ( .A(n31), .B(n1243), .ZN(n1117) );
  XNOR2_X1 U1914 ( .A(n55), .B(n1248), .ZN(n1038) );
  XNOR2_X1 U1915 ( .A(n31), .B(n1247), .ZN(n1121) );
  XNOR2_X1 U1916 ( .A(n31), .B(n1249), .ZN(n1123) );
  XNOR2_X1 U1917 ( .A(n19), .B(n1244), .ZN(n1160) );
  XNOR2_X1 U1918 ( .A(n55), .B(n1247), .ZN(n1037) );
  XNOR2_X1 U1919 ( .A(n1421), .B(n55), .ZN(n1040) );
  XNOR2_X1 U1920 ( .A(n31), .B(n1385), .ZN(n1116) );
  XNOR2_X1 U1921 ( .A(n19), .B(n1248), .ZN(n1164) );
  XNOR2_X1 U1922 ( .A(n19), .B(n1247), .ZN(n1163) );
  XNOR2_X1 U1923 ( .A(n1444), .B(n1417), .ZN(n1115) );
  XNOR2_X1 U1924 ( .A(n31), .B(n1250), .ZN(n1124) );
  XNOR2_X1 U1925 ( .A(n19), .B(n1255), .ZN(n1171) );
  XNOR2_X1 U1926 ( .A(n13), .B(n1251), .ZN(n1188) );
  XNOR2_X1 U1927 ( .A(n7), .B(n1246), .ZN(n1204) );
  XNOR2_X1 U1928 ( .A(n13), .B(n1246), .ZN(n1183) );
  XNOR2_X1 U1929 ( .A(n31), .B(n1248), .ZN(n1122) );
  XNOR2_X1 U1930 ( .A(n7), .B(n1241), .ZN(n1199) );
  XNOR2_X1 U1931 ( .A(n13), .B(n1252), .ZN(n1189) );
  XNOR2_X1 U1932 ( .A(n55), .B(n1258), .ZN(n1048) );
  XNOR2_X1 U1933 ( .A(n31), .B(n1251), .ZN(n1125) );
  XNOR2_X1 U1934 ( .A(n7), .B(n1242), .ZN(n1200) );
  XNOR2_X1 U1935 ( .A(n13), .B(n1245), .ZN(n1182) );
  XNOR2_X1 U1936 ( .A(n7), .B(n1250), .ZN(n1208) );
  XNOR2_X1 U1937 ( .A(n55), .B(n1249), .ZN(n1039) );
  XNOR2_X1 U1938 ( .A(n13), .B(n1247), .ZN(n1184) );
  XNOR2_X1 U1939 ( .A(n19), .B(n1254), .ZN(n1170) );
  XNOR2_X1 U1940 ( .A(n31), .B(n1252), .ZN(n1126) );
  XNOR2_X1 U1941 ( .A(n19), .B(n1249), .ZN(n1165) );
  XNOR2_X1 U1942 ( .A(n7), .B(n1247), .ZN(n1205) );
  XNOR2_X1 U1943 ( .A(n13), .B(n1244), .ZN(n1181) );
  XNOR2_X1 U1944 ( .A(n7), .B(n1243), .ZN(n1201) );
  XNOR2_X1 U1945 ( .A(n1415), .B(n1251), .ZN(n1209) );
  XNOR2_X1 U1946 ( .A(n19), .B(n1251), .ZN(n1167) );
  XNOR2_X1 U1947 ( .A(n31), .B(n1253), .ZN(n1127) );
  XNOR2_X1 U1948 ( .A(n19), .B(n1246), .ZN(n1162) );
  XNOR2_X1 U1949 ( .A(n31), .B(n1254), .ZN(n1128) );
  XNOR2_X1 U1950 ( .A(n13), .B(n1250), .ZN(n1187) );
  XNOR2_X1 U1951 ( .A(n19), .B(n1250), .ZN(n1166) );
  XNOR2_X1 U1952 ( .A(n19), .B(n1257), .ZN(n1173) );
  XNOR2_X1 U1953 ( .A(n7), .B(n1244), .ZN(n1202) );
  XNOR2_X1 U1954 ( .A(n31), .B(n1255), .ZN(n1129) );
  XNOR2_X1 U1955 ( .A(n1257), .B(n31), .ZN(n1131) );
  XNOR2_X1 U1956 ( .A(n55), .B(n1246), .ZN(n1036) );
  XNOR2_X1 U1957 ( .A(n7), .B(n1253), .ZN(n1211) );
  XNOR2_X1 U1958 ( .A(n7), .B(n1245), .ZN(n1203) );
  XNOR2_X1 U1959 ( .A(n13), .B(n1249), .ZN(n1186) );
  XNOR2_X1 U1960 ( .A(n19), .B(n1245), .ZN(n1161) );
  XNOR2_X1 U1961 ( .A(n19), .B(n1252), .ZN(n1168) );
  XNOR2_X1 U1962 ( .A(n31), .B(n1256), .ZN(n1130) );
  XNOR2_X1 U1963 ( .A(n13), .B(n1248), .ZN(n1185) );
  XNOR2_X1 U1964 ( .A(n19), .B(n1258), .ZN(n1174) );
  XNOR2_X1 U1965 ( .A(n19), .B(n1253), .ZN(n1169) );
  XNOR2_X1 U1966 ( .A(n31), .B(n1258), .ZN(n1132) );
  XNOR2_X1 U1967 ( .A(n7), .B(n1249), .ZN(n1207) );
  XNOR2_X1 U1968 ( .A(n1415), .B(n1254), .ZN(n1212) );
  XNOR2_X1 U1969 ( .A(n19), .B(n1256), .ZN(n1172) );
  XNOR2_X1 U1970 ( .A(n13), .B(n1258), .ZN(n1195) );
  XNOR2_X1 U1971 ( .A(n13), .B(n1257), .ZN(n1194) );
  XNOR2_X1 U1972 ( .A(n7), .B(n1248), .ZN(n1206) );
  XNOR2_X1 U1973 ( .A(n13), .B(n1253), .ZN(n1190) );
  XNOR2_X1 U1974 ( .A(n13), .B(n1254), .ZN(n1191) );
  XNOR2_X1 U1975 ( .A(n7), .B(n1252), .ZN(n1210) );
  XNOR2_X1 U1976 ( .A(n13), .B(n1255), .ZN(n1192) );
  XNOR2_X1 U1977 ( .A(n13), .B(n1256), .ZN(n1193) );
  XNOR2_X1 U1978 ( .A(n7), .B(n1256), .ZN(n1214) );
  XNOR2_X1 U1979 ( .A(n7), .B(n1257), .ZN(n1215) );
  XNOR2_X1 U1980 ( .A(n7), .B(n1255), .ZN(n1213) );
  XNOR2_X1 U1981 ( .A(n7), .B(n1258), .ZN(n1216) );
  XNOR2_X1 U1982 ( .A(n55), .B(n1244), .ZN(n1034) );
  XNOR2_X1 U1983 ( .A(n55), .B(n1245), .ZN(n1035) );
  XNOR2_X1 U1984 ( .A(n55), .B(n1243), .ZN(n1033) );
  XNOR2_X1 U1985 ( .A(n55), .B(n1242), .ZN(n1032) );
  XNOR2_X1 U1986 ( .A(n55), .B(n1417), .ZN(n1031) );
  OAI22_X1 U1987 ( .A1(n5), .A2(n1238), .B1(n1237), .B2(n4), .ZN(n1029) );
  BUF_X1 U1988 ( .A(n1288), .Z(n9) );
  XNOR2_X1 U1989 ( .A(n19), .B(n1240), .ZN(n1156) );
  XNOR2_X1 U1990 ( .A(n13), .B(n1240), .ZN(n1177) );
  XNOR2_X1 U1991 ( .A(n1444), .B(n1419), .ZN(n1114) );
  XNOR2_X1 U1992 ( .A(n7), .B(n1240), .ZN(n1198) );
  XNOR2_X1 U1993 ( .A(n55), .B(n1442), .ZN(n1030) );
  BUF_X1 U1994 ( .A(n1288), .Z(n10) );
  BUF_X1 U1995 ( .A(n1281), .Z(n52) );
  BUF_X1 U1996 ( .A(n1271), .Z(n54) );
  BUF_X2 U1997 ( .A(n1279), .Z(n6) );
  BUF_X1 U1998 ( .A(n1278), .Z(n11) );
  OAI22_X1 U1999 ( .A1(n59), .A2(n1049), .B1(n1481), .B2(n1438), .ZN(n848) );
  OAI22_X1 U2000 ( .A1(n60), .A2(n1290), .B1(n1050), .B2(n58), .ZN(n820) );
  XNOR2_X1 U2001 ( .A(n55), .B(n1420), .ZN(n1049) );
  OAI22_X1 U2002 ( .A1(n23), .A2(n1175), .B1(n1443), .B2(n1174), .ZN(n968) );
  OAI22_X1 U2003 ( .A1(n24), .A2(n1296), .B1(n1176), .B2(n1443), .ZN(n826) );
  XNOR2_X1 U2004 ( .A(n19), .B(n1492), .ZN(n1175) );
  INV_X1 U2005 ( .A(n49), .ZN(n1291) );
  INV_X1 U2006 ( .A(n37), .ZN(n1293) );
  OAI22_X1 U2007 ( .A1(n11), .A2(n1298), .B1(n1218), .B2(n10), .ZN(n828) );
  OR2_X1 U2008 ( .A1(n1420), .A2(n1298), .ZN(n1218) );
  INV_X1 U2009 ( .A(n7), .ZN(n1298) );
  BUF_X2 U2010 ( .A(n1274), .Z(n35) );
  INV_X1 U2011 ( .A(n31), .ZN(n1294) );
  INV_X1 U2012 ( .A(n19), .ZN(n1296) );
  INV_X1 U2013 ( .A(n13), .ZN(n1297) );
  INV_X1 U2014 ( .A(n55), .ZN(n1290) );
  INV_X1 U2015 ( .A(n25), .ZN(n1295) );
  XNOR2_X1 U2016 ( .A(a[2]), .B(a[1]), .ZN(n1288) );
  XNOR2_X1 U2017 ( .A(a[16]), .B(a[15]), .ZN(n1281) );
  BUF_X4 U2018 ( .A(a[5]), .Z(n13) );
  BUF_X4 U2019 ( .A(a[7]), .Z(n19) );
  BUF_X4 U2020 ( .A(a[11]), .Z(n31) );
  BUF_X4 U2021 ( .A(a[3]), .Z(n7) );
  CLKBUF_X3 U2022 ( .A(b[8]), .Z(n1251) );
  CLKBUF_X3 U2023 ( .A(b[3]), .Z(n1256) );
  NAND2_X1 U2024 ( .A1(n1268), .A2(n1288), .ZN(n1278) );
  NAND2_X1 U2025 ( .A1(n767), .A2(n772), .ZN(n384) );
  CLKBUF_X1 U2026 ( .A(n43), .Z(n1489) );
  BUF_X2 U2027 ( .A(n291), .Z(n64) );
  INV_X1 U2028 ( .A(n303), .ZN(n302) );
  OAI22_X1 U2029 ( .A1(n54), .A2(n1052), .B1(n52), .B2(n1051), .ZN(n454) );
  INV_X1 U2030 ( .A(n361), .ZN(n436) );
  OAI21_X1 U2031 ( .B1(n361), .B2(n365), .A(n362), .ZN(n360) );
  NOR2_X1 U2032 ( .A1(n361), .A2(n364), .ZN(n359) );
  NAND2_X1 U2033 ( .A1(n294), .A2(n310), .ZN(n292) );
  AOI21_X1 U2034 ( .B1(n340), .B2(n321), .A(n322), .ZN(n320) );
  OAI21_X1 U2035 ( .B1(n341), .B2(n358), .A(n342), .ZN(n340) );
  AOI21_X1 U2036 ( .B1(n349), .B2(n1457), .A(n344), .ZN(n342) );
  XNOR2_X1 U2037 ( .A(n319), .B(n86), .ZN(product[19]) );
  OAI21_X1 U2038 ( .B1(n251), .B2(n276), .A(n252), .ZN(n250) );
  NAND2_X1 U2039 ( .A1(n1265), .A2(n1285), .ZN(n1275) );
  OAI22_X1 U2040 ( .A1(n41), .A2(n1104), .B1(n39), .B2(n1103), .ZN(n900) );
  NAND2_X1 U2041 ( .A1(n1263), .A2(n1283), .ZN(n1273) );
  XNOR2_X1 U2042 ( .A(n25), .B(n1420), .ZN(n1154) );
  XNOR2_X1 U2043 ( .A(n25), .B(n1254), .ZN(n1149) );
  XNOR2_X1 U2044 ( .A(n25), .B(n1258), .ZN(n1153) );
  XNOR2_X1 U2045 ( .A(n25), .B(n1257), .ZN(n1152) );
  XNOR2_X1 U2046 ( .A(n1256), .B(n1435), .ZN(n1151) );
  XNOR2_X1 U2047 ( .A(n1435), .B(n1255), .ZN(n1150) );
  XNOR2_X1 U2048 ( .A(n1435), .B(n1250), .ZN(n1145) );
  XNOR2_X1 U2049 ( .A(n25), .B(n1246), .ZN(n1141) );
  XNOR2_X1 U2050 ( .A(n1435), .B(n1247), .ZN(n1142) );
  XNOR2_X1 U2051 ( .A(n25), .B(n1253), .ZN(n1148) );
  XNOR2_X1 U2052 ( .A(n1435), .B(n1245), .ZN(n1140) );
  XNOR2_X1 U2053 ( .A(n1435), .B(n1249), .ZN(n1144) );
  XNOR2_X1 U2054 ( .A(n1435), .B(n1248), .ZN(n1143) );
  XNOR2_X1 U2055 ( .A(n25), .B(n1244), .ZN(n1139) );
  XNOR2_X1 U2056 ( .A(n1435), .B(n1252), .ZN(n1147) );
  XNOR2_X1 U2057 ( .A(n1435), .B(n1251), .ZN(n1146) );
  XNOR2_X1 U2058 ( .A(n1435), .B(n1243), .ZN(n1138) );
  XNOR2_X1 U2059 ( .A(n25), .B(n1240), .ZN(n1135) );
  XNOR2_X1 U2060 ( .A(n1435), .B(n1385), .ZN(n1137) );
  XNOR2_X1 U2061 ( .A(n1435), .B(n1241), .ZN(n1136) );
  OAI21_X1 U2062 ( .B1(n217), .B2(n121), .A(n122), .ZN(n120) );
  OAI21_X1 U2063 ( .B1(n217), .B2(n192), .A(n193), .ZN(n187) );
  NOR2_X1 U2064 ( .A1(n229), .A2(n220), .ZN(n218) );
  INV_X1 U2065 ( .A(a[0]), .ZN(n1289) );
  NAND2_X1 U2066 ( .A1(n1269), .A2(n1289), .ZN(n1279) );
  BUF_X2 U2067 ( .A(n1289), .Z(n4) );
  INV_X1 U2068 ( .A(n817), .ZN(n1010) );
  INV_X1 U2069 ( .A(n1454), .ZN(n280) );
  INV_X1 U2070 ( .A(n289), .ZN(n287) );
  OAI21_X1 U2071 ( .B1(n339), .B2(n326), .A(n1482), .ZN(n325) );
  OAI21_X1 U2072 ( .B1(n327), .B2(n323), .A(n324), .ZN(n322) );
  XNOR2_X1 U2073 ( .A(n1440), .B(n1243), .ZN(n1096) );
  XNOR2_X1 U2074 ( .A(n1440), .B(n1419), .ZN(n1093) );
  XNOR2_X1 U2075 ( .A(n37), .B(n1253), .ZN(n1106) );
  XNOR2_X1 U2076 ( .A(n1440), .B(n1385), .ZN(n1095) );
  XNOR2_X1 U2077 ( .A(n1440), .B(n1417), .ZN(n1094) );
  XNOR2_X1 U2078 ( .A(n37), .B(n1252), .ZN(n1105) );
  XNOR2_X1 U2079 ( .A(n37), .B(n1249), .ZN(n1102) );
  XNOR2_X1 U2080 ( .A(n37), .B(n1254), .ZN(n1107) );
  XNOR2_X1 U2081 ( .A(n1386), .B(n1245), .ZN(n1098) );
  XNOR2_X1 U2082 ( .A(n37), .B(n1257), .ZN(n1110) );
  XNOR2_X1 U2083 ( .A(n1386), .B(n1244), .ZN(n1097) );
  XNOR2_X1 U2084 ( .A(n1256), .B(n37), .ZN(n1109) );
  XNOR2_X1 U2085 ( .A(n37), .B(n1491), .ZN(n1112) );
  XNOR2_X1 U2086 ( .A(n37), .B(n1255), .ZN(n1108) );
  XNOR2_X1 U2087 ( .A(n37), .B(n1258), .ZN(n1111) );
  XNOR2_X1 U2088 ( .A(n1386), .B(n1248), .ZN(n1101) );
  XNOR2_X1 U2089 ( .A(n37), .B(n1247), .ZN(n1100) );
  XNOR2_X1 U2090 ( .A(n37), .B(n1246), .ZN(n1099) );
  XNOR2_X1 U2091 ( .A(n37), .B(n1251), .ZN(n1104) );
  XNOR2_X1 U2092 ( .A(n37), .B(n1250), .ZN(n1103) );
  XNOR2_X1 U2093 ( .A(a[14]), .B(a[13]), .ZN(n1282) );
  BUF_X4 U2094 ( .A(a[13]), .Z(n37) );
  XNOR2_X1 U2095 ( .A(n385), .B(n97), .ZN(product[8]) );
  NAND2_X1 U2096 ( .A1(n1266), .A2(n1286), .ZN(n1276) );
  AOI21_X1 U2097 ( .B1(n357), .B2(n348), .A(n349), .ZN(n347) );
  NAND2_X1 U2098 ( .A1(n348), .A2(n1457), .ZN(n341) );
  AOI21_X1 U2099 ( .B1(n283), .B2(n249), .A(n250), .ZN(n248) );
  OAI21_X1 U2100 ( .B1(n284), .B2(n290), .A(n285), .ZN(n283) );
  BUF_X2 U2101 ( .A(n1277), .Z(n18) );
  NAND2_X1 U2102 ( .A1(n1267), .A2(n1287), .ZN(n1277) );
  XOR2_X1 U2103 ( .A(n388), .B(n98), .Z(product[7]) );
  OAI21_X1 U2104 ( .B1(n296), .B2(n304), .A(n297), .ZN(n295) );
  NOR2_X1 U2105 ( .A1(n1478), .A2(n303), .ZN(n294) );
  INV_X1 U2106 ( .A(n1446), .ZN(n426) );
  XOR2_X1 U2107 ( .A(n157), .B(n70), .Z(product[35]) );
  OAI21_X1 U2108 ( .B1(n292), .B2(n320), .A(n293), .ZN(n291) );
  BUF_X2 U2109 ( .A(n291), .Z(n63) );
  XNOR2_X1 U2110 ( .A(n49), .B(n1243), .ZN(n1054) );
  XNOR2_X1 U2111 ( .A(n49), .B(n1385), .ZN(n1053) );
  XNOR2_X1 U2112 ( .A(n49), .B(n1247), .ZN(n1058) );
  XNOR2_X1 U2113 ( .A(n49), .B(n1246), .ZN(n1057) );
  XNOR2_X1 U2114 ( .A(n49), .B(n1244), .ZN(n1055) );
  XNOR2_X1 U2115 ( .A(n49), .B(n1245), .ZN(n1056) );
  XNOR2_X1 U2116 ( .A(n49), .B(n1491), .ZN(n1070) );
  XNOR2_X1 U2117 ( .A(n49), .B(n1253), .ZN(n1064) );
  XNOR2_X1 U2118 ( .A(n49), .B(n1257), .ZN(n1068) );
  XNOR2_X1 U2119 ( .A(n49), .B(n1256), .ZN(n1067) );
  XNOR2_X1 U2120 ( .A(n49), .B(n1258), .ZN(n1069) );
  XNOR2_X1 U2121 ( .A(n49), .B(n1248), .ZN(n1059) );
  XNOR2_X1 U2122 ( .A(n49), .B(n1252), .ZN(n1063) );
  XNOR2_X1 U2123 ( .A(n49), .B(n1251), .ZN(n1062) );
  XNOR2_X1 U2124 ( .A(n49), .B(n1250), .ZN(n1061) );
  XNOR2_X1 U2125 ( .A(n49), .B(n1249), .ZN(n1060) );
  XNOR2_X1 U2126 ( .A(n49), .B(n1255), .ZN(n1066) );
  XNOR2_X1 U2127 ( .A(n49), .B(n1254), .ZN(n1065) );
  XNOR2_X1 U2128 ( .A(n49), .B(n1417), .ZN(n1052) );
  XNOR2_X1 U2129 ( .A(n49), .B(n1442), .ZN(n1051) );
  XNOR2_X1 U2130 ( .A(a[18]), .B(a[17]), .ZN(n1280) );
  BUF_X4 U2131 ( .A(a[17]), .Z(n49) );
  NOR2_X1 U2132 ( .A1(n251), .A2(n275), .ZN(n249) );
  NAND2_X1 U2133 ( .A1(n1480), .A2(n1471), .ZN(n251) );
  AOI21_X1 U2134 ( .B1(n6), .B2(n4), .A(n1219), .ZN(n817) );
  XNOR2_X1 U2135 ( .A(n1384), .B(n1251), .ZN(n1230) );
  XNOR2_X1 U2136 ( .A(n1384), .B(n1252), .ZN(n1231) );
  XNOR2_X1 U2137 ( .A(n1384), .B(n1248), .ZN(n1227) );
  XNOR2_X1 U2138 ( .A(n1384), .B(n1250), .ZN(n1229) );
  XNOR2_X1 U2139 ( .A(n1384), .B(n1249), .ZN(n1228) );
  XNOR2_X1 U2140 ( .A(n1), .B(n1242), .ZN(n1221) );
  XNOR2_X1 U2141 ( .A(n1), .B(n1241), .ZN(n1220) );
  XNOR2_X1 U2142 ( .A(n1384), .B(n1247), .ZN(n1226) );
  XNOR2_X1 U2143 ( .A(n1384), .B(n1246), .ZN(n1225) );
  XNOR2_X1 U2144 ( .A(n1384), .B(n1253), .ZN(n1232) );
  XNOR2_X1 U2145 ( .A(n1384), .B(n1254), .ZN(n1233) );
  XNOR2_X1 U2146 ( .A(n1384), .B(n1245), .ZN(n1224) );
  XNOR2_X1 U2147 ( .A(n1), .B(n1244), .ZN(n1223) );
  XNOR2_X1 U2148 ( .A(n1), .B(n1243), .ZN(n1222) );
  XNOR2_X1 U2149 ( .A(n1384), .B(n1492), .ZN(n1238) );
  XNOR2_X1 U2150 ( .A(n1384), .B(n1256), .ZN(n1235) );
  XNOR2_X1 U2151 ( .A(n1384), .B(n1255), .ZN(n1234) );
  XNOR2_X1 U2152 ( .A(n1), .B(n1240), .ZN(n1219) );
  XNOR2_X1 U2153 ( .A(n1384), .B(n1258), .ZN(n1237) );
  XNOR2_X1 U2154 ( .A(n1384), .B(n1257), .ZN(n1236) );
  OAI22_X1 U2155 ( .A1(n1390), .A2(n1237), .B1(n1236), .B2(n4), .ZN(n1028) );
  XOR2_X1 U2156 ( .A(a[8]), .B(a[9]), .Z(n1265) );
  XNOR2_X1 U2157 ( .A(a[10]), .B(a[9]), .ZN(n1284) );
  XNOR2_X1 U2158 ( .A(a[4]), .B(a[3]), .ZN(n1287) );
  XOR2_X1 U2159 ( .A(a[2]), .B(a[3]), .Z(n1268) );
  XNOR2_X1 U2160 ( .A(a[8]), .B(a[7]), .ZN(n1285) );
  XOR2_X1 U2161 ( .A(a[6]), .B(a[7]), .Z(n1266) );
  XOR2_X1 U2162 ( .A(a[4]), .B(a[5]), .Z(n1267) );
  XNOR2_X1 U2163 ( .A(a[6]), .B(a[5]), .ZN(n1286) );
  XOR2_X1 U2164 ( .A(a[18]), .B(a[19]), .Z(n1260) );
  AOI21_X1 U2165 ( .B1(n1448), .B2(n106), .A(n107), .ZN(n105) );
  AOI21_X1 U2166 ( .B1(n64), .B2(n115), .A(n116), .ZN(n114) );
  AOI21_X1 U2167 ( .B1(n64), .B2(n128), .A(n129), .ZN(n127) );
  AOI21_X1 U2168 ( .B1(n64), .B2(n199), .A(n200), .ZN(n198) );
  AOI21_X1 U2169 ( .B1(n64), .B2(n182), .A(n183), .ZN(n181) );
  AOI21_X1 U2170 ( .B1(n63), .B2(n210), .A(n211), .ZN(n209) );
  AOI21_X1 U2171 ( .B1(n64), .B2(n169), .A(n170), .ZN(n168) );
  AOI21_X1 U2172 ( .B1(n64), .B2(n143), .A(n144), .ZN(n142) );
  AOI21_X1 U2173 ( .B1(n64), .B2(n158), .A(n159), .ZN(n157) );
  XOR2_X1 U2174 ( .A(a[10]), .B(a[11]), .Z(n1264) );
  XNOR2_X1 U2175 ( .A(a[11]), .B(a[12]), .ZN(n1283) );
  XOR2_X1 U2176 ( .A(a[14]), .B(a[15]), .Z(n1262) );
  NOR2_X1 U2177 ( .A1(n350), .A2(n355), .ZN(n348) );
  OAI21_X1 U2178 ( .B1(n350), .B2(n356), .A(n351), .ZN(n349) );
  XOR2_X1 U2179 ( .A(a[12]), .B(a[13]), .Z(n1263) );
  XNOR2_X1 U2180 ( .A(n99), .B(n393), .ZN(product[6]) );
  AOI21_X1 U2181 ( .B1(n63), .B2(n223), .A(n224), .ZN(n222) );
  AOI21_X1 U2182 ( .B1(n64), .B2(n232), .A(n233), .ZN(n231) );
  AOI21_X1 U2183 ( .B1(n64), .B2(n245), .A(n246), .ZN(n244) );
  XNOR2_X1 U2184 ( .A(n64), .B(n82), .ZN(product[23]) );
  AOI21_X1 U2185 ( .B1(n63), .B2(n1454), .A(n279), .ZN(n277) );
  AOI21_X1 U2186 ( .B1(n63), .B2(n287), .A(n288), .ZN(n286) );
  AOI21_X1 U2187 ( .B1(n63), .B2(n258), .A(n259), .ZN(n257) );
  AOI21_X1 U2188 ( .B1(n63), .B2(n269), .A(n270), .ZN(n268) );
  XOR2_X1 U2189 ( .A(a[16]), .B(a[17]), .Z(n1261) );
  NOR2_X1 U2190 ( .A1(n289), .A2(n1475), .ZN(n282) );
  XOR2_X1 U2191 ( .A(a[0]), .B(a[1]), .Z(n1269) );
endmodule


module datapath_DW_mult_tc_13 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n15, n16, n17, n18,
         n19, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34, n35,
         n36, n37, n40, n41, n42, n43, n45, n46, n47, n48, n49, n51, n52, n53,
         n54, n55, n57, n58, n59, n60, n61, n63, n64, n66, n67, n68, n69, n70,
         n71, n72, n73, n82, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n105, n106, n107, n108,
         n109, n111, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n124, n126, n127, n128, n129, n130, n131, n134, n135, n136,
         n137, n139, n141, n142, n143, n144, n145, n146, n149, n150, n151,
         n152, n154, n156, n157, n158, n159, n160, n161, n165, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n190, n191, n192,
         n193, n195, n197, n198, n199, n200, n201, n202, n206, n208, n209,
         n210, n211, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n264, n265, n266, n267, n268, n269, n270, n273, n274, n275, n276,
         n277, n280, n281, n282, n283, n284, n285, n286, n288, n289, n290,
         n291, n292, n293, n294, n295, n297, n298, n299, n300, n302, n303,
         n304, n305, n306, n309, n310, n311, n313, n314, n316, n317, n318,
         n319, n320, n321, n322, n324, n325, n326, n327, n331, n332, n336,
         n337, n338, n339, n340, n341, n342, n344, n346, n347, n348, n349,
         n350, n351, n352, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n371, n373, n374,
         n376, n378, n379, n380, n382, n384, n385, n386, n387, n388, n390,
         n392, n393, n394, n395, n396, n398, n400, n401, n402, n403, n404,
         n405, n406, n407, n409, n418, n424, n425, n426, n428, n429, n432,
         n434, n435, n436, n437, n441, n443, n445, n446, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n793, n794, n796, n797, n799, n800, n802, n803, n805, n806, n808,
         n809, n811, n812, n814, n815, n817, n818, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1549, n1550;
  assign product[39] = n105;

  FA_X1 U488 ( .A(n831), .B(n454), .CI(n850), .CO(n450), .S(n451) );
  FA_X1 U489 ( .A(n455), .B(n832), .CI(n458), .CO(n452), .S(n453) );
  FA_X1 U491 ( .A(n462), .B(n833), .CI(n459), .CO(n456), .S(n457) );
  FA_X1 U492 ( .A(n851), .B(n464), .CI(n870), .CO(n458), .S(n459) );
  FA_X1 U493 ( .A(n463), .B(n470), .CI(n468), .CO(n460), .S(n461) );
  FA_X1 U494 ( .A(n834), .B(n852), .CI(n465), .CO(n462), .S(n463) );
  FA_X1 U496 ( .A(n474), .B(n471), .CI(n469), .CO(n466), .S(n467) );
  FA_X1 U497 ( .A(n478), .B(n871), .CI(n476), .CO(n468), .S(n469) );
  FA_X1 U498 ( .A(n853), .B(n835), .CI(n890), .CO(n470), .S(n471) );
  FA_X1 U499 ( .A(n475), .B(n477), .CI(n482), .CO(n472), .S(n473) );
  FA_X1 U500 ( .A(n486), .B(n479), .CI(n484), .CO(n474), .S(n475) );
  FA_X1 U501 ( .A(n836), .B(n854), .CI(n872), .CO(n476), .S(n477) );
  FA_X1 U503 ( .A(n490), .B(n492), .CI(n483), .CO(n480), .S(n481) );
  FA_X1 U504 ( .A(n485), .B(n494), .CI(n487), .CO(n482), .S(n483) );
  FA_X1 U505 ( .A(n855), .B(n496), .CI(n873), .CO(n484), .S(n485) );
  FA_X1 U506 ( .A(n891), .B(n837), .CI(n910), .CO(n486), .S(n487) );
  FA_X1 U507 ( .A(n500), .B(n493), .CI(n491), .CO(n488), .S(n489) );
  FA_X1 U508 ( .A(n495), .B(n504), .CI(n502), .CO(n490), .S(n491) );
  FA_X1 U509 ( .A(n497), .B(n874), .CI(n506), .CO(n492), .S(n493) );
  FA_X1 U510 ( .A(n892), .B(n856), .CI(n838), .CO(n494), .S(n495) );
  FA_X1 U512 ( .A(n510), .B(n503), .CI(n501), .CO(n498), .S(n499) );
  FA_X1 U513 ( .A(n507), .B(n505), .CI(n512), .CO(n500), .S(n501) );
  FA_X1 U514 ( .A(n516), .B(n893), .CI(n514), .CO(n502), .S(n503) );
  FA_X1 U515 ( .A(n857), .B(n911), .CI(n875), .CO(n504), .S(n505) );
  FA_X1 U516 ( .A(n518), .B(n839), .CI(n930), .CO(n506), .S(n507) );
  FA_X1 U517 ( .A(n522), .B(n513), .CI(n511), .CO(n508), .S(n509) );
  FA_X1 U518 ( .A(n526), .B(n515), .CI(n524), .CO(n510), .S(n511) );
  FA_X1 U519 ( .A(n528), .B(n530), .CI(n517), .CO(n512), .S(n513) );
  FA_X1 U520 ( .A(n840), .B(n858), .CI(n519), .CO(n514), .S(n515) );
  FA_X1 U521 ( .A(n912), .B(n876), .CI(n894), .CO(n516), .S(n517) );
  FA_X1 U523 ( .A(n523), .B(n525), .CI(n534), .CO(n520), .S(n521) );
  FA_X1 U524 ( .A(n527), .B(n538), .CI(n536), .CO(n522), .S(n523) );
  FA_X1 U525 ( .A(n529), .B(n540), .CI(n531), .CO(n524), .S(n525) );
  FA_X1 U526 ( .A(n877), .B(n895), .CI(n542), .CO(n526), .S(n527) );
  FA_X1 U527 ( .A(n859), .B(n931), .CI(n913), .CO(n528), .S(n529) );
  FA_X1 U528 ( .A(n544), .B(n841), .CI(n950), .CO(n530), .S(n531) );
  FA_X1 U529 ( .A(n535), .B(n537), .CI(n548), .CO(n532), .S(n533) );
  FA_X1 U530 ( .A(n539), .B(n552), .CI(n550), .CO(n534), .S(n535) );
  FA_X1 U531 ( .A(n541), .B(n554), .CI(n543), .CO(n536), .S(n537) );
  FA_X1 U532 ( .A(n558), .B(n545), .CI(n556), .CO(n538), .S(n539) );
  FA_X1 U533 ( .A(n896), .B(n932), .CI(n914), .CO(n540), .S(n541) );
  FA_X1 U534 ( .A(n878), .B(n842), .CI(n860), .CO(n542), .S(n543) );
  FA_X1 U536 ( .A(n562), .B(n551), .CI(n549), .CO(n546), .S(n547) );
  FA_X1 U537 ( .A(n553), .B(n566), .CI(n564), .CO(n548), .S(n549) );
  FA_X1 U538 ( .A(n559), .B(n557), .CI(n568), .CO(n550), .S(n551) );
  FA_X1 U539 ( .A(n570), .B(n572), .CI(n555), .CO(n552), .S(n553) );
  FA_X1 U540 ( .A(n879), .B(n915), .CI(n897), .CO(n554), .S(n555) );
  FA_X1 U541 ( .A(n861), .B(n951), .CI(n933), .CO(n556), .S(n557) );
  FA_X1 U542 ( .A(n574), .B(n843), .CI(n970), .CO(n558), .S(n559) );
  FA_X1 U543 ( .A(n578), .B(n565), .CI(n563), .CO(n560), .S(n561) );
  FA_X1 U544 ( .A(n567), .B(n582), .CI(n580), .CO(n562), .S(n563) );
  FA_X1 U546 ( .A(n586), .B(n588), .CI(n571), .CO(n566), .S(n567) );
  FA_X1 U548 ( .A(n844), .B(n916), .CI(n862), .CO(n570), .S(n571) );
  FA_X1 U549 ( .A(n952), .B(n880), .CI(n934), .CO(n572), .S(n573) );
  FA_X1 U552 ( .A(n583), .B(n598), .CI(n596), .CO(n578), .S(n579) );
  FA_X1 U553 ( .A(n600), .B(n591), .CI(n585), .CO(n580), .S(n581) );
  FA_X1 U554 ( .A(n587), .B(n602), .CI(n589), .CO(n582), .S(n583) );
  FA_X1 U555 ( .A(n606), .B(n917), .CI(n604), .CO(n584), .S(n585) );
  FA_X1 U556 ( .A(n881), .B(n935), .CI(n899), .CO(n586), .S(n587) );
  FA_X1 U557 ( .A(n608), .B(n953), .CI(n863), .CO(n588), .S(n589) );
  FA_X1 U559 ( .A(n612), .B(n597), .CI(n595), .CO(n592), .S(n593) );
  FA_X1 U560 ( .A(n599), .B(n616), .CI(n614), .CO(n594), .S(n595) );
  FA_X1 U561 ( .A(n618), .B(n603), .CI(n601), .CO(n596), .S(n597) );
  FA_X1 U562 ( .A(n605), .B(n620), .CI(n607), .CO(n598), .S(n599) );
  FA_X1 U563 ( .A(n624), .B(n626), .CI(n622), .CO(n600), .S(n601) );
  FA_X1 U564 ( .A(n918), .B(n936), .CI(n609), .CO(n602), .S(n603) );
  FA_X1 U565 ( .A(n954), .B(n864), .CI(n882), .CO(n604), .S(n605) );
  FA_X1 U566 ( .A(n972), .B(n900), .CI(n846), .CO(n606), .S(n607) );
  FA_X1 U569 ( .A(n617), .B(n634), .CI(n632), .CO(n612), .S(n613) );
  FA_X1 U571 ( .A(n623), .B(n638), .CI(n625), .CO(n616), .S(n617) );
  FA_X1 U572 ( .A(n627), .B(n642), .CI(n640), .CO(n618), .S(n619) );
  FA_X1 U573 ( .A(n955), .B(n973), .CI(n644), .CO(n620), .S(n621) );
  FA_X1 U574 ( .A(n991), .B(n901), .CI(n883), .CO(n622), .S(n623) );
  FA_X1 U575 ( .A(n847), .B(n919), .CI(n1010), .CO(n624), .S(n625) );
  FA_X1 U580 ( .A(n654), .B(n643), .CI(n652), .CO(n632), .S(n633) );
  FA_X1 U581 ( .A(n639), .B(n656), .CI(n641), .CO(n634), .S(n635) );
  FA_X1 U583 ( .A(n920), .B(n992), .CI(n974), .CO(n638), .S(n639) );
  FA_X1 U584 ( .A(n956), .B(n902), .CI(n1011), .CO(n640), .S(n641) );
  HA_X1 U586 ( .A(n820), .B(n848), .CO(n644), .S(n645) );
  FA_X1 U588 ( .A(n653), .B(n655), .CI(n666), .CO(n648), .S(n649) );
  FA_X1 U589 ( .A(n670), .B(n659), .CI(n668), .CO(n650), .S(n651) );
  FA_X1 U590 ( .A(n661), .B(n672), .CI(n657), .CO(n652), .S(n653) );
  FA_X1 U591 ( .A(n676), .B(n957), .CI(n674), .CO(n654), .S(n655) );
  FA_X1 U592 ( .A(n921), .B(n975), .CI(n939), .CO(n656), .S(n657) );
  FA_X1 U593 ( .A(n867), .B(n993), .CI(n903), .CO(n658), .S(n659) );
  FA_X1 U594 ( .A(n849), .B(n1012), .CI(n885), .CO(n660), .S(n661) );
  FA_X1 U595 ( .A(n667), .B(n680), .CI(n665), .CO(n662), .S(n663) );
  FA_X1 U596 ( .A(n669), .B(n671), .CI(n682), .CO(n664), .S(n665) );
  FA_X1 U597 ( .A(n675), .B(n673), .CI(n684), .CO(n666), .S(n667) );
  FA_X1 U598 ( .A(n688), .B(n690), .CI(n686), .CO(n668), .S(n669) );
  FA_X1 U599 ( .A(n958), .B(n976), .CI(n677), .CO(n670), .S(n671) );
  FA_X1 U600 ( .A(n886), .B(n904), .CI(n922), .CO(n672), .S(n673) );
  FA_X1 U601 ( .A(n1013), .B(n940), .CI(n994), .CO(n674), .S(n675) );
  HA_X1 U602 ( .A(n821), .B(n868), .CO(n676), .S(n677) );
  FA_X1 U604 ( .A(n696), .B(n698), .CI(n685), .CO(n680), .S(n681) );
  FA_X1 U605 ( .A(n689), .B(n691), .CI(n687), .CO(n682), .S(n683) );
  FA_X1 U606 ( .A(n702), .B(n704), .CI(n700), .CO(n684), .S(n685) );
  FA_X1 U607 ( .A(n941), .B(n977), .CI(n959), .CO(n686), .S(n687) );
  FA_X1 U608 ( .A(n995), .B(n887), .CI(n923), .CO(n688), .S(n689) );
  FA_X1 U609 ( .A(n905), .B(n869), .CI(n1014), .CO(n690), .S(n691) );
  FA_X1 U610 ( .A(n697), .B(n708), .CI(n695), .CO(n692), .S(n693) );
  FA_X1 U611 ( .A(n710), .B(n703), .CI(n699), .CO(n694), .S(n695) );
  FA_X1 U612 ( .A(n712), .B(n714), .CI(n701), .CO(n696), .S(n697) );
  FA_X1 U613 ( .A(n705), .B(n996), .CI(n716), .CO(n698), .S(n699) );
  FA_X1 U614 ( .A(n1015), .B(n942), .CI(n978), .CO(n700), .S(n701) );
  FA_X1 U615 ( .A(n960), .B(n924), .CI(n906), .CO(n702), .S(n703) );
  HA_X1 U616 ( .A(n822), .B(n888), .CO(n704), .S(n705) );
  FA_X1 U617 ( .A(n711), .B(n720), .CI(n709), .CO(n706), .S(n707) );
  FA_X1 U618 ( .A(n713), .B(n715), .CI(n722), .CO(n708), .S(n709) );
  FA_X1 U619 ( .A(n724), .B(n726), .CI(n717), .CO(n710), .S(n711) );
  FA_X1 U620 ( .A(n961), .B(n979), .CI(n728), .CO(n712), .S(n713) );
  FA_X1 U621 ( .A(n907), .B(n997), .CI(n943), .CO(n714), .S(n715) );
  FA_X1 U622 ( .A(n889), .B(n1016), .CI(n925), .CO(n716), .S(n717) );
  FA_X1 U623 ( .A(n732), .B(n723), .CI(n721), .CO(n718), .S(n719) );
  FA_X1 U624 ( .A(n727), .B(n725), .CI(n734), .CO(n720), .S(n721) );
  FA_X1 U625 ( .A(n738), .B(n729), .CI(n736), .CO(n722), .S(n723) );
  FA_X1 U626 ( .A(n926), .B(n980), .CI(n944), .CO(n724), .S(n725) );
  FA_X1 U627 ( .A(n1017), .B(n962), .CI(n998), .CO(n726), .S(n727) );
  HA_X1 U628 ( .A(n908), .B(n823), .CO(n728), .S(n729) );
  FA_X1 U629 ( .A(n735), .B(n742), .CI(n733), .CO(n730), .S(n731) );
  FA_X1 U630 ( .A(n737), .B(n739), .CI(n744), .CO(n732), .S(n733) );
  FA_X1 U631 ( .A(n748), .B(n981), .CI(n746), .CO(n734), .S(n735) );
  FA_X1 U632 ( .A(n927), .B(n999), .CI(n963), .CO(n736), .S(n737) );
  FA_X1 U633 ( .A(n945), .B(n909), .CI(n1018), .CO(n738), .S(n739) );
  FA_X1 U634 ( .A(n752), .B(n745), .CI(n743), .CO(n740), .S(n741) );
  FA_X1 U635 ( .A(n754), .B(n756), .CI(n747), .CO(n742), .S(n743) );
  FA_X1 U636 ( .A(n964), .B(n1000), .CI(n749), .CO(n744), .S(n745) );
  FA_X1 U637 ( .A(n946), .B(n982), .CI(n1019), .CO(n746), .S(n747) );
  HA_X1 U638 ( .A(n824), .B(n928), .CO(n748), .S(n749) );
  FA_X1 U639 ( .A(n760), .B(n755), .CI(n753), .CO(n750), .S(n751) );
  FA_X1 U640 ( .A(n762), .B(n764), .CI(n757), .CO(n752), .S(n753) );
  FA_X1 U641 ( .A(n947), .B(n1001), .CI(n983), .CO(n754), .S(n755) );
  FA_X1 U642 ( .A(n965), .B(n929), .CI(n1020), .CO(n756), .S(n757) );
  FA_X1 U643 ( .A(n763), .B(n768), .CI(n761), .CO(n758), .S(n759) );
  FA_X1 U644 ( .A(n765), .B(n1021), .CI(n770), .CO(n760), .S(n761) );
  FA_X1 U645 ( .A(n966), .B(n984), .CI(n1002), .CO(n762), .S(n763) );
  HA_X1 U646 ( .A(n825), .B(n948), .CO(n764), .S(n765) );
  FA_X1 U647 ( .A(n771), .B(n774), .CI(n769), .CO(n766), .S(n767) );
  FA_X1 U648 ( .A(n967), .B(n1003), .CI(n776), .CO(n768), .S(n769) );
  FA_X1 U649 ( .A(n985), .B(n949), .CI(n1022), .CO(n770), .S(n771) );
  FA_X1 U650 ( .A(n780), .B(n777), .CI(n775), .CO(n772), .S(n773) );
  FA_X1 U651 ( .A(n986), .B(n1023), .CI(n1004), .CO(n774), .S(n775) );
  HA_X1 U652 ( .A(n826), .B(n968), .CO(n776), .S(n777) );
  FA_X1 U653 ( .A(n784), .B(n987), .CI(n781), .CO(n778), .S(n779) );
  FA_X1 U654 ( .A(n1024), .B(n969), .CI(n1005), .CO(n780), .S(n781) );
  FA_X1 U655 ( .A(n1006), .B(n1025), .CI(n785), .CO(n782), .S(n783) );
  HA_X1 U656 ( .A(n827), .B(n988), .CO(n784), .S(n785) );
  FA_X1 U657 ( .A(n1007), .B(n989), .CI(n1026), .CO(n786), .S(n787) );
  HA_X1 U658 ( .A(n1008), .B(n1027), .CO(n788), .S(n789) );
  XNOR2_X1 U1180 ( .A(n314), .B(n1383), .ZN(product[20]) );
  AND2_X1 U1181 ( .A1(n428), .A2(n313), .ZN(n1383) );
  XNOR2_X1 U1182 ( .A(n268), .B(n1384), .ZN(product[26]) );
  AND2_X1 U1183 ( .A1(n264), .A2(n267), .ZN(n1384) );
  CLKBUF_X1 U1184 ( .A(n289), .Z(n1385) );
  NOR2_X1 U1185 ( .A1(n251), .A2(n275), .ZN(n1386) );
  NOR2_X2 U1186 ( .A1(n533), .A2(n546), .ZN(n275) );
  XNOR2_X1 U1187 ( .A(n1257), .B(n43), .ZN(n1387) );
  OAI22_X1 U1188 ( .A1(n1490), .A2(n1087), .B1(n46), .B2(n1086), .ZN(n1388) );
  CLKBUF_X3 U1189 ( .A(b[12]), .Z(n1247) );
  CLKBUF_X3 U1190 ( .A(b[16]), .Z(n1243) );
  BUF_X2 U1191 ( .A(n1246), .Z(n1389) );
  CLKBUF_X1 U1192 ( .A(n1282), .Z(n46) );
  BUF_X1 U1193 ( .A(b[4]), .Z(n1390) );
  CLKBUF_X1 U1194 ( .A(b[4]), .Z(n1255) );
  BUF_X1 U1195 ( .A(n1273), .Z(n41) );
  CLKBUF_X3 U1196 ( .A(b[15]), .Z(n1244) );
  CLKBUF_X3 U1197 ( .A(n1273), .Z(n1486) );
  CLKBUF_X3 U1198 ( .A(n1273), .Z(n42) );
  BUF_X4 U1199 ( .A(n1274), .Z(n36) );
  CLKBUF_X3 U1200 ( .A(n247), .Z(n1475) );
  CLKBUF_X3 U1201 ( .A(b[3]), .Z(n1256) );
  CLKBUF_X3 U1202 ( .A(b[2]), .Z(n1257) );
  CLKBUF_X3 U1203 ( .A(n291), .Z(n64) );
  XOR2_X1 U1204 ( .A(n866), .B(n938), .Z(n1391) );
  XOR2_X1 U1205 ( .A(n1388), .B(n1391), .Z(n643) );
  NAND2_X1 U1206 ( .A1(n884), .A2(n866), .ZN(n1392) );
  NAND2_X1 U1207 ( .A1(n884), .A2(n938), .ZN(n1393) );
  NAND2_X1 U1208 ( .A1(n866), .A2(n938), .ZN(n1394) );
  NAND3_X1 U1209 ( .A1(n1392), .A2(n1393), .A3(n1394), .ZN(n642) );
  XOR2_X1 U1210 ( .A(n637), .B(n635), .Z(n1395) );
  XOR2_X1 U1211 ( .A(n650), .B(n1395), .Z(n631) );
  NAND2_X1 U1212 ( .A1(n650), .A2(n637), .ZN(n1396) );
  NAND2_X1 U1213 ( .A1(n650), .A2(n635), .ZN(n1397) );
  NAND2_X1 U1214 ( .A1(n637), .A2(n635), .ZN(n1398) );
  NAND3_X1 U1215 ( .A1(n1396), .A2(n1397), .A3(n1398), .ZN(n630) );
  XOR2_X1 U1216 ( .A(n621), .B(n636), .Z(n1399) );
  XOR2_X1 U1217 ( .A(n619), .B(n1399), .Z(n615) );
  NAND2_X1 U1218 ( .A1(n619), .A2(n621), .ZN(n1400) );
  NAND2_X1 U1219 ( .A1(n619), .A2(n636), .ZN(n1401) );
  NAND2_X1 U1220 ( .A1(n621), .A2(n636), .ZN(n1402) );
  NAND3_X1 U1221 ( .A1(n1400), .A2(n1401), .A3(n1402), .ZN(n614) );
  NAND3_X2 U1222 ( .A1(n1449), .A2(n1450), .A3(n1451), .ZN(n636) );
  BUF_X1 U1223 ( .A(n22), .Z(n1481) );
  BUF_X2 U1224 ( .A(b[19]), .Z(n1240) );
  OR2_X1 U1225 ( .A1(n779), .A2(n782), .ZN(n1403) );
  OR2_X1 U1226 ( .A1(n787), .A2(n788), .ZN(n1404) );
  CLKBUF_X1 U1227 ( .A(n1446), .Z(n22) );
  BUF_X1 U1228 ( .A(n22), .Z(n1480) );
  XOR2_X1 U1229 ( .A(n664), .B(n651), .Z(n1405) );
  XOR2_X1 U1230 ( .A(n649), .B(n1405), .Z(n647) );
  NAND2_X1 U1231 ( .A1(n649), .A2(n664), .ZN(n1406) );
  NAND2_X1 U1232 ( .A1(n649), .A2(n651), .ZN(n1407) );
  NAND2_X1 U1233 ( .A1(n664), .A2(n651), .ZN(n1408) );
  NAND3_X1 U1234 ( .A1(n1406), .A2(n1407), .A3(n1408), .ZN(n646) );
  CLKBUF_X1 U1235 ( .A(n1180), .Z(n1409) );
  BUF_X1 U1236 ( .A(n1276), .Z(n24) );
  OR2_X1 U1237 ( .A1(n759), .A2(n766), .ZN(n1410) );
  XOR2_X1 U1238 ( .A(n648), .B(n633), .Z(n1411) );
  XOR2_X1 U1239 ( .A(n631), .B(n1411), .Z(n629) );
  NAND2_X1 U1240 ( .A1(n631), .A2(n648), .ZN(n1412) );
  NAND2_X1 U1241 ( .A1(n631), .A2(n633), .ZN(n1413) );
  NAND2_X1 U1242 ( .A1(n648), .A2(n633), .ZN(n1414) );
  NAND3_X1 U1243 ( .A1(n1412), .A2(n1413), .A3(n1414), .ZN(n628) );
  CLKBUF_X3 U1244 ( .A(b[1]), .Z(n1258) );
  CLKBUF_X1 U1245 ( .A(n1283), .Z(n1477) );
  CLKBUF_X3 U1246 ( .A(b[6]), .Z(n1253) );
  AOI21_X1 U1247 ( .B1(n1536), .B2(n336), .A(n1479), .ZN(n1415) );
  OR2_X2 U1248 ( .A1(n663), .A2(n678), .ZN(n1536) );
  BUF_X1 U1249 ( .A(n1279), .Z(n6) );
  BUF_X1 U1250 ( .A(n1278), .Z(n12) );
  BUF_X2 U1251 ( .A(b[14]), .Z(n1245) );
  OAI22_X1 U1252 ( .A1(n60), .A2(n1031), .B1(n58), .B2(n1030), .ZN(n448) );
  BUF_X2 U1253 ( .A(n61), .Z(n1550) );
  NOR2_X1 U1254 ( .A1(n577), .A2(n592), .ZN(n1416) );
  NOR2_X1 U1255 ( .A1(n577), .A2(n592), .ZN(n1532) );
  BUF_X2 U1256 ( .A(n1272), .Z(n1490) );
  OR2_X1 U1257 ( .A1(n473), .A2(n480), .ZN(n1417) );
  OR2_X1 U1258 ( .A1(n453), .A2(n456), .ZN(n1418) );
  OR2_X1 U1259 ( .A1(n467), .A2(n472), .ZN(n1419) );
  OR2_X1 U1260 ( .A1(n830), .A2(n448), .ZN(n1420) );
  OR2_X1 U1261 ( .A1(n452), .A2(n451), .ZN(n1421) );
  OR2_X1 U1262 ( .A1(n450), .A2(n449), .ZN(n1422) );
  OR2_X1 U1263 ( .A1(n751), .A2(n758), .ZN(n1423) );
  OR2_X1 U1264 ( .A1(n457), .A2(n460), .ZN(n1424) );
  OR2_X1 U1265 ( .A1(n767), .A2(n772), .ZN(n1425) );
  OR2_X1 U1266 ( .A1(n1029), .A2(n829), .ZN(n1426) );
  CLKBUF_X1 U1267 ( .A(n358), .Z(n1427) );
  CLKBUF_X1 U1268 ( .A(n282), .Z(n1428) );
  CLKBUF_X1 U1269 ( .A(n1501), .Z(n1429) );
  CLKBUF_X1 U1270 ( .A(n350), .Z(n1430) );
  CLKBUF_X3 U1271 ( .A(a[9]), .Z(n1488) );
  BUF_X1 U1272 ( .A(a[9]), .Z(n25) );
  CLKBUF_X1 U1273 ( .A(n64), .Z(n1431) );
  CLKBUF_X1 U1274 ( .A(n1099), .Z(n1432) );
  CLKBUF_X1 U1275 ( .A(n1282), .Z(n45) );
  CLKBUF_X1 U1276 ( .A(n1282), .Z(n1461) );
  CLKBUF_X3 U1277 ( .A(b[10]), .Z(n1249) );
  CLKBUF_X1 U1278 ( .A(b[17]), .Z(n1437) );
  BUF_X2 U1279 ( .A(n1276), .Z(n1433) );
  XNOR2_X1 U1280 ( .A(n43), .B(n1258), .ZN(n1434) );
  XNOR2_X1 U1281 ( .A(n19), .B(n1250), .ZN(n1435) );
  XNOR2_X1 U1282 ( .A(a[9]), .B(a[10]), .ZN(n1436) );
  CLKBUF_X1 U1283 ( .A(b[17]), .Z(n1438) );
  CLKBUF_X1 U1284 ( .A(b[17]), .Z(n1242) );
  BUF_X1 U1285 ( .A(n1279), .Z(n1439) );
  BUF_X1 U1286 ( .A(n1279), .Z(n1440) );
  NOR2_X1 U1287 ( .A1(n303), .A2(n1532), .ZN(n1441) );
  NOR2_X1 U1288 ( .A1(n509), .A2(n520), .ZN(n255) );
  BUF_X1 U1289 ( .A(n28), .Z(n1473) );
  BUF_X2 U1290 ( .A(b[13]), .Z(n1246) );
  BUF_X1 U1291 ( .A(n1436), .Z(n34) );
  CLKBUF_X2 U1292 ( .A(n1436), .Z(n33) );
  XNOR2_X1 U1293 ( .A(n613), .B(n1442), .ZN(n611) );
  XNOR2_X1 U1294 ( .A(n630), .B(n615), .ZN(n1442) );
  XNOR2_X1 U1295 ( .A(n25), .B(n1241), .ZN(n1443) );
  OR2_X2 U1296 ( .A1(n693), .A2(n706), .ZN(n1444) );
  CLKBUF_X1 U1297 ( .A(n1060), .Z(n1445) );
  XNOR2_X1 U1298 ( .A(a[6]), .B(a[5]), .ZN(n1446) );
  NOR2_X1 U1299 ( .A1(n707), .A2(n718), .ZN(n1447) );
  XOR2_X1 U1300 ( .A(n658), .B(n645), .Z(n1448) );
  XOR2_X1 U1301 ( .A(n660), .B(n1448), .Z(n637) );
  NAND2_X1 U1302 ( .A1(n660), .A2(n658), .ZN(n1449) );
  NAND2_X1 U1303 ( .A1(n660), .A2(n645), .ZN(n1450) );
  NAND2_X1 U1304 ( .A1(n658), .A2(n645), .ZN(n1451) );
  CLKBUF_X1 U1305 ( .A(n1241), .Z(n1452) );
  BUF_X2 U1306 ( .A(n1469), .Z(n1501) );
  BUF_X2 U1307 ( .A(n1277), .Z(n17) );
  XNOR2_X1 U1308 ( .A(n681), .B(n1453), .ZN(n679) );
  XNOR2_X1 U1309 ( .A(n694), .B(n683), .ZN(n1453) );
  NAND2_X1 U1310 ( .A1(n613), .A2(n630), .ZN(n1454) );
  NAND2_X1 U1311 ( .A1(n613), .A2(n615), .ZN(n1455) );
  NAND2_X1 U1312 ( .A1(n630), .A2(n615), .ZN(n1456) );
  NAND3_X1 U1313 ( .A1(n1454), .A2(n1455), .A3(n1456), .ZN(n610) );
  BUF_X2 U1314 ( .A(n10), .Z(n1457) );
  CLKBUF_X1 U1315 ( .A(n10), .Z(n1458) );
  CLKBUF_X3 U1316 ( .A(n1275), .Z(n1484) );
  CLKBUF_X3 U1317 ( .A(b[8]), .Z(n1251) );
  CLKBUF_X1 U1318 ( .A(n1251), .Z(n1459) );
  CLKBUF_X1 U1319 ( .A(n1531), .Z(n1470) );
  BUF_X1 U1320 ( .A(n1272), .Z(n47) );
  BUF_X2 U1321 ( .A(b[18]), .Z(n1241) );
  BUF_X2 U1322 ( .A(n1271), .Z(n1460) );
  CLKBUF_X1 U1323 ( .A(n1271), .Z(n53) );
  CLKBUF_X1 U1324 ( .A(n304), .Z(n1462) );
  XNOR2_X1 U1325 ( .A(n7), .B(n1245), .ZN(n1463) );
  INV_X1 U1326 ( .A(n1479), .ZN(n331) );
  CLKBUF_X1 U1327 ( .A(n1281), .Z(n52) );
  CLKBUF_X2 U1328 ( .A(n1281), .Z(n51) );
  CLKBUF_X1 U1329 ( .A(n1536), .Z(n1464) );
  CLKBUF_X3 U1330 ( .A(n1277), .Z(n1472) );
  CLKBUF_X1 U1331 ( .A(n303), .Z(n1465) );
  CLKBUF_X1 U1332 ( .A(n311), .Z(n1466) );
  CLKBUF_X1 U1333 ( .A(n1278), .Z(n1467) );
  BUF_X2 U1334 ( .A(n1278), .Z(n11) );
  CLKBUF_X1 U1335 ( .A(n1204), .Z(n1468) );
  AOI21_X1 U1336 ( .B1(n283), .B2(n1386), .A(n250), .ZN(n1469) );
  XNOR2_X1 U1337 ( .A(n1256), .B(n49), .ZN(n1471) );
  BUF_X2 U1338 ( .A(n28), .Z(n1474) );
  CLKBUF_X1 U1339 ( .A(n247), .Z(n66) );
  CLKBUF_X1 U1340 ( .A(n1283), .Z(n1476) );
  XNOR2_X1 U1341 ( .A(n25), .B(n1248), .ZN(n1478) );
  AND2_X1 U1342 ( .A1(n663), .A2(n678), .ZN(n1479) );
  CLKBUF_X1 U1343 ( .A(n7), .Z(n1482) );
  XNOR2_X1 U1344 ( .A(n49), .B(n1257), .ZN(n1483) );
  CLKBUF_X3 U1345 ( .A(n27), .Z(n1485) );
  BUF_X1 U1346 ( .A(n1285), .Z(n27) );
  BUF_X1 U1347 ( .A(a[9]), .Z(n1487) );
  CLKBUF_X1 U1348 ( .A(n19), .Z(n1489) );
  CLKBUF_X1 U1349 ( .A(n43), .Z(n1491) );
  XNOR2_X1 U1350 ( .A(n277), .B(n1492), .ZN(product[25]) );
  AND2_X1 U1351 ( .A1(n273), .A2(n276), .ZN(n1492) );
  CLKBUF_X1 U1352 ( .A(n37), .Z(n1493) );
  CLKBUF_X1 U1353 ( .A(a[5]), .Z(n1494) );
  OAI22_X1 U1354 ( .A1(n23), .A2(n1157), .B1(n1481), .B2(n1156), .ZN(n1495) );
  INV_X1 U1355 ( .A(n1428), .ZN(n280) );
  XNOR2_X1 U1356 ( .A(n579), .B(n1496), .ZN(n577) );
  XNOR2_X1 U1357 ( .A(n594), .B(n581), .ZN(n1496) );
  XOR2_X1 U1358 ( .A(n569), .B(n573), .Z(n1497) );
  XOR2_X1 U1359 ( .A(n1497), .B(n584), .Z(n565) );
  NAND2_X1 U1360 ( .A1(n584), .A2(n569), .ZN(n1498) );
  NAND2_X1 U1361 ( .A1(n584), .A2(n573), .ZN(n1499) );
  NAND2_X1 U1362 ( .A1(n569), .A2(n573), .ZN(n1500) );
  NAND3_X1 U1363 ( .A1(n1498), .A2(n1499), .A3(n1500), .ZN(n564) );
  NAND2_X1 U1364 ( .A1(n579), .A2(n594), .ZN(n1502) );
  NAND2_X1 U1365 ( .A1(n579), .A2(n581), .ZN(n1503) );
  NAND2_X1 U1366 ( .A1(n594), .A2(n581), .ZN(n1504) );
  NAND3_X1 U1367 ( .A1(n1502), .A2(n1503), .A3(n1504), .ZN(n576) );
  NOR2_X1 U1368 ( .A1(n561), .A2(n576), .ZN(n289) );
  CLKBUF_X1 U1369 ( .A(a[5]), .Z(n13) );
  CLKBUF_X1 U1370 ( .A(n31), .Z(n1505) );
  NOR2_X1 U1371 ( .A1(n593), .A2(n610), .ZN(n303) );
  XOR2_X1 U1372 ( .A(n845), .B(n971), .Z(n1506) );
  XOR2_X1 U1373 ( .A(n1506), .B(n990), .Z(n591) );
  NAND2_X1 U1374 ( .A1(n845), .A2(n971), .ZN(n1507) );
  NAND2_X1 U1375 ( .A1(n845), .A2(n990), .ZN(n1508) );
  NAND2_X1 U1376 ( .A1(n971), .A2(n990), .ZN(n1509) );
  NAND3_X1 U1377 ( .A1(n1507), .A2(n1508), .A3(n1509), .ZN(n590) );
  XOR2_X1 U1378 ( .A(n575), .B(n898), .Z(n1510) );
  XOR2_X1 U1379 ( .A(n1510), .B(n590), .Z(n569) );
  NAND2_X1 U1380 ( .A1(n575), .A2(n898), .ZN(n1511) );
  NAND2_X1 U1381 ( .A1(n575), .A2(n590), .ZN(n1512) );
  NAND2_X1 U1382 ( .A1(n898), .A2(n590), .ZN(n1513) );
  NAND3_X1 U1383 ( .A1(n1511), .A2(n1512), .A3(n1513), .ZN(n568) );
  BUF_X2 U1384 ( .A(n1280), .Z(n57) );
  CLKBUF_X1 U1385 ( .A(n1280), .Z(n58) );
  BUF_X2 U1386 ( .A(n1270), .Z(n60) );
  BUF_X2 U1387 ( .A(n291), .Z(n63) );
  XNOR2_X1 U1388 ( .A(n222), .B(n1514), .ZN(product[30]) );
  AND2_X1 U1389 ( .A1(n418), .A2(n221), .ZN(n1514) );
  XNOR2_X1 U1390 ( .A(n209), .B(n1515), .ZN(product[31]) );
  AND2_X1 U1391 ( .A1(n1417), .A2(n208), .ZN(n1515) );
  CLKBUF_X1 U1392 ( .A(n290), .Z(n1516) );
  OR2_X1 U1393 ( .A1(n266), .A2(n255), .ZN(n251) );
  NOR2_X1 U1394 ( .A1(n547), .A2(n560), .ZN(n1517) );
  NOR2_X1 U1395 ( .A1(n547), .A2(n560), .ZN(n284) );
  CLKBUF_X1 U1396 ( .A(n340), .Z(n1518) );
  CLKBUF_X1 U1397 ( .A(n49), .Z(n1519) );
  XNOR2_X1 U1398 ( .A(n55), .B(n1390), .ZN(n1520) );
  CLKBUF_X1 U1399 ( .A(n1488), .Z(n1521) );
  CLKBUF_X1 U1400 ( .A(n1257), .Z(n1522) );
  CLKBUF_X3 U1401 ( .A(n61), .Z(n1523) );
  XNOR2_X1 U1402 ( .A(n1528), .B(n1437), .ZN(n1524) );
  XNOR2_X1 U1403 ( .A(n55), .B(n1256), .ZN(n1525) );
  BUF_X4 U1404 ( .A(a[19]), .Z(n55) );
  CLKBUF_X1 U1405 ( .A(n1288), .Z(n9) );
  CLKBUF_X3 U1406 ( .A(n61), .Z(n1549) );
  OR2_X1 U1407 ( .A1(n1470), .A2(n317), .ZN(n1526) );
  CLKBUF_X1 U1408 ( .A(n1240), .Z(n1527) );
  BUF_X1 U1409 ( .A(n1285), .Z(n28) );
  CLKBUF_X3 U1410 ( .A(a[5]), .Z(n1528) );
  BUF_X2 U1411 ( .A(n1277), .Z(n18) );
  CLKBUF_X3 U1412 ( .A(b[7]), .Z(n1252) );
  NOR2_X1 U1413 ( .A1(n647), .A2(n662), .ZN(n1529) );
  OAI21_X1 U1414 ( .B1(n284), .B2(n290), .A(n285), .ZN(n1530) );
  OAI22_X1 U1415 ( .A1(n1460), .A2(n1471), .B1(n51), .B2(n1066), .ZN(n865) );
  BUF_X1 U1416 ( .A(b[0]), .Z(n61) );
  CLKBUF_X3 U1417 ( .A(b[11]), .Z(n1248) );
  NOR2_X1 U1418 ( .A1(n611), .A2(n628), .ZN(n1531) );
  NAND2_X1 U1419 ( .A1(n1263), .A2(n1283), .ZN(n1273) );
  BUF_X1 U1420 ( .A(n1103), .Z(n1533) );
  BUF_X2 U1421 ( .A(n1270), .Z(n59) );
  OR2_X1 U1422 ( .A1(n647), .A2(n662), .ZN(n1534) );
  CLKBUF_X1 U1423 ( .A(n1429), .Z(n1535) );
  NAND2_X1 U1424 ( .A1(n1262), .A2(n1282), .ZN(n1272) );
  NAND2_X1 U1425 ( .A1(n681), .A2(n694), .ZN(n1537) );
  NAND2_X1 U1426 ( .A1(n681), .A2(n683), .ZN(n1538) );
  NAND2_X1 U1427 ( .A1(n694), .A2(n683), .ZN(n1539) );
  NAND3_X1 U1428 ( .A1(n1537), .A2(n1538), .A3(n1539), .ZN(n678) );
  CLKBUF_X3 U1429 ( .A(b[5]), .Z(n1254) );
  CLKBUF_X1 U1430 ( .A(n320), .Z(n1540) );
  CLKBUF_X1 U1431 ( .A(n1256), .Z(n1541) );
  CLKBUF_X3 U1432 ( .A(b[9]), .Z(n1250) );
  NOR2_X1 U1433 ( .A1(n629), .A2(n646), .ZN(n317) );
  BUF_X2 U1434 ( .A(n1276), .Z(n23) );
  INV_X1 U1435 ( .A(n1530), .ZN(n281) );
  XNOR2_X1 U1436 ( .A(n257), .B(n1542), .ZN(product[27]) );
  AND2_X1 U1437 ( .A1(n253), .A2(n256), .ZN(n1542) );
  XNOR2_X1 U1438 ( .A(n298), .B(n1543), .ZN(product[22]) );
  AND2_X1 U1439 ( .A1(n426), .A2(n297), .ZN(n1543) );
  XNOR2_X1 U1440 ( .A(n286), .B(n1544), .ZN(product[24]) );
  AND2_X1 U1441 ( .A1(n424), .A2(n285), .ZN(n1544) );
  XNOR2_X1 U1442 ( .A(n305), .B(n1545), .ZN(product[21]) );
  AND2_X1 U1443 ( .A1(n302), .A2(n1462), .ZN(n1545) );
  AOI21_X1 U1444 ( .B1(n1536), .B2(n336), .A(n1479), .ZN(n327) );
  XNOR2_X1 U1445 ( .A(n231), .B(n1546), .ZN(product[29]) );
  AND2_X1 U1446 ( .A1(n227), .A2(n230), .ZN(n1546) );
  XNOR2_X1 U1447 ( .A(n244), .B(n1547), .ZN(product[28]) );
  AND2_X1 U1448 ( .A1(n240), .A2(n243), .ZN(n1547) );
  NOR2_X1 U1449 ( .A1(n707), .A2(n718), .ZN(n350) );
  NOR2_X1 U1450 ( .A1(n679), .A2(n692), .ZN(n337) );
  NAND2_X1 U1451 ( .A1(n629), .A2(n646), .ZN(n318) );
  NAND2_X1 U1452 ( .A1(n533), .A2(n546), .ZN(n276) );
  NAND2_X1 U1453 ( .A1(n593), .A2(n610), .ZN(n304) );
  NOR2_X1 U1454 ( .A1(n461), .A2(n466), .ZN(n179) );
  NOR2_X1 U1455 ( .A1(n489), .A2(n498), .ZN(n229) );
  NOR2_X1 U1456 ( .A1(n741), .A2(n750), .ZN(n364) );
  NOR2_X1 U1457 ( .A1(n499), .A2(n508), .ZN(n242) );
  NOR2_X1 U1458 ( .A1(n1028), .A2(n1009), .ZN(n406) );
  NOR2_X1 U1459 ( .A1(n773), .A2(n778), .ZN(n386) );
  NOR2_X1 U1460 ( .A1(n789), .A2(n828), .ZN(n402) );
  AND2_X1 U1461 ( .A1(n1426), .A2(n409), .ZN(product[1]) );
  BUF_X2 U1462 ( .A(n1446), .Z(n21) );
  BUF_X2 U1463 ( .A(n1287), .Z(n15) );
  BUF_X2 U1464 ( .A(n1287), .Z(n16) );
  BUF_X4 U1465 ( .A(a[1]), .Z(n1) );
  NAND2_X1 U1466 ( .A1(n1260), .A2(n1280), .ZN(n1270) );
  NAND2_X1 U1467 ( .A1(n1266), .A2(n1286), .ZN(n1276) );
  NAND2_X1 U1468 ( .A1(n1261), .A2(n1281), .ZN(n1271) );
  NAND2_X1 U1469 ( .A1(n1267), .A2(n1287), .ZN(n1277) );
  INV_X1 U1470 ( .A(a[0]), .ZN(n1289) );
  NOR2_X1 U1471 ( .A1(n280), .A2(n260), .ZN(n258) );
  NOR2_X1 U1472 ( .A1(n280), .A2(n275), .ZN(n269) );
  NAND2_X1 U1473 ( .A1(n214), .A2(n134), .ZN(n130) );
  INV_X1 U1474 ( .A(n186), .ZN(n184) );
  INV_X1 U1475 ( .A(n173), .ZN(n171) );
  INV_X1 U1476 ( .A(n1475), .ZN(n245) );
  INV_X1 U1477 ( .A(n1526), .ZN(n306) );
  NOR2_X1 U1478 ( .A1(n216), .A2(n175), .ZN(n173) );
  NOR2_X1 U1479 ( .A1(n216), .A2(n192), .ZN(n186) );
  OAI21_X1 U1480 ( .B1(n281), .B2(n260), .A(n261), .ZN(n259) );
  AOI21_X1 U1481 ( .B1(n274), .B2(n264), .A(n265), .ZN(n261) );
  INV_X1 U1482 ( .A(n187), .ZN(n185) );
  INV_X1 U1483 ( .A(n216), .ZN(n214) );
  NAND2_X1 U1484 ( .A1(n1536), .A2(n432), .ZN(n326) );
  OAI21_X1 U1485 ( .B1(n281), .B2(n275), .A(n276), .ZN(n270) );
  NAND2_X1 U1486 ( .A1(n273), .A2(n264), .ZN(n260) );
  INV_X1 U1487 ( .A(n1466), .ZN(n309) );
  NOR2_X1 U1488 ( .A1(n1526), .A2(n1465), .ZN(n299) );
  INV_X1 U1489 ( .A(n192), .ZN(n190) );
  NAND2_X1 U1490 ( .A1(n186), .A2(n149), .ZN(n145) );
  NAND2_X1 U1491 ( .A1(n214), .A2(n1417), .ZN(n201) );
  INV_X1 U1492 ( .A(n119), .ZN(n117) );
  INV_X1 U1493 ( .A(n1501), .ZN(n246) );
  NAND2_X1 U1494 ( .A1(n429), .A2(n318), .ZN(n86) );
  INV_X1 U1495 ( .A(n317), .ZN(n429) );
  XOR2_X1 U1496 ( .A(n339), .B(n89), .Z(product[16]) );
  NAND2_X1 U1497 ( .A1(n432), .A2(n338), .ZN(n89) );
  INV_X1 U1498 ( .A(n337), .ZN(n432) );
  OAI21_X1 U1499 ( .B1(n318), .B2(n1531), .A(n313), .ZN(n311) );
  NOR2_X1 U1500 ( .A1(n317), .A2(n1531), .ZN(n310) );
  AOI21_X1 U1501 ( .B1(n319), .B2(n429), .A(n316), .ZN(n314) );
  INV_X1 U1502 ( .A(n1470), .ZN(n428) );
  NOR2_X1 U1503 ( .A1(n303), .A2(n1532), .ZN(n294) );
  NAND2_X1 U1504 ( .A1(n348), .A2(n1444), .ZN(n341) );
  INV_X1 U1505 ( .A(n346), .ZN(n344) );
  NAND2_X1 U1506 ( .A1(n425), .A2(n1516), .ZN(n82) );
  INV_X1 U1507 ( .A(n1385), .ZN(n425) );
  INV_X1 U1508 ( .A(n1517), .ZN(n424) );
  AOI21_X1 U1509 ( .B1(n311), .B2(n1441), .A(n295), .ZN(n293) );
  NAND2_X1 U1510 ( .A1(n294), .A2(n310), .ZN(n292) );
  OAI21_X1 U1511 ( .B1(n217), .B2(n192), .A(n193), .ZN(n187) );
  NAND2_X1 U1512 ( .A1(n218), .A2(n240), .ZN(n216) );
  NOR2_X1 U1513 ( .A1(n216), .A2(n121), .ZN(n119) );
  INV_X1 U1514 ( .A(n1532), .ZN(n426) );
  XOR2_X1 U1515 ( .A(n347), .B(n90), .Z(product[15]) );
  NAND2_X1 U1516 ( .A1(n1444), .A2(n346), .ZN(n90) );
  AOI21_X1 U1517 ( .B1(n340), .B2(n321), .A(n322), .ZN(n320) );
  NOR2_X1 U1518 ( .A1(n1529), .A2(n326), .ZN(n321) );
  OAI21_X1 U1519 ( .B1(n327), .B2(n1529), .A(n324), .ZN(n322) );
  AOI21_X1 U1520 ( .B1(n283), .B2(n1386), .A(n250), .ZN(n248) );
  OAI21_X1 U1521 ( .B1(n251), .B2(n276), .A(n252), .ZN(n250) );
  AOI21_X1 U1522 ( .B1(n253), .B2(n265), .A(n254), .ZN(n252) );
  AOI21_X1 U1523 ( .B1(n215), .B2(n1417), .A(n206), .ZN(n202) );
  INV_X1 U1524 ( .A(n174), .ZN(n172) );
  XOR2_X1 U1525 ( .A(n352), .B(n91), .Z(product[14]) );
  NAND2_X1 U1526 ( .A1(n434), .A2(n351), .ZN(n91) );
  AOI21_X1 U1527 ( .B1(n357), .B2(n435), .A(n354), .ZN(n352) );
  INV_X1 U1528 ( .A(n1430), .ZN(n434) );
  INV_X1 U1529 ( .A(n255), .ZN(n253) );
  INV_X1 U1530 ( .A(n266), .ZN(n264) );
  XNOR2_X1 U1531 ( .A(n332), .B(n88), .ZN(product[17]) );
  NAND2_X1 U1532 ( .A1(n1464), .A2(n331), .ZN(n88) );
  OAI21_X1 U1533 ( .B1(n339), .B2(n337), .A(n338), .ZN(n332) );
  INV_X1 U1534 ( .A(n217), .ZN(n215) );
  NAND2_X1 U1535 ( .A1(n190), .A2(n177), .ZN(n175) );
  INV_X1 U1536 ( .A(n267), .ZN(n265) );
  OAI21_X1 U1537 ( .B1(n309), .B2(n1465), .A(n1462), .ZN(n300) );
  INV_X1 U1538 ( .A(n275), .ZN(n273) );
  INV_X1 U1539 ( .A(n338), .ZN(n336) );
  INV_X1 U1540 ( .A(n276), .ZN(n274) );
  NAND2_X1 U1541 ( .A1(n1417), .A2(n1419), .ZN(n192) );
  INV_X1 U1542 ( .A(n193), .ZN(n191) );
  INV_X1 U1543 ( .A(n367), .ZN(n366) );
  INV_X1 U1544 ( .A(n256), .ZN(n254) );
  NAND2_X1 U1545 ( .A1(n240), .A2(n227), .ZN(n225) );
  XNOR2_X1 U1546 ( .A(n325), .B(n87), .ZN(product[18]) );
  OAI21_X1 U1547 ( .B1(n339), .B2(n326), .A(n1415), .ZN(n325) );
  NAND2_X1 U1548 ( .A1(n1534), .A2(n324), .ZN(n87) );
  NAND2_X1 U1549 ( .A1(n173), .A2(n1424), .ZN(n160) );
  INV_X1 U1550 ( .A(n318), .ZN(n316) );
  INV_X1 U1551 ( .A(n1516), .ZN(n288) );
  XOR2_X1 U1552 ( .A(n198), .B(n73), .Z(product[32]) );
  NAND2_X1 U1553 ( .A1(n1419), .A2(n197), .ZN(n73) );
  AOI21_X1 U1554 ( .B1(n218), .B2(n241), .A(n219), .ZN(n217) );
  XNOR2_X1 U1555 ( .A(n357), .B(n92), .ZN(product[13]) );
  NAND2_X1 U1556 ( .A1(n435), .A2(n356), .ZN(n92) );
  INV_X1 U1557 ( .A(n355), .ZN(n435) );
  XNOR2_X1 U1558 ( .A(n363), .B(n93), .ZN(product[12]) );
  NAND2_X1 U1559 ( .A1(n436), .A2(n362), .ZN(n93) );
  OAI21_X1 U1560 ( .B1(n366), .B2(n364), .A(n365), .ZN(n363) );
  INV_X1 U1561 ( .A(n361), .ZN(n436) );
  XNOR2_X1 U1562 ( .A(n379), .B(n96), .ZN(product[9]) );
  NAND2_X1 U1563 ( .A1(n1410), .A2(n378), .ZN(n96) );
  XOR2_X1 U1564 ( .A(n181), .B(n72), .Z(product[33]) );
  NAND2_X1 U1565 ( .A1(n177), .A2(n180), .ZN(n72) );
  NOR2_X1 U1566 ( .A1(n350), .A2(n355), .ZN(n348) );
  AOI21_X1 U1567 ( .B1(n1419), .B2(n206), .A(n195), .ZN(n193) );
  INV_X1 U1568 ( .A(n197), .ZN(n195) );
  NAND2_X1 U1569 ( .A1(n561), .A2(n576), .ZN(n290) );
  NAND2_X1 U1570 ( .A1(n679), .A2(n692), .ZN(n338) );
  OAI21_X1 U1571 ( .B1(n217), .B2(n175), .A(n176), .ZN(n174) );
  AOI21_X1 U1572 ( .B1(n191), .B2(n177), .A(n178), .ZN(n176) );
  INV_X1 U1573 ( .A(n180), .ZN(n178) );
  AOI21_X1 U1574 ( .B1(n241), .B2(n227), .A(n228), .ZN(n226) );
  INV_X1 U1575 ( .A(n230), .ZN(n228) );
  AOI21_X1 U1576 ( .B1(n187), .B2(n149), .A(n150), .ZN(n146) );
  AOI21_X1 U1577 ( .B1(n174), .B2(n1424), .A(n165), .ZN(n161) );
  AOI21_X1 U1578 ( .B1(n215), .B2(n134), .A(n135), .ZN(n131) );
  INV_X1 U1579 ( .A(n120), .ZN(n118) );
  INV_X1 U1580 ( .A(n380), .ZN(n379) );
  NAND2_X1 U1581 ( .A1(n693), .A2(n706), .ZN(n346) );
  NAND2_X1 U1582 ( .A1(n647), .A2(n662), .ZN(n324) );
  NOR2_X1 U1583 ( .A1(n179), .A2(n151), .ZN(n149) );
  NAND2_X1 U1584 ( .A1(n611), .A2(n628), .ZN(n313) );
  INV_X1 U1585 ( .A(n179), .ZN(n177) );
  NAND2_X1 U1586 ( .A1(n1424), .A2(n1418), .ZN(n151) );
  NAND2_X1 U1587 ( .A1(n577), .A2(n592), .ZN(n297) );
  NAND2_X1 U1588 ( .A1(n547), .A2(n560), .ZN(n285) );
  NAND2_X1 U1589 ( .A1(n707), .A2(n718), .ZN(n351) );
  INV_X1 U1590 ( .A(n242), .ZN(n240) );
  OAI21_X1 U1591 ( .B1(n368), .B2(n380), .A(n369), .ZN(n367) );
  NAND2_X1 U1592 ( .A1(n1423), .A2(n1410), .ZN(n368) );
  AOI21_X1 U1593 ( .B1(n1423), .B2(n376), .A(n371), .ZN(n369) );
  INV_X1 U1594 ( .A(n243), .ZN(n241) );
  INV_X1 U1595 ( .A(n378), .ZN(n376) );
  INV_X1 U1596 ( .A(n208), .ZN(n206) );
  XOR2_X1 U1597 ( .A(n366), .B(n94), .Z(product[11]) );
  NAND2_X1 U1598 ( .A1(n437), .A2(n365), .ZN(n94) );
  INV_X1 U1599 ( .A(n364), .ZN(n437) );
  XOR2_X1 U1600 ( .A(n374), .B(n95), .Z(product[10]) );
  AOI21_X1 U1601 ( .B1(n379), .B2(n1410), .A(n376), .ZN(n374) );
  NAND2_X1 U1602 ( .A1(n1423), .A2(n373), .ZN(n95) );
  NAND2_X1 U1603 ( .A1(n119), .A2(n1420), .ZN(n108) );
  INV_X1 U1604 ( .A(n356), .ZN(n354) );
  INV_X1 U1605 ( .A(n373), .ZN(n371) );
  NAND2_X1 U1606 ( .A1(n1403), .A2(n392), .ZN(n99) );
  XOR2_X1 U1607 ( .A(n168), .B(n71), .Z(product[34]) );
  NAND2_X1 U1608 ( .A1(n1424), .A2(n167), .ZN(n71) );
  XOR2_X1 U1609 ( .A(n142), .B(n69), .Z(product[36]) );
  NAND2_X1 U1610 ( .A1(n1421), .A2(n141), .ZN(n69) );
  XOR2_X1 U1611 ( .A(n127), .B(n68), .Z(product[37]) );
  NAND2_X1 U1612 ( .A1(n1422), .A2(n126), .ZN(n68) );
  XOR2_X1 U1613 ( .A(n114), .B(n67), .Z(product[38]) );
  NAND2_X1 U1614 ( .A1(n1420), .A2(n113), .ZN(n67) );
  XOR2_X1 U1615 ( .A(n157), .B(n70), .Z(product[35]) );
  NAND2_X1 U1616 ( .A1(n1418), .A2(n156), .ZN(n70) );
  INV_X1 U1617 ( .A(n392), .ZN(n390) );
  NOR2_X1 U1618 ( .A1(n731), .A2(n740), .ZN(n361) );
  AOI21_X1 U1619 ( .B1(n385), .B2(n1425), .A(n382), .ZN(n380) );
  INV_X1 U1620 ( .A(n384), .ZN(n382) );
  NOR2_X1 U1621 ( .A1(n719), .A2(n730), .ZN(n355) );
  OAI21_X1 U1622 ( .B1(n217), .B2(n121), .A(n122), .ZN(n120) );
  AOI21_X1 U1623 ( .B1(n135), .B2(n1422), .A(n124), .ZN(n122) );
  INV_X1 U1624 ( .A(n126), .ZN(n124) );
  NAND2_X1 U1625 ( .A1(n461), .A2(n466), .ZN(n180) );
  OAI21_X1 U1626 ( .B1(n193), .B2(n136), .A(n137), .ZN(n135) );
  AOI21_X1 U1627 ( .B1(n150), .B2(n1421), .A(n139), .ZN(n137) );
  INV_X1 U1628 ( .A(n141), .ZN(n139) );
  NAND2_X1 U1629 ( .A1(n443), .A2(n395), .ZN(n100) );
  NAND2_X1 U1630 ( .A1(n489), .A2(n498), .ZN(n230) );
  NAND2_X1 U1631 ( .A1(n719), .A2(n730), .ZN(n356) );
  NAND2_X1 U1632 ( .A1(n741), .A2(n750), .ZN(n365) );
  AOI21_X1 U1633 ( .B1(n120), .B2(n1420), .A(n111), .ZN(n109) );
  INV_X1 U1634 ( .A(n113), .ZN(n111) );
  NAND2_X1 U1635 ( .A1(n499), .A2(n508), .ZN(n243) );
  NAND2_X1 U1636 ( .A1(n759), .A2(n766), .ZN(n378) );
  NAND2_X1 U1637 ( .A1(n751), .A2(n758), .ZN(n373) );
  NAND2_X1 U1638 ( .A1(n473), .A2(n480), .ZN(n208) );
  NAND2_X1 U1639 ( .A1(n467), .A2(n472), .ZN(n197) );
  NAND2_X1 U1640 ( .A1(n481), .A2(n488), .ZN(n221) );
  INV_X1 U1641 ( .A(n167), .ZN(n165) );
  NAND2_X1 U1642 ( .A1(n441), .A2(n387), .ZN(n98) );
  INV_X1 U1643 ( .A(n386), .ZN(n441) );
  NAND2_X1 U1644 ( .A1(n1425), .A2(n384), .ZN(n97) );
  OAI21_X1 U1645 ( .B1(n151), .B2(n180), .A(n152), .ZN(n150) );
  AOI21_X1 U1646 ( .B1(n165), .B2(n1418), .A(n154), .ZN(n152) );
  INV_X1 U1647 ( .A(n156), .ZN(n154) );
  XOR2_X1 U1648 ( .A(n102), .B(n404), .Z(product[3]) );
  NAND2_X1 U1649 ( .A1(n445), .A2(n403), .ZN(n102) );
  INV_X1 U1650 ( .A(n402), .ZN(n445) );
  XOR2_X1 U1651 ( .A(n103), .B(n409), .Z(product[2]) );
  NAND2_X1 U1652 ( .A1(n446), .A2(n407), .ZN(n103) );
  INV_X1 U1653 ( .A(n406), .ZN(n446) );
  XNOR2_X1 U1654 ( .A(n101), .B(n401), .ZN(product[4]) );
  NAND2_X1 U1655 ( .A1(n1404), .A2(n400), .ZN(n101) );
  OAI21_X1 U1656 ( .B1(n402), .B2(n404), .A(n403), .ZN(n401) );
  NAND2_X1 U1657 ( .A1(n830), .A2(n448), .ZN(n113) );
  INV_X1 U1658 ( .A(n448), .ZN(n449) );
  AOI21_X1 U1659 ( .B1(n1404), .B2(n401), .A(n398), .ZN(n396) );
  INV_X1 U1660 ( .A(n400), .ZN(n398) );
  NAND2_X1 U1661 ( .A1(n1028), .A2(n1009), .ZN(n407) );
  INV_X1 U1662 ( .A(n478), .ZN(n479) );
  OR2_X1 U1663 ( .A1(n937), .A2(n865), .ZN(n626) );
  XNOR2_X1 U1664 ( .A(n937), .B(n865), .ZN(n627) );
  INV_X1 U1665 ( .A(n1495), .ZN(n545) );
  NAND2_X1 U1666 ( .A1(n457), .A2(n460), .ZN(n167) );
  NAND2_X1 U1667 ( .A1(n452), .A2(n451), .ZN(n141) );
  NAND2_X1 U1668 ( .A1(n450), .A2(n449), .ZN(n126) );
  NAND2_X1 U1669 ( .A1(n767), .A2(n772), .ZN(n384) );
  NAND2_X1 U1670 ( .A1(n779), .A2(n782), .ZN(n392) );
  NAND2_X1 U1671 ( .A1(n453), .A2(n456), .ZN(n156) );
  NAND2_X1 U1672 ( .A1(n773), .A2(n778), .ZN(n387) );
  NAND2_X1 U1673 ( .A1(n783), .A2(n786), .ZN(n395) );
  INV_X1 U1674 ( .A(n405), .ZN(n404) );
  OAI21_X1 U1675 ( .B1(n406), .B2(n409), .A(n407), .ZN(n405) );
  OAI22_X1 U1676 ( .A1(n36), .A2(n1115), .B1(n34), .B2(n1114), .ZN(n496) );
  OAI22_X1 U1677 ( .A1(n1460), .A2(n1052), .B1(n52), .B2(n1051), .ZN(n454) );
  OAI22_X1 U1678 ( .A1(n1439), .A2(n1237), .B1(n1236), .B2(n3), .ZN(n1028) );
  OAI22_X1 U1679 ( .A1(n29), .A2(n1443), .B1(n1474), .B2(n1135), .ZN(n518) );
  OAI22_X1 U1680 ( .A1(n42), .A2(n1094), .B1(n1476), .B2(n1093), .ZN(n478) );
  OAI22_X1 U1681 ( .A1(n1490), .A2(n1073), .B1(n1461), .B2(n1072), .ZN(n464)
         );
  OAI22_X1 U1682 ( .A1(n29), .A2(n1478), .B1(n1474), .B2(n1142), .ZN(n937) );
  OAI22_X1 U1683 ( .A1(n24), .A2(n1157), .B1(n1481), .B2(n1156), .ZN(n544) );
  OAI22_X1 U1684 ( .A1(n18), .A2(n1178), .B1(n16), .B2(n1177), .ZN(n574) );
  OAI22_X1 U1685 ( .A1(n11), .A2(n1199), .B1(n1198), .B2(n1458), .ZN(n608) );
  OAI22_X1 U1686 ( .A1(n48), .A2(n1292), .B1(n1092), .B2(n45), .ZN(n822) );
  OAI22_X1 U1687 ( .A1(n48), .A2(n1091), .B1(n1461), .B2(n1434), .ZN(n888) );
  OR2_X1 U1688 ( .A1(n1523), .A2(n1292), .ZN(n1092) );
  OAI22_X1 U1689 ( .A1(n29), .A2(n1295), .B1(n1155), .B2(n1485), .ZN(n825) );
  OAI22_X1 U1690 ( .A1(n1484), .A2(n1154), .B1(n1485), .B2(n1153), .ZN(n948)
         );
  OR2_X1 U1691 ( .A1(n1549), .A2(n1295), .ZN(n1155) );
  AOI21_X1 U1692 ( .B1(n1486), .B2(n1476), .A(n1093), .ZN(n799) );
  OAI22_X1 U1693 ( .A1(n60), .A2(n1032), .B1(n58), .B2(n1031), .ZN(n831) );
  INV_X1 U1694 ( .A(n793), .ZN(n850) );
  AOI21_X1 U1695 ( .B1(n54), .B2(n52), .A(n1051), .ZN(n793) );
  OAI22_X1 U1696 ( .A1(n60), .A2(n1034), .B1(n58), .B2(n1033), .ZN(n833) );
  OAI22_X1 U1697 ( .A1(n1467), .A2(n1216), .B1(n9), .B2(n1215), .ZN(n1007) );
  AND2_X1 U1698 ( .A1(n1550), .A2(n812), .ZN(n989) );
  OAI22_X1 U1699 ( .A1(n1440), .A2(n1235), .B1(n1234), .B2(n3), .ZN(n1026) );
  OAI22_X1 U1700 ( .A1(n11), .A2(n1463), .B1(n1457), .B2(n1202), .ZN(n994) );
  OAI22_X1 U1701 ( .A1(n1484), .A2(n1146), .B1(n1485), .B2(n1145), .ZN(n940)
         );
  OAI22_X1 U1702 ( .A1(n1440), .A2(n1222), .B1(n1221), .B2(n4), .ZN(n1013) );
  OAI22_X1 U1703 ( .A1(n1484), .A2(n1140), .B1(n1485), .B2(n1139), .ZN(n934)
         );
  OAI22_X1 U1704 ( .A1(n1490), .A2(n1083), .B1(n1461), .B2(n1082), .ZN(n880)
         );
  OAI22_X1 U1705 ( .A1(n23), .A2(n1159), .B1(n1480), .B2(n1158), .ZN(n952) );
  OAI22_X1 U1706 ( .A1(n29), .A2(n1145), .B1(n1474), .B2(n1144), .ZN(n939) );
  OAI22_X1 U1707 ( .A1(n35), .A2(n1126), .B1(n33), .B2(n1125), .ZN(n921) );
  OAI22_X1 U1708 ( .A1(n18), .A2(n1183), .B1(n16), .B2(n1182), .ZN(n975) );
  OAI22_X1 U1709 ( .A1(n1484), .A2(n1152), .B1(n1485), .B2(n1151), .ZN(n946)
         );
  OAI22_X1 U1710 ( .A1(n1439), .A2(n1228), .B1(n1227), .B2(n4), .ZN(n1019) );
  OAI22_X1 U1711 ( .A1(n1472), .A2(n1190), .B1(n15), .B2(n1189), .ZN(n982) );
  OAI22_X1 U1712 ( .A1(n30), .A2(n1151), .B1(n1473), .B2(n1150), .ZN(n945) );
  AND2_X1 U1713 ( .A1(n1549), .A2(n800), .ZN(n909) );
  OAI22_X1 U1714 ( .A1(n1439), .A2(n1227), .B1(n1226), .B2(n4), .ZN(n1018) );
  OAI22_X1 U1715 ( .A1(n1484), .A2(n1148), .B1(n1473), .B2(n1147), .ZN(n942)
         );
  OAI22_X1 U1716 ( .A1(n1440), .A2(n1224), .B1(n1223), .B2(n4), .ZN(n1015) );
  OAI22_X1 U1717 ( .A1(n17), .A2(n1186), .B1(n16), .B2(n1185), .ZN(n978) );
  OAI22_X1 U1718 ( .A1(n36), .A2(n1132), .B1(n33), .B2(n1131), .ZN(n927) );
  OAI22_X1 U1719 ( .A1(n11), .A2(n1208), .B1(n9), .B2(n1207), .ZN(n999) );
  OAI22_X1 U1720 ( .A1(n1433), .A2(n1170), .B1(n21), .B2(n1169), .ZN(n963) );
  OAI22_X1 U1721 ( .A1(n29), .A2(n1153), .B1(n1485), .B2(n1152), .ZN(n947) );
  OAI22_X1 U1722 ( .A1(n1467), .A2(n1210), .B1(n9), .B2(n1209), .ZN(n1001) );
  OAI22_X1 U1723 ( .A1(n17), .A2(n1191), .B1(n15), .B2(n1190), .ZN(n983) );
  OAI22_X1 U1724 ( .A1(n42), .A2(n1096), .B1(n40), .B2(n1095), .ZN(n892) );
  OAI22_X1 U1725 ( .A1(n54), .A2(n1058), .B1(n52), .B2(n1057), .ZN(n856) );
  OAI22_X1 U1726 ( .A1(n60), .A2(n1039), .B1(n58), .B2(n1038), .ZN(n838) );
  AOI21_X1 U1727 ( .B1(n6), .B2(n4), .A(n1219), .ZN(n817) );
  AOI21_X1 U1728 ( .B1(n12), .B2(n1457), .A(n1198), .ZN(n814) );
  AOI21_X1 U1729 ( .B1(n36), .B2(n34), .A(n1114), .ZN(n802) );
  OAI22_X1 U1730 ( .A1(n1460), .A2(n1291), .B1(n1071), .B2(n52), .ZN(n821) );
  OAI22_X1 U1731 ( .A1(n1460), .A2(n1070), .B1(n51), .B2(n1069), .ZN(n868) );
  OR2_X1 U1732 ( .A1(n1550), .A2(n1291), .ZN(n1071) );
  NAND2_X1 U1733 ( .A1(n1029), .A2(n829), .ZN(n409) );
  OAI22_X1 U1734 ( .A1(n17), .A2(n1195), .B1(n15), .B2(n1194), .ZN(n987) );
  OAI22_X1 U1735 ( .A1(n11), .A2(n1215), .B1(n9), .B2(n1214), .ZN(n1006) );
  OAI22_X1 U1736 ( .A1(n1439), .A2(n1234), .B1(n1233), .B2(n3), .ZN(n1025) );
  OAI22_X1 U1737 ( .A1(n60), .A2(n1033), .B1(n58), .B2(n1032), .ZN(n832) );
  INV_X1 U1738 ( .A(n454), .ZN(n455) );
  NAND2_X1 U1739 ( .A1(n789), .A2(n828), .ZN(n403) );
  AND2_X1 U1740 ( .A1(n1549), .A2(n815), .ZN(n1009) );
  INV_X1 U1741 ( .A(n9), .ZN(n815) );
  INV_X1 U1742 ( .A(n805), .ZN(n930) );
  OAI22_X1 U1743 ( .A1(n59), .A2(n1040), .B1(n58), .B2(n1039), .ZN(n839) );
  AOI21_X1 U1744 ( .B1(n29), .B2(n1485), .A(n1135), .ZN(n805) );
  OAI22_X1 U1745 ( .A1(n35), .A2(n1119), .B1(n34), .B2(n1118), .ZN(n914) );
  OAI22_X1 U1746 ( .A1(n30), .A2(n1138), .B1(n1474), .B2(n1137), .ZN(n932) );
  OAI22_X1 U1747 ( .A1(n41), .A2(n1100), .B1(n1477), .B2(n1099), .ZN(n896) );
  OAI22_X1 U1748 ( .A1(n36), .A2(n1125), .B1(n33), .B2(n1124), .ZN(n920) );
  OAI22_X1 U1749 ( .A1(n11), .A2(n1201), .B1(n1457), .B2(n1200), .ZN(n992) );
  OAI22_X1 U1750 ( .A1(n17), .A2(n1182), .B1(n16), .B2(n1181), .ZN(n974) );
  OAI22_X1 U1751 ( .A1(n35), .A2(n1118), .B1(n34), .B2(n1117), .ZN(n913) );
  OAI22_X1 U1752 ( .A1(n30), .A2(n1137), .B1(n1473), .B2(n1136), .ZN(n931) );
  OAI22_X1 U1753 ( .A1(n53), .A2(n1061), .B1(n1060), .B2(n51), .ZN(n859) );
  OAI22_X1 U1754 ( .A1(n35), .A2(n1128), .B1(n33), .B2(n1127), .ZN(n923) );
  OAI22_X1 U1755 ( .A1(n1204), .A2(n12), .B1(n1203), .B2(n10), .ZN(n995) );
  OAI22_X1 U1756 ( .A1(n1090), .A2(n47), .B1(n45), .B2(n1089), .ZN(n887) );
  OAI22_X1 U1757 ( .A1(n1490), .A2(n1080), .B1(n46), .B2(n1079), .ZN(n877) );
  OAI22_X1 U1758 ( .A1(n42), .A2(n1432), .B1(n1476), .B2(n1098), .ZN(n895) );
  AND2_X1 U1759 ( .A1(n1523), .A2(n791), .ZN(n849) );
  OAI22_X1 U1760 ( .A1(n6), .A2(n1221), .B1(n1220), .B2(n4), .ZN(n1012) );
  OAI22_X1 U1761 ( .A1(n47), .A2(n1088), .B1(n1087), .B2(n45), .ZN(n885) );
  OAI22_X1 U1762 ( .A1(n29), .A2(n1141), .B1(n1140), .B2(n1485), .ZN(n935) );
  OAI22_X1 U1763 ( .A1(n1486), .A2(n1533), .B1(n1476), .B2(n1102), .ZN(n899)
         );
  OAI22_X1 U1764 ( .A1(n48), .A2(n1084), .B1(n46), .B2(n1083), .ZN(n881) );
  OAI22_X1 U1765 ( .A1(n48), .A2(n1076), .B1(n1461), .B2(n1075), .ZN(n873) );
  OAI22_X1 U1766 ( .A1(n1460), .A2(n1057), .B1(n52), .B2(n1056), .ZN(n855) );
  OAI22_X1 U1767 ( .A1(n1433), .A2(n1162), .B1(n1481), .B2(n1161), .ZN(n955)
         );
  OAI22_X1 U1768 ( .A1(n1472), .A2(n1181), .B1(n16), .B2(n1409), .ZN(n973) );
  OAI22_X1 U1769 ( .A1(n1433), .A2(n1165), .B1(n21), .B2(n1164), .ZN(n958) );
  OAI22_X1 U1770 ( .A1(n1472), .A2(n1184), .B1(n16), .B2(n1183), .ZN(n976) );
  OAI22_X1 U1771 ( .A1(n1490), .A2(n1077), .B1(n1461), .B2(n1076), .ZN(n874)
         );
  INV_X1 U1772 ( .A(n496), .ZN(n497) );
  AND2_X1 U1773 ( .A1(n1550), .A2(n794), .ZN(n869) );
  OAI22_X1 U1774 ( .A1(n1223), .A2(n6), .B1(n1222), .B2(n4), .ZN(n1014) );
  OAI22_X1 U1775 ( .A1(n41), .A2(n1109), .B1(n1108), .B2(n1477), .ZN(n905) );
  OAI22_X1 U1776 ( .A1(n29), .A2(n1139), .B1(n1485), .B2(n1138), .ZN(n933) );
  OAI22_X1 U1777 ( .A1(n1460), .A2(n1063), .B1(n51), .B2(n1062), .ZN(n861) );
  OAI22_X1 U1778 ( .A1(n23), .A2(n1158), .B1(n1481), .B2(n1157), .ZN(n951) );
  OAI22_X1 U1779 ( .A1(n1467), .A2(n1202), .B1(n1458), .B2(n1201), .ZN(n993)
         );
  OAI22_X1 U1780 ( .A1(n42), .A2(n1107), .B1(n40), .B2(n1106), .ZN(n903) );
  OAI22_X1 U1781 ( .A1(n1460), .A2(n1069), .B1(n51), .B2(n1483), .ZN(n867) );
  OAI22_X1 U1782 ( .A1(n36), .A2(n1116), .B1(n34), .B2(n1115), .ZN(n911) );
  OAI22_X1 U1783 ( .A1(n1490), .A2(n1078), .B1(n46), .B2(n1077), .ZN(n875) );
  OAI22_X1 U1784 ( .A1(n1460), .A2(n1059), .B1(n52), .B2(n1058), .ZN(n857) );
  INV_X1 U1785 ( .A(n1485), .ZN(n806) );
  INV_X1 U1786 ( .A(n45), .ZN(n797) );
  INV_X1 U1787 ( .A(n1477), .ZN(n800) );
  OAI22_X1 U1788 ( .A1(n1484), .A2(n1150), .B1(n1485), .B2(n1149), .ZN(n944)
         );
  OAI22_X1 U1789 ( .A1(n36), .A2(n1131), .B1(n33), .B2(n1130), .ZN(n926) );
  OAI22_X1 U1790 ( .A1(n1472), .A2(n1188), .B1(n15), .B2(n1187), .ZN(n980) );
  OAI22_X1 U1791 ( .A1(n1144), .A2(n30), .B1(n1143), .B2(n27), .ZN(n938) );
  OAI22_X1 U1792 ( .A1(n1490), .A2(n1087), .B1(n46), .B2(n1086), .ZN(n884) );
  OAI22_X1 U1793 ( .A1(n1483), .A2(n53), .B1(n1067), .B2(n51), .ZN(n866) );
  OAI22_X1 U1794 ( .A1(n36), .A2(n1117), .B1(n34), .B2(n1116), .ZN(n912) );
  OAI22_X1 U1795 ( .A1(n42), .A2(n1098), .B1(n1476), .B2(n1097), .ZN(n894) );
  OAI22_X1 U1796 ( .A1(n48), .A2(n1079), .B1(n1461), .B2(n1078), .ZN(n876) );
  OAI22_X1 U1797 ( .A1(n36), .A2(n1122), .B1(n34), .B2(n1121), .ZN(n917) );
  OAI22_X1 U1798 ( .A1(n18), .A2(n1180), .B1(n16), .B2(n1524), .ZN(n972) );
  OAI22_X1 U1799 ( .A1(n1047), .A2(n59), .B1(n57), .B2(n1525), .ZN(n846) );
  OAI22_X1 U1800 ( .A1(n1486), .A2(n1104), .B1(n1477), .B2(n1103), .ZN(n900)
         );
  OAI22_X1 U1801 ( .A1(n23), .A2(n1164), .B1(n21), .B2(n1163), .ZN(n957) );
  OAI22_X1 U1802 ( .A1(n1129), .A2(n35), .B1(n33), .B2(n1128), .ZN(n924) );
  OAI22_X1 U1803 ( .A1(n1486), .A2(n1110), .B1(n1476), .B2(n1109), .ZN(n906)
         );
  OAI22_X1 U1804 ( .A1(n24), .A2(n1167), .B1(n1166), .B2(n21), .ZN(n960) );
  OAI22_X1 U1805 ( .A1(n5), .A2(n1230), .B1(n1229), .B2(n3), .ZN(n1021) );
  OAI22_X1 U1806 ( .A1(n11), .A2(n1211), .B1(n9), .B2(n1210), .ZN(n1002) );
  OAI22_X1 U1807 ( .A1(n1433), .A2(n1173), .B1(n21), .B2(n1172), .ZN(n966) );
  OAI22_X1 U1808 ( .A1(n17), .A2(n1192), .B1(n15), .B2(n1191), .ZN(n984) );
  OAI22_X1 U1809 ( .A1(n1124), .A2(n35), .B1(n1123), .B2(n33), .ZN(n919) );
  INV_X1 U1810 ( .A(n817), .ZN(n1010) );
  OAI22_X1 U1811 ( .A1(n59), .A2(n1048), .B1(n1047), .B2(n57), .ZN(n847) );
  OAI22_X1 U1812 ( .A1(n59), .A2(n1044), .B1(n57), .B2(n1043), .ZN(n843) );
  INV_X1 U1813 ( .A(n811), .ZN(n970) );
  AOI21_X1 U1814 ( .B1(n18), .B2(n16), .A(n1177), .ZN(n811) );
  OAI22_X1 U1815 ( .A1(n23), .A2(n1168), .B1(n21), .B2(n1167), .ZN(n961) );
  OAI22_X1 U1816 ( .A1(n1472), .A2(n1187), .B1(n15), .B2(n1186), .ZN(n979) );
  INV_X1 U1817 ( .A(n802), .ZN(n910) );
  OAI22_X1 U1818 ( .A1(n60), .A2(n1038), .B1(n58), .B2(n1037), .ZN(n837) );
  OAI22_X1 U1819 ( .A1(n1486), .A2(n1095), .B1(n40), .B2(n1094), .ZN(n891) );
  OAI22_X1 U1820 ( .A1(n1467), .A2(n1212), .B1(n9), .B2(n1211), .ZN(n1003) );
  OAI22_X1 U1821 ( .A1(n1433), .A2(n1174), .B1(n21), .B2(n1173), .ZN(n967) );
  OAI22_X1 U1822 ( .A1(n30), .A2(n1147), .B1(n1474), .B2(n1146), .ZN(n941) );
  OAI22_X1 U1823 ( .A1(n23), .A2(n1435), .B1(n21), .B2(n1165), .ZN(n959) );
  OAI22_X1 U1824 ( .A1(n18), .A2(n1185), .B1(n16), .B2(n1184), .ZN(n977) );
  OAI22_X1 U1825 ( .A1(n11), .A2(n1213), .B1(n9), .B2(n1212), .ZN(n1004) );
  OAI22_X1 U1826 ( .A1(n1440), .A2(n1232), .B1(n1231), .B2(n3), .ZN(n1023) );
  OAI22_X1 U1827 ( .A1(n17), .A2(n1194), .B1(n15), .B2(n1193), .ZN(n986) );
  OAI22_X1 U1828 ( .A1(n11), .A2(n1214), .B1(n9), .B2(n1213), .ZN(n1005) );
  AND2_X1 U1829 ( .A1(n1549), .A2(n809), .ZN(n969) );
  OAI22_X1 U1830 ( .A1(n1439), .A2(n1233), .B1(n1232), .B2(n3), .ZN(n1024) );
  OAI22_X1 U1831 ( .A1(n48), .A2(n1074), .B1(n46), .B2(n1073), .ZN(n871) );
  OAI22_X1 U1832 ( .A1(n1460), .A2(n1062), .B1(n51), .B2(n1061), .ZN(n860) );
  OAI22_X1 U1833 ( .A1(n48), .A2(n1081), .B1(n45), .B2(n1080), .ZN(n878) );
  OAI22_X1 U1834 ( .A1(n59), .A2(n1043), .B1(n57), .B2(n1042), .ZN(n842) );
  OAI22_X1 U1835 ( .A1(n36), .A2(n1121), .B1(n34), .B2(n1120), .ZN(n916) );
  OAI22_X1 U1836 ( .A1(n1460), .A2(n1064), .B1(n51), .B2(n1063), .ZN(n862) );
  OAI22_X1 U1837 ( .A1(n59), .A2(n1520), .B1(n57), .B2(n1044), .ZN(n844) );
  AND2_X1 U1838 ( .A1(n1523), .A2(n803), .ZN(n929) );
  OAI22_X1 U1839 ( .A1(n1439), .A2(n1229), .B1(n1228), .B2(n3), .ZN(n1020) );
  OAI22_X1 U1840 ( .A1(n24), .A2(n1172), .B1(n21), .B2(n1171), .ZN(n965) );
  OAI22_X1 U1841 ( .A1(n5), .A2(n1220), .B1(n1219), .B2(n4), .ZN(n1011) );
  OAI22_X1 U1842 ( .A1(n42), .A2(n1106), .B1(n1477), .B2(n1105), .ZN(n902) );
  OAI22_X1 U1843 ( .A1(n24), .A2(n1163), .B1(n1480), .B2(n1162), .ZN(n956) );
  OAI22_X1 U1844 ( .A1(n36), .A2(n1120), .B1(n34), .B2(n1119), .ZN(n915) );
  OAI22_X1 U1845 ( .A1(n1486), .A2(n1101), .B1(n1476), .B2(n1100), .ZN(n897)
         );
  OAI22_X1 U1846 ( .A1(n1490), .A2(n1082), .B1(n46), .B2(n1081), .ZN(n879) );
  OAI22_X1 U1847 ( .A1(n1484), .A2(n1149), .B1(n1485), .B2(n1148), .ZN(n943)
         );
  OAI22_X1 U1848 ( .A1(n1467), .A2(n1206), .B1(n1457), .B2(n1205), .ZN(n997)
         );
  OAI22_X1 U1849 ( .A1(n42), .A2(n1111), .B1(n40), .B2(n1110), .ZN(n907) );
  OAI22_X1 U1850 ( .A1(n54), .A2(n1065), .B1(n51), .B2(n1064), .ZN(n863) );
  OAI22_X1 U1851 ( .A1(n1433), .A2(n1160), .B1(n1481), .B2(n1159), .ZN(n953)
         );
  OAI22_X1 U1852 ( .A1(n11), .A2(n1205), .B1(n1458), .B2(n1468), .ZN(n996) );
  OAI22_X1 U1853 ( .A1(n1467), .A2(n1207), .B1(n1458), .B2(n1206), .ZN(n998)
         );
  OAI22_X1 U1854 ( .A1(n5), .A2(n1226), .B1(n1225), .B2(n4), .ZN(n1017) );
  OAI22_X1 U1855 ( .A1(n23), .A2(n1169), .B1(n21), .B2(n1168), .ZN(n962) );
  OAI22_X1 U1856 ( .A1(n59), .A2(n1042), .B1(n57), .B2(n1041), .ZN(n841) );
  INV_X1 U1857 ( .A(n808), .ZN(n950) );
  AOI21_X1 U1858 ( .B1(n24), .B2(n1480), .A(n1156), .ZN(n808) );
  OAI22_X1 U1859 ( .A1(n1484), .A2(n1142), .B1(n1485), .B2(n1141), .ZN(n936)
         );
  OAI22_X1 U1860 ( .A1(n36), .A2(n1123), .B1(n34), .B2(n1122), .ZN(n918) );
  INV_X1 U1861 ( .A(n608), .ZN(n609) );
  OAI22_X1 U1862 ( .A1(n36), .A2(n1127), .B1(n33), .B2(n1126), .ZN(n922) );
  OAI22_X1 U1863 ( .A1(n1490), .A2(n1387), .B1(n1461), .B2(n1088), .ZN(n886)
         );
  OAI22_X1 U1864 ( .A1(n42), .A2(n1108), .B1(n40), .B2(n1107), .ZN(n904) );
  OAI22_X1 U1865 ( .A1(n1460), .A2(n1055), .B1(n52), .B2(n1054), .ZN(n853) );
  OAI22_X1 U1866 ( .A1(n60), .A2(n1036), .B1(n58), .B2(n1035), .ZN(n835) );
  INV_X1 U1867 ( .A(n799), .ZN(n890) );
  OAI22_X1 U1868 ( .A1(n48), .A2(n1085), .B1(n1461), .B2(n1084), .ZN(n882) );
  OAI22_X1 U1869 ( .A1(n54), .A2(n1066), .B1(n51), .B2(n1065), .ZN(n864) );
  OAI22_X1 U1870 ( .A1(n1433), .A2(n1161), .B1(n21), .B2(n1160), .ZN(n954) );
  OAI22_X1 U1871 ( .A1(n11), .A2(n1200), .B1(n1457), .B2(n1199), .ZN(n991) );
  OAI22_X1 U1872 ( .A1(n1490), .A2(n1086), .B1(n46), .B2(n1085), .ZN(n883) );
  OAI22_X1 U1873 ( .A1(n1486), .A2(n1105), .B1(n40), .B2(n1104), .ZN(n901) );
  OAI22_X1 U1874 ( .A1(n48), .A2(n1075), .B1(n1461), .B2(n1074), .ZN(n872) );
  OAI22_X1 U1875 ( .A1(n60), .A2(n1037), .B1(n58), .B2(n1036), .ZN(n836) );
  OAI22_X1 U1876 ( .A1(n1460), .A2(n1056), .B1(n52), .B2(n1055), .ZN(n854) );
  INV_X1 U1877 ( .A(n814), .ZN(n990) );
  OAI22_X1 U1878 ( .A1(n59), .A2(n1046), .B1(n57), .B2(n1520), .ZN(n845) );
  OAI22_X1 U1879 ( .A1(n17), .A2(n1179), .B1(n1178), .B2(n16), .ZN(n971) );
  OAI22_X1 U1880 ( .A1(n1486), .A2(n1102), .B1(n40), .B2(n1101), .ZN(n898) );
  INV_X1 U1881 ( .A(n574), .ZN(n575) );
  INV_X1 U1882 ( .A(n518), .ZN(n519) );
  OAI22_X1 U1883 ( .A1(n59), .A2(n1041), .B1(n57), .B2(n1040), .ZN(n840) );
  OAI22_X1 U1884 ( .A1(n54), .A2(n1445), .B1(n52), .B2(n1059), .ZN(n858) );
  OAI22_X1 U1885 ( .A1(n11), .A2(n1209), .B1(n9), .B2(n1208), .ZN(n1000) );
  OAI22_X1 U1886 ( .A1(n23), .A2(n1171), .B1(n21), .B2(n1170), .ZN(n964) );
  OAI22_X1 U1887 ( .A1(n1472), .A2(n1189), .B1(n15), .B2(n1188), .ZN(n981) );
  OAI22_X1 U1888 ( .A1(n1486), .A2(n1097), .B1(n40), .B2(n1096), .ZN(n893) );
  OAI22_X1 U1889 ( .A1(n35), .A2(n1130), .B1(n33), .B2(n1129), .ZN(n925) );
  AND2_X1 U1890 ( .A1(n1523), .A2(n797), .ZN(n889) );
  OAI22_X1 U1891 ( .A1(n1440), .A2(n1225), .B1(n1224), .B2(n4), .ZN(n1016) );
  AND2_X1 U1892 ( .A1(n1523), .A2(n806), .ZN(n949) );
  OAI22_X1 U1893 ( .A1(n5), .A2(n1231), .B1(n1230), .B2(n3), .ZN(n1022) );
  OAI22_X1 U1894 ( .A1(n1472), .A2(n1193), .B1(n15), .B2(n1192), .ZN(n985) );
  NAND2_X1 U1895 ( .A1(n787), .A2(n788), .ZN(n400) );
  OAI22_X1 U1896 ( .A1(n41), .A2(n1293), .B1(n1113), .B2(n1477), .ZN(n823) );
  OAI22_X1 U1897 ( .A1(n1486), .A2(n1112), .B1(n1477), .B2(n1111), .ZN(n908)
         );
  OR2_X1 U1898 ( .A1(n1523), .A2(n1293), .ZN(n1113) );
  INV_X1 U1899 ( .A(n790), .ZN(n830) );
  AOI21_X1 U1900 ( .B1(n60), .B2(n58), .A(n1030), .ZN(n790) );
  OAI22_X1 U1901 ( .A1(n54), .A2(n1054), .B1(n52), .B2(n1053), .ZN(n852) );
  OAI22_X1 U1902 ( .A1(n60), .A2(n1035), .B1(n58), .B2(n1034), .ZN(n834) );
  INV_X1 U1903 ( .A(n464), .ZN(n465) );
  OR2_X1 U1904 ( .A1(n1549), .A2(n1290), .ZN(n1050) );
  OR2_X1 U1905 ( .A1(n1550), .A2(n1296), .ZN(n1176) );
  OR2_X1 U1906 ( .A1(n1549), .A2(n1297), .ZN(n1197) );
  OR2_X1 U1907 ( .A1(n1549), .A2(n1294), .ZN(n1134) );
  OAI22_X1 U1908 ( .A1(n54), .A2(n1053), .B1(n52), .B2(n1052), .ZN(n851) );
  INV_X1 U1909 ( .A(n796), .ZN(n870) );
  AOI21_X1 U1910 ( .B1(n48), .B2(n46), .A(n1072), .ZN(n796) );
  INV_X1 U1911 ( .A(n57), .ZN(n791) );
  INV_X1 U1912 ( .A(n33), .ZN(n803) );
  INV_X1 U1913 ( .A(n51), .ZN(n794) );
  INV_X1 U1914 ( .A(n21), .ZN(n809) );
  INV_X1 U1915 ( .A(n15), .ZN(n812) );
  AND2_X1 U1916 ( .A1(n1523), .A2(n818), .ZN(product[0]) );
  INV_X1 U1917 ( .A(n3), .ZN(n818) );
  OAI22_X1 U1918 ( .A1(n12), .A2(n1217), .B1(n9), .B2(n1216), .ZN(n1008) );
  OAI22_X1 U1919 ( .A1(n5), .A2(n1236), .B1(n1235), .B2(n3), .ZN(n1027) );
  XNOR2_X1 U1920 ( .A(n7), .B(n1549), .ZN(n1217) );
  OAI22_X1 U1921 ( .A1(n11), .A2(n1298), .B1(n1218), .B2(n1457), .ZN(n828) );
  OR2_X1 U1922 ( .A1(n1550), .A2(n1298), .ZN(n1218) );
  INV_X1 U1923 ( .A(n1482), .ZN(n1298) );
  OAI22_X1 U1924 ( .A1(n1440), .A2(n1299), .B1(n1239), .B2(n4), .ZN(n829) );
  INV_X1 U1925 ( .A(n1), .ZN(n1299) );
  OAI22_X1 U1926 ( .A1(n5), .A2(n1238), .B1(n1237), .B2(n3), .ZN(n1029) );
  XNOR2_X1 U1927 ( .A(n1528), .B(n1438), .ZN(n1179) );
  XNOR2_X1 U1928 ( .A(n1528), .B(n1241), .ZN(n1178) );
  XNOR2_X1 U1929 ( .A(n7), .B(n1438), .ZN(n1200) );
  XNOR2_X1 U1930 ( .A(n13), .B(n1245), .ZN(n1182) );
  XNOR2_X1 U1931 ( .A(n13), .B(n1246), .ZN(n1183) );
  XNOR2_X1 U1932 ( .A(n7), .B(n1241), .ZN(n1199) );
  XNOR2_X1 U1933 ( .A(n13), .B(n1247), .ZN(n1184) );
  XNOR2_X1 U1934 ( .A(n7), .B(n1243), .ZN(n1201) );
  XNOR2_X1 U1935 ( .A(n1528), .B(n1243), .ZN(n1180) );
  XNOR2_X1 U1936 ( .A(n7), .B(n1246), .ZN(n1204) );
  XNOR2_X1 U1937 ( .A(n1494), .B(n1244), .ZN(n1181) );
  XNOR2_X1 U1938 ( .A(n7), .B(n1247), .ZN(n1205) );
  XNOR2_X1 U1939 ( .A(n7), .B(n1245), .ZN(n1203) );
  XNOR2_X1 U1940 ( .A(n1494), .B(n1248), .ZN(n1185) );
  XNOR2_X1 U1941 ( .A(n7), .B(n1244), .ZN(n1202) );
  XNOR2_X1 U1942 ( .A(n1528), .B(n1249), .ZN(n1186) );
  XNOR2_X1 U1943 ( .A(n1494), .B(n1251), .ZN(n1188) );
  XNOR2_X1 U1944 ( .A(n1250), .B(n1528), .ZN(n1187) );
  XNOR2_X1 U1945 ( .A(n1528), .B(n1252), .ZN(n1189) );
  XNOR2_X1 U1946 ( .A(n1250), .B(n7), .ZN(n1208) );
  XNOR2_X1 U1947 ( .A(n7), .B(n1248), .ZN(n1206) );
  XNOR2_X1 U1948 ( .A(n1482), .B(n1459), .ZN(n1209) );
  XNOR2_X1 U1949 ( .A(n7), .B(n1253), .ZN(n1211) );
  XNOR2_X1 U1950 ( .A(n7), .B(n1249), .ZN(n1207) );
  XNOR2_X1 U1951 ( .A(n1528), .B(n1254), .ZN(n1191) );
  XNOR2_X1 U1952 ( .A(n7), .B(n1252), .ZN(n1210) );
  XNOR2_X1 U1953 ( .A(n1528), .B(n1390), .ZN(n1192) );
  XNOR2_X1 U1954 ( .A(n1494), .B(n1522), .ZN(n1194) );
  XNOR2_X1 U1955 ( .A(n1528), .B(n1253), .ZN(n1190) );
  XNOR2_X1 U1956 ( .A(n1482), .B(n1254), .ZN(n1212) );
  XNOR2_X1 U1957 ( .A(n1528), .B(n1541), .ZN(n1193) );
  XNOR2_X1 U1958 ( .A(n1494), .B(n1258), .ZN(n1195) );
  XNOR2_X1 U1959 ( .A(n7), .B(n1256), .ZN(n1214) );
  XNOR2_X1 U1960 ( .A(n7), .B(n1390), .ZN(n1213) );
  XNOR2_X1 U1961 ( .A(n7), .B(n1257), .ZN(n1215) );
  XNOR2_X1 U1962 ( .A(n7), .B(n1258), .ZN(n1216) );
  XNOR2_X1 U1963 ( .A(n55), .B(n1258), .ZN(n1048) );
  XNOR2_X1 U1964 ( .A(n31), .B(n1248), .ZN(n1122) );
  XNOR2_X1 U1965 ( .A(n19), .B(n1241), .ZN(n1157) );
  XNOR2_X1 U1966 ( .A(n31), .B(n1247), .ZN(n1121) );
  XNOR2_X1 U1967 ( .A(n55), .B(n1257), .ZN(n1047) );
  XNOR2_X1 U1968 ( .A(n31), .B(n1249), .ZN(n1123) );
  XNOR2_X1 U1969 ( .A(n55), .B(n1256), .ZN(n1046) );
  XNOR2_X1 U1970 ( .A(n1250), .B(n31), .ZN(n1124) );
  XNOR2_X1 U1971 ( .A(n19), .B(n1247), .ZN(n1163) );
  XNOR2_X1 U1972 ( .A(n19), .B(n1244), .ZN(n1160) );
  XNOR2_X1 U1973 ( .A(n1489), .B(n1248), .ZN(n1164) );
  XNOR2_X1 U1974 ( .A(n55), .B(n1252), .ZN(n1042) );
  XNOR2_X1 U1975 ( .A(n55), .B(n1253), .ZN(n1043) );
  XNOR2_X1 U1976 ( .A(n55), .B(n1251), .ZN(n1041) );
  XNOR2_X1 U1977 ( .A(n31), .B(n1244), .ZN(n1118) );
  XNOR2_X1 U1978 ( .A(n55), .B(n1254), .ZN(n1044) );
  XNOR2_X1 U1979 ( .A(n31), .B(n1245), .ZN(n1119) );
  XNOR2_X1 U1980 ( .A(n1251), .B(n31), .ZN(n1125) );
  XNOR2_X1 U1981 ( .A(n19), .B(n1437), .ZN(n1158) );
  XNOR2_X1 U1982 ( .A(n31), .B(n1246), .ZN(n1120) );
  XNOR2_X1 U1983 ( .A(n31), .B(n1243), .ZN(n1117) );
  XNOR2_X1 U1984 ( .A(n19), .B(n1243), .ZN(n1159) );
  XNOR2_X1 U1985 ( .A(n31), .B(n1252), .ZN(n1126) );
  XNOR2_X1 U1986 ( .A(n19), .B(n1249), .ZN(n1165) );
  XNOR2_X1 U1987 ( .A(n19), .B(n1245), .ZN(n1161) );
  XNOR2_X1 U1988 ( .A(n31), .B(n1253), .ZN(n1127) );
  XNOR2_X1 U1989 ( .A(n19), .B(n1250), .ZN(n1166) );
  XNOR2_X1 U1990 ( .A(n19), .B(n1246), .ZN(n1162) );
  XNOR2_X1 U1991 ( .A(n31), .B(n1254), .ZN(n1128) );
  XNOR2_X1 U1992 ( .A(n1250), .B(n55), .ZN(n1040) );
  XNOR2_X1 U1993 ( .A(n19), .B(n1251), .ZN(n1167) );
  XNOR2_X1 U1994 ( .A(n19), .B(n1390), .ZN(n1171) );
  XNOR2_X1 U1995 ( .A(n31), .B(n1437), .ZN(n1116) );
  XNOR2_X1 U1996 ( .A(n31), .B(n1255), .ZN(n1129) );
  XNOR2_X1 U1997 ( .A(n19), .B(n1252), .ZN(n1168) );
  XNOR2_X1 U1998 ( .A(n19), .B(n1254), .ZN(n1170) );
  XNOR2_X1 U1999 ( .A(n19), .B(n1257), .ZN(n1173) );
  XNOR2_X1 U2000 ( .A(n31), .B(n1257), .ZN(n1131) );
  XNOR2_X1 U2001 ( .A(n31), .B(n1256), .ZN(n1130) );
  XNOR2_X1 U2002 ( .A(n19), .B(n1253), .ZN(n1169) );
  XNOR2_X1 U2003 ( .A(n19), .B(n1256), .ZN(n1172) );
  XNOR2_X1 U2004 ( .A(n31), .B(n1258), .ZN(n1132) );
  XNOR2_X1 U2005 ( .A(n19), .B(n1258), .ZN(n1174) );
  XNOR2_X1 U2006 ( .A(n1505), .B(n1241), .ZN(n1115) );
  XNOR2_X1 U2007 ( .A(n55), .B(n1249), .ZN(n1039) );
  XNOR2_X1 U2008 ( .A(n55), .B(n1248), .ZN(n1038) );
  XNOR2_X1 U2009 ( .A(n55), .B(n1247), .ZN(n1037) );
  XNOR2_X1 U2010 ( .A(n55), .B(n1244), .ZN(n1034) );
  XNOR2_X1 U2011 ( .A(n55), .B(n1389), .ZN(n1036) );
  XNOR2_X1 U2012 ( .A(n55), .B(n1245), .ZN(n1035) );
  XNOR2_X1 U2013 ( .A(n55), .B(n1243), .ZN(n1033) );
  XNOR2_X1 U2014 ( .A(n55), .B(n1437), .ZN(n1032) );
  XNOR2_X1 U2015 ( .A(n55), .B(n1452), .ZN(n1031) );
  XNOR2_X1 U2016 ( .A(n13), .B(n1240), .ZN(n1177) );
  XNOR2_X1 U2017 ( .A(n7), .B(n1240), .ZN(n1198) );
  XNOR2_X1 U2018 ( .A(n19), .B(n1240), .ZN(n1156) );
  XNOR2_X1 U2019 ( .A(n1505), .B(n1240), .ZN(n1114) );
  XNOR2_X1 U2020 ( .A(n55), .B(n1527), .ZN(n1030) );
  BUF_X1 U2021 ( .A(n1288), .Z(n10) );
  BUF_X2 U2022 ( .A(n1274), .Z(n35) );
  BUF_X1 U2023 ( .A(n1279), .Z(n5) );
  OAI22_X1 U2024 ( .A1(n36), .A2(n1133), .B1(n33), .B2(n1132), .ZN(n928) );
  OAI22_X1 U2025 ( .A1(n36), .A2(n1294), .B1(n1134), .B2(n34), .ZN(n824) );
  XNOR2_X1 U2026 ( .A(n31), .B(n1523), .ZN(n1133) );
  OAI22_X1 U2027 ( .A1(n1472), .A2(n1196), .B1(n15), .B2(n1195), .ZN(n988) );
  OAI22_X1 U2028 ( .A1(n17), .A2(n1297), .B1(n1197), .B2(n16), .ZN(n827) );
  XNOR2_X1 U2029 ( .A(n1528), .B(n1523), .ZN(n1196) );
  OAI22_X1 U2030 ( .A1(n59), .A2(n1049), .B1(n57), .B2(n1048), .ZN(n848) );
  OAI22_X1 U2031 ( .A1(n60), .A2(n1290), .B1(n1050), .B2(n57), .ZN(n820) );
  XNOR2_X1 U2032 ( .A(n55), .B(n1550), .ZN(n1049) );
  OAI22_X1 U2033 ( .A1(n23), .A2(n1175), .B1(n21), .B2(n1174), .ZN(n968) );
  OAI22_X1 U2034 ( .A1(n1433), .A2(n1296), .B1(n1176), .B2(n21), .ZN(n826) );
  XNOR2_X1 U2035 ( .A(n1489), .B(n1550), .ZN(n1175) );
  INV_X1 U2036 ( .A(n43), .ZN(n1292) );
  INV_X1 U2037 ( .A(n49), .ZN(n1291) );
  INV_X1 U2038 ( .A(n1487), .ZN(n1295) );
  BUF_X2 U2039 ( .A(n1272), .Z(n48) );
  INV_X1 U2040 ( .A(n1494), .ZN(n1297) );
  INV_X1 U2041 ( .A(n31), .ZN(n1294) );
  INV_X1 U2042 ( .A(n19), .ZN(n1296) );
  INV_X1 U2043 ( .A(n55), .ZN(n1290) );
  BUF_X1 U2044 ( .A(n1289), .Z(n3) );
  BUF_X1 U2045 ( .A(n1289), .Z(n4) );
  BUF_X1 U2046 ( .A(n1271), .Z(n54) );
  INV_X1 U2047 ( .A(n37), .ZN(n1293) );
  XNOR2_X1 U2048 ( .A(a[6]), .B(a[5]), .ZN(n1286) );
  XNOR2_X1 U2049 ( .A(a[4]), .B(a[3]), .ZN(n1287) );
  XNOR2_X1 U2050 ( .A(a[16]), .B(a[15]), .ZN(n1281) );
  XNOR2_X1 U2051 ( .A(a[1]), .B(a[2]), .ZN(n1288) );
  BUF_X4 U2052 ( .A(a[3]), .Z(n7) );
  BUF_X4 U2053 ( .A(a[11]), .Z(n31) );
  BUF_X4 U2054 ( .A(a[7]), .Z(n19) );
  BUF_X4 U2055 ( .A(a[13]), .Z(n37) );
  NAND2_X1 U2056 ( .A1(n1268), .A2(n1288), .ZN(n1278) );
  NAND2_X1 U2057 ( .A1(n1269), .A2(n1289), .ZN(n1279) );
  INV_X1 U2058 ( .A(n220), .ZN(n418) );
  OAI21_X1 U2059 ( .B1(n230), .B2(n220), .A(n221), .ZN(n219) );
  NOR2_X1 U2060 ( .A1(n481), .A2(n488), .ZN(n220) );
  BUF_X2 U2061 ( .A(n1275), .Z(n30) );
  BUF_X1 U2062 ( .A(n1275), .Z(n29) );
  NAND2_X1 U2063 ( .A1(n1285), .A2(n1265), .ZN(n1275) );
  CLKBUF_X1 U2064 ( .A(n1283), .Z(n40) );
  NOR2_X1 U2065 ( .A1(n192), .A2(n136), .ZN(n134) );
  NAND2_X1 U2066 ( .A1(n149), .A2(n1421), .ZN(n136) );
  NAND2_X1 U2067 ( .A1(n509), .A2(n520), .ZN(n256) );
  NOR2_X1 U2068 ( .A1(n229), .A2(n220), .ZN(n218) );
  INV_X1 U2069 ( .A(n229), .ZN(n227) );
  NOR2_X1 U2070 ( .A1(n783), .A2(n786), .ZN(n394) );
  OAI21_X1 U2071 ( .B1(n394), .B2(n396), .A(n395), .ZN(n393) );
  INV_X1 U2072 ( .A(n394), .ZN(n443) );
  XNOR2_X1 U2073 ( .A(n1487), .B(n1389), .ZN(n1141) );
  XNOR2_X1 U2074 ( .A(n1521), .B(n1550), .ZN(n1154) );
  XNOR2_X1 U2075 ( .A(n1488), .B(n1244), .ZN(n1139) );
  XNOR2_X1 U2076 ( .A(n1488), .B(n1245), .ZN(n1140) );
  XNOR2_X1 U2077 ( .A(n1487), .B(n1257), .ZN(n1152) );
  XNOR2_X1 U2078 ( .A(n1488), .B(n1256), .ZN(n1151) );
  XNOR2_X1 U2079 ( .A(n1390), .B(n1487), .ZN(n1150) );
  XNOR2_X1 U2080 ( .A(n1487), .B(n1247), .ZN(n1142) );
  XNOR2_X1 U2081 ( .A(n1487), .B(n1258), .ZN(n1153) );
  XNOR2_X1 U2082 ( .A(n1488), .B(n1254), .ZN(n1149) );
  XNOR2_X1 U2083 ( .A(n1250), .B(n1488), .ZN(n1145) );
  XNOR2_X1 U2084 ( .A(n25), .B(n1248), .ZN(n1143) );
  XNOR2_X1 U2085 ( .A(n1487), .B(n1243), .ZN(n1138) );
  XNOR2_X1 U2086 ( .A(n25), .B(n1249), .ZN(n1144) );
  XNOR2_X1 U2087 ( .A(n1488), .B(n1242), .ZN(n1137) );
  XNOR2_X1 U2088 ( .A(n1487), .B(n1253), .ZN(n1148) );
  XNOR2_X1 U2089 ( .A(n1488), .B(n1252), .ZN(n1147) );
  XNOR2_X1 U2090 ( .A(n1488), .B(n1251), .ZN(n1146) );
  XNOR2_X1 U2091 ( .A(n25), .B(n1241), .ZN(n1136) );
  XNOR2_X1 U2092 ( .A(n1488), .B(n1240), .ZN(n1135) );
  XNOR2_X1 U2093 ( .A(a[9]), .B(a[10]), .ZN(n1284) );
  NOR2_X1 U2094 ( .A1(n1475), .A2(n108), .ZN(n106) );
  NOR2_X1 U2095 ( .A1(n1475), .A2(n117), .ZN(n115) );
  NOR2_X1 U2096 ( .A1(n1475), .A2(n184), .ZN(n182) );
  NOR2_X1 U2097 ( .A1(n1475), .A2(n225), .ZN(n223) );
  NOR2_X1 U2098 ( .A1(n66), .A2(n242), .ZN(n232) );
  NOR2_X1 U2099 ( .A1(n1475), .A2(n171), .ZN(n169) );
  NOR2_X1 U2100 ( .A1(n1475), .A2(n160), .ZN(n158) );
  NOR2_X1 U2101 ( .A1(n1475), .A2(n201), .ZN(n199) );
  NOR2_X1 U2102 ( .A1(n1475), .A2(n145), .ZN(n143) );
  NOR2_X1 U2103 ( .A1(n1475), .A2(n130), .ZN(n128) );
  NOR2_X1 U2104 ( .A1(n66), .A2(n216), .ZN(n210) );
  OAI21_X1 U2105 ( .B1(n284), .B2(n290), .A(n285), .ZN(n283) );
  XNOR2_X1 U2106 ( .A(n1491), .B(n1245), .ZN(n1077) );
  XNOR2_X1 U2107 ( .A(n1491), .B(n1244), .ZN(n1076) );
  XNOR2_X1 U2108 ( .A(n43), .B(n1251), .ZN(n1083) );
  XNOR2_X1 U2109 ( .A(n43), .B(n1254), .ZN(n1086) );
  XNOR2_X1 U2110 ( .A(n43), .B(n1243), .ZN(n1075) );
  XNOR2_X1 U2111 ( .A(n1491), .B(n1437), .ZN(n1074) );
  XNOR2_X1 U2112 ( .A(n1250), .B(n43), .ZN(n1082) );
  XNOR2_X1 U2113 ( .A(n43), .B(n1249), .ZN(n1081) );
  XNOR2_X1 U2114 ( .A(n43), .B(n1248), .ZN(n1080) );
  XNOR2_X1 U2115 ( .A(n43), .B(n1550), .ZN(n1091) );
  XNOR2_X1 U2116 ( .A(n1491), .B(n1241), .ZN(n1073) );
  XNOR2_X1 U2117 ( .A(n1256), .B(n43), .ZN(n1088) );
  XNOR2_X1 U2118 ( .A(n43), .B(n1253), .ZN(n1085) );
  XNOR2_X1 U2119 ( .A(n43), .B(n1252), .ZN(n1084) );
  XNOR2_X1 U2120 ( .A(n43), .B(n1247), .ZN(n1079) );
  XNOR2_X1 U2121 ( .A(n1491), .B(n1527), .ZN(n1072) );
  XNOR2_X1 U2122 ( .A(n43), .B(n1255), .ZN(n1087) );
  XNOR2_X1 U2123 ( .A(n43), .B(n1246), .ZN(n1078) );
  XNOR2_X1 U2124 ( .A(n43), .B(n1258), .ZN(n1090) );
  XNOR2_X1 U2125 ( .A(n1257), .B(n43), .ZN(n1089) );
  BUF_X4 U2126 ( .A(a[15]), .Z(n43) );
  NOR2_X1 U2127 ( .A1(n521), .A2(n532), .ZN(n266) );
  NAND2_X1 U2128 ( .A1(n521), .A2(n532), .ZN(n267) );
  NOR2_X1 U2129 ( .A1(n251), .A2(n275), .ZN(n249) );
  NAND2_X1 U2130 ( .A1(n282), .A2(n249), .ZN(n247) );
  XNOR2_X1 U2131 ( .A(n1519), .B(n1243), .ZN(n1054) );
  XNOR2_X1 U2132 ( .A(n1519), .B(n1438), .ZN(n1053) );
  XNOR2_X1 U2133 ( .A(n49), .B(n1247), .ZN(n1058) );
  XNOR2_X1 U2134 ( .A(n49), .B(n1389), .ZN(n1057) );
  XNOR2_X1 U2135 ( .A(n49), .B(n1245), .ZN(n1056) );
  XNOR2_X1 U2136 ( .A(n1519), .B(n1244), .ZN(n1055) );
  XNOR2_X1 U2137 ( .A(n49), .B(n1248), .ZN(n1059) );
  XNOR2_X1 U2138 ( .A(n49), .B(n1549), .ZN(n1070) );
  XNOR2_X1 U2139 ( .A(n1256), .B(n49), .ZN(n1067) );
  XNOR2_X1 U2140 ( .A(n49), .B(n1253), .ZN(n1064) );
  XNOR2_X1 U2141 ( .A(n49), .B(n1258), .ZN(n1069) );
  XNOR2_X1 U2142 ( .A(n49), .B(n1252), .ZN(n1063) );
  XNOR2_X1 U2143 ( .A(n49), .B(n1251), .ZN(n1062) );
  XNOR2_X1 U2144 ( .A(n1250), .B(n49), .ZN(n1061) );
  XNOR2_X1 U2145 ( .A(n49), .B(n1249), .ZN(n1060) );
  XNOR2_X1 U2146 ( .A(n1519), .B(n1241), .ZN(n1052) );
  XNOR2_X1 U2147 ( .A(n1519), .B(n1527), .ZN(n1051) );
  XNOR2_X1 U2148 ( .A(n49), .B(n1390), .ZN(n1066) );
  XNOR2_X1 U2149 ( .A(n49), .B(n1254), .ZN(n1065) );
  XNOR2_X1 U2150 ( .A(a[18]), .B(a[17]), .ZN(n1280) );
  BUF_X4 U2151 ( .A(a[17]), .Z(n49) );
  AOI21_X1 U2152 ( .B1(n1431), .B2(n106), .A(n107), .ZN(n105) );
  AOI21_X1 U2153 ( .B1(n64), .B2(n115), .A(n116), .ZN(n114) );
  AOI21_X1 U2154 ( .B1(n64), .B2(n182), .A(n183), .ZN(n181) );
  AOI21_X1 U2155 ( .B1(n64), .B2(n169), .A(n170), .ZN(n168) );
  AOI21_X1 U2156 ( .B1(n64), .B2(n158), .A(n159), .ZN(n157) );
  AOI21_X1 U2157 ( .B1(n64), .B2(n143), .A(n144), .ZN(n142) );
  AOI21_X1 U2158 ( .B1(n64), .B2(n128), .A(n129), .ZN(n127) );
  AOI21_X1 U2159 ( .B1(n64), .B2(n199), .A(n200), .ZN(n198) );
  AOI21_X1 U2160 ( .B1(n63), .B2(n269), .A(n270), .ZN(n268) );
  AOI21_X1 U2161 ( .B1(n63), .B2(n232), .A(n233), .ZN(n231) );
  XNOR2_X1 U2162 ( .A(n64), .B(n82), .ZN(product[23]) );
  AOI21_X1 U2163 ( .B1(n64), .B2(n245), .A(n246), .ZN(n244) );
  AOI21_X1 U2164 ( .B1(n63), .B2(n258), .A(n259), .ZN(n257) );
  AOI21_X1 U2165 ( .B1(n64), .B2(n425), .A(n288), .ZN(n286) );
  AOI21_X1 U2166 ( .B1(n63), .B2(n223), .A(n224), .ZN(n222) );
  XNOR2_X1 U2167 ( .A(n1493), .B(n1243), .ZN(n1096) );
  XNOR2_X1 U2168 ( .A(n1493), .B(n1240), .ZN(n1093) );
  XNOR2_X1 U2169 ( .A(n1493), .B(n1438), .ZN(n1095) );
  XNOR2_X1 U2170 ( .A(n1493), .B(n1241), .ZN(n1094) );
  XNOR2_X1 U2171 ( .A(n37), .B(n1253), .ZN(n1106) );
  XNOR2_X1 U2172 ( .A(n37), .B(n1245), .ZN(n1098) );
  XNOR2_X1 U2173 ( .A(n37), .B(n1249), .ZN(n1102) );
  XNOR2_X1 U2174 ( .A(n37), .B(n1244), .ZN(n1097) );
  XNOR2_X1 U2175 ( .A(n37), .B(n1254), .ZN(n1107) );
  XNOR2_X1 U2176 ( .A(n37), .B(n1252), .ZN(n1105) );
  XNOR2_X1 U2177 ( .A(n37), .B(n1248), .ZN(n1101) );
  XNOR2_X1 U2178 ( .A(n37), .B(n1247), .ZN(n1100) );
  XNOR2_X1 U2179 ( .A(n37), .B(n1246), .ZN(n1099) );
  XNOR2_X1 U2180 ( .A(n37), .B(n1255), .ZN(n1108) );
  XNOR2_X1 U2181 ( .A(n37), .B(n1257), .ZN(n1110) );
  XNOR2_X1 U2182 ( .A(n1256), .B(n37), .ZN(n1109) );
  XNOR2_X1 U2183 ( .A(n37), .B(n1549), .ZN(n1112) );
  XNOR2_X1 U2184 ( .A(n37), .B(n1251), .ZN(n1104) );
  XNOR2_X1 U2185 ( .A(n1250), .B(n37), .ZN(n1103) );
  XNOR2_X1 U2186 ( .A(n37), .B(n1258), .ZN(n1111) );
  AOI21_X1 U2187 ( .B1(n63), .B2(n210), .A(n211), .ZN(n209) );
  XNOR2_X1 U2188 ( .A(n319), .B(n86), .ZN(product[19]) );
  AOI21_X1 U2189 ( .B1(n299), .B2(n319), .A(n300), .ZN(n298) );
  XNOR2_X1 U2190 ( .A(n385), .B(n97), .ZN(product[8]) );
  AOI21_X1 U2191 ( .B1(n319), .B2(n306), .A(n1466), .ZN(n305) );
  XNOR2_X1 U2192 ( .A(n1), .B(n1248), .ZN(n1227) );
  XNOR2_X1 U2193 ( .A(n1), .B(n1459), .ZN(n1230) );
  XNOR2_X1 U2194 ( .A(n1), .B(n1252), .ZN(n1231) );
  XNOR2_X1 U2195 ( .A(n1), .B(n1247), .ZN(n1226) );
  XNOR2_X1 U2196 ( .A(n1), .B(n1246), .ZN(n1225) );
  XNOR2_X1 U2197 ( .A(n1), .B(n1254), .ZN(n1233) );
  XNOR2_X1 U2198 ( .A(n1250), .B(n1), .ZN(n1229) );
  XNOR2_X1 U2199 ( .A(n1), .B(n1390), .ZN(n1234) );
  XNOR2_X1 U2200 ( .A(n1), .B(n1253), .ZN(n1232) );
  XNOR2_X1 U2201 ( .A(n1), .B(n1242), .ZN(n1221) );
  XNOR2_X1 U2202 ( .A(n1), .B(n1249), .ZN(n1228) );
  XNOR2_X1 U2203 ( .A(n1), .B(n1241), .ZN(n1220) );
  XNOR2_X1 U2204 ( .A(n1), .B(n1245), .ZN(n1224) );
  XNOR2_X1 U2205 ( .A(n1), .B(n1523), .ZN(n1238) );
  XNOR2_X1 U2206 ( .A(n1), .B(n1240), .ZN(n1219) );
  XNOR2_X1 U2207 ( .A(n1), .B(n1244), .ZN(n1223) );
  XNOR2_X1 U2208 ( .A(n1), .B(n1541), .ZN(n1235) );
  XNOR2_X1 U2209 ( .A(n1), .B(n1243), .ZN(n1222) );
  XNOR2_X1 U2210 ( .A(n1), .B(n1258), .ZN(n1237) );
  XNOR2_X1 U2211 ( .A(n1), .B(n1522), .ZN(n1236) );
  OAI21_X1 U2212 ( .B1(n1535), .B2(n108), .A(n109), .ZN(n107) );
  OAI21_X1 U2213 ( .B1(n1535), .B2(n117), .A(n118), .ZN(n116) );
  OAI21_X1 U2214 ( .B1(n248), .B2(n242), .A(n243), .ZN(n233) );
  OAI21_X1 U2215 ( .B1(n1501), .B2(n171), .A(n172), .ZN(n170) );
  OAI21_X1 U2216 ( .B1(n1501), .B2(n160), .A(n161), .ZN(n159) );
  OAI21_X1 U2217 ( .B1(n1429), .B2(n145), .A(n146), .ZN(n144) );
  OAI21_X1 U2218 ( .B1(n248), .B2(n225), .A(n226), .ZN(n224) );
  OAI21_X1 U2219 ( .B1(n1429), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U2220 ( .B1(n1501), .B2(n201), .A(n202), .ZN(n200) );
  OAI21_X1 U2221 ( .B1(n1501), .B2(n184), .A(n185), .ZN(n183) );
  OAI21_X1 U2222 ( .B1(n248), .B2(n216), .A(n217), .ZN(n211) );
  NAND2_X1 U2223 ( .A1(n1264), .A2(n1284), .ZN(n1274) );
  XOR2_X1 U2224 ( .A(a[10]), .B(a[11]), .Z(n1264) );
  XNOR2_X1 U2225 ( .A(a[11]), .B(a[12]), .ZN(n1283) );
  OAI21_X1 U2226 ( .B1(n1416), .B2(n304), .A(n297), .ZN(n295) );
  XOR2_X1 U2227 ( .A(a[18]), .B(a[19]), .Z(n1260) );
  INV_X1 U2228 ( .A(n1465), .ZN(n302) );
  OAI21_X1 U2229 ( .B1(n320), .B2(n292), .A(n293), .ZN(n291) );
  INV_X1 U2230 ( .A(n1540), .ZN(n319) );
  NOR2_X1 U2231 ( .A1(n361), .A2(n364), .ZN(n359) );
  OAI21_X1 U2232 ( .B1(n361), .B2(n365), .A(n362), .ZN(n360) );
  NAND2_X1 U2233 ( .A1(n731), .A2(n740), .ZN(n362) );
  INV_X1 U2234 ( .A(n1518), .ZN(n339) );
  XNOR2_X1 U2235 ( .A(a[8]), .B(a[7]), .ZN(n1285) );
  XOR2_X1 U2236 ( .A(a[6]), .B(a[7]), .Z(n1266) );
  XOR2_X1 U2237 ( .A(a[14]), .B(a[15]), .Z(n1262) );
  XNOR2_X1 U2238 ( .A(a[13]), .B(a[14]), .ZN(n1282) );
  XOR2_X1 U2239 ( .A(a[12]), .B(a[13]), .Z(n1263) );
  NAND2_X1 U2240 ( .A1(n134), .A2(n1422), .ZN(n121) );
  XOR2_X1 U2241 ( .A(a[2]), .B(a[3]), .Z(n1268) );
  OAI21_X1 U2242 ( .B1(n341), .B2(n358), .A(n342), .ZN(n340) );
  XOR2_X1 U2243 ( .A(a[9]), .B(a[8]), .Z(n1265) );
  NOR2_X1 U2244 ( .A1(n289), .A2(n1517), .ZN(n282) );
  XOR2_X1 U2245 ( .A(n388), .B(n98), .Z(product[7]) );
  OAI21_X1 U2246 ( .B1(n388), .B2(n386), .A(n387), .ZN(n385) );
  XOR2_X1 U2247 ( .A(a[4]), .B(a[5]), .Z(n1267) );
  AOI21_X1 U2248 ( .B1(n357), .B2(n348), .A(n349), .ZN(n347) );
  AOI21_X1 U2249 ( .B1(n349), .B2(n1444), .A(n344), .ZN(n342) );
  OAI21_X1 U2250 ( .B1(n1447), .B2(n356), .A(n351), .ZN(n349) );
  XOR2_X1 U2251 ( .A(a[16]), .B(a[17]), .Z(n1261) );
  XNOR2_X1 U2252 ( .A(n99), .B(n393), .ZN(product[6]) );
  INV_X1 U2253 ( .A(n1427), .ZN(n357) );
  AOI21_X1 U2254 ( .B1(n1403), .B2(n393), .A(n390), .ZN(n388) );
  XOR2_X1 U2255 ( .A(a[0]), .B(a[1]), .Z(n1269) );
  XOR2_X1 U2256 ( .A(n100), .B(n396), .Z(product[5]) );
  AOI21_X1 U2257 ( .B1(n367), .B2(n359), .A(n360), .ZN(n358) );
  AOI21_X1 U2258 ( .B1(n63), .B2(n1428), .A(n1530), .ZN(n277) );
  OR2_X1 U2259 ( .A1(n1550), .A2(n1299), .ZN(n1239) );
endmodule


module datapath_DW_mult_tc_14 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n15, n16, n17, n18,
         n21, n22, n23, n24, n25, n27, n29, n30, n31, n33, n34, n35, n36, n37,
         n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n51, n52, n53, n54,
         n55, n57, n58, n59, n60, n61, n63, n64, n65, n67, n68, n69, n70, n71,
         n72, n73, n82, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n105, n106, n107, n108, n109,
         n111, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n124, n126, n127, n128, n129, n130, n131, n134, n135, n136, n137,
         n139, n141, n142, n143, n144, n145, n146, n149, n150, n151, n152,
         n154, n156, n157, n158, n159, n160, n161, n165, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n190, n191, n192, n193,
         n195, n197, n198, n199, n200, n201, n202, n206, n208, n209, n210,
         n211, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n255, n256, n257, n258, n259, n260, n261, n264, n266, n267,
         n268, n269, n270, n273, n274, n275, n276, n277, n279, n280, n281,
         n282, n283, n284, n285, n286, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n303, n304, n305,
         n306, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n332, n333,
         n334, n336, n338, n339, n340, n341, n342, n344, n346, n347, n348,
         n349, n350, n351, n352, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n371, n373,
         n374, n376, n378, n379, n380, n382, n384, n385, n386, n387, n388,
         n390, n392, n393, n394, n395, n396, n398, n400, n401, n402, n403,
         n404, n405, n406, n407, n409, n418, n421, n424, n425, n428, n430,
         n434, n435, n436, n437, n441, n443, n445, n446, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n793,
         n794, n796, n797, n799, n800, n802, n803, n805, n806, n808, n809,
         n811, n812, n814, n815, n817, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1494, n1495;
  assign product[39] = n105;

  FA_X1 U488 ( .A(n831), .B(n454), .CI(n850), .CO(n450), .S(n451) );
  FA_X1 U489 ( .A(n455), .B(n832), .CI(n458), .CO(n452), .S(n453) );
  FA_X1 U491 ( .A(n462), .B(n833), .CI(n459), .CO(n456), .S(n457) );
  FA_X1 U492 ( .A(n851), .B(n464), .CI(n870), .CO(n458), .S(n459) );
  FA_X1 U493 ( .A(n463), .B(n470), .CI(n468), .CO(n460), .S(n461) );
  FA_X1 U494 ( .A(n834), .B(n852), .CI(n465), .CO(n462), .S(n463) );
  FA_X1 U496 ( .A(n474), .B(n471), .CI(n469), .CO(n466), .S(n467) );
  FA_X1 U497 ( .A(n478), .B(n871), .CI(n476), .CO(n468), .S(n469) );
  FA_X1 U498 ( .A(n853), .B(n835), .CI(n890), .CO(n470), .S(n471) );
  FA_X1 U499 ( .A(n475), .B(n477), .CI(n482), .CO(n472), .S(n473) );
  FA_X1 U500 ( .A(n486), .B(n479), .CI(n484), .CO(n474), .S(n475) );
  FA_X1 U501 ( .A(n836), .B(n854), .CI(n872), .CO(n476), .S(n477) );
  FA_X1 U503 ( .A(n490), .B(n492), .CI(n483), .CO(n480), .S(n481) );
  FA_X1 U504 ( .A(n485), .B(n494), .CI(n487), .CO(n482), .S(n483) );
  FA_X1 U505 ( .A(n855), .B(n496), .CI(n873), .CO(n484), .S(n485) );
  FA_X1 U506 ( .A(n891), .B(n837), .CI(n910), .CO(n486), .S(n487) );
  FA_X1 U507 ( .A(n500), .B(n493), .CI(n491), .CO(n488), .S(n489) );
  FA_X1 U508 ( .A(n495), .B(n504), .CI(n502), .CO(n490), .S(n491) );
  FA_X1 U509 ( .A(n497), .B(n874), .CI(n506), .CO(n492), .S(n493) );
  FA_X1 U510 ( .A(n892), .B(n856), .CI(n838), .CO(n494), .S(n495) );
  FA_X1 U512 ( .A(n510), .B(n503), .CI(n501), .CO(n498), .S(n499) );
  FA_X1 U513 ( .A(n507), .B(n505), .CI(n512), .CO(n500), .S(n501) );
  FA_X1 U514 ( .A(n516), .B(n893), .CI(n514), .CO(n502), .S(n503) );
  FA_X1 U515 ( .A(n857), .B(n911), .CI(n875), .CO(n504), .S(n505) );
  FA_X1 U516 ( .A(n518), .B(n839), .CI(n930), .CO(n506), .S(n507) );
  FA_X1 U517 ( .A(n522), .B(n513), .CI(n511), .CO(n508), .S(n509) );
  FA_X1 U518 ( .A(n526), .B(n515), .CI(n524), .CO(n510), .S(n511) );
  FA_X1 U519 ( .A(n528), .B(n530), .CI(n517), .CO(n512), .S(n513) );
  FA_X1 U520 ( .A(n840), .B(n858), .CI(n519), .CO(n514), .S(n515) );
  FA_X1 U521 ( .A(n912), .B(n876), .CI(n894), .CO(n516), .S(n517) );
  FA_X1 U523 ( .A(n525), .B(n534), .CI(n523), .CO(n520), .S(n521) );
  FA_X1 U524 ( .A(n527), .B(n538), .CI(n536), .CO(n522), .S(n523) );
  FA_X1 U525 ( .A(n529), .B(n540), .CI(n531), .CO(n524), .S(n525) );
  FA_X1 U526 ( .A(n877), .B(n895), .CI(n542), .CO(n526), .S(n527) );
  FA_X1 U527 ( .A(n859), .B(n913), .CI(n931), .CO(n528), .S(n529) );
  FA_X1 U528 ( .A(n544), .B(n841), .CI(n950), .CO(n530), .S(n531) );
  FA_X1 U529 ( .A(n548), .B(n537), .CI(n535), .CO(n532), .S(n533) );
  FA_X1 U530 ( .A(n539), .B(n552), .CI(n550), .CO(n534), .S(n535) );
  FA_X1 U531 ( .A(n541), .B(n554), .CI(n543), .CO(n536), .S(n537) );
  FA_X1 U532 ( .A(n558), .B(n545), .CI(n556), .CO(n538), .S(n539) );
  FA_X1 U533 ( .A(n896), .B(n932), .CI(n914), .CO(n540), .S(n541) );
  FA_X1 U534 ( .A(n842), .B(n878), .CI(n860), .CO(n542), .S(n543) );
  FA_X1 U536 ( .A(n562), .B(n551), .CI(n549), .CO(n546), .S(n547) );
  FA_X1 U537 ( .A(n553), .B(n566), .CI(n564), .CO(n548), .S(n549) );
  FA_X1 U538 ( .A(n559), .B(n557), .CI(n568), .CO(n550), .S(n551) );
  FA_X1 U539 ( .A(n570), .B(n572), .CI(n555), .CO(n552), .S(n553) );
  FA_X1 U540 ( .A(n879), .B(n915), .CI(n897), .CO(n554), .S(n555) );
  FA_X1 U541 ( .A(n861), .B(n951), .CI(n933), .CO(n556), .S(n557) );
  FA_X1 U542 ( .A(n574), .B(n843), .CI(n970), .CO(n558), .S(n559) );
  FA_X1 U543 ( .A(n578), .B(n565), .CI(n563), .CO(n560), .S(n561) );
  FA_X1 U544 ( .A(n567), .B(n582), .CI(n580), .CO(n562), .S(n563) );
  FA_X1 U546 ( .A(n586), .B(n588), .CI(n571), .CO(n566), .S(n567) );
  FA_X1 U548 ( .A(n844), .B(n916), .CI(n862), .CO(n570), .S(n571) );
  FA_X1 U549 ( .A(n952), .B(n880), .CI(n934), .CO(n572), .S(n573) );
  FA_X1 U552 ( .A(n583), .B(n598), .CI(n596), .CO(n578), .S(n579) );
  FA_X1 U553 ( .A(n600), .B(n591), .CI(n585), .CO(n580), .S(n581) );
  FA_X1 U554 ( .A(n587), .B(n602), .CI(n589), .CO(n582), .S(n583) );
  FA_X1 U555 ( .A(n606), .B(n917), .CI(n604), .CO(n584), .S(n585) );
  FA_X1 U556 ( .A(n881), .B(n935), .CI(n899), .CO(n586), .S(n587) );
  FA_X1 U557 ( .A(n608), .B(n953), .CI(n863), .CO(n588), .S(n589) );
  FA_X1 U558 ( .A(n845), .B(n971), .CI(n990), .CO(n590), .S(n591) );
  FA_X1 U559 ( .A(n612), .B(n597), .CI(n595), .CO(n592), .S(n593) );
  FA_X1 U560 ( .A(n599), .B(n616), .CI(n614), .CO(n594), .S(n595) );
  FA_X1 U561 ( .A(n618), .B(n603), .CI(n601), .CO(n596), .S(n597) );
  FA_X1 U562 ( .A(n605), .B(n607), .CI(n620), .CO(n598), .S(n599) );
  FA_X1 U563 ( .A(n624), .B(n626), .CI(n622), .CO(n600), .S(n601) );
  FA_X1 U564 ( .A(n918), .B(n936), .CI(n609), .CO(n602), .S(n603) );
  FA_X1 U565 ( .A(n954), .B(n864), .CI(n882), .CO(n604), .S(n605) );
  FA_X1 U569 ( .A(n617), .B(n634), .CI(n632), .CO(n612), .S(n613) );
  FA_X1 U570 ( .A(n636), .B(n621), .CI(n619), .CO(n614), .S(n615) );
  FA_X1 U571 ( .A(n623), .B(n638), .CI(n625), .CO(n616), .S(n617) );
  FA_X1 U572 ( .A(n642), .B(n627), .CI(n640), .CO(n618), .S(n619) );
  FA_X1 U573 ( .A(n955), .B(n973), .CI(n644), .CO(n620), .S(n621) );
  FA_X1 U574 ( .A(n991), .B(n901), .CI(n883), .CO(n622), .S(n623) );
  FA_X1 U575 ( .A(n847), .B(n919), .CI(n1010), .CO(n624), .S(n625) );
  FA_X1 U578 ( .A(n648), .B(n633), .CI(n631), .CO(n628), .S(n629) );
  FA_X1 U579 ( .A(n650), .B(n637), .CI(n635), .CO(n630), .S(n631) );
  FA_X1 U580 ( .A(n654), .B(n643), .CI(n652), .CO(n632), .S(n633) );
  FA_X1 U581 ( .A(n639), .B(n656), .CI(n641), .CO(n634), .S(n635) );
  FA_X1 U582 ( .A(n660), .B(n645), .CI(n658), .CO(n636), .S(n637) );
  FA_X1 U583 ( .A(n920), .B(n992), .CI(n974), .CO(n638), .S(n639) );
  FA_X1 U584 ( .A(n1011), .B(n956), .CI(n902), .CO(n640), .S(n641) );
  HA_X1 U586 ( .A(n820), .B(n848), .CO(n644), .S(n645) );
  FA_X1 U587 ( .A(n664), .B(n651), .CI(n649), .CO(n646), .S(n647) );
  FA_X1 U588 ( .A(n653), .B(n655), .CI(n666), .CO(n648), .S(n649) );
  FA_X1 U589 ( .A(n670), .B(n659), .CI(n668), .CO(n650), .S(n651) );
  FA_X1 U590 ( .A(n661), .B(n672), .CI(n657), .CO(n652), .S(n653) );
  FA_X1 U591 ( .A(n676), .B(n957), .CI(n674), .CO(n654), .S(n655) );
  FA_X1 U592 ( .A(n921), .B(n975), .CI(n939), .CO(n656), .S(n657) );
  FA_X1 U593 ( .A(n867), .B(n993), .CI(n903), .CO(n658), .S(n659) );
  FA_X1 U594 ( .A(n885), .B(n849), .CI(n1012), .CO(n660), .S(n661) );
  FA_X1 U595 ( .A(n667), .B(n680), .CI(n665), .CO(n662), .S(n663) );
  FA_X1 U596 ( .A(n669), .B(n671), .CI(n682), .CO(n664), .S(n665) );
  FA_X1 U597 ( .A(n675), .B(n673), .CI(n684), .CO(n666), .S(n667) );
  FA_X1 U598 ( .A(n690), .B(n686), .CI(n688), .CO(n668), .S(n669) );
  FA_X1 U599 ( .A(n958), .B(n976), .CI(n677), .CO(n670), .S(n671) );
  FA_X1 U600 ( .A(n886), .B(n904), .CI(n922), .CO(n672), .S(n673) );
  FA_X1 U601 ( .A(n1013), .B(n940), .CI(n994), .CO(n674), .S(n675) );
  HA_X1 U602 ( .A(n821), .B(n868), .CO(n676), .S(n677) );
  FA_X1 U603 ( .A(n694), .B(n683), .CI(n681), .CO(n678), .S(n679) );
  FA_X1 U604 ( .A(n685), .B(n698), .CI(n696), .CO(n680), .S(n681) );
  FA_X1 U605 ( .A(n689), .B(n691), .CI(n687), .CO(n682), .S(n683) );
  FA_X1 U606 ( .A(n702), .B(n1401), .CI(n700), .CO(n684), .S(n685) );
  FA_X1 U607 ( .A(n959), .B(n977), .CI(n941), .CO(n686), .S(n687) );
  FA_X1 U608 ( .A(n887), .B(n995), .CI(n923), .CO(n688), .S(n689) );
  FA_X1 U609 ( .A(n869), .B(n905), .CI(n1014), .CO(n690), .S(n691) );
  FA_X1 U610 ( .A(n697), .B(n708), .CI(n695), .CO(n692), .S(n693) );
  FA_X1 U611 ( .A(n710), .B(n703), .CI(n699), .CO(n694), .S(n695) );
  FA_X1 U612 ( .A(n701), .B(n714), .CI(n712), .CO(n696), .S(n697) );
  FA_X1 U613 ( .A(n705), .B(n996), .CI(n716), .CO(n698), .S(n699) );
  FA_X1 U614 ( .A(n1015), .B(n978), .CI(n942), .CO(n700), .S(n701) );
  FA_X1 U615 ( .A(n924), .B(n906), .CI(n960), .CO(n702), .S(n703) );
  FA_X1 U617 ( .A(n711), .B(n720), .CI(n709), .CO(n706), .S(n707) );
  FA_X1 U618 ( .A(n713), .B(n715), .CI(n722), .CO(n708), .S(n709) );
  FA_X1 U619 ( .A(n724), .B(n726), .CI(n717), .CO(n710), .S(n711) );
  FA_X1 U620 ( .A(n961), .B(n979), .CI(n728), .CO(n712), .S(n713) );
  FA_X1 U621 ( .A(n907), .B(n997), .CI(n943), .CO(n714), .S(n715) );
  FA_X1 U622 ( .A(n925), .B(n889), .CI(n1016), .CO(n716), .S(n717) );
  FA_X1 U623 ( .A(n732), .B(n723), .CI(n721), .CO(n718), .S(n719) );
  FA_X1 U624 ( .A(n727), .B(n725), .CI(n734), .CO(n720), .S(n721) );
  FA_X1 U625 ( .A(n738), .B(n729), .CI(n736), .CO(n722), .S(n723) );
  FA_X1 U626 ( .A(n926), .B(n980), .CI(n944), .CO(n724), .S(n725) );
  FA_X1 U627 ( .A(n1017), .B(n962), .CI(n998), .CO(n726), .S(n727) );
  HA_X1 U628 ( .A(n908), .B(n823), .CO(n728), .S(n729) );
  FA_X1 U629 ( .A(n735), .B(n742), .CI(n733), .CO(n730), .S(n731) );
  FA_X1 U630 ( .A(n737), .B(n739), .CI(n744), .CO(n732), .S(n733) );
  FA_X1 U631 ( .A(n748), .B(n981), .CI(n746), .CO(n734), .S(n735) );
  FA_X1 U632 ( .A(n927), .B(n999), .CI(n963), .CO(n736), .S(n737) );
  FA_X1 U633 ( .A(n945), .B(n909), .CI(n1018), .CO(n738), .S(n739) );
  FA_X1 U634 ( .A(n752), .B(n745), .CI(n743), .CO(n740), .S(n741) );
  FA_X1 U635 ( .A(n754), .B(n756), .CI(n747), .CO(n742), .S(n743) );
  FA_X1 U636 ( .A(n964), .B(n1000), .CI(n749), .CO(n744), .S(n745) );
  FA_X1 U637 ( .A(n946), .B(n982), .CI(n1019), .CO(n746), .S(n747) );
  HA_X1 U638 ( .A(n824), .B(n928), .CO(n748), .S(n749) );
  FA_X1 U639 ( .A(n760), .B(n755), .CI(n753), .CO(n750), .S(n751) );
  FA_X1 U640 ( .A(n762), .B(n764), .CI(n757), .CO(n752), .S(n753) );
  FA_X1 U641 ( .A(n947), .B(n1001), .CI(n983), .CO(n754), .S(n755) );
  FA_X1 U642 ( .A(n965), .B(n929), .CI(n1020), .CO(n756), .S(n757) );
  FA_X1 U643 ( .A(n763), .B(n768), .CI(n761), .CO(n758), .S(n759) );
  FA_X1 U644 ( .A(n765), .B(n1021), .CI(n770), .CO(n760), .S(n761) );
  FA_X1 U645 ( .A(n966), .B(n984), .CI(n1002), .CO(n762), .S(n763) );
  HA_X1 U646 ( .A(n825), .B(n948), .CO(n764), .S(n765) );
  FA_X1 U647 ( .A(n771), .B(n774), .CI(n769), .CO(n766), .S(n767) );
  FA_X1 U648 ( .A(n967), .B(n1003), .CI(n776), .CO(n768), .S(n769) );
  FA_X1 U649 ( .A(n985), .B(n949), .CI(n1022), .CO(n770), .S(n771) );
  FA_X1 U650 ( .A(n780), .B(n777), .CI(n775), .CO(n772), .S(n773) );
  FA_X1 U651 ( .A(n986), .B(n1023), .CI(n1004), .CO(n774), .S(n775) );
  HA_X1 U652 ( .A(n826), .B(n968), .CO(n776), .S(n777) );
  FA_X1 U653 ( .A(n784), .B(n987), .CI(n781), .CO(n778), .S(n779) );
  FA_X1 U654 ( .A(n1024), .B(n969), .CI(n1005), .CO(n780), .S(n781) );
  FA_X1 U655 ( .A(n1006), .B(n1025), .CI(n785), .CO(n782), .S(n783) );
  HA_X1 U656 ( .A(n827), .B(n988), .CO(n784), .S(n785) );
  FA_X1 U657 ( .A(n1026), .B(n989), .CI(n1007), .CO(n786), .S(n787) );
  HA_X1 U658 ( .A(n1008), .B(n1027), .CO(n788), .S(n789) );
  BUF_X1 U1180 ( .A(b[3]), .Z(n1488) );
  CLKBUF_X3 U1181 ( .A(b[18]), .Z(n1241) );
  CLKBUF_X3 U1182 ( .A(b[11]), .Z(n1248) );
  CLKBUF_X2 U1183 ( .A(b[7]), .Z(n1252) );
  CLKBUF_X3 U1184 ( .A(b[16]), .Z(n1243) );
  CLKBUF_X1 U1185 ( .A(b[2]), .Z(n1257) );
  CLKBUF_X3 U1186 ( .A(b[13]), .Z(n1246) );
  CLKBUF_X1 U1187 ( .A(b[9]), .Z(n1489) );
  CLKBUF_X3 U1188 ( .A(b[15]), .Z(n1244) );
  CLKBUF_X3 U1189 ( .A(b[14]), .Z(n1245) );
  CLKBUF_X3 U1190 ( .A(b[6]), .Z(n1253) );
  CLKBUF_X3 U1191 ( .A(b[17]), .Z(n1242) );
  CLKBUF_X1 U1192 ( .A(b[2]), .Z(n1486) );
  AND2_X1 U1193 ( .A1(n521), .A2(n532), .ZN(n1383) );
  BUF_X1 U1194 ( .A(n248), .Z(n1448) );
  INV_X1 U1195 ( .A(n1383), .ZN(n267) );
  BUF_X1 U1196 ( .A(n1484), .Z(n1458) );
  BUF_X2 U1197 ( .A(a[7]), .Z(n1471) );
  NAND2_X2 U1198 ( .A1(n282), .A2(n249), .ZN(n247) );
  BUF_X2 U1199 ( .A(n1275), .Z(n30) );
  CLKBUF_X3 U1200 ( .A(n1277), .Z(n17) );
  OR2_X2 U1201 ( .A1(n663), .A2(n678), .ZN(n1482) );
  CLKBUF_X3 U1202 ( .A(b[4]), .Z(n1255) );
  BUF_X1 U1203 ( .A(n1279), .Z(n6) );
  BUF_X1 U1204 ( .A(n1272), .Z(n47) );
  BUF_X2 U1205 ( .A(n1281), .Z(n51) );
  BUF_X2 U1206 ( .A(n1468), .Z(n1415) );
  BUF_X2 U1207 ( .A(n1468), .Z(n1414) );
  BUF_X2 U1208 ( .A(a[5]), .Z(n1467) );
  BUF_X2 U1209 ( .A(n1273), .Z(n42) );
  CLKBUF_X3 U1210 ( .A(n1273), .Z(n41) );
  XOR2_X1 U1211 ( .A(n866), .B(n938), .Z(n1384) );
  XOR2_X1 U1212 ( .A(n884), .B(n1384), .Z(n643) );
  NAND2_X1 U1213 ( .A1(n884), .A2(n866), .ZN(n1385) );
  NAND2_X1 U1214 ( .A1(n884), .A2(n938), .ZN(n1386) );
  NAND2_X1 U1215 ( .A1(n866), .A2(n938), .ZN(n1387) );
  NAND3_X1 U1216 ( .A1(n1385), .A2(n1386), .A3(n1387), .ZN(n642) );
  INV_X1 U1217 ( .A(n1422), .ZN(n256) );
  OR2_X1 U1218 ( .A1(n473), .A2(n480), .ZN(n1388) );
  OR2_X1 U1219 ( .A1(n759), .A2(n766), .ZN(n1389) );
  OR2_X1 U1220 ( .A1(n453), .A2(n456), .ZN(n1390) );
  OR2_X1 U1221 ( .A1(n467), .A2(n472), .ZN(n1391) );
  OR2_X1 U1222 ( .A1(n830), .A2(n448), .ZN(n1392) );
  OR2_X1 U1223 ( .A1(n452), .A2(n451), .ZN(n1393) );
  OR2_X1 U1224 ( .A1(n450), .A2(n449), .ZN(n1394) );
  OR2_X1 U1225 ( .A1(n751), .A2(n758), .ZN(n1395) );
  OR2_X1 U1226 ( .A1(n457), .A2(n460), .ZN(n1396) );
  OR2_X1 U1227 ( .A1(n767), .A2(n772), .ZN(n1397) );
  OR2_X1 U1228 ( .A1(n779), .A2(n782), .ZN(n1398) );
  OR2_X1 U1229 ( .A1(n787), .A2(n788), .ZN(n1399) );
  AND2_X1 U1230 ( .A1(n663), .A2(n678), .ZN(n1400) );
  AND2_X1 U1231 ( .A1(n822), .A2(n888), .ZN(n1401) );
  BUF_X2 U1232 ( .A(n1285), .Z(n27) );
  OR2_X1 U1233 ( .A1(n1029), .A2(n829), .ZN(n1402) );
  OR2_X1 U1234 ( .A1(n577), .A2(n592), .ZN(n1403) );
  CLKBUF_X1 U1235 ( .A(n1286), .Z(n21) );
  BUF_X1 U1236 ( .A(n1271), .Z(n53) );
  INV_X1 U1237 ( .A(n1400), .ZN(n1404) );
  CLKBUF_X1 U1238 ( .A(b[9]), .Z(n1250) );
  CLKBUF_X1 U1239 ( .A(a[15]), .Z(n1468) );
  XNOR2_X1 U1240 ( .A(n1467), .B(n1248), .ZN(n1405) );
  INV_X2 U1241 ( .A(n1290), .ZN(n1406) );
  CLKBUF_X3 U1242 ( .A(a[19]), .Z(n55) );
  CLKBUF_X1 U1243 ( .A(b[19]), .Z(n1484) );
  XNOR2_X1 U1244 ( .A(n13), .B(n1247), .ZN(n1407) );
  BUF_X2 U1245 ( .A(a[5]), .Z(n13) );
  BUF_X2 U1246 ( .A(n1271), .Z(n1408) );
  NOR2_X1 U1247 ( .A1(n647), .A2(n662), .ZN(n1409) );
  NOR2_X1 U1248 ( .A1(n647), .A2(n662), .ZN(n323) );
  CLKBUF_X1 U1249 ( .A(n1492), .Z(n1410) );
  BUF_X1 U1250 ( .A(n1274), .Z(n1411) );
  BUF_X1 U1251 ( .A(n1274), .Z(n1412) );
  BUF_X2 U1252 ( .A(n1283), .Z(n39) );
  CLKBUF_X1 U1253 ( .A(n1468), .Z(n1413) );
  CLKBUF_X1 U1254 ( .A(n1448), .Z(n1416) );
  CLKBUF_X1 U1255 ( .A(n1281), .Z(n52) );
  XOR2_X1 U1256 ( .A(n630), .B(n615), .Z(n1417) );
  XOR2_X1 U1257 ( .A(n613), .B(n1417), .Z(n611) );
  NAND2_X1 U1258 ( .A1(n613), .A2(n630), .ZN(n1418) );
  NAND2_X1 U1259 ( .A1(n613), .A2(n615), .ZN(n1419) );
  NAND2_X1 U1260 ( .A1(n630), .A2(n615), .ZN(n1420) );
  NAND3_X1 U1261 ( .A1(n1418), .A2(n1419), .A3(n1420), .ZN(n610) );
  BUF_X2 U1262 ( .A(n1282), .Z(n45) );
  CLKBUF_X1 U1263 ( .A(n304), .Z(n1421) );
  OAI22_X1 U1264 ( .A1(n60), .A2(n1031), .B1(n58), .B2(n1030), .ZN(n448) );
  CLKBUF_X2 U1265 ( .A(n1287), .Z(n16) );
  BUF_X1 U1266 ( .A(n1287), .Z(n15) );
  CLKBUF_X3 U1267 ( .A(n1278), .Z(n1451) );
  CLKBUF_X1 U1268 ( .A(b[8]), .Z(n1487) );
  BUF_X4 U1269 ( .A(a[17]), .Z(n49) );
  AND2_X1 U1270 ( .A1(n509), .A2(n520), .ZN(n1422) );
  INV_X1 U1271 ( .A(n316), .ZN(n1423) );
  XOR2_X1 U1272 ( .A(n575), .B(n898), .Z(n1424) );
  XOR2_X1 U1273 ( .A(n1424), .B(n590), .Z(n569) );
  XOR2_X1 U1274 ( .A(n584), .B(n573), .Z(n1425) );
  XOR2_X1 U1275 ( .A(n1425), .B(n569), .Z(n565) );
  NAND2_X1 U1276 ( .A1(n575), .A2(n898), .ZN(n1426) );
  NAND2_X1 U1277 ( .A1(n575), .A2(n590), .ZN(n1427) );
  NAND2_X1 U1278 ( .A1(n898), .A2(n590), .ZN(n1428) );
  NAND3_X1 U1279 ( .A1(n1428), .A2(n1427), .A3(n1426), .ZN(n568) );
  NAND2_X1 U1280 ( .A1(n584), .A2(n573), .ZN(n1429) );
  NAND2_X1 U1281 ( .A1(n584), .A2(n569), .ZN(n1430) );
  NAND2_X1 U1282 ( .A1(n573), .A2(n569), .ZN(n1431) );
  NAND3_X1 U1283 ( .A1(n1429), .A2(n1430), .A3(n1431), .ZN(n564) );
  BUF_X2 U1284 ( .A(n1272), .Z(n1432) );
  XNOR2_X1 U1285 ( .A(n579), .B(n1433), .ZN(n577) );
  XNOR2_X1 U1286 ( .A(n594), .B(n581), .ZN(n1433) );
  NAND2_X1 U1287 ( .A1(n579), .A2(n594), .ZN(n1434) );
  NAND2_X1 U1288 ( .A1(n579), .A2(n581), .ZN(n1435) );
  NAND2_X1 U1289 ( .A1(n594), .A2(n581), .ZN(n1436) );
  NAND3_X1 U1290 ( .A1(n1434), .A2(n1435), .A3(n1436), .ZN(n576) );
  OR2_X1 U1291 ( .A1(n693), .A2(n706), .ZN(n1437) );
  CLKBUF_X1 U1292 ( .A(a[15]), .Z(n43) );
  CLKBUF_X3 U1293 ( .A(n1280), .Z(n57) );
  BUF_X1 U1294 ( .A(n248), .Z(n65) );
  CLKBUF_X1 U1295 ( .A(n340), .Z(n1438) );
  CLKBUF_X1 U1296 ( .A(n7), .Z(n1439) );
  XNOR2_X1 U1297 ( .A(n314), .B(n1440), .ZN(product[20]) );
  AND2_X1 U1298 ( .A1(n428), .A2(n313), .ZN(n1440) );
  OR2_X1 U1299 ( .A1(n312), .A2(n317), .ZN(n1441) );
  BUF_X1 U1300 ( .A(n291), .Z(n63) );
  XNOR2_X1 U1301 ( .A(n298), .B(n1442), .ZN(product[22]) );
  AND2_X1 U1302 ( .A1(n1403), .A2(n297), .ZN(n1442) );
  BUF_X2 U1303 ( .A(n1284), .Z(n33) );
  BUF_X1 U1304 ( .A(n1284), .Z(n34) );
  OAI22_X1 U1305 ( .A1(n48), .A2(n1292), .B1(n1092), .B2(n46), .ZN(n822) );
  BUF_X2 U1306 ( .A(n1279), .Z(n1443) );
  BUF_X4 U1307 ( .A(a[1]), .Z(n1444) );
  CLKBUF_X1 U1308 ( .A(a[1]), .Z(n1) );
  NOR2_X1 U1309 ( .A1(n296), .A2(n303), .ZN(n1445) );
  XNOR2_X1 U1310 ( .A(n305), .B(n1446), .ZN(product[21]) );
  AND2_X1 U1311 ( .A1(n1473), .A2(n1421), .ZN(n1446) );
  CLKBUF_X1 U1312 ( .A(n311), .Z(n1447) );
  BUF_X1 U1313 ( .A(b[3]), .Z(n1256) );
  OR2_X1 U1314 ( .A1(n509), .A2(n520), .ZN(n1449) );
  XNOR2_X1 U1315 ( .A(n244), .B(n1450), .ZN(product[28]) );
  AND2_X1 U1316 ( .A1(n240), .A2(n243), .ZN(n1450) );
  CLKBUF_X1 U1317 ( .A(n1278), .Z(n12) );
  XNOR2_X1 U1318 ( .A(n13), .B(n1241), .ZN(n1452) );
  CLKBUF_X1 U1319 ( .A(n1288), .Z(n9) );
  XNOR2_X1 U1320 ( .A(n1453), .B(n846), .ZN(n607) );
  XNOR2_X1 U1321 ( .A(n900), .B(n972), .ZN(n1453) );
  CLKBUF_X1 U1322 ( .A(n320), .Z(n1454) );
  CLKBUF_X1 U1323 ( .A(n31), .Z(n1455) );
  CLKBUF_X1 U1324 ( .A(n49), .Z(n1456) );
  NOR2_X1 U1325 ( .A1(n611), .A2(n628), .ZN(n1457) );
  NOR2_X1 U1326 ( .A1(n611), .A2(n628), .ZN(n312) );
  BUF_X2 U1327 ( .A(n1285), .Z(n1459) );
  CLKBUF_X1 U1328 ( .A(n1282), .Z(n46) );
  XNOR2_X1 U1329 ( .A(n286), .B(n1460), .ZN(product[24]) );
  AND2_X1 U1330 ( .A1(n424), .A2(n285), .ZN(n1460) );
  BUF_X1 U1331 ( .A(b[0]), .Z(n61) );
  XNOR2_X1 U1332 ( .A(n222), .B(n1461), .ZN(product[30]) );
  AND2_X1 U1333 ( .A1(n418), .A2(n221), .ZN(n1461) );
  XOR2_X1 U1334 ( .A(n822), .B(n888), .Z(n705) );
  BUF_X2 U1335 ( .A(n1274), .Z(n35) );
  NOR2_X2 U1336 ( .A1(n731), .A2(n740), .ZN(n361) );
  CLKBUF_X1 U1337 ( .A(n1416), .Z(n1462) );
  CLKBUF_X3 U1338 ( .A(b[12]), .Z(n1247) );
  XNOR2_X1 U1339 ( .A(n277), .B(n1463), .ZN(product[25]) );
  AND2_X1 U1340 ( .A1(n273), .A2(n276), .ZN(n1463) );
  XNOR2_X1 U1341 ( .A(n268), .B(n1464), .ZN(product[26]) );
  AND2_X1 U1342 ( .A1(n264), .A2(n267), .ZN(n1464) );
  XNOR2_X1 U1343 ( .A(n257), .B(n1465), .ZN(product[27]) );
  AND2_X1 U1344 ( .A1(n421), .A2(n256), .ZN(n1465) );
  CLKBUF_X1 U1345 ( .A(n593), .Z(n1466) );
  OR2_X1 U1346 ( .A1(n266), .A2(n255), .ZN(n251) );
  OAI22_X1 U1347 ( .A1(n42), .A2(n1094), .B1(n40), .B2(n1093), .ZN(n478) );
  NAND2_X1 U1348 ( .A1(n1267), .A2(n1287), .ZN(n1277) );
  CLKBUF_X3 U1349 ( .A(a[13]), .Z(n1469) );
  CLKBUF_X1 U1350 ( .A(a[13]), .Z(n37) );
  BUF_X1 U1351 ( .A(a[7]), .Z(n1470) );
  BUF_X1 U1352 ( .A(n1110), .Z(n1472) );
  BUF_X2 U1353 ( .A(n1286), .Z(n22) );
  BUF_X2 U1354 ( .A(n1276), .Z(n24) );
  OR2_X1 U1355 ( .A1(n1466), .A2(n610), .ZN(n1473) );
  BUF_X1 U1356 ( .A(n1275), .Z(n1474) );
  BUF_X1 U1357 ( .A(n1275), .Z(n1475) );
  CLKBUF_X1 U1358 ( .A(b[19]), .Z(n1240) );
  NOR2_X1 U1359 ( .A1(n577), .A2(n592), .ZN(n1476) );
  NOR2_X1 U1360 ( .A1(n577), .A2(n592), .ZN(n296) );
  NAND2_X1 U1361 ( .A1(n846), .A2(n900), .ZN(n1477) );
  NAND2_X1 U1362 ( .A1(n846), .A2(n972), .ZN(n1478) );
  NAND2_X1 U1363 ( .A1(n900), .A2(n972), .ZN(n1479) );
  NAND3_X1 U1364 ( .A1(n1477), .A2(n1478), .A3(n1479), .ZN(n606) );
  BUF_X2 U1365 ( .A(n1270), .Z(n59) );
  BUF_X2 U1366 ( .A(n1277), .Z(n18) );
  BUF_X4 U1367 ( .A(a[3]), .Z(n7) );
  CLKBUF_X1 U1368 ( .A(b[8]), .Z(n1251) );
  NAND2_X1 U1369 ( .A1(n1266), .A2(n1286), .ZN(n1276) );
  CLKBUF_X3 U1370 ( .A(n1276), .Z(n23) );
  OR2_X2 U1371 ( .A1(n692), .A2(n679), .ZN(n1480) );
  CLKBUF_X1 U1372 ( .A(n336), .Z(n1481) );
  BUF_X4 U1373 ( .A(a[9]), .Z(n25) );
  CLKBUF_X3 U1374 ( .A(b[5]), .Z(n1254) );
  BUF_X4 U1375 ( .A(a[11]), .Z(n31) );
  CLKBUF_X3 U1376 ( .A(b[10]), .Z(n1249) );
  CLKBUF_X3 U1377 ( .A(b[1]), .Z(n1258) );
  BUF_X4 U1378 ( .A(n61), .Z(n1494) );
  XNOR2_X1 U1379 ( .A(n231), .B(n1483), .ZN(product[29]) );
  AND2_X1 U1380 ( .A1(n227), .A2(n230), .ZN(n1483) );
  XNOR2_X1 U1381 ( .A(n209), .B(n1485), .ZN(product[31]) );
  AND2_X1 U1382 ( .A1(n1388), .A2(n208), .ZN(n1485) );
  AOI21_X1 U1383 ( .B1(n1482), .B2(n1481), .A(n1400), .ZN(n1490) );
  BUF_X1 U1384 ( .A(n291), .Z(n1491) );
  BUF_X1 U1385 ( .A(n291), .Z(n1492) );
  NOR2_X1 U1386 ( .A1(n629), .A2(n646), .ZN(n317) );
  NOR2_X1 U1387 ( .A1(n533), .A2(n546), .ZN(n275) );
  NOR2_X1 U1388 ( .A1(n547), .A2(n560), .ZN(n284) );
  NOR2_X1 U1389 ( .A1(n461), .A2(n466), .ZN(n179) );
  NOR2_X1 U1390 ( .A1(n489), .A2(n498), .ZN(n229) );
  NOR2_X1 U1391 ( .A1(n719), .A2(n730), .ZN(n355) );
  NOR2_X1 U1392 ( .A1(n741), .A2(n750), .ZN(n364) );
  NOR2_X1 U1393 ( .A1(n481), .A2(n488), .ZN(n220) );
  NOR2_X1 U1394 ( .A1(n499), .A2(n508), .ZN(n242) );
  NOR2_X1 U1395 ( .A1(n1028), .A2(n1009), .ZN(n406) );
  NOR2_X1 U1396 ( .A1(n773), .A2(n778), .ZN(n386) );
  AND2_X1 U1397 ( .A1(n1402), .A2(n409), .ZN(product[1]) );
  BUF_X1 U1398 ( .A(n1270), .Z(n60) );
  NAND2_X1 U1399 ( .A1(n1284), .A2(n1264), .ZN(n1274) );
  NAND2_X1 U1400 ( .A1(n1269), .A2(n1289), .ZN(n1279) );
  INV_X1 U1401 ( .A(a[0]), .ZN(n1289) );
  NAND2_X1 U1402 ( .A1(n1282), .A2(n1262), .ZN(n1272) );
  NAND2_X1 U1403 ( .A1(n1261), .A2(n1281), .ZN(n1271) );
  NOR2_X1 U1404 ( .A1(n280), .A2(n275), .ZN(n269) );
  NOR2_X1 U1405 ( .A1(n280), .A2(n260), .ZN(n258) );
  NAND2_X1 U1406 ( .A1(n214), .A2(n134), .ZN(n130) );
  INV_X1 U1407 ( .A(n1441), .ZN(n306) );
  INV_X1 U1408 ( .A(n186), .ZN(n184) );
  INV_X1 U1409 ( .A(n173), .ZN(n171) );
  INV_X1 U1410 ( .A(n247), .ZN(n245) );
  INV_X1 U1411 ( .A(n281), .ZN(n279) );
  BUF_X1 U1412 ( .A(n291), .Z(n64) );
  INV_X1 U1413 ( .A(n282), .ZN(n280) );
  INV_X1 U1414 ( .A(n1438), .ZN(n339) );
  NOR2_X1 U1415 ( .A1(n216), .A2(n175), .ZN(n173) );
  NOR2_X1 U1416 ( .A1(n216), .A2(n192), .ZN(n186) );
  INV_X1 U1417 ( .A(n187), .ZN(n185) );
  INV_X1 U1418 ( .A(n1447), .ZN(n309) );
  INV_X1 U1419 ( .A(n283), .ZN(n281) );
  INV_X1 U1420 ( .A(n216), .ZN(n214) );
  NAND2_X1 U1421 ( .A1(n273), .A2(n264), .ZN(n260) );
  OAI21_X1 U1422 ( .B1(n281), .B2(n275), .A(n276), .ZN(n270) );
  OAI21_X1 U1423 ( .B1(n281), .B2(n260), .A(n261), .ZN(n259) );
  AOI21_X1 U1424 ( .B1(n274), .B2(n264), .A(n1383), .ZN(n261) );
  NOR2_X1 U1425 ( .A1(n1441), .A2(n301), .ZN(n299) );
  NAND2_X1 U1426 ( .A1(n1482), .A2(n1480), .ZN(n326) );
  INV_X1 U1427 ( .A(n192), .ZN(n190) );
  INV_X1 U1428 ( .A(n119), .ZN(n117) );
  NAND2_X1 U1429 ( .A1(n186), .A2(n149), .ZN(n145) );
  INV_X1 U1430 ( .A(n1480), .ZN(n333) );
  INV_X1 U1431 ( .A(n1481), .ZN(n334) );
  NAND2_X1 U1432 ( .A1(n214), .A2(n1388), .ZN(n201) );
  INV_X1 U1433 ( .A(n1448), .ZN(n246) );
  NAND2_X1 U1434 ( .A1(n315), .A2(n1423), .ZN(n86) );
  XOR2_X1 U1435 ( .A(n339), .B(n89), .Z(product[16]) );
  NAND2_X1 U1436 ( .A1(n1480), .A2(n338), .ZN(n89) );
  XOR2_X1 U1437 ( .A(n347), .B(n90), .Z(product[15]) );
  NAND2_X1 U1438 ( .A1(n1437), .A2(n346), .ZN(n90) );
  XNOR2_X1 U1439 ( .A(n325), .B(n87), .ZN(product[18]) );
  NAND2_X1 U1440 ( .A1(n430), .A2(n324), .ZN(n87) );
  OAI21_X1 U1441 ( .B1(n339), .B2(n326), .A(n1490), .ZN(n325) );
  INV_X1 U1442 ( .A(n1409), .ZN(n430) );
  INV_X1 U1443 ( .A(n284), .ZN(n424) );
  INV_X1 U1444 ( .A(n255), .ZN(n421) );
  NOR2_X1 U1445 ( .A1(n296), .A2(n303), .ZN(n294) );
  AOI21_X1 U1446 ( .B1(n1445), .B2(n311), .A(n295), .ZN(n293) );
  NAND2_X1 U1447 ( .A1(n294), .A2(n310), .ZN(n292) );
  NOR2_X1 U1448 ( .A1(n216), .A2(n121), .ZN(n119) );
  NAND2_X1 U1449 ( .A1(n425), .A2(n290), .ZN(n82) );
  INV_X1 U1450 ( .A(n289), .ZN(n425) );
  OAI21_X1 U1451 ( .B1(n284), .B2(n290), .A(n285), .ZN(n283) );
  INV_X1 U1452 ( .A(n217), .ZN(n215) );
  OAI21_X1 U1453 ( .B1(n341), .B2(n358), .A(n342), .ZN(n340) );
  XNOR2_X1 U1454 ( .A(n332), .B(n88), .ZN(product[17]) );
  NAND2_X1 U1455 ( .A1(n1482), .A2(n1404), .ZN(n88) );
  OAI21_X1 U1456 ( .B1(n339), .B2(n333), .A(n334), .ZN(n332) );
  NAND2_X1 U1457 ( .A1(n218), .A2(n240), .ZN(n216) );
  AOI21_X1 U1458 ( .B1(n215), .B2(n1388), .A(n206), .ZN(n202) );
  INV_X1 U1459 ( .A(n174), .ZN(n172) );
  XOR2_X1 U1460 ( .A(n352), .B(n91), .Z(product[14]) );
  NAND2_X1 U1461 ( .A1(n434), .A2(n351), .ZN(n91) );
  AOI21_X1 U1462 ( .B1(n357), .B2(n435), .A(n354), .ZN(n352) );
  INV_X1 U1463 ( .A(n350), .ZN(n434) );
  AOI21_X1 U1464 ( .B1(n283), .B2(n249), .A(n250), .ZN(n248) );
  OAI21_X1 U1465 ( .B1(n251), .B2(n276), .A(n252), .ZN(n250) );
  AOI21_X1 U1466 ( .B1(n1449), .B2(n1383), .A(n1422), .ZN(n252) );
  INV_X1 U1467 ( .A(n358), .ZN(n357) );
  NOR2_X1 U1468 ( .A1(n251), .A2(n275), .ZN(n249) );
  INV_X1 U1469 ( .A(n380), .ZN(n379) );
  NOR2_X1 U1470 ( .A1(n192), .A2(n136), .ZN(n134) );
  INV_X1 U1471 ( .A(n275), .ZN(n273) );
  OAI21_X1 U1472 ( .B1(n309), .B2(n301), .A(n1421), .ZN(n300) );
  NAND2_X1 U1473 ( .A1(n1388), .A2(n1391), .ZN(n192) );
  NAND2_X1 U1474 ( .A1(n190), .A2(n177), .ZN(n175) );
  INV_X1 U1475 ( .A(n276), .ZN(n274) );
  INV_X1 U1476 ( .A(n266), .ZN(n264) );
  INV_X1 U1477 ( .A(n1473), .ZN(n301) );
  INV_X1 U1478 ( .A(n193), .ZN(n191) );
  INV_X1 U1479 ( .A(n367), .ZN(n366) );
  INV_X1 U1480 ( .A(n317), .ZN(n315) );
  NAND2_X1 U1481 ( .A1(n240), .A2(n227), .ZN(n225) );
  NAND2_X1 U1482 ( .A1(n173), .A2(n1396), .ZN(n160) );
  AOI21_X1 U1483 ( .B1(n1482), .B2(n336), .A(n1400), .ZN(n327) );
  INV_X1 U1484 ( .A(n290), .ZN(n288) );
  INV_X1 U1485 ( .A(n318), .ZN(n316) );
  INV_X1 U1486 ( .A(n346), .ZN(n344) );
  XOR2_X1 U1487 ( .A(n181), .B(n72), .Z(product[33]) );
  NAND2_X1 U1488 ( .A1(n177), .A2(n180), .ZN(n72) );
  XOR2_X1 U1489 ( .A(n374), .B(n95), .Z(product[10]) );
  NAND2_X1 U1490 ( .A1(n1395), .A2(n373), .ZN(n95) );
  AOI21_X1 U1491 ( .B1(n379), .B2(n1389), .A(n376), .ZN(n374) );
  XNOR2_X1 U1492 ( .A(n357), .B(n92), .ZN(product[13]) );
  NAND2_X1 U1493 ( .A1(n435), .A2(n356), .ZN(n92) );
  INV_X1 U1494 ( .A(n355), .ZN(n435) );
  XNOR2_X1 U1495 ( .A(n363), .B(n93), .ZN(product[12]) );
  NAND2_X1 U1496 ( .A1(n436), .A2(n362), .ZN(n93) );
  OAI21_X1 U1497 ( .B1(n366), .B2(n364), .A(n365), .ZN(n363) );
  INV_X1 U1498 ( .A(n361), .ZN(n436) );
  XNOR2_X1 U1499 ( .A(n379), .B(n96), .ZN(product[9]) );
  NAND2_X1 U1500 ( .A1(n1389), .A2(n378), .ZN(n96) );
  OAI21_X1 U1501 ( .B1(n217), .B2(n175), .A(n176), .ZN(n174) );
  AOI21_X1 U1502 ( .B1(n191), .B2(n177), .A(n178), .ZN(n176) );
  INV_X1 U1503 ( .A(n180), .ZN(n178) );
  AOI21_X1 U1504 ( .B1(n187), .B2(n149), .A(n150), .ZN(n146) );
  AOI21_X1 U1505 ( .B1(n215), .B2(n134), .A(n135), .ZN(n131) );
  INV_X1 U1506 ( .A(n120), .ZN(n118) );
  AOI21_X1 U1507 ( .B1(n174), .B2(n1396), .A(n165), .ZN(n161) );
  NOR2_X1 U1508 ( .A1(n521), .A2(n532), .ZN(n266) );
  AOI21_X1 U1509 ( .B1(n385), .B2(n1397), .A(n382), .ZN(n380) );
  INV_X1 U1510 ( .A(n384), .ZN(n382) );
  OAI21_X1 U1511 ( .B1(n368), .B2(n380), .A(n369), .ZN(n367) );
  NAND2_X1 U1512 ( .A1(n1395), .A2(n1389), .ZN(n368) );
  AOI21_X1 U1513 ( .B1(n1395), .B2(n376), .A(n371), .ZN(n369) );
  AOI21_X1 U1514 ( .B1(n1391), .B2(n206), .A(n195), .ZN(n193) );
  INV_X1 U1515 ( .A(n197), .ZN(n195) );
  INV_X1 U1516 ( .A(n220), .ZN(n418) );
  AOI21_X1 U1517 ( .B1(n218), .B2(n241), .A(n219), .ZN(n217) );
  OAI21_X1 U1518 ( .B1(n230), .B2(n220), .A(n221), .ZN(n219) );
  NOR2_X1 U1519 ( .A1(n593), .A2(n610), .ZN(n303) );
  XOR2_X1 U1520 ( .A(n198), .B(n73), .Z(product[32]) );
  NAND2_X1 U1521 ( .A1(n1391), .A2(n197), .ZN(n73) );
  NOR2_X1 U1522 ( .A1(n561), .A2(n576), .ZN(n289) );
  NOR2_X1 U1523 ( .A1(n229), .A2(n220), .ZN(n218) );
  NOR2_X1 U1524 ( .A1(n179), .A2(n151), .ZN(n149) );
  NOR2_X1 U1525 ( .A1(n707), .A2(n718), .ZN(n350) );
  NOR2_X1 U1526 ( .A1(n509), .A2(n520), .ZN(n255) );
  AOI21_X1 U1527 ( .B1(n241), .B2(n227), .A(n228), .ZN(n226) );
  INV_X1 U1528 ( .A(n230), .ZN(n228) );
  NAND2_X1 U1529 ( .A1(n561), .A2(n576), .ZN(n290) );
  NAND2_X1 U1530 ( .A1(n533), .A2(n546), .ZN(n276) );
  NAND2_X1 U1531 ( .A1(n629), .A2(n646), .ZN(n318) );
  NAND2_X1 U1532 ( .A1(n593), .A2(n610), .ZN(n304) );
  NAND2_X1 U1533 ( .A1(n679), .A2(n692), .ZN(n338) );
  NAND2_X1 U1534 ( .A1(n693), .A2(n706), .ZN(n346) );
  NAND2_X1 U1535 ( .A1(n547), .A2(n560), .ZN(n285) );
  INV_X1 U1536 ( .A(n179), .ZN(n177) );
  INV_X1 U1537 ( .A(n229), .ZN(n227) );
  NAND2_X1 U1538 ( .A1(n149), .A2(n1393), .ZN(n136) );
  NAND2_X1 U1539 ( .A1(n577), .A2(n592), .ZN(n297) );
  NAND2_X1 U1540 ( .A1(n707), .A2(n718), .ZN(n351) );
  NAND2_X1 U1541 ( .A1(n1396), .A2(n1390), .ZN(n151) );
  INV_X1 U1542 ( .A(n242), .ZN(n240) );
  NAND2_X1 U1543 ( .A1(n611), .A2(n628), .ZN(n313) );
  NAND2_X1 U1544 ( .A1(n647), .A2(n662), .ZN(n324) );
  INV_X1 U1545 ( .A(n243), .ZN(n241) );
  INV_X1 U1546 ( .A(n208), .ZN(n206) );
  NAND2_X1 U1547 ( .A1(n119), .A2(n1392), .ZN(n108) );
  INV_X1 U1548 ( .A(n378), .ZN(n376) );
  AOI21_X1 U1549 ( .B1(n1410), .B2(n106), .A(n107), .ZN(n105) );
  XOR2_X1 U1550 ( .A(n366), .B(n94), .Z(product[11]) );
  NAND2_X1 U1551 ( .A1(n437), .A2(n365), .ZN(n94) );
  INV_X1 U1552 ( .A(n364), .ZN(n437) );
  INV_X1 U1553 ( .A(n356), .ZN(n354) );
  INV_X1 U1554 ( .A(n373), .ZN(n371) );
  AOI21_X1 U1555 ( .B1(n135), .B2(n1394), .A(n124), .ZN(n122) );
  INV_X1 U1556 ( .A(n126), .ZN(n124) );
  XOR2_X1 U1557 ( .A(n168), .B(n71), .Z(product[34]) );
  NAND2_X1 U1558 ( .A1(n1396), .A2(n167), .ZN(n71) );
  XOR2_X1 U1559 ( .A(n114), .B(n67), .Z(product[38]) );
  NAND2_X1 U1560 ( .A1(n1392), .A2(n113), .ZN(n67) );
  AOI21_X1 U1561 ( .B1(n64), .B2(n115), .A(n116), .ZN(n114) );
  XOR2_X1 U1562 ( .A(n100), .B(n396), .Z(product[5]) );
  NAND2_X1 U1563 ( .A1(n443), .A2(n395), .ZN(n100) );
  XOR2_X1 U1564 ( .A(n142), .B(n69), .Z(product[36]) );
  NAND2_X1 U1565 ( .A1(n1393), .A2(n141), .ZN(n69) );
  AOI21_X1 U1566 ( .B1(n1410), .B2(n143), .A(n144), .ZN(n142) );
  XOR2_X1 U1567 ( .A(n127), .B(n68), .Z(product[37]) );
  NAND2_X1 U1568 ( .A1(n1394), .A2(n126), .ZN(n68) );
  AOI21_X1 U1569 ( .B1(n1410), .B2(n128), .A(n129), .ZN(n127) );
  AOI21_X1 U1570 ( .B1(n1398), .B2(n393), .A(n390), .ZN(n388) );
  INV_X1 U1571 ( .A(n392), .ZN(n390) );
  XOR2_X1 U1572 ( .A(n157), .B(n70), .Z(product[35]) );
  NAND2_X1 U1573 ( .A1(n1390), .A2(n156), .ZN(n70) );
  AOI21_X1 U1574 ( .B1(n64), .B2(n158), .A(n159), .ZN(n157) );
  OAI21_X1 U1575 ( .B1(n394), .B2(n396), .A(n395), .ZN(n393) );
  OAI21_X1 U1576 ( .B1(n193), .B2(n136), .A(n137), .ZN(n135) );
  AOI21_X1 U1577 ( .B1(n150), .B2(n1393), .A(n139), .ZN(n137) );
  INV_X1 U1578 ( .A(n141), .ZN(n139) );
  OAI21_X1 U1579 ( .B1(n151), .B2(n180), .A(n152), .ZN(n150) );
  AOI21_X1 U1580 ( .B1(n165), .B2(n1390), .A(n154), .ZN(n152) );
  INV_X1 U1581 ( .A(n156), .ZN(n154) );
  OAI21_X1 U1582 ( .B1(n388), .B2(n386), .A(n387), .ZN(n385) );
  NAND2_X1 U1583 ( .A1(n461), .A2(n466), .ZN(n180) );
  NAND2_X1 U1584 ( .A1(n489), .A2(n498), .ZN(n230) );
  AOI21_X1 U1585 ( .B1(n120), .B2(n1392), .A(n111), .ZN(n109) );
  INV_X1 U1586 ( .A(n113), .ZN(n111) );
  NAND2_X1 U1587 ( .A1(n719), .A2(n730), .ZN(n356) );
  NAND2_X1 U1588 ( .A1(n741), .A2(n750), .ZN(n365) );
  NAND2_X1 U1589 ( .A1(n499), .A2(n508), .ZN(n243) );
  NAND2_X1 U1590 ( .A1(n473), .A2(n480), .ZN(n208) );
  NAND2_X1 U1591 ( .A1(n751), .A2(n758), .ZN(n373) );
  NAND2_X1 U1592 ( .A1(n467), .A2(n472), .ZN(n197) );
  NAND2_X1 U1593 ( .A1(n481), .A2(n488), .ZN(n221) );
  NAND2_X1 U1594 ( .A1(n759), .A2(n766), .ZN(n378) );
  NAND2_X1 U1595 ( .A1(n731), .A2(n740), .ZN(n362) );
  INV_X1 U1596 ( .A(n167), .ZN(n165) );
  NAND2_X1 U1597 ( .A1(n441), .A2(n387), .ZN(n98) );
  INV_X1 U1598 ( .A(n386), .ZN(n441) );
  NAND2_X1 U1599 ( .A1(n1398), .A2(n392), .ZN(n99) );
  NAND2_X1 U1600 ( .A1(n1399), .A2(n400), .ZN(n101) );
  INV_X1 U1601 ( .A(n400), .ZN(n398) );
  XOR2_X1 U1602 ( .A(n102), .B(n404), .Z(product[3]) );
  NAND2_X1 U1603 ( .A1(n445), .A2(n403), .ZN(n102) );
  INV_X1 U1604 ( .A(n402), .ZN(n445) );
  XOR2_X1 U1605 ( .A(n103), .B(n409), .Z(product[2]) );
  NAND2_X1 U1606 ( .A1(n446), .A2(n407), .ZN(n103) );
  INV_X1 U1607 ( .A(n406), .ZN(n446) );
  OAI21_X1 U1608 ( .B1(n402), .B2(n404), .A(n403), .ZN(n401) );
  NAND2_X1 U1609 ( .A1(n830), .A2(n448), .ZN(n113) );
  INV_X1 U1610 ( .A(n448), .ZN(n449) );
  INV_X1 U1611 ( .A(n405), .ZN(n404) );
  OAI21_X1 U1612 ( .B1(n406), .B2(n409), .A(n407), .ZN(n405) );
  NAND2_X1 U1613 ( .A1(n1028), .A2(n1009), .ZN(n407) );
  INV_X1 U1614 ( .A(n478), .ZN(n479) );
  OR2_X1 U1615 ( .A1(n937), .A2(n865), .ZN(n626) );
  XNOR2_X1 U1616 ( .A(n937), .B(n865), .ZN(n627) );
  INV_X1 U1617 ( .A(n544), .ZN(n545) );
  NAND2_X1 U1618 ( .A1(n457), .A2(n460), .ZN(n167) );
  NAND2_X1 U1619 ( .A1(n779), .A2(n782), .ZN(n392) );
  NAND2_X1 U1620 ( .A1(n453), .A2(n456), .ZN(n156) );
  NAND2_X1 U1621 ( .A1(n452), .A2(n451), .ZN(n141) );
  NAND2_X1 U1622 ( .A1(n450), .A2(n449), .ZN(n126) );
  NAND2_X1 U1623 ( .A1(n773), .A2(n778), .ZN(n387) );
  NAND2_X1 U1624 ( .A1(n783), .A2(n786), .ZN(n395) );
  OAI22_X1 U1625 ( .A1(n5), .A2(n1237), .B1(n1236), .B2(n3), .ZN(n1028) );
  OAI22_X1 U1626 ( .A1(n24), .A2(n1157), .B1(n22), .B2(n1156), .ZN(n544) );
  OAI22_X1 U1627 ( .A1(n18), .A2(n1452), .B1(n16), .B2(n1177), .ZN(n574) );
  OAI22_X1 U1628 ( .A1(n1475), .A2(n1136), .B1(n1459), .B2(n1135), .ZN(n518)
         );
  OAI22_X1 U1629 ( .A1(n30), .A2(n1143), .B1(n1459), .B2(n1142), .ZN(n937) );
  OAI22_X1 U1630 ( .A1(n1451), .A2(n1199), .B1(n10), .B2(n1198), .ZN(n608) );
  OAI22_X1 U1631 ( .A1(n1432), .A2(n1073), .B1(n46), .B2(n1072), .ZN(n464) );
  OAI22_X1 U1632 ( .A1(n1408), .A2(n1052), .B1(n52), .B2(n1051), .ZN(n454) );
  OAI22_X1 U1633 ( .A1(n36), .A2(n1115), .B1(n34), .B2(n1114), .ZN(n496) );
  OAI22_X1 U1634 ( .A1(n1408), .A2(n1067), .B1(n51), .B2(n1066), .ZN(n865) );
  OAI22_X1 U1635 ( .A1(n24), .A2(n1296), .B1(n1176), .B2(n22), .ZN(n826) );
  OAI22_X1 U1636 ( .A1(n23), .A2(n1175), .B1(n21), .B2(n1174), .ZN(n968) );
  OR2_X1 U1637 ( .A1(n1494), .A2(n1296), .ZN(n1176) );
  OAI22_X1 U1638 ( .A1(n1408), .A2(n1065), .B1(n51), .B2(n1064), .ZN(n863) );
  OAI22_X1 U1639 ( .A1(n24), .A2(n1160), .B1(n22), .B2(n1159), .ZN(n953) );
  OAI22_X1 U1640 ( .A1(n41), .A2(n1106), .B1(n39), .B2(n1105), .ZN(n902) );
  OAI22_X1 U1641 ( .A1(n1443), .A2(n1220), .B1(n1219), .B2(n4), .ZN(n1011) );
  OAI22_X1 U1642 ( .A1(n24), .A2(n1163), .B1(n22), .B2(n1162), .ZN(n956) );
  OAI22_X1 U1643 ( .A1(n17), .A2(n1195), .B1(n15), .B2(n1194), .ZN(n987) );
  OAI22_X1 U1644 ( .A1(n60), .A2(n1034), .B1(n58), .B2(n1033), .ZN(n833) );
  OAI22_X1 U1645 ( .A1(n60), .A2(n1033), .B1(n58), .B2(n1032), .ZN(n832) );
  INV_X1 U1646 ( .A(n454), .ZN(n455) );
  OAI22_X1 U1647 ( .A1(n1451), .A2(n1216), .B1(n9), .B2(n1215), .ZN(n1007) );
  AND2_X1 U1648 ( .A1(n1495), .A2(n812), .ZN(n989) );
  OAI22_X1 U1649 ( .A1(n1443), .A2(n1235), .B1(n1234), .B2(n3), .ZN(n1026) );
  OAI22_X1 U1650 ( .A1(n1474), .A2(n1295), .B1(n1155), .B2(n1459), .ZN(n825)
         );
  OAI22_X1 U1651 ( .A1(n29), .A2(n1154), .B1(n27), .B2(n1153), .ZN(n948) );
  OR2_X1 U1652 ( .A1(n1495), .A2(n1295), .ZN(n1155) );
  OAI22_X1 U1653 ( .A1(n1474), .A2(n1152), .B1(n27), .B2(n1151), .ZN(n946) );
  OAI22_X1 U1654 ( .A1(n1443), .A2(n1228), .B1(n1227), .B2(n4), .ZN(n1019) );
  OAI22_X1 U1655 ( .A1(n17), .A2(n1190), .B1(n15), .B2(n1189), .ZN(n982) );
  OAI22_X1 U1656 ( .A1(n17), .A2(n1297), .B1(n1197), .B2(n16), .ZN(n827) );
  OAI22_X1 U1657 ( .A1(n17), .A2(n1196), .B1(n15), .B2(n1195), .ZN(n988) );
  OR2_X1 U1658 ( .A1(n1494), .A2(n1297), .ZN(n1197) );
  OAI22_X1 U1659 ( .A1(n30), .A2(n1139), .B1(n1459), .B2(n1138), .ZN(n933) );
  OAI22_X1 U1660 ( .A1(n24), .A2(n1158), .B1(n22), .B2(n1157), .ZN(n951) );
  OAI22_X1 U1661 ( .A1(n54), .A2(n1063), .B1(n51), .B2(n1062), .ZN(n861) );
  OAI22_X1 U1662 ( .A1(n30), .A2(n1142), .B1(n1459), .B2(n1141), .ZN(n936) );
  INV_X1 U1663 ( .A(n608), .ZN(n609) );
  OAI22_X1 U1664 ( .A1(n1411), .A2(n1123), .B1(n34), .B2(n1122), .ZN(n918) );
  OAI22_X1 U1665 ( .A1(n1475), .A2(n1153), .B1(n27), .B2(n1152), .ZN(n947) );
  OAI22_X1 U1666 ( .A1(n11), .A2(n1210), .B1(n9), .B2(n1209), .ZN(n1001) );
  OAI22_X1 U1667 ( .A1(n17), .A2(n1191), .B1(n15), .B2(n1190), .ZN(n983) );
  OAI22_X1 U1668 ( .A1(n1451), .A2(n1213), .B1(n9), .B2(n1212), .ZN(n1004) );
  OAI22_X1 U1669 ( .A1(n17), .A2(n1194), .B1(n15), .B2(n1193), .ZN(n986) );
  OAI22_X1 U1670 ( .A1(n5), .A2(n1232), .B1(n1231), .B2(n3), .ZN(n1023) );
  OAI22_X1 U1671 ( .A1(n1474), .A2(n1140), .B1(n1459), .B2(n1139), .ZN(n934)
         );
  OAI22_X1 U1672 ( .A1(n24), .A2(n1159), .B1(n22), .B2(n1158), .ZN(n952) );
  OAI22_X1 U1673 ( .A1(n1432), .A2(n1083), .B1(n45), .B2(n1082), .ZN(n880) );
  OAI22_X1 U1674 ( .A1(n59), .A2(n1041), .B1(n57), .B2(n1040), .ZN(n840) );
  INV_X1 U1675 ( .A(n518), .ZN(n519) );
  OAI22_X1 U1676 ( .A1(n54), .A2(n1060), .B1(n52), .B2(n1059), .ZN(n858) );
  OAI22_X1 U1677 ( .A1(n42), .A2(n1098), .B1(n40), .B2(n1097), .ZN(n894) );
  OAI22_X1 U1678 ( .A1(n1411), .A2(n1117), .B1(n34), .B2(n1116), .ZN(n912) );
  OAI22_X1 U1679 ( .A1(n1432), .A2(n1079), .B1(n46), .B2(n1078), .ZN(n876) );
  OAI22_X1 U1680 ( .A1(n60), .A2(n1037), .B1(n58), .B2(n1036), .ZN(n836) );
  OAI22_X1 U1681 ( .A1(n1432), .A2(n1075), .B1(n46), .B2(n1074), .ZN(n872) );
  OAI22_X1 U1682 ( .A1(n1408), .A2(n1056), .B1(n52), .B2(n1055), .ZN(n854) );
  OAI22_X1 U1683 ( .A1(n1432), .A2(n1091), .B1(n45), .B2(n1090), .ZN(n888) );
  OR2_X1 U1684 ( .A1(n1495), .A2(n1292), .ZN(n1092) );
  NOR2_X1 U1685 ( .A1(n789), .A2(n828), .ZN(n402) );
  AND2_X1 U1686 ( .A1(n1495), .A2(n800), .ZN(n909) );
  OAI22_X1 U1687 ( .A1(n30), .A2(n1151), .B1(n27), .B2(n1150), .ZN(n945) );
  OAI22_X1 U1688 ( .A1(n5), .A2(n1227), .B1(n1226), .B2(n4), .ZN(n1018) );
  AOI21_X1 U1689 ( .B1(n42), .B2(n40), .A(n1093), .ZN(n799) );
  AOI21_X1 U1690 ( .B1(n6), .B2(n4), .A(n1219), .ZN(n817) );
  AOI21_X1 U1691 ( .B1(n1411), .B2(n34), .A(n1114), .ZN(n802) );
  AOI21_X1 U1692 ( .B1(n12), .B2(n10), .A(n1198), .ZN(n814) );
  OAI22_X1 U1693 ( .A1(n53), .A2(n1291), .B1(n1071), .B2(n52), .ZN(n821) );
  OAI22_X1 U1694 ( .A1(n1408), .A2(n1070), .B1(n51), .B2(n1069), .ZN(n868) );
  OR2_X1 U1695 ( .A1(n1495), .A2(n1291), .ZN(n1071) );
  NAND2_X1 U1696 ( .A1(n1029), .A2(n829), .ZN(n409) );
  OAI22_X1 U1697 ( .A1(n11), .A2(n1215), .B1(n9), .B2(n1214), .ZN(n1006) );
  OAI22_X1 U1698 ( .A1(n1443), .A2(n1234), .B1(n1233), .B2(n3), .ZN(n1025) );
  AND2_X1 U1699 ( .A1(n1495), .A2(n815), .ZN(n1009) );
  INV_X1 U1700 ( .A(n9), .ZN(n815) );
  OAI22_X1 U1701 ( .A1(n29), .A2(n1137), .B1(n1459), .B2(n1136), .ZN(n931) );
  OAI22_X1 U1702 ( .A1(n35), .A2(n1118), .B1(n34), .B2(n1117), .ZN(n913) );
  OAI22_X1 U1703 ( .A1(n53), .A2(n1061), .B1(n51), .B2(n1060), .ZN(n859) );
  OAI22_X1 U1704 ( .A1(n42), .A2(n1100), .B1(n40), .B2(n1099), .ZN(n896) );
  OAI22_X1 U1705 ( .A1(n1474), .A2(n1138), .B1(n1459), .B2(n1137), .ZN(n932)
         );
  OAI22_X1 U1706 ( .A1(n35), .A2(n1119), .B1(n34), .B2(n1118), .ZN(n914) );
  OAI22_X1 U1707 ( .A1(n1475), .A2(n1146), .B1(n27), .B2(n1145), .ZN(n940) );
  OAI22_X1 U1708 ( .A1(n1451), .A2(n1203), .B1(n10), .B2(n1202), .ZN(n994) );
  OAI22_X1 U1709 ( .A1(n1443), .A2(n1222), .B1(n1221), .B2(n4), .ZN(n1013) );
  OAI22_X1 U1710 ( .A1(n42), .A2(n1099), .B1(n40), .B2(n1098), .ZN(n895) );
  OAI22_X1 U1711 ( .A1(n48), .A2(n1080), .B1(n46), .B2(n1079), .ZN(n877) );
  OAI22_X1 U1712 ( .A1(n1408), .A2(n1057), .B1(n52), .B2(n1056), .ZN(n855) );
  OAI22_X1 U1713 ( .A1(n1432), .A2(n1076), .B1(n46), .B2(n1075), .ZN(n873) );
  OAI22_X1 U1714 ( .A1(n41), .A2(n1103), .B1(n39), .B2(n1102), .ZN(n899) );
  OAI22_X1 U1715 ( .A1(n29), .A2(n1141), .B1(n1459), .B2(n1140), .ZN(n935) );
  OAI22_X1 U1716 ( .A1(n48), .A2(n1084), .B1(n45), .B2(n1083), .ZN(n881) );
  AND2_X1 U1717 ( .A1(n1495), .A2(n791), .ZN(n849) );
  OAI22_X1 U1718 ( .A1(n6), .A2(n1221), .B1(n1220), .B2(n4), .ZN(n1012) );
  OAI22_X1 U1719 ( .A1(n47), .A2(n1088), .B1(n1087), .B2(n45), .ZN(n885) );
  OAI22_X1 U1720 ( .A1(n11), .A2(n1201), .B1(n10), .B2(n1200), .ZN(n992) );
  OAI22_X1 U1721 ( .A1(n17), .A2(n1182), .B1(n16), .B2(n1181), .ZN(n974) );
  OAI22_X1 U1722 ( .A1(n1412), .A2(n1125), .B1(n33), .B2(n1124), .ZN(n920) );
  OAI22_X1 U1723 ( .A1(n41), .A2(n1108), .B1(n39), .B2(n1107), .ZN(n904) );
  OAI22_X1 U1724 ( .A1(n1412), .A2(n1127), .B1(n33), .B2(n1126), .ZN(n922) );
  OAI22_X1 U1725 ( .A1(n1432), .A2(n1089), .B1(n45), .B2(n1088), .ZN(n886) );
  OAI22_X1 U1726 ( .A1(n48), .A2(n1077), .B1(n46), .B2(n1076), .ZN(n874) );
  INV_X1 U1727 ( .A(n496), .ZN(n497) );
  OAI22_X1 U1728 ( .A1(n1408), .A2(n1059), .B1(n52), .B2(n1058), .ZN(n857) );
  OAI22_X1 U1729 ( .A1(n36), .A2(n1116), .B1(n34), .B2(n1115), .ZN(n911) );
  OAI22_X1 U1730 ( .A1(n48), .A2(n1078), .B1(n46), .B2(n1077), .ZN(n875) );
  OAI22_X1 U1731 ( .A1(n41), .A2(n1107), .B1(n39), .B2(n1106), .ZN(n903) );
  OAI22_X1 U1732 ( .A1(n1451), .A2(n1202), .B1(n10), .B2(n1201), .ZN(n993) );
  OAI22_X1 U1733 ( .A1(n1408), .A2(n1069), .B1(n51), .B2(n1068), .ZN(n867) );
  INV_X1 U1734 ( .A(n15), .ZN(n812) );
  INV_X1 U1735 ( .A(n21), .ZN(n809) );
  OAI22_X1 U1736 ( .A1(n1475), .A2(n1147), .B1(n27), .B2(n1146), .ZN(n941) );
  OAI22_X1 U1737 ( .A1(n23), .A2(n1166), .B1(n22), .B2(n1165), .ZN(n959) );
  OAI22_X1 U1738 ( .A1(n18), .A2(n1185), .B1(n16), .B2(n1184), .ZN(n977) );
  OAI22_X1 U1739 ( .A1(n59), .A2(n1047), .B1(n57), .B2(n1046), .ZN(n846) );
  OAI22_X1 U1740 ( .A1(n41), .A2(n1104), .B1(n39), .B2(n1103), .ZN(n900) );
  OAI22_X1 U1741 ( .A1(n18), .A2(n1180), .B1(n16), .B2(n1179), .ZN(n972) );
  OAI22_X1 U1742 ( .A1(n1412), .A2(n1122), .B1(n34), .B2(n1121), .ZN(n917) );
  OAI22_X1 U1743 ( .A1(n24), .A2(n1164), .B1(n22), .B2(n1163), .ZN(n957) );
  OAI22_X1 U1744 ( .A1(n59), .A2(n1045), .B1(n57), .B2(n1044), .ZN(n844) );
  OAI22_X1 U1745 ( .A1(n1408), .A2(n1064), .B1(n51), .B2(n1063), .ZN(n862) );
  OAI22_X1 U1746 ( .A1(n36), .A2(n1121), .B1(n34), .B2(n1120), .ZN(n916) );
  OAI22_X1 U1747 ( .A1(n17), .A2(n1407), .B1(n16), .B2(n1183), .ZN(n976) );
  OAI22_X1 U1748 ( .A1(n24), .A2(n1165), .B1(n22), .B2(n1164), .ZN(n958) );
  OAI22_X1 U1749 ( .A1(n11), .A2(n1211), .B1(n9), .B2(n1210), .ZN(n1002) );
  OAI22_X1 U1750 ( .A1(n17), .A2(n1192), .B1(n15), .B2(n1191), .ZN(n984) );
  OAI22_X1 U1751 ( .A1(n23), .A2(n1173), .B1(n21), .B2(n1172), .ZN(n966) );
  OAI22_X1 U1752 ( .A1(n30), .A2(n1144), .B1(n27), .B2(n1143), .ZN(n938) );
  OAI22_X1 U1753 ( .A1(n47), .A2(n1087), .B1(n45), .B2(n1086), .ZN(n884) );
  OAI22_X1 U1754 ( .A1(n53), .A2(n1068), .B1(n1067), .B2(n51), .ZN(n866) );
  OAI22_X1 U1755 ( .A1(n1110), .A2(n41), .B1(n39), .B2(n1109), .ZN(n906) );
  OAI22_X1 U1756 ( .A1(n1129), .A2(n35), .B1(n33), .B2(n1128), .ZN(n924) );
  OAI22_X1 U1757 ( .A1(n23), .A2(n1167), .B1(n21), .B2(n1166), .ZN(n960) );
  OAI22_X1 U1758 ( .A1(n1475), .A2(n1150), .B1(n27), .B2(n1149), .ZN(n944) );
  OAI22_X1 U1759 ( .A1(n17), .A2(n1188), .B1(n15), .B2(n1187), .ZN(n980) );
  OAI22_X1 U1760 ( .A1(n1412), .A2(n1131), .B1(n33), .B2(n1130), .ZN(n926) );
  OAI22_X1 U1761 ( .A1(n42), .A2(n1095), .B1(n40), .B2(n1094), .ZN(n891) );
  OAI22_X1 U1762 ( .A1(n60), .A2(n1038), .B1(n58), .B2(n1037), .ZN(n837) );
  INV_X1 U1763 ( .A(n802), .ZN(n910) );
  OAI22_X1 U1764 ( .A1(n59), .A2(n1044), .B1(n57), .B2(n1043), .ZN(n843) );
  INV_X1 U1765 ( .A(n811), .ZN(n970) );
  AOI21_X1 U1766 ( .B1(n18), .B2(n16), .A(n1177), .ZN(n811) );
  OAI22_X1 U1767 ( .A1(n17), .A2(n1187), .B1(n15), .B2(n1186), .ZN(n979) );
  OAI22_X1 U1768 ( .A1(n23), .A2(n1168), .B1(n21), .B2(n1167), .ZN(n961) );
  OAI22_X1 U1769 ( .A1(n1451), .A2(n1212), .B1(n9), .B2(n1211), .ZN(n1003) );
  OAI22_X1 U1770 ( .A1(n23), .A2(n1174), .B1(n21), .B2(n1173), .ZN(n967) );
  OAI22_X1 U1771 ( .A1(n59), .A2(n1042), .B1(n57), .B2(n1041), .ZN(n841) );
  INV_X1 U1772 ( .A(n808), .ZN(n950) );
  AOI21_X1 U1773 ( .B1(n24), .B2(n22), .A(n1156), .ZN(n808) );
  OAI22_X1 U1774 ( .A1(n1451), .A2(n1214), .B1(n9), .B2(n1213), .ZN(n1005) );
  AND2_X1 U1775 ( .A1(n1495), .A2(n809), .ZN(n969) );
  OAI22_X1 U1776 ( .A1(n5), .A2(n1233), .B1(n1232), .B2(n3), .ZN(n1024) );
  OAI22_X1 U1777 ( .A1(n5), .A2(n1230), .B1(n1229), .B2(n3), .ZN(n1021) );
  OAI22_X1 U1778 ( .A1(n11), .A2(n1205), .B1(n10), .B2(n1204), .ZN(n996) );
  OAI22_X1 U1779 ( .A1(n42), .A2(n1101), .B1(n40), .B2(n1100), .ZN(n897) );
  OAI22_X1 U1780 ( .A1(n1432), .A2(n1082), .B1(n45), .B2(n1081), .ZN(n879) );
  OAI22_X1 U1781 ( .A1(n1412), .A2(n1120), .B1(n34), .B2(n1119), .ZN(n915) );
  AND2_X1 U1782 ( .A1(n1495), .A2(n803), .ZN(n929) );
  OAI22_X1 U1783 ( .A1(n1443), .A2(n1229), .B1(n1228), .B2(n3), .ZN(n1020) );
  OAI22_X1 U1784 ( .A1(n23), .A2(n1172), .B1(n21), .B2(n1171), .ZN(n965) );
  OAI22_X1 U1785 ( .A1(n29), .A2(n1145), .B1(n27), .B2(n1144), .ZN(n939) );
  OAI22_X1 U1786 ( .A1(n18), .A2(n1183), .B1(n16), .B2(n1182), .ZN(n975) );
  OAI22_X1 U1787 ( .A1(n36), .A2(n1126), .B1(n33), .B2(n1125), .ZN(n921) );
  OAI22_X1 U1788 ( .A1(n59), .A2(n1043), .B1(n57), .B2(n1042), .ZN(n842) );
  OAI22_X1 U1789 ( .A1(n1408), .A2(n1062), .B1(n51), .B2(n1061), .ZN(n860) );
  OAI22_X1 U1790 ( .A1(n1432), .A2(n1081), .B1(n46), .B2(n1080), .ZN(n878) );
  AND2_X1 U1791 ( .A1(n1495), .A2(n797), .ZN(n889) );
  OAI22_X1 U1792 ( .A1(n5), .A2(n1225), .B1(n1224), .B2(n4), .ZN(n1016) );
  OAI22_X1 U1793 ( .A1(n1411), .A2(n1130), .B1(n1129), .B2(n33), .ZN(n925) );
  OAI22_X1 U1794 ( .A1(n60), .A2(n1039), .B1(n58), .B2(n1038), .ZN(n838) );
  OAI22_X1 U1795 ( .A1(n42), .A2(n1096), .B1(n40), .B2(n1095), .ZN(n892) );
  OAI22_X1 U1796 ( .A1(n54), .A2(n1058), .B1(n52), .B2(n1057), .ZN(n856) );
  OAI22_X1 U1797 ( .A1(n1451), .A2(n1207), .B1(n10), .B2(n1206), .ZN(n998) );
  OAI22_X1 U1798 ( .A1(n1443), .A2(n1226), .B1(n1225), .B2(n4), .ZN(n1017) );
  OAI22_X1 U1799 ( .A1(n23), .A2(n1169), .B1(n21), .B2(n1168), .ZN(n962) );
  OAI22_X1 U1800 ( .A1(n41), .A2(n1109), .B1(n1108), .B2(n39), .ZN(n905) );
  AND2_X1 U1801 ( .A1(n1495), .A2(n794), .ZN(n869) );
  OAI22_X1 U1802 ( .A1(n6), .A2(n1223), .B1(n1222), .B2(n4), .ZN(n1014) );
  OAI22_X1 U1803 ( .A1(n29), .A2(n1149), .B1(n27), .B2(n1148), .ZN(n943) );
  OAI22_X1 U1804 ( .A1(n41), .A2(n1111), .B1(n39), .B2(n1472), .ZN(n907) );
  OAI22_X1 U1805 ( .A1(n1451), .A2(n1206), .B1(n10), .B2(n1205), .ZN(n997) );
  OAI22_X1 U1806 ( .A1(n60), .A2(n1036), .B1(n58), .B2(n1035), .ZN(n835) );
  INV_X1 U1807 ( .A(n799), .ZN(n890) );
  OAI22_X1 U1808 ( .A1(n1408), .A2(n1055), .B1(n52), .B2(n1054), .ZN(n853) );
  OAI22_X1 U1809 ( .A1(n17), .A2(n1181), .B1(n16), .B2(n1180), .ZN(n973) );
  OAI22_X1 U1810 ( .A1(n24), .A2(n1162), .B1(n22), .B2(n1161), .ZN(n955) );
  OAI22_X1 U1811 ( .A1(n1432), .A2(n1074), .B1(n46), .B2(n1073), .ZN(n871) );
  OAI22_X1 U1812 ( .A1(n11), .A2(n1208), .B1(n9), .B2(n1207), .ZN(n999) );
  OAI22_X1 U1813 ( .A1(n23), .A2(n1170), .B1(n21), .B2(n1169), .ZN(n963) );
  OAI22_X1 U1814 ( .A1(n1411), .A2(n1132), .B1(n33), .B2(n1131), .ZN(n927) );
  OAI22_X1 U1815 ( .A1(n1474), .A2(n1148), .B1(n27), .B2(n1147), .ZN(n942) );
  OAI22_X1 U1816 ( .A1(n18), .A2(n1186), .B1(n16), .B2(n1405), .ZN(n978) );
  OAI22_X1 U1817 ( .A1(n1443), .A2(n1224), .B1(n1223), .B2(n4), .ZN(n1015) );
  OAI22_X1 U1818 ( .A1(n42), .A2(n1097), .B1(n40), .B2(n1096), .ZN(n893) );
  OAI22_X1 U1819 ( .A1(n1451), .A2(n1209), .B1(n9), .B2(n1208), .ZN(n1000) );
  OAI22_X1 U1820 ( .A1(n23), .A2(n1171), .B1(n21), .B2(n1170), .ZN(n964) );
  OAI22_X1 U1821 ( .A1(n42), .A2(n1102), .B1(n40), .B2(n1101), .ZN(n898) );
  INV_X1 U1822 ( .A(n574), .ZN(n575) );
  OAI22_X1 U1823 ( .A1(n17), .A2(n1189), .B1(n15), .B2(n1188), .ZN(n981) );
  OAI22_X1 U1824 ( .A1(n59), .A2(n1046), .B1(n1045), .B2(n57), .ZN(n845) );
  INV_X1 U1825 ( .A(n814), .ZN(n990) );
  OAI22_X1 U1826 ( .A1(n18), .A2(n1179), .B1(n16), .B2(n1178), .ZN(n971) );
  OAI22_X1 U1827 ( .A1(n41), .A2(n1105), .B1(n39), .B2(n1104), .ZN(n901) );
  OAI22_X1 U1828 ( .A1(n1451), .A2(n1200), .B1(n10), .B2(n1199), .ZN(n991) );
  OAI22_X1 U1829 ( .A1(n1432), .A2(n1086), .B1(n45), .B2(n1085), .ZN(n883) );
  OAI22_X1 U1830 ( .A1(n48), .A2(n1085), .B1(n45), .B2(n1084), .ZN(n882) );
  OAI22_X1 U1831 ( .A1(n24), .A2(n1161), .B1(n22), .B2(n1160), .ZN(n954) );
  OAI22_X1 U1832 ( .A1(n53), .A2(n1066), .B1(n1065), .B2(n51), .ZN(n864) );
  OAI22_X1 U1833 ( .A1(n12), .A2(n1204), .B1(n10), .B2(n1203), .ZN(n995) );
  OAI22_X1 U1834 ( .A1(n35), .A2(n1128), .B1(n33), .B2(n1127), .ZN(n923) );
  OAI22_X1 U1835 ( .A1(n47), .A2(n1090), .B1(n45), .B2(n1089), .ZN(n887) );
  AND2_X1 U1836 ( .A1(n1495), .A2(n806), .ZN(n949) );
  OAI22_X1 U1837 ( .A1(n1443), .A2(n1231), .B1(n1230), .B2(n3), .ZN(n1022) );
  OAI22_X1 U1838 ( .A1(n17), .A2(n1193), .B1(n15), .B2(n1192), .ZN(n985) );
  NAND2_X1 U1839 ( .A1(n787), .A2(n788), .ZN(n400) );
  OAI22_X1 U1840 ( .A1(n60), .A2(n1290), .B1(n1050), .B2(n58), .ZN(n820) );
  OAI22_X1 U1841 ( .A1(n59), .A2(n1049), .B1(n57), .B2(n1048), .ZN(n848) );
  OR2_X1 U1842 ( .A1(n1494), .A2(n1290), .ZN(n1050) );
  OAI22_X1 U1843 ( .A1(n42), .A2(n1293), .B1(n1113), .B2(n40), .ZN(n823) );
  OAI22_X1 U1844 ( .A1(n41), .A2(n1112), .B1(n39), .B2(n1111), .ZN(n908) );
  OR2_X1 U1845 ( .A1(n1495), .A2(n1293), .ZN(n1113) );
  INV_X1 U1846 ( .A(n790), .ZN(n830) );
  AOI21_X1 U1847 ( .B1(n60), .B2(n58), .A(n1030), .ZN(n790) );
  INV_X1 U1848 ( .A(n27), .ZN(n806) );
  OAI22_X1 U1849 ( .A1(n60), .A2(n1035), .B1(n58), .B2(n1034), .ZN(n834) );
  OAI22_X1 U1850 ( .A1(n54), .A2(n1054), .B1(n52), .B2(n1053), .ZN(n852) );
  INV_X1 U1851 ( .A(n464), .ZN(n465) );
  OR2_X1 U1852 ( .A1(n1495), .A2(n1294), .ZN(n1134) );
  OAI22_X1 U1853 ( .A1(n59), .A2(n1040), .B1(n57), .B2(n1039), .ZN(n839) );
  INV_X1 U1854 ( .A(n805), .ZN(n930) );
  AOI21_X1 U1855 ( .B1(n30), .B2(n1459), .A(n1135), .ZN(n805) );
  OAI22_X1 U1856 ( .A1(n54), .A2(n1053), .B1(n52), .B2(n1052), .ZN(n851) );
  INV_X1 U1857 ( .A(n796), .ZN(n870) );
  AOI21_X1 U1858 ( .B1(n48), .B2(n46), .A(n1072), .ZN(n796) );
  OAI22_X1 U1859 ( .A1(n60), .A2(n1032), .B1(n58), .B2(n1031), .ZN(n831) );
  INV_X1 U1860 ( .A(n793), .ZN(n850) );
  AOI21_X1 U1861 ( .B1(n54), .B2(n52), .A(n1051), .ZN(n793) );
  OAI22_X1 U1862 ( .A1(n1048), .A2(n59), .B1(n1047), .B2(n57), .ZN(n847) );
  OAI22_X1 U1863 ( .A1(n35), .A2(n1124), .B1(n33), .B2(n1123), .ZN(n919) );
  INV_X1 U1864 ( .A(n817), .ZN(n1010) );
  INV_X1 U1865 ( .A(n45), .ZN(n797) );
  INV_X1 U1866 ( .A(n39), .ZN(n800) );
  INV_X1 U1867 ( .A(n51), .ZN(n794) );
  INV_X1 U1868 ( .A(n33), .ZN(n803) );
  INV_X1 U1869 ( .A(n57), .ZN(n791) );
  AND2_X1 U1870 ( .A1(n1495), .A2(a[0]), .ZN(product[0]) );
  INV_X1 U1871 ( .A(n1444), .ZN(n1299) );
  OAI22_X1 U1872 ( .A1(n11), .A2(n1298), .B1(n1218), .B2(n10), .ZN(n828) );
  OR2_X1 U1873 ( .A1(n1494), .A2(n1298), .ZN(n1218) );
  INV_X1 U1874 ( .A(n1439), .ZN(n1298) );
  OAI22_X1 U1875 ( .A1(n1443), .A2(n1238), .B1(n1237), .B2(n3), .ZN(n1029) );
  OAI22_X1 U1876 ( .A1(n1451), .A2(n1217), .B1(n9), .B2(n1216), .ZN(n1008) );
  OAI22_X1 U1877 ( .A1(n1443), .A2(n1236), .B1(n1235), .B2(n3), .ZN(n1027) );
  XNOR2_X1 U1878 ( .A(n7), .B(n1494), .ZN(n1217) );
  OAI22_X1 U1879 ( .A1(n36), .A2(n1133), .B1(n33), .B2(n1132), .ZN(n928) );
  OAI22_X1 U1880 ( .A1(n1411), .A2(n1294), .B1(n1134), .B2(n34), .ZN(n824) );
  XNOR2_X1 U1881 ( .A(n31), .B(n1494), .ZN(n1133) );
  XNOR2_X1 U1882 ( .A(n7), .B(n1245), .ZN(n1203) );
  XNOR2_X1 U1883 ( .A(n7), .B(n1246), .ZN(n1204) );
  XNOR2_X1 U1884 ( .A(n31), .B(n1243), .ZN(n1117) );
  XNOR2_X1 U1885 ( .A(n31), .B(n1254), .ZN(n1128) );
  XNOR2_X1 U1886 ( .A(n31), .B(n1253), .ZN(n1127) );
  XNOR2_X1 U1887 ( .A(n31), .B(n1255), .ZN(n1129) );
  XNOR2_X1 U1888 ( .A(n31), .B(n1249), .ZN(n1123) );
  XNOR2_X1 U1889 ( .A(n31), .B(n1244), .ZN(n1118) );
  XNOR2_X1 U1890 ( .A(n31), .B(n1489), .ZN(n1124) );
  XNOR2_X1 U1891 ( .A(n31), .B(n1245), .ZN(n1119) );
  XNOR2_X1 U1892 ( .A(n31), .B(n1246), .ZN(n1120) );
  XNOR2_X1 U1893 ( .A(n7), .B(n1486), .ZN(n1215) );
  XNOR2_X1 U1894 ( .A(n7), .B(n1258), .ZN(n1216) );
  XNOR2_X1 U1895 ( .A(n31), .B(n1251), .ZN(n1125) );
  XNOR2_X1 U1896 ( .A(n7), .B(n1255), .ZN(n1213) );
  XNOR2_X1 U1897 ( .A(n7), .B(n1242), .ZN(n1200) );
  XNOR2_X1 U1898 ( .A(n7), .B(n1488), .ZN(n1214) );
  XNOR2_X1 U1899 ( .A(n7), .B(n1252), .ZN(n1210) );
  XNOR2_X1 U1900 ( .A(n7), .B(n1241), .ZN(n1199) );
  XNOR2_X1 U1901 ( .A(n7), .B(n1243), .ZN(n1201) );
  XNOR2_X1 U1902 ( .A(n7), .B(n1253), .ZN(n1211) );
  XNOR2_X1 U1903 ( .A(n31), .B(n1488), .ZN(n1130) );
  XNOR2_X1 U1904 ( .A(n31), .B(n1247), .ZN(n1121) );
  XNOR2_X1 U1905 ( .A(n31), .B(n1242), .ZN(n1116) );
  XNOR2_X1 U1906 ( .A(n31), .B(n1252), .ZN(n1126) );
  XNOR2_X1 U1907 ( .A(n7), .B(n1244), .ZN(n1202) );
  XNOR2_X1 U1908 ( .A(n31), .B(n1486), .ZN(n1131) );
  XNOR2_X1 U1909 ( .A(n7), .B(n1248), .ZN(n1206) );
  XNOR2_X1 U1910 ( .A(n7), .B(n1249), .ZN(n1207) );
  XNOR2_X1 U1911 ( .A(n1455), .B(n1241), .ZN(n1115) );
  XNOR2_X1 U1912 ( .A(n31), .B(n1258), .ZN(n1132) );
  XNOR2_X1 U1913 ( .A(n31), .B(n1248), .ZN(n1122) );
  XNOR2_X1 U1914 ( .A(n7), .B(n1247), .ZN(n1205) );
  XNOR2_X1 U1915 ( .A(n7), .B(n1250), .ZN(n1208) );
  XNOR2_X1 U1916 ( .A(n1439), .B(n1487), .ZN(n1209) );
  XNOR2_X1 U1917 ( .A(n1439), .B(n1254), .ZN(n1212) );
  XNOR2_X1 U1918 ( .A(n7), .B(n1240), .ZN(n1198) );
  XNOR2_X1 U1919 ( .A(n1455), .B(n1458), .ZN(n1114) );
  BUF_X1 U1920 ( .A(n1283), .Z(n40) );
  BUF_X1 U1921 ( .A(n1288), .Z(n10) );
  BUF_X1 U1922 ( .A(n1280), .Z(n58) );
  BUF_X1 U1923 ( .A(n1275), .Z(n29) );
  BUF_X1 U1924 ( .A(n1278), .Z(n11) );
  BUF_X1 U1925 ( .A(n61), .Z(n1495) );
  INV_X1 U1926 ( .A(n31), .ZN(n1294) );
  BUF_X1 U1927 ( .A(n1289), .Z(n3) );
  BUF_X1 U1928 ( .A(n1289), .Z(n4) );
  BUF_X1 U1929 ( .A(n1272), .Z(n48) );
  BUF_X1 U1930 ( .A(n1274), .Z(n36) );
  BUF_X1 U1931 ( .A(n1271), .Z(n54) );
  INV_X1 U1932 ( .A(n49), .ZN(n1291) );
  INV_X1 U1933 ( .A(n25), .ZN(n1295) );
  INV_X1 U1934 ( .A(n43), .ZN(n1292) );
  INV_X1 U1935 ( .A(n37), .ZN(n1293) );
  INV_X1 U1936 ( .A(n55), .ZN(n1290) );
  INV_X1 U1937 ( .A(n1467), .ZN(n1297) );
  INV_X1 U1938 ( .A(n1471), .ZN(n1296) );
  BUF_X1 U1939 ( .A(n1279), .Z(n5) );
  XNOR2_X1 U1940 ( .A(a[15]), .B(a[16]), .ZN(n1281) );
  XNOR2_X1 U1941 ( .A(a[10]), .B(a[9]), .ZN(n1284) );
  XNOR2_X1 U1942 ( .A(a[2]), .B(a[1]), .ZN(n1288) );
  XNOR2_X1 U1943 ( .A(a[17]), .B(a[18]), .ZN(n1280) );
  NAND2_X1 U1944 ( .A1(n1268), .A2(n1288), .ZN(n1278) );
  AOI21_X1 U1945 ( .B1(n367), .B2(n359), .A(n360), .ZN(n358) );
  NAND2_X1 U1946 ( .A1(n1265), .A2(n1285), .ZN(n1275) );
  XNOR2_X1 U1947 ( .A(a[8]), .B(a[7]), .ZN(n1285) );
  NOR2_X1 U1948 ( .A1(n1409), .A2(n326), .ZN(n321) );
  OAI21_X1 U1949 ( .B1(n327), .B2(n323), .A(n324), .ZN(n322) );
  XNOR2_X1 U1950 ( .A(n385), .B(n97), .ZN(product[8]) );
  XNOR2_X1 U1951 ( .A(n1467), .B(n1487), .ZN(n1188) );
  XNOR2_X1 U1952 ( .A(n1467), .B(n1250), .ZN(n1187) );
  XNOR2_X1 U1953 ( .A(n1467), .B(n1486), .ZN(n1194) );
  XNOR2_X1 U1954 ( .A(n1467), .B(n1253), .ZN(n1190) );
  XNOR2_X1 U1955 ( .A(n1467), .B(n1494), .ZN(n1196) );
  XNOR2_X1 U1956 ( .A(n1467), .B(n1252), .ZN(n1189) );
  XNOR2_X1 U1957 ( .A(n1467), .B(n1488), .ZN(n1193) );
  XNOR2_X1 U1958 ( .A(n1467), .B(n1258), .ZN(n1195) );
  XNOR2_X1 U1959 ( .A(n1467), .B(n1244), .ZN(n1181) );
  XNOR2_X1 U1960 ( .A(n13), .B(n1246), .ZN(n1183) );
  XNOR2_X1 U1961 ( .A(n13), .B(n1245), .ZN(n1182) );
  XNOR2_X1 U1962 ( .A(n1467), .B(n1255), .ZN(n1192) );
  XNOR2_X1 U1963 ( .A(n1467), .B(n1254), .ZN(n1191) );
  XNOR2_X1 U1964 ( .A(n1467), .B(n1249), .ZN(n1186) );
  XNOR2_X1 U1965 ( .A(n13), .B(n1243), .ZN(n1180) );
  XNOR2_X1 U1966 ( .A(n1242), .B(n13), .ZN(n1179) );
  XNOR2_X1 U1967 ( .A(n13), .B(n1241), .ZN(n1178) );
  XNOR2_X1 U1968 ( .A(n1467), .B(n1248), .ZN(n1185) );
  XNOR2_X1 U1969 ( .A(n13), .B(n1247), .ZN(n1184) );
  XNOR2_X1 U1970 ( .A(n1467), .B(n1484), .ZN(n1177) );
  NOR2_X1 U1971 ( .A1(n247), .A2(n117), .ZN(n115) );
  NOR2_X1 U1972 ( .A1(n247), .A2(n108), .ZN(n106) );
  NOR2_X1 U1973 ( .A1(n247), .A2(n201), .ZN(n199) );
  NOR2_X1 U1974 ( .A1(n247), .A2(n130), .ZN(n128) );
  NOR2_X1 U1975 ( .A1(n247), .A2(n171), .ZN(n169) );
  NOR2_X1 U1976 ( .A1(n247), .A2(n160), .ZN(n158) );
  NOR2_X1 U1977 ( .A1(n247), .A2(n145), .ZN(n143) );
  NOR2_X1 U1978 ( .A1(n247), .A2(n242), .ZN(n232) );
  NOR2_X1 U1979 ( .A1(n247), .A2(n184), .ZN(n182) );
  NOR2_X1 U1980 ( .A1(n247), .A2(n216), .ZN(n210) );
  NOR2_X1 U1981 ( .A1(n247), .A2(n225), .ZN(n223) );
  AOI21_X1 U1982 ( .B1(n349), .B2(n1437), .A(n344), .ZN(n342) );
  XNOR2_X1 U1983 ( .A(n1469), .B(n1243), .ZN(n1096) );
  XNOR2_X1 U1984 ( .A(n1469), .B(n1242), .ZN(n1095) );
  XNOR2_X1 U1985 ( .A(n1469), .B(n1245), .ZN(n1098) );
  XNOR2_X1 U1986 ( .A(n1469), .B(n1249), .ZN(n1102) );
  XNOR2_X1 U1987 ( .A(n1469), .B(n1244), .ZN(n1097) );
  XNOR2_X1 U1988 ( .A(n1469), .B(n1253), .ZN(n1106) );
  XNOR2_X1 U1989 ( .A(n1469), .B(n1248), .ZN(n1101) );
  XNOR2_X1 U1990 ( .A(n1469), .B(n1254), .ZN(n1107) );
  XNOR2_X1 U1991 ( .A(n1469), .B(n1252), .ZN(n1105) );
  XNOR2_X1 U1992 ( .A(n1469), .B(n1494), .ZN(n1112) );
  XNOR2_X1 U1993 ( .A(n1469), .B(n1247), .ZN(n1100) );
  XNOR2_X1 U1994 ( .A(n37), .B(n1246), .ZN(n1099) );
  XNOR2_X1 U1995 ( .A(n1469), .B(n1258), .ZN(n1111) );
  XNOR2_X1 U1996 ( .A(n37), .B(n1255), .ZN(n1108) );
  XNOR2_X1 U1997 ( .A(n37), .B(n1257), .ZN(n1110) );
  XNOR2_X1 U1998 ( .A(n1469), .B(n1251), .ZN(n1104) );
  XNOR2_X1 U1999 ( .A(n37), .B(n1256), .ZN(n1109) );
  XNOR2_X1 U2000 ( .A(n37), .B(n1489), .ZN(n1103) );
  XNOR2_X1 U2001 ( .A(n1469), .B(n1241), .ZN(n1094) );
  XNOR2_X1 U2002 ( .A(n1469), .B(n1458), .ZN(n1093) );
  OAI21_X1 U2003 ( .B1(n1476), .B2(n304), .A(n297), .ZN(n295) );
  XNOR2_X1 U2004 ( .A(n1406), .B(n1458), .ZN(n1030) );
  XNOR2_X1 U2005 ( .A(n1406), .B(n1241), .ZN(n1031) );
  XNOR2_X1 U2006 ( .A(n1406), .B(n1242), .ZN(n1032) );
  XNOR2_X1 U2007 ( .A(n1406), .B(n1243), .ZN(n1033) );
  XNOR2_X1 U2008 ( .A(n55), .B(n1249), .ZN(n1039) );
  XNOR2_X1 U2009 ( .A(n1406), .B(n1245), .ZN(n1035) );
  XNOR2_X1 U2010 ( .A(n1406), .B(n1244), .ZN(n1034) );
  XNOR2_X1 U2011 ( .A(n55), .B(n1248), .ZN(n1038) );
  XNOR2_X1 U2012 ( .A(n55), .B(n1250), .ZN(n1040) );
  XNOR2_X1 U2013 ( .A(n55), .B(n1247), .ZN(n1037) );
  XNOR2_X1 U2014 ( .A(n1406), .B(n1246), .ZN(n1036) );
  XNOR2_X1 U2015 ( .A(n55), .B(n1494), .ZN(n1049) );
  XNOR2_X1 U2016 ( .A(n55), .B(n1254), .ZN(n1044) );
  XNOR2_X1 U2017 ( .A(n55), .B(n1253), .ZN(n1043) );
  XNOR2_X1 U2018 ( .A(n55), .B(n1252), .ZN(n1042) );
  XNOR2_X1 U2019 ( .A(n55), .B(n1487), .ZN(n1041) );
  XNOR2_X1 U2020 ( .A(n55), .B(n1255), .ZN(n1045) );
  XNOR2_X1 U2021 ( .A(n55), .B(n1256), .ZN(n1046) );
  XNOR2_X1 U2022 ( .A(n55), .B(n1258), .ZN(n1048) );
  XNOR2_X1 U2023 ( .A(n55), .B(n1257), .ZN(n1047) );
  NAND2_X1 U2024 ( .A1(n1397), .A2(n384), .ZN(n97) );
  XNOR2_X1 U2025 ( .A(n1470), .B(n1248), .ZN(n1164) );
  XNOR2_X1 U2026 ( .A(n1470), .B(n1254), .ZN(n1170) );
  XNOR2_X1 U2027 ( .A(n1471), .B(n1494), .ZN(n1175) );
  XNOR2_X1 U2028 ( .A(n1470), .B(n1258), .ZN(n1174) );
  XNOR2_X1 U2029 ( .A(n1471), .B(n1242), .ZN(n1158) );
  XNOR2_X1 U2030 ( .A(n1471), .B(n1253), .ZN(n1169) );
  XNOR2_X1 U2031 ( .A(n1470), .B(n1252), .ZN(n1168) );
  XNOR2_X1 U2032 ( .A(n1470), .B(n1243), .ZN(n1159) );
  XNOR2_X1 U2033 ( .A(n1471), .B(n1486), .ZN(n1173) );
  XNOR2_X1 U2034 ( .A(n1470), .B(n1245), .ZN(n1161) );
  XNOR2_X1 U2035 ( .A(n1470), .B(n1244), .ZN(n1160) );
  XNOR2_X1 U2036 ( .A(n1471), .B(n1247), .ZN(n1163) );
  XNOR2_X1 U2037 ( .A(n1470), .B(n1246), .ZN(n1162) );
  XNOR2_X1 U2038 ( .A(n1471), .B(n1249), .ZN(n1165) );
  XNOR2_X1 U2039 ( .A(n1471), .B(n1241), .ZN(n1157) );
  XNOR2_X1 U2040 ( .A(n1471), .B(n1487), .ZN(n1167) );
  XNOR2_X1 U2041 ( .A(n1471), .B(n1488), .ZN(n1172) );
  XNOR2_X1 U2042 ( .A(n1471), .B(n1489), .ZN(n1166) );
  XNOR2_X1 U2043 ( .A(n1471), .B(n1255), .ZN(n1171) );
  XNOR2_X1 U2044 ( .A(n1471), .B(n1240), .ZN(n1156) );
  INV_X1 U2045 ( .A(n338), .ZN(n336) );
  INV_X1 U2046 ( .A(n1454), .ZN(n319) );
  XNOR2_X1 U2047 ( .A(n1415), .B(n1245), .ZN(n1077) );
  XNOR2_X1 U2048 ( .A(n1414), .B(n1244), .ZN(n1076) );
  XNOR2_X1 U2049 ( .A(n1414), .B(n1242), .ZN(n1074) );
  XNOR2_X1 U2050 ( .A(n1415), .B(n1243), .ZN(n1075) );
  XNOR2_X1 U2051 ( .A(n1414), .B(n1247), .ZN(n1079) );
  XNOR2_X1 U2052 ( .A(n1415), .B(n1246), .ZN(n1078) );
  XNOR2_X1 U2053 ( .A(n1414), .B(n1241), .ZN(n1073) );
  XNOR2_X1 U2054 ( .A(n1415), .B(n1494), .ZN(n1091) );
  XNOR2_X1 U2055 ( .A(n1415), .B(n1458), .ZN(n1072) );
  XNOR2_X1 U2056 ( .A(n1415), .B(n1250), .ZN(n1082) );
  XNOR2_X1 U2057 ( .A(n1414), .B(n1251), .ZN(n1083) );
  XNOR2_X1 U2058 ( .A(n1415), .B(n1249), .ZN(n1081) );
  XNOR2_X1 U2059 ( .A(n1413), .B(n1248), .ZN(n1080) );
  XNOR2_X1 U2060 ( .A(n43), .B(n1488), .ZN(n1088) );
  XNOR2_X1 U2061 ( .A(n1414), .B(n1253), .ZN(n1085) );
  XNOR2_X1 U2062 ( .A(n1414), .B(n1252), .ZN(n1084) );
  XNOR2_X1 U2063 ( .A(n43), .B(n1255), .ZN(n1087) );
  XNOR2_X1 U2064 ( .A(n43), .B(n1254), .ZN(n1086) );
  XNOR2_X1 U2065 ( .A(n43), .B(n1258), .ZN(n1090) );
  XNOR2_X1 U2066 ( .A(n43), .B(n1257), .ZN(n1089) );
  AOI21_X1 U2067 ( .B1(n357), .B2(n348), .A(n349), .ZN(n347) );
  AOI21_X1 U2068 ( .B1(n340), .B2(n321), .A(n322), .ZN(n320) );
  NAND2_X1 U2069 ( .A1(n348), .A2(n1437), .ZN(n341) );
  NAND2_X1 U2070 ( .A1(n767), .A2(n772), .ZN(n384) );
  XNOR2_X1 U2071 ( .A(n25), .B(n1244), .ZN(n1139) );
  XNOR2_X1 U2072 ( .A(n25), .B(n1254), .ZN(n1149) );
  XNOR2_X1 U2073 ( .A(n25), .B(n1246), .ZN(n1141) );
  XNOR2_X1 U2074 ( .A(n25), .B(n1250), .ZN(n1145) );
  XNOR2_X1 U2075 ( .A(n25), .B(n1245), .ZN(n1140) );
  XNOR2_X1 U2076 ( .A(n25), .B(n1494), .ZN(n1154) );
  XNOR2_X1 U2077 ( .A(n25), .B(n1243), .ZN(n1138) );
  XNOR2_X1 U2078 ( .A(n25), .B(n1247), .ZN(n1142) );
  XNOR2_X1 U2079 ( .A(n25), .B(n1484), .ZN(n1135) );
  XNOR2_X1 U2080 ( .A(n25), .B(n1255), .ZN(n1150) );
  XNOR2_X1 U2081 ( .A(n25), .B(n1486), .ZN(n1152) );
  XNOR2_X1 U2082 ( .A(n25), .B(n1258), .ZN(n1153) );
  XNOR2_X1 U2083 ( .A(n25), .B(n1256), .ZN(n1151) );
  XNOR2_X1 U2084 ( .A(n25), .B(n1242), .ZN(n1137) );
  XNOR2_X1 U2085 ( .A(n25), .B(n1253), .ZN(n1148) );
  XNOR2_X1 U2086 ( .A(n25), .B(n1249), .ZN(n1144) );
  XNOR2_X1 U2087 ( .A(n25), .B(n1248), .ZN(n1143) );
  XNOR2_X1 U2088 ( .A(n25), .B(n1241), .ZN(n1136) );
  XNOR2_X1 U2089 ( .A(n25), .B(n1252), .ZN(n1147) );
  XNOR2_X1 U2090 ( .A(n25), .B(n1251), .ZN(n1146) );
  XNOR2_X1 U2091 ( .A(n1456), .B(n1458), .ZN(n1051) );
  XNOR2_X1 U2092 ( .A(n1456), .B(n1247), .ZN(n1058) );
  XNOR2_X1 U2093 ( .A(n1456), .B(n1243), .ZN(n1054) );
  XNOR2_X1 U2094 ( .A(n49), .B(n1246), .ZN(n1057) );
  XNOR2_X1 U2095 ( .A(n1456), .B(n1242), .ZN(n1053) );
  XNOR2_X1 U2096 ( .A(n49), .B(n1245), .ZN(n1056) );
  XNOR2_X1 U2097 ( .A(n1456), .B(n1241), .ZN(n1052) );
  XNOR2_X1 U2098 ( .A(n1456), .B(n1244), .ZN(n1055) );
  XNOR2_X1 U2099 ( .A(n49), .B(n1248), .ZN(n1059) );
  XNOR2_X1 U2100 ( .A(n49), .B(n1253), .ZN(n1064) );
  XNOR2_X1 U2101 ( .A(n49), .B(n1252), .ZN(n1063) );
  XNOR2_X1 U2102 ( .A(n49), .B(n1487), .ZN(n1062) );
  XNOR2_X1 U2103 ( .A(n49), .B(n1494), .ZN(n1070) );
  XNOR2_X1 U2104 ( .A(n49), .B(n1489), .ZN(n1061) );
  XNOR2_X1 U2105 ( .A(n49), .B(n1255), .ZN(n1066) );
  XNOR2_X1 U2106 ( .A(n49), .B(n1254), .ZN(n1065) );
  XNOR2_X1 U2107 ( .A(n49), .B(n1258), .ZN(n1069) );
  XNOR2_X1 U2108 ( .A(n49), .B(n1249), .ZN(n1060) );
  XNOR2_X1 U2109 ( .A(n49), .B(n1257), .ZN(n1068) );
  XNOR2_X1 U2110 ( .A(n49), .B(n1256), .ZN(n1067) );
  AOI21_X1 U2111 ( .B1(n319), .B2(n315), .A(n316), .ZN(n314) );
  XNOR2_X1 U2112 ( .A(n319), .B(n86), .ZN(product[19]) );
  AOI21_X1 U2113 ( .B1(n299), .B2(n319), .A(n300), .ZN(n298) );
  AOI21_X1 U2114 ( .B1(n319), .B2(n306), .A(n1447), .ZN(n305) );
  NOR2_X1 U2115 ( .A1(n350), .A2(n355), .ZN(n348) );
  OAI21_X1 U2116 ( .B1(n350), .B2(n356), .A(n351), .ZN(n349) );
  AOI21_X1 U2117 ( .B1(n1491), .B2(n210), .A(n211), .ZN(n209) );
  AOI21_X1 U2118 ( .B1(n63), .B2(n199), .A(n200), .ZN(n198) );
  OAI21_X1 U2119 ( .B1(n217), .B2(n121), .A(n122), .ZN(n120) );
  OAI21_X1 U2120 ( .B1(n217), .B2(n192), .A(n193), .ZN(n187) );
  OAI21_X1 U2121 ( .B1(n1457), .B2(n318), .A(n313), .ZN(n311) );
  NOR2_X1 U2122 ( .A1(n312), .A2(n317), .ZN(n310) );
  INV_X1 U2123 ( .A(n312), .ZN(n428) );
  OAI21_X1 U2124 ( .B1(n1462), .B2(n108), .A(n109), .ZN(n107) );
  OAI21_X1 U2125 ( .B1(n1462), .B2(n117), .A(n118), .ZN(n116) );
  OAI21_X1 U2126 ( .B1(n1416), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U2127 ( .B1(n1416), .B2(n145), .A(n146), .ZN(n144) );
  OAI21_X1 U2128 ( .B1(n65), .B2(n216), .A(n217), .ZN(n211) );
  OAI21_X1 U2129 ( .B1(n1448), .B2(n184), .A(n185), .ZN(n183) );
  OAI21_X1 U2130 ( .B1(n1448), .B2(n171), .A(n172), .ZN(n170) );
  OAI21_X1 U2131 ( .B1(n242), .B2(n65), .A(n243), .ZN(n233) );
  OAI21_X1 U2132 ( .B1(n1448), .B2(n160), .A(n161), .ZN(n159) );
  OAI21_X1 U2133 ( .B1(n1448), .B2(n201), .A(n202), .ZN(n200) );
  OAI21_X1 U2134 ( .B1(n65), .B2(n225), .A(n226), .ZN(n224) );
  NAND2_X1 U2135 ( .A1(n1260), .A2(n1280), .ZN(n1270) );
  XNOR2_X1 U2136 ( .A(n101), .B(n401), .ZN(product[4]) );
  AOI21_X1 U2137 ( .B1(n1399), .B2(n401), .A(n398), .ZN(n396) );
  XNOR2_X1 U2138 ( .A(n1444), .B(n1246), .ZN(n1225) );
  XNOR2_X1 U2139 ( .A(n1444), .B(n1251), .ZN(n1230) );
  XNOR2_X1 U2140 ( .A(n1444), .B(n1252), .ZN(n1231) );
  XNOR2_X1 U2141 ( .A(n1), .B(n1245), .ZN(n1224) );
  XNOR2_X1 U2142 ( .A(n1444), .B(n1247), .ZN(n1226) );
  XNOR2_X1 U2143 ( .A(n1444), .B(n1248), .ZN(n1227) );
  XNOR2_X1 U2144 ( .A(n1), .B(n1244), .ZN(n1223) );
  XNOR2_X1 U2145 ( .A(n1), .B(n1243), .ZN(n1222) );
  XNOR2_X1 U2146 ( .A(n1444), .B(n1242), .ZN(n1221) );
  XNOR2_X1 U2147 ( .A(n1), .B(n1241), .ZN(n1220) );
  XNOR2_X1 U2148 ( .A(n1444), .B(n1254), .ZN(n1233) );
  XNOR2_X1 U2149 ( .A(n1444), .B(n1253), .ZN(n1232) );
  XNOR2_X1 U2150 ( .A(n1444), .B(n1250), .ZN(n1229) );
  XNOR2_X1 U2151 ( .A(n1444), .B(n1255), .ZN(n1234) );
  XNOR2_X1 U2152 ( .A(n1444), .B(n1256), .ZN(n1235) );
  XNOR2_X1 U2153 ( .A(n1444), .B(n1249), .ZN(n1228) );
  XNOR2_X1 U2154 ( .A(n1444), .B(n1494), .ZN(n1238) );
  XNOR2_X1 U2155 ( .A(n1), .B(n1240), .ZN(n1219) );
  XNOR2_X1 U2156 ( .A(n1444), .B(n1258), .ZN(n1237) );
  XNOR2_X1 U2157 ( .A(n1444), .B(n1486), .ZN(n1236) );
  XOR2_X1 U2158 ( .A(n388), .B(n98), .Z(product[7]) );
  XOR2_X1 U2159 ( .A(a[18]), .B(a[19]), .Z(n1260) );
  AOI21_X1 U2160 ( .B1(n64), .B2(n182), .A(n183), .ZN(n181) );
  XNOR2_X1 U2161 ( .A(n99), .B(n393), .ZN(product[6]) );
  XOR2_X1 U2162 ( .A(a[4]), .B(a[5]), .Z(n1267) );
  XNOR2_X1 U2163 ( .A(a[6]), .B(a[5]), .ZN(n1286) );
  XOR2_X1 U2164 ( .A(a[7]), .B(a[6]), .Z(n1266) );
  NOR2_X1 U2165 ( .A1(n361), .A2(n364), .ZN(n359) );
  OAI21_X1 U2166 ( .B1(n361), .B2(n365), .A(n362), .ZN(n360) );
  XNOR2_X1 U2167 ( .A(a[11]), .B(a[12]), .ZN(n1283) );
  XOR2_X1 U2168 ( .A(a[11]), .B(a[10]), .Z(n1264) );
  NAND2_X1 U2169 ( .A1(n1263), .A2(n1283), .ZN(n1273) );
  XOR2_X1 U2170 ( .A(a[15]), .B(a[14]), .Z(n1262) );
  XNOR2_X1 U2171 ( .A(a[3]), .B(a[4]), .ZN(n1287) );
  XOR2_X1 U2172 ( .A(a[2]), .B(a[3]), .Z(n1268) );
  AOI21_X1 U2173 ( .B1(n64), .B2(n169), .A(n170), .ZN(n168) );
  XNOR2_X1 U2174 ( .A(a[13]), .B(a[14]), .ZN(n1282) );
  XOR2_X1 U2175 ( .A(a[12]), .B(a[13]), .Z(n1263) );
  NAND2_X1 U2176 ( .A1(n134), .A2(n1394), .ZN(n121) );
  AOI21_X1 U2177 ( .B1(n63), .B2(n232), .A(n233), .ZN(n231) );
  AOI21_X1 U2178 ( .B1(n1492), .B2(n223), .A(n224), .ZN(n222) );
  AOI21_X1 U2179 ( .B1(n1492), .B2(n245), .A(n246), .ZN(n244) );
  XNOR2_X1 U2180 ( .A(n1492), .B(n82), .ZN(product[23]) );
  AOI21_X1 U2181 ( .B1(n1491), .B2(n258), .A(n259), .ZN(n257) );
  AOI21_X1 U2182 ( .B1(n63), .B2(n269), .A(n270), .ZN(n268) );
  AOI21_X1 U2183 ( .B1(n64), .B2(n425), .A(n288), .ZN(n286) );
  NOR2_X1 U2184 ( .A1(n289), .A2(n284), .ZN(n282) );
  INV_X1 U2185 ( .A(n394), .ZN(n443) );
  NOR2_X1 U2186 ( .A1(n783), .A2(n786), .ZN(n394) );
  XOR2_X1 U2187 ( .A(a[8]), .B(a[9]), .Z(n1265) );
  NAND2_X1 U2188 ( .A1(n789), .A2(n828), .ZN(n403) );
  OAI21_X1 U2189 ( .B1(n292), .B2(n320), .A(n293), .ZN(n291) );
  XOR2_X1 U2190 ( .A(a[16]), .B(a[17]), .Z(n1261) );
  XOR2_X1 U2191 ( .A(a[0]), .B(a[1]), .Z(n1269) );
  OAI22_X1 U2192 ( .A1(n5), .A2(n1299), .B1(n1239), .B2(n4), .ZN(n829) );
  OR2_X1 U2193 ( .A1(n1495), .A2(n1299), .ZN(n1239) );
  AOI21_X1 U2194 ( .B1(n1491), .B2(n282), .A(n279), .ZN(n277) );
endmodule


module datapath_DW_mult_tc_15 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n3, n4, n5, n6, n7, n9, n10, n12, n13, n15, n16, n17, n18, n19,
         n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34, n35, n36,
         n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n51, n52, n53,
         n54, n57, n58, n59, n60, n61, n63, n64, n65, n66, n67, n68, n69, n70,
         n72, n82, n83, n84, n85, n86, n87, n88, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n105, n106, n107, n108,
         n109, n111, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n124, n126, n127, n128, n129, n130, n131, n134, n135, n136,
         n137, n139, n141, n142, n143, n144, n145, n146, n149, n150, n151,
         n152, n154, n156, n157, n158, n159, n160, n161, n165, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n190, n191, n192,
         n193, n195, n197, n198, n199, n200, n201, n202, n206, n208, n209,
         n210, n211, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n254, n256, n257, n258, n259, n260, n261, n262, n263,
         n265, n267, n268, n269, n270, n273, n274, n275, n276, n277, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n329, n331, n332, n333, n334, n336, n338, n339,
         n340, n341, n342, n344, n346, n347, n348, n349, n350, n351, n352,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n376,
         n378, n379, n380, n382, n384, n385, n386, n387, n388, n390, n392,
         n393, n394, n395, n396, n398, n400, n401, n402, n403, n404, n405,
         n406, n407, n409, n418, n424, n426, n428, n430, n434, n435, n436,
         n437, n438, n441, n443, n445, n446, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n793, n794,
         n796, n797, n799, n800, n802, n803, n805, n806, n808, n809, n811,
         n812, n814, n815, n817, n818, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1480, n1481;
  assign product[39] = n105;

  FA_X1 U488 ( .A(n831), .B(n454), .CI(n850), .CO(n450), .S(n451) );
  FA_X1 U489 ( .A(n455), .B(n832), .CI(n458), .CO(n452), .S(n453) );
  FA_X1 U491 ( .A(n462), .B(n833), .CI(n459), .CO(n456), .S(n457) );
  FA_X1 U492 ( .A(n851), .B(n464), .CI(n870), .CO(n458), .S(n459) );
  FA_X1 U493 ( .A(n463), .B(n470), .CI(n468), .CO(n460), .S(n461) );
  FA_X1 U494 ( .A(n834), .B(n852), .CI(n465), .CO(n462), .S(n463) );
  FA_X1 U496 ( .A(n474), .B(n471), .CI(n469), .CO(n466), .S(n467) );
  FA_X1 U497 ( .A(n478), .B(n871), .CI(n476), .CO(n468), .S(n469) );
  FA_X1 U498 ( .A(n853), .B(n835), .CI(n890), .CO(n470), .S(n471) );
  FA_X1 U499 ( .A(n475), .B(n477), .CI(n482), .CO(n472), .S(n473) );
  FA_X1 U500 ( .A(n486), .B(n479), .CI(n484), .CO(n474), .S(n475) );
  FA_X1 U501 ( .A(n836), .B(n854), .CI(n872), .CO(n476), .S(n477) );
  FA_X1 U503 ( .A(n490), .B(n492), .CI(n483), .CO(n480), .S(n481) );
  FA_X1 U504 ( .A(n485), .B(n494), .CI(n487), .CO(n482), .S(n483) );
  FA_X1 U505 ( .A(n855), .B(n496), .CI(n873), .CO(n484), .S(n485) );
  FA_X1 U506 ( .A(n891), .B(n837), .CI(n910), .CO(n486), .S(n487) );
  FA_X1 U507 ( .A(n500), .B(n493), .CI(n491), .CO(n488), .S(n489) );
  FA_X1 U508 ( .A(n495), .B(n504), .CI(n502), .CO(n490), .S(n491) );
  FA_X1 U509 ( .A(n497), .B(n874), .CI(n506), .CO(n492), .S(n493) );
  FA_X1 U510 ( .A(n892), .B(n856), .CI(n838), .CO(n494), .S(n495) );
  FA_X1 U512 ( .A(n510), .B(n503), .CI(n501), .CO(n498), .S(n499) );
  FA_X1 U513 ( .A(n507), .B(n505), .CI(n512), .CO(n500), .S(n501) );
  FA_X1 U514 ( .A(n516), .B(n893), .CI(n514), .CO(n502), .S(n503) );
  FA_X1 U515 ( .A(n857), .B(n911), .CI(n875), .CO(n504), .S(n505) );
  FA_X1 U516 ( .A(n518), .B(n839), .CI(n930), .CO(n506), .S(n507) );
  FA_X1 U517 ( .A(n522), .B(n513), .CI(n511), .CO(n508), .S(n509) );
  FA_X1 U518 ( .A(n526), .B(n515), .CI(n524), .CO(n510), .S(n511) );
  FA_X1 U519 ( .A(n528), .B(n530), .CI(n517), .CO(n512), .S(n513) );
  FA_X1 U520 ( .A(n840), .B(n858), .CI(n519), .CO(n514), .S(n515) );
  FA_X1 U521 ( .A(n912), .B(n876), .CI(n894), .CO(n516), .S(n517) );
  FA_X1 U523 ( .A(n525), .B(n534), .CI(n523), .CO(n520), .S(n521) );
  FA_X1 U524 ( .A(n527), .B(n538), .CI(n536), .CO(n522), .S(n523) );
  FA_X1 U525 ( .A(n529), .B(n540), .CI(n531), .CO(n524), .S(n525) );
  FA_X1 U526 ( .A(n877), .B(n895), .CI(n542), .CO(n526), .S(n527) );
  FA_X1 U527 ( .A(n859), .B(n931), .CI(n913), .CO(n528), .S(n529) );
  FA_X1 U528 ( .A(n544), .B(n841), .CI(n950), .CO(n530), .S(n531) );
  FA_X1 U529 ( .A(n535), .B(n537), .CI(n548), .CO(n532), .S(n533) );
  FA_X1 U530 ( .A(n539), .B(n552), .CI(n550), .CO(n534), .S(n535) );
  FA_X1 U531 ( .A(n541), .B(n554), .CI(n543), .CO(n536), .S(n537) );
  FA_X1 U532 ( .A(n558), .B(n545), .CI(n556), .CO(n538), .S(n539) );
  FA_X1 U533 ( .A(n896), .B(n932), .CI(n914), .CO(n540), .S(n541) );
  FA_X1 U534 ( .A(n842), .B(n878), .CI(n860), .CO(n542), .S(n543) );
  FA_X1 U536 ( .A(n562), .B(n551), .CI(n549), .CO(n546), .S(n547) );
  FA_X1 U537 ( .A(n553), .B(n566), .CI(n564), .CO(n548), .S(n549) );
  FA_X1 U538 ( .A(n559), .B(n557), .CI(n568), .CO(n550), .S(n551) );
  FA_X1 U539 ( .A(n570), .B(n572), .CI(n555), .CO(n552), .S(n553) );
  FA_X1 U540 ( .A(n879), .B(n915), .CI(n897), .CO(n554), .S(n555) );
  FA_X1 U541 ( .A(n861), .B(n951), .CI(n933), .CO(n556), .S(n557) );
  FA_X1 U542 ( .A(n574), .B(n843), .CI(n970), .CO(n558), .S(n559) );
  FA_X1 U543 ( .A(n578), .B(n565), .CI(n563), .CO(n560), .S(n561) );
  FA_X1 U544 ( .A(n567), .B(n582), .CI(n580), .CO(n562), .S(n563) );
  FA_X1 U545 ( .A(n584), .B(n573), .CI(n569), .CO(n564), .S(n565) );
  FA_X1 U546 ( .A(n586), .B(n588), .CI(n571), .CO(n566), .S(n567) );
  FA_X1 U547 ( .A(n575), .B(n898), .CI(n590), .CO(n568), .S(n569) );
  FA_X1 U548 ( .A(n844), .B(n916), .CI(n862), .CO(n570), .S(n571) );
  FA_X1 U549 ( .A(n952), .B(n880), .CI(n934), .CO(n572), .S(n573) );
  FA_X1 U551 ( .A(n594), .B(n581), .CI(n579), .CO(n576), .S(n577) );
  FA_X1 U552 ( .A(n583), .B(n598), .CI(n596), .CO(n578), .S(n579) );
  FA_X1 U553 ( .A(n600), .B(n591), .CI(n585), .CO(n580), .S(n581) );
  FA_X1 U554 ( .A(n587), .B(n602), .CI(n589), .CO(n582), .S(n583) );
  FA_X1 U555 ( .A(n606), .B(n917), .CI(n604), .CO(n584), .S(n585) );
  FA_X1 U556 ( .A(n881), .B(n935), .CI(n899), .CO(n586), .S(n587) );
  FA_X1 U557 ( .A(n608), .B(n953), .CI(n863), .CO(n588), .S(n589) );
  FA_X1 U558 ( .A(n971), .B(n845), .CI(n990), .CO(n590), .S(n591) );
  FA_X1 U559 ( .A(n612), .B(n597), .CI(n595), .CO(n592), .S(n593) );
  FA_X1 U560 ( .A(n599), .B(n616), .CI(n614), .CO(n594), .S(n595) );
  FA_X1 U561 ( .A(n618), .B(n603), .CI(n601), .CO(n596), .S(n597) );
  FA_X1 U562 ( .A(n605), .B(n620), .CI(n607), .CO(n598), .S(n599) );
  FA_X1 U563 ( .A(n626), .B(n624), .CI(n622), .CO(n600), .S(n601) );
  FA_X1 U564 ( .A(n918), .B(n936), .CI(n609), .CO(n602), .S(n603) );
  FA_X1 U565 ( .A(n882), .B(n864), .CI(n954), .CO(n604), .S(n605) );
  FA_X1 U569 ( .A(n617), .B(n634), .CI(n632), .CO(n612), .S(n613) );
  FA_X1 U570 ( .A(n636), .B(n621), .CI(n619), .CO(n614), .S(n615) );
  FA_X1 U571 ( .A(n623), .B(n638), .CI(n625), .CO(n616), .S(n617) );
  FA_X1 U572 ( .A(n627), .B(n642), .CI(n640), .CO(n618), .S(n619) );
  FA_X1 U573 ( .A(n955), .B(n973), .CI(n644), .CO(n620), .S(n621) );
  FA_X1 U574 ( .A(n991), .B(n901), .CI(n883), .CO(n622), .S(n623) );
  FA_X1 U575 ( .A(n919), .B(n847), .CI(n1010), .CO(n624), .S(n625) );
  FA_X1 U578 ( .A(n648), .B(n633), .CI(n631), .CO(n628), .S(n629) );
  FA_X1 U579 ( .A(n635), .B(n637), .CI(n650), .CO(n630), .S(n631) );
  FA_X1 U580 ( .A(n654), .B(n643), .CI(n652), .CO(n632), .S(n633) );
  FA_X1 U581 ( .A(n639), .B(n656), .CI(n641), .CO(n634), .S(n635) );
  FA_X1 U582 ( .A(n660), .B(n645), .CI(n658), .CO(n636), .S(n637) );
  FA_X1 U583 ( .A(n920), .B(n992), .CI(n974), .CO(n638), .S(n639) );
  FA_X1 U584 ( .A(n1011), .B(n956), .CI(n902), .CO(n640), .S(n641) );
  FA_X1 U585 ( .A(n866), .B(n884), .CI(n938), .CO(n642), .S(n643) );
  HA_X1 U586 ( .A(n820), .B(n848), .CO(n644), .S(n645) );
  FA_X1 U587 ( .A(n664), .B(n651), .CI(n649), .CO(n646), .S(n647) );
  FA_X1 U588 ( .A(n666), .B(n655), .CI(n653), .CO(n648), .S(n649) );
  FA_X1 U589 ( .A(n670), .B(n659), .CI(n668), .CO(n650), .S(n651) );
  FA_X1 U590 ( .A(n661), .B(n672), .CI(n657), .CO(n652), .S(n653) );
  FA_X1 U591 ( .A(n676), .B(n957), .CI(n674), .CO(n654), .S(n655) );
  FA_X1 U592 ( .A(n921), .B(n975), .CI(n939), .CO(n656), .S(n657) );
  FA_X1 U593 ( .A(n867), .B(n993), .CI(n903), .CO(n658), .S(n659) );
  FA_X1 U594 ( .A(n849), .B(n885), .CI(n1012), .CO(n660), .S(n661) );
  FA_X1 U595 ( .A(n667), .B(n680), .CI(n665), .CO(n662), .S(n663) );
  FA_X1 U596 ( .A(n682), .B(n671), .CI(n669), .CO(n664), .S(n665) );
  FA_X1 U597 ( .A(n675), .B(n673), .CI(n684), .CO(n666), .S(n667) );
  FA_X1 U598 ( .A(n686), .B(n690), .CI(n688), .CO(n668), .S(n669) );
  FA_X1 U599 ( .A(n958), .B(n976), .CI(n677), .CO(n670), .S(n671) );
  FA_X1 U600 ( .A(n886), .B(n904), .CI(n922), .CO(n672), .S(n673) );
  FA_X1 U601 ( .A(n1013), .B(n940), .CI(n994), .CO(n674), .S(n675) );
  HA_X1 U602 ( .A(n821), .B(n868), .CO(n676), .S(n677) );
  FA_X1 U603 ( .A(n694), .B(n683), .CI(n681), .CO(n678), .S(n679) );
  FA_X1 U604 ( .A(n685), .B(n698), .CI(n696), .CO(n680), .S(n681) );
  FA_X1 U605 ( .A(n689), .B(n691), .CI(n687), .CO(n682), .S(n683) );
  FA_X1 U606 ( .A(n702), .B(n704), .CI(n700), .CO(n684), .S(n685) );
  FA_X1 U607 ( .A(n941), .B(n959), .CI(n977), .CO(n686), .S(n687) );
  FA_X1 U608 ( .A(n887), .B(n923), .CI(n995), .CO(n688), .S(n689) );
  FA_X1 U609 ( .A(n869), .B(n1014), .CI(n905), .CO(n690), .S(n691) );
  FA_X1 U610 ( .A(n697), .B(n708), .CI(n695), .CO(n692), .S(n693) );
  FA_X1 U611 ( .A(n710), .B(n703), .CI(n699), .CO(n694), .S(n695) );
  FA_X1 U612 ( .A(n712), .B(n714), .CI(n701), .CO(n696), .S(n697) );
  FA_X1 U613 ( .A(n705), .B(n996), .CI(n716), .CO(n698), .S(n699) );
  FA_X1 U614 ( .A(n1015), .B(n942), .CI(n978), .CO(n700), .S(n701) );
  HA_X1 U616 ( .A(n822), .B(n888), .CO(n704), .S(n705) );
  FA_X1 U617 ( .A(n711), .B(n720), .CI(n709), .CO(n706), .S(n707) );
  FA_X1 U618 ( .A(n713), .B(n715), .CI(n722), .CO(n708), .S(n709) );
  FA_X1 U619 ( .A(n724), .B(n726), .CI(n717), .CO(n710), .S(n711) );
  FA_X1 U620 ( .A(n961), .B(n979), .CI(n728), .CO(n712), .S(n713) );
  FA_X1 U621 ( .A(n907), .B(n997), .CI(n943), .CO(n714), .S(n715) );
  FA_X1 U622 ( .A(n889), .B(n925), .CI(n1016), .CO(n716), .S(n717) );
  FA_X1 U623 ( .A(n732), .B(n723), .CI(n721), .CO(n718), .S(n719) );
  FA_X1 U624 ( .A(n727), .B(n725), .CI(n734), .CO(n720), .S(n721) );
  FA_X1 U625 ( .A(n738), .B(n729), .CI(n736), .CO(n722), .S(n723) );
  FA_X1 U626 ( .A(n926), .B(n980), .CI(n944), .CO(n724), .S(n725) );
  FA_X1 U627 ( .A(n1017), .B(n962), .CI(n998), .CO(n726), .S(n727) );
  HA_X1 U628 ( .A(n823), .B(n908), .CO(n728), .S(n729) );
  FA_X1 U629 ( .A(n735), .B(n742), .CI(n733), .CO(n730), .S(n731) );
  FA_X1 U630 ( .A(n737), .B(n739), .CI(n744), .CO(n732), .S(n733) );
  FA_X1 U631 ( .A(n748), .B(n981), .CI(n746), .CO(n734), .S(n735) );
  FA_X1 U632 ( .A(n927), .B(n999), .CI(n963), .CO(n736), .S(n737) );
  FA_X1 U633 ( .A(n945), .B(n909), .CI(n1018), .CO(n738), .S(n739) );
  FA_X1 U634 ( .A(n752), .B(n745), .CI(n743), .CO(n740), .S(n741) );
  FA_X1 U635 ( .A(n754), .B(n756), .CI(n747), .CO(n742), .S(n743) );
  FA_X1 U636 ( .A(n964), .B(n1000), .CI(n749), .CO(n744), .S(n745) );
  FA_X1 U637 ( .A(n946), .B(n982), .CI(n1019), .CO(n746), .S(n747) );
  HA_X1 U638 ( .A(n824), .B(n928), .CO(n748), .S(n749) );
  FA_X1 U639 ( .A(n760), .B(n755), .CI(n753), .CO(n750), .S(n751) );
  FA_X1 U640 ( .A(n762), .B(n764), .CI(n757), .CO(n752), .S(n753) );
  FA_X1 U641 ( .A(n947), .B(n1001), .CI(n983), .CO(n754), .S(n755) );
  FA_X1 U642 ( .A(n965), .B(n929), .CI(n1020), .CO(n756), .S(n757) );
  FA_X1 U643 ( .A(n763), .B(n768), .CI(n761), .CO(n758), .S(n759) );
  FA_X1 U644 ( .A(n765), .B(n1021), .CI(n770), .CO(n760), .S(n761) );
  FA_X1 U645 ( .A(n966), .B(n984), .CI(n1002), .CO(n762), .S(n763) );
  HA_X1 U646 ( .A(n825), .B(n948), .CO(n764), .S(n765) );
  FA_X1 U647 ( .A(n771), .B(n774), .CI(n769), .CO(n766), .S(n767) );
  FA_X1 U648 ( .A(n967), .B(n1003), .CI(n776), .CO(n768), .S(n769) );
  FA_X1 U649 ( .A(n985), .B(n949), .CI(n1022), .CO(n770), .S(n771) );
  FA_X1 U650 ( .A(n780), .B(n777), .CI(n775), .CO(n772), .S(n773) );
  FA_X1 U651 ( .A(n986), .B(n1023), .CI(n1004), .CO(n774), .S(n775) );
  HA_X1 U652 ( .A(n826), .B(n968), .CO(n776), .S(n777) );
  FA_X1 U653 ( .A(n784), .B(n987), .CI(n781), .CO(n778), .S(n779) );
  FA_X1 U654 ( .A(n1024), .B(n969), .CI(n1005), .CO(n780), .S(n781) );
  FA_X1 U655 ( .A(n1006), .B(n1025), .CI(n785), .CO(n782), .S(n783) );
  HA_X1 U656 ( .A(n827), .B(n988), .CO(n784), .S(n785) );
  FA_X1 U657 ( .A(n1026), .B(n989), .CI(n1007), .CO(n786), .S(n787) );
  HA_X1 U658 ( .A(n1008), .B(n1027), .CO(n788), .S(n789) );
  BUF_X2 U1180 ( .A(n1277), .Z(n1383) );
  OAI21_X1 U1181 ( .B1(n284), .B2(n290), .A(n285), .ZN(n1384) );
  INV_X1 U1182 ( .A(n1298), .ZN(n1385) );
  CLKBUF_X3 U1183 ( .A(b[18]), .Z(n1241) );
  CLKBUF_X2 U1184 ( .A(b[11]), .Z(n1248) );
  CLKBUF_X3 U1185 ( .A(b[7]), .Z(n1252) );
  CLKBUF_X3 U1186 ( .A(b[9]), .Z(n1250) );
  CLKBUF_X3 U1187 ( .A(n1277), .Z(n17) );
  CLKBUF_X3 U1188 ( .A(b[15]), .Z(n1244) );
  CLKBUF_X3 U1189 ( .A(n1279), .Z(n1441) );
  CLKBUF_X1 U1190 ( .A(n1279), .Z(n5) );
  CLKBUF_X3 U1191 ( .A(b[14]), .Z(n1245) );
  CLKBUF_X3 U1192 ( .A(b[16]), .Z(n1243) );
  CLKBUF_X3 U1193 ( .A(n291), .Z(n64) );
  CLKBUF_X3 U1194 ( .A(b[17]), .Z(n1242) );
  CLKBUF_X3 U1195 ( .A(b[2]), .Z(n1257) );
  BUF_X2 U1196 ( .A(a[15]), .Z(n1447) );
  BUF_X2 U1197 ( .A(n1270), .Z(n59) );
  BUF_X2 U1198 ( .A(n1276), .Z(n24) );
  BUF_X2 U1199 ( .A(n1386), .Z(n1458) );
  CLKBUF_X3 U1200 ( .A(b[13]), .Z(n1246) );
  AOI21_X1 U1201 ( .B1(n1384), .B2(n249), .A(n250), .ZN(n1386) );
  CLKBUF_X3 U1202 ( .A(b[1]), .Z(n1258) );
  CLKBUF_X1 U1203 ( .A(n1161), .Z(n1387) );
  CLKBUF_X1 U1204 ( .A(b[4]), .Z(n1388) );
  CLKBUF_X1 U1205 ( .A(b[4]), .Z(n1389) );
  CLKBUF_X1 U1206 ( .A(b[4]), .Z(n1255) );
  CLKBUF_X3 U1207 ( .A(b[6]), .Z(n1253) );
  CLKBUF_X3 U1208 ( .A(b[10]), .Z(n1249) );
  BUF_X2 U1209 ( .A(a[11]), .Z(n1448) );
  OAI22_X1 U1210 ( .A1(n60), .A2(n1031), .B1(n58), .B2(n1030), .ZN(n448) );
  BUF_X1 U1211 ( .A(n247), .Z(n66) );
  OR2_X1 U1212 ( .A1(n473), .A2(n480), .ZN(n1390) );
  OR2_X1 U1213 ( .A1(n453), .A2(n456), .ZN(n1391) );
  OR2_X1 U1214 ( .A1(n467), .A2(n472), .ZN(n1392) );
  OR2_X1 U1215 ( .A1(n830), .A2(n448), .ZN(n1393) );
  OR2_X1 U1216 ( .A1(n452), .A2(n451), .ZN(n1394) );
  OR2_X1 U1217 ( .A1(n759), .A2(n766), .ZN(n1395) );
  OR2_X1 U1218 ( .A1(n450), .A2(n449), .ZN(n1396) );
  OR2_X1 U1219 ( .A1(n457), .A2(n460), .ZN(n1397) );
  OR2_X1 U1220 ( .A1(n767), .A2(n772), .ZN(n1398) );
  OR2_X1 U1221 ( .A1(n779), .A2(n782), .ZN(n1399) );
  OR2_X1 U1222 ( .A1(n787), .A2(n788), .ZN(n1400) );
  BUF_X2 U1223 ( .A(a[5]), .Z(n1445) );
  CLKBUF_X2 U1224 ( .A(a[5]), .Z(n13) );
  NOR2_X1 U1225 ( .A1(n461), .A2(n466), .ZN(n179) );
  NOR2_X1 U1226 ( .A1(n561), .A2(n576), .ZN(n289) );
  OR2_X1 U1227 ( .A1(n1029), .A2(n829), .ZN(n1401) );
  NOR2_X1 U1228 ( .A1(n533), .A2(n546), .ZN(n275) );
  CLKBUF_X1 U1229 ( .A(a[0]), .Z(n1402) );
  CLKBUF_X1 U1230 ( .A(n331), .Z(n1403) );
  OR2_X1 U1231 ( .A1(n693), .A2(n706), .ZN(n1404) );
  NOR2_X1 U1232 ( .A1(n1466), .A2(n326), .ZN(n1405) );
  XNOR2_X1 U1233 ( .A(n1), .B(n1243), .ZN(n1406) );
  BUF_X1 U1234 ( .A(n1285), .Z(n27) );
  NOR2_X1 U1235 ( .A1(n593), .A2(n610), .ZN(n1407) );
  CLKBUF_X1 U1236 ( .A(n1240), .Z(n1408) );
  CLKBUF_X1 U1237 ( .A(n304), .Z(n1409) );
  CLKBUF_X1 U1238 ( .A(n340), .Z(n1410) );
  CLKBUF_X3 U1239 ( .A(n1272), .Z(n1411) );
  CLKBUF_X1 U1240 ( .A(n1272), .Z(n47) );
  BUF_X2 U1241 ( .A(n1274), .Z(n1412) );
  CLKBUF_X1 U1242 ( .A(n1274), .Z(n35) );
  OR2_X2 U1243 ( .A1(n509), .A2(n520), .ZN(n1413) );
  XNOR2_X1 U1244 ( .A(n31), .B(n1253), .ZN(n1414) );
  CLKBUF_X1 U1245 ( .A(n1281), .Z(n51) );
  CLKBUF_X2 U1246 ( .A(n1281), .Z(n52) );
  BUF_X2 U1247 ( .A(a[19]), .Z(n1429) );
  BUF_X1 U1248 ( .A(a[19]), .Z(n1428) );
  BUF_X1 U1249 ( .A(n1286), .Z(n22) );
  BUF_X1 U1250 ( .A(n1286), .Z(n21) );
  BUF_X1 U1251 ( .A(n1278), .Z(n12) );
  BUF_X2 U1252 ( .A(n1421), .Z(n10) );
  BUF_X2 U1253 ( .A(b[19]), .Z(n1240) );
  CLKBUF_X2 U1254 ( .A(n1284), .Z(n33) );
  BUF_X1 U1255 ( .A(n1284), .Z(n34) );
  OR2_X1 U1256 ( .A1(n663), .A2(n678), .ZN(n1443) );
  XOR2_X1 U1257 ( .A(n906), .B(n960), .Z(n1415) );
  XOR2_X1 U1258 ( .A(n924), .B(n1415), .Z(n703) );
  NAND2_X1 U1259 ( .A1(n924), .A2(n906), .ZN(n1416) );
  NAND2_X1 U1260 ( .A1(n924), .A2(n960), .ZN(n1417) );
  NAND2_X1 U1261 ( .A1(n906), .A2(n960), .ZN(n1418) );
  NAND3_X1 U1262 ( .A1(n1416), .A2(n1417), .A3(n1418), .ZN(n702) );
  CLKBUF_X1 U1263 ( .A(n317), .Z(n1419) );
  BUF_X2 U1264 ( .A(a[9]), .Z(n25) );
  XNOR2_X1 U1265 ( .A(n1429), .B(n1388), .ZN(n1420) );
  XNOR2_X1 U1266 ( .A(a[1]), .B(a[2]), .ZN(n1421) );
  XNOR2_X1 U1267 ( .A(n13), .B(n1241), .ZN(n1422) );
  XNOR2_X1 U1268 ( .A(n286), .B(n1423), .ZN(product[24]) );
  AND2_X1 U1269 ( .A1(n424), .A2(n285), .ZN(n1423) );
  CLKBUF_X1 U1270 ( .A(n63), .Z(n1424) );
  BUF_X1 U1271 ( .A(n1285), .Z(n28) );
  XNOR2_X1 U1272 ( .A(n13), .B(n1242), .ZN(n1425) );
  CLKBUF_X1 U1273 ( .A(n296), .Z(n1426) );
  XNOR2_X1 U1274 ( .A(n7), .B(n1240), .ZN(n1427) );
  CLKBUF_X3 U1275 ( .A(a[1]), .Z(n1442) );
  BUF_X2 U1276 ( .A(a[1]), .Z(n1) );
  CLKBUF_X1 U1277 ( .A(n1282), .Z(n46) );
  BUF_X1 U1278 ( .A(n1282), .Z(n45) );
  OR2_X1 U1279 ( .A1(n692), .A2(n679), .ZN(n1430) );
  XNOR2_X1 U1280 ( .A(n613), .B(n1431), .ZN(n611) );
  XNOR2_X1 U1281 ( .A(n630), .B(n615), .ZN(n1431) );
  NOR2_X1 U1282 ( .A1(n296), .A2(n1407), .ZN(n1432) );
  BUF_X2 U1283 ( .A(n247), .Z(n1433) );
  CLKBUF_X1 U1284 ( .A(n1407), .Z(n1434) );
  XNOR2_X1 U1285 ( .A(n1), .B(n1240), .ZN(n1435) );
  CLKBUF_X1 U1286 ( .A(n1280), .Z(n58) );
  CLKBUF_X2 U1287 ( .A(n1280), .Z(n57) );
  CLKBUF_X1 U1288 ( .A(n37), .Z(n1436) );
  XNOR2_X1 U1289 ( .A(n43), .B(n1255), .ZN(n1437) );
  XNOR2_X1 U1290 ( .A(n1428), .B(n1258), .ZN(n1438) );
  CLKBUF_X1 U1291 ( .A(n1421), .Z(n9) );
  XNOR2_X1 U1292 ( .A(n31), .B(n1249), .ZN(n1439) );
  BUF_X2 U1293 ( .A(a[11]), .Z(n31) );
  CLKBUF_X3 U1294 ( .A(a[9]), .Z(n1440) );
  CLKBUF_X1 U1295 ( .A(n1279), .Z(n6) );
  CLKBUF_X1 U1296 ( .A(n1257), .Z(n1444) );
  XNOR2_X1 U1297 ( .A(n1428), .B(n1256), .ZN(n1446) );
  CLKBUF_X1 U1298 ( .A(a[15]), .Z(n43) );
  CLKBUF_X3 U1299 ( .A(n61), .Z(n1481) );
  OAI22_X1 U1300 ( .A1(n24), .A2(n1157), .B1(n22), .B2(n1156), .ZN(n1449) );
  XNOR2_X1 U1301 ( .A(n1257), .B(n1429), .ZN(n1450) );
  CLKBUF_X3 U1302 ( .A(n61), .Z(n1451) );
  XNOR2_X1 U1303 ( .A(n244), .B(n1452), .ZN(product[28]) );
  AND2_X1 U1304 ( .A1(n240), .A2(n243), .ZN(n1452) );
  XNOR2_X1 U1305 ( .A(n268), .B(n1453), .ZN(product[26]) );
  AND2_X1 U1306 ( .A1(n262), .A2(n267), .ZN(n1453) );
  AOI21_X1 U1307 ( .B1(n1405), .B2(n340), .A(n322), .ZN(n1454) );
  XNOR2_X1 U1308 ( .A(n209), .B(n1455), .ZN(product[31]) );
  AND2_X1 U1309 ( .A1(n1390), .A2(n208), .ZN(n1455) );
  XNOR2_X1 U1310 ( .A(n231), .B(n1456), .ZN(product[29]) );
  AND2_X1 U1311 ( .A1(n227), .A2(n230), .ZN(n1456) );
  XNOR2_X1 U1312 ( .A(n277), .B(n1457), .ZN(product[25]) );
  AND2_X1 U1313 ( .A1(n273), .A2(n276), .ZN(n1457) );
  BUF_X1 U1314 ( .A(n1278), .Z(n1459) );
  BUF_X2 U1315 ( .A(n1278), .Z(n1460) );
  NOR2_X1 U1316 ( .A1(n577), .A2(n592), .ZN(n1461) );
  NAND2_X1 U1317 ( .A1(n613), .A2(n630), .ZN(n1462) );
  NAND2_X1 U1318 ( .A1(n613), .A2(n615), .ZN(n1463) );
  NAND2_X1 U1319 ( .A1(n630), .A2(n615), .ZN(n1464) );
  NAND3_X1 U1320 ( .A1(n1462), .A2(n1463), .A3(n1464), .ZN(n610) );
  XNOR2_X1 U1321 ( .A(n222), .B(n1465), .ZN(product[30]) );
  AND2_X1 U1322 ( .A1(n418), .A2(n221), .ZN(n1465) );
  NOR2_X1 U1323 ( .A1(n647), .A2(n662), .ZN(n1466) );
  NOR2_X1 U1324 ( .A1(n647), .A2(n662), .ZN(n323) );
  CLKBUF_X1 U1325 ( .A(n1240), .Z(n1467) );
  XOR2_X1 U1326 ( .A(n900), .B(n972), .Z(n1468) );
  XOR2_X1 U1327 ( .A(n846), .B(n1468), .Z(n607) );
  NAND2_X1 U1328 ( .A1(n846), .A2(n900), .ZN(n1469) );
  NAND2_X1 U1329 ( .A1(n846), .A2(n972), .ZN(n1470) );
  NAND2_X1 U1330 ( .A1(n900), .A2(n972), .ZN(n1471) );
  NAND3_X1 U1331 ( .A1(n1469), .A2(n1470), .A3(n1471), .ZN(n606) );
  INV_X1 U1332 ( .A(n338), .ZN(n1472) );
  NOR2_X2 U1333 ( .A1(n547), .A2(n560), .ZN(n284) );
  BUF_X4 U1334 ( .A(a[13]), .Z(n37) );
  CLKBUF_X3 U1335 ( .A(b[8]), .Z(n1251) );
  OR2_X1 U1336 ( .A1(n521), .A2(n532), .ZN(n1473) );
  BUF_X2 U1337 ( .A(n248), .Z(n65) );
  CLKBUF_X3 U1338 ( .A(b[12]), .Z(n1247) );
  NOR2_X1 U1339 ( .A1(n629), .A2(n646), .ZN(n317) );
  BUF_X2 U1340 ( .A(n1277), .Z(n18) );
  CLKBUF_X3 U1341 ( .A(b[5]), .Z(n1254) );
  AOI21_X1 U1342 ( .B1(n1443), .B2(n336), .A(n329), .ZN(n1474) );
  XNOR2_X1 U1343 ( .A(n257), .B(n1475), .ZN(product[27]) );
  AND2_X1 U1344 ( .A1(n1413), .A2(n256), .ZN(n1475) );
  BUF_X1 U1345 ( .A(b[0]), .Z(n61) );
  CLKBUF_X3 U1346 ( .A(b[3]), .Z(n1256) );
  NAND2_X1 U1347 ( .A1(n1266), .A2(n1286), .ZN(n1276) );
  NAND2_X1 U1348 ( .A1(n1263), .A2(n1283), .ZN(n1273) );
  NOR2_X1 U1349 ( .A1(n216), .A2(n192), .ZN(n186) );
  XNOR2_X1 U1350 ( .A(n339), .B(n1476), .ZN(product[16]) );
  AND2_X1 U1351 ( .A1(n1430), .A2(n338), .ZN(n1476) );
  XNOR2_X1 U1352 ( .A(n198), .B(n1477), .ZN(product[32]) );
  AND2_X1 U1353 ( .A1(n1392), .A2(n197), .ZN(n1477) );
  NOR2_X1 U1354 ( .A1(n611), .A2(n628), .ZN(n312) );
  XNOR2_X1 U1355 ( .A(n168), .B(n1478), .ZN(product[34]) );
  AND2_X1 U1356 ( .A1(n1397), .A2(n167), .ZN(n1478) );
  NOR2_X1 U1357 ( .A1(n489), .A2(n498), .ZN(n229) );
  NOR2_X1 U1358 ( .A1(n707), .A2(n718), .ZN(n350) );
  NOR2_X1 U1359 ( .A1(n481), .A2(n488), .ZN(n220) );
  NOR2_X1 U1360 ( .A1(n741), .A2(n750), .ZN(n364) );
  NOR2_X1 U1361 ( .A1(n499), .A2(n508), .ZN(n242) );
  NAND2_X1 U1362 ( .A1(n461), .A2(n466), .ZN(n180) );
  NOR2_X1 U1363 ( .A1(n773), .A2(n778), .ZN(n386) );
  NOR2_X1 U1364 ( .A1(n789), .A2(n828), .ZN(n402) );
  AND2_X1 U1365 ( .A1(n1401), .A2(n409), .ZN(product[1]) );
  CLKBUF_X3 U1366 ( .A(n61), .Z(n1480) );
  BUF_X2 U1367 ( .A(n1287), .Z(n15) );
  BUF_X2 U1368 ( .A(n1287), .Z(n16) );
  BUF_X2 U1369 ( .A(n1275), .Z(n29) );
  BUF_X2 U1370 ( .A(n1276), .Z(n23) );
  BUF_X2 U1371 ( .A(n1273), .Z(n42) );
  BUF_X2 U1372 ( .A(n1273), .Z(n41) );
  INV_X1 U1373 ( .A(n1402), .ZN(n1289) );
  NAND2_X1 U1374 ( .A1(n1268), .A2(n1421), .ZN(n1278) );
  NAND2_X1 U1375 ( .A1(n1267), .A2(n1287), .ZN(n1277) );
  NAND2_X1 U1376 ( .A1(n1269), .A2(n1289), .ZN(n1279) );
  NOR2_X1 U1377 ( .A1(n280), .A2(n275), .ZN(n269) );
  NOR2_X1 U1378 ( .A1(n280), .A2(n260), .ZN(n258) );
  NAND2_X1 U1379 ( .A1(n214), .A2(n134), .ZN(n130) );
  INV_X1 U1380 ( .A(n308), .ZN(n306) );
  INV_X1 U1381 ( .A(n186), .ZN(n184) );
  INV_X1 U1382 ( .A(n173), .ZN(n171) );
  INV_X1 U1383 ( .A(n1433), .ZN(n245) );
  INV_X1 U1384 ( .A(n309), .ZN(n307) );
  INV_X1 U1385 ( .A(n281), .ZN(n279) );
  INV_X1 U1386 ( .A(n187), .ZN(n185) );
  INV_X1 U1387 ( .A(n282), .ZN(n280) );
  NOR2_X1 U1388 ( .A1(n216), .A2(n175), .ZN(n173) );
  INV_X1 U1389 ( .A(n1410), .ZN(n339) );
  INV_X1 U1390 ( .A(n311), .ZN(n309) );
  INV_X1 U1391 ( .A(n216), .ZN(n214) );
  INV_X1 U1392 ( .A(n1384), .ZN(n281) );
  NAND2_X1 U1393 ( .A1(n1443), .A2(n1430), .ZN(n326) );
  NAND2_X1 U1394 ( .A1(n273), .A2(n262), .ZN(n260) );
  OAI21_X1 U1395 ( .B1(n281), .B2(n275), .A(n276), .ZN(n270) );
  OAI21_X1 U1396 ( .B1(n281), .B2(n260), .A(n261), .ZN(n259) );
  AOI21_X1 U1397 ( .B1(n274), .B2(n262), .A(n265), .ZN(n261) );
  NAND2_X1 U1398 ( .A1(n1473), .A2(n1413), .ZN(n251) );
  NOR2_X1 U1399 ( .A1(n308), .A2(n1434), .ZN(n299) );
  INV_X1 U1400 ( .A(n192), .ZN(n190) );
  INV_X1 U1401 ( .A(n263), .ZN(n262) );
  INV_X1 U1402 ( .A(n1473), .ZN(n263) );
  NAND2_X1 U1403 ( .A1(n186), .A2(n149), .ZN(n145) );
  INV_X1 U1404 ( .A(n1430), .ZN(n333) );
  NAND2_X1 U1405 ( .A1(n214), .A2(n1390), .ZN(n201) );
  INV_X1 U1406 ( .A(n336), .ZN(n334) );
  INV_X1 U1407 ( .A(n119), .ZN(n117) );
  NAND2_X1 U1408 ( .A1(n315), .A2(n318), .ZN(n86) );
  XOR2_X1 U1409 ( .A(n347), .B(n90), .Z(product[15]) );
  NAND2_X1 U1410 ( .A1(n1404), .A2(n346), .ZN(n90) );
  XNOR2_X1 U1411 ( .A(n325), .B(n87), .ZN(product[18]) );
  OAI21_X1 U1412 ( .B1(n339), .B2(n326), .A(n1474), .ZN(n325) );
  NAND2_X1 U1413 ( .A1(n430), .A2(n324), .ZN(n87) );
  INV_X1 U1414 ( .A(n1466), .ZN(n430) );
  NAND2_X1 U1415 ( .A1(n218), .A2(n240), .ZN(n216) );
  INV_X1 U1416 ( .A(n284), .ZN(n424) );
  NOR2_X1 U1417 ( .A1(n1466), .A2(n326), .ZN(n321) );
  OAI21_X1 U1418 ( .B1(n284), .B2(n290), .A(n285), .ZN(n283) );
  NAND2_X1 U1419 ( .A1(n287), .A2(n290), .ZN(n82) );
  XOR2_X1 U1420 ( .A(n314), .B(n85), .Z(product[20]) );
  NAND2_X1 U1421 ( .A1(n428), .A2(n313), .ZN(n85) );
  INV_X1 U1422 ( .A(n312), .ZN(n428) );
  OAI21_X1 U1423 ( .B1(n217), .B2(n192), .A(n193), .ZN(n187) );
  XNOR2_X1 U1424 ( .A(n332), .B(n88), .ZN(product[17]) );
  NAND2_X1 U1425 ( .A1(n1443), .A2(n1403), .ZN(n88) );
  OAI21_X1 U1426 ( .B1(n339), .B2(n333), .A(n334), .ZN(n332) );
  NOR2_X1 U1427 ( .A1(n216), .A2(n121), .ZN(n119) );
  AOI21_X1 U1428 ( .B1(n1443), .B2(n1472), .A(n329), .ZN(n327) );
  INV_X1 U1429 ( .A(n331), .ZN(n329) );
  XOR2_X1 U1430 ( .A(n298), .B(n83), .Z(product[22]) );
  NAND2_X1 U1431 ( .A1(n426), .A2(n297), .ZN(n83) );
  XOR2_X1 U1432 ( .A(n305), .B(n84), .Z(product[21]) );
  NAND2_X1 U1433 ( .A1(n302), .A2(n1409), .ZN(n84) );
  AOI21_X1 U1434 ( .B1(n1413), .B2(n265), .A(n254), .ZN(n252) );
  NOR2_X1 U1435 ( .A1(n192), .A2(n136), .ZN(n134) );
  INV_X1 U1436 ( .A(n174), .ZN(n172) );
  AOI21_X1 U1437 ( .B1(n215), .B2(n1390), .A(n206), .ZN(n202) );
  INV_X1 U1438 ( .A(n217), .ZN(n215) );
  INV_X1 U1439 ( .A(n275), .ZN(n273) );
  NAND2_X1 U1440 ( .A1(n190), .A2(n177), .ZN(n175) );
  INV_X1 U1441 ( .A(n338), .ZN(n336) );
  NAND2_X1 U1442 ( .A1(n1390), .A2(n1392), .ZN(n192) );
  OAI21_X1 U1443 ( .B1(n309), .B2(n1434), .A(n1409), .ZN(n300) );
  NOR2_X1 U1444 ( .A1(n251), .A2(n275), .ZN(n249) );
  INV_X1 U1445 ( .A(n267), .ZN(n265) );
  INV_X1 U1446 ( .A(n276), .ZN(n274) );
  INV_X1 U1447 ( .A(n193), .ZN(n191) );
  INV_X1 U1448 ( .A(n256), .ZN(n254) );
  NAND2_X1 U1449 ( .A1(n240), .A2(n227), .ZN(n225) );
  NAND2_X1 U1450 ( .A1(n173), .A2(n1397), .ZN(n160) );
  INV_X1 U1451 ( .A(n289), .ZN(n287) );
  INV_X1 U1452 ( .A(n1419), .ZN(n315) );
  INV_X1 U1453 ( .A(n290), .ZN(n288) );
  INV_X1 U1454 ( .A(n346), .ZN(n344) );
  INV_X1 U1455 ( .A(n318), .ZN(n316) );
  XOR2_X1 U1456 ( .A(n352), .B(n91), .Z(product[14]) );
  NAND2_X1 U1457 ( .A1(n434), .A2(n351), .ZN(n91) );
  INV_X1 U1458 ( .A(n350), .ZN(n434) );
  XOR2_X1 U1459 ( .A(n374), .B(n95), .Z(product[10]) );
  NAND2_X1 U1460 ( .A1(n438), .A2(n373), .ZN(n95) );
  AOI21_X1 U1461 ( .B1(n379), .B2(n1395), .A(n376), .ZN(n374) );
  INV_X1 U1462 ( .A(n372), .ZN(n438) );
  AOI21_X1 U1463 ( .B1(n218), .B2(n241), .A(n219), .ZN(n217) );
  XNOR2_X1 U1464 ( .A(n363), .B(n93), .ZN(product[12]) );
  NAND2_X1 U1465 ( .A1(n436), .A2(n362), .ZN(n93) );
  OAI21_X1 U1466 ( .B1(n366), .B2(n364), .A(n365), .ZN(n363) );
  INV_X1 U1467 ( .A(n361), .ZN(n436) );
  XNOR2_X1 U1468 ( .A(n357), .B(n92), .ZN(product[13]) );
  NAND2_X1 U1469 ( .A1(n435), .A2(n356), .ZN(n92) );
  INV_X1 U1470 ( .A(n355), .ZN(n435) );
  XNOR2_X1 U1471 ( .A(n379), .B(n96), .ZN(product[9]) );
  NAND2_X1 U1472 ( .A1(n1395), .A2(n378), .ZN(n96) );
  INV_X1 U1473 ( .A(n220), .ZN(n418) );
  NOR2_X1 U1474 ( .A1(n229), .A2(n220), .ZN(n218) );
  AOI21_X1 U1475 ( .B1(n1392), .B2(n206), .A(n195), .ZN(n193) );
  INV_X1 U1476 ( .A(n197), .ZN(n195) );
  XOR2_X1 U1477 ( .A(n181), .B(n72), .Z(product[33]) );
  NAND2_X1 U1478 ( .A1(n177), .A2(n180), .ZN(n72) );
  AOI21_X1 U1479 ( .B1(n63), .B2(n182), .A(n183), .ZN(n181) );
  OAI21_X1 U1480 ( .B1(n217), .B2(n175), .A(n176), .ZN(n174) );
  AOI21_X1 U1481 ( .B1(n191), .B2(n177), .A(n178), .ZN(n176) );
  INV_X1 U1482 ( .A(n180), .ZN(n178) );
  NAND2_X1 U1483 ( .A1(n561), .A2(n576), .ZN(n290) );
  NOR2_X1 U1484 ( .A1(n593), .A2(n610), .ZN(n303) );
  NOR2_X1 U1485 ( .A1(n179), .A2(n151), .ZN(n149) );
  NAND2_X1 U1486 ( .A1(n663), .A2(n678), .ZN(n331) );
  AOI21_X1 U1487 ( .B1(n174), .B2(n1397), .A(n165), .ZN(n161) );
  AOI21_X1 U1488 ( .B1(n241), .B2(n227), .A(n228), .ZN(n226) );
  INV_X1 U1489 ( .A(n230), .ZN(n228) );
  INV_X1 U1490 ( .A(n120), .ZN(n118) );
  AOI21_X1 U1491 ( .B1(n187), .B2(n149), .A(n150), .ZN(n146) );
  AOI21_X1 U1492 ( .B1(n215), .B2(n134), .A(n135), .ZN(n131) );
  OAI21_X1 U1493 ( .B1(n368), .B2(n380), .A(n369), .ZN(n367) );
  NAND2_X1 U1494 ( .A1(n370), .A2(n1395), .ZN(n368) );
  AOI21_X1 U1495 ( .B1(n370), .B2(n376), .A(n371), .ZN(n369) );
  INV_X1 U1496 ( .A(n372), .ZN(n370) );
  OAI21_X1 U1497 ( .B1(n350), .B2(n356), .A(n351), .ZN(n349) );
  INV_X1 U1498 ( .A(n208), .ZN(n206) );
  NAND2_X1 U1499 ( .A1(n533), .A2(n546), .ZN(n276) );
  NAND2_X1 U1500 ( .A1(n629), .A2(n646), .ZN(n318) );
  NAND2_X1 U1501 ( .A1(n593), .A2(n610), .ZN(n304) );
  INV_X1 U1502 ( .A(n380), .ZN(n379) );
  NAND2_X1 U1503 ( .A1(n693), .A2(n706), .ZN(n346) );
  NAND2_X1 U1504 ( .A1(n521), .A2(n532), .ZN(n267) );
  NAND2_X1 U1505 ( .A1(n547), .A2(n560), .ZN(n285) );
  INV_X1 U1506 ( .A(n179), .ZN(n177) );
  NAND2_X1 U1507 ( .A1(n1397), .A2(n1391), .ZN(n151) );
  NAND2_X1 U1508 ( .A1(n149), .A2(n1394), .ZN(n136) );
  NAND2_X1 U1509 ( .A1(n134), .A2(n1396), .ZN(n121) );
  NAND2_X1 U1510 ( .A1(n647), .A2(n662), .ZN(n324) );
  NAND2_X1 U1511 ( .A1(n611), .A2(n628), .ZN(n313) );
  INV_X1 U1512 ( .A(n229), .ZN(n227) );
  NAND2_X1 U1513 ( .A1(n577), .A2(n592), .ZN(n297) );
  INV_X1 U1514 ( .A(n242), .ZN(n240) );
  INV_X1 U1515 ( .A(n243), .ZN(n241) );
  INV_X1 U1516 ( .A(n378), .ZN(n376) );
  AOI21_X1 U1517 ( .B1(n1424), .B2(n106), .A(n107), .ZN(n105) );
  XOR2_X1 U1518 ( .A(n366), .B(n94), .Z(product[11]) );
  NAND2_X1 U1519 ( .A1(n437), .A2(n365), .ZN(n94) );
  INV_X1 U1520 ( .A(n364), .ZN(n437) );
  NAND2_X1 U1521 ( .A1(n119), .A2(n1393), .ZN(n108) );
  INV_X1 U1522 ( .A(n373), .ZN(n371) );
  INV_X1 U1523 ( .A(n356), .ZN(n354) );
  NAND2_X1 U1524 ( .A1(n1399), .A2(n392), .ZN(n99) );
  XOR2_X1 U1525 ( .A(n114), .B(n67), .Z(product[38]) );
  NAND2_X1 U1526 ( .A1(n1393), .A2(n113), .ZN(n67) );
  XOR2_X1 U1527 ( .A(n100), .B(n396), .Z(product[5]) );
  NAND2_X1 U1528 ( .A1(n443), .A2(n395), .ZN(n100) );
  INV_X1 U1529 ( .A(n394), .ZN(n443) );
  XNOR2_X1 U1530 ( .A(n385), .B(n97), .ZN(product[8]) );
  NAND2_X1 U1531 ( .A1(n1398), .A2(n384), .ZN(n97) );
  NAND2_X1 U1532 ( .A1(n1391), .A2(n156), .ZN(n70) );
  OAI21_X1 U1533 ( .B1(n388), .B2(n386), .A(n387), .ZN(n385) );
  XOR2_X1 U1534 ( .A(n127), .B(n68), .Z(product[37]) );
  NAND2_X1 U1535 ( .A1(n1396), .A2(n126), .ZN(n68) );
  OAI21_X1 U1536 ( .B1(n394), .B2(n396), .A(n395), .ZN(n393) );
  NAND2_X1 U1537 ( .A1(n489), .A2(n498), .ZN(n230) );
  XOR2_X1 U1538 ( .A(n142), .B(n69), .Z(product[36]) );
  NAND2_X1 U1539 ( .A1(n1394), .A2(n141), .ZN(n69) );
  NOR2_X1 U1540 ( .A1(n719), .A2(n730), .ZN(n355) );
  AOI21_X1 U1541 ( .B1(n385), .B2(n1398), .A(n382), .ZN(n380) );
  INV_X1 U1542 ( .A(n384), .ZN(n382) );
  NOR2_X1 U1543 ( .A1(n731), .A2(n740), .ZN(n361) );
  OAI21_X1 U1544 ( .B1(n151), .B2(n180), .A(n152), .ZN(n150) );
  AOI21_X1 U1545 ( .B1(n165), .B2(n1391), .A(n154), .ZN(n152) );
  INV_X1 U1546 ( .A(n156), .ZN(n154) );
  OAI21_X1 U1547 ( .B1(n193), .B2(n136), .A(n137), .ZN(n135) );
  AOI21_X1 U1548 ( .B1(n150), .B2(n1394), .A(n139), .ZN(n137) );
  INV_X1 U1549 ( .A(n141), .ZN(n139) );
  OAI21_X1 U1550 ( .B1(n217), .B2(n121), .A(n122), .ZN(n120) );
  AOI21_X1 U1551 ( .B1(n135), .B2(n1396), .A(n124), .ZN(n122) );
  INV_X1 U1552 ( .A(n126), .ZN(n124) );
  NOR2_X1 U1553 ( .A1(n751), .A2(n758), .ZN(n372) );
  NAND2_X1 U1554 ( .A1(n719), .A2(n730), .ZN(n356) );
  NAND2_X1 U1555 ( .A1(n741), .A2(n750), .ZN(n365) );
  AOI21_X1 U1556 ( .B1(n120), .B2(n1393), .A(n111), .ZN(n109) );
  INV_X1 U1557 ( .A(n113), .ZN(n111) );
  NAND2_X1 U1558 ( .A1(n467), .A2(n472), .ZN(n197) );
  NAND2_X1 U1559 ( .A1(n499), .A2(n508), .ZN(n243) );
  NAND2_X1 U1560 ( .A1(n759), .A2(n766), .ZN(n378) );
  NAND2_X1 U1561 ( .A1(n751), .A2(n758), .ZN(n373) );
  NAND2_X1 U1562 ( .A1(n707), .A2(n718), .ZN(n351) );
  NAND2_X1 U1563 ( .A1(n731), .A2(n740), .ZN(n362) );
  NAND2_X1 U1564 ( .A1(n481), .A2(n488), .ZN(n221) );
  INV_X1 U1565 ( .A(n167), .ZN(n165) );
  AOI21_X1 U1566 ( .B1(n1399), .B2(n393), .A(n390), .ZN(n388) );
  INV_X1 U1567 ( .A(n392), .ZN(n390) );
  NAND2_X1 U1568 ( .A1(n441), .A2(n387), .ZN(n98) );
  INV_X1 U1569 ( .A(n386), .ZN(n441) );
  XOR2_X1 U1570 ( .A(n102), .B(n404), .Z(product[3]) );
  NAND2_X1 U1571 ( .A1(n445), .A2(n403), .ZN(n102) );
  INV_X1 U1572 ( .A(n402), .ZN(n445) );
  XOR2_X1 U1573 ( .A(n103), .B(n409), .Z(product[2]) );
  NAND2_X1 U1574 ( .A1(n446), .A2(n407), .ZN(n103) );
  INV_X1 U1575 ( .A(n406), .ZN(n446) );
  XNOR2_X1 U1576 ( .A(n101), .B(n401), .ZN(product[4]) );
  NAND2_X1 U1577 ( .A1(n1400), .A2(n400), .ZN(n101) );
  NOR2_X1 U1578 ( .A1(n1028), .A2(n1009), .ZN(n406) );
  OAI21_X1 U1579 ( .B1(n402), .B2(n404), .A(n403), .ZN(n401) );
  AOI21_X1 U1580 ( .B1(n1400), .B2(n401), .A(n398), .ZN(n396) );
  INV_X1 U1581 ( .A(n400), .ZN(n398) );
  NAND2_X1 U1582 ( .A1(n830), .A2(n448), .ZN(n113) );
  NOR2_X1 U1583 ( .A1(n783), .A2(n786), .ZN(n394) );
  INV_X1 U1584 ( .A(n448), .ZN(n449) );
  INV_X1 U1585 ( .A(n1449), .ZN(n545) );
  INV_X1 U1586 ( .A(n478), .ZN(n479) );
  OR2_X1 U1587 ( .A1(n937), .A2(n865), .ZN(n626) );
  XNOR2_X1 U1588 ( .A(n937), .B(n865), .ZN(n627) );
  NAND2_X1 U1589 ( .A1(n457), .A2(n460), .ZN(n167) );
  NAND2_X1 U1590 ( .A1(n779), .A2(n782), .ZN(n392) );
  NAND2_X1 U1591 ( .A1(n452), .A2(n451), .ZN(n141) );
  NAND2_X1 U1592 ( .A1(n450), .A2(n449), .ZN(n126) );
  NAND2_X1 U1593 ( .A1(n453), .A2(n456), .ZN(n156) );
  NAND2_X1 U1594 ( .A1(n767), .A2(n772), .ZN(n384) );
  NAND2_X1 U1595 ( .A1(n773), .A2(n778), .ZN(n387) );
  NAND2_X1 U1596 ( .A1(n783), .A2(n786), .ZN(n395) );
  INV_X1 U1597 ( .A(n405), .ZN(n404) );
  OAI21_X1 U1598 ( .B1(n406), .B2(n409), .A(n407), .ZN(n405) );
  OAI22_X1 U1599 ( .A1(n36), .A2(n1115), .B1(n34), .B2(n1114), .ZN(n496) );
  OAI22_X1 U1600 ( .A1(n30), .A2(n1143), .B1(n28), .B2(n1142), .ZN(n937) );
  OAI22_X1 U1601 ( .A1(n42), .A2(n1094), .B1(n40), .B2(n1093), .ZN(n478) );
  OAI22_X1 U1602 ( .A1(n24), .A2(n1157), .B1(n21), .B2(n1156), .ZN(n544) );
  OAI22_X1 U1603 ( .A1(n1459), .A2(n1199), .B1(n10), .B2(n1427), .ZN(n608) );
  OAI22_X1 U1604 ( .A1(n17), .A2(n1422), .B1(n16), .B2(n1177), .ZN(n574) );
  OAI22_X1 U1605 ( .A1(n1411), .A2(n1073), .B1(n46), .B2(n1072), .ZN(n464) );
  OAI22_X1 U1606 ( .A1(n30), .A2(n1136), .B1(n28), .B2(n1135), .ZN(n518) );
  OAI22_X1 U1607 ( .A1(n53), .A2(n1067), .B1(n52), .B2(n1066), .ZN(n865) );
  OAI22_X1 U1608 ( .A1(n60), .A2(n1032), .B1(n58), .B2(n1031), .ZN(n831) );
  INV_X1 U1609 ( .A(n793), .ZN(n850) );
  AOI21_X1 U1610 ( .B1(n54), .B2(n52), .A(n1051), .ZN(n793) );
  OAI22_X1 U1611 ( .A1(n60), .A2(n1034), .B1(n58), .B2(n1033), .ZN(n833) );
  OAI22_X1 U1612 ( .A1(n1460), .A2(n1215), .B1(n9), .B2(n1214), .ZN(n1006) );
  OAI22_X1 U1613 ( .A1(n1441), .A2(n1234), .B1(n1233), .B2(n3), .ZN(n1025) );
  OAI22_X1 U1614 ( .A1(n1383), .A2(n1195), .B1(n15), .B2(n1194), .ZN(n987) );
  AND2_X1 U1615 ( .A1(n1481), .A2(n812), .ZN(n989) );
  OAI22_X1 U1616 ( .A1(n1459), .A2(n1216), .B1(n9), .B2(n1215), .ZN(n1007) );
  OAI22_X1 U1617 ( .A1(n1441), .A2(n1235), .B1(n1234), .B2(n3), .ZN(n1026) );
  OAI22_X1 U1618 ( .A1(n5), .A2(n1237), .B1(n1236), .B2(n3), .ZN(n1028) );
  OAI22_X1 U1619 ( .A1(n30), .A2(n1295), .B1(n1155), .B2(n28), .ZN(n825) );
  OAI22_X1 U1620 ( .A1(n29), .A2(n1154), .B1(n27), .B2(n1153), .ZN(n948) );
  OR2_X1 U1621 ( .A1(n1451), .A2(n1295), .ZN(n1155) );
  OAI22_X1 U1622 ( .A1(n30), .A2(n1140), .B1(n28), .B2(n1139), .ZN(n934) );
  OAI22_X1 U1623 ( .A1(n1411), .A2(n1083), .B1(n46), .B2(n1082), .ZN(n880) );
  OAI22_X1 U1624 ( .A1(n24), .A2(n1159), .B1(n22), .B2(n1158), .ZN(n952) );
  OAI22_X1 U1625 ( .A1(n60), .A2(n1420), .B1(n57), .B2(n1044), .ZN(n844) );
  OAI22_X1 U1626 ( .A1(n36), .A2(n1121), .B1(n34), .B2(n1120), .ZN(n916) );
  OAI22_X1 U1627 ( .A1(n53), .A2(n1064), .B1(n52), .B2(n1063), .ZN(n862) );
  OAI22_X1 U1628 ( .A1(n59), .A2(n1043), .B1(n57), .B2(n1042), .ZN(n842) );
  OAI22_X1 U1629 ( .A1(n1411), .A2(n1081), .B1(n46), .B2(n1080), .ZN(n878) );
  OAI22_X1 U1630 ( .A1(n53), .A2(n1062), .B1(n52), .B2(n1061), .ZN(n860) );
  OAI22_X1 U1631 ( .A1(n29), .A2(n1147), .B1(n27), .B2(n1146), .ZN(n941) );
  OAI22_X1 U1632 ( .A1(n23), .A2(n1166), .B1(n21), .B2(n1165), .ZN(n959) );
  OAI22_X1 U1633 ( .A1(n1383), .A2(n1185), .B1(n16), .B2(n1184), .ZN(n977) );
  OAI22_X1 U1634 ( .A1(n48), .A2(n1086), .B1(n45), .B2(n1085), .ZN(n883) );
  OAI22_X1 U1635 ( .A1(n1460), .A2(n1200), .B1(n10), .B2(n1199), .ZN(n991) );
  OAI22_X1 U1636 ( .A1(n41), .A2(n1105), .B1(n39), .B2(n1104), .ZN(n901) );
  OAI22_X1 U1637 ( .A1(n1412), .A2(n1132), .B1(n33), .B2(n1131), .ZN(n927) );
  OAI22_X1 U1638 ( .A1(n23), .A2(n1170), .B1(n22), .B2(n1169), .ZN(n963) );
  OAI22_X1 U1639 ( .A1(n1460), .A2(n1208), .B1(n9), .B2(n1207), .ZN(n999) );
  AND2_X1 U1640 ( .A1(n1481), .A2(n791), .ZN(n849) );
  OAI22_X1 U1641 ( .A1(n47), .A2(n1088), .B1(n45), .B2(n1437), .ZN(n885) );
  OAI22_X1 U1642 ( .A1(n1441), .A2(n1221), .B1(n1220), .B2(n4), .ZN(n1012) );
  OAI22_X1 U1643 ( .A1(n29), .A2(n1151), .B1(n27), .B2(n1150), .ZN(n945) );
  AND2_X1 U1644 ( .A1(n1451), .A2(n800), .ZN(n909) );
  OAI22_X1 U1645 ( .A1(n1441), .A2(n1227), .B1(n1226), .B2(n4), .ZN(n1018) );
  OAI22_X1 U1646 ( .A1(n53), .A2(n1069), .B1(n52), .B2(n1068), .ZN(n867) );
  OAI22_X1 U1647 ( .A1(n1459), .A2(n1202), .B1(n10), .B2(n1201), .ZN(n993) );
  OAI22_X1 U1648 ( .A1(n41), .A2(n1107), .B1(n40), .B2(n1106), .ZN(n903) );
  OAI22_X1 U1649 ( .A1(n29), .A2(n1146), .B1(n27), .B2(n1145), .ZN(n940) );
  OAI22_X1 U1650 ( .A1(n5), .A2(n1406), .B1(n1221), .B2(n4), .ZN(n1013) );
  OAI22_X1 U1651 ( .A1(n1460), .A2(n1203), .B1(n10), .B2(n1202), .ZN(n994) );
  AOI21_X1 U1652 ( .B1(n6), .B2(n4), .A(n1219), .ZN(n817) );
  AOI21_X1 U1653 ( .B1(n42), .B2(n40), .A(n1093), .ZN(n799) );
  AOI21_X1 U1654 ( .B1(n1412), .B2(n34), .A(n1114), .ZN(n802) );
  AOI21_X1 U1655 ( .B1(n12), .B2(n10), .A(n1198), .ZN(n814) );
  INV_X1 U1656 ( .A(n790), .ZN(n830) );
  AOI21_X1 U1657 ( .B1(n60), .B2(n58), .A(n1030), .ZN(n790) );
  OAI22_X1 U1658 ( .A1(n54), .A2(n1291), .B1(n1071), .B2(n52), .ZN(n821) );
  OAI22_X1 U1659 ( .A1(n53), .A2(n1070), .B1(n51), .B2(n1069), .ZN(n868) );
  OR2_X1 U1660 ( .A1(n1480), .A2(n1291), .ZN(n1071) );
  OAI22_X1 U1661 ( .A1(n60), .A2(n1033), .B1(n58), .B2(n1032), .ZN(n832) );
  INV_X1 U1662 ( .A(n454), .ZN(n455) );
  NAND2_X1 U1663 ( .A1(n1029), .A2(n829), .ZN(n409) );
  NAND2_X1 U1664 ( .A1(n789), .A2(n828), .ZN(n403) );
  AND2_X1 U1665 ( .A1(n1451), .A2(n818), .ZN(product[0]) );
  INV_X1 U1666 ( .A(n3), .ZN(n818) );
  OAI22_X1 U1667 ( .A1(n60), .A2(n1040), .B1(n57), .B2(n1039), .ZN(n839) );
  INV_X1 U1668 ( .A(n805), .ZN(n930) );
  AOI21_X1 U1669 ( .B1(n30), .B2(n28), .A(n1135), .ZN(n805) );
  OAI22_X1 U1670 ( .A1(n35), .A2(n1128), .B1(n1127), .B2(n33), .ZN(n923) );
  OAI22_X1 U1671 ( .A1(n47), .A2(n1090), .B1(n1089), .B2(n45), .ZN(n887) );
  OAI22_X1 U1672 ( .A1(n12), .A2(n1204), .B1(n10), .B2(n1203), .ZN(n995) );
  OAI22_X1 U1673 ( .A1(n1412), .A2(n1125), .B1(n33), .B2(n1124), .ZN(n920) );
  OAI22_X1 U1674 ( .A1(n1459), .A2(n1201), .B1(n10), .B2(n1200), .ZN(n992) );
  OAI22_X1 U1675 ( .A1(n1383), .A2(n1182), .B1(n16), .B2(n1181), .ZN(n974) );
  OAI22_X1 U1676 ( .A1(n48), .A2(n1076), .B1(n46), .B2(n1075), .ZN(n873) );
  OAI22_X1 U1677 ( .A1(n54), .A2(n1057), .B1(n52), .B2(n1056), .ZN(n855) );
  OAI22_X1 U1678 ( .A1(n36), .A2(n1118), .B1(n34), .B2(n1117), .ZN(n913) );
  OAI22_X1 U1679 ( .A1(n30), .A2(n1137), .B1(n1136), .B2(n28), .ZN(n931) );
  OAI22_X1 U1680 ( .A1(n53), .A2(n1061), .B1(n51), .B2(n1060), .ZN(n859) );
  OAI22_X1 U1681 ( .A1(n1412), .A2(n1119), .B1(n34), .B2(n1118), .ZN(n914) );
  OAI22_X1 U1682 ( .A1(n30), .A2(n1138), .B1(n28), .B2(n1137), .ZN(n932) );
  OAI22_X1 U1683 ( .A1(n42), .A2(n1100), .B1(n39), .B2(n1099), .ZN(n896) );
  OAI22_X1 U1684 ( .A1(n1411), .A2(n1080), .B1(n46), .B2(n1079), .ZN(n877) );
  OAI22_X1 U1685 ( .A1(n42), .A2(n1099), .B1(n40), .B2(n1098), .ZN(n895) );
  OAI22_X1 U1686 ( .A1(n60), .A2(n1036), .B1(n58), .B2(n1035), .ZN(n835) );
  OAI22_X1 U1687 ( .A1(n54), .A2(n1055), .B1(n52), .B2(n1054), .ZN(n853) );
  INV_X1 U1688 ( .A(n799), .ZN(n890) );
  OAI22_X1 U1689 ( .A1(n24), .A2(n1162), .B1(n22), .B2(n1387), .ZN(n955) );
  OAI22_X1 U1690 ( .A1(n17), .A2(n1181), .B1(n16), .B2(n1180), .ZN(n973) );
  OAI22_X1 U1691 ( .A1(n1412), .A2(n1414), .B1(n33), .B2(n1126), .ZN(n922) );
  OAI22_X1 U1692 ( .A1(n48), .A2(n1089), .B1(n45), .B2(n1088), .ZN(n886) );
  OAI22_X1 U1693 ( .A1(n41), .A2(n1108), .B1(n40), .B2(n1107), .ZN(n904) );
  OAI22_X1 U1694 ( .A1(n1411), .A2(n1078), .B1(n46), .B2(n1077), .ZN(n875) );
  OAI22_X1 U1695 ( .A1(n36), .A2(n1116), .B1(n34), .B2(n1115), .ZN(n911) );
  OAI22_X1 U1696 ( .A1(n54), .A2(n1059), .B1(n52), .B2(n1058), .ZN(n857) );
  OAI22_X1 U1697 ( .A1(n24), .A2(n1165), .B1(n22), .B2(n1164), .ZN(n958) );
  OAI22_X1 U1698 ( .A1(n17), .A2(n1184), .B1(n16), .B2(n1183), .ZN(n976) );
  OAI22_X1 U1699 ( .A1(n1460), .A2(n1209), .B1(n9), .B2(n1208), .ZN(n1000) );
  OAI22_X1 U1700 ( .A1(n23), .A2(n1171), .B1(n22), .B2(n1170), .ZN(n964) );
  OAI22_X1 U1701 ( .A1(n24), .A2(n1164), .B1(n22), .B2(n1163), .ZN(n957) );
  OAI22_X1 U1702 ( .A1(n48), .A2(n1077), .B1(n46), .B2(n1076), .ZN(n874) );
  INV_X1 U1703 ( .A(n496), .ZN(n497) );
  AND2_X1 U1704 ( .A1(n1481), .A2(n794), .ZN(n869) );
  OAI22_X1 U1705 ( .A1(n6), .A2(n1223), .B1(n1222), .B2(n4), .ZN(n1014) );
  OAI22_X1 U1706 ( .A1(n41), .A2(n1109), .B1(n39), .B2(n1108), .ZN(n905) );
  OAI22_X1 U1707 ( .A1(n30), .A2(n1139), .B1(n28), .B2(n1138), .ZN(n933) );
  OAI22_X1 U1708 ( .A1(n53), .A2(n1063), .B1(n52), .B2(n1062), .ZN(n861) );
  OAI22_X1 U1709 ( .A1(n24), .A2(n1158), .B1(n22), .B2(n1157), .ZN(n951) );
  INV_X1 U1710 ( .A(n51), .ZN(n794) );
  OAI22_X1 U1711 ( .A1(n1129), .A2(n36), .B1(n33), .B2(n1128), .ZN(n924) );
  OAI22_X1 U1712 ( .A1(n41), .A2(n1110), .B1(n39), .B2(n1109), .ZN(n906) );
  OAI22_X1 U1713 ( .A1(n23), .A2(n1167), .B1(n21), .B2(n1166), .ZN(n960) );
  OAI22_X1 U1714 ( .A1(n1437), .A2(n47), .B1(n45), .B2(n1086), .ZN(n884) );
  OAI22_X1 U1715 ( .A1(n1144), .A2(n30), .B1(n28), .B2(n1143), .ZN(n938) );
  OAI22_X1 U1716 ( .A1(n53), .A2(n1068), .B1(n1067), .B2(n51), .ZN(n866) );
  OAI22_X1 U1717 ( .A1(n29), .A2(n1150), .B1(n27), .B2(n1149), .ZN(n944) );
  OAI22_X1 U1718 ( .A1(n36), .A2(n1131), .B1(n33), .B2(n1130), .ZN(n926) );
  OAI22_X1 U1719 ( .A1(n17), .A2(n1188), .B1(n15), .B2(n1187), .ZN(n980) );
  OAI22_X1 U1720 ( .A1(n1412), .A2(n1122), .B1(n34), .B2(n1121), .ZN(n917) );
  OAI22_X1 U1721 ( .A1(n59), .A2(n1450), .B1(n57), .B2(n1446), .ZN(n846) );
  OAI22_X1 U1722 ( .A1(n18), .A2(n1180), .B1(n16), .B2(n1179), .ZN(n972) );
  OAI22_X1 U1723 ( .A1(n41), .A2(n1104), .B1(n1103), .B2(n39), .ZN(n900) );
  OAI22_X1 U1724 ( .A1(n1411), .A2(n1084), .B1(n45), .B2(n1083), .ZN(n881) );
  OAI22_X1 U1725 ( .A1(n30), .A2(n1141), .B1(n28), .B2(n1140), .ZN(n935) );
  OAI22_X1 U1726 ( .A1(n41), .A2(n1103), .B1(n40), .B2(n1102), .ZN(n899) );
  OAI22_X1 U1727 ( .A1(n29), .A2(n1153), .B1(n27), .B2(n1152), .ZN(n947) );
  OAI22_X1 U1728 ( .A1(n1383), .A2(n1191), .B1(n15), .B2(n1190), .ZN(n983) );
  OAI22_X1 U1729 ( .A1(n1460), .A2(n1210), .B1(n9), .B2(n1209), .ZN(n1001) );
  OAI22_X1 U1730 ( .A1(n1460), .A2(n1211), .B1(n9), .B2(n1210), .ZN(n1002) );
  OAI22_X1 U1731 ( .A1(n23), .A2(n1173), .B1(n22), .B2(n1172), .ZN(n966) );
  OAI22_X1 U1732 ( .A1(n17), .A2(n1192), .B1(n15), .B2(n1191), .ZN(n984) );
  OAI22_X1 U1733 ( .A1(n23), .A2(n1168), .B1(n22), .B2(n1167), .ZN(n961) );
  OAI22_X1 U1734 ( .A1(n17), .A2(n1187), .B1(n15), .B2(n1186), .ZN(n979) );
  OAI22_X1 U1735 ( .A1(n60), .A2(n1035), .B1(n58), .B2(n1034), .ZN(n834) );
  OAI22_X1 U1736 ( .A1(n54), .A2(n1054), .B1(n52), .B2(n1053), .ZN(n852) );
  INV_X1 U1737 ( .A(n464), .ZN(n465) );
  OAI22_X1 U1738 ( .A1(n60), .A2(n1038), .B1(n58), .B2(n1037), .ZN(n837) );
  INV_X1 U1739 ( .A(n802), .ZN(n910) );
  OAI22_X1 U1740 ( .A1(n42), .A2(n1095), .B1(n40), .B2(n1094), .ZN(n891) );
  OAI22_X1 U1741 ( .A1(n54), .A2(n1053), .B1(n52), .B2(n1052), .ZN(n851) );
  INV_X1 U1742 ( .A(n796), .ZN(n870) );
  AOI21_X1 U1743 ( .B1(n48), .B2(n46), .A(n1072), .ZN(n796) );
  OAI22_X1 U1744 ( .A1(n1459), .A2(n1212), .B1(n9), .B2(n1211), .ZN(n1003) );
  OAI22_X1 U1745 ( .A1(n23), .A2(n1174), .B1(n22), .B2(n1173), .ZN(n967) );
  OAI22_X1 U1746 ( .A1(n1411), .A2(n1082), .B1(n45), .B2(n1081), .ZN(n879) );
  OAI22_X1 U1747 ( .A1(n36), .A2(n1120), .B1(n34), .B2(n1119), .ZN(n915) );
  OAI22_X1 U1748 ( .A1(n42), .A2(n1101), .B1(n40), .B2(n1100), .ZN(n897) );
  OAI22_X1 U1749 ( .A1(n48), .A2(n1079), .B1(n46), .B2(n1078), .ZN(n876) );
  OAI22_X1 U1750 ( .A1(n36), .A2(n1117), .B1(n34), .B2(n1116), .ZN(n912) );
  OAI22_X1 U1751 ( .A1(n42), .A2(n1098), .B1(n40), .B2(n1097), .ZN(n894) );
  OAI22_X1 U1752 ( .A1(n5), .A2(n1232), .B1(n1231), .B2(n3), .ZN(n1023) );
  OAI22_X1 U1753 ( .A1(n1459), .A2(n1213), .B1(n9), .B2(n1212), .ZN(n1004) );
  OAI22_X1 U1754 ( .A1(n1383), .A2(n1194), .B1(n15), .B2(n1193), .ZN(n986) );
  AND2_X1 U1755 ( .A1(n1480), .A2(n809), .ZN(n969) );
  OAI22_X1 U1756 ( .A1(n5), .A2(n1233), .B1(n1232), .B2(n3), .ZN(n1024) );
  OAI22_X1 U1757 ( .A1(n1459), .A2(n1214), .B1(n9), .B2(n1213), .ZN(n1005) );
  OAI22_X1 U1758 ( .A1(n1460), .A2(n1205), .B1(n10), .B2(n1204), .ZN(n996) );
  OAI22_X1 U1759 ( .A1(n1411), .A2(n1074), .B1(n46), .B2(n1073), .ZN(n871) );
  OAI22_X1 U1760 ( .A1(n5), .A2(n1230), .B1(n1229), .B2(n3), .ZN(n1021) );
  AND2_X1 U1761 ( .A1(n1480), .A2(n797), .ZN(n889) );
  OAI22_X1 U1762 ( .A1(n35), .A2(n1130), .B1(n33), .B2(n1129), .ZN(n925) );
  OAI22_X1 U1763 ( .A1(n5), .A2(n1225), .B1(n1224), .B2(n4), .ZN(n1016) );
  OAI22_X1 U1764 ( .A1(n29), .A2(n1145), .B1(n27), .B2(n1144), .ZN(n939) );
  OAI22_X1 U1765 ( .A1(n36), .A2(n1126), .B1(n33), .B2(n1125), .ZN(n921) );
  OAI22_X1 U1766 ( .A1(n1383), .A2(n1183), .B1(n16), .B2(n1182), .ZN(n975) );
  OAI22_X1 U1767 ( .A1(n29), .A2(n1152), .B1(n27), .B2(n1151), .ZN(n946) );
  OAI22_X1 U1768 ( .A1(n5), .A2(n1228), .B1(n1227), .B2(n4), .ZN(n1019) );
  OAI22_X1 U1769 ( .A1(n1383), .A2(n1190), .B1(n15), .B2(n1189), .ZN(n982) );
  AND2_X1 U1770 ( .A1(n1451), .A2(n803), .ZN(n929) );
  OAI22_X1 U1771 ( .A1(n1441), .A2(n1229), .B1(n1228), .B2(n3), .ZN(n1020) );
  OAI22_X1 U1772 ( .A1(n23), .A2(n1172), .B1(n21), .B2(n1171), .ZN(n965) );
  OAI22_X1 U1773 ( .A1(n53), .A2(n1065), .B1(n52), .B2(n1064), .ZN(n863) );
  OAI22_X1 U1774 ( .A1(n24), .A2(n1160), .B1(n22), .B2(n1159), .ZN(n953) );
  OAI22_X1 U1775 ( .A1(n29), .A2(n1149), .B1(n27), .B2(n1148), .ZN(n943) );
  OAI22_X1 U1776 ( .A1(n1460), .A2(n1206), .B1(n10), .B2(n1205), .ZN(n997) );
  OAI22_X1 U1777 ( .A1(n41), .A2(n1111), .B1(n40), .B2(n1110), .ZN(n907) );
  OAI22_X1 U1778 ( .A1(n60), .A2(n1039), .B1(n58), .B2(n1038), .ZN(n838) );
  OAI22_X1 U1779 ( .A1(n54), .A2(n1058), .B1(n52), .B2(n1057), .ZN(n856) );
  OAI22_X1 U1780 ( .A1(n42), .A2(n1096), .B1(n40), .B2(n1095), .ZN(n892) );
  OAI22_X1 U1781 ( .A1(n1460), .A2(n1207), .B1(n10), .B2(n1206), .ZN(n998) );
  OAI22_X1 U1782 ( .A1(n1441), .A2(n1226), .B1(n1225), .B2(n4), .ZN(n1017) );
  OAI22_X1 U1783 ( .A1(n23), .A2(n1169), .B1(n21), .B2(n1168), .ZN(n962) );
  OAI22_X1 U1784 ( .A1(n59), .A2(n1042), .B1(n57), .B2(n1041), .ZN(n841) );
  INV_X1 U1785 ( .A(n808), .ZN(n950) );
  AOI21_X1 U1786 ( .B1(n24), .B2(n21), .A(n1156), .ZN(n808) );
  OAI22_X1 U1787 ( .A1(n29), .A2(n1148), .B1(n27), .B2(n1147), .ZN(n942) );
  OAI22_X1 U1788 ( .A1(n1441), .A2(n1224), .B1(n1223), .B2(n4), .ZN(n1015) );
  OAI22_X1 U1789 ( .A1(n1383), .A2(n1186), .B1(n16), .B2(n1185), .ZN(n978) );
  OAI22_X1 U1790 ( .A1(n1441), .A2(n1220), .B1(n1435), .B2(n4), .ZN(n1011) );
  OAI22_X1 U1791 ( .A1(n41), .A2(n1106), .B1(n40), .B2(n1105), .ZN(n902) );
  OAI22_X1 U1792 ( .A1(n24), .A2(n1163), .B1(n21), .B2(n1162), .ZN(n956) );
  OAI22_X1 U1793 ( .A1(n48), .A2(n1075), .B1(n46), .B2(n1074), .ZN(n872) );
  OAI22_X1 U1794 ( .A1(n60), .A2(n1037), .B1(n58), .B2(n1036), .ZN(n836) );
  OAI22_X1 U1795 ( .A1(n54), .A2(n1056), .B1(n52), .B2(n1055), .ZN(n854) );
  OAI22_X1 U1796 ( .A1(n42), .A2(n1097), .B1(n40), .B2(n1096), .ZN(n893) );
  OAI22_X1 U1797 ( .A1(n1411), .A2(n1085), .B1(n45), .B2(n1084), .ZN(n882) );
  OAI22_X1 U1798 ( .A1(n53), .A2(n1066), .B1(n51), .B2(n1065), .ZN(n864) );
  OAI22_X1 U1799 ( .A1(n24), .A2(n1161), .B1(n21), .B2(n1160), .ZN(n954) );
  OAI22_X1 U1800 ( .A1(n42), .A2(n1102), .B1(n40), .B2(n1101), .ZN(n898) );
  INV_X1 U1801 ( .A(n574), .ZN(n575) );
  OAI22_X1 U1802 ( .A1(n1046), .A2(n59), .B1(n1045), .B2(n57), .ZN(n845) );
  OAI22_X1 U1803 ( .A1(n1425), .A2(n18), .B1(n1178), .B2(n16), .ZN(n971) );
  INV_X1 U1804 ( .A(n814), .ZN(n990) );
  OAI22_X1 U1805 ( .A1(n17), .A2(n1189), .B1(n15), .B2(n1188), .ZN(n981) );
  OAI22_X1 U1806 ( .A1(n60), .A2(n1041), .B1(n57), .B2(n1040), .ZN(n840) );
  OAI22_X1 U1807 ( .A1(n54), .A2(n1060), .B1(n52), .B2(n1059), .ZN(n858) );
  AND2_X1 U1808 ( .A1(n1451), .A2(n806), .ZN(n949) );
  OAI22_X1 U1809 ( .A1(n1441), .A2(n1231), .B1(n1230), .B2(n3), .ZN(n1022) );
  OAI22_X1 U1810 ( .A1(n1383), .A2(n1193), .B1(n15), .B2(n1192), .ZN(n985) );
  NAND2_X1 U1811 ( .A1(n787), .A2(n788), .ZN(n400) );
  AND2_X1 U1812 ( .A1(n1480), .A2(n815), .ZN(n1009) );
  INV_X1 U1813 ( .A(n9), .ZN(n815) );
  OAI22_X1 U1814 ( .A1(n1412), .A2(n1439), .B1(n34), .B2(n1122), .ZN(n918) );
  OAI22_X1 U1815 ( .A1(n30), .A2(n1142), .B1(n28), .B2(n1141), .ZN(n936) );
  INV_X1 U1816 ( .A(n608), .ZN(n609) );
  OR2_X1 U1817 ( .A1(n1480), .A2(n1290), .ZN(n1050) );
  OR2_X1 U1818 ( .A1(n1480), .A2(n1297), .ZN(n1197) );
  OR2_X1 U1819 ( .A1(n1480), .A2(n1296), .ZN(n1176) );
  OR2_X1 U1820 ( .A1(n1451), .A2(n1293), .ZN(n1113) );
  OR2_X1 U1821 ( .A1(n1481), .A2(n1292), .ZN(n1092) );
  OR2_X1 U1822 ( .A1(n1481), .A2(n1294), .ZN(n1134) );
  OAI22_X1 U1823 ( .A1(n1048), .A2(n59), .B1(n1047), .B2(n57), .ZN(n847) );
  OAI22_X1 U1824 ( .A1(n1124), .A2(n35), .B1(n1439), .B2(n33), .ZN(n919) );
  INV_X1 U1825 ( .A(n817), .ZN(n1010) );
  OAI22_X1 U1826 ( .A1(n60), .A2(n1044), .B1(n57), .B2(n1043), .ZN(n843) );
  INV_X1 U1827 ( .A(n811), .ZN(n970) );
  AOI21_X1 U1828 ( .B1(n1383), .B2(n16), .A(n1177), .ZN(n811) );
  INV_X1 U1829 ( .A(n57), .ZN(n791) );
  INV_X1 U1830 ( .A(n33), .ZN(n803) );
  INV_X1 U1831 ( .A(n39), .ZN(n800) );
  INV_X1 U1832 ( .A(n15), .ZN(n812) );
  INV_X1 U1833 ( .A(n21), .ZN(n809) );
  INV_X1 U1834 ( .A(n27), .ZN(n806) );
  INV_X1 U1835 ( .A(n45), .ZN(n797) );
  OAI22_X1 U1836 ( .A1(n1441), .A2(n1236), .B1(n1235), .B2(n3), .ZN(n1027) );
  OAI22_X1 U1837 ( .A1(n1460), .A2(n1217), .B1(n9), .B2(n1216), .ZN(n1008) );
  XNOR2_X1 U1838 ( .A(n1385), .B(n1451), .ZN(n1217) );
  OAI22_X1 U1839 ( .A1(n1459), .A2(n1298), .B1(n1218), .B2(n10), .ZN(n828) );
  OR2_X1 U1840 ( .A1(n1481), .A2(n1298), .ZN(n1218) );
  INV_X1 U1841 ( .A(n7), .ZN(n1298) );
  OAI22_X1 U1842 ( .A1(n1441), .A2(n1299), .B1(n1239), .B2(n4), .ZN(n829) );
  OR2_X1 U1843 ( .A1(n1451), .A2(n1299), .ZN(n1239) );
  INV_X1 U1844 ( .A(n1442), .ZN(n1299) );
  OAI22_X1 U1845 ( .A1(n1441), .A2(n1238), .B1(n1237), .B2(n3), .ZN(n1029) );
  OAI22_X1 U1846 ( .A1(n48), .A2(n1091), .B1(n45), .B2(n1090), .ZN(n888) );
  OAI22_X1 U1847 ( .A1(n48), .A2(n1292), .B1(n1092), .B2(n46), .ZN(n822) );
  XNOR2_X1 U1848 ( .A(n1447), .B(n1480), .ZN(n1091) );
  OAI22_X1 U1849 ( .A1(n36), .A2(n1133), .B1(n33), .B2(n1132), .ZN(n928) );
  OAI22_X1 U1850 ( .A1(n1412), .A2(n1294), .B1(n1134), .B2(n34), .ZN(n824) );
  XNOR2_X1 U1851 ( .A(n1448), .B(n1481), .ZN(n1133) );
  XNOR2_X1 U1852 ( .A(n37), .B(n1258), .ZN(n1111) );
  XNOR2_X1 U1853 ( .A(n7), .B(n1246), .ZN(n1204) );
  XNOR2_X1 U1854 ( .A(n7), .B(n1247), .ZN(n1205) );
  XNOR2_X1 U1855 ( .A(n1436), .B(n1241), .ZN(n1094) );
  XNOR2_X1 U1856 ( .A(n1256), .B(n37), .ZN(n1109) );
  XNOR2_X1 U1857 ( .A(n31), .B(n1254), .ZN(n1128) );
  XNOR2_X1 U1858 ( .A(n37), .B(n1257), .ZN(n1110) );
  XNOR2_X1 U1859 ( .A(n31), .B(n1255), .ZN(n1129) );
  XNOR2_X1 U1860 ( .A(n1445), .B(n1246), .ZN(n1183) );
  XNOR2_X1 U1861 ( .A(n13), .B(n1248), .ZN(n1185) );
  XNOR2_X1 U1862 ( .A(n13), .B(n1247), .ZN(n1184) );
  XNOR2_X1 U1863 ( .A(n37), .B(n1255), .ZN(n1108) );
  XNOR2_X1 U1864 ( .A(n31), .B(n1253), .ZN(n1127) );
  XNOR2_X1 U1865 ( .A(n1436), .B(n1242), .ZN(n1095) );
  XNOR2_X1 U1866 ( .A(n37), .B(n1254), .ZN(n1107) );
  XNOR2_X1 U1867 ( .A(n1448), .B(n1252), .ZN(n1126) );
  XNOR2_X1 U1868 ( .A(n7), .B(n1245), .ZN(n1203) );
  XNOR2_X1 U1869 ( .A(n13), .B(n1243), .ZN(n1180) );
  XNOR2_X1 U1870 ( .A(n13), .B(n1245), .ZN(n1182) );
  XNOR2_X1 U1871 ( .A(n1448), .B(n1251), .ZN(n1125) );
  XNOR2_X1 U1872 ( .A(n7), .B(n1244), .ZN(n1202) );
  XNOR2_X1 U1873 ( .A(n1250), .B(n31), .ZN(n1124) );
  XNOR2_X1 U1874 ( .A(n1445), .B(n1244), .ZN(n1181) );
  XNOR2_X1 U1875 ( .A(n7), .B(n1248), .ZN(n1206) );
  XNOR2_X1 U1876 ( .A(n1448), .B(n1256), .ZN(n1130) );
  XNOR2_X1 U1877 ( .A(n1448), .B(n1248), .ZN(n1122) );
  XNOR2_X1 U1878 ( .A(n1445), .B(n1249), .ZN(n1186) );
  XNOR2_X1 U1879 ( .A(n1436), .B(n1243), .ZN(n1096) );
  XNOR2_X1 U1880 ( .A(n7), .B(n1243), .ZN(n1201) );
  XNOR2_X1 U1881 ( .A(n37), .B(n1244), .ZN(n1097) );
  XNOR2_X1 U1882 ( .A(n7), .B(n1242), .ZN(n1200) );
  XNOR2_X1 U1883 ( .A(n37), .B(n1251), .ZN(n1104) );
  XNOR2_X1 U1884 ( .A(n1448), .B(n1247), .ZN(n1121) );
  XNOR2_X1 U1885 ( .A(n37), .B(n1252), .ZN(n1105) );
  XNOR2_X1 U1886 ( .A(n37), .B(n1253), .ZN(n1106) );
  XNOR2_X1 U1887 ( .A(n1448), .B(n1241), .ZN(n1115) );
  XNOR2_X1 U1888 ( .A(n1445), .B(n1251), .ZN(n1188) );
  XNOR2_X1 U1889 ( .A(n37), .B(n1246), .ZN(n1099) );
  XNOR2_X1 U1890 ( .A(n13), .B(n1242), .ZN(n1179) );
  XNOR2_X1 U1891 ( .A(n37), .B(n1248), .ZN(n1101) );
  XNOR2_X1 U1892 ( .A(n7), .B(n1241), .ZN(n1199) );
  XNOR2_X1 U1893 ( .A(n37), .B(n1245), .ZN(n1098) );
  XNOR2_X1 U1894 ( .A(n13), .B(n1241), .ZN(n1178) );
  XNOR2_X1 U1895 ( .A(n37), .B(n1250), .ZN(n1103) );
  XNOR2_X1 U1896 ( .A(n37), .B(n1249), .ZN(n1102) );
  XNOR2_X1 U1897 ( .A(n1448), .B(n1244), .ZN(n1118) );
  XNOR2_X1 U1898 ( .A(n31), .B(n1243), .ZN(n1117) );
  XNOR2_X1 U1899 ( .A(n1448), .B(n1245), .ZN(n1119) );
  XNOR2_X1 U1900 ( .A(n37), .B(n1247), .ZN(n1100) );
  XNOR2_X1 U1901 ( .A(n1448), .B(n1257), .ZN(n1131) );
  XNOR2_X1 U1902 ( .A(n1445), .B(n1252), .ZN(n1189) );
  XNOR2_X1 U1903 ( .A(n1448), .B(n1242), .ZN(n1116) );
  XNOR2_X1 U1904 ( .A(n1250), .B(n1445), .ZN(n1187) );
  XNOR2_X1 U1905 ( .A(n1448), .B(n1246), .ZN(n1120) );
  XNOR2_X1 U1906 ( .A(n7), .B(n1249), .ZN(n1207) );
  XNOR2_X1 U1907 ( .A(n1385), .B(n1251), .ZN(n1209) );
  XNOR2_X1 U1908 ( .A(n7), .B(n1250), .ZN(n1208) );
  XNOR2_X1 U1909 ( .A(n1445), .B(n1253), .ZN(n1190) );
  XNOR2_X1 U1910 ( .A(n1448), .B(n1258), .ZN(n1132) );
  XNOR2_X1 U1911 ( .A(n1445), .B(n1254), .ZN(n1191) );
  XNOR2_X1 U1912 ( .A(n7), .B(n1252), .ZN(n1210) );
  XNOR2_X1 U1913 ( .A(n7), .B(n1253), .ZN(n1211) );
  XNOR2_X1 U1914 ( .A(n1445), .B(n1388), .ZN(n1192) );
  XNOR2_X1 U1915 ( .A(n7), .B(n1258), .ZN(n1216) );
  XNOR2_X1 U1916 ( .A(n7), .B(n1257), .ZN(n1215) );
  XNOR2_X1 U1917 ( .A(n7), .B(n1389), .ZN(n1213) );
  XNOR2_X1 U1918 ( .A(n7), .B(n1256), .ZN(n1214) );
  XNOR2_X1 U1919 ( .A(n1385), .B(n1254), .ZN(n1212) );
  XNOR2_X1 U1920 ( .A(n1445), .B(n1258), .ZN(n1195) );
  XNOR2_X1 U1921 ( .A(n1445), .B(n1256), .ZN(n1193) );
  XNOR2_X1 U1922 ( .A(n13), .B(n1444), .ZN(n1194) );
  XNOR2_X1 U1923 ( .A(n1429), .B(n1244), .ZN(n1034) );
  XNOR2_X1 U1924 ( .A(n1447), .B(n1241), .ZN(n1073) );
  XNOR2_X1 U1925 ( .A(n1428), .B(n1243), .ZN(n1033) );
  XNOR2_X1 U1926 ( .A(n1447), .B(n1242), .ZN(n1074) );
  XNOR2_X1 U1927 ( .A(n1428), .B(n1245), .ZN(n1035) );
  XNOR2_X1 U1928 ( .A(n1428), .B(n1246), .ZN(n1036) );
  XNOR2_X1 U1929 ( .A(n19), .B(n1250), .ZN(n1166) );
  XNOR2_X1 U1930 ( .A(n43), .B(n1258), .ZN(n1090) );
  XNOR2_X1 U1931 ( .A(n19), .B(n1248), .ZN(n1164) );
  XNOR2_X1 U1932 ( .A(n19), .B(n1249), .ZN(n1165) );
  XNOR2_X1 U1933 ( .A(n43), .B(n1257), .ZN(n1089) );
  XNOR2_X1 U1934 ( .A(n1429), .B(n1247), .ZN(n1037) );
  XNOR2_X1 U1935 ( .A(n43), .B(n1256), .ZN(n1088) );
  XNOR2_X1 U1936 ( .A(n19), .B(n1247), .ZN(n1163) );
  XNOR2_X1 U1937 ( .A(n1428), .B(n1248), .ZN(n1038) );
  XNOR2_X1 U1938 ( .A(n1447), .B(n1244), .ZN(n1076) );
  XNOR2_X1 U1939 ( .A(n19), .B(n1245), .ZN(n1161) );
  XNOR2_X1 U1940 ( .A(n1429), .B(n1242), .ZN(n1032) );
  XNOR2_X1 U1941 ( .A(n19), .B(n1251), .ZN(n1167) );
  XNOR2_X1 U1942 ( .A(n1429), .B(n1258), .ZN(n1048) );
  XNOR2_X1 U1943 ( .A(n1447), .B(n1243), .ZN(n1075) );
  XNOR2_X1 U1944 ( .A(n1257), .B(n1429), .ZN(n1047) );
  XNOR2_X1 U1945 ( .A(n19), .B(n1246), .ZN(n1162) );
  XNOR2_X1 U1946 ( .A(n1447), .B(n1253), .ZN(n1085) );
  XNOR2_X1 U1947 ( .A(n43), .B(n1254), .ZN(n1086) );
  XNOR2_X1 U1948 ( .A(n1447), .B(n1245), .ZN(n1077) );
  XNOR2_X1 U1949 ( .A(n19), .B(n1241), .ZN(n1157) );
  XNOR2_X1 U1950 ( .A(n1428), .B(n1256), .ZN(n1046) );
  XNOR2_X1 U1951 ( .A(n1447), .B(n1247), .ZN(n1079) );
  XNOR2_X1 U1952 ( .A(n19), .B(n1244), .ZN(n1160) );
  XNOR2_X1 U1953 ( .A(n1447), .B(n1248), .ZN(n1080) );
  XNOR2_X1 U1954 ( .A(n1429), .B(n1251), .ZN(n1041) );
  XNOR2_X1 U1955 ( .A(n1428), .B(n1252), .ZN(n1042) );
  XNOR2_X1 U1956 ( .A(n1429), .B(n1389), .ZN(n1045) );
  XNOR2_X1 U1957 ( .A(n1429), .B(n1249), .ZN(n1039) );
  XNOR2_X1 U1958 ( .A(n1447), .B(n1252), .ZN(n1084) );
  XNOR2_X1 U1959 ( .A(n1428), .B(n1254), .ZN(n1044) );
  XNOR2_X1 U1960 ( .A(n1429), .B(n1253), .ZN(n1043) );
  XNOR2_X1 U1961 ( .A(n19), .B(n1243), .ZN(n1159) );
  XNOR2_X1 U1962 ( .A(n1428), .B(n1250), .ZN(n1040) );
  XNOR2_X1 U1963 ( .A(n1447), .B(n1250), .ZN(n1082) );
  XNOR2_X1 U1964 ( .A(n19), .B(n1242), .ZN(n1158) );
  XNOR2_X1 U1965 ( .A(n1447), .B(n1246), .ZN(n1078) );
  XNOR2_X1 U1966 ( .A(n1447), .B(n1251), .ZN(n1083) );
  XNOR2_X1 U1967 ( .A(n1447), .B(n1249), .ZN(n1081) );
  XNOR2_X1 U1968 ( .A(n19), .B(n1253), .ZN(n1169) );
  XNOR2_X1 U1969 ( .A(n19), .B(n1252), .ZN(n1168) );
  XNOR2_X1 U1970 ( .A(n19), .B(n1388), .ZN(n1171) );
  XNOR2_X1 U1971 ( .A(n19), .B(n1254), .ZN(n1170) );
  XNOR2_X1 U1972 ( .A(n19), .B(n1256), .ZN(n1172) );
  XNOR2_X1 U1973 ( .A(n19), .B(n1257), .ZN(n1173) );
  XNOR2_X1 U1974 ( .A(n19), .B(n1258), .ZN(n1174) );
  XNOR2_X1 U1975 ( .A(n1429), .B(n1241), .ZN(n1031) );
  BUF_X1 U1976 ( .A(n1283), .Z(n39) );
  XNOR2_X1 U1977 ( .A(n1436), .B(n1408), .ZN(n1093) );
  XNOR2_X1 U1978 ( .A(n1240), .B(n1448), .ZN(n1114) );
  XNOR2_X1 U1979 ( .A(n1445), .B(n1240), .ZN(n1177) );
  XNOR2_X1 U1980 ( .A(n1240), .B(n7), .ZN(n1198) );
  XNOR2_X1 U1981 ( .A(n1447), .B(n1467), .ZN(n1072) );
  XNOR2_X1 U1982 ( .A(n19), .B(n1240), .ZN(n1156) );
  XNOR2_X1 U1983 ( .A(n1428), .B(n1467), .ZN(n1030) );
  BUF_X1 U1984 ( .A(n1283), .Z(n40) );
  BUF_X2 U1985 ( .A(n1270), .Z(n60) );
  BUF_X2 U1986 ( .A(n1274), .Z(n36) );
  BUF_X2 U1987 ( .A(n1275), .Z(n30) );
  BUF_X2 U1988 ( .A(n1272), .Z(n48) );
  OAI22_X1 U1989 ( .A1(n1383), .A2(n1196), .B1(n15), .B2(n1195), .ZN(n988) );
  OAI22_X1 U1990 ( .A1(n1383), .A2(n1297), .B1(n1197), .B2(n16), .ZN(n827) );
  XNOR2_X1 U1991 ( .A(n1445), .B(n1451), .ZN(n1196) );
  OAI22_X1 U1992 ( .A1(n1112), .A2(n41), .B1(n39), .B2(n1111), .ZN(n908) );
  OAI22_X1 U1993 ( .A1(n42), .A2(n1293), .B1(n1113), .B2(n39), .ZN(n823) );
  XNOR2_X1 U1994 ( .A(n37), .B(n1451), .ZN(n1112) );
  OAI22_X1 U1995 ( .A1(n59), .A2(n1049), .B1(n57), .B2(n1438), .ZN(n848) );
  OAI22_X1 U1996 ( .A1(n60), .A2(n1290), .B1(n1050), .B2(n58), .ZN(n820) );
  XNOR2_X1 U1997 ( .A(n1429), .B(n1481), .ZN(n1049) );
  OAI22_X1 U1998 ( .A1(n23), .A2(n1175), .B1(n22), .B2(n1174), .ZN(n968) );
  OAI22_X1 U1999 ( .A1(n24), .A2(n1296), .B1(n1176), .B2(n22), .ZN(n826) );
  XNOR2_X1 U2000 ( .A(n19), .B(n1481), .ZN(n1175) );
  INV_X1 U2001 ( .A(n49), .ZN(n1291) );
  INV_X1 U2002 ( .A(n1440), .ZN(n1295) );
  BUF_X2 U2003 ( .A(n1271), .Z(n53) );
  INV_X1 U2004 ( .A(n37), .ZN(n1293) );
  INV_X1 U2005 ( .A(n1448), .ZN(n1294) );
  INV_X1 U2006 ( .A(n1445), .ZN(n1297) );
  INV_X1 U2007 ( .A(n43), .ZN(n1292) );
  INV_X1 U2008 ( .A(n19), .ZN(n1296) );
  INV_X1 U2009 ( .A(n1429), .ZN(n1290) );
  BUF_X1 U2010 ( .A(n1289), .Z(n3) );
  BUF_X1 U2011 ( .A(n1289), .Z(n4) );
  XNOR2_X1 U2012 ( .A(a[11]), .B(a[12]), .ZN(n1283) );
  XNOR2_X1 U2013 ( .A(a[6]), .B(a[5]), .ZN(n1286) );
  XNOR2_X1 U2014 ( .A(a[4]), .B(a[3]), .ZN(n1287) );
  BUF_X4 U2015 ( .A(a[3]), .Z(n7) );
  BUF_X4 U2016 ( .A(a[7]), .Z(n19) );
  XNOR2_X1 U2017 ( .A(a[14]), .B(a[13]), .ZN(n1282) );
  NAND2_X1 U2018 ( .A1(n1265), .A2(n1285), .ZN(n1275) );
  XNOR2_X1 U2019 ( .A(a[8]), .B(a[7]), .ZN(n1285) );
  NAND2_X1 U2020 ( .A1(n1261), .A2(n1281), .ZN(n1271) );
  XNOR2_X1 U2021 ( .A(a[15]), .B(a[16]), .ZN(n1281) );
  OAI21_X1 U2022 ( .B1(n1461), .B2(n304), .A(n297), .ZN(n295) );
  INV_X1 U2023 ( .A(n1426), .ZN(n426) );
  NOR2_X1 U2024 ( .A1(n577), .A2(n592), .ZN(n296) );
  AOI21_X1 U2025 ( .B1(n349), .B2(n1404), .A(n344), .ZN(n342) );
  NOR2_X1 U2026 ( .A1(n296), .A2(n303), .ZN(n294) );
  INV_X1 U2027 ( .A(n1434), .ZN(n302) );
  XNOR2_X1 U2028 ( .A(n1440), .B(n1240), .ZN(n1135) );
  XNOR2_X1 U2029 ( .A(n1440), .B(n1244), .ZN(n1139) );
  XNOR2_X1 U2030 ( .A(n25), .B(n1241), .ZN(n1136) );
  XNOR2_X1 U2031 ( .A(n1440), .B(n1246), .ZN(n1141) );
  XNOR2_X1 U2032 ( .A(n1440), .B(n1480), .ZN(n1154) );
  XNOR2_X1 U2033 ( .A(n1440), .B(n1254), .ZN(n1149) );
  XNOR2_X1 U2034 ( .A(n1440), .B(n1250), .ZN(n1145) );
  XNOR2_X1 U2035 ( .A(n1440), .B(n1245), .ZN(n1140) );
  XNOR2_X1 U2036 ( .A(n25), .B(n1388), .ZN(n1150) );
  XNOR2_X1 U2037 ( .A(n1440), .B(n1257), .ZN(n1152) );
  XNOR2_X1 U2038 ( .A(n1440), .B(n1243), .ZN(n1138) );
  XNOR2_X1 U2039 ( .A(n25), .B(n1256), .ZN(n1151) );
  XNOR2_X1 U2040 ( .A(n1440), .B(n1258), .ZN(n1153) );
  XNOR2_X1 U2041 ( .A(n25), .B(n1251), .ZN(n1146) );
  XNOR2_X1 U2042 ( .A(n25), .B(n1242), .ZN(n1137) );
  XNOR2_X1 U2043 ( .A(n1440), .B(n1247), .ZN(n1142) );
  XNOR2_X1 U2044 ( .A(n25), .B(n1249), .ZN(n1144) );
  XNOR2_X1 U2045 ( .A(n25), .B(n1248), .ZN(n1143) );
  XNOR2_X1 U2046 ( .A(n1440), .B(n1253), .ZN(n1148) );
  XNOR2_X1 U2047 ( .A(n1440), .B(n1252), .ZN(n1147) );
  XNOR2_X1 U2048 ( .A(a[10]), .B(a[9]), .ZN(n1284) );
  OAI21_X1 U2049 ( .B1(n341), .B2(n358), .A(n342), .ZN(n340) );
  INV_X1 U2050 ( .A(n518), .ZN(n519) );
  NAND2_X1 U2051 ( .A1(n509), .A2(n520), .ZN(n256) );
  INV_X1 U2052 ( .A(n65), .ZN(n246) );
  AOI21_X1 U2053 ( .B1(n340), .B2(n321), .A(n322), .ZN(n320) );
  OAI21_X1 U2054 ( .B1(n327), .B2(n323), .A(n324), .ZN(n322) );
  AOI21_X1 U2055 ( .B1(n357), .B2(n435), .A(n354), .ZN(n352) );
  XOR2_X1 U2056 ( .A(n157), .B(n70), .Z(product[35]) );
  NOR2_X1 U2057 ( .A1(n312), .A2(n317), .ZN(n310) );
  NAND2_X1 U2058 ( .A1(n294), .A2(n310), .ZN(n292) );
  INV_X1 U2059 ( .A(n310), .ZN(n308) );
  AOI21_X1 U2060 ( .B1(n283), .B2(n249), .A(n250), .ZN(n248) );
  BUF_X2 U2061 ( .A(n291), .Z(n63) );
  AOI21_X1 U2062 ( .B1(n1432), .B2(n311), .A(n295), .ZN(n293) );
  OAI21_X1 U2063 ( .B1(n312), .B2(n318), .A(n313), .ZN(n311) );
  INV_X1 U2064 ( .A(n1454), .ZN(n319) );
  OAI21_X1 U2065 ( .B1(n320), .B2(n292), .A(n293), .ZN(n291) );
  XNOR2_X1 U2066 ( .A(n49), .B(n1247), .ZN(n1058) );
  XNOR2_X1 U2067 ( .A(n49), .B(n1243), .ZN(n1054) );
  XNOR2_X1 U2068 ( .A(n49), .B(n1246), .ZN(n1057) );
  XNOR2_X1 U2069 ( .A(n49), .B(n1242), .ZN(n1053) );
  XNOR2_X1 U2070 ( .A(n49), .B(n1245), .ZN(n1056) );
  XNOR2_X1 U2071 ( .A(n49), .B(n1244), .ZN(n1055) );
  XNOR2_X1 U2072 ( .A(n49), .B(n1248), .ZN(n1059) );
  XNOR2_X1 U2073 ( .A(n49), .B(n1253), .ZN(n1064) );
  XNOR2_X1 U2074 ( .A(n49), .B(n1252), .ZN(n1063) );
  XNOR2_X1 U2075 ( .A(n49), .B(n1249), .ZN(n1060) );
  XNOR2_X1 U2076 ( .A(n49), .B(n1251), .ZN(n1062) );
  XNOR2_X1 U2077 ( .A(n49), .B(n1250), .ZN(n1061) );
  XNOR2_X1 U2078 ( .A(n49), .B(n1451), .ZN(n1070) );
  XNOR2_X1 U2079 ( .A(n49), .B(n1254), .ZN(n1065) );
  XNOR2_X1 U2080 ( .A(n49), .B(n1389), .ZN(n1066) );
  XNOR2_X1 U2081 ( .A(n49), .B(n1257), .ZN(n1068) );
  XNOR2_X1 U2082 ( .A(n49), .B(n1256), .ZN(n1067) );
  XNOR2_X1 U2083 ( .A(n49), .B(n1258), .ZN(n1069) );
  XNOR2_X1 U2084 ( .A(n49), .B(n1241), .ZN(n1052) );
  XNOR2_X1 U2085 ( .A(n49), .B(n1467), .ZN(n1051) );
  XNOR2_X1 U2086 ( .A(a[18]), .B(a[17]), .ZN(n1280) );
  BUF_X4 U2087 ( .A(a[17]), .Z(n49) );
  AOI21_X1 U2088 ( .B1(n63), .B2(n169), .A(n170), .ZN(n168) );
  OAI21_X1 U2089 ( .B1(n230), .B2(n220), .A(n221), .ZN(n219) );
  AOI21_X1 U2090 ( .B1(n1424), .B2(n115), .A(n116), .ZN(n114) );
  OAI21_X1 U2091 ( .B1(n251), .B2(n276), .A(n252), .ZN(n250) );
  AOI21_X1 U2092 ( .B1(n63), .B2(n128), .A(n129), .ZN(n127) );
  AOI21_X1 U2093 ( .B1(n63), .B2(n199), .A(n200), .ZN(n198) );
  AOI21_X1 U2094 ( .B1(n63), .B2(n158), .A(n159), .ZN(n157) );
  XNOR2_X1 U2095 ( .A(n63), .B(n82), .ZN(product[23]) );
  AOI21_X1 U2096 ( .B1(n64), .B2(n258), .A(n259), .ZN(n257) );
  AOI21_X1 U2097 ( .B1(n64), .B2(n287), .A(n288), .ZN(n286) );
  AOI21_X1 U2098 ( .B1(n63), .B2(n245), .A(n246), .ZN(n244) );
  AOI21_X1 U2099 ( .B1(n64), .B2(n269), .A(n270), .ZN(n268) );
  AOI21_X1 U2100 ( .B1(n64), .B2(n282), .A(n279), .ZN(n277) );
  AOI21_X1 U2101 ( .B1(n63), .B2(n223), .A(n224), .ZN(n222) );
  NAND2_X1 U2102 ( .A1(n679), .A2(n692), .ZN(n338) );
  AOI21_X1 U2103 ( .B1(n64), .B2(n210), .A(n211), .ZN(n209) );
  NOR2_X1 U2104 ( .A1(n1433), .A2(n108), .ZN(n106) );
  NOR2_X1 U2105 ( .A1(n1433), .A2(n117), .ZN(n115) );
  NOR2_X1 U2106 ( .A1(n1433), .A2(n145), .ZN(n143) );
  NOR2_X1 U2107 ( .A1(n1433), .A2(n130), .ZN(n128) );
  NOR2_X1 U2108 ( .A1(n1433), .A2(n201), .ZN(n199) );
  NOR2_X1 U2109 ( .A1(n1433), .A2(n171), .ZN(n169) );
  NOR2_X1 U2110 ( .A1(n1433), .A2(n184), .ZN(n182) );
  NOR2_X1 U2111 ( .A1(n1433), .A2(n160), .ZN(n158) );
  NOR2_X1 U2112 ( .A1(n66), .A2(n216), .ZN(n210) );
  NOR2_X1 U2113 ( .A1(n66), .A2(n225), .ZN(n223) );
  NOR2_X1 U2114 ( .A1(n66), .A2(n242), .ZN(n232) );
  NAND2_X1 U2115 ( .A1(n1260), .A2(n1280), .ZN(n1270) );
  NAND2_X1 U2116 ( .A1(n1264), .A2(n1284), .ZN(n1274) );
  AOI21_X1 U2117 ( .B1(n63), .B2(n143), .A(n144), .ZN(n142) );
  INV_X1 U2118 ( .A(n358), .ZN(n357) );
  XNOR2_X1 U2119 ( .A(n1442), .B(n1248), .ZN(n1227) );
  XNOR2_X1 U2120 ( .A(n1442), .B(n1251), .ZN(n1230) );
  XNOR2_X1 U2121 ( .A(n1442), .B(n1252), .ZN(n1231) );
  XNOR2_X1 U2122 ( .A(n1442), .B(n1247), .ZN(n1226) );
  XNOR2_X1 U2123 ( .A(n1), .B(n1246), .ZN(n1225) );
  XNOR2_X1 U2124 ( .A(n1), .B(n1245), .ZN(n1224) );
  XNOR2_X1 U2125 ( .A(n1), .B(n1242), .ZN(n1221) );
  XNOR2_X1 U2126 ( .A(n1442), .B(n1389), .ZN(n1234) );
  XNOR2_X1 U2127 ( .A(n1442), .B(n1254), .ZN(n1233) );
  XNOR2_X1 U2128 ( .A(n1), .B(n1241), .ZN(n1220) );
  XNOR2_X1 U2129 ( .A(n1), .B(n1244), .ZN(n1223) );
  XNOR2_X1 U2130 ( .A(n1), .B(n1253), .ZN(n1232) );
  XNOR2_X1 U2131 ( .A(n1442), .B(n1480), .ZN(n1238) );
  XNOR2_X1 U2132 ( .A(n1), .B(n1243), .ZN(n1222) );
  XNOR2_X1 U2133 ( .A(n1), .B(n1250), .ZN(n1229) );
  XNOR2_X1 U2134 ( .A(n1), .B(n1249), .ZN(n1228) );
  XNOR2_X1 U2135 ( .A(n1442), .B(n1258), .ZN(n1237) );
  XNOR2_X1 U2136 ( .A(n1442), .B(n1257), .ZN(n1236) );
  XNOR2_X1 U2137 ( .A(n1442), .B(n1256), .ZN(n1235) );
  XNOR2_X1 U2138 ( .A(n1), .B(n1240), .ZN(n1219) );
  NAND2_X1 U2139 ( .A1(n473), .A2(n480), .ZN(n208) );
  AOI21_X1 U2140 ( .B1(n299), .B2(n319), .A(n300), .ZN(n298) );
  XNOR2_X1 U2141 ( .A(n319), .B(n86), .ZN(product[19]) );
  AOI21_X1 U2142 ( .B1(n319), .B2(n306), .A(n307), .ZN(n305) );
  AOI21_X1 U2143 ( .B1(n319), .B2(n315), .A(n316), .ZN(n314) );
  NAND2_X1 U2144 ( .A1(n1262), .A2(n1282), .ZN(n1272) );
  XOR2_X1 U2145 ( .A(n388), .B(n98), .Z(product[7]) );
  INV_X1 U2146 ( .A(n367), .ZN(n366) );
  AOI21_X1 U2147 ( .B1(n367), .B2(n359), .A(n360), .ZN(n358) );
  OAI21_X1 U2148 ( .B1(n1458), .B2(n108), .A(n109), .ZN(n107) );
  OAI21_X1 U2149 ( .B1(n65), .B2(n117), .A(n118), .ZN(n116) );
  OAI21_X1 U2150 ( .B1(n1458), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U2151 ( .B1(n1458), .B2(n145), .A(n146), .ZN(n144) );
  OAI21_X1 U2152 ( .B1(n1458), .B2(n201), .A(n202), .ZN(n200) );
  OAI21_X1 U2153 ( .B1(n1458), .B2(n171), .A(n172), .ZN(n170) );
  OAI21_X1 U2154 ( .B1(n65), .B2(n216), .A(n217), .ZN(n211) );
  OAI21_X1 U2155 ( .B1(n1458), .B2(n160), .A(n161), .ZN(n159) );
  OAI21_X1 U2156 ( .B1(n1458), .B2(n184), .A(n185), .ZN(n183) );
  OAI21_X1 U2157 ( .B1(n65), .B2(n225), .A(n226), .ZN(n224) );
  OAI21_X1 U2158 ( .B1(n65), .B2(n242), .A(n243), .ZN(n233) );
  OAI22_X1 U2159 ( .A1(n54), .A2(n1052), .B1(n52), .B2(n1051), .ZN(n454) );
  BUF_X2 U2160 ( .A(n1271), .Z(n54) );
  NAND2_X1 U2161 ( .A1(n1028), .A2(n1009), .ZN(n407) );
  AOI21_X1 U2162 ( .B1(n64), .B2(n232), .A(n233), .ZN(n231) );
  NAND2_X1 U2163 ( .A1(n282), .A2(n249), .ZN(n247) );
  OAI21_X1 U2164 ( .B1(n361), .B2(n365), .A(n362), .ZN(n360) );
  NOR2_X1 U2165 ( .A1(n361), .A2(n364), .ZN(n359) );
  XOR2_X1 U2166 ( .A(a[11]), .B(a[10]), .Z(n1264) );
  AOI21_X1 U2167 ( .B1(n357), .B2(n348), .A(n349), .ZN(n347) );
  NAND2_X1 U2168 ( .A1(n348), .A2(n1404), .ZN(n341) );
  NOR2_X1 U2169 ( .A1(n350), .A2(n355), .ZN(n348) );
  XOR2_X1 U2170 ( .A(a[18]), .B(a[19]), .Z(n1260) );
  XOR2_X1 U2171 ( .A(a[15]), .B(a[14]), .Z(n1262) );
  XOR2_X1 U2172 ( .A(a[8]), .B(a[9]), .Z(n1265) );
  XOR2_X1 U2173 ( .A(a[12]), .B(a[13]), .Z(n1263) );
  XOR2_X1 U2174 ( .A(a[2]), .B(a[3]), .Z(n1268) );
  XOR2_X1 U2175 ( .A(a[6]), .B(a[7]), .Z(n1266) );
  XOR2_X1 U2176 ( .A(a[16]), .B(a[17]), .Z(n1261) );
  XNOR2_X1 U2177 ( .A(n99), .B(n393), .ZN(product[6]) );
  XOR2_X1 U2178 ( .A(a[4]), .B(a[5]), .Z(n1267) );
  NOR2_X1 U2179 ( .A1(n289), .A2(n284), .ZN(n282) );
  XOR2_X1 U2180 ( .A(a[0]), .B(a[1]), .Z(n1269) );
endmodule


module datapath_DW01_add_8 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n43, n44, n46, n48, n50, n52, n53, n54, n55,
         n56, n57, n59, n61, n62, n63, n64, n65, n68, n70, n71, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n94, n95, n96, n97, n98, n99, n100, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n125, n126, n127, n128, n129,
         n130, n131, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n179, n180,
         n181, n182, n183, n184, n185, n186, n188, n189, n190, n191, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n246, n247, n248, n249, n252, n253, n254, n255, n256,
         n257, n258, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n275, n276, n277, n278, n279, n280,
         n283, n284, n285, n286, n287, n289, n290, n291, n292, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n353, n358,
         n360, n361, n366, n368, n370, n372, n374, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n570, n571;

  BUF_X1 U437 ( .A(n105), .Z(n520) );
  NOR2_X1 U438 ( .A1(B[33]), .A2(A[33]), .ZN(n98) );
  CLKBUF_X1 U439 ( .A(n115), .Z(n521) );
  CLKBUF_X1 U440 ( .A(n219), .Z(n522) );
  CLKBUF_X1 U441 ( .A(n55), .Z(n523) );
  NOR2_X2 U442 ( .A1(B[23]), .A2(A[23]), .ZN(n202) );
  AND2_X1 U443 ( .A1(n54), .A2(n530), .ZN(n524) );
  NOR2_X1 U444 ( .A1(n147), .A2(n138), .ZN(n525) );
  CLKBUF_X1 U445 ( .A(B[29]), .Z(n526) );
  NOR2_X1 U446 ( .A1(B[35]), .A2(A[35]), .ZN(n82) );
  NOR2_X1 U447 ( .A1(n189), .A2(n182), .ZN(n527) );
  NOR2_X1 U448 ( .A1(B[29]), .A2(A[29]), .ZN(n528) );
  OR2_X1 U449 ( .A1(A[37]), .A2(B[37]), .ZN(n529) );
  OR2_X1 U450 ( .A1(A[38]), .A2(B[38]), .ZN(n530) );
  OR2_X1 U451 ( .A1(A[36]), .A2(B[36]), .ZN(n531) );
  NOR2_X1 U452 ( .A1(A[34]), .A2(B[34]), .ZN(n89) );
  INV_X1 U453 ( .A(n146), .ZN(n532) );
  CLKBUF_X1 U454 ( .A(n180), .Z(n556) );
  OAI21_X1 U455 ( .B1(n98), .B2(n104), .A(n99), .ZN(n533) );
  OR2_X1 U456 ( .A1(B[30]), .A2(A[30]), .ZN(n534) );
  NAND2_X1 U457 ( .A1(n543), .A2(n527), .ZN(n535) );
  CLKBUF_X1 U458 ( .A(n126), .Z(n536) );
  AOI21_X1 U459 ( .B1(n80), .B2(n533), .A(n81), .ZN(n537) );
  NOR2_X1 U460 ( .A1(n125), .A2(n540), .ZN(n538) );
  CLKBUF_X1 U461 ( .A(n182), .Z(n539) );
  NOR2_X1 U462 ( .A1(B[31]), .A2(A[31]), .ZN(n540) );
  CLKBUF_X1 U463 ( .A(B[31]), .Z(n541) );
  BUF_X1 U464 ( .A(n520), .Z(n548) );
  NOR2_X1 U465 ( .A1(n236), .A2(n198), .ZN(n542) );
  NOR2_X1 U466 ( .A1(n160), .A2(n169), .ZN(n543) );
  NOR2_X1 U467 ( .A1(B[25]), .A2(A[25]), .ZN(n544) );
  OR2_X1 U468 ( .A1(n541), .A2(A[31]), .ZN(n545) );
  BUF_X1 U469 ( .A(n220), .Z(n546) );
  CLKBUF_X1 U470 ( .A(n137), .Z(n547) );
  CLKBUF_X1 U471 ( .A(n181), .Z(n549) );
  NOR2_X1 U472 ( .A1(n110), .A2(n156), .ZN(n550) );
  CLKBUF_X1 U473 ( .A(B[21]), .Z(n551) );
  OR2_X1 U474 ( .A1(A[29]), .A2(n526), .ZN(n552) );
  CLKBUF_X1 U475 ( .A(n209), .Z(n553) );
  CLKBUF_X1 U476 ( .A(n546), .Z(n554) );
  NOR2_X1 U477 ( .A1(B[27]), .A2(A[27]), .ZN(n555) );
  CLKBUF_X1 U478 ( .A(n189), .Z(n557) );
  NOR2_X1 U479 ( .A1(B[30]), .A2(A[30]), .ZN(n125) );
  CLKBUF_X1 U480 ( .A(n147), .Z(n558) );
  XNOR2_X1 U481 ( .A(n91), .B(n559), .ZN(SUM[34]) );
  AND2_X1 U482 ( .A1(n88), .A2(n90), .ZN(n559) );
  BUF_X1 U483 ( .A(n157), .Z(n560) );
  CLKBUF_X1 U484 ( .A(n160), .Z(n561) );
  XNOR2_X1 U485 ( .A(n71), .B(n562), .ZN(SUM[36]) );
  AND2_X1 U486 ( .A1(n531), .A2(n70), .ZN(n562) );
  XNOR2_X1 U487 ( .A(n84), .B(n563), .ZN(SUM[35]) );
  AND2_X1 U488 ( .A1(n358), .A2(n83), .ZN(n563) );
  XNOR2_X1 U489 ( .A(n62), .B(n564), .ZN(SUM[37]) );
  AND2_X1 U490 ( .A1(n529), .A2(n61), .ZN(n564) );
  XNOR2_X1 U491 ( .A(n53), .B(n565), .ZN(SUM[38]) );
  AND2_X1 U492 ( .A1(n530), .A2(n52), .ZN(n565) );
  XNOR2_X1 U493 ( .A(n100), .B(n566), .ZN(SUM[33]) );
  AND2_X1 U494 ( .A1(n360), .A2(n99), .ZN(n566) );
  XNOR2_X1 U495 ( .A(n44), .B(n567), .ZN(SUM[39]) );
  AND2_X1 U496 ( .A1(n571), .A2(n43), .ZN(n567) );
  BUF_X1 U497 ( .A(n105), .Z(n568) );
  INV_X1 U498 ( .A(n534), .ZN(n123) );
  NOR2_X1 U499 ( .A1(A[4]), .A2(B[4]), .ZN(n337) );
  NOR2_X1 U500 ( .A1(A[12]), .A2(B[12]), .ZN(n290) );
  NOR2_X1 U501 ( .A1(A[10]), .A2(B[10]), .ZN(n306) );
  NOR2_X1 U502 ( .A1(A[16]), .A2(B[16]), .ZN(n261) );
  NOR2_X1 U503 ( .A1(A[18]), .A2(B[18]), .ZN(n247) );
  NOR2_X1 U504 ( .A1(A[14]), .A2(B[14]), .ZN(n276) );
  NOR2_X1 U505 ( .A1(A[6]), .A2(B[6]), .ZN(n327) );
  NOR2_X1 U506 ( .A1(A[7]), .A2(B[7]), .ZN(n324) );
  NOR2_X1 U507 ( .A1(A[11]), .A2(B[11]), .ZN(n301) );
  NOR2_X1 U508 ( .A1(A[17]), .A2(B[17]), .ZN(n256) );
  NOR2_X1 U509 ( .A1(A[9]), .A2(B[9]), .ZN(n313) );
  NOR2_X1 U510 ( .A1(A[5]), .A2(B[5]), .ZN(n332) );
  NOR2_X1 U511 ( .A1(A[15]), .A2(B[15]), .ZN(n271) );
  NOR2_X1 U512 ( .A1(A[3]), .A2(B[3]), .ZN(n343) );
  NOR2_X1 U513 ( .A1(A[8]), .A2(B[8]), .ZN(n316) );
  NOR2_X1 U514 ( .A1(A[2]), .A2(B[2]), .ZN(n346) );
  NOR2_X1 U515 ( .A1(A[1]), .A2(B[1]), .ZN(n350) );
  INV_X1 U516 ( .A(n236), .ZN(n230) );
  INV_X1 U517 ( .A(n195), .ZN(n193) );
  INV_X1 U518 ( .A(n215), .ZN(n213) );
  INV_X1 U519 ( .A(n214), .ZN(n212) );
  INV_X1 U520 ( .A(n556), .ZN(n174) );
  INV_X1 U521 ( .A(n535), .ZN(n154) );
  INV_X1 U522 ( .A(n154), .ZN(n152) );
  NAND2_X1 U523 ( .A1(n154), .A2(n525), .ZN(n130) );
  INV_X1 U524 ( .A(n94), .ZN(n92) );
  OAI21_X1 U525 ( .B1(n318), .B2(n297), .A(n298), .ZN(n292) );
  INV_X1 U526 ( .A(n264), .ZN(n263) );
  NOR2_X1 U527 ( .A1(n110), .A2(n535), .ZN(n108) );
  NOR2_X1 U528 ( .A1(n78), .A2(n56), .ZN(n54) );
  NAND2_X1 U529 ( .A1(n230), .A2(n216), .ZN(n214) );
  INV_X1 U530 ( .A(n78), .ZN(n76) );
  INV_X1 U531 ( .A(n297), .ZN(n295) );
  NAND2_X1 U532 ( .A1(n556), .A2(n167), .ZN(n165) );
  AOI21_X1 U533 ( .B1(n339), .B2(n330), .A(n331), .ZN(n329) );
  NOR2_X1 U534 ( .A1(n78), .A2(n65), .ZN(n63) );
  OAI21_X1 U535 ( .B1(n537), .B2(n65), .A(n70), .ZN(n64) );
  INV_X1 U536 ( .A(n531), .ZN(n65) );
  INV_X1 U537 ( .A(n48), .ZN(n46) );
  INV_X1 U538 ( .A(n197), .ZN(n195) );
  AOI21_X1 U539 ( .B1(n319), .B2(n265), .A(n266), .ZN(n264) );
  NOR2_X1 U540 ( .A1(n297), .A2(n267), .ZN(n265) );
  OAI21_X1 U541 ( .B1(n298), .B2(n267), .A(n268), .ZN(n266) );
  NAND2_X1 U542 ( .A1(n283), .A2(n269), .ZN(n267) );
  OAI21_X1 U543 ( .B1(n318), .B2(n279), .A(n280), .ZN(n278) );
  NAND2_X1 U544 ( .A1(n295), .A2(n283), .ZN(n279) );
  AOI21_X1 U545 ( .B1(n296), .B2(n283), .A(n284), .ZN(n280) );
  OAI21_X1 U546 ( .B1(n318), .B2(n309), .A(n310), .ZN(n308) );
  INV_X1 U547 ( .A(n312), .ZN(n310) );
  INV_X1 U548 ( .A(n311), .ZN(n309) );
  BUF_X1 U549 ( .A(n105), .Z(n1) );
  INV_X1 U550 ( .A(n319), .ZN(n318) );
  AOI21_X1 U551 ( .B1(n235), .B2(n216), .A(n522), .ZN(n215) );
  NAND2_X1 U552 ( .A1(n121), .A2(n154), .ZN(n119) );
  INV_X1 U553 ( .A(n547), .ZN(n135) );
  INV_X1 U554 ( .A(n525), .ZN(n134) );
  INV_X1 U555 ( .A(n237), .ZN(n235) );
  INV_X1 U556 ( .A(n533), .ZN(n95) );
  NOR2_X1 U557 ( .A1(n134), .A2(n123), .ZN(n121) );
  NAND2_X1 U558 ( .A1(n311), .A2(n299), .ZN(n297) );
  INV_X1 U559 ( .A(n340), .ZN(n339) );
  NAND2_X1 U560 ( .A1(n254), .A2(n238), .ZN(n236) );
  INV_X1 U561 ( .A(n255), .ZN(n253) );
  INV_X1 U562 ( .A(n254), .ZN(n252) );
  INV_X1 U563 ( .A(n217), .ZN(n216) );
  INV_X1 U564 ( .A(n298), .ZN(n296) );
  INV_X1 U565 ( .A(n549), .ZN(n179) );
  INV_X1 U566 ( .A(n349), .ZN(n348) );
  NAND2_X1 U567 ( .A1(n531), .A2(n529), .ZN(n56) );
  NOR2_X1 U568 ( .A1(n290), .A2(n285), .ZN(n283) );
  AOI21_X1 U569 ( .B1(n529), .B2(n68), .A(n59), .ZN(n57) );
  INV_X1 U570 ( .A(n61), .ZN(n59) );
  NOR2_X1 U571 ( .A1(n252), .A2(n247), .ZN(n243) );
  OAI21_X1 U572 ( .B1(n253), .B2(n247), .A(n248), .ZN(n244) );
  AOI21_X1 U573 ( .B1(n299), .B2(n312), .A(n300), .ZN(n298) );
  OAI21_X1 U574 ( .B1(n301), .B2(n307), .A(n302), .ZN(n300) );
  AOI21_X1 U575 ( .B1(n341), .B2(n349), .A(n342), .ZN(n340) );
  NOR2_X1 U576 ( .A1(n346), .A2(n343), .ZN(n341) );
  OAI21_X1 U577 ( .B1(n343), .B2(n347), .A(n344), .ZN(n342) );
  AOI21_X1 U578 ( .B1(n55), .B2(n530), .A(n50), .ZN(n48) );
  INV_X1 U579 ( .A(n52), .ZN(n50) );
  AOI21_X1 U580 ( .B1(n238), .B2(n255), .A(n239), .ZN(n237) );
  OAI21_X1 U581 ( .B1(n313), .B2(n317), .A(n314), .ZN(n312) );
  OAI21_X1 U582 ( .B1(n332), .B2(n338), .A(n333), .ZN(n331) );
  OAI21_X1 U583 ( .B1(n350), .B2(n353), .A(n351), .ZN(n349) );
  OAI21_X1 U584 ( .B1(n340), .B2(n320), .A(n321), .ZN(n319) );
  AOI21_X1 U585 ( .B1(n322), .B2(n331), .A(n323), .ZN(n321) );
  NAND2_X1 U586 ( .A1(n330), .A2(n322), .ZN(n320) );
  OAI21_X1 U587 ( .B1(n324), .B2(n328), .A(n325), .ZN(n323) );
  NOR2_X1 U588 ( .A1(n214), .A2(n553), .ZN(n205) );
  NOR2_X1 U589 ( .A1(n236), .A2(n225), .ZN(n223) );
  OAI21_X1 U590 ( .B1(n237), .B2(n225), .A(n228), .ZN(n224) );
  INV_X1 U591 ( .A(n226), .ZN(n225) );
  INV_X1 U592 ( .A(n104), .ZN(n102) );
  NOR2_X1 U593 ( .A1(n94), .A2(n87), .ZN(n85) );
  OAI21_X1 U594 ( .B1(n95), .B2(n87), .A(n90), .ZN(n86) );
  INV_X1 U595 ( .A(n88), .ZN(n87) );
  INV_X1 U596 ( .A(n262), .ZN(n260) );
  NOR2_X1 U597 ( .A1(n327), .A2(n324), .ZN(n322) );
  OAI21_X1 U598 ( .B1(n98), .B2(n104), .A(n99), .ZN(n97) );
  NOR2_X1 U599 ( .A1(n276), .A2(n271), .ZN(n269) );
  NOR2_X1 U600 ( .A1(n306), .A2(n301), .ZN(n299) );
  NOR2_X1 U601 ( .A1(n337), .A2(n332), .ZN(n330) );
  OAI21_X1 U602 ( .B1(n256), .B2(n262), .A(n257), .ZN(n255) );
  OAI21_X1 U603 ( .B1(n135), .B2(n123), .A(n536), .ZN(n122) );
  INV_X1 U604 ( .A(n148), .ZN(n146) );
  NOR2_X1 U605 ( .A1(n261), .A2(n256), .ZN(n254) );
  NOR2_X1 U606 ( .A1(n316), .A2(n313), .ZN(n311) );
  AOI21_X1 U607 ( .B1(n269), .B2(n284), .A(n270), .ZN(n268) );
  OAI21_X1 U608 ( .B1(n271), .B2(n277), .A(n272), .ZN(n270) );
  AOI21_X1 U609 ( .B1(n278), .B2(n379), .A(n275), .ZN(n273) );
  INV_X1 U610 ( .A(n277), .ZN(n275) );
  AOI21_X1 U611 ( .B1(n308), .B2(n383), .A(n305), .ZN(n303) );
  INV_X1 U612 ( .A(n307), .ZN(n305) );
  AOI21_X1 U613 ( .B1(n339), .B2(n389), .A(n336), .ZN(n334) );
  INV_X1 U614 ( .A(n338), .ZN(n336) );
  AOI21_X1 U615 ( .B1(n292), .B2(n381), .A(n289), .ZN(n287) );
  INV_X1 U616 ( .A(n291), .ZN(n289) );
  INV_X1 U617 ( .A(n169), .ZN(n167) );
  OAI21_X1 U618 ( .B1(n318), .B2(n316), .A(n317), .ZN(n315) );
  AOI21_X1 U619 ( .B1(n549), .B2(n167), .A(n168), .ZN(n166) );
  INV_X1 U620 ( .A(n170), .ZN(n168) );
  INV_X1 U621 ( .A(n103), .ZN(n361) );
  INV_X1 U622 ( .A(n70), .ZN(n68) );
  INV_X1 U623 ( .A(n240), .ZN(n374) );
  INV_X1 U624 ( .A(n247), .ZN(n246) );
  INV_X1 U625 ( .A(n89), .ZN(n88) );
  INV_X1 U626 ( .A(n227), .ZN(n226) );
  INV_X1 U627 ( .A(n561), .ZN(n366) );
  INV_X1 U628 ( .A(n539), .ZN(n368) );
  INV_X1 U629 ( .A(n327), .ZN(n387) );
  INV_X1 U630 ( .A(n316), .ZN(n385) );
  INV_X1 U631 ( .A(n346), .ZN(n391) );
  INV_X1 U632 ( .A(n256), .ZN(n376) );
  INV_X1 U633 ( .A(n271), .ZN(n378) );
  INV_X1 U634 ( .A(n261), .ZN(n377) );
  INV_X1 U635 ( .A(n301), .ZN(n382) );
  INV_X1 U636 ( .A(n332), .ZN(n388) );
  INV_X1 U637 ( .A(n313), .ZN(n384) );
  INV_X1 U638 ( .A(n276), .ZN(n379) );
  INV_X1 U639 ( .A(n337), .ZN(n389) );
  INV_X1 U640 ( .A(n306), .ZN(n383) );
  NAND2_X1 U641 ( .A1(n386), .A2(n325), .ZN(n34) );
  INV_X1 U642 ( .A(n324), .ZN(n386) );
  INV_X1 U643 ( .A(n290), .ZN(n381) );
  NAND2_X1 U644 ( .A1(n390), .A2(n344), .ZN(n38) );
  INV_X1 U645 ( .A(n343), .ZN(n390) );
  INV_X1 U646 ( .A(n98), .ZN(n360) );
  INV_X1 U647 ( .A(n350), .ZN(n392) );
  INV_X1 U648 ( .A(n202), .ZN(n370) );
  INV_X1 U649 ( .A(n82), .ZN(n358) );
  INV_X1 U650 ( .A(n554), .ZN(n372) );
  INV_X1 U651 ( .A(n285), .ZN(n380) );
  NOR2_X1 U652 ( .A1(B[26]), .A2(A[26]), .ZN(n169) );
  NOR2_X1 U653 ( .A1(B[20]), .A2(A[20]), .ZN(n227) );
  NOR2_X1 U654 ( .A1(B[21]), .A2(A[21]), .ZN(n220) );
  NOR2_X1 U655 ( .A1(B[31]), .A2(A[31]), .ZN(n114) );
  NOR2_X1 U656 ( .A1(B[25]), .A2(A[25]), .ZN(n182) );
  NOR2_X1 U657 ( .A1(B[27]), .A2(A[27]), .ZN(n160) );
  NAND2_X1 U658 ( .A1(A[32]), .A2(B[32]), .ZN(n104) );
  NAND2_X1 U659 ( .A1(A[34]), .A2(B[34]), .ZN(n90) );
  NAND2_X1 U660 ( .A1(n372), .A2(n221), .ZN(n20) );
  NAND2_X1 U661 ( .A1(n368), .A2(n183), .ZN(n16) );
  NOR2_X1 U662 ( .A1(A[13]), .A2(B[13]), .ZN(n285) );
  NAND2_X1 U663 ( .A1(A[37]), .A2(B[37]), .ZN(n61) );
  NAND2_X1 U664 ( .A1(n377), .A2(n262), .ZN(n25) );
  NAND2_X1 U665 ( .A1(A[6]), .A2(B[6]), .ZN(n328) );
  XOR2_X1 U666 ( .A(n329), .B(n35), .Z(SUM[6]) );
  NAND2_X1 U667 ( .A1(n387), .A2(n328), .ZN(n35) );
  XOR2_X1 U668 ( .A(n242), .B(n22), .Z(SUM[19]) );
  NAND2_X1 U669 ( .A1(n374), .A2(n241), .ZN(n22) );
  XOR2_X1 U670 ( .A(n171), .B(n15), .Z(SUM[26]) );
  NAND2_X1 U671 ( .A1(A[16]), .A2(B[16]), .ZN(n262) );
  NAND2_X1 U672 ( .A1(A[24]), .A2(B[24]), .ZN(n190) );
  NAND2_X1 U673 ( .A1(A[8]), .A2(B[8]), .ZN(n317) );
  NAND2_X1 U674 ( .A1(A[14]), .A2(B[14]), .ZN(n277) );
  NAND2_X1 U675 ( .A1(A[10]), .A2(B[10]), .ZN(n307) );
  NAND2_X1 U676 ( .A1(A[4]), .A2(B[4]), .ZN(n338) );
  NAND2_X1 U677 ( .A1(A[2]), .A2(B[2]), .ZN(n347) );
  XOR2_X1 U678 ( .A(n191), .B(n17), .Z(SUM[24]) );
  NAND2_X1 U679 ( .A1(n188), .A2(n190), .ZN(n17) );
  XOR2_X1 U680 ( .A(n211), .B(n19), .Z(SUM[22]) );
  NAND2_X1 U681 ( .A1(n208), .A2(n210), .ZN(n19) );
  XOR2_X1 U682 ( .A(n162), .B(n14), .Z(SUM[27]) );
  NAND2_X1 U683 ( .A1(n366), .A2(n161), .ZN(n14) );
  XOR2_X1 U684 ( .A(n140), .B(n12), .Z(SUM[29]) );
  NAND2_X1 U685 ( .A1(n552), .A2(n139), .ZN(n12) );
  NAND2_X1 U686 ( .A1(n545), .A2(n521), .ZN(n10) );
  NAND2_X1 U687 ( .A1(n370), .A2(n203), .ZN(n18) );
  NAND2_X1 U688 ( .A1(n145), .A2(n532), .ZN(n13) );
  NAND2_X1 U689 ( .A1(n534), .A2(n536), .ZN(n11) );
  NAND2_X1 U690 ( .A1(n361), .A2(n104), .ZN(n9) );
  XOR2_X1 U691 ( .A(n249), .B(n23), .Z(SUM[18]) );
  NAND2_X1 U692 ( .A1(n246), .A2(n248), .ZN(n23) );
  XOR2_X1 U693 ( .A(n229), .B(n21), .Z(SUM[20]) );
  NAND2_X1 U694 ( .A1(n226), .A2(n228), .ZN(n21) );
  NAND2_X1 U695 ( .A1(n376), .A2(n257), .ZN(n24) );
  XOR2_X1 U696 ( .A(n273), .B(n26), .Z(SUM[15]) );
  NAND2_X1 U697 ( .A1(n378), .A2(n272), .ZN(n26) );
  XNOR2_X1 U698 ( .A(n308), .B(n31), .ZN(SUM[10]) );
  NAND2_X1 U699 ( .A1(n383), .A2(n307), .ZN(n31) );
  XNOR2_X1 U700 ( .A(n315), .B(n32), .ZN(SUM[9]) );
  NAND2_X1 U701 ( .A1(n384), .A2(n314), .ZN(n32) );
  XOR2_X1 U702 ( .A(n40), .B(n353), .Z(SUM[1]) );
  NAND2_X1 U703 ( .A1(n392), .A2(n351), .ZN(n40) );
  XOR2_X1 U704 ( .A(n348), .B(n39), .Z(SUM[2]) );
  NAND2_X1 U705 ( .A1(n391), .A2(n347), .ZN(n39) );
  XNOR2_X1 U706 ( .A(n345), .B(n38), .ZN(SUM[3]) );
  OAI21_X1 U707 ( .B1(n348), .B2(n346), .A(n347), .ZN(n345) );
  XNOR2_X1 U708 ( .A(n339), .B(n37), .ZN(SUM[4]) );
  NAND2_X1 U709 ( .A1(n389), .A2(n338), .ZN(n37) );
  XOR2_X1 U710 ( .A(n334), .B(n36), .Z(SUM[5]) );
  NAND2_X1 U711 ( .A1(n388), .A2(n333), .ZN(n36) );
  XOR2_X1 U712 ( .A(n318), .B(n33), .Z(SUM[8]) );
  NAND2_X1 U713 ( .A1(n385), .A2(n317), .ZN(n33) );
  XNOR2_X1 U714 ( .A(n326), .B(n34), .ZN(SUM[7]) );
  OAI21_X1 U715 ( .B1(n329), .B2(n327), .A(n328), .ZN(n326) );
  AND2_X1 U716 ( .A1(n570), .A2(n353), .ZN(SUM[0]) );
  NAND2_X1 U717 ( .A1(A[7]), .A2(B[7]), .ZN(n325) );
  NAND2_X1 U718 ( .A1(A[0]), .A2(B[0]), .ZN(n353) );
  NAND2_X1 U719 ( .A1(A[18]), .A2(B[18]), .ZN(n248) );
  NAND2_X1 U720 ( .A1(A[12]), .A2(B[12]), .ZN(n291) );
  NAND2_X1 U721 ( .A1(A[15]), .A2(B[15]), .ZN(n272) );
  NAND2_X1 U722 ( .A1(A[17]), .A2(B[17]), .ZN(n257) );
  XNOR2_X1 U723 ( .A(n278), .B(n27), .ZN(SUM[14]) );
  NAND2_X1 U724 ( .A1(n379), .A2(n277), .ZN(n27) );
  XNOR2_X1 U725 ( .A(n292), .B(n29), .ZN(SUM[12]) );
  NAND2_X1 U726 ( .A1(n381), .A2(n291), .ZN(n29) );
  NAND2_X1 U727 ( .A1(A[23]), .A2(B[23]), .ZN(n203) );
  NAND2_X1 U728 ( .A1(A[11]), .A2(B[11]), .ZN(n302) );
  NAND2_X1 U729 ( .A1(A[9]), .A2(B[9]), .ZN(n314) );
  NAND2_X1 U730 ( .A1(A[1]), .A2(B[1]), .ZN(n351) );
  NAND2_X1 U731 ( .A1(A[5]), .A2(B[5]), .ZN(n333) );
  NAND2_X1 U732 ( .A1(A[3]), .A2(B[3]), .ZN(n344) );
  NAND2_X1 U733 ( .A1(A[38]), .A2(B[38]), .ZN(n52) );
  NAND2_X1 U734 ( .A1(A[13]), .A2(B[13]), .ZN(n286) );
  NAND2_X1 U735 ( .A1(B[22]), .A2(A[22]), .ZN(n210) );
  NAND2_X1 U736 ( .A1(A[39]), .A2(B[39]), .ZN(n43) );
  XOR2_X1 U737 ( .A(n287), .B(n28), .Z(SUM[13]) );
  NAND2_X1 U738 ( .A1(n380), .A2(n286), .ZN(n28) );
  XOR2_X1 U739 ( .A(n303), .B(n30), .Z(SUM[11]) );
  NAND2_X1 U740 ( .A1(n382), .A2(n302), .ZN(n30) );
  OR2_X1 U741 ( .A1(A[0]), .A2(B[0]), .ZN(n570) );
  OR2_X1 U742 ( .A1(A[39]), .A2(B[39]), .ZN(n571) );
  NAND2_X1 U743 ( .A1(A[35]), .A2(B[35]), .ZN(n83) );
  INV_X1 U744 ( .A(n560), .ZN(n155) );
  NAND2_X1 U745 ( .A1(A[21]), .A2(n551), .ZN(n221) );
  INV_X1 U746 ( .A(n558), .ZN(n145) );
  NAND2_X1 U747 ( .A1(n167), .A2(n170), .ZN(n15) );
  OAI21_X1 U748 ( .B1(n544), .B2(n190), .A(n183), .ZN(n181) );
  XOR2_X1 U749 ( .A(n222), .B(n20), .Z(SUM[21]) );
  NOR2_X1 U750 ( .A1(n247), .A2(n240), .ZN(n238) );
  OAI21_X1 U751 ( .B1(n240), .B2(n248), .A(n241), .ZN(n239) );
  NAND2_X1 U752 ( .A1(A[19]), .A2(B[19]), .ZN(n241) );
  NOR2_X1 U753 ( .A1(A[19]), .A2(B[19]), .ZN(n240) );
  INV_X1 U754 ( .A(n218), .ZN(n217) );
  NOR2_X1 U755 ( .A1(n227), .A2(n220), .ZN(n218) );
  INV_X1 U756 ( .A(n542), .ZN(n194) );
  NOR2_X1 U757 ( .A1(n236), .A2(n198), .ZN(n196) );
  INV_X1 U758 ( .A(n537), .ZN(n77) );
  NAND2_X1 U759 ( .A1(A[33]), .A2(B[33]), .ZN(n99) );
  AOI21_X1 U760 ( .B1(n197), .B2(n108), .A(n109), .ZN(n107) );
  NAND2_X1 U761 ( .A1(A[36]), .A2(B[36]), .ZN(n70) );
  XOR2_X1 U762 ( .A(n204), .B(n18), .Z(SUM[23]) );
  OAI21_X1 U763 ( .B1(n215), .B2(n553), .A(n210), .ZN(n206) );
  NOR2_X1 U764 ( .A1(n89), .A2(n82), .ZN(n80) );
  XNOR2_X1 U765 ( .A(n263), .B(n25), .ZN(SUM[16]) );
  XOR2_X1 U766 ( .A(n258), .B(n24), .Z(SUM[17]) );
  AOI21_X1 U767 ( .B1(n263), .B2(n185), .A(n186), .ZN(n184) );
  AOI21_X1 U768 ( .B1(n263), .B2(n377), .A(n260), .ZN(n258) );
  AOI21_X1 U769 ( .B1(n263), .B2(n254), .A(n255), .ZN(n249) );
  AOI21_X1 U770 ( .B1(n263), .B2(n230), .A(n235), .ZN(n229) );
  AOI21_X1 U771 ( .B1(n263), .B2(n212), .A(n213), .ZN(n211) );
  AOI21_X1 U772 ( .B1(n263), .B2(n542), .A(n193), .ZN(n191) );
  AOI21_X1 U773 ( .B1(n263), .B2(n243), .A(n244), .ZN(n242) );
  AOI21_X1 U774 ( .B1(n263), .B2(n205), .A(n206), .ZN(n204) );
  AOI21_X1 U775 ( .B1(n263), .B2(n223), .A(n224), .ZN(n222) );
  AOI21_X1 U776 ( .B1(n263), .B2(n163), .A(n164), .ZN(n162) );
  OAI21_X1 U777 ( .B1(n285), .B2(n291), .A(n286), .ZN(n284) );
  NOR2_X1 U778 ( .A1(A[32]), .A2(B[32]), .ZN(n103) );
  XOR2_X1 U779 ( .A(n116), .B(n10), .Z(SUM[31]) );
  AOI21_X1 U780 ( .B1(n155), .B2(n525), .A(n547), .ZN(n131) );
  AOI21_X1 U781 ( .B1(n121), .B2(n155), .A(n122), .ZN(n120) );
  AOI21_X1 U782 ( .B1(n155), .B2(n145), .A(n146), .ZN(n144) );
  NAND2_X1 U783 ( .A1(B[27]), .A2(A[27]), .ZN(n161) );
  AOI21_X1 U784 ( .B1(n263), .B2(n172), .A(n173), .ZN(n171) );
  AOI21_X1 U785 ( .B1(n263), .B2(n141), .A(n142), .ZN(n140) );
  OAI21_X1 U786 ( .B1(n264), .B2(n106), .A(n107), .ZN(n105) );
  INV_X1 U787 ( .A(n557), .ZN(n188) );
  NOR2_X1 U788 ( .A1(n182), .A2(n189), .ZN(n180) );
  OAI21_X1 U789 ( .B1(n237), .B2(n198), .A(n199), .ZN(n197) );
  NAND2_X1 U790 ( .A1(A[20]), .A2(B[20]), .ZN(n228) );
  AOI21_X1 U791 ( .B1(n80), .B2(n97), .A(n81), .ZN(n79) );
  XOR2_X1 U792 ( .A(n149), .B(n13), .Z(SUM[28]) );
  AOI21_X1 U793 ( .B1(n263), .B2(n150), .A(n151), .ZN(n149) );
  NAND2_X1 U794 ( .A1(B[25]), .A2(A[25]), .ZN(n183) );
  XOR2_X1 U795 ( .A(n127), .B(n11), .Z(SUM[30]) );
  AOI21_X1 U796 ( .B1(n263), .B2(n128), .A(n129), .ZN(n127) );
  NOR2_X1 U797 ( .A1(n209), .A2(n202), .ZN(n200) );
  NAND2_X1 U798 ( .A1(n218), .A2(n200), .ZN(n198) );
  AOI21_X1 U799 ( .B1(n219), .B2(n200), .A(n201), .ZN(n199) );
  INV_X1 U800 ( .A(n553), .ZN(n208) );
  NOR2_X1 U801 ( .A1(B[22]), .A2(A[22]), .ZN(n209) );
  NAND2_X1 U802 ( .A1(n154), .A2(n145), .ZN(n143) );
  INV_X1 U803 ( .A(n96), .ZN(n94) );
  NAND2_X1 U804 ( .A1(n96), .A2(n80), .ZN(n78) );
  AOI21_X1 U805 ( .B1(n263), .B2(n117), .A(n118), .ZN(n116) );
  NOR2_X1 U806 ( .A1(n147), .A2(n138), .ZN(n136) );
  NAND2_X1 U807 ( .A1(n550), .A2(n196), .ZN(n106) );
  NAND2_X1 U808 ( .A1(B[31]), .A2(A[31]), .ZN(n115) );
  XOR2_X1 U809 ( .A(n184), .B(n16), .Z(SUM[25]) );
  NOR2_X1 U810 ( .A1(n194), .A2(n557), .ZN(n185) );
  NOR2_X1 U811 ( .A1(n194), .A2(n174), .ZN(n172) );
  NOR2_X1 U812 ( .A1(n194), .A2(n165), .ZN(n163) );
  NOR2_X1 U813 ( .A1(n194), .A2(n152), .ZN(n150) );
  NOR2_X1 U814 ( .A1(n194), .A2(n143), .ZN(n141) );
  NOR2_X1 U815 ( .A1(n194), .A2(n130), .ZN(n128) );
  NOR2_X1 U816 ( .A1(n194), .A2(n119), .ZN(n117) );
  OAI21_X1 U817 ( .B1(n546), .B2(n228), .A(n221), .ZN(n219) );
  OAI21_X1 U818 ( .B1(n82), .B2(n90), .A(n83), .ZN(n81) );
  OAI21_X1 U819 ( .B1(n195), .B2(n557), .A(n190), .ZN(n186) );
  OAI21_X1 U820 ( .B1(n195), .B2(n174), .A(n179), .ZN(n173) );
  OAI21_X1 U821 ( .B1(n195), .B2(n165), .A(n166), .ZN(n164) );
  OAI21_X1 U822 ( .B1(n195), .B2(n152), .A(n560), .ZN(n151) );
  OAI21_X1 U823 ( .B1(n195), .B2(n143), .A(n144), .ZN(n142) );
  OAI21_X1 U824 ( .B1(n195), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U825 ( .B1(n119), .B2(n195), .A(n120), .ZN(n118) );
  OAI21_X1 U826 ( .B1(n202), .B2(n210), .A(n203), .ZN(n201) );
  NOR2_X1 U827 ( .A1(B[24]), .A2(A[24]), .ZN(n189) );
  OAI21_X1 U828 ( .B1(n79), .B2(n56), .A(n57), .ZN(n55) );
  NOR2_X1 U829 ( .A1(n103), .A2(n98), .ZN(n96) );
  AOI21_X1 U830 ( .B1(n158), .B2(n181), .A(n159), .ZN(n157) );
  NAND2_X1 U831 ( .A1(n543), .A2(n180), .ZN(n156) );
  NOR2_X1 U832 ( .A1(n160), .A2(n169), .ZN(n158) );
  NAND2_X1 U833 ( .A1(B[26]), .A2(A[26]), .ZN(n170) );
  NAND2_X1 U834 ( .A1(B[28]), .A2(A[28]), .ZN(n148) );
  NOR2_X1 U835 ( .A1(B[28]), .A2(A[28]), .ZN(n147) );
  NAND2_X1 U836 ( .A1(B[29]), .A2(A[29]), .ZN(n139) );
  NOR2_X1 U837 ( .A1(B[29]), .A2(A[29]), .ZN(n138) );
  OAI21_X1 U838 ( .B1(n157), .B2(n110), .A(n111), .ZN(n109) );
  OAI21_X1 U839 ( .B1(n555), .B2(n170), .A(n161), .ZN(n159) );
  AOI21_X1 U840 ( .B1(n137), .B2(n112), .A(n113), .ZN(n111) );
  NAND2_X1 U841 ( .A1(n136), .A2(n538), .ZN(n110) );
  NOR2_X1 U842 ( .A1(n540), .A2(n125), .ZN(n112) );
  NAND2_X1 U843 ( .A1(B[30]), .A2(A[30]), .ZN(n126) );
  XNOR2_X1 U844 ( .A(n548), .B(n9), .ZN(SUM[32]) );
  AOI21_X1 U845 ( .B1(n1), .B2(n54), .A(n523), .ZN(n53) );
  AOI21_X1 U846 ( .B1(n520), .B2(n63), .A(n64), .ZN(n62) );
  AOI21_X1 U847 ( .B1(n1), .B2(n76), .A(n77), .ZN(n71) );
  AOI21_X1 U848 ( .B1(n1), .B2(n92), .A(n533), .ZN(n91) );
  AOI21_X1 U849 ( .B1(n568), .B2(n361), .A(n102), .ZN(n100) );
  AOI21_X1 U850 ( .B1(n520), .B2(n524), .A(n46), .ZN(n44) );
  AOI21_X1 U851 ( .B1(n568), .B2(n85), .A(n86), .ZN(n84) );
  OAI21_X1 U852 ( .B1(n528), .B2(n148), .A(n139), .ZN(n137) );
  OAI21_X1 U853 ( .B1(n114), .B2(n126), .A(n115), .ZN(n113) );
endmodule


module datapath_DW01_add_9 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n9, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n43, n44, n46, n48, n50, n52, n53, n54, n55, n56, n57, n59, n61,
         n62, n63, n64, n65, n68, n70, n71, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n93, n94, n95, n96,
         n97, n98, n99, n100, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n195, n196, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n226, n227, n228, n229, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n246,
         n247, n248, n249, n252, n253, n254, n255, n256, n257, n258, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n275, n276, n277, n278, n279, n280, n283, n284, n285,
         n286, n287, n289, n290, n291, n292, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n353, n358, n360, n361, n362,
         n364, n370, n372, n374, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569;

  NOR2_X1 U437 ( .A1(n189), .A2(n182), .ZN(n520) );
  BUF_X1 U438 ( .A(n105), .Z(n521) );
  CLKBUF_X1 U439 ( .A(n157), .Z(n541) );
  XNOR2_X1 U440 ( .A(n149), .B(n522), .ZN(SUM[28]) );
  AND2_X1 U441 ( .A1(n145), .A2(n148), .ZN(n522) );
  NOR2_X1 U442 ( .A1(n156), .A2(n110), .ZN(n523) );
  XNOR2_X1 U443 ( .A(n140), .B(n524), .ZN(SUM[29]) );
  AND2_X1 U444 ( .A1(n364), .A2(n139), .ZN(n524) );
  BUF_X1 U445 ( .A(n552), .Z(n567) );
  CLKBUF_X1 U446 ( .A(n181), .Z(n525) );
  OR2_X1 U447 ( .A1(A[37]), .A2(B[37]), .ZN(n526) );
  OR2_X1 U448 ( .A1(A[36]), .A2(B[36]), .ZN(n527) );
  OR2_X1 U449 ( .A1(A[38]), .A2(B[38]), .ZN(n528) );
  AND2_X1 U450 ( .A1(n532), .A2(n353), .ZN(SUM[0]) );
  OR2_X1 U451 ( .A1(n537), .A2(n567), .ZN(n530) );
  AND2_X1 U452 ( .A1(n54), .A2(n528), .ZN(n531) );
  OR2_X1 U453 ( .A1(A[0]), .A2(B[0]), .ZN(n532) );
  CLKBUF_X1 U454 ( .A(n161), .Z(n533) );
  NOR2_X1 U455 ( .A1(A[30]), .A2(B[30]), .ZN(n534) );
  CLKBUF_X1 U456 ( .A(n137), .Z(n535) );
  XNOR2_X1 U457 ( .A(n127), .B(n536), .ZN(SUM[30]) );
  AND2_X1 U458 ( .A1(n124), .A2(n538), .ZN(n536) );
  CLKBUF_X1 U459 ( .A(n147), .Z(n537) );
  CLKBUF_X1 U460 ( .A(n126), .Z(n538) );
  OAI21_X1 U461 ( .B1(n237), .B2(n198), .A(n199), .ZN(n539) );
  CLKBUF_X1 U462 ( .A(n558), .Z(n540) );
  OR2_X2 U463 ( .A1(n236), .A2(n198), .ZN(n542) );
  CLKBUF_X1 U464 ( .A(n227), .Z(n543) );
  XNOR2_X1 U465 ( .A(n116), .B(n544), .ZN(SUM[31]) );
  AND2_X1 U466 ( .A1(n362), .A2(n115), .ZN(n544) );
  NOR2_X1 U467 ( .A1(n160), .A2(n169), .ZN(n545) );
  NOR2_X1 U468 ( .A1(B[25]), .A2(A[25]), .ZN(n546) );
  CLKBUF_X1 U469 ( .A(B[25]), .Z(n547) );
  NOR2_X1 U470 ( .A1(B[27]), .A2(A[27]), .ZN(n548) );
  CLKBUF_X1 U471 ( .A(n169), .Z(n549) );
  CLKBUF_X1 U472 ( .A(n534), .Z(n550) );
  CLKBUF_X1 U473 ( .A(B[27]), .Z(n551) );
  NOR2_X1 U474 ( .A1(B[29]), .A2(A[29]), .ZN(n552) );
  NOR2_X1 U475 ( .A1(n114), .A2(n534), .ZN(n553) );
  CLKBUF_X1 U476 ( .A(n209), .Z(n554) );
  CLKBUF_X1 U477 ( .A(n220), .Z(n555) );
  OR2_X1 U478 ( .A1(A[25]), .A2(n547), .ZN(n556) );
  OR2_X1 U479 ( .A1(A[27]), .A2(n551), .ZN(n557) );
  NOR2_X1 U480 ( .A1(B[31]), .A2(A[31]), .ZN(n558) );
  XNOR2_X1 U481 ( .A(n71), .B(n559), .ZN(SUM[36]) );
  AND2_X1 U482 ( .A1(n527), .A2(n70), .ZN(n559) );
  XNOR2_X1 U483 ( .A(n100), .B(n560), .ZN(SUM[33]) );
  AND2_X1 U484 ( .A1(n360), .A2(n99), .ZN(n560) );
  XNOR2_X1 U485 ( .A(n53), .B(n561), .ZN(SUM[38]) );
  AND2_X1 U486 ( .A1(n528), .A2(n52), .ZN(n561) );
  XNOR2_X1 U487 ( .A(n62), .B(n562), .ZN(SUM[37]) );
  AND2_X1 U488 ( .A1(n526), .A2(n61), .ZN(n562) );
  XNOR2_X1 U489 ( .A(n91), .B(n563), .ZN(SUM[34]) );
  AND2_X1 U490 ( .A1(n88), .A2(n90), .ZN(n563) );
  XNOR2_X1 U491 ( .A(n84), .B(n564), .ZN(SUM[35]) );
  AND2_X1 U492 ( .A1(n358), .A2(n83), .ZN(n564) );
  XNOR2_X1 U493 ( .A(n44), .B(n565), .ZN(SUM[39]) );
  AND2_X1 U494 ( .A1(n569), .A2(n43), .ZN(n565) );
  CLKBUF_X1 U495 ( .A(n156), .Z(n566) );
  BUF_X1 U496 ( .A(n105), .Z(n568) );
  NOR2_X1 U497 ( .A1(A[4]), .A2(B[4]), .ZN(n337) );
  NOR2_X1 U498 ( .A1(A[18]), .A2(B[18]), .ZN(n247) );
  NOR2_X1 U499 ( .A1(A[12]), .A2(B[12]), .ZN(n290) );
  NOR2_X1 U500 ( .A1(A[10]), .A2(B[10]), .ZN(n306) );
  NOR2_X1 U501 ( .A1(A[16]), .A2(B[16]), .ZN(n261) );
  NOR2_X1 U502 ( .A1(A[14]), .A2(B[14]), .ZN(n276) );
  NOR2_X1 U503 ( .A1(A[6]), .A2(B[6]), .ZN(n327) );
  NOR2_X1 U504 ( .A1(A[7]), .A2(B[7]), .ZN(n324) );
  NOR2_X1 U505 ( .A1(A[17]), .A2(B[17]), .ZN(n256) );
  NOR2_X1 U506 ( .A1(A[11]), .A2(B[11]), .ZN(n301) );
  NOR2_X1 U507 ( .A1(A[13]), .A2(B[13]), .ZN(n285) );
  NOR2_X1 U508 ( .A1(A[9]), .A2(B[9]), .ZN(n313) );
  NOR2_X1 U509 ( .A1(A[5]), .A2(B[5]), .ZN(n332) );
  NOR2_X1 U510 ( .A1(A[3]), .A2(B[3]), .ZN(n343) );
  NOR2_X1 U511 ( .A1(A[8]), .A2(B[8]), .ZN(n316) );
  NOR2_X1 U512 ( .A1(A[2]), .A2(B[2]), .ZN(n346) );
  NOR2_X1 U513 ( .A1(A[1]), .A2(B[1]), .ZN(n350) );
  INV_X1 U514 ( .A(n542), .ZN(n192) );
  INV_X1 U515 ( .A(n195), .ZN(n193) );
  INV_X1 U516 ( .A(n566), .ZN(n154) );
  NOR2_X1 U517 ( .A1(n78), .A2(n56), .ZN(n54) );
  NAND2_X1 U518 ( .A1(n154), .A2(n132), .ZN(n130) );
  INV_X1 U519 ( .A(n95), .ZN(n93) );
  INV_X1 U520 ( .A(n215), .ZN(n213) );
  INV_X1 U521 ( .A(n214), .ZN(n212) );
  OAI21_X1 U522 ( .B1(n318), .B2(n297), .A(n298), .ZN(n292) );
  INV_X1 U523 ( .A(n264), .ZN(n263) );
  AOI21_X1 U524 ( .B1(n155), .B2(n132), .A(n535), .ZN(n131) );
  NAND2_X1 U525 ( .A1(n234), .A2(n216), .ZN(n214) );
  NOR2_X1 U526 ( .A1(n236), .A2(n198), .ZN(n196) );
  INV_X1 U527 ( .A(n530), .ZN(n132) );
  INV_X1 U528 ( .A(n78), .ZN(n76) );
  INV_X1 U529 ( .A(n236), .ZN(n234) );
  INV_X1 U530 ( .A(n297), .ZN(n295) );
  INV_X1 U531 ( .A(n154), .ZN(n152) );
  INV_X1 U532 ( .A(n155), .ZN(n153) );
  NAND2_X1 U533 ( .A1(n154), .A2(n145), .ZN(n143) );
  INV_X1 U534 ( .A(n541), .ZN(n155) );
  AOI21_X1 U535 ( .B1(n339), .B2(n330), .A(n331), .ZN(n329) );
  AOI21_X1 U536 ( .B1(n235), .B2(n216), .A(n219), .ZN(n215) );
  INV_X1 U537 ( .A(n48), .ZN(n46) );
  NOR2_X1 U538 ( .A1(n78), .A2(n65), .ZN(n63) );
  OAI21_X1 U539 ( .B1(n75), .B2(n65), .A(n70), .ZN(n64) );
  INV_X1 U540 ( .A(n527), .ZN(n65) );
  AOI21_X1 U541 ( .B1(n319), .B2(n265), .A(n266), .ZN(n264) );
  NOR2_X1 U542 ( .A1(n297), .A2(n267), .ZN(n265) );
  OAI21_X1 U543 ( .B1(n298), .B2(n267), .A(n268), .ZN(n266) );
  NAND2_X1 U544 ( .A1(n283), .A2(n269), .ZN(n267) );
  OAI21_X1 U545 ( .B1(n318), .B2(n279), .A(n280), .ZN(n278) );
  AOI21_X1 U546 ( .B1(n296), .B2(n283), .A(n284), .ZN(n280) );
  NAND2_X1 U547 ( .A1(n295), .A2(n283), .ZN(n279) );
  OAI21_X1 U548 ( .B1(n318), .B2(n309), .A(n310), .ZN(n308) );
  INV_X1 U549 ( .A(n312), .ZN(n310) );
  INV_X1 U550 ( .A(n311), .ZN(n309) );
  INV_X1 U551 ( .A(n319), .ZN(n318) );
  NAND2_X1 U552 ( .A1(n121), .A2(n154), .ZN(n119) );
  NAND2_X1 U553 ( .A1(n520), .A2(n167), .ZN(n165) );
  INV_X1 U554 ( .A(n96), .ZN(n94) );
  INV_X1 U555 ( .A(n97), .ZN(n95) );
  BUF_X1 U556 ( .A(n105), .Z(n1) );
  NOR2_X1 U557 ( .A1(n530), .A2(n550), .ZN(n121) );
  INV_X1 U558 ( .A(n535), .ZN(n135) );
  NAND2_X1 U559 ( .A1(n254), .A2(n238), .ZN(n236) );
  NAND2_X1 U560 ( .A1(n311), .A2(n299), .ZN(n297) );
  INV_X1 U561 ( .A(n340), .ZN(n339) );
  INV_X1 U562 ( .A(n255), .ZN(n253) );
  INV_X1 U563 ( .A(n254), .ZN(n252) );
  INV_X1 U564 ( .A(n298), .ZN(n296) );
  INV_X1 U565 ( .A(n525), .ZN(n179) );
  INV_X1 U566 ( .A(n349), .ZN(n348) );
  INV_X1 U567 ( .A(n77), .ZN(n75) );
  INV_X1 U568 ( .A(n79), .ZN(n77) );
  INV_X1 U569 ( .A(n520), .ZN(n178) );
  INV_X1 U570 ( .A(n237), .ZN(n235) );
  NAND2_X1 U571 ( .A1(n527), .A2(n526), .ZN(n56) );
  INV_X1 U572 ( .A(n217), .ZN(n216) );
  INV_X1 U573 ( .A(n218), .ZN(n217) );
  INV_X1 U574 ( .A(n52), .ZN(n50) );
  NOR2_X1 U575 ( .A1(n276), .A2(n271), .ZN(n269) );
  NOR2_X1 U576 ( .A1(n247), .A2(n240), .ZN(n238) );
  NOR2_X1 U577 ( .A1(n236), .A2(n543), .ZN(n223) );
  OAI21_X1 U578 ( .B1(n237), .B2(n543), .A(n228), .ZN(n224) );
  INV_X1 U579 ( .A(n262), .ZN(n260) );
  NOR2_X1 U580 ( .A1(n252), .A2(n247), .ZN(n243) );
  OAI21_X1 U581 ( .B1(n253), .B2(n247), .A(n248), .ZN(n244) );
  AOI21_X1 U582 ( .B1(n299), .B2(n312), .A(n300), .ZN(n298) );
  OAI21_X1 U583 ( .B1(n301), .B2(n307), .A(n302), .ZN(n300) );
  AOI21_X1 U584 ( .B1(n341), .B2(n349), .A(n342), .ZN(n340) );
  NOR2_X1 U585 ( .A1(n346), .A2(n343), .ZN(n341) );
  OAI21_X1 U586 ( .B1(n343), .B2(n347), .A(n344), .ZN(n342) );
  AOI21_X1 U587 ( .B1(n526), .B2(n68), .A(n59), .ZN(n57) );
  INV_X1 U588 ( .A(n61), .ZN(n59) );
  OAI21_X1 U589 ( .B1(n98), .B2(n104), .A(n99), .ZN(n97) );
  NOR2_X1 U590 ( .A1(n147), .A2(n138), .ZN(n136) );
  AOI21_X1 U591 ( .B1(n80), .B2(n97), .A(n81), .ZN(n79) );
  OAI21_X1 U592 ( .B1(n256), .B2(n262), .A(n257), .ZN(n255) );
  OAI21_X1 U593 ( .B1(n313), .B2(n317), .A(n314), .ZN(n312) );
  OAI21_X1 U594 ( .B1(n332), .B2(n338), .A(n333), .ZN(n331) );
  OAI21_X1 U595 ( .B1(n285), .B2(n291), .A(n286), .ZN(n284) );
  OAI21_X1 U596 ( .B1(n350), .B2(n353), .A(n351), .ZN(n349) );
  OAI21_X1 U597 ( .B1(n340), .B2(n320), .A(n321), .ZN(n319) );
  AOI21_X1 U598 ( .B1(n322), .B2(n331), .A(n323), .ZN(n321) );
  NAND2_X1 U599 ( .A1(n330), .A2(n322), .ZN(n320) );
  OAI21_X1 U600 ( .B1(n324), .B2(n328), .A(n325), .ZN(n323) );
  INV_X1 U601 ( .A(n104), .ZN(n102) );
  NOR2_X1 U602 ( .A1(n94), .A2(n87), .ZN(n85) );
  OAI21_X1 U603 ( .B1(n95), .B2(n87), .A(n90), .ZN(n86) );
  INV_X1 U604 ( .A(n88), .ZN(n87) );
  NOR2_X1 U605 ( .A1(n214), .A2(n554), .ZN(n205) );
  NOR2_X1 U606 ( .A1(n327), .A2(n324), .ZN(n322) );
  AOI21_X1 U607 ( .B1(n238), .B2(n255), .A(n239), .ZN(n237) );
  NOR2_X1 U608 ( .A1(n306), .A2(n301), .ZN(n299) );
  NOR2_X1 U609 ( .A1(n337), .A2(n332), .ZN(n330) );
  OAI21_X1 U610 ( .B1(n135), .B2(n550), .A(n538), .ZN(n122) );
  NOR2_X1 U611 ( .A1(n261), .A2(n256), .ZN(n254) );
  NOR2_X1 U612 ( .A1(n316), .A2(n313), .ZN(n311) );
  NOR2_X1 U613 ( .A1(n290), .A2(n285), .ZN(n283) );
  AOI21_X1 U614 ( .B1(n269), .B2(n284), .A(n270), .ZN(n268) );
  NOR2_X1 U615 ( .A1(n189), .A2(n182), .ZN(n180) );
  INV_X1 U616 ( .A(n188), .ZN(n187) );
  AOI21_X1 U617 ( .B1(n292), .B2(n381), .A(n289), .ZN(n287) );
  INV_X1 U618 ( .A(n291), .ZN(n289) );
  AOI21_X1 U619 ( .B1(n308), .B2(n383), .A(n305), .ZN(n303) );
  INV_X1 U620 ( .A(n307), .ZN(n305) );
  AOI21_X1 U621 ( .B1(n339), .B2(n389), .A(n336), .ZN(n334) );
  INV_X1 U622 ( .A(n338), .ZN(n336) );
  AOI21_X1 U623 ( .B1(n278), .B2(n379), .A(n275), .ZN(n273) );
  INV_X1 U624 ( .A(n277), .ZN(n275) );
  INV_X1 U625 ( .A(n549), .ZN(n167) );
  INV_X1 U626 ( .A(n189), .ZN(n188) );
  AOI21_X1 U627 ( .B1(n155), .B2(n145), .A(n146), .ZN(n144) );
  INV_X1 U628 ( .A(n148), .ZN(n146) );
  OAI21_X1 U629 ( .B1(n329), .B2(n327), .A(n328), .ZN(n326) );
  OAI21_X1 U630 ( .B1(n318), .B2(n316), .A(n317), .ZN(n315) );
  OAI21_X1 U631 ( .B1(n348), .B2(n346), .A(n347), .ZN(n345) );
  AOI21_X1 U632 ( .B1(n525), .B2(n167), .A(n168), .ZN(n166) );
  INV_X1 U633 ( .A(n103), .ZN(n361) );
  INV_X1 U634 ( .A(n70), .ZN(n68) );
  INV_X1 U635 ( .A(n540), .ZN(n362) );
  INV_X1 U636 ( .A(n247), .ZN(n246) );
  INV_X1 U637 ( .A(n89), .ZN(n88) );
  INV_X1 U638 ( .A(n256), .ZN(n376) );
  NAND2_X1 U639 ( .A1(n387), .A2(n328), .ZN(n35) );
  INV_X1 U640 ( .A(n327), .ZN(n387) );
  NAND2_X1 U641 ( .A1(n386), .A2(n325), .ZN(n34) );
  INV_X1 U642 ( .A(n324), .ZN(n386) );
  NAND2_X1 U643 ( .A1(n389), .A2(n338), .ZN(n37) );
  INV_X1 U644 ( .A(n337), .ZN(n389) );
  NAND2_X1 U645 ( .A1(n381), .A2(n291), .ZN(n29) );
  INV_X1 U646 ( .A(n290), .ZN(n381) );
  NAND2_X1 U647 ( .A1(n383), .A2(n307), .ZN(n31) );
  INV_X1 U648 ( .A(n306), .ZN(n383) );
  NAND2_X1 U649 ( .A1(n385), .A2(n317), .ZN(n33) );
  INV_X1 U650 ( .A(n316), .ZN(n385) );
  NAND2_X1 U651 ( .A1(n391), .A2(n347), .ZN(n39) );
  INV_X1 U652 ( .A(n346), .ZN(n391) );
  NAND2_X1 U653 ( .A1(n379), .A2(n277), .ZN(n27) );
  INV_X1 U654 ( .A(n276), .ZN(n379) );
  INV_X1 U655 ( .A(n567), .ZN(n364) );
  NAND2_X1 U656 ( .A1(n390), .A2(n344), .ZN(n38) );
  INV_X1 U657 ( .A(n343), .ZN(n390) );
  NAND2_X1 U658 ( .A1(n384), .A2(n314), .ZN(n32) );
  INV_X1 U659 ( .A(n313), .ZN(n384) );
  INV_X1 U660 ( .A(n98), .ZN(n360) );
  NAND2_X1 U661 ( .A1(n382), .A2(n302), .ZN(n30) );
  INV_X1 U662 ( .A(n301), .ZN(n382) );
  NAND2_X1 U663 ( .A1(n388), .A2(n333), .ZN(n36) );
  INV_X1 U664 ( .A(n332), .ZN(n388) );
  NAND2_X1 U665 ( .A1(n380), .A2(n286), .ZN(n28) );
  INV_X1 U666 ( .A(n285), .ZN(n380) );
  NAND2_X1 U667 ( .A1(n392), .A2(n351), .ZN(n40) );
  INV_X1 U668 ( .A(n350), .ZN(n392) );
  NAND2_X1 U669 ( .A1(n378), .A2(n272), .ZN(n26) );
  INV_X1 U670 ( .A(n271), .ZN(n378) );
  NAND2_X1 U671 ( .A1(n377), .A2(n262), .ZN(n25) );
  INV_X1 U672 ( .A(n261), .ZN(n377) );
  INV_X1 U673 ( .A(n82), .ZN(n358) );
  INV_X1 U674 ( .A(n555), .ZN(n372) );
  INV_X1 U675 ( .A(n202), .ZN(n370) );
  INV_X1 U676 ( .A(n240), .ZN(n374) );
  NOR2_X1 U677 ( .A1(B[25]), .A2(A[25]), .ZN(n182) );
  NOR2_X1 U678 ( .A1(B[29]), .A2(A[29]), .ZN(n138) );
  NOR2_X1 U679 ( .A1(A[26]), .A2(B[26]), .ZN(n169) );
  NOR2_X1 U680 ( .A1(A[34]), .A2(B[34]), .ZN(n89) );
  NOR2_X1 U681 ( .A1(A[33]), .A2(B[33]), .ZN(n98) );
  NOR2_X1 U682 ( .A1(A[21]), .A2(B[21]), .ZN(n220) );
  NOR2_X1 U683 ( .A1(B[23]), .A2(A[23]), .ZN(n202) );
  NOR2_X1 U684 ( .A1(A[35]), .A2(B[35]), .ZN(n82) );
  NAND2_X1 U685 ( .A1(B[28]), .A2(A[28]), .ZN(n148) );
  NOR2_X1 U686 ( .A1(A[19]), .A2(B[19]), .ZN(n240) );
  NOR2_X1 U687 ( .A1(A[15]), .A2(B[15]), .ZN(n271) );
  NAND2_X1 U688 ( .A1(A[37]), .A2(B[37]), .ZN(n61) );
  NAND2_X1 U689 ( .A1(A[6]), .A2(B[6]), .ZN(n328) );
  XOR2_X1 U690 ( .A(n222), .B(n20), .Z(SUM[21]) );
  NAND2_X1 U691 ( .A1(n372), .A2(n221), .ZN(n20) );
  XOR2_X1 U692 ( .A(n162), .B(n14), .Z(SUM[27]) );
  NAND2_X1 U693 ( .A1(n557), .A2(n533), .ZN(n14) );
  XOR2_X1 U694 ( .A(n229), .B(n21), .Z(SUM[20]) );
  NAND2_X1 U695 ( .A1(n226), .A2(n228), .ZN(n21) );
  XOR2_X1 U696 ( .A(n171), .B(n15), .Z(SUM[26]) );
  NAND2_X1 U697 ( .A1(B[22]), .A2(A[22]), .ZN(n210) );
  NAND2_X1 U698 ( .A1(A[8]), .A2(B[8]), .ZN(n317) );
  NAND2_X1 U699 ( .A1(A[4]), .A2(B[4]), .ZN(n338) );
  NAND2_X1 U700 ( .A1(A[7]), .A2(B[7]), .ZN(n325) );
  NAND2_X1 U701 ( .A1(A[12]), .A2(B[12]), .ZN(n291) );
  NAND2_X1 U702 ( .A1(A[16]), .A2(B[16]), .ZN(n262) );
  NAND2_X1 U703 ( .A1(A[10]), .A2(B[10]), .ZN(n307) );
  NAND2_X1 U704 ( .A1(A[2]), .A2(B[2]), .ZN(n347) );
  NAND2_X1 U705 ( .A1(A[0]), .A2(B[0]), .ZN(n353) );
  NAND2_X1 U706 ( .A1(A[18]), .A2(B[18]), .ZN(n248) );
  NAND2_X1 U707 ( .A1(A[38]), .A2(B[38]), .ZN(n52) );
  NAND2_X1 U708 ( .A1(A[17]), .A2(B[17]), .ZN(n257) );
  NAND2_X1 U709 ( .A1(A[14]), .A2(B[14]), .ZN(n277) );
  NAND2_X1 U710 ( .A1(B[20]), .A2(A[20]), .ZN(n228) );
  NAND2_X1 U711 ( .A1(A[11]), .A2(B[11]), .ZN(n302) );
  NAND2_X1 U712 ( .A1(A[13]), .A2(B[13]), .ZN(n286) );
  NAND2_X1 U713 ( .A1(A[9]), .A2(B[9]), .ZN(n314) );
  NAND2_X1 U714 ( .A1(A[1]), .A2(B[1]), .ZN(n351) );
  NAND2_X1 U715 ( .A1(A[3]), .A2(B[3]), .ZN(n344) );
  NAND2_X1 U716 ( .A1(A[5]), .A2(B[5]), .ZN(n333) );
  NAND2_X1 U717 ( .A1(A[19]), .A2(B[19]), .ZN(n241) );
  NAND2_X1 U718 ( .A1(A[39]), .A2(B[39]), .ZN(n43) );
  NAND2_X1 U719 ( .A1(A[15]), .A2(B[15]), .ZN(n272) );
  XOR2_X1 U720 ( .A(n191), .B(n17), .Z(SUM[24]) );
  NAND2_X1 U721 ( .A1(n188), .A2(n190), .ZN(n17) );
  XOR2_X1 U722 ( .A(n184), .B(n16), .Z(SUM[25]) );
  NAND2_X1 U723 ( .A1(n556), .A2(n183), .ZN(n16) );
  NAND2_X1 U724 ( .A1(n361), .A2(n104), .ZN(n9) );
  NAND2_X1 U725 ( .A1(n208), .A2(n210), .ZN(n19) );
  NAND2_X1 U726 ( .A1(n370), .A2(n203), .ZN(n18) );
  XNOR2_X1 U727 ( .A(n278), .B(n27), .ZN(SUM[14]) );
  XOR2_X1 U728 ( .A(n40), .B(n353), .Z(SUM[1]) );
  XOR2_X1 U729 ( .A(n348), .B(n39), .Z(SUM[2]) );
  XNOR2_X1 U730 ( .A(n345), .B(n38), .ZN(SUM[3]) );
  XNOR2_X1 U731 ( .A(n339), .B(n37), .ZN(SUM[4]) );
  XOR2_X1 U732 ( .A(n334), .B(n36), .Z(SUM[5]) );
  XOR2_X1 U733 ( .A(n329), .B(n35), .Z(SUM[6]) );
  XOR2_X1 U734 ( .A(n258), .B(n24), .Z(SUM[17]) );
  NAND2_X1 U735 ( .A1(n376), .A2(n257), .ZN(n24) );
  XOR2_X1 U736 ( .A(n249), .B(n23), .Z(SUM[18]) );
  NAND2_X1 U737 ( .A1(n246), .A2(n248), .ZN(n23) );
  XOR2_X1 U738 ( .A(n242), .B(n22), .Z(SUM[19]) );
  NAND2_X1 U739 ( .A1(n374), .A2(n241), .ZN(n22) );
  XOR2_X1 U740 ( .A(n273), .B(n26), .Z(SUM[15]) );
  XOR2_X1 U741 ( .A(n287), .B(n28), .Z(SUM[13]) );
  XNOR2_X1 U742 ( .A(n292), .B(n29), .ZN(SUM[12]) );
  XOR2_X1 U743 ( .A(n303), .B(n30), .Z(SUM[11]) );
  XNOR2_X1 U744 ( .A(n308), .B(n31), .ZN(SUM[10]) );
  XNOR2_X1 U745 ( .A(n315), .B(n32), .ZN(SUM[9]) );
  XOR2_X1 U746 ( .A(n318), .B(n33), .Z(SUM[8]) );
  XNOR2_X1 U747 ( .A(n326), .B(n34), .ZN(SUM[7]) );
  OR2_X1 U748 ( .A1(A[39]), .A2(B[39]), .ZN(n569) );
  NOR2_X1 U749 ( .A1(n227), .A2(n220), .ZN(n218) );
  INV_X1 U750 ( .A(n543), .ZN(n226) );
  NOR2_X1 U751 ( .A1(B[20]), .A2(A[20]), .ZN(n227) );
  NAND2_X1 U752 ( .A1(n167), .A2(n170), .ZN(n15) );
  INV_X1 U753 ( .A(n170), .ZN(n168) );
  OAI21_X1 U754 ( .B1(n190), .B2(n546), .A(n183), .ZN(n181) );
  NAND2_X1 U755 ( .A1(A[34]), .A2(B[34]), .ZN(n90) );
  INV_X1 U756 ( .A(n550), .ZN(n124) );
  NAND2_X1 U757 ( .A1(A[23]), .A2(B[23]), .ZN(n203) );
  NAND2_X1 U758 ( .A1(A[35]), .A2(B[35]), .ZN(n83) );
  INV_X1 U759 ( .A(n554), .ZN(n208) );
  NAND2_X1 U760 ( .A1(A[33]), .A2(B[33]), .ZN(n99) );
  NAND2_X1 U761 ( .A1(A[36]), .A2(B[36]), .ZN(n70) );
  NOR2_X1 U762 ( .A1(n169), .A2(n160), .ZN(n158) );
  AOI21_X1 U763 ( .B1(n55), .B2(n528), .A(n50), .ZN(n48) );
  OAI21_X1 U764 ( .B1(n79), .B2(n56), .A(n57), .ZN(n55) );
  NAND2_X1 U765 ( .A1(B[31]), .A2(A[31]), .ZN(n115) );
  NOR2_X1 U766 ( .A1(A[31]), .A2(B[31]), .ZN(n114) );
  INV_X1 U767 ( .A(n537), .ZN(n145) );
  XOR2_X1 U768 ( .A(n211), .B(n19), .Z(SUM[22]) );
  OAI21_X1 U769 ( .B1(n215), .B2(n554), .A(n210), .ZN(n206) );
  OAI21_X1 U770 ( .B1(n240), .B2(n248), .A(n241), .ZN(n239) );
  NOR2_X1 U771 ( .A1(A[32]), .A2(B[32]), .ZN(n103) );
  NAND2_X1 U772 ( .A1(A[32]), .A2(B[32]), .ZN(n104) );
  NAND2_X1 U773 ( .A1(n218), .A2(n200), .ZN(n198) );
  NAND2_X1 U774 ( .A1(A[21]), .A2(B[21]), .ZN(n221) );
  XOR2_X1 U775 ( .A(n204), .B(n18), .Z(SUM[23]) );
  XNOR2_X1 U776 ( .A(n263), .B(n25), .ZN(SUM[16]) );
  AOI21_X1 U777 ( .B1(n263), .B2(n254), .A(n255), .ZN(n249) );
  AOI21_X1 U778 ( .B1(n263), .B2(n243), .A(n244), .ZN(n242) );
  AOI21_X1 U779 ( .B1(n263), .B2(n234), .A(n235), .ZN(n229) );
  AOI21_X1 U780 ( .B1(n263), .B2(n223), .A(n224), .ZN(n222) );
  AOI21_X1 U781 ( .B1(n263), .B2(n212), .A(n213), .ZN(n211) );
  AOI21_X1 U782 ( .B1(n263), .B2(n205), .A(n206), .ZN(n204) );
  AOI21_X1 U783 ( .B1(n263), .B2(n192), .A(n193), .ZN(n191) );
  AOI21_X1 U784 ( .B1(n263), .B2(n185), .A(n186), .ZN(n184) );
  AOI21_X1 U785 ( .B1(n263), .B2(n172), .A(n173), .ZN(n171) );
  AOI21_X1 U786 ( .B1(n263), .B2(n163), .A(n164), .ZN(n162) );
  AOI21_X1 U787 ( .B1(n263), .B2(n377), .A(n260), .ZN(n258) );
  OAI21_X1 U788 ( .B1(n271), .B2(n277), .A(n272), .ZN(n270) );
  AOI21_X1 U789 ( .B1(n263), .B2(n150), .A(n151), .ZN(n149) );
  NOR2_X1 U790 ( .A1(n156), .A2(n110), .ZN(n108) );
  NAND2_X1 U791 ( .A1(A[26]), .A2(B[26]), .ZN(n170) );
  AOI21_X1 U792 ( .B1(n263), .B2(n117), .A(n118), .ZN(n116) );
  NAND2_X1 U793 ( .A1(B[30]), .A2(A[30]), .ZN(n126) );
  NOR2_X1 U794 ( .A1(B[30]), .A2(A[30]), .ZN(n125) );
  INV_X1 U795 ( .A(n539), .ZN(n195) );
  AOI21_X1 U796 ( .B1(n263), .B2(n128), .A(n129), .ZN(n127) );
  NAND2_X1 U797 ( .A1(B[25]), .A2(A[25]), .ZN(n183) );
  AOI21_X1 U798 ( .B1(n263), .B2(n141), .A(n142), .ZN(n140) );
  AOI21_X1 U799 ( .B1(n158), .B2(n181), .A(n159), .ZN(n157) );
  NOR2_X1 U800 ( .A1(A[24]), .A2(B[24]), .ZN(n189) );
  NAND2_X1 U801 ( .A1(A[24]), .A2(B[24]), .ZN(n190) );
  OAI21_X1 U802 ( .B1(n106), .B2(n264), .A(n107), .ZN(n105) );
  AOI21_X1 U803 ( .B1(n200), .B2(n219), .A(n201), .ZN(n199) );
  OAI21_X1 U804 ( .B1(n202), .B2(n210), .A(n203), .ZN(n201) );
  NOR2_X1 U805 ( .A1(n209), .A2(n202), .ZN(n200) );
  NOR2_X1 U806 ( .A1(n542), .A2(n119), .ZN(n117) );
  NOR2_X1 U807 ( .A1(n542), .A2(n187), .ZN(n185) );
  NOR2_X1 U808 ( .A1(n542), .A2(n178), .ZN(n172) );
  NOR2_X1 U809 ( .A1(n542), .A2(n165), .ZN(n163) );
  NOR2_X1 U810 ( .A1(n542), .A2(n152), .ZN(n150) );
  NOR2_X1 U811 ( .A1(n542), .A2(n143), .ZN(n141) );
  NOR2_X1 U812 ( .A1(n542), .A2(n130), .ZN(n128) );
  NOR2_X1 U813 ( .A1(B[22]), .A2(A[22]), .ZN(n209) );
  OAI21_X1 U814 ( .B1(n195), .B2(n178), .A(n179), .ZN(n173) );
  OAI21_X1 U815 ( .B1(n195), .B2(n152), .A(n153), .ZN(n151) );
  OAI21_X1 U816 ( .B1(n195), .B2(n165), .A(n166), .ZN(n164) );
  OAI21_X1 U817 ( .B1(n195), .B2(n143), .A(n144), .ZN(n142) );
  OAI21_X1 U818 ( .B1(n195), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U819 ( .B1(n195), .B2(n119), .A(n120), .ZN(n118) );
  OAI21_X1 U820 ( .B1(n195), .B2(n187), .A(n190), .ZN(n186) );
  OAI21_X1 U821 ( .B1(n220), .B2(n228), .A(n221), .ZN(n219) );
  AOI21_X1 U822 ( .B1(n121), .B2(n155), .A(n122), .ZN(n120) );
  NAND2_X1 U823 ( .A1(n180), .A2(n545), .ZN(n156) );
  NOR2_X1 U824 ( .A1(n89), .A2(n82), .ZN(n80) );
  OAI21_X1 U825 ( .B1(n82), .B2(n90), .A(n83), .ZN(n81) );
  NAND2_X1 U826 ( .A1(n96), .A2(n80), .ZN(n78) );
  NOR2_X1 U827 ( .A1(n103), .A2(n98), .ZN(n96) );
  AOI21_X1 U828 ( .B1(n523), .B2(n539), .A(n109), .ZN(n107) );
  NAND2_X1 U829 ( .A1(n108), .A2(n196), .ZN(n106) );
  OAI21_X1 U830 ( .B1(n548), .B2(n170), .A(n161), .ZN(n159) );
  NAND2_X1 U831 ( .A1(B[27]), .A2(A[27]), .ZN(n161) );
  NOR2_X1 U832 ( .A1(A[27]), .A2(B[27]), .ZN(n160) );
  OAI21_X1 U833 ( .B1(n157), .B2(n110), .A(n111), .ZN(n109) );
  NOR2_X1 U834 ( .A1(B[28]), .A2(A[28]), .ZN(n147) );
  AOI21_X1 U835 ( .B1(n553), .B2(n137), .A(n113), .ZN(n111) );
  NAND2_X1 U836 ( .A1(n112), .A2(n136), .ZN(n110) );
  NOR2_X1 U837 ( .A1(n114), .A2(n125), .ZN(n112) );
  XNOR2_X1 U838 ( .A(n1), .B(n9), .ZN(SUM[32]) );
  AOI21_X1 U839 ( .B1(n521), .B2(n531), .A(n46), .ZN(n44) );
  AOI21_X1 U840 ( .B1(n568), .B2(n76), .A(n77), .ZN(n71) );
  AOI21_X1 U841 ( .B1(n1), .B2(n96), .A(n93), .ZN(n91) );
  AOI21_X1 U842 ( .B1(n568), .B2(n63), .A(n64), .ZN(n62) );
  AOI21_X1 U843 ( .B1(n521), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U844 ( .B1(n521), .B2(n54), .A(n55), .ZN(n53) );
  AOI21_X1 U845 ( .B1(n568), .B2(n361), .A(n102), .ZN(n100) );
  OAI21_X1 U846 ( .B1(n552), .B2(n148), .A(n139), .ZN(n137) );
  NAND2_X1 U847 ( .A1(B[29]), .A2(A[29]), .ZN(n139) );
  OAI21_X1 U848 ( .B1(n558), .B2(n126), .A(n115), .ZN(n113) );
endmodule


module datapath_DW01_add_10 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n43, n44, n46, n48, n50, n52, n53, n54, n55, n56,
         n57, n59, n61, n62, n63, n64, n67, n68, n69, n70, n71, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n226, n227, n228, n229, n230, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n246, n247,
         n248, n249, n252, n253, n254, n255, n256, n257, n258, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n275, n276, n277, n278, n279, n280, n283, n284, n285, n286,
         n287, n289, n290, n291, n292, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n353, n358, n360, n361, n362, n364,
         n366, n368, n370, n372, n374, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n551, n552, n553;

  INV_X1 U437 ( .A(n197), .ZN(n520) );
  NOR2_X1 U438 ( .A1(n110), .A2(n156), .ZN(n521) );
  NOR2_X1 U439 ( .A1(A[19]), .A2(B[19]), .ZN(n240) );
  NOR2_X1 U440 ( .A1(n247), .A2(n240), .ZN(n238) );
  OAI21_X1 U441 ( .B1(n79), .B2(n56), .A(n57), .ZN(n522) );
  CLKBUF_X1 U442 ( .A(B[32]), .Z(n523) );
  OR2_X1 U443 ( .A1(A[37]), .A2(B[37]), .ZN(n524) );
  OR2_X1 U444 ( .A1(A[38]), .A2(B[38]), .ZN(n525) );
  NOR2_X1 U445 ( .A1(n189), .A2(n531), .ZN(n526) );
  NOR2_X1 U446 ( .A1(A[20]), .A2(B[20]), .ZN(n227) );
  AND2_X1 U447 ( .A1(n54), .A2(n525), .ZN(n527) );
  NOR2_X1 U448 ( .A1(A[18]), .A2(B[18]), .ZN(n247) );
  CLKBUF_X1 U449 ( .A(n147), .Z(n528) );
  NOR2_X1 U450 ( .A1(A[33]), .A2(B[33]), .ZN(n529) );
  NOR2_X1 U451 ( .A1(A[35]), .A2(B[35]), .ZN(n530) );
  CLKBUF_X1 U452 ( .A(n182), .Z(n531) );
  NOR2_X1 U453 ( .A1(n160), .A2(n169), .ZN(n532) );
  CLKBUF_X1 U454 ( .A(n160), .Z(n533) );
  OR2_X1 U455 ( .A1(n147), .A2(n138), .ZN(n534) );
  NOR2_X1 U456 ( .A1(n125), .A2(n537), .ZN(n535) );
  NOR2_X1 U457 ( .A1(A[29]), .A2(B[29]), .ZN(n536) );
  NOR2_X1 U458 ( .A1(B[31]), .A2(A[31]), .ZN(n537) );
  CLKBUF_X1 U459 ( .A(n169), .Z(n538) );
  NOR2_X1 U460 ( .A1(A[27]), .A2(B[27]), .ZN(n539) );
  OAI21_X1 U461 ( .B1(n106), .B2(n264), .A(n107), .ZN(n540) );
  OAI21_X1 U462 ( .B1(n106), .B2(n264), .A(n107), .ZN(n105) );
  CLKBUF_X1 U463 ( .A(n181), .Z(n541) );
  NOR2_X1 U464 ( .A1(A[25]), .A2(B[25]), .ZN(n542) );
  XNOR2_X1 U465 ( .A(n62), .B(n543), .ZN(SUM[37]) );
  AND2_X1 U466 ( .A1(n524), .A2(n61), .ZN(n543) );
  XNOR2_X1 U467 ( .A(n71), .B(n544), .ZN(SUM[36]) );
  AND2_X1 U468 ( .A1(n67), .A2(n70), .ZN(n544) );
  XNOR2_X1 U469 ( .A(n84), .B(n545), .ZN(SUM[35]) );
  AND2_X1 U470 ( .A1(n358), .A2(n83), .ZN(n545) );
  XNOR2_X1 U471 ( .A(n91), .B(n546), .ZN(SUM[34]) );
  AND2_X1 U472 ( .A1(n88), .A2(n90), .ZN(n546) );
  XNOR2_X1 U473 ( .A(n100), .B(n547), .ZN(SUM[33]) );
  AND2_X1 U474 ( .A1(n360), .A2(n99), .ZN(n547) );
  XNOR2_X1 U475 ( .A(n53), .B(n548), .ZN(SUM[38]) );
  AND2_X1 U476 ( .A1(n525), .A2(n52), .ZN(n548) );
  CLKBUF_X1 U477 ( .A(n536), .Z(n549) );
  AOI21_X1 U478 ( .B1(n238), .B2(n255), .A(n239), .ZN(n237) );
  NOR2_X1 U479 ( .A1(A[4]), .A2(B[4]), .ZN(n337) );
  NOR2_X1 U480 ( .A1(A[10]), .A2(B[10]), .ZN(n306) );
  NOR2_X1 U481 ( .A1(A[12]), .A2(B[12]), .ZN(n290) );
  NOR2_X1 U482 ( .A1(A[16]), .A2(B[16]), .ZN(n261) );
  NOR2_X1 U483 ( .A1(A[6]), .A2(B[6]), .ZN(n327) );
  NOR2_X1 U484 ( .A1(A[7]), .A2(B[7]), .ZN(n324) );
  NOR2_X1 U485 ( .A1(A[13]), .A2(B[13]), .ZN(n285) );
  NOR2_X1 U486 ( .A1(A[11]), .A2(B[11]), .ZN(n301) );
  NOR2_X1 U487 ( .A1(A[9]), .A2(B[9]), .ZN(n313) );
  NOR2_X1 U488 ( .A1(A[5]), .A2(B[5]), .ZN(n332) );
  NOR2_X1 U489 ( .A1(A[3]), .A2(B[3]), .ZN(n343) );
  NOR2_X1 U490 ( .A1(A[8]), .A2(B[8]), .ZN(n316) );
  NOR2_X1 U491 ( .A1(A[2]), .A2(B[2]), .ZN(n346) );
  NOR2_X1 U492 ( .A1(A[1]), .A2(B[1]), .ZN(n350) );
  OR2_X1 U493 ( .A1(A[39]), .A2(B[39]), .ZN(n553) );
  INV_X1 U494 ( .A(n236), .ZN(n230) );
  INV_X1 U495 ( .A(n214), .ZN(n212) );
  INV_X1 U496 ( .A(n215), .ZN(n213) );
  INV_X1 U497 ( .A(n520), .ZN(n193) );
  INV_X1 U498 ( .A(n526), .ZN(n174) );
  NAND2_X1 U499 ( .A1(n154), .A2(n132), .ZN(n130) );
  INV_X1 U500 ( .A(n94), .ZN(n92) );
  INV_X1 U501 ( .A(n95), .ZN(n93) );
  INV_X1 U502 ( .A(n156), .ZN(n154) );
  OAI21_X1 U503 ( .B1(n318), .B2(n297), .A(n298), .ZN(n292) );
  INV_X1 U504 ( .A(n264), .ZN(n263) );
  NOR2_X1 U505 ( .A1(n78), .A2(n56), .ZN(n54) );
  AOI21_X1 U506 ( .B1(n155), .B2(n132), .A(n133), .ZN(n131) );
  INV_X1 U507 ( .A(n135), .ZN(n133) );
  NAND2_X1 U508 ( .A1(n230), .A2(n216), .ZN(n214) );
  NOR2_X1 U509 ( .A1(n236), .A2(n198), .ZN(n196) );
  INV_X1 U510 ( .A(n534), .ZN(n132) );
  INV_X1 U511 ( .A(n76), .ZN(n74) );
  INV_X1 U512 ( .A(n297), .ZN(n295) );
  NAND2_X1 U513 ( .A1(n121), .A2(n154), .ZN(n119) );
  NAND2_X1 U514 ( .A1(n526), .A2(n167), .ZN(n165) );
  AOI21_X1 U515 ( .B1(n339), .B2(n330), .A(n331), .ZN(n329) );
  NOR2_X1 U516 ( .A1(n74), .A2(n69), .ZN(n63) );
  INV_X1 U517 ( .A(n197), .ZN(n195) );
  AOI21_X1 U518 ( .B1(n319), .B2(n265), .A(n266), .ZN(n264) );
  OAI21_X1 U519 ( .B1(n298), .B2(n267), .A(n268), .ZN(n266) );
  NOR2_X1 U520 ( .A1(n297), .A2(n267), .ZN(n265) );
  AOI21_X1 U521 ( .B1(n269), .B2(n284), .A(n270), .ZN(n268) );
  OAI21_X1 U522 ( .B1(n318), .B2(n279), .A(n280), .ZN(n278) );
  AOI21_X1 U523 ( .B1(n296), .B2(n283), .A(n284), .ZN(n280) );
  NAND2_X1 U524 ( .A1(n295), .A2(n283), .ZN(n279) );
  OAI21_X1 U525 ( .B1(n318), .B2(n309), .A(n310), .ZN(n308) );
  INV_X1 U526 ( .A(n312), .ZN(n310) );
  INV_X1 U527 ( .A(n311), .ZN(n309) );
  INV_X1 U528 ( .A(n79), .ZN(n77) );
  AOI21_X1 U529 ( .B1(n235), .B2(n216), .A(n219), .ZN(n215) );
  INV_X1 U530 ( .A(n319), .ZN(n318) );
  NAND2_X1 U531 ( .A1(n154), .A2(n145), .ZN(n143) );
  INV_X1 U532 ( .A(n96), .ZN(n94) );
  INV_X1 U533 ( .A(n137), .ZN(n135) );
  INV_X1 U534 ( .A(n97), .ZN(n95) );
  INV_X1 U535 ( .A(n157), .ZN(n155) );
  INV_X1 U536 ( .A(n255), .ZN(n253) );
  NAND2_X1 U537 ( .A1(n254), .A2(n238), .ZN(n236) );
  NOR2_X1 U538 ( .A1(n534), .A2(n123), .ZN(n121) );
  NAND2_X1 U539 ( .A1(n283), .A2(n269), .ZN(n267) );
  NAND2_X1 U540 ( .A1(n311), .A2(n299), .ZN(n297) );
  INV_X1 U541 ( .A(n340), .ZN(n339) );
  INV_X1 U542 ( .A(n254), .ZN(n252) );
  INV_X1 U543 ( .A(n237), .ZN(n235) );
  INV_X1 U544 ( .A(n298), .ZN(n296) );
  INV_X1 U545 ( .A(n349), .ZN(n348) );
  INV_X1 U546 ( .A(n217), .ZN(n216) );
  INV_X1 U547 ( .A(n218), .ZN(n217) );
  NAND2_X1 U548 ( .A1(n67), .A2(n524), .ZN(n56) );
  INV_X1 U549 ( .A(n48), .ZN(n46) );
  NOR2_X1 U550 ( .A1(n276), .A2(n271), .ZN(n269) );
  NOR2_X1 U551 ( .A1(n261), .A2(n256), .ZN(n254) );
  INV_X1 U552 ( .A(n262), .ZN(n260) );
  NOR2_X1 U553 ( .A1(n252), .A2(n247), .ZN(n243) );
  OAI21_X1 U554 ( .B1(n253), .B2(n247), .A(n248), .ZN(n244) );
  AOI21_X1 U555 ( .B1(n299), .B2(n312), .A(n300), .ZN(n298) );
  OAI21_X1 U556 ( .B1(n301), .B2(n307), .A(n302), .ZN(n300) );
  AOI21_X1 U557 ( .B1(n341), .B2(n349), .A(n342), .ZN(n340) );
  NOR2_X1 U558 ( .A1(n346), .A2(n343), .ZN(n341) );
  OAI21_X1 U559 ( .B1(n343), .B2(n347), .A(n344), .ZN(n342) );
  AOI21_X1 U560 ( .B1(n524), .B2(n68), .A(n59), .ZN(n57) );
  INV_X1 U561 ( .A(n61), .ZN(n59) );
  OAI21_X1 U562 ( .B1(n332), .B2(n338), .A(n333), .ZN(n331) );
  AOI21_X1 U563 ( .B1(n80), .B2(n97), .A(n81), .ZN(n79) );
  OAI21_X1 U564 ( .B1(n313), .B2(n317), .A(n314), .ZN(n312) );
  OAI21_X1 U565 ( .B1(n285), .B2(n291), .A(n286), .ZN(n284) );
  OAI21_X1 U566 ( .B1(n350), .B2(n353), .A(n351), .ZN(n349) );
  OAI21_X1 U567 ( .B1(n340), .B2(n320), .A(n321), .ZN(n319) );
  AOI21_X1 U568 ( .B1(n322), .B2(n331), .A(n323), .ZN(n321) );
  NAND2_X1 U569 ( .A1(n330), .A2(n322), .ZN(n320) );
  OAI21_X1 U570 ( .B1(n324), .B2(n328), .A(n325), .ZN(n323) );
  NOR2_X1 U571 ( .A1(n94), .A2(n87), .ZN(n85) );
  OAI21_X1 U572 ( .B1(n95), .B2(n87), .A(n90), .ZN(n86) );
  INV_X1 U573 ( .A(n88), .ZN(n87) );
  NOR2_X1 U574 ( .A1(n236), .A2(n227), .ZN(n223) );
  OAI21_X1 U575 ( .B1(n237), .B2(n227), .A(n228), .ZN(n224) );
  INV_X1 U576 ( .A(n188), .ZN(n187) );
  NOR2_X1 U577 ( .A1(n327), .A2(n324), .ZN(n322) );
  NOR2_X1 U578 ( .A1(n337), .A2(n332), .ZN(n330) );
  NOR2_X1 U579 ( .A1(n316), .A2(n313), .ZN(n311) );
  NOR2_X1 U580 ( .A1(n306), .A2(n301), .ZN(n299) );
  OAI21_X1 U581 ( .B1(n135), .B2(n123), .A(n126), .ZN(n122) );
  INV_X1 U582 ( .A(n148), .ZN(n146) );
  NOR2_X1 U583 ( .A1(n290), .A2(n285), .ZN(n283) );
  NOR2_X1 U584 ( .A1(n227), .A2(n220), .ZN(n218) );
  AOI21_X1 U585 ( .B1(n292), .B2(n381), .A(n289), .ZN(n287) );
  INV_X1 U586 ( .A(n291), .ZN(n289) );
  AOI21_X1 U587 ( .B1(n308), .B2(n383), .A(n305), .ZN(n303) );
  INV_X1 U588 ( .A(n307), .ZN(n305) );
  AOI21_X1 U589 ( .B1(n278), .B2(n379), .A(n275), .ZN(n273) );
  INV_X1 U590 ( .A(n277), .ZN(n275) );
  XOR2_X1 U591 ( .A(n329), .B(n35), .Z(SUM[6]) );
  NAND2_X1 U592 ( .A1(n387), .A2(n328), .ZN(n35) );
  INV_X1 U593 ( .A(n227), .ZN(n226) );
  INV_X1 U594 ( .A(n69), .ZN(n67) );
  INV_X1 U595 ( .A(n209), .ZN(n208) );
  NOR2_X1 U596 ( .A1(n209), .A2(n202), .ZN(n200) );
  OAI21_X1 U597 ( .B1(n318), .B2(n316), .A(n317), .ZN(n315) );
  AOI21_X1 U598 ( .B1(n541), .B2(n167), .A(n168), .ZN(n166) );
  INV_X1 U599 ( .A(n170), .ZN(n168) );
  INV_X1 U600 ( .A(n189), .ZN(n188) );
  INV_X1 U601 ( .A(n202), .ZN(n370) );
  INV_X1 U602 ( .A(n220), .ZN(n372) );
  INV_X1 U603 ( .A(n537), .ZN(n362) );
  INV_X1 U604 ( .A(n103), .ZN(n361) );
  INV_X1 U605 ( .A(n124), .ZN(n123) );
  INV_X1 U606 ( .A(n125), .ZN(n124) );
  INV_X1 U607 ( .A(n70), .ZN(n68) );
  INV_X1 U608 ( .A(n247), .ZN(n246) );
  INV_X1 U609 ( .A(n89), .ZN(n88) );
  INV_X1 U610 ( .A(n530), .ZN(n358) );
  NOR2_X1 U611 ( .A1(n214), .A2(n207), .ZN(n205) );
  INV_X1 U612 ( .A(n208), .ZN(n207) );
  INV_X1 U613 ( .A(n327), .ZN(n387) );
  INV_X1 U614 ( .A(n316), .ZN(n385) );
  INV_X1 U615 ( .A(n346), .ZN(n391) );
  INV_X1 U616 ( .A(n285), .ZN(n380) );
  INV_X1 U617 ( .A(n337), .ZN(n389) );
  INV_X1 U618 ( .A(n301), .ZN(n382) );
  INV_X1 U619 ( .A(n313), .ZN(n384) );
  INV_X1 U620 ( .A(n290), .ZN(n381) );
  INV_X1 U621 ( .A(n306), .ZN(n383) );
  NAND2_X1 U622 ( .A1(n386), .A2(n325), .ZN(n34) );
  INV_X1 U623 ( .A(n324), .ZN(n386) );
  NAND2_X1 U624 ( .A1(n388), .A2(n333), .ZN(n36) );
  INV_X1 U625 ( .A(n332), .ZN(n388) );
  INV_X1 U626 ( .A(n240), .ZN(n374) );
  NAND2_X1 U627 ( .A1(n390), .A2(n344), .ZN(n38) );
  INV_X1 U628 ( .A(n343), .ZN(n390) );
  XOR2_X1 U629 ( .A(n287), .B(n28), .Z(SUM[13]) );
  NAND2_X1 U630 ( .A1(n380), .A2(n286), .ZN(n28) );
  XNOR2_X1 U631 ( .A(n292), .B(n29), .ZN(SUM[12]) );
  NAND2_X1 U632 ( .A1(n381), .A2(n291), .ZN(n29) );
  XOR2_X1 U633 ( .A(n303), .B(n30), .Z(SUM[11]) );
  NAND2_X1 U634 ( .A1(n382), .A2(n302), .ZN(n30) );
  INV_X1 U635 ( .A(n350), .ZN(n392) );
  NAND2_X1 U636 ( .A1(n378), .A2(n272), .ZN(n26) );
  INV_X1 U637 ( .A(n271), .ZN(n378) );
  INV_X1 U638 ( .A(n533), .ZN(n366) );
  INV_X1 U639 ( .A(n529), .ZN(n360) );
  INV_X1 U640 ( .A(n531), .ZN(n368) );
  INV_X1 U641 ( .A(n338), .ZN(n336) );
  NAND2_X1 U642 ( .A1(n377), .A2(n262), .ZN(n25) );
  INV_X1 U643 ( .A(n261), .ZN(n377) );
  XNOR2_X1 U644 ( .A(n278), .B(n27), .ZN(SUM[14]) );
  NAND2_X1 U645 ( .A1(n379), .A2(n277), .ZN(n27) );
  XOR2_X1 U646 ( .A(n40), .B(n353), .Z(SUM[1]) );
  NAND2_X1 U647 ( .A1(n392), .A2(n351), .ZN(n40) );
  XNOR2_X1 U648 ( .A(n345), .B(n38), .ZN(SUM[3]) );
  OAI21_X1 U649 ( .B1(n348), .B2(n346), .A(n347), .ZN(n345) );
  XNOR2_X1 U650 ( .A(n339), .B(n37), .ZN(SUM[4]) );
  NAND2_X1 U651 ( .A1(n389), .A2(n338), .ZN(n37) );
  XNOR2_X1 U652 ( .A(n308), .B(n31), .ZN(SUM[10]) );
  NAND2_X1 U653 ( .A1(n383), .A2(n307), .ZN(n31) );
  XNOR2_X1 U654 ( .A(n315), .B(n32), .ZN(SUM[9]) );
  NAND2_X1 U655 ( .A1(n384), .A2(n314), .ZN(n32) );
  XOR2_X1 U656 ( .A(n318), .B(n33), .Z(SUM[8]) );
  NAND2_X1 U657 ( .A1(n385), .A2(n317), .ZN(n33) );
  XNOR2_X1 U658 ( .A(n326), .B(n34), .ZN(SUM[7]) );
  OAI21_X1 U659 ( .B1(n329), .B2(n327), .A(n328), .ZN(n326) );
  XOR2_X1 U660 ( .A(n334), .B(n36), .Z(SUM[5]) );
  AOI21_X1 U661 ( .B1(n339), .B2(n389), .A(n336), .ZN(n334) );
  AND2_X1 U662 ( .A1(n551), .A2(n353), .ZN(SUM[0]) );
  XOR2_X1 U663 ( .A(n348), .B(n39), .Z(SUM[2]) );
  NAND2_X1 U664 ( .A1(n391), .A2(n347), .ZN(n39) );
  INV_X1 U665 ( .A(n52), .ZN(n50) );
  OR2_X1 U666 ( .A1(A[0]), .A2(B[0]), .ZN(n551) );
  NOR2_X1 U667 ( .A1(A[34]), .A2(B[34]), .ZN(n89) );
  NOR2_X1 U668 ( .A1(B[25]), .A2(A[25]), .ZN(n182) );
  NOR2_X1 U669 ( .A1(A[33]), .A2(B[33]), .ZN(n98) );
  NOR2_X1 U670 ( .A1(B[27]), .A2(A[27]), .ZN(n160) );
  NOR2_X1 U671 ( .A1(A[36]), .A2(B[36]), .ZN(n69) );
  NOR2_X1 U672 ( .A1(A[17]), .A2(B[17]), .ZN(n256) );
  NOR2_X1 U673 ( .A1(A[35]), .A2(B[35]), .ZN(n82) );
  NAND2_X1 U674 ( .A1(n368), .A2(n183), .ZN(n16) );
  NAND2_X1 U675 ( .A1(n364), .A2(n139), .ZN(n12) );
  NAND2_X1 U676 ( .A1(n145), .A2(n148), .ZN(n13) );
  NOR2_X1 U677 ( .A1(A[15]), .A2(B[15]), .ZN(n271) );
  NAND2_X1 U678 ( .A1(A[36]), .A2(B[36]), .ZN(n70) );
  NAND2_X1 U679 ( .A1(A[37]), .A2(B[37]), .ZN(n61) );
  NAND2_X1 U680 ( .A1(A[6]), .A2(B[6]), .ZN(n328) );
  NAND2_X1 U681 ( .A1(A[8]), .A2(B[8]), .ZN(n317) );
  XOR2_X1 U682 ( .A(n211), .B(n19), .Z(SUM[22]) );
  NAND2_X1 U683 ( .A1(n208), .A2(n210), .ZN(n19) );
  XOR2_X1 U684 ( .A(n191), .B(n17), .Z(SUM[24]) );
  NAND2_X1 U685 ( .A1(n188), .A2(n190), .ZN(n17) );
  XOR2_X1 U686 ( .A(n229), .B(n21), .Z(SUM[20]) );
  NAND2_X1 U687 ( .A1(n226), .A2(n228), .ZN(n21) );
  NAND2_X1 U688 ( .A1(A[4]), .A2(B[4]), .ZN(n338) );
  NAND2_X1 U689 ( .A1(A[5]), .A2(B[5]), .ZN(n333) );
  NAND2_X1 U690 ( .A1(A[7]), .A2(B[7]), .ZN(n325) );
  NAND2_X1 U691 ( .A1(A[12]), .A2(B[12]), .ZN(n291) );
  NAND2_X1 U692 ( .A1(A[10]), .A2(B[10]), .ZN(n307) );
  NAND2_X1 U693 ( .A1(A[2]), .A2(B[2]), .ZN(n347) );
  NAND2_X1 U694 ( .A1(A[0]), .A2(B[0]), .ZN(n353) );
  NAND2_X1 U695 ( .A1(A[18]), .A2(B[18]), .ZN(n248) );
  NAND2_X1 U696 ( .A1(A[16]), .A2(B[16]), .ZN(n262) );
  NAND2_X1 U697 ( .A1(A[38]), .A2(B[38]), .ZN(n52) );
  NAND2_X1 U698 ( .A1(A[26]), .A2(B[26]), .ZN(n170) );
  NAND2_X1 U699 ( .A1(A[34]), .A2(B[34]), .ZN(n90) );
  NAND2_X1 U700 ( .A1(A[14]), .A2(B[14]), .ZN(n277) );
  NAND2_X1 U701 ( .A1(A[13]), .A2(B[13]), .ZN(n286) );
  NAND2_X1 U702 ( .A1(A[11]), .A2(B[11]), .ZN(n302) );
  NAND2_X1 U703 ( .A1(A[9]), .A2(B[9]), .ZN(n314) );
  NAND2_X1 U704 ( .A1(A[3]), .A2(B[3]), .ZN(n344) );
  NAND2_X1 U705 ( .A1(A[1]), .A2(B[1]), .ZN(n351) );
  NAND2_X1 U706 ( .A1(A[39]), .A2(B[39]), .ZN(n43) );
  NAND2_X1 U707 ( .A1(A[15]), .A2(B[15]), .ZN(n272) );
  NAND2_X1 U708 ( .A1(A[17]), .A2(B[17]), .ZN(n257) );
  XNOR2_X1 U709 ( .A(n44), .B(n552), .ZN(SUM[39]) );
  AND2_X1 U710 ( .A1(n553), .A2(n43), .ZN(n552) );
  XOR2_X1 U711 ( .A(n116), .B(n10), .Z(SUM[31]) );
  NAND2_X1 U712 ( .A1(n362), .A2(n115), .ZN(n10) );
  NAND2_X1 U713 ( .A1(n372), .A2(n221), .ZN(n20) );
  XOR2_X1 U714 ( .A(n171), .B(n15), .Z(SUM[26]) );
  NAND2_X1 U715 ( .A1(n167), .A2(n170), .ZN(n15) );
  XOR2_X1 U716 ( .A(n162), .B(n14), .Z(SUM[27]) );
  NAND2_X1 U717 ( .A1(n366), .A2(n161), .ZN(n14) );
  XOR2_X1 U718 ( .A(n258), .B(n24), .Z(SUM[17]) );
  NAND2_X1 U719 ( .A1(n376), .A2(n257), .ZN(n24) );
  XOR2_X1 U720 ( .A(n249), .B(n23), .Z(SUM[18]) );
  NAND2_X1 U721 ( .A1(n246), .A2(n248), .ZN(n23) );
  XOR2_X1 U722 ( .A(n242), .B(n22), .Z(SUM[19]) );
  NAND2_X1 U723 ( .A1(n374), .A2(n241), .ZN(n22) );
  NAND2_X1 U724 ( .A1(n124), .A2(n126), .ZN(n11) );
  NAND2_X1 U725 ( .A1(n370), .A2(n203), .ZN(n18) );
  XOR2_X1 U726 ( .A(n273), .B(n26), .Z(SUM[15]) );
  NAND2_X1 U727 ( .A1(A[22]), .A2(B[22]), .ZN(n210) );
  NOR2_X1 U728 ( .A1(A[22]), .A2(B[22]), .ZN(n209) );
  INV_X1 U729 ( .A(n549), .ZN(n364) );
  INV_X1 U730 ( .A(n276), .ZN(n379) );
  NOR2_X1 U731 ( .A1(A[14]), .A2(B[14]), .ZN(n276) );
  NOR2_X1 U732 ( .A1(B[30]), .A2(A[30]), .ZN(n125) );
  NOR2_X1 U733 ( .A1(B[31]), .A2(A[31]), .ZN(n114) );
  INV_X1 U734 ( .A(n541), .ZN(n179) );
  AOI21_X1 U735 ( .B1(n532), .B2(n181), .A(n159), .ZN(n157) );
  INV_X1 U736 ( .A(n538), .ZN(n167) );
  NAND2_X1 U737 ( .A1(A[20]), .A2(B[20]), .ZN(n228) );
  AOI21_X1 U738 ( .B1(n200), .B2(n219), .A(n201), .ZN(n199) );
  OAI21_X1 U739 ( .B1(n75), .B2(n69), .A(n70), .ZN(n64) );
  INV_X1 U740 ( .A(n77), .ZN(n75) );
  OAI21_X1 U741 ( .B1(n98), .B2(n104), .A(n99), .ZN(n97) );
  INV_X1 U742 ( .A(n104), .ZN(n102) );
  NAND2_X1 U743 ( .A1(n361), .A2(n104), .ZN(n9) );
  NAND2_X1 U744 ( .A1(A[32]), .A2(B[32]), .ZN(n104) );
  NOR2_X1 U745 ( .A1(A[32]), .A2(n523), .ZN(n103) );
  OAI21_X1 U746 ( .B1(n256), .B2(n262), .A(n257), .ZN(n255) );
  INV_X1 U747 ( .A(n256), .ZN(n376) );
  XOR2_X1 U748 ( .A(n222), .B(n20), .Z(SUM[21]) );
  NAND2_X1 U749 ( .A1(A[35]), .A2(B[35]), .ZN(n83) );
  NAND2_X1 U750 ( .A1(n218), .A2(n200), .ZN(n198) );
  NAND2_X1 U751 ( .A1(A[21]), .A2(B[21]), .ZN(n221) );
  NOR2_X1 U752 ( .A1(A[21]), .A2(B[21]), .ZN(n220) );
  XOR2_X1 U753 ( .A(n204), .B(n18), .Z(SUM[23]) );
  OAI21_X1 U754 ( .B1(n215), .B2(n207), .A(n210), .ZN(n206) );
  OAI21_X1 U755 ( .B1(n240), .B2(n248), .A(n241), .ZN(n239) );
  NAND2_X1 U756 ( .A1(A[19]), .A2(B[19]), .ZN(n241) );
  NAND2_X1 U757 ( .A1(A[33]), .A2(B[33]), .ZN(n99) );
  NOR2_X1 U758 ( .A1(A[24]), .A2(B[24]), .ZN(n189) );
  NAND2_X1 U759 ( .A1(A[24]), .A2(B[24]), .ZN(n190) );
  XOR2_X1 U760 ( .A(n127), .B(n11), .Z(SUM[30]) );
  INV_X1 U761 ( .A(n528), .ZN(n145) );
  XNOR2_X1 U762 ( .A(n263), .B(n25), .ZN(SUM[16]) );
  AOI21_X1 U763 ( .B1(n263), .B2(n150), .A(n151), .ZN(n149) );
  AOI21_X1 U764 ( .B1(n263), .B2(n185), .A(n186), .ZN(n184) );
  AOI21_X1 U765 ( .B1(n263), .B2(n377), .A(n260), .ZN(n258) );
  AOI21_X1 U766 ( .B1(n263), .B2(n254), .A(n255), .ZN(n249) );
  AOI21_X1 U767 ( .B1(n263), .B2(n243), .A(n244), .ZN(n242) );
  AOI21_X1 U768 ( .B1(n263), .B2(n223), .A(n224), .ZN(n222) );
  AOI21_X1 U769 ( .B1(n263), .B2(n212), .A(n213), .ZN(n211) );
  AOI21_X1 U770 ( .B1(n263), .B2(n205), .A(n206), .ZN(n204) );
  AOI21_X1 U771 ( .B1(n263), .B2(n192), .A(n193), .ZN(n191) );
  AOI21_X1 U772 ( .B1(n263), .B2(n230), .A(n235), .ZN(n229) );
  OAI21_X1 U773 ( .B1(n271), .B2(n277), .A(n272), .ZN(n270) );
  AOI21_X1 U774 ( .B1(n263), .B2(n163), .A(n164), .ZN(n162) );
  NAND2_X1 U775 ( .A1(A[23]), .A2(B[23]), .ZN(n203) );
  NOR2_X1 U776 ( .A1(A[23]), .A2(B[23]), .ZN(n202) );
  AOI21_X1 U777 ( .B1(n263), .B2(n172), .A(n173), .ZN(n171) );
  XOR2_X1 U778 ( .A(n184), .B(n16), .Z(SUM[25]) );
  INV_X1 U779 ( .A(n194), .ZN(n192) );
  NAND2_X1 U780 ( .A1(B[25]), .A2(A[25]), .ZN(n183) );
  OAI21_X1 U781 ( .B1(n237), .B2(n198), .A(n199), .ZN(n197) );
  XOR2_X1 U782 ( .A(n149), .B(n13), .Z(SUM[28]) );
  INV_X1 U783 ( .A(n155), .ZN(n153) );
  AOI21_X1 U784 ( .B1(n55), .B2(n525), .A(n50), .ZN(n48) );
  OAI21_X1 U785 ( .B1(n79), .B2(n56), .A(n57), .ZN(n55) );
  INV_X1 U786 ( .A(n78), .ZN(n76) );
  NOR2_X1 U787 ( .A1(B[26]), .A2(A[26]), .ZN(n169) );
  INV_X1 U788 ( .A(n154), .ZN(n152) );
  INV_X1 U789 ( .A(n196), .ZN(n194) );
  AOI21_X1 U790 ( .B1(n263), .B2(n117), .A(n118), .ZN(n116) );
  AOI21_X1 U791 ( .B1(n263), .B2(n128), .A(n129), .ZN(n127) );
  NAND2_X1 U792 ( .A1(B[27]), .A2(A[27]), .ZN(n161) );
  XOR2_X1 U793 ( .A(n140), .B(n12), .Z(SUM[29]) );
  AOI21_X1 U794 ( .B1(n263), .B2(n141), .A(n142), .ZN(n140) );
  NAND2_X1 U795 ( .A1(B[31]), .A2(A[31]), .ZN(n115) );
  AOI21_X1 U796 ( .B1(n155), .B2(n145), .A(n146), .ZN(n144) );
  NOR2_X1 U797 ( .A1(n89), .A2(n530), .ZN(n80) );
  NOR2_X1 U798 ( .A1(n194), .A2(n152), .ZN(n150) );
  NOR2_X1 U799 ( .A1(n194), .A2(n143), .ZN(n141) );
  NOR2_X1 U800 ( .A1(n194), .A2(n130), .ZN(n128) );
  NOR2_X1 U801 ( .A1(n194), .A2(n119), .ZN(n117) );
  NOR2_X1 U802 ( .A1(n194), .A2(n174), .ZN(n172) );
  NOR2_X1 U803 ( .A1(n194), .A2(n165), .ZN(n163) );
  NOR2_X1 U804 ( .A1(n194), .A2(n187), .ZN(n185) );
  OAI21_X1 U805 ( .B1(n202), .B2(n210), .A(n203), .ZN(n201) );
  OAI21_X1 U806 ( .B1(n195), .B2(n152), .A(n153), .ZN(n151) );
  OAI21_X1 U807 ( .B1(n520), .B2(n143), .A(n144), .ZN(n142) );
  OAI21_X1 U808 ( .B1(n520), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U809 ( .B1(n195), .B2(n119), .A(n120), .ZN(n118) );
  OAI21_X1 U810 ( .B1(n195), .B2(n187), .A(n190), .ZN(n186) );
  OAI21_X1 U811 ( .B1(n520), .B2(n174), .A(n179), .ZN(n173) );
  OAI21_X1 U812 ( .B1(n195), .B2(n165), .A(n166), .ZN(n164) );
  OAI21_X1 U813 ( .B1(n220), .B2(n228), .A(n221), .ZN(n219) );
  NOR2_X1 U814 ( .A1(n110), .A2(n156), .ZN(n108) );
  NOR2_X1 U815 ( .A1(n160), .A2(n169), .ZN(n158) );
  NAND2_X1 U816 ( .A1(n96), .A2(n80), .ZN(n78) );
  OAI21_X1 U817 ( .B1(n82), .B2(n90), .A(n83), .ZN(n81) );
  NAND2_X1 U818 ( .A1(n158), .A2(n180), .ZN(n156) );
  NOR2_X1 U819 ( .A1(n189), .A2(n182), .ZN(n180) );
  NOR2_X1 U820 ( .A1(n103), .A2(n529), .ZN(n96) );
  AOI21_X1 U821 ( .B1(n121), .B2(n155), .A(n122), .ZN(n120) );
  NAND2_X1 U822 ( .A1(B[30]), .A2(A[30]), .ZN(n126) );
  NOR2_X1 U823 ( .A1(n138), .A2(n147), .ZN(n136) );
  NAND2_X1 U824 ( .A1(A[28]), .A2(B[28]), .ZN(n148) );
  NOR2_X1 U825 ( .A1(B[28]), .A2(A[28]), .ZN(n147) );
  AOI21_X1 U826 ( .B1(n521), .B2(n197), .A(n109), .ZN(n107) );
  NAND2_X1 U827 ( .A1(n108), .A2(n196), .ZN(n106) );
  NAND2_X1 U828 ( .A1(B[29]), .A2(A[29]), .ZN(n139) );
  NOR2_X1 U829 ( .A1(B[29]), .A2(A[29]), .ZN(n138) );
  OAI21_X1 U830 ( .B1(n157), .B2(n110), .A(n111), .ZN(n109) );
  OAI21_X1 U831 ( .B1(n539), .B2(n170), .A(n161), .ZN(n159) );
  AOI21_X1 U832 ( .B1(n535), .B2(n137), .A(n113), .ZN(n111) );
  NAND2_X1 U833 ( .A1(n112), .A2(n136), .ZN(n110) );
  NOR2_X1 U834 ( .A1(n114), .A2(n125), .ZN(n112) );
  OAI21_X1 U835 ( .B1(n542), .B2(n190), .A(n183), .ZN(n181) );
  XNOR2_X1 U836 ( .A(n105), .B(n9), .ZN(SUM[32]) );
  AOI21_X1 U837 ( .B1(n540), .B2(n527), .A(n46), .ZN(n44) );
  AOI21_X1 U838 ( .B1(n540), .B2(n76), .A(n77), .ZN(n71) );
  AOI21_X1 U839 ( .B1(n105), .B2(n92), .A(n93), .ZN(n91) );
  AOI21_X1 U840 ( .B1(n105), .B2(n63), .A(n64), .ZN(n62) );
  AOI21_X1 U841 ( .B1(n105), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U842 ( .B1(n540), .B2(n54), .A(n522), .ZN(n53) );
  AOI21_X1 U843 ( .B1(n540), .B2(n361), .A(n102), .ZN(n100) );
  OAI21_X1 U844 ( .B1(n536), .B2(n148), .A(n139), .ZN(n137) );
  OAI21_X1 U845 ( .B1(n114), .B2(n126), .A(n115), .ZN(n113) );
endmodule


module datapath_DW01_add_11 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n9, n11, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n43, n44, n46, n48, n50, n52, n53, n54, n55, n56, n57, n59,
         n61, n62, n63, n64, n65, n68, n70, n71, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n179, n180,
         n181, n182, n183, n184, n185, n186, n188, n189, n190, n191, n192,
         n193, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n208, n209, n210, n211, n212, n213, n214, n215, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n233, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n246, n247, n248, n249, n252, n253, n254, n255, n256, n257,
         n258, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n275, n276, n277, n278, n279, n280, n283,
         n284, n285, n286, n287, n289, n290, n291, n292, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n353, n360, n361,
         n362, n364, n366, n370, n372, n374, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n565;

  NOR2_X1 U437 ( .A1(n156), .A2(n110), .ZN(n520) );
  CLKBUF_X1 U438 ( .A(B[27]), .Z(n521) );
  NOR2_X1 U439 ( .A1(n521), .A2(A[27]), .ZN(n522) );
  BUF_X1 U440 ( .A(n137), .Z(n554) );
  OR2_X1 U441 ( .A1(A[37]), .A2(B[37]), .ZN(n523) );
  OR2_X1 U442 ( .A1(A[36]), .A2(B[36]), .ZN(n524) );
  OR2_X1 U443 ( .A1(A[38]), .A2(B[38]), .ZN(n525) );
  CLKBUF_X1 U444 ( .A(n180), .Z(n526) );
  XNOR2_X1 U445 ( .A(n140), .B(n527), .ZN(SUM[29]) );
  AND2_X1 U446 ( .A1(n364), .A2(n139), .ZN(n527) );
  BUF_X1 U447 ( .A(n98), .Z(n528) );
  OR2_X1 U448 ( .A1(A[35]), .A2(B[35]), .ZN(n529) );
  AOI21_X1 U449 ( .B1(n158), .B2(n181), .A(n159), .ZN(n530) );
  CLKBUF_X1 U450 ( .A(n218), .Z(n531) );
  XNOR2_X1 U451 ( .A(n116), .B(n532), .ZN(SUM[31]) );
  AND2_X1 U452 ( .A1(n362), .A2(n115), .ZN(n532) );
  OAI21_X1 U453 ( .B1(n237), .B2(n198), .A(n199), .ZN(n533) );
  INV_X1 U454 ( .A(n197), .ZN(n534) );
  NOR2_X1 U455 ( .A1(n557), .A2(n169), .ZN(n535) );
  CLKBUF_X1 U456 ( .A(n169), .Z(n536) );
  CLKBUF_X1 U457 ( .A(n147), .Z(n537) );
  BUF_X1 U458 ( .A(n558), .Z(n541) );
  XNOR2_X1 U459 ( .A(n53), .B(n538), .ZN(SUM[38]) );
  AND2_X1 U460 ( .A1(n525), .A2(n52), .ZN(n538) );
  NOR2_X1 U461 ( .A1(B[29]), .A2(A[29]), .ZN(n539) );
  CLKBUF_X1 U462 ( .A(n209), .Z(n540) );
  XNOR2_X1 U463 ( .A(n100), .B(n542), .ZN(SUM[33]) );
  AND2_X1 U464 ( .A1(n360), .A2(n99), .ZN(n542) );
  XNOR2_X1 U465 ( .A(n44), .B(n543), .ZN(SUM[39]) );
  AND2_X1 U466 ( .A1(n565), .A2(n43), .ZN(n543) );
  XNOR2_X1 U467 ( .A(n62), .B(n544), .ZN(SUM[37]) );
  AND2_X1 U468 ( .A1(n523), .A2(n61), .ZN(n544) );
  XNOR2_X1 U469 ( .A(n84), .B(n545), .ZN(SUM[35]) );
  AND2_X1 U470 ( .A1(n529), .A2(n83), .ZN(n545) );
  CLKBUF_X1 U471 ( .A(n189), .Z(n546) );
  CLKBUF_X1 U472 ( .A(B[25]), .Z(n547) );
  OR2_X2 U473 ( .A1(n236), .A2(n198), .ZN(n548) );
  CLKBUF_X1 U474 ( .A(B[21]), .Z(n549) );
  NOR2_X1 U475 ( .A1(n125), .A2(n114), .ZN(n550) );
  CLKBUF_X1 U476 ( .A(n559), .Z(n551) );
  XNOR2_X1 U477 ( .A(n71), .B(n552), .ZN(SUM[36]) );
  AND2_X1 U478 ( .A1(n524), .A2(n70), .ZN(n552) );
  XNOR2_X1 U479 ( .A(n91), .B(n553), .ZN(SUM[34]) );
  AND2_X1 U480 ( .A1(n88), .A2(n90), .ZN(n553) );
  CLKBUF_X1 U481 ( .A(n181), .Z(n555) );
  OR2_X1 U482 ( .A1(n147), .A2(n138), .ZN(n556) );
  NOR2_X1 U483 ( .A1(A[27]), .A2(B[27]), .ZN(n557) );
  OAI21_X1 U484 ( .B1(n106), .B2(n264), .A(n107), .ZN(n558) );
  OAI21_X1 U485 ( .B1(n106), .B2(n264), .A(n107), .ZN(n105) );
  CLKBUF_X1 U486 ( .A(n539), .Z(n560) );
  NOR2_X1 U487 ( .A1(B[31]), .A2(A[31]), .ZN(n559) );
  OR2_X1 U488 ( .A1(A[25]), .A2(n547), .ZN(n561) );
  INV_X1 U489 ( .A(n48), .ZN(n46) );
  NOR2_X1 U490 ( .A1(A[4]), .A2(B[4]), .ZN(n337) );
  NOR2_X1 U491 ( .A1(A[12]), .A2(B[12]), .ZN(n290) );
  NOR2_X1 U492 ( .A1(A[10]), .A2(B[10]), .ZN(n306) );
  NOR2_X1 U493 ( .A1(A[16]), .A2(B[16]), .ZN(n261) );
  NOR2_X1 U494 ( .A1(A[6]), .A2(B[6]), .ZN(n327) );
  NOR2_X1 U495 ( .A1(A[11]), .A2(B[11]), .ZN(n301) );
  NOR2_X1 U496 ( .A1(A[13]), .A2(B[13]), .ZN(n285) );
  NOR2_X1 U497 ( .A1(A[5]), .A2(B[5]), .ZN(n332) );
  NOR2_X1 U498 ( .A1(A[9]), .A2(B[9]), .ZN(n313) );
  NOR2_X1 U499 ( .A1(A[7]), .A2(B[7]), .ZN(n324) );
  NOR2_X1 U500 ( .A1(A[3]), .A2(B[3]), .ZN(n343) );
  NOR2_X1 U501 ( .A1(A[8]), .A2(B[8]), .ZN(n316) );
  NOR2_X1 U502 ( .A1(A[2]), .A2(B[2]), .ZN(n346) );
  NOR2_X1 U503 ( .A1(A[1]), .A2(B[1]), .ZN(n350) );
  INV_X1 U504 ( .A(n236), .ZN(n230) );
  INV_X1 U505 ( .A(n526), .ZN(n174) );
  INV_X1 U506 ( .A(n548), .ZN(n192) );
  INV_X1 U507 ( .A(n534), .ZN(n193) );
  INV_X1 U508 ( .A(n215), .ZN(n213) );
  INV_X1 U509 ( .A(n214), .ZN(n212) );
  NOR2_X1 U510 ( .A1(n236), .A2(n198), .ZN(n196) );
  INV_X1 U511 ( .A(n156), .ZN(n154) );
  INV_X1 U512 ( .A(n94), .ZN(n92) );
  INV_X1 U513 ( .A(n95), .ZN(n93) );
  OAI21_X1 U514 ( .B1(n318), .B2(n297), .A(n298), .ZN(n292) );
  INV_X1 U515 ( .A(n264), .ZN(n263) );
  INV_X1 U516 ( .A(n154), .ZN(n152) );
  NAND2_X1 U517 ( .A1(n154), .A2(n132), .ZN(n130) );
  NOR2_X1 U518 ( .A1(n78), .A2(n56), .ZN(n54) );
  NAND2_X1 U519 ( .A1(n230), .A2(n531), .ZN(n214) );
  INV_X1 U520 ( .A(n297), .ZN(n295) );
  INV_X1 U521 ( .A(n235), .ZN(n233) );
  INV_X1 U522 ( .A(n556), .ZN(n132) );
  INV_X1 U523 ( .A(n78), .ZN(n76) );
  NAND2_X1 U524 ( .A1(n526), .A2(n167), .ZN(n165) );
  AOI21_X1 U525 ( .B1(n339), .B2(n330), .A(n331), .ZN(n329) );
  NOR2_X1 U526 ( .A1(n78), .A2(n65), .ZN(n63) );
  OAI21_X1 U527 ( .B1(n75), .B2(n65), .A(n70), .ZN(n64) );
  INV_X1 U528 ( .A(n524), .ZN(n65) );
  AND2_X1 U529 ( .A1(n54), .A2(n525), .ZN(n562) );
  AOI21_X1 U530 ( .B1(n319), .B2(n265), .A(n266), .ZN(n264) );
  NOR2_X1 U531 ( .A1(n297), .A2(n267), .ZN(n265) );
  OAI21_X1 U532 ( .B1(n298), .B2(n267), .A(n268), .ZN(n266) );
  NAND2_X1 U533 ( .A1(n283), .A2(n269), .ZN(n267) );
  OAI21_X1 U534 ( .B1(n318), .B2(n279), .A(n280), .ZN(n278) );
  AOI21_X1 U535 ( .B1(n296), .B2(n283), .A(n284), .ZN(n280) );
  NAND2_X1 U536 ( .A1(n295), .A2(n283), .ZN(n279) );
  OAI21_X1 U537 ( .B1(n318), .B2(n309), .A(n310), .ZN(n308) );
  INV_X1 U538 ( .A(n312), .ZN(n310) );
  INV_X1 U539 ( .A(n311), .ZN(n309) );
  INV_X1 U540 ( .A(n319), .ZN(n318) );
  AOI21_X1 U541 ( .B1(n235), .B2(n531), .A(n219), .ZN(n215) );
  NAND2_X1 U542 ( .A1(n154), .A2(n145), .ZN(n143) );
  INV_X1 U543 ( .A(n96), .ZN(n94) );
  INV_X1 U544 ( .A(n554), .ZN(n135) );
  INV_X1 U545 ( .A(n97), .ZN(n95) );
  INV_X1 U546 ( .A(n255), .ZN(n253) );
  NAND2_X1 U547 ( .A1(n254), .A2(n238), .ZN(n236) );
  NAND2_X1 U548 ( .A1(n311), .A2(n299), .ZN(n297) );
  INV_X1 U549 ( .A(n340), .ZN(n339) );
  NOR2_X1 U550 ( .A1(n556), .A2(n123), .ZN(n121) );
  INV_X1 U551 ( .A(n254), .ZN(n252) );
  INV_X1 U552 ( .A(n237), .ZN(n235) );
  INV_X1 U553 ( .A(n77), .ZN(n75) );
  INV_X1 U554 ( .A(n298), .ZN(n296) );
  NAND2_X1 U555 ( .A1(n524), .A2(n523), .ZN(n56) );
  INV_X1 U556 ( .A(n349), .ZN(n348) );
  NOR2_X1 U557 ( .A1(n276), .A2(n271), .ZN(n269) );
  NOR2_X1 U558 ( .A1(n247), .A2(n240), .ZN(n238) );
  NOR2_X1 U559 ( .A1(n261), .A2(n256), .ZN(n254) );
  AOI21_X1 U560 ( .B1(n523), .B2(n68), .A(n59), .ZN(n57) );
  INV_X1 U561 ( .A(n61), .ZN(n59) );
  NOR2_X1 U562 ( .A1(n214), .A2(n540), .ZN(n205) );
  NOR2_X1 U563 ( .A1(n252), .A2(n247), .ZN(n243) );
  OAI21_X1 U564 ( .B1(n253), .B2(n247), .A(n248), .ZN(n244) );
  AOI21_X1 U565 ( .B1(n299), .B2(n312), .A(n300), .ZN(n298) );
  OAI21_X1 U566 ( .B1(n301), .B2(n307), .A(n302), .ZN(n300) );
  AOI21_X1 U567 ( .B1(n341), .B2(n349), .A(n342), .ZN(n340) );
  NOR2_X1 U568 ( .A1(n346), .A2(n343), .ZN(n341) );
  OAI21_X1 U569 ( .B1(n343), .B2(n347), .A(n344), .ZN(n342) );
  OAI21_X1 U570 ( .B1(n332), .B2(n338), .A(n333), .ZN(n331) );
  OAI21_X1 U571 ( .B1(n313), .B2(n317), .A(n314), .ZN(n312) );
  OAI21_X1 U572 ( .B1(n285), .B2(n291), .A(n286), .ZN(n284) );
  OAI21_X1 U573 ( .B1(n350), .B2(n353), .A(n351), .ZN(n349) );
  OAI21_X1 U574 ( .B1(n340), .B2(n320), .A(n321), .ZN(n319) );
  AOI21_X1 U575 ( .B1(n322), .B2(n331), .A(n323), .ZN(n321) );
  NAND2_X1 U576 ( .A1(n330), .A2(n322), .ZN(n320) );
  OAI21_X1 U577 ( .B1(n324), .B2(n328), .A(n325), .ZN(n323) );
  NOR2_X1 U578 ( .A1(n236), .A2(n225), .ZN(n223) );
  OAI21_X1 U579 ( .B1(n233), .B2(n225), .A(n228), .ZN(n224) );
  INV_X1 U580 ( .A(n226), .ZN(n225) );
  INV_X1 U581 ( .A(n104), .ZN(n102) );
  NOR2_X1 U582 ( .A1(n94), .A2(n87), .ZN(n85) );
  OAI21_X1 U583 ( .B1(n95), .B2(n87), .A(n90), .ZN(n86) );
  INV_X1 U584 ( .A(n88), .ZN(n87) );
  INV_X1 U585 ( .A(n262), .ZN(n260) );
  AOI21_X1 U586 ( .B1(n238), .B2(n255), .A(n239), .ZN(n237) );
  NOR2_X1 U587 ( .A1(n327), .A2(n324), .ZN(n322) );
  NOR2_X1 U588 ( .A1(n337), .A2(n332), .ZN(n330) );
  NOR2_X1 U589 ( .A1(n306), .A2(n301), .ZN(n299) );
  OAI21_X1 U590 ( .B1(n135), .B2(n123), .A(n126), .ZN(n122) );
  INV_X1 U591 ( .A(n148), .ZN(n146) );
  NOR2_X1 U592 ( .A1(n316), .A2(n313), .ZN(n311) );
  NOR2_X1 U593 ( .A1(n290), .A2(n285), .ZN(n283) );
  AOI21_X1 U594 ( .B1(n55), .B2(n525), .A(n50), .ZN(n48) );
  INV_X1 U595 ( .A(n52), .ZN(n50) );
  AOI21_X1 U596 ( .B1(n269), .B2(n284), .A(n270), .ZN(n268) );
  AOI21_X1 U597 ( .B1(n292), .B2(n381), .A(n289), .ZN(n287) );
  INV_X1 U598 ( .A(n291), .ZN(n289) );
  AOI21_X1 U599 ( .B1(n308), .B2(n383), .A(n305), .ZN(n303) );
  INV_X1 U600 ( .A(n307), .ZN(n305) );
  AOI21_X1 U601 ( .B1(n278), .B2(n379), .A(n275), .ZN(n273) );
  INV_X1 U602 ( .A(n277), .ZN(n275) );
  OAI21_X1 U603 ( .B1(n318), .B2(n316), .A(n317), .ZN(n315) );
  INV_X1 U604 ( .A(n227), .ZN(n226) );
  INV_X1 U605 ( .A(n546), .ZN(n188) );
  AOI21_X1 U606 ( .B1(n555), .B2(n167), .A(n168), .ZN(n166) );
  INV_X1 U607 ( .A(n170), .ZN(n168) );
  INV_X1 U608 ( .A(n271), .ZN(n378) );
  INV_X1 U609 ( .A(n522), .ZN(n366) );
  INV_X1 U610 ( .A(n70), .ZN(n68) );
  INV_X1 U611 ( .A(n124), .ZN(n123) );
  INV_X1 U612 ( .A(n89), .ZN(n88) );
  INV_X1 U613 ( .A(n560), .ZN(n364) );
  INV_X1 U614 ( .A(n327), .ZN(n387) );
  INV_X1 U615 ( .A(n346), .ZN(n391) );
  INV_X1 U616 ( .A(n316), .ZN(n385) );
  INV_X1 U617 ( .A(n285), .ZN(n380) );
  INV_X1 U618 ( .A(n301), .ZN(n382) );
  INV_X1 U619 ( .A(n313), .ZN(n384) );
  INV_X1 U620 ( .A(n290), .ZN(n381) );
  INV_X1 U621 ( .A(n337), .ZN(n389) );
  INV_X1 U622 ( .A(n306), .ZN(n383) );
  NAND2_X1 U623 ( .A1(n386), .A2(n325), .ZN(n34) );
  INV_X1 U624 ( .A(n324), .ZN(n386) );
  INV_X1 U625 ( .A(n261), .ZN(n377) );
  NAND2_X1 U626 ( .A1(n388), .A2(n333), .ZN(n36) );
  INV_X1 U627 ( .A(n332), .ZN(n388) );
  NAND2_X1 U628 ( .A1(n390), .A2(n344), .ZN(n38) );
  INV_X1 U629 ( .A(n343), .ZN(n390) );
  INV_X1 U630 ( .A(n103), .ZN(n361) );
  INV_X1 U631 ( .A(n350), .ZN(n392) );
  INV_X1 U632 ( .A(n338), .ZN(n336) );
  INV_X1 U633 ( .A(n551), .ZN(n362) );
  INV_X1 U634 ( .A(n220), .ZN(n372) );
  INV_X1 U635 ( .A(n202), .ZN(n370) );
  OR2_X1 U636 ( .A1(A[0]), .A2(B[0]), .ZN(n563) );
  NOR2_X1 U637 ( .A1(A[32]), .A2(B[32]), .ZN(n103) );
  NOR2_X1 U638 ( .A1(A[34]), .A2(B[34]), .ZN(n89) );
  NOR2_X1 U639 ( .A1(B[21]), .A2(A[21]), .ZN(n220) );
  NOR2_X1 U640 ( .A1(A[23]), .A2(B[23]), .ZN(n202) );
  NOR2_X1 U641 ( .A1(B[31]), .A2(A[31]), .ZN(n114) );
  NOR2_X1 U642 ( .A1(A[17]), .A2(B[17]), .ZN(n256) );
  NOR2_X1 U643 ( .A1(A[19]), .A2(B[19]), .ZN(n240) );
  NOR2_X1 U644 ( .A1(A[30]), .A2(B[30]), .ZN(n125) );
  NOR2_X1 U645 ( .A1(A[18]), .A2(B[18]), .ZN(n247) );
  NOR2_X1 U646 ( .A1(B[25]), .A2(A[25]), .ZN(n182) );
  NOR2_X1 U647 ( .A1(B[29]), .A2(A[29]), .ZN(n138) );
  NAND2_X1 U648 ( .A1(A[30]), .A2(B[30]), .ZN(n126) );
  NAND2_X1 U649 ( .A1(A[32]), .A2(B[32]), .ZN(n104) );
  NAND2_X1 U650 ( .A1(A[34]), .A2(B[34]), .ZN(n90) );
  NAND2_X1 U651 ( .A1(n124), .A2(n126), .ZN(n11) );
  NAND2_X1 U652 ( .A1(n372), .A2(n221), .ZN(n20) );
  NAND2_X1 U653 ( .A1(n376), .A2(n257), .ZN(n24) );
  NOR2_X1 U654 ( .A1(A[26]), .A2(B[26]), .ZN(n169) );
  NAND2_X1 U655 ( .A1(n226), .A2(n228), .ZN(n21) );
  NOR2_X1 U656 ( .A1(B[22]), .A2(A[22]), .ZN(n209) );
  NOR2_X1 U657 ( .A1(A[35]), .A2(B[35]), .ZN(n82) );
  NOR2_X1 U658 ( .A1(A[33]), .A2(B[33]), .ZN(n98) );
  NAND2_X1 U659 ( .A1(A[2]), .A2(B[2]), .ZN(n347) );
  NAND2_X1 U660 ( .A1(n377), .A2(n262), .ZN(n25) );
  NAND2_X1 U661 ( .A1(A[6]), .A2(B[6]), .ZN(n328) );
  XOR2_X1 U662 ( .A(n329), .B(n35), .Z(SUM[6]) );
  NAND2_X1 U663 ( .A1(n387), .A2(n328), .ZN(n35) );
  XOR2_X1 U664 ( .A(n204), .B(n18), .Z(SUM[23]) );
  NAND2_X1 U665 ( .A1(n370), .A2(n203), .ZN(n18) );
  XOR2_X1 U666 ( .A(n162), .B(n14), .Z(SUM[27]) );
  NAND2_X1 U667 ( .A1(n366), .A2(n161), .ZN(n14) );
  XOR2_X1 U668 ( .A(n249), .B(n23), .Z(SUM[18]) );
  NAND2_X1 U669 ( .A1(n246), .A2(n248), .ZN(n23) );
  XOR2_X1 U670 ( .A(n242), .B(n22), .Z(SUM[19]) );
  NAND2_X1 U671 ( .A1(n374), .A2(n241), .ZN(n22) );
  XOR2_X1 U672 ( .A(n191), .B(n17), .Z(SUM[24]) );
  NAND2_X1 U673 ( .A1(n188), .A2(n190), .ZN(n17) );
  XOR2_X1 U674 ( .A(n211), .B(n19), .Z(SUM[22]) );
  NAND2_X1 U675 ( .A1(n208), .A2(n210), .ZN(n19) );
  NAND2_X1 U676 ( .A1(A[8]), .A2(B[8]), .ZN(n317) );
  NAND2_X1 U677 ( .A1(A[12]), .A2(B[12]), .ZN(n291) );
  NAND2_X1 U678 ( .A1(A[10]), .A2(B[10]), .ZN(n307) );
  NAND2_X1 U679 ( .A1(A[4]), .A2(B[4]), .ZN(n338) );
  XOR2_X1 U680 ( .A(n184), .B(n16), .Z(SUM[25]) );
  NAND2_X1 U681 ( .A1(n561), .A2(n183), .ZN(n16) );
  XOR2_X1 U682 ( .A(n171), .B(n15), .Z(SUM[26]) );
  NAND2_X1 U683 ( .A1(n167), .A2(n170), .ZN(n15) );
  NAND2_X1 U684 ( .A1(n361), .A2(n104), .ZN(n9) );
  XNOR2_X1 U685 ( .A(n292), .B(n29), .ZN(SUM[12]) );
  NAND2_X1 U686 ( .A1(n381), .A2(n291), .ZN(n29) );
  XNOR2_X1 U687 ( .A(n308), .B(n31), .ZN(SUM[10]) );
  NAND2_X1 U688 ( .A1(n383), .A2(n307), .ZN(n31) );
  XNOR2_X1 U689 ( .A(n315), .B(n32), .ZN(SUM[9]) );
  NAND2_X1 U690 ( .A1(n384), .A2(n314), .ZN(n32) );
  XOR2_X1 U691 ( .A(n40), .B(n353), .Z(SUM[1]) );
  NAND2_X1 U692 ( .A1(n392), .A2(n351), .ZN(n40) );
  XNOR2_X1 U693 ( .A(n345), .B(n38), .ZN(SUM[3]) );
  OAI21_X1 U694 ( .B1(n348), .B2(n346), .A(n347), .ZN(n345) );
  XNOR2_X1 U695 ( .A(n339), .B(n37), .ZN(SUM[4]) );
  NAND2_X1 U696 ( .A1(n389), .A2(n338), .ZN(n37) );
  XOR2_X1 U697 ( .A(n318), .B(n33), .Z(SUM[8]) );
  NAND2_X1 U698 ( .A1(n385), .A2(n317), .ZN(n33) );
  XOR2_X1 U699 ( .A(n334), .B(n36), .Z(SUM[5]) );
  AOI21_X1 U700 ( .B1(n339), .B2(n389), .A(n336), .ZN(n334) );
  XNOR2_X1 U701 ( .A(n326), .B(n34), .ZN(SUM[7]) );
  OAI21_X1 U702 ( .B1(n329), .B2(n327), .A(n328), .ZN(n326) );
  AND2_X1 U703 ( .A1(n563), .A2(n353), .ZN(SUM[0]) );
  XOR2_X1 U704 ( .A(n348), .B(n39), .Z(SUM[2]) );
  NAND2_X1 U705 ( .A1(n391), .A2(n347), .ZN(n39) );
  NAND2_X1 U706 ( .A1(A[5]), .A2(B[5]), .ZN(n333) );
  NAND2_X1 U707 ( .A1(A[7]), .A2(B[7]), .ZN(n325) );
  NAND2_X1 U708 ( .A1(A[0]), .A2(B[0]), .ZN(n353) );
  NAND2_X1 U709 ( .A1(A[16]), .A2(B[16]), .ZN(n262) );
  NAND2_X1 U710 ( .A1(B[26]), .A2(A[26]), .ZN(n170) );
  XNOR2_X1 U711 ( .A(n278), .B(n27), .ZN(SUM[14]) );
  NAND2_X1 U712 ( .A1(n379), .A2(n277), .ZN(n27) );
  NAND2_X1 U713 ( .A1(A[38]), .A2(B[38]), .ZN(n52) );
  NAND2_X1 U714 ( .A1(A[11]), .A2(B[11]), .ZN(n302) );
  NAND2_X1 U715 ( .A1(A[13]), .A2(B[13]), .ZN(n286) );
  NAND2_X1 U716 ( .A1(A[9]), .A2(B[9]), .ZN(n314) );
  NAND2_X1 U717 ( .A1(A[1]), .A2(B[1]), .ZN(n351) );
  NAND2_X1 U718 ( .A1(A[3]), .A2(B[3]), .ZN(n344) );
  NAND2_X1 U719 ( .A1(A[18]), .A2(B[18]), .ZN(n248) );
  NAND2_X1 U720 ( .A1(A[14]), .A2(B[14]), .ZN(n277) );
  NAND2_X1 U721 ( .A1(A[37]), .A2(B[37]), .ZN(n61) );
  NAND2_X1 U722 ( .A1(A[36]), .A2(B[36]), .ZN(n70) );
  NAND2_X1 U723 ( .A1(A[39]), .A2(B[39]), .ZN(n43) );
  NAND2_X1 U724 ( .A1(A[17]), .A2(B[17]), .ZN(n257) );
  NAND2_X1 U725 ( .A1(A[19]), .A2(B[19]), .ZN(n241) );
  NAND2_X1 U726 ( .A1(A[35]), .A2(B[35]), .ZN(n83) );
  XOR2_X1 U727 ( .A(n149), .B(n13), .Z(SUM[28]) );
  XOR2_X1 U728 ( .A(n273), .B(n26), .Z(SUM[15]) );
  NAND2_X1 U729 ( .A1(n378), .A2(n272), .ZN(n26) );
  XOR2_X1 U730 ( .A(n287), .B(n28), .Z(SUM[13]) );
  NAND2_X1 U731 ( .A1(n380), .A2(n286), .ZN(n28) );
  XOR2_X1 U732 ( .A(n303), .B(n30), .Z(SUM[11]) );
  NAND2_X1 U733 ( .A1(n382), .A2(n302), .ZN(n30) );
  OR2_X1 U734 ( .A1(A[39]), .A2(B[39]), .ZN(n565) );
  NAND2_X1 U735 ( .A1(A[23]), .A2(B[23]), .ZN(n203) );
  NAND2_X1 U736 ( .A1(A[15]), .A2(B[15]), .ZN(n272) );
  NOR2_X1 U737 ( .A1(A[15]), .A2(B[15]), .ZN(n271) );
  INV_X1 U738 ( .A(n247), .ZN(n246) );
  INV_X1 U739 ( .A(n276), .ZN(n379) );
  NOR2_X1 U740 ( .A1(A[14]), .A2(B[14]), .ZN(n276) );
  NAND2_X1 U741 ( .A1(A[20]), .A2(B[20]), .ZN(n228) );
  NOR2_X1 U742 ( .A1(A[20]), .A2(B[20]), .ZN(n227) );
  NOR2_X1 U743 ( .A1(n209), .A2(n202), .ZN(n200) );
  INV_X1 U744 ( .A(n540), .ZN(n208) );
  INV_X1 U745 ( .A(n528), .ZN(n360) );
  NOR2_X1 U746 ( .A1(n103), .A2(n528), .ZN(n96) );
  OAI21_X1 U747 ( .B1(n98), .B2(n104), .A(n99), .ZN(n97) );
  NAND2_X1 U748 ( .A1(B[27]), .A2(A[27]), .ZN(n161) );
  NOR2_X1 U749 ( .A1(B[27]), .A2(A[27]), .ZN(n160) );
  INV_X1 U750 ( .A(n125), .ZN(n124) );
  XOR2_X1 U751 ( .A(n229), .B(n21), .Z(SUM[20]) );
  OAI21_X1 U752 ( .B1(n256), .B2(n262), .A(n257), .ZN(n255) );
  INV_X1 U753 ( .A(n256), .ZN(n376) );
  NAND2_X1 U754 ( .A1(A[24]), .A2(B[24]), .ZN(n190) );
  NOR2_X1 U755 ( .A1(B[24]), .A2(A[24]), .ZN(n189) );
  XOR2_X1 U756 ( .A(n222), .B(n20), .Z(SUM[21]) );
  OAI21_X1 U757 ( .B1(n240), .B2(n248), .A(n241), .ZN(n239) );
  INV_X1 U758 ( .A(n240), .ZN(n374) );
  XOR2_X1 U759 ( .A(n127), .B(n11), .Z(SUM[30]) );
  INV_X1 U760 ( .A(n537), .ZN(n145) );
  NAND2_X1 U761 ( .A1(n145), .A2(n148), .ZN(n13) );
  OAI21_X1 U762 ( .B1(n138), .B2(n148), .A(n139), .ZN(n137) );
  OAI21_X1 U763 ( .B1(n237), .B2(n198), .A(n199), .ZN(n197) );
  NAND2_X1 U764 ( .A1(A[22]), .A2(B[22]), .ZN(n210) );
  XNOR2_X1 U765 ( .A(n263), .B(n25), .ZN(SUM[16]) );
  XOR2_X1 U766 ( .A(n258), .B(n24), .Z(SUM[17]) );
  AOI21_X1 U767 ( .B1(n263), .B2(n141), .A(n142), .ZN(n140) );
  AOI21_X1 U768 ( .B1(n263), .B2(n377), .A(n260), .ZN(n258) );
  AOI21_X1 U769 ( .B1(n263), .B2(n254), .A(n255), .ZN(n249) );
  AOI21_X1 U770 ( .B1(n263), .B2(n230), .A(n235), .ZN(n229) );
  AOI21_X1 U771 ( .B1(n263), .B2(n212), .A(n213), .ZN(n211) );
  AOI21_X1 U772 ( .B1(n263), .B2(n243), .A(n244), .ZN(n242) );
  AOI21_X1 U773 ( .B1(n263), .B2(n223), .A(n224), .ZN(n222) );
  AOI21_X1 U774 ( .B1(n263), .B2(n205), .A(n206), .ZN(n204) );
  AOI21_X1 U775 ( .B1(n263), .B2(n192), .A(n193), .ZN(n191) );
  AOI21_X1 U776 ( .B1(n263), .B2(n172), .A(n173), .ZN(n171) );
  AOI21_X1 U777 ( .B1(n263), .B2(n163), .A(n164), .ZN(n162) );
  OAI21_X1 U778 ( .B1(n271), .B2(n277), .A(n272), .ZN(n270) );
  INV_X1 U779 ( .A(n79), .ZN(n77) );
  OAI21_X1 U780 ( .B1(n215), .B2(n540), .A(n210), .ZN(n206) );
  NAND2_X1 U781 ( .A1(n200), .A2(n218), .ZN(n198) );
  NOR2_X1 U782 ( .A1(n227), .A2(n220), .ZN(n218) );
  AOI21_X1 U783 ( .B1(n263), .B2(n117), .A(n118), .ZN(n116) );
  NOR2_X1 U784 ( .A1(B[28]), .A2(A[28]), .ZN(n147) );
  NAND2_X1 U785 ( .A1(B[28]), .A2(A[28]), .ZN(n148) );
  INV_X1 U786 ( .A(n197), .ZN(n195) );
  AOI21_X1 U787 ( .B1(n263), .B2(n185), .A(n186), .ZN(n184) );
  OAI21_X1 U788 ( .B1(n220), .B2(n228), .A(n221), .ZN(n219) );
  NAND2_X1 U789 ( .A1(A[21]), .A2(n549), .ZN(n221) );
  AOI21_X1 U790 ( .B1(n263), .B2(n150), .A(n151), .ZN(n149) );
  NAND2_X1 U791 ( .A1(B[25]), .A2(A[25]), .ZN(n183) );
  AOI21_X1 U792 ( .B1(n137), .B2(n550), .A(n113), .ZN(n111) );
  AOI21_X1 U793 ( .B1(n263), .B2(n128), .A(n129), .ZN(n127) );
  NAND2_X1 U794 ( .A1(B[31]), .A2(A[31]), .ZN(n115) );
  NOR2_X1 U795 ( .A1(n169), .A2(n557), .ZN(n158) );
  INV_X1 U796 ( .A(n536), .ZN(n167) );
  NOR2_X1 U797 ( .A1(n548), .A2(n143), .ZN(n141) );
  NOR2_X1 U798 ( .A1(n548), .A2(n546), .ZN(n185) );
  NOR2_X1 U799 ( .A1(n548), .A2(n174), .ZN(n172) );
  NOR2_X1 U800 ( .A1(n548), .A2(n165), .ZN(n163) );
  NOR2_X1 U801 ( .A1(n548), .A2(n152), .ZN(n150) );
  NOR2_X1 U802 ( .A1(n548), .A2(n130), .ZN(n128) );
  AOI21_X1 U803 ( .B1(n219), .B2(n200), .A(n201), .ZN(n199) );
  AOI21_X1 U804 ( .B1(n80), .B2(n97), .A(n81), .ZN(n79) );
  NAND2_X1 U805 ( .A1(n96), .A2(n80), .ZN(n78) );
  OAI21_X1 U806 ( .B1(n195), .B2(n143), .A(n144), .ZN(n142) );
  OAI21_X1 U807 ( .B1(n195), .B2(n546), .A(n190), .ZN(n186) );
  OAI21_X1 U808 ( .B1(n534), .B2(n174), .A(n179), .ZN(n173) );
  OAI21_X1 U809 ( .B1(n195), .B2(n165), .A(n166), .ZN(n164) );
  OAI21_X1 U810 ( .B1(n534), .B2(n152), .A(n530), .ZN(n151) );
  OAI21_X1 U811 ( .B1(n195), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U812 ( .B1(n202), .B2(n210), .A(n203), .ZN(n201) );
  NOR2_X1 U813 ( .A1(n89), .A2(n82), .ZN(n80) );
  OAI21_X1 U814 ( .B1(n82), .B2(n90), .A(n83), .ZN(n81) );
  NOR2_X1 U815 ( .A1(n548), .A2(n119), .ZN(n117) );
  NOR2_X1 U816 ( .A1(n114), .A2(n125), .ZN(n112) );
  AOI21_X1 U817 ( .B1(n158), .B2(n181), .A(n159), .ZN(n157) );
  INV_X1 U818 ( .A(n555), .ZN(n179) );
  INV_X1 U819 ( .A(n530), .ZN(n155) );
  AOI21_X1 U820 ( .B1(n155), .B2(n132), .A(n554), .ZN(n131) );
  AOI21_X1 U821 ( .B1(n155), .B2(n145), .A(n146), .ZN(n144) );
  NOR2_X1 U822 ( .A1(n156), .A2(n110), .ZN(n108) );
  NAND2_X1 U823 ( .A1(n180), .A2(n535), .ZN(n156) );
  OAI21_X1 U824 ( .B1(n79), .B2(n56), .A(n57), .ZN(n55) );
  NAND2_X1 U825 ( .A1(A[33]), .A2(B[33]), .ZN(n99) );
  AOI21_X1 U826 ( .B1(n121), .B2(n155), .A(n122), .ZN(n120) );
  NAND2_X1 U827 ( .A1(n121), .A2(n154), .ZN(n119) );
  NAND2_X1 U828 ( .A1(n136), .A2(n112), .ZN(n110) );
  OAI21_X1 U829 ( .B1(n195), .B2(n119), .A(n120), .ZN(n118) );
  OAI21_X1 U830 ( .B1(n157), .B2(n110), .A(n111), .ZN(n109) );
  OAI21_X1 U831 ( .B1(n160), .B2(n170), .A(n161), .ZN(n159) );
  NOR2_X1 U832 ( .A1(n182), .A2(n189), .ZN(n180) );
  OAI21_X1 U833 ( .B1(n182), .B2(n190), .A(n183), .ZN(n181) );
  XNOR2_X1 U834 ( .A(n541), .B(n9), .ZN(SUM[32]) );
  AOI21_X1 U835 ( .B1(n105), .B2(n54), .A(n55), .ZN(n53) );
  AOI21_X1 U836 ( .B1(n105), .B2(n76), .A(n77), .ZN(n71) );
  AOI21_X1 U837 ( .B1(n105), .B2(n92), .A(n93), .ZN(n91) );
  AOI21_X1 U838 ( .B1(n105), .B2(n361), .A(n102), .ZN(n100) );
  AOI21_X1 U839 ( .B1(n558), .B2(n562), .A(n46), .ZN(n44) );
  AOI21_X1 U840 ( .B1(n558), .B2(n63), .A(n64), .ZN(n62) );
  AOI21_X1 U841 ( .B1(n558), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U842 ( .B1(n533), .B2(n108), .A(n109), .ZN(n107) );
  NAND2_X1 U843 ( .A1(n520), .A2(n196), .ZN(n106) );
  NOR2_X1 U844 ( .A1(n147), .A2(n539), .ZN(n136) );
  NAND2_X1 U845 ( .A1(B[29]), .A2(A[29]), .ZN(n139) );
  OAI21_X1 U846 ( .B1(n559), .B2(n126), .A(n115), .ZN(n113) );
endmodule


module datapath_DW01_add_12 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n9, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n43, n44, n46, n48, n50, n52, n53, n54, n55, n56, n57, n59,
         n61, n62, n63, n64, n67, n68, n69, n70, n71, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n93, n94,
         n95, n96, n97, n98, n99, n100, n102, n103, n104, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n125, n126, n127, n128, n129, n130, n131,
         n132, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n176, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n208, n209, n210, n211, n212, n213, n214, n215, n218,
         n219, n220, n221, n222, n223, n224, n226, n227, n228, n229, n230,
         n233, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n246, n247, n248, n249, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n275, n276, n277, n278, n279, n280, n283,
         n284, n285, n286, n287, n289, n290, n291, n292, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n353, n358, n360,
         n361, n362, n364, n365, n366, n368, n370, n372, n374, n376, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n520, n521, n522, n523, n524, n525, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560;

  INV_X1 U437 ( .A(n197), .ZN(n520) );
  CLKBUF_X1 U438 ( .A(n147), .Z(n521) );
  CLKBUF_X1 U439 ( .A(n218), .Z(n522) );
  NOR2_X1 U440 ( .A1(n247), .A2(n240), .ZN(n238) );
  NOR2_X1 U441 ( .A1(A[17]), .A2(B[17]), .ZN(n256) );
  NOR2_X1 U442 ( .A1(A[13]), .A2(B[13]), .ZN(n285) );
  NOR2_X1 U443 ( .A1(A[11]), .A2(B[11]), .ZN(n301) );
  OR2_X1 U444 ( .A1(A[37]), .A2(B[37]), .ZN(n523) );
  OR2_X1 U445 ( .A1(A[38]), .A2(B[38]), .ZN(n524) );
  OR2_X1 U446 ( .A1(A[30]), .A2(B[30]), .ZN(n525) );
  AND2_X1 U447 ( .A1(n528), .A2(n353), .ZN(SUM[0]) );
  NOR2_X1 U448 ( .A1(A[16]), .A2(B[16]), .ZN(n261) );
  NOR2_X1 U449 ( .A1(A[18]), .A2(B[18]), .ZN(n247) );
  AND2_X1 U450 ( .A1(n54), .A2(n524), .ZN(n527) );
  OR2_X1 U451 ( .A1(A[0]), .A2(B[0]), .ZN(n528) );
  XNOR2_X1 U452 ( .A(n127), .B(n529), .ZN(SUM[30]) );
  AND2_X1 U453 ( .A1(n525), .A2(n126), .ZN(n529) );
  XNOR2_X1 U454 ( .A(n140), .B(n530), .ZN(SUM[29]) );
  AND2_X1 U455 ( .A1(n364), .A2(n139), .ZN(n530) );
  NOR2_X1 U456 ( .A1(A[33]), .A2(B[33]), .ZN(n531) );
  NOR2_X1 U457 ( .A1(A[35]), .A2(B[35]), .ZN(n532) );
  XNOR2_X1 U458 ( .A(n116), .B(n533), .ZN(SUM[31]) );
  AND2_X1 U459 ( .A1(n362), .A2(n115), .ZN(n533) );
  CLKBUF_X1 U460 ( .A(n169), .Z(n534) );
  CLKBUF_X1 U461 ( .A(n227), .Z(n535) );
  CLKBUF_X1 U462 ( .A(n559), .Z(n536) );
  BUF_X1 U463 ( .A(n541), .Z(n1) );
  OR2_X1 U464 ( .A1(n189), .A2(n182), .ZN(n537) );
  CLKBUF_X1 U465 ( .A(n181), .Z(n538) );
  NOR2_X1 U466 ( .A1(n160), .A2(n169), .ZN(n539) );
  OAI21_X1 U467 ( .B1(n106), .B2(n264), .A(n107), .ZN(n540) );
  OAI21_X1 U468 ( .B1(n106), .B2(n264), .A(n107), .ZN(n541) );
  CLKBUF_X1 U469 ( .A(n209), .Z(n542) );
  NOR2_X1 U470 ( .A1(B[25]), .A2(A[25]), .ZN(n543) );
  NOR2_X1 U471 ( .A1(n125), .A2(n547), .ZN(n544) );
  CLKBUF_X1 U472 ( .A(n137), .Z(n545) );
  NOR2_X1 U473 ( .A1(A[27]), .A2(B[27]), .ZN(n546) );
  NOR2_X1 U474 ( .A1(A[31]), .A2(B[31]), .ZN(n547) );
  XNOR2_X1 U475 ( .A(n44), .B(n548), .ZN(SUM[39]) );
  AND2_X1 U476 ( .A1(n560), .A2(n43), .ZN(n548) );
  XNOR2_X1 U477 ( .A(n62), .B(n549), .ZN(SUM[37]) );
  AND2_X1 U478 ( .A1(n523), .A2(n61), .ZN(n549) );
  XNOR2_X1 U479 ( .A(n71), .B(n550), .ZN(SUM[36]) );
  AND2_X1 U480 ( .A1(n67), .A2(n70), .ZN(n550) );
  XNOR2_X1 U481 ( .A(n84), .B(n551), .ZN(SUM[35]) );
  AND2_X1 U482 ( .A1(n358), .A2(n83), .ZN(n551) );
  XNOR2_X1 U483 ( .A(n91), .B(n552), .ZN(SUM[34]) );
  AND2_X1 U484 ( .A1(n88), .A2(n90), .ZN(n552) );
  XNOR2_X1 U485 ( .A(n100), .B(n553), .ZN(SUM[33]) );
  AND2_X1 U486 ( .A1(n360), .A2(n99), .ZN(n553) );
  XNOR2_X1 U487 ( .A(n53), .B(n554), .ZN(SUM[38]) );
  AND2_X1 U488 ( .A1(n524), .A2(n52), .ZN(n554) );
  CLKBUF_X1 U489 ( .A(n543), .Z(n555) );
  CLKBUF_X1 U490 ( .A(n160), .Z(n556) );
  CLKBUF_X1 U491 ( .A(n156), .Z(n557) );
  NOR2_X1 U492 ( .A1(B[25]), .A2(A[25]), .ZN(n182) );
  NOR2_X1 U493 ( .A1(B[27]), .A2(A[27]), .ZN(n160) );
  OR2_X1 U494 ( .A1(n147), .A2(n138), .ZN(n558) );
  NOR2_X1 U495 ( .A1(B[29]), .A2(A[29]), .ZN(n559) );
  AOI21_X1 U496 ( .B1(n299), .B2(n312), .A(n300), .ZN(n298) );
  NOR2_X1 U497 ( .A1(n306), .A2(n301), .ZN(n299) );
  OAI21_X1 U498 ( .B1(n285), .B2(n291), .A(n286), .ZN(n284) );
  NOR2_X1 U499 ( .A1(n261), .A2(n256), .ZN(n254) );
  NOR2_X1 U500 ( .A1(n290), .A2(n285), .ZN(n283) );
  NOR2_X1 U501 ( .A1(A[10]), .A2(B[10]), .ZN(n306) );
  NOR2_X1 U502 ( .A1(A[12]), .A2(B[12]), .ZN(n290) );
  NOR2_X1 U503 ( .A1(A[4]), .A2(B[4]), .ZN(n337) );
  NOR2_X1 U504 ( .A1(A[14]), .A2(B[14]), .ZN(n276) );
  NOR2_X1 U505 ( .A1(A[6]), .A2(B[6]), .ZN(n327) );
  NOR2_X1 U506 ( .A1(A[7]), .A2(B[7]), .ZN(n324) );
  NOR2_X1 U507 ( .A1(A[35]), .A2(B[35]), .ZN(n82) );
  NOR2_X1 U508 ( .A1(A[9]), .A2(B[9]), .ZN(n313) );
  NOR2_X1 U509 ( .A1(A[5]), .A2(B[5]), .ZN(n332) );
  NOR2_X1 U510 ( .A1(A[3]), .A2(B[3]), .ZN(n343) );
  NOR2_X1 U511 ( .A1(A[8]), .A2(B[8]), .ZN(n316) );
  NOR2_X1 U512 ( .A1(A[2]), .A2(B[2]), .ZN(n346) );
  NOR2_X1 U513 ( .A1(A[1]), .A2(B[1]), .ZN(n350) );
  INV_X1 U514 ( .A(n236), .ZN(n230) );
  INV_X1 U515 ( .A(n215), .ZN(n213) );
  INV_X1 U516 ( .A(n214), .ZN(n212) );
  INV_X1 U517 ( .A(n557), .ZN(n154) );
  INV_X1 U518 ( .A(n95), .ZN(n93) );
  INV_X1 U519 ( .A(n194), .ZN(n192) );
  OAI21_X1 U520 ( .B1(n318), .B2(n297), .A(n298), .ZN(n292) );
  INV_X1 U521 ( .A(n264), .ZN(n263) );
  NAND2_X1 U522 ( .A1(n154), .A2(n132), .ZN(n130) );
  NOR2_X1 U523 ( .A1(n78), .A2(n56), .ZN(n54) );
  AOI21_X1 U524 ( .B1(n155), .B2(n132), .A(n545), .ZN(n131) );
  NAND2_X1 U525 ( .A1(n230), .A2(n522), .ZN(n214) );
  INV_X1 U526 ( .A(n558), .ZN(n132) );
  INV_X1 U527 ( .A(n297), .ZN(n295) );
  INV_X1 U528 ( .A(n235), .ZN(n233) );
  INV_X1 U529 ( .A(n78), .ZN(n76) );
  NAND2_X1 U530 ( .A1(n176), .A2(n167), .ZN(n165) );
  AOI21_X1 U531 ( .B1(n235), .B2(n522), .A(n219), .ZN(n215) );
  AOI21_X1 U532 ( .B1(n339), .B2(n330), .A(n331), .ZN(n329) );
  OAI21_X1 U533 ( .B1(n75), .B2(n69), .A(n70), .ZN(n64) );
  NOR2_X1 U534 ( .A1(n78), .A2(n69), .ZN(n63) );
  INV_X1 U535 ( .A(n48), .ZN(n46) );
  AOI21_X1 U536 ( .B1(n319), .B2(n265), .A(n266), .ZN(n264) );
  OAI21_X1 U537 ( .B1(n298), .B2(n267), .A(n268), .ZN(n266) );
  NOR2_X1 U538 ( .A1(n297), .A2(n267), .ZN(n265) );
  AOI21_X1 U539 ( .B1(n269), .B2(n284), .A(n270), .ZN(n268) );
  OAI21_X1 U540 ( .B1(n318), .B2(n279), .A(n280), .ZN(n278) );
  AOI21_X1 U541 ( .B1(n296), .B2(n283), .A(n284), .ZN(n280) );
  NAND2_X1 U542 ( .A1(n295), .A2(n283), .ZN(n279) );
  OAI21_X1 U543 ( .B1(n318), .B2(n309), .A(n310), .ZN(n308) );
  INV_X1 U544 ( .A(n312), .ZN(n310) );
  INV_X1 U545 ( .A(n311), .ZN(n309) );
  NOR2_X1 U546 ( .A1(n558), .A2(n123), .ZN(n121) );
  INV_X1 U547 ( .A(n319), .ZN(n318) );
  NAND2_X1 U548 ( .A1(n154), .A2(n365), .ZN(n143) );
  NAND2_X1 U549 ( .A1(n121), .A2(n154), .ZN(n119) );
  INV_X1 U550 ( .A(n97), .ZN(n95) );
  INV_X1 U551 ( .A(n157), .ZN(n155) );
  NAND2_X1 U552 ( .A1(n283), .A2(n269), .ZN(n267) );
  NAND2_X1 U553 ( .A1(n311), .A2(n299), .ZN(n297) );
  INV_X1 U554 ( .A(n340), .ZN(n339) );
  INV_X1 U555 ( .A(n255), .ZN(n253) );
  INV_X1 U556 ( .A(n254), .ZN(n252) );
  INV_X1 U557 ( .A(n96), .ZN(n94) );
  NAND2_X1 U558 ( .A1(n254), .A2(n238), .ZN(n236) );
  INV_X1 U559 ( .A(n298), .ZN(n296) );
  INV_X1 U560 ( .A(n349), .ZN(n348) );
  INV_X1 U561 ( .A(n538), .ZN(n179) );
  INV_X1 U562 ( .A(n537), .ZN(n176) );
  INV_X1 U563 ( .A(n237), .ZN(n235) );
  NAND2_X1 U564 ( .A1(n67), .A2(n523), .ZN(n56) );
  INV_X1 U565 ( .A(n77), .ZN(n75) );
  NOR2_X1 U566 ( .A1(n276), .A2(n271), .ZN(n269) );
  NOR2_X1 U567 ( .A1(n236), .A2(n535), .ZN(n223) );
  OAI21_X1 U568 ( .B1(n233), .B2(n535), .A(n228), .ZN(n224) );
  INV_X1 U569 ( .A(n188), .ZN(n187) );
  INV_X1 U570 ( .A(n262), .ZN(n260) );
  INV_X1 U571 ( .A(n261), .ZN(n259) );
  NOR2_X1 U572 ( .A1(n252), .A2(n247), .ZN(n243) );
  OAI21_X1 U573 ( .B1(n253), .B2(n247), .A(n248), .ZN(n244) );
  OAI21_X1 U574 ( .B1(n543), .B2(n190), .A(n183), .ZN(n181) );
  AOI21_X1 U575 ( .B1(n158), .B2(n181), .A(n159), .ZN(n157) );
  OAI21_X1 U576 ( .B1(n301), .B2(n307), .A(n302), .ZN(n300) );
  AOI21_X1 U577 ( .B1(n341), .B2(n349), .A(n342), .ZN(n340) );
  NOR2_X1 U578 ( .A1(n346), .A2(n343), .ZN(n341) );
  OAI21_X1 U579 ( .B1(n343), .B2(n347), .A(n344), .ZN(n342) );
  AOI21_X1 U580 ( .B1(n523), .B2(n68), .A(n59), .ZN(n57) );
  INV_X1 U581 ( .A(n61), .ZN(n59) );
  NOR2_X1 U582 ( .A1(n103), .A2(n531), .ZN(n96) );
  OAI21_X1 U583 ( .B1(n256), .B2(n262), .A(n257), .ZN(n255) );
  OAI21_X1 U584 ( .B1(n313), .B2(n317), .A(n314), .ZN(n312) );
  OAI21_X1 U585 ( .B1(n332), .B2(n338), .A(n333), .ZN(n331) );
  OAI21_X1 U586 ( .B1(n350), .B2(n353), .A(n351), .ZN(n349) );
  OAI21_X1 U587 ( .B1(n340), .B2(n320), .A(n321), .ZN(n319) );
  AOI21_X1 U588 ( .B1(n322), .B2(n331), .A(n323), .ZN(n321) );
  NAND2_X1 U589 ( .A1(n330), .A2(n322), .ZN(n320) );
  OAI21_X1 U590 ( .B1(n324), .B2(n328), .A(n325), .ZN(n323) );
  INV_X1 U591 ( .A(n104), .ZN(n102) );
  NOR2_X1 U592 ( .A1(n94), .A2(n87), .ZN(n85) );
  OAI21_X1 U593 ( .B1(n95), .B2(n87), .A(n90), .ZN(n86) );
  INV_X1 U594 ( .A(n88), .ZN(n87) );
  NOR2_X1 U595 ( .A1(n327), .A2(n324), .ZN(n322) );
  AOI21_X1 U596 ( .B1(n238), .B2(n255), .A(n239), .ZN(n237) );
  NOR2_X1 U597 ( .A1(n316), .A2(n313), .ZN(n311) );
  OAI21_X1 U598 ( .B1(n98), .B2(n104), .A(n99), .ZN(n97) );
  NOR2_X1 U599 ( .A1(n337), .A2(n332), .ZN(n330) );
  AOI21_X1 U600 ( .B1(n292), .B2(n381), .A(n289), .ZN(n287) );
  INV_X1 U601 ( .A(n291), .ZN(n289) );
  AOI21_X1 U602 ( .B1(n308), .B2(n383), .A(n305), .ZN(n303) );
  INV_X1 U603 ( .A(n307), .ZN(n305) );
  AOI21_X1 U604 ( .B1(n339), .B2(n389), .A(n336), .ZN(n334) );
  INV_X1 U605 ( .A(n338), .ZN(n336) );
  AOI21_X1 U606 ( .B1(n278), .B2(n379), .A(n275), .ZN(n273) );
  INV_X1 U607 ( .A(n277), .ZN(n275) );
  INV_X1 U608 ( .A(n69), .ZN(n67) );
  NOR2_X1 U609 ( .A1(n89), .A2(n532), .ZN(n80) );
  OAI21_X1 U610 ( .B1(n318), .B2(n316), .A(n317), .ZN(n315) );
  OAI21_X1 U611 ( .B1(n329), .B2(n327), .A(n328), .ZN(n326) );
  AOI21_X1 U612 ( .B1(n538), .B2(n167), .A(n168), .ZN(n166) );
  INV_X1 U613 ( .A(n170), .ZN(n168) );
  OAI21_X1 U614 ( .B1(n348), .B2(n346), .A(n347), .ZN(n345) );
  AOI21_X1 U615 ( .B1(n155), .B2(n365), .A(n146), .ZN(n144) );
  INV_X1 U616 ( .A(n148), .ZN(n146) );
  INV_X1 U617 ( .A(n189), .ZN(n188) );
  AOI21_X1 U618 ( .B1(n121), .B2(n155), .A(n122), .ZN(n120) );
  OAI21_X1 U619 ( .B1(n135), .B2(n123), .A(n126), .ZN(n122) );
  INV_X1 U620 ( .A(n521), .ZN(n365) );
  INV_X1 U621 ( .A(n536), .ZN(n364) );
  INV_X1 U622 ( .A(n89), .ZN(n88) );
  INV_X1 U623 ( .A(n70), .ZN(n68) );
  INV_X1 U624 ( .A(n247), .ZN(n246) );
  INV_X1 U625 ( .A(n525), .ZN(n123) );
  INV_X1 U626 ( .A(n535), .ZN(n226) );
  INV_X1 U627 ( .A(n555), .ZN(n368) );
  OAI21_X1 U628 ( .B1(n215), .B2(n542), .A(n210), .ZN(n206) );
  NOR2_X1 U629 ( .A1(n214), .A2(n542), .ZN(n205) );
  INV_X1 U630 ( .A(n256), .ZN(n376) );
  NAND2_X1 U631 ( .A1(n387), .A2(n328), .ZN(n35) );
  INV_X1 U632 ( .A(n327), .ZN(n387) );
  NAND2_X1 U633 ( .A1(n385), .A2(n317), .ZN(n33) );
  INV_X1 U634 ( .A(n316), .ZN(n385) );
  INV_X1 U635 ( .A(n531), .ZN(n360) );
  NAND2_X1 U636 ( .A1(n386), .A2(n325), .ZN(n34) );
  INV_X1 U637 ( .A(n324), .ZN(n386) );
  NAND2_X1 U638 ( .A1(n381), .A2(n291), .ZN(n29) );
  INV_X1 U639 ( .A(n290), .ZN(n381) );
  NAND2_X1 U640 ( .A1(n383), .A2(n307), .ZN(n31) );
  INV_X1 U641 ( .A(n306), .ZN(n383) );
  NAND2_X1 U642 ( .A1(n389), .A2(n338), .ZN(n37) );
  INV_X1 U643 ( .A(n337), .ZN(n389) );
  NAND2_X1 U644 ( .A1(n391), .A2(n347), .ZN(n39) );
  INV_X1 U645 ( .A(n346), .ZN(n391) );
  NAND2_X1 U646 ( .A1(n379), .A2(n277), .ZN(n27) );
  INV_X1 U647 ( .A(n276), .ZN(n379) );
  NAND2_X1 U648 ( .A1(n390), .A2(n344), .ZN(n38) );
  INV_X1 U649 ( .A(n343), .ZN(n390) );
  NAND2_X1 U650 ( .A1(n384), .A2(n314), .ZN(n32) );
  INV_X1 U651 ( .A(n313), .ZN(n384) );
  NAND2_X1 U652 ( .A1(n380), .A2(n286), .ZN(n28) );
  INV_X1 U653 ( .A(n285), .ZN(n380) );
  NAND2_X1 U654 ( .A1(n382), .A2(n302), .ZN(n30) );
  INV_X1 U655 ( .A(n301), .ZN(n382) );
  NAND2_X1 U656 ( .A1(n388), .A2(n333), .ZN(n36) );
  INV_X1 U657 ( .A(n332), .ZN(n388) );
  NAND2_X1 U658 ( .A1(n392), .A2(n351), .ZN(n40) );
  INV_X1 U659 ( .A(n350), .ZN(n392) );
  INV_X1 U660 ( .A(n202), .ZN(n370) );
  INV_X1 U661 ( .A(n532), .ZN(n358) );
  NAND2_X1 U662 ( .A1(n259), .A2(n262), .ZN(n25) );
  INV_X1 U663 ( .A(n547), .ZN(n362) );
  INV_X1 U664 ( .A(n556), .ZN(n366) );
  NAND2_X1 U665 ( .A1(n361), .A2(n104), .ZN(n9) );
  INV_X1 U666 ( .A(n103), .ZN(n361) );
  INV_X1 U667 ( .A(n271), .ZN(n378) );
  INV_X1 U668 ( .A(n220), .ZN(n372) );
  INV_X1 U669 ( .A(n52), .ZN(n50) );
  NOR2_X1 U670 ( .A1(A[32]), .A2(B[32]), .ZN(n103) );
  NOR2_X1 U671 ( .A1(A[34]), .A2(B[34]), .ZN(n89) );
  NOR2_X1 U672 ( .A1(A[33]), .A2(B[33]), .ZN(n98) );
  NOR2_X1 U673 ( .A1(B[20]), .A2(A[20]), .ZN(n227) );
  NOR2_X1 U674 ( .A1(A[30]), .A2(B[30]), .ZN(n125) );
  NOR2_X1 U675 ( .A1(B[31]), .A2(A[31]), .ZN(n114) );
  NAND2_X1 U676 ( .A1(A[34]), .A2(B[34]), .ZN(n90) );
  NAND2_X1 U677 ( .A1(n188), .A2(n190), .ZN(n17) );
  NAND2_X1 U678 ( .A1(n365), .A2(n148), .ZN(n13) );
  NOR2_X1 U679 ( .A1(A[15]), .A2(B[15]), .ZN(n271) );
  NOR2_X1 U680 ( .A1(A[23]), .A2(B[23]), .ZN(n202) );
  NAND2_X1 U681 ( .A1(A[37]), .A2(B[37]), .ZN(n61) );
  NOR2_X1 U682 ( .A1(A[21]), .A2(B[21]), .ZN(n220) );
  NOR2_X1 U683 ( .A1(A[36]), .A2(B[36]), .ZN(n69) );
  NAND2_X1 U684 ( .A1(A[8]), .A2(B[8]), .ZN(n317) );
  NAND2_X1 U685 ( .A1(A[6]), .A2(B[6]), .ZN(n328) );
  XOR2_X1 U686 ( .A(n329), .B(n35), .Z(SUM[6]) );
  XOR2_X1 U687 ( .A(n162), .B(n14), .Z(SUM[27]) );
  NAND2_X1 U688 ( .A1(n366), .A2(n161), .ZN(n14) );
  XOR2_X1 U689 ( .A(n242), .B(n22), .Z(SUM[19]) );
  NAND2_X1 U690 ( .A1(n374), .A2(n241), .ZN(n22) );
  XOR2_X1 U691 ( .A(n211), .B(n19), .Z(SUM[22]) );
  NAND2_X1 U692 ( .A1(n208), .A2(n210), .ZN(n19) );
  XOR2_X1 U693 ( .A(n184), .B(n16), .Z(SUM[25]) );
  NAND2_X1 U694 ( .A1(n368), .A2(n183), .ZN(n16) );
  NAND2_X1 U695 ( .A1(A[4]), .A2(B[4]), .ZN(n338) );
  NAND2_X1 U696 ( .A1(A[7]), .A2(B[7]), .ZN(n325) );
  NAND2_X1 U697 ( .A1(A[12]), .A2(B[12]), .ZN(n291) );
  NAND2_X1 U698 ( .A1(A[10]), .A2(B[10]), .ZN(n307) );
  NAND2_X1 U699 ( .A1(A[16]), .A2(B[16]), .ZN(n262) );
  NAND2_X1 U700 ( .A1(A[2]), .A2(B[2]), .ZN(n347) );
  NAND2_X1 U701 ( .A1(A[0]), .A2(B[0]), .ZN(n353) );
  NAND2_X1 U702 ( .A1(A[18]), .A2(B[18]), .ZN(n248) );
  NAND2_X1 U703 ( .A1(A[32]), .A2(B[32]), .ZN(n104) );
  NAND2_X1 U704 ( .A1(A[23]), .A2(B[23]), .ZN(n203) );
  NAND2_X1 U705 ( .A1(A[36]), .A2(B[36]), .ZN(n70) );
  NAND2_X1 U706 ( .A1(A[38]), .A2(B[38]), .ZN(n52) );
  NAND2_X1 U707 ( .A1(A[17]), .A2(B[17]), .ZN(n257) );
  NAND2_X1 U708 ( .A1(A[14]), .A2(B[14]), .ZN(n277) );
  NAND2_X1 U709 ( .A1(A[13]), .A2(B[13]), .ZN(n286) );
  NAND2_X1 U710 ( .A1(A[11]), .A2(B[11]), .ZN(n302) );
  NAND2_X1 U711 ( .A1(A[9]), .A2(B[9]), .ZN(n314) );
  NAND2_X1 U712 ( .A1(A[5]), .A2(B[5]), .ZN(n333) );
  NAND2_X1 U713 ( .A1(A[1]), .A2(B[1]), .ZN(n351) );
  NAND2_X1 U714 ( .A1(A[3]), .A2(B[3]), .ZN(n344) );
  NAND2_X1 U715 ( .A1(B[22]), .A2(A[22]), .ZN(n210) );
  NAND2_X1 U716 ( .A1(A[21]), .A2(B[21]), .ZN(n221) );
  NAND2_X1 U717 ( .A1(A[15]), .A2(B[15]), .ZN(n272) );
  NAND2_X1 U718 ( .A1(A[39]), .A2(B[39]), .ZN(n43) );
  NAND2_X1 U719 ( .A1(A[33]), .A2(B[33]), .ZN(n99) );
  NAND2_X1 U720 ( .A1(B[31]), .A2(A[31]), .ZN(n115) );
  XOR2_X1 U721 ( .A(n222), .B(n20), .Z(SUM[21]) );
  NAND2_X1 U722 ( .A1(n372), .A2(n221), .ZN(n20) );
  XOR2_X1 U723 ( .A(n204), .B(n18), .Z(SUM[23]) );
  NAND2_X1 U724 ( .A1(n370), .A2(n203), .ZN(n18) );
  XOR2_X1 U725 ( .A(n258), .B(n24), .Z(SUM[17]) );
  NAND2_X1 U726 ( .A1(n376), .A2(n257), .ZN(n24) );
  XOR2_X1 U727 ( .A(n249), .B(n23), .Z(SUM[18]) );
  NAND2_X1 U728 ( .A1(n246), .A2(n248), .ZN(n23) );
  XOR2_X1 U729 ( .A(n229), .B(n21), .Z(SUM[20]) );
  NAND2_X1 U730 ( .A1(n226), .A2(n228), .ZN(n21) );
  XOR2_X1 U731 ( .A(n171), .B(n15), .Z(SUM[26]) );
  NAND2_X1 U732 ( .A1(n167), .A2(n170), .ZN(n15) );
  XOR2_X1 U733 ( .A(n273), .B(n26), .Z(SUM[15]) );
  NAND2_X1 U734 ( .A1(n378), .A2(n272), .ZN(n26) );
  XOR2_X1 U735 ( .A(n287), .B(n28), .Z(SUM[13]) );
  XNOR2_X1 U736 ( .A(n278), .B(n27), .ZN(SUM[14]) );
  XNOR2_X1 U737 ( .A(n292), .B(n29), .ZN(SUM[12]) );
  XOR2_X1 U738 ( .A(n303), .B(n30), .Z(SUM[11]) );
  XNOR2_X1 U739 ( .A(n308), .B(n31), .ZN(SUM[10]) );
  XNOR2_X1 U740 ( .A(n315), .B(n32), .ZN(SUM[9]) );
  XOR2_X1 U741 ( .A(n40), .B(n353), .Z(SUM[1]) );
  XNOR2_X1 U742 ( .A(n345), .B(n38), .ZN(SUM[3]) );
  XNOR2_X1 U743 ( .A(n339), .B(n37), .ZN(SUM[4]) );
  XOR2_X1 U744 ( .A(n318), .B(n33), .Z(SUM[8]) );
  XNOR2_X1 U745 ( .A(n326), .B(n34), .ZN(SUM[7]) );
  XOR2_X1 U746 ( .A(n334), .B(n36), .Z(SUM[5]) );
  XOR2_X1 U747 ( .A(n348), .B(n39), .Z(SUM[2]) );
  OR2_X1 U748 ( .A1(A[39]), .A2(B[39]), .ZN(n560) );
  INV_X1 U749 ( .A(n542), .ZN(n208) );
  NOR2_X1 U750 ( .A1(n209), .A2(n202), .ZN(n200) );
  NOR2_X1 U751 ( .A1(B[22]), .A2(A[22]), .ZN(n209) );
  NOR2_X1 U752 ( .A1(A[19]), .A2(B[19]), .ZN(n240) );
  NAND2_X1 U753 ( .A1(A[19]), .A2(B[19]), .ZN(n241) );
  OAI21_X1 U754 ( .B1(n240), .B2(n248), .A(n241), .ZN(n239) );
  INV_X1 U755 ( .A(n240), .ZN(n374) );
  INV_X1 U756 ( .A(n79), .ZN(n77) );
  AOI21_X1 U757 ( .B1(n80), .B2(n97), .A(n81), .ZN(n79) );
  AOI21_X1 U758 ( .B1(n55), .B2(n524), .A(n50), .ZN(n48) );
  INV_X1 U759 ( .A(n545), .ZN(n135) );
  NOR2_X1 U760 ( .A1(n138), .A2(n147), .ZN(n136) );
  INV_X1 U761 ( .A(n534), .ZN(n167) );
  XNOR2_X1 U762 ( .A(n263), .B(n25), .ZN(SUM[16]) );
  AOI21_X1 U763 ( .B1(n263), .B2(n192), .A(n193), .ZN(n191) );
  AOI21_X1 U764 ( .B1(n263), .B2(n150), .A(n151), .ZN(n149) );
  AOI21_X1 U765 ( .B1(n263), .B2(n254), .A(n255), .ZN(n249) );
  AOI21_X1 U766 ( .B1(n263), .B2(n243), .A(n244), .ZN(n242) );
  AOI21_X1 U767 ( .B1(n263), .B2(n230), .A(n235), .ZN(n229) );
  AOI21_X1 U768 ( .B1(n263), .B2(n223), .A(n224), .ZN(n222) );
  AOI21_X1 U769 ( .B1(n263), .B2(n212), .A(n213), .ZN(n211) );
  AOI21_X1 U770 ( .B1(n263), .B2(n205), .A(n206), .ZN(n204) );
  AOI21_X1 U771 ( .B1(n263), .B2(n172), .A(n173), .ZN(n171) );
  AOI21_X1 U772 ( .B1(n263), .B2(n259), .A(n260), .ZN(n258) );
  OAI21_X1 U773 ( .B1(n271), .B2(n277), .A(n272), .ZN(n270) );
  XOR2_X1 U774 ( .A(n191), .B(n17), .Z(SUM[24]) );
  NOR2_X1 U775 ( .A1(n236), .A2(n198), .ZN(n196) );
  NAND2_X1 U776 ( .A1(A[24]), .A2(B[24]), .ZN(n190) );
  NOR2_X1 U777 ( .A1(A[24]), .A2(B[24]), .ZN(n189) );
  OAI21_X1 U778 ( .B1(n79), .B2(n56), .A(n57), .ZN(n55) );
  NAND2_X1 U779 ( .A1(A[35]), .A2(B[35]), .ZN(n83) );
  NOR2_X1 U780 ( .A1(n110), .A2(n156), .ZN(n108) );
  NAND2_X1 U781 ( .A1(B[27]), .A2(A[27]), .ZN(n161) );
  NOR2_X1 U782 ( .A1(n189), .A2(n182), .ZN(n180) );
  INV_X1 U783 ( .A(n155), .ZN(n153) );
  NAND2_X1 U784 ( .A1(n218), .A2(n200), .ZN(n198) );
  NOR2_X1 U785 ( .A1(n227), .A2(n220), .ZN(n218) );
  OAI21_X1 U786 ( .B1(n237), .B2(n198), .A(n199), .ZN(n197) );
  AOI21_X1 U787 ( .B1(n263), .B2(n163), .A(n164), .ZN(n162) );
  NAND2_X1 U788 ( .A1(A[25]), .A2(B[25]), .ZN(n183) );
  INV_X1 U789 ( .A(n520), .ZN(n193) );
  AOI21_X1 U790 ( .B1(n200), .B2(n219), .A(n201), .ZN(n199) );
  NAND2_X1 U791 ( .A1(A[20]), .A2(B[20]), .ZN(n228) );
  XOR2_X1 U792 ( .A(n149), .B(n13), .Z(SUM[28]) );
  INV_X1 U793 ( .A(n154), .ZN(n152) );
  INV_X1 U794 ( .A(n196), .ZN(n194) );
  INV_X1 U795 ( .A(n197), .ZN(n195) );
  AOI21_X1 U796 ( .B1(n263), .B2(n128), .A(n129), .ZN(n127) );
  NAND2_X1 U797 ( .A1(B[28]), .A2(A[28]), .ZN(n148) );
  NOR2_X1 U798 ( .A1(B[28]), .A2(A[28]), .ZN(n147) );
  AOI21_X1 U799 ( .B1(n263), .B2(n141), .A(n142), .ZN(n140) );
  AOI21_X1 U800 ( .B1(n263), .B2(n185), .A(n186), .ZN(n184) );
  OAI21_X1 U801 ( .B1(n220), .B2(n228), .A(n221), .ZN(n219) );
  NAND2_X1 U802 ( .A1(n96), .A2(n80), .ZN(n78) );
  AOI21_X1 U803 ( .B1(n263), .B2(n117), .A(n118), .ZN(n116) );
  NOR2_X1 U804 ( .A1(n194), .A2(n537), .ZN(n172) );
  NOR2_X1 U805 ( .A1(n194), .A2(n165), .ZN(n163) );
  NOR2_X1 U806 ( .A1(n194), .A2(n152), .ZN(n150) );
  NOR2_X1 U807 ( .A1(n194), .A2(n143), .ZN(n141) );
  NOR2_X1 U808 ( .A1(n194), .A2(n130), .ZN(n128) );
  NOR2_X1 U809 ( .A1(n194), .A2(n119), .ZN(n117) );
  NOR2_X1 U810 ( .A1(n194), .A2(n187), .ZN(n185) );
  OAI21_X1 U811 ( .B1(n195), .B2(n187), .A(n190), .ZN(n186) );
  OAI21_X1 U812 ( .B1(n195), .B2(n537), .A(n179), .ZN(n173) );
  OAI21_X1 U813 ( .B1(n195), .B2(n152), .A(n153), .ZN(n151) );
  OAI21_X1 U814 ( .B1(n195), .B2(n165), .A(n166), .ZN(n164) );
  OAI21_X1 U815 ( .B1(n520), .B2(n143), .A(n144), .ZN(n142) );
  OAI21_X1 U816 ( .B1(n520), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U817 ( .B1(n520), .B2(n119), .A(n120), .ZN(n118) );
  OAI21_X1 U818 ( .B1(n202), .B2(n210), .A(n203), .ZN(n201) );
  OAI21_X1 U819 ( .B1(n82), .B2(n90), .A(n83), .ZN(n81) );
  NAND2_X1 U820 ( .A1(n180), .A2(n539), .ZN(n156) );
  NOR2_X1 U821 ( .A1(n160), .A2(n169), .ZN(n158) );
  NAND2_X1 U822 ( .A1(A[26]), .A2(B[26]), .ZN(n170) );
  NOR2_X1 U823 ( .A1(A[26]), .A2(B[26]), .ZN(n169) );
  AOI21_X1 U824 ( .B1(n108), .B2(n197), .A(n109), .ZN(n107) );
  NAND2_X1 U825 ( .A1(n108), .A2(n196), .ZN(n106) );
  OAI21_X1 U826 ( .B1(n546), .B2(n170), .A(n161), .ZN(n159) );
  OAI21_X1 U827 ( .B1(n157), .B2(n110), .A(n111), .ZN(n109) );
  AOI21_X1 U828 ( .B1(n137), .B2(n544), .A(n113), .ZN(n111) );
  NAND2_X1 U829 ( .A1(n136), .A2(n112), .ZN(n110) );
  NAND2_X1 U830 ( .A1(A[30]), .A2(B[30]), .ZN(n126) );
  NOR2_X1 U831 ( .A1(n125), .A2(n114), .ZN(n112) );
  XNOR2_X1 U832 ( .A(n1), .B(n9), .ZN(SUM[32]) );
  AOI21_X1 U833 ( .B1(n540), .B2(n527), .A(n46), .ZN(n44) );
  AOI21_X1 U834 ( .B1(n540), .B2(n76), .A(n77), .ZN(n71) );
  AOI21_X1 U835 ( .B1(n540), .B2(n96), .A(n93), .ZN(n91) );
  AOI21_X1 U836 ( .B1(n541), .B2(n63), .A(n64), .ZN(n62) );
  AOI21_X1 U837 ( .B1(n541), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U838 ( .B1(n541), .B2(n54), .A(n55), .ZN(n53) );
  AOI21_X1 U839 ( .B1(n540), .B2(n361), .A(n102), .ZN(n100) );
  OAI21_X1 U840 ( .B1(n559), .B2(n148), .A(n139), .ZN(n137) );
  NAND2_X1 U841 ( .A1(B[29]), .A2(A[29]), .ZN(n139) );
  NOR2_X1 U842 ( .A1(A[29]), .A2(B[29]), .ZN(n138) );
  OAI21_X1 U843 ( .B1(n114), .B2(n126), .A(n115), .ZN(n113) );
endmodule


module datapath_DW01_add_13 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n9, n10, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n43, n44, n46, n48, n50, n52, n53, n54, n55, n56, n57,
         n59, n61, n62, n63, n64, n67, n68, n69, n70, n71, n72, n75, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n88, n89, n90, n91, n93, n94,
         n95, n96, n97, n98, n99, n100, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n179, n180,
         n181, n182, n183, n184, n185, n186, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n218, n219, n220, n221, n222, n223, n224, n226, n227, n228,
         n229, n230, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n246, n247, n248, n249, n252, n253, n254, n255, n256, n257,
         n258, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n275, n276, n277, n278, n279, n280, n283,
         n284, n285, n286, n287, n289, n290, n291, n292, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n353, n358, n360,
         n361, n362, n364, n368, n370, n372, n374, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n520, n521, n522, n523, n524, n525, n526, n527, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554;

  OAI21_X1 U437 ( .B1(n106), .B2(n264), .A(n107), .ZN(n520) );
  OAI21_X1 U438 ( .B1(n106), .B2(n264), .A(n107), .ZN(n105) );
  CLKBUF_X1 U439 ( .A(n157), .Z(n533) );
  CLKBUF_X1 U440 ( .A(n137), .Z(n535) );
  CLKBUF_X1 U441 ( .A(n147), .Z(n521) );
  OAI21_X1 U442 ( .B1(n182), .B2(n190), .A(n183), .ZN(n522) );
  CLKBUF_X1 U443 ( .A(n190), .Z(n523) );
  NOR2_X1 U444 ( .A1(n169), .A2(n160), .ZN(n524) );
  NOR2_X1 U445 ( .A1(B[27]), .A2(A[27]), .ZN(n525) );
  NOR2_X1 U446 ( .A1(n247), .A2(n240), .ZN(n238) );
  NOR2_X1 U447 ( .A1(A[11]), .A2(B[11]), .ZN(n301) );
  OR2_X1 U448 ( .A1(A[37]), .A2(B[37]), .ZN(n526) );
  OR2_X1 U449 ( .A1(A[38]), .A2(B[38]), .ZN(n527) );
  AND2_X1 U450 ( .A1(n530), .A2(n353), .ZN(SUM[0]) );
  AND2_X1 U451 ( .A1(n54), .A2(n527), .ZN(n529) );
  OR2_X1 U452 ( .A1(A[0]), .A2(B[0]), .ZN(n530) );
  NOR2_X1 U453 ( .A1(n209), .A2(n202), .ZN(n200) );
  CLKBUF_X1 U454 ( .A(n218), .Z(n531) );
  CLKBUF_X1 U455 ( .A(n125), .Z(n532) );
  NOR2_X1 U456 ( .A1(A[25]), .A2(B[25]), .ZN(n534) );
  OR2_X1 U457 ( .A1(A[27]), .A2(B[27]), .ZN(n536) );
  NOR2_X1 U458 ( .A1(n156), .A2(n110), .ZN(n537) );
  CLKBUF_X1 U459 ( .A(n227), .Z(n538) );
  NOR2_X1 U460 ( .A1(A[29]), .A2(B[29]), .ZN(n539) );
  CLKBUF_X1 U461 ( .A(n114), .Z(n540) );
  CLKBUF_X1 U462 ( .A(n189), .Z(n541) );
  CLKBUF_X1 U463 ( .A(n169), .Z(n542) );
  CLKBUF_X1 U464 ( .A(n522), .Z(n543) );
  CLKBUF_X1 U465 ( .A(n180), .Z(n544) );
  NOR2_X1 U466 ( .A1(B[27]), .A2(A[27]), .ZN(n160) );
  XNOR2_X1 U467 ( .A(n71), .B(n545), .ZN(SUM[36]) );
  AND2_X1 U468 ( .A1(n67), .A2(n70), .ZN(n545) );
  XNOR2_X1 U469 ( .A(n100), .B(n546), .ZN(SUM[33]) );
  AND2_X1 U470 ( .A1(n360), .A2(n99), .ZN(n546) );
  XNOR2_X1 U471 ( .A(n62), .B(n547), .ZN(SUM[37]) );
  AND2_X1 U472 ( .A1(n526), .A2(n61), .ZN(n547) );
  XNOR2_X1 U473 ( .A(n84), .B(n548), .ZN(SUM[35]) );
  AND2_X1 U474 ( .A1(n358), .A2(n83), .ZN(n548) );
  XNOR2_X1 U475 ( .A(n44), .B(n549), .ZN(SUM[39]) );
  AND2_X1 U476 ( .A1(n554), .A2(n43), .ZN(n549) );
  XNOR2_X1 U477 ( .A(n53), .B(n550), .ZN(SUM[38]) );
  AND2_X1 U478 ( .A1(n527), .A2(n52), .ZN(n550) );
  XNOR2_X1 U479 ( .A(n91), .B(n551), .ZN(SUM[34]) );
  AND2_X1 U480 ( .A1(n88), .A2(n90), .ZN(n551) );
  OR2_X1 U481 ( .A1(n521), .A2(n138), .ZN(n552) );
  NOR2_X1 U482 ( .A1(A[24]), .A2(B[24]), .ZN(n189) );
  NOR2_X1 U483 ( .A1(n147), .A2(n138), .ZN(n136) );
  INV_X1 U484 ( .A(n156), .ZN(n154) );
  NOR2_X1 U485 ( .A1(A[28]), .A2(B[28]), .ZN(n147) );
  NOR2_X1 U486 ( .A1(A[25]), .A2(B[25]), .ZN(n182) );
  INV_X2 U487 ( .A(n264), .ZN(n263) );
  AOI21_X1 U488 ( .B1(n238), .B2(n255), .A(n239), .ZN(n237) );
  AOI21_X1 U489 ( .B1(n299), .B2(n312), .A(n300), .ZN(n298) );
  NOR2_X1 U490 ( .A1(n306), .A2(n301), .ZN(n299) );
  OAI21_X1 U491 ( .B1(n237), .B2(n198), .A(n199), .ZN(n197) );
  NOR2_X1 U492 ( .A1(A[18]), .A2(B[18]), .ZN(n247) );
  NOR2_X1 U493 ( .A1(A[10]), .A2(B[10]), .ZN(n306) );
  NOR2_X1 U494 ( .A1(A[4]), .A2(B[4]), .ZN(n337) );
  NOR2_X1 U495 ( .A1(A[16]), .A2(B[16]), .ZN(n261) );
  NOR2_X1 U496 ( .A1(A[14]), .A2(B[14]), .ZN(n276) );
  NOR2_X1 U497 ( .A1(A[12]), .A2(B[12]), .ZN(n290) );
  NOR2_X1 U498 ( .A1(A[6]), .A2(B[6]), .ZN(n327) );
  NOR2_X1 U499 ( .A1(A[7]), .A2(B[7]), .ZN(n324) );
  NOR2_X1 U500 ( .A1(A[13]), .A2(B[13]), .ZN(n285) );
  NOR2_X1 U501 ( .A1(A[9]), .A2(B[9]), .ZN(n313) );
  NOR2_X1 U502 ( .A1(A[5]), .A2(B[5]), .ZN(n332) );
  NOR2_X1 U503 ( .A1(A[3]), .A2(B[3]), .ZN(n343) );
  NOR2_X1 U504 ( .A1(A[8]), .A2(B[8]), .ZN(n316) );
  NOR2_X1 U505 ( .A1(A[2]), .A2(B[2]), .ZN(n346) );
  NOR2_X1 U506 ( .A1(A[1]), .A2(B[1]), .ZN(n350) );
  INV_X1 U507 ( .A(n196), .ZN(n194) );
  INV_X1 U508 ( .A(n236), .ZN(n230) );
  NAND2_X1 U509 ( .A1(n154), .A2(n132), .ZN(n130) );
  INV_X1 U510 ( .A(n154), .ZN(n152) );
  INV_X1 U511 ( .A(n544), .ZN(n174) );
  INV_X1 U512 ( .A(n194), .ZN(n192) );
  INV_X1 U513 ( .A(n195), .ZN(n193) );
  INV_X1 U514 ( .A(n215), .ZN(n213) );
  INV_X1 U515 ( .A(n214), .ZN(n212) );
  NOR2_X1 U516 ( .A1(n78), .A2(n56), .ZN(n54) );
  INV_X1 U517 ( .A(n95), .ZN(n93) );
  INV_X1 U518 ( .A(n78), .ZN(n72) );
  OAI21_X1 U519 ( .B1(n318), .B2(n297), .A(n298), .ZN(n292) );
  NOR2_X1 U520 ( .A1(n236), .A2(n198), .ZN(n196) );
  AOI21_X1 U521 ( .B1(n155), .B2(n132), .A(n535), .ZN(n131) );
  NAND2_X1 U522 ( .A1(n230), .A2(n531), .ZN(n214) );
  INV_X1 U523 ( .A(n552), .ZN(n132) );
  INV_X1 U524 ( .A(n297), .ZN(n295) );
  INV_X1 U525 ( .A(n155), .ZN(n153) );
  INV_X1 U526 ( .A(n533), .ZN(n155) );
  AOI21_X1 U527 ( .B1(n339), .B2(n330), .A(n331), .ZN(n329) );
  AOI21_X1 U528 ( .B1(n235), .B2(n531), .A(n219), .ZN(n215) );
  NOR2_X1 U529 ( .A1(n78), .A2(n69), .ZN(n63) );
  OAI21_X1 U530 ( .B1(n75), .B2(n69), .A(n70), .ZN(n64) );
  INV_X1 U531 ( .A(n48), .ZN(n46) );
  AOI21_X1 U532 ( .B1(n55), .B2(n527), .A(n50), .ZN(n48) );
  NAND2_X1 U533 ( .A1(n121), .A2(n154), .ZN(n119) );
  NAND2_X1 U534 ( .A1(n154), .A2(n145), .ZN(n143) );
  AOI21_X1 U535 ( .B1(n319), .B2(n265), .A(n266), .ZN(n264) );
  NOR2_X1 U536 ( .A1(n297), .A2(n267), .ZN(n265) );
  OAI21_X1 U537 ( .B1(n298), .B2(n267), .A(n268), .ZN(n266) );
  NAND2_X1 U538 ( .A1(n283), .A2(n269), .ZN(n267) );
  OAI21_X1 U539 ( .B1(n318), .B2(n279), .A(n280), .ZN(n278) );
  AOI21_X1 U540 ( .B1(n296), .B2(n283), .A(n284), .ZN(n280) );
  NAND2_X1 U541 ( .A1(n295), .A2(n283), .ZN(n279) );
  OAI21_X1 U542 ( .B1(n318), .B2(n309), .A(n310), .ZN(n308) );
  INV_X1 U543 ( .A(n312), .ZN(n310) );
  INV_X1 U544 ( .A(n311), .ZN(n309) );
  NOR2_X1 U545 ( .A1(n552), .A2(n532), .ZN(n121) );
  INV_X1 U546 ( .A(n319), .ZN(n318) );
  NAND2_X1 U547 ( .A1(n254), .A2(n238), .ZN(n236) );
  NAND2_X1 U548 ( .A1(n544), .A2(n167), .ZN(n165) );
  INV_X1 U549 ( .A(n535), .ZN(n135) );
  INV_X1 U550 ( .A(n96), .ZN(n94) );
  INV_X1 U551 ( .A(n254), .ZN(n252) );
  NAND2_X1 U552 ( .A1(n218), .A2(n200), .ZN(n198) );
  INV_X1 U553 ( .A(n197), .ZN(n195) );
  NAND2_X1 U554 ( .A1(n311), .A2(n299), .ZN(n297) );
  INV_X1 U555 ( .A(n340), .ZN(n339) );
  INV_X1 U556 ( .A(n255), .ZN(n253) );
  INV_X1 U557 ( .A(n97), .ZN(n95) );
  INV_X1 U558 ( .A(n77), .ZN(n75) );
  INV_X1 U559 ( .A(n298), .ZN(n296) );
  INV_X1 U560 ( .A(n349), .ZN(n348) );
  INV_X1 U561 ( .A(n543), .ZN(n179) );
  INV_X1 U562 ( .A(n237), .ZN(n235) );
  NAND2_X1 U563 ( .A1(n67), .A2(n526), .ZN(n56) );
  OAI21_X1 U564 ( .B1(n256), .B2(n262), .A(n257), .ZN(n255) );
  NOR2_X1 U565 ( .A1(n276), .A2(n271), .ZN(n269) );
  NOR2_X1 U566 ( .A1(n227), .A2(n220), .ZN(n218) );
  AOI21_X1 U567 ( .B1(n526), .B2(n68), .A(n59), .ZN(n57) );
  INV_X1 U568 ( .A(n61), .ZN(n59) );
  NOR2_X1 U569 ( .A1(n236), .A2(n538), .ZN(n223) );
  OAI21_X1 U570 ( .B1(n237), .B2(n538), .A(n228), .ZN(n224) );
  INV_X1 U571 ( .A(n262), .ZN(n260) );
  NOR2_X1 U572 ( .A1(n252), .A2(n247), .ZN(n243) );
  OAI21_X1 U573 ( .B1(n253), .B2(n247), .A(n248), .ZN(n244) );
  OAI21_X1 U574 ( .B1(n182), .B2(n190), .A(n183), .ZN(n181) );
  OAI21_X1 U575 ( .B1(n98), .B2(n104), .A(n99), .ZN(n97) );
  OAI21_X1 U576 ( .B1(n301), .B2(n307), .A(n302), .ZN(n300) );
  AOI21_X1 U577 ( .B1(n341), .B2(n349), .A(n342), .ZN(n340) );
  NOR2_X1 U578 ( .A1(n346), .A2(n343), .ZN(n341) );
  OAI21_X1 U579 ( .B1(n343), .B2(n347), .A(n344), .ZN(n342) );
  OAI21_X1 U580 ( .B1(n332), .B2(n338), .A(n333), .ZN(n331) );
  AOI21_X1 U581 ( .B1(n181), .B2(n524), .A(n159), .ZN(n157) );
  OAI21_X1 U582 ( .B1(n313), .B2(n317), .A(n314), .ZN(n312) );
  OAI21_X1 U583 ( .B1(n285), .B2(n291), .A(n286), .ZN(n284) );
  OAI21_X1 U584 ( .B1(n350), .B2(n353), .A(n351), .ZN(n349) );
  OAI21_X1 U585 ( .B1(n340), .B2(n320), .A(n321), .ZN(n319) );
  AOI21_X1 U586 ( .B1(n322), .B2(n331), .A(n323), .ZN(n321) );
  NAND2_X1 U587 ( .A1(n330), .A2(n322), .ZN(n320) );
  OAI21_X1 U588 ( .B1(n324), .B2(n328), .A(n325), .ZN(n323) );
  NOR2_X1 U589 ( .A1(n94), .A2(n89), .ZN(n85) );
  OAI21_X1 U590 ( .B1(n95), .B2(n89), .A(n90), .ZN(n86) );
  INV_X1 U591 ( .A(n104), .ZN(n102) );
  NOR2_X1 U592 ( .A1(n327), .A2(n324), .ZN(n322) );
  NOR2_X1 U593 ( .A1(n337), .A2(n332), .ZN(n330) );
  NOR2_X1 U594 ( .A1(n316), .A2(n313), .ZN(n311) );
  NOR2_X1 U595 ( .A1(n290), .A2(n285), .ZN(n283) );
  AOI21_X1 U596 ( .B1(n269), .B2(n284), .A(n270), .ZN(n268) );
  AOI21_X1 U597 ( .B1(n292), .B2(n381), .A(n289), .ZN(n287) );
  INV_X1 U598 ( .A(n291), .ZN(n289) );
  AOI21_X1 U599 ( .B1(n308), .B2(n383), .A(n305), .ZN(n303) );
  INV_X1 U600 ( .A(n307), .ZN(n305) );
  AOI21_X1 U601 ( .B1(n339), .B2(n389), .A(n336), .ZN(n334) );
  INV_X1 U602 ( .A(n338), .ZN(n336) );
  AOI21_X1 U603 ( .B1(n278), .B2(n379), .A(n275), .ZN(n273) );
  INV_X1 U604 ( .A(n277), .ZN(n275) );
  INV_X1 U605 ( .A(n542), .ZN(n167) );
  INV_X1 U606 ( .A(n521), .ZN(n145) );
  INV_X1 U607 ( .A(n69), .ZN(n67) );
  INV_X1 U608 ( .A(n209), .ZN(n208) );
  NOR2_X1 U609 ( .A1(n89), .A2(n82), .ZN(n80) );
  OAI21_X1 U610 ( .B1(n318), .B2(n316), .A(n317), .ZN(n315) );
  OAI21_X1 U611 ( .B1(n329), .B2(n327), .A(n328), .ZN(n326) );
  OAI21_X1 U612 ( .B1(n348), .B2(n346), .A(n347), .ZN(n345) );
  AOI21_X1 U613 ( .B1(n121), .B2(n155), .A(n122), .ZN(n120) );
  OAI21_X1 U614 ( .B1(n135), .B2(n532), .A(n126), .ZN(n122) );
  AOI21_X1 U615 ( .B1(n155), .B2(n145), .A(n146), .ZN(n144) );
  INV_X1 U616 ( .A(n148), .ZN(n146) );
  AOI21_X1 U617 ( .B1(n543), .B2(n167), .A(n168), .ZN(n166) );
  INV_X1 U618 ( .A(n170), .ZN(n168) );
  INV_X1 U619 ( .A(n539), .ZN(n364) );
  INV_X1 U620 ( .A(n70), .ZN(n68) );
  INV_X1 U621 ( .A(n247), .ZN(n246) );
  INV_X1 U622 ( .A(n89), .ZN(n88) );
  INV_X1 U623 ( .A(n541), .ZN(n188) );
  INV_X1 U624 ( .A(n534), .ZN(n368) );
  NOR2_X1 U625 ( .A1(n214), .A2(n207), .ZN(n205) );
  INV_X1 U626 ( .A(n208), .ZN(n207) );
  NAND2_X1 U627 ( .A1(n387), .A2(n328), .ZN(n35) );
  INV_X1 U628 ( .A(n327), .ZN(n387) );
  NAND2_X1 U629 ( .A1(n385), .A2(n317), .ZN(n33) );
  INV_X1 U630 ( .A(n316), .ZN(n385) );
  NAND2_X1 U631 ( .A1(n386), .A2(n325), .ZN(n34) );
  INV_X1 U632 ( .A(n324), .ZN(n386) );
  NAND2_X1 U633 ( .A1(n378), .A2(n272), .ZN(n26) );
  INV_X1 U634 ( .A(n271), .ZN(n378) );
  NAND2_X1 U635 ( .A1(n389), .A2(n338), .ZN(n37) );
  INV_X1 U636 ( .A(n337), .ZN(n389) );
  NAND2_X1 U637 ( .A1(n381), .A2(n291), .ZN(n29) );
  INV_X1 U638 ( .A(n290), .ZN(n381) );
  NAND2_X1 U639 ( .A1(n383), .A2(n307), .ZN(n31) );
  INV_X1 U640 ( .A(n306), .ZN(n383) );
  NAND2_X1 U641 ( .A1(n388), .A2(n333), .ZN(n36) );
  INV_X1 U642 ( .A(n332), .ZN(n388) );
  NAND2_X1 U643 ( .A1(n391), .A2(n347), .ZN(n39) );
  INV_X1 U644 ( .A(n346), .ZN(n391) );
  NAND2_X1 U645 ( .A1(n379), .A2(n277), .ZN(n27) );
  INV_X1 U646 ( .A(n276), .ZN(n379) );
  INV_X1 U647 ( .A(n220), .ZN(n372) );
  INV_X1 U648 ( .A(n202), .ZN(n370) );
  NAND2_X1 U649 ( .A1(n390), .A2(n344), .ZN(n38) );
  INV_X1 U650 ( .A(n343), .ZN(n390) );
  NAND2_X1 U651 ( .A1(n384), .A2(n314), .ZN(n32) );
  INV_X1 U652 ( .A(n313), .ZN(n384) );
  INV_X1 U653 ( .A(n98), .ZN(n360) );
  NAND2_X1 U654 ( .A1(n382), .A2(n302), .ZN(n30) );
  INV_X1 U655 ( .A(n301), .ZN(n382) );
  NAND2_X1 U656 ( .A1(n380), .A2(n286), .ZN(n28) );
  INV_X1 U657 ( .A(n285), .ZN(n380) );
  NAND2_X1 U658 ( .A1(n392), .A2(n351), .ZN(n40) );
  INV_X1 U659 ( .A(n350), .ZN(n392) );
  INV_X1 U660 ( .A(n540), .ZN(n362) );
  NAND2_X1 U661 ( .A1(n377), .A2(n262), .ZN(n25) );
  INV_X1 U662 ( .A(n261), .ZN(n377) );
  INV_X1 U663 ( .A(n82), .ZN(n358) );
  INV_X1 U664 ( .A(n103), .ZN(n361) );
  INV_X1 U665 ( .A(n256), .ZN(n376) );
  INV_X1 U666 ( .A(n52), .ZN(n50) );
  NOR2_X1 U667 ( .A1(A[21]), .A2(B[21]), .ZN(n220) );
  NOR2_X1 U668 ( .A1(A[23]), .A2(B[23]), .ZN(n202) );
  NOR2_X1 U669 ( .A1(B[26]), .A2(A[26]), .ZN(n169) );
  NOR2_X1 U670 ( .A1(A[33]), .A2(B[33]), .ZN(n98) );
  NOR2_X1 U671 ( .A1(B[31]), .A2(A[31]), .ZN(n114) );
  NOR2_X1 U672 ( .A1(A[20]), .A2(B[20]), .ZN(n227) );
  NOR2_X1 U673 ( .A1(A[34]), .A2(B[34]), .ZN(n89) );
  NAND2_X1 U674 ( .A1(B[26]), .A2(A[26]), .ZN(n170) );
  NAND2_X1 U675 ( .A1(n362), .A2(n115), .ZN(n10) );
  NAND2_X1 U676 ( .A1(n364), .A2(n139), .ZN(n12) );
  NOR2_X1 U677 ( .A1(A[35]), .A2(B[35]), .ZN(n82) );
  NOR2_X1 U678 ( .A1(A[32]), .A2(B[32]), .ZN(n103) );
  NOR2_X1 U679 ( .A1(A[17]), .A2(B[17]), .ZN(n256) );
  NOR2_X1 U680 ( .A1(A[36]), .A2(B[36]), .ZN(n69) );
  NAND2_X1 U681 ( .A1(A[24]), .A2(B[24]), .ZN(n190) );
  NAND2_X1 U682 ( .A1(A[6]), .A2(B[6]), .ZN(n328) );
  NAND2_X1 U683 ( .A1(A[8]), .A2(B[8]), .ZN(n317) );
  XOR2_X1 U684 ( .A(n329), .B(n35), .Z(SUM[6]) );
  XOR2_X1 U685 ( .A(n229), .B(n21), .Z(SUM[20]) );
  NAND2_X1 U686 ( .A1(n226), .A2(n228), .ZN(n21) );
  XOR2_X1 U687 ( .A(n242), .B(n22), .Z(SUM[19]) );
  NAND2_X1 U688 ( .A1(n374), .A2(n241), .ZN(n22) );
  NAND2_X1 U689 ( .A1(A[32]), .A2(B[32]), .ZN(n104) );
  NAND2_X1 U690 ( .A1(A[4]), .A2(B[4]), .ZN(n338) );
  NAND2_X1 U691 ( .A1(A[5]), .A2(B[5]), .ZN(n333) );
  NAND2_X1 U692 ( .A1(A[7]), .A2(B[7]), .ZN(n325) );
  NAND2_X1 U693 ( .A1(A[12]), .A2(B[12]), .ZN(n291) );
  NAND2_X1 U694 ( .A1(A[10]), .A2(B[10]), .ZN(n307) );
  NAND2_X1 U695 ( .A1(A[2]), .A2(B[2]), .ZN(n347) );
  NAND2_X1 U696 ( .A1(A[34]), .A2(B[34]), .ZN(n90) );
  NAND2_X1 U697 ( .A1(A[16]), .A2(B[16]), .ZN(n262) );
  NAND2_X1 U698 ( .A1(A[0]), .A2(B[0]), .ZN(n353) );
  NAND2_X1 U699 ( .A1(A[36]), .A2(B[36]), .ZN(n70) );
  NAND2_X1 U700 ( .A1(A[37]), .A2(B[37]), .ZN(n61) );
  NAND2_X1 U701 ( .A1(A[38]), .A2(B[38]), .ZN(n52) );
  NAND2_X1 U702 ( .A1(A[18]), .A2(B[18]), .ZN(n248) );
  NAND2_X1 U703 ( .A1(A[14]), .A2(B[14]), .ZN(n277) );
  NAND2_X1 U704 ( .A1(A[20]), .A2(B[20]), .ZN(n228) );
  NAND2_X1 U705 ( .A1(A[35]), .A2(B[35]), .ZN(n83) );
  NAND2_X1 U706 ( .A1(A[17]), .A2(B[17]), .ZN(n257) );
  NAND2_X1 U707 ( .A1(A[11]), .A2(B[11]), .ZN(n302) );
  NAND2_X1 U708 ( .A1(A[13]), .A2(B[13]), .ZN(n286) );
  NAND2_X1 U709 ( .A1(A[9]), .A2(B[9]), .ZN(n314) );
  NAND2_X1 U710 ( .A1(A[3]), .A2(B[3]), .ZN(n344) );
  NAND2_X1 U711 ( .A1(A[1]), .A2(B[1]), .ZN(n351) );
  NAND2_X1 U712 ( .A1(A[39]), .A2(B[39]), .ZN(n43) );
  NAND2_X1 U713 ( .A1(A[19]), .A2(B[19]), .ZN(n241) );
  NAND2_X1 U714 ( .A1(A[21]), .A2(B[21]), .ZN(n221) );
  XNOR2_X1 U715 ( .A(n127), .B(n553), .ZN(SUM[30]) );
  AND2_X1 U716 ( .A1(n124), .A2(n126), .ZN(n553) );
  XOR2_X1 U717 ( .A(n149), .B(n13), .Z(SUM[28]) );
  NAND2_X1 U718 ( .A1(n145), .A2(n148), .ZN(n13) );
  NAND2_X1 U719 ( .A1(n361), .A2(n104), .ZN(n9) );
  XNOR2_X1 U720 ( .A(n278), .B(n27), .ZN(SUM[14]) );
  XOR2_X1 U721 ( .A(n40), .B(n353), .Z(SUM[1]) );
  XOR2_X1 U722 ( .A(n348), .B(n39), .Z(SUM[2]) );
  XOR2_X1 U723 ( .A(n184), .B(n16), .Z(SUM[25]) );
  NAND2_X1 U724 ( .A1(n368), .A2(n183), .ZN(n16) );
  XOR2_X1 U725 ( .A(n171), .B(n15), .Z(SUM[26]) );
  NAND2_X1 U726 ( .A1(n167), .A2(n170), .ZN(n15) );
  XOR2_X1 U727 ( .A(n162), .B(n14), .Z(SUM[27]) );
  NAND2_X1 U728 ( .A1(n536), .A2(n161), .ZN(n14) );
  XOR2_X1 U729 ( .A(n222), .B(n20), .Z(SUM[21]) );
  NAND2_X1 U730 ( .A1(n372), .A2(n221), .ZN(n20) );
  XOR2_X1 U731 ( .A(n191), .B(n17), .Z(SUM[24]) );
  NAND2_X1 U732 ( .A1(n188), .A2(n523), .ZN(n17) );
  XOR2_X1 U733 ( .A(n211), .B(n19), .Z(SUM[22]) );
  NAND2_X1 U734 ( .A1(n208), .A2(n210), .ZN(n19) );
  NAND2_X1 U735 ( .A1(n370), .A2(n203), .ZN(n18) );
  XOR2_X1 U736 ( .A(n258), .B(n24), .Z(SUM[17]) );
  NAND2_X1 U737 ( .A1(n376), .A2(n257), .ZN(n24) );
  XOR2_X1 U738 ( .A(n249), .B(n23), .Z(SUM[18]) );
  NAND2_X1 U739 ( .A1(n246), .A2(n248), .ZN(n23) );
  XOR2_X1 U740 ( .A(n273), .B(n26), .Z(SUM[15]) );
  XOR2_X1 U741 ( .A(n287), .B(n28), .Z(SUM[13]) );
  XNOR2_X1 U742 ( .A(n292), .B(n29), .ZN(SUM[12]) );
  XOR2_X1 U743 ( .A(n303), .B(n30), .Z(SUM[11]) );
  XNOR2_X1 U744 ( .A(n308), .B(n31), .ZN(SUM[10]) );
  XNOR2_X1 U745 ( .A(n315), .B(n32), .ZN(SUM[9]) );
  XNOR2_X1 U746 ( .A(n345), .B(n38), .ZN(SUM[3]) );
  XNOR2_X1 U747 ( .A(n339), .B(n37), .ZN(SUM[4]) );
  XOR2_X1 U748 ( .A(n318), .B(n33), .Z(SUM[8]) );
  XNOR2_X1 U749 ( .A(n326), .B(n34), .ZN(SUM[7]) );
  XOR2_X1 U750 ( .A(n334), .B(n36), .Z(SUM[5]) );
  OR2_X1 U751 ( .A1(A[39]), .A2(B[39]), .ZN(n554) );
  NAND2_X1 U752 ( .A1(B[31]), .A2(A[31]), .ZN(n115) );
  NAND2_X1 U753 ( .A1(A[22]), .A2(B[22]), .ZN(n210) );
  NOR2_X1 U754 ( .A1(A[22]), .A2(B[22]), .ZN(n209) );
  INV_X1 U755 ( .A(n538), .ZN(n226) );
  OAI21_X1 U756 ( .B1(n240), .B2(n248), .A(n241), .ZN(n239) );
  INV_X1 U757 ( .A(n240), .ZN(n374) );
  NOR2_X1 U758 ( .A1(A[19]), .A2(B[19]), .ZN(n240) );
  XOR2_X1 U759 ( .A(n140), .B(n12), .Z(SUM[29]) );
  NOR2_X1 U760 ( .A1(n189), .A2(n534), .ZN(n180) );
  XOR2_X1 U761 ( .A(n204), .B(n18), .Z(SUM[23]) );
  OAI21_X1 U762 ( .B1(n215), .B2(n207), .A(n210), .ZN(n206) );
  NOR2_X1 U763 ( .A1(n261), .A2(n256), .ZN(n254) );
  XNOR2_X1 U764 ( .A(n263), .B(n25), .ZN(SUM[16]) );
  AOI21_X1 U765 ( .B1(n263), .B2(n254), .A(n255), .ZN(n249) );
  AOI21_X1 U766 ( .B1(n263), .B2(n243), .A(n244), .ZN(n242) );
  AOI21_X1 U767 ( .B1(n263), .B2(n230), .A(n235), .ZN(n229) );
  AOI21_X1 U768 ( .B1(n263), .B2(n223), .A(n224), .ZN(n222) );
  AOI21_X1 U769 ( .B1(n263), .B2(n212), .A(n213), .ZN(n211) );
  AOI21_X1 U770 ( .B1(n263), .B2(n205), .A(n206), .ZN(n204) );
  AOI21_X1 U771 ( .B1(n263), .B2(n192), .A(n193), .ZN(n191) );
  AOI21_X1 U772 ( .B1(n263), .B2(n377), .A(n260), .ZN(n258) );
  OAI21_X1 U773 ( .B1(n271), .B2(n277), .A(n272), .ZN(n270) );
  NAND2_X1 U774 ( .A1(A[15]), .A2(B[15]), .ZN(n272) );
  NOR2_X1 U775 ( .A1(A[15]), .A2(B[15]), .ZN(n271) );
  XOR2_X1 U776 ( .A(n116), .B(n10), .Z(SUM[31]) );
  INV_X1 U777 ( .A(n532), .ZN(n124) );
  AOI21_X1 U778 ( .B1(n263), .B2(n163), .A(n164), .ZN(n162) );
  INV_X1 U779 ( .A(n79), .ZN(n77) );
  OAI21_X1 U780 ( .B1(n79), .B2(n56), .A(n57), .ZN(n55) );
  NAND2_X1 U781 ( .A1(A[33]), .A2(B[33]), .ZN(n99) );
  AOI21_X1 U782 ( .B1(n263), .B2(n172), .A(n173), .ZN(n171) );
  AOI21_X1 U783 ( .B1(n200), .B2(n219), .A(n201), .ZN(n199) );
  AOI21_X1 U784 ( .B1(n263), .B2(n150), .A(n151), .ZN(n149) );
  AOI21_X1 U785 ( .B1(n263), .B2(n185), .A(n186), .ZN(n184) );
  AOI21_X1 U786 ( .B1(n80), .B2(n97), .A(n81), .ZN(n79) );
  NAND2_X1 U787 ( .A1(n96), .A2(n80), .ZN(n78) );
  AOI21_X1 U788 ( .B1(n263), .B2(n128), .A(n129), .ZN(n127) );
  NAND2_X1 U789 ( .A1(A[28]), .A2(B[28]), .ZN(n148) );
  AOI21_X1 U790 ( .B1(n263), .B2(n141), .A(n142), .ZN(n140) );
  NAND2_X1 U791 ( .A1(B[27]), .A2(A[27]), .ZN(n161) );
  AOI21_X1 U792 ( .B1(n263), .B2(n117), .A(n118), .ZN(n116) );
  NAND2_X1 U793 ( .A1(A[29]), .A2(B[29]), .ZN(n139) );
  NOR2_X1 U794 ( .A1(A[29]), .A2(B[29]), .ZN(n138) );
  NOR2_X1 U795 ( .A1(n194), .A2(n174), .ZN(n172) );
  NOR2_X1 U796 ( .A1(n194), .A2(n165), .ZN(n163) );
  NOR2_X1 U797 ( .A1(n194), .A2(n152), .ZN(n150) );
  NOR2_X1 U798 ( .A1(n194), .A2(n143), .ZN(n141) );
  NOR2_X1 U799 ( .A1(n194), .A2(n130), .ZN(n128) );
  NOR2_X1 U800 ( .A1(n194), .A2(n119), .ZN(n117) );
  NOR2_X1 U801 ( .A1(n194), .A2(n541), .ZN(n185) );
  OAI21_X1 U802 ( .B1(n220), .B2(n228), .A(n221), .ZN(n219) );
  OAI21_X1 U803 ( .B1(n195), .B2(n541), .A(n523), .ZN(n186) );
  OAI21_X1 U804 ( .B1(n195), .B2(n174), .A(n179), .ZN(n173) );
  OAI21_X1 U805 ( .B1(n195), .B2(n165), .A(n166), .ZN(n164) );
  OAI21_X1 U806 ( .B1(n195), .B2(n143), .A(n144), .ZN(n142) );
  OAI21_X1 U807 ( .B1(n195), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U808 ( .B1(n195), .B2(n119), .A(n120), .ZN(n118) );
  OAI21_X1 U809 ( .B1(n195), .B2(n152), .A(n153), .ZN(n151) );
  OAI21_X1 U810 ( .B1(n202), .B2(n210), .A(n203), .ZN(n201) );
  NAND2_X1 U811 ( .A1(A[23]), .A2(B[23]), .ZN(n203) );
  OAI21_X1 U812 ( .B1(n82), .B2(n90), .A(n83), .ZN(n81) );
  NOR2_X1 U813 ( .A1(n103), .A2(n98), .ZN(n96) );
  NOR2_X1 U814 ( .A1(n156), .A2(n110), .ZN(n108) );
  NAND2_X1 U815 ( .A1(A[25]), .A2(B[25]), .ZN(n183) );
  NAND2_X1 U816 ( .A1(n180), .A2(n158), .ZN(n156) );
  NOR2_X1 U817 ( .A1(n169), .A2(n160), .ZN(n158) );
  AOI21_X1 U818 ( .B1(n197), .B2(n537), .A(n109), .ZN(n107) );
  NAND2_X1 U819 ( .A1(n108), .A2(n196), .ZN(n106) );
  OAI21_X1 U820 ( .B1(n157), .B2(n110), .A(n111), .ZN(n109) );
  OAI21_X1 U821 ( .B1(n525), .B2(n170), .A(n161), .ZN(n159) );
  AOI21_X1 U822 ( .B1(n137), .B2(n112), .A(n113), .ZN(n111) );
  NAND2_X1 U823 ( .A1(n112), .A2(n136), .ZN(n110) );
  NAND2_X1 U824 ( .A1(B[30]), .A2(A[30]), .ZN(n126) );
  NOR2_X1 U825 ( .A1(n114), .A2(n125), .ZN(n112) );
  NOR2_X1 U826 ( .A1(B[30]), .A2(A[30]), .ZN(n125) );
  XNOR2_X1 U827 ( .A(n520), .B(n9), .ZN(SUM[32]) );
  AOI21_X1 U828 ( .B1(n520), .B2(n529), .A(n46), .ZN(n44) );
  AOI21_X1 U829 ( .B1(n520), .B2(n72), .A(n77), .ZN(n71) );
  AOI21_X1 U830 ( .B1(n520), .B2(n96), .A(n93), .ZN(n91) );
  AOI21_X1 U831 ( .B1(n105), .B2(n63), .A(n64), .ZN(n62) );
  AOI21_X1 U832 ( .B1(n105), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U833 ( .B1(n105), .B2(n54), .A(n55), .ZN(n53) );
  AOI21_X1 U834 ( .B1(n105), .B2(n361), .A(n102), .ZN(n100) );
  OAI21_X1 U835 ( .B1(n539), .B2(n148), .A(n139), .ZN(n137) );
  OAI21_X1 U836 ( .B1(n114), .B2(n126), .A(n115), .ZN(n113) );
endmodule


module datapath_DW01_add_14 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n43, n44, n46, n48, n50, n52, n53, n54, n55, n56,
         n57, n59, n61, n62, n63, n64, n65, n68, n70, n71, n72, n75, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n88, n89, n90, n91, n93, n94,
         n95, n96, n97, n98, n99, n100, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n125, n126, n127, n128, n129, n130,
         n131, n132, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n179, n180,
         n181, n182, n183, n184, n185, n186, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n233, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n246, n247, n248, n249, n252, n253, n254,
         n255, n256, n257, n258, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n275, n276, n277, n278,
         n279, n280, n283, n284, n285, n286, n287, n289, n290, n291, n292,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n353, n360, n361, n362, n364, n366, n368, n370, n372, n374, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n556, n557;

  OR2_X1 U437 ( .A1(A[35]), .A2(B[35]), .ZN(n520) );
  OAI21_X1 U438 ( .B1(n106), .B2(n264), .A(n107), .ZN(n521) );
  OAI21_X1 U439 ( .B1(n106), .B2(n264), .A(n107), .ZN(n105) );
  CLKBUF_X1 U440 ( .A(n182), .Z(n532) );
  OR2_X1 U441 ( .A1(A[37]), .A2(B[37]), .ZN(n522) );
  OR2_X1 U442 ( .A1(A[36]), .A2(B[36]), .ZN(n523) );
  OR2_X1 U443 ( .A1(A[38]), .A2(B[38]), .ZN(n524) );
  OR2_X1 U444 ( .A1(n529), .A2(n138), .ZN(n525) );
  NOR2_X1 U445 ( .A1(n198), .A2(n236), .ZN(n196) );
  NOR2_X1 U446 ( .A1(n537), .A2(n169), .ZN(n526) );
  CLKBUF_X1 U447 ( .A(n537), .Z(n527) );
  CLKBUF_X1 U448 ( .A(n190), .Z(n528) );
  NOR2_X1 U449 ( .A1(A[28]), .A2(B[28]), .ZN(n529) );
  CLKBUF_X1 U450 ( .A(B[30]), .Z(n530) );
  NOR2_X1 U451 ( .A1(B[31]), .A2(A[31]), .ZN(n531) );
  BUF_X1 U452 ( .A(n549), .Z(n533) );
  CLKBUF_X1 U453 ( .A(n148), .Z(n534) );
  CLKBUF_X1 U454 ( .A(n209), .Z(n535) );
  NOR2_X1 U455 ( .A1(B[25]), .A2(A[25]), .ZN(n536) );
  NOR2_X1 U456 ( .A1(B[25]), .A2(A[25]), .ZN(n182) );
  NOR2_X1 U457 ( .A1(B[27]), .A2(A[27]), .ZN(n537) );
  NOR2_X1 U458 ( .A1(B[27]), .A2(A[27]), .ZN(n160) );
  NOR2_X1 U459 ( .A1(A[31]), .A2(B[31]), .ZN(n538) );
  NOR2_X1 U460 ( .A1(B[31]), .A2(A[31]), .ZN(n114) );
  OAI21_X1 U461 ( .B1(n190), .B2(n532), .A(n183), .ZN(n539) );
  CLKBUF_X1 U462 ( .A(n180), .Z(n540) );
  CLKBUF_X1 U463 ( .A(n189), .Z(n541) );
  NOR2_X1 U464 ( .A1(n110), .A2(n156), .ZN(n542) );
  XNOR2_X1 U465 ( .A(n44), .B(n543), .ZN(SUM[39]) );
  AND2_X1 U466 ( .A1(n557), .A2(n43), .ZN(n543) );
  XNOR2_X1 U467 ( .A(n71), .B(n544), .ZN(SUM[36]) );
  AND2_X1 U468 ( .A1(n523), .A2(n70), .ZN(n544) );
  XNOR2_X1 U469 ( .A(n84), .B(n545), .ZN(SUM[35]) );
  AND2_X1 U470 ( .A1(n520), .A2(n83), .ZN(n545) );
  XNOR2_X1 U471 ( .A(n53), .B(n546), .ZN(SUM[38]) );
  AND2_X1 U472 ( .A1(n524), .A2(n52), .ZN(n546) );
  XNOR2_X1 U473 ( .A(n91), .B(n547), .ZN(SUM[34]) );
  AND2_X1 U474 ( .A1(n88), .A2(n90), .ZN(n547) );
  XNOR2_X1 U475 ( .A(n100), .B(n548), .ZN(SUM[33]) );
  AND2_X1 U476 ( .A1(n360), .A2(n99), .ZN(n548) );
  NOR2_X1 U477 ( .A1(B[29]), .A2(A[29]), .ZN(n549) );
  OAI21_X1 U478 ( .B1(n533), .B2(n148), .A(n139), .ZN(n550) );
  NOR2_X1 U479 ( .A1(n538), .A2(n125), .ZN(n551) );
  OR2_X1 U480 ( .A1(n530), .A2(A[30]), .ZN(n552) );
  XNOR2_X1 U481 ( .A(n62), .B(n553), .ZN(SUM[37]) );
  AND2_X1 U482 ( .A1(n522), .A2(n61), .ZN(n553) );
  INV_X1 U483 ( .A(n48), .ZN(n46) );
  NOR2_X1 U484 ( .A1(A[4]), .A2(B[4]), .ZN(n337) );
  NOR2_X1 U485 ( .A1(A[10]), .A2(B[10]), .ZN(n306) );
  NOR2_X1 U486 ( .A1(A[12]), .A2(B[12]), .ZN(n290) );
  NOR2_X1 U487 ( .A1(A[16]), .A2(B[16]), .ZN(n261) );
  NOR2_X1 U488 ( .A1(A[14]), .A2(B[14]), .ZN(n276) );
  NOR2_X1 U489 ( .A1(A[6]), .A2(B[6]), .ZN(n327) );
  NOR2_X1 U490 ( .A1(A[7]), .A2(B[7]), .ZN(n324) );
  NOR2_X1 U491 ( .A1(A[11]), .A2(B[11]), .ZN(n301) );
  NOR2_X1 U492 ( .A1(A[13]), .A2(B[13]), .ZN(n285) );
  NOR2_X1 U493 ( .A1(A[9]), .A2(B[9]), .ZN(n313) );
  NOR2_X1 U494 ( .A1(A[3]), .A2(B[3]), .ZN(n343) );
  NOR2_X1 U495 ( .A1(A[5]), .A2(B[5]), .ZN(n332) );
  NOR2_X1 U496 ( .A1(A[8]), .A2(B[8]), .ZN(n316) );
  NOR2_X1 U497 ( .A1(A[2]), .A2(B[2]), .ZN(n346) );
  NOR2_X1 U498 ( .A1(A[1]), .A2(B[1]), .ZN(n350) );
  INV_X1 U499 ( .A(n236), .ZN(n230) );
  INV_X1 U500 ( .A(n154), .ZN(n152) );
  NAND2_X1 U501 ( .A1(n154), .A2(n132), .ZN(n130) );
  INV_X1 U502 ( .A(n540), .ZN(n174) );
  INV_X1 U503 ( .A(n155), .ZN(n153) );
  INV_X1 U504 ( .A(n194), .ZN(n192) );
  INV_X1 U505 ( .A(n156), .ZN(n154) );
  INV_X1 U506 ( .A(n95), .ZN(n93) );
  INV_X1 U507 ( .A(n214), .ZN(n212) );
  INV_X1 U508 ( .A(n215), .ZN(n213) );
  OAI21_X1 U509 ( .B1(n318), .B2(n297), .A(n298), .ZN(n292) );
  INV_X1 U510 ( .A(n264), .ZN(n263) );
  NOR2_X1 U511 ( .A1(n78), .A2(n56), .ZN(n54) );
  NAND2_X1 U512 ( .A1(n230), .A2(n216), .ZN(n214) );
  INV_X1 U513 ( .A(n235), .ZN(n233) );
  INV_X1 U514 ( .A(n297), .ZN(n295) );
  INV_X1 U515 ( .A(n525), .ZN(n132) );
  INV_X1 U516 ( .A(n78), .ZN(n72) );
  AOI21_X1 U517 ( .B1(n339), .B2(n330), .A(n331), .ZN(n329) );
  NAND2_X1 U518 ( .A1(n121), .A2(n154), .ZN(n119) );
  AND2_X1 U519 ( .A1(n54), .A2(n524), .ZN(n554) );
  NOR2_X1 U520 ( .A1(n78), .A2(n65), .ZN(n63) );
  OAI21_X1 U521 ( .B1(n75), .B2(n65), .A(n70), .ZN(n64) );
  INV_X1 U522 ( .A(n523), .ZN(n65) );
  AOI21_X1 U523 ( .B1(n319), .B2(n265), .A(n266), .ZN(n264) );
  OAI21_X1 U524 ( .B1(n298), .B2(n267), .A(n268), .ZN(n266) );
  NOR2_X1 U525 ( .A1(n297), .A2(n267), .ZN(n265) );
  AOI21_X1 U526 ( .B1(n269), .B2(n284), .A(n270), .ZN(n268) );
  OAI21_X1 U527 ( .B1(n318), .B2(n279), .A(n280), .ZN(n278) );
  AOI21_X1 U528 ( .B1(n296), .B2(n283), .A(n284), .ZN(n280) );
  NAND2_X1 U529 ( .A1(n295), .A2(n283), .ZN(n279) );
  OAI21_X1 U530 ( .B1(n318), .B2(n309), .A(n310), .ZN(n308) );
  INV_X1 U531 ( .A(n312), .ZN(n310) );
  INV_X1 U532 ( .A(n311), .ZN(n309) );
  INV_X1 U533 ( .A(n319), .ZN(n318) );
  AOI21_X1 U534 ( .B1(n235), .B2(n216), .A(n219), .ZN(n215) );
  NAND2_X1 U535 ( .A1(n254), .A2(n238), .ZN(n236) );
  INV_X1 U536 ( .A(n96), .ZN(n94) );
  INV_X1 U537 ( .A(n550), .ZN(n135) );
  NOR2_X1 U538 ( .A1(n525), .A2(n123), .ZN(n121) );
  INV_X1 U539 ( .A(n254), .ZN(n252) );
  NAND2_X1 U540 ( .A1(n283), .A2(n269), .ZN(n267) );
  NAND2_X1 U541 ( .A1(n311), .A2(n299), .ZN(n297) );
  INV_X1 U542 ( .A(n255), .ZN(n253) );
  INV_X1 U543 ( .A(n340), .ZN(n339) );
  INV_X1 U544 ( .A(n237), .ZN(n235) );
  INV_X1 U545 ( .A(n77), .ZN(n75) );
  INV_X1 U546 ( .A(n298), .ZN(n296) );
  INV_X1 U547 ( .A(n539), .ZN(n179) );
  NAND2_X1 U548 ( .A1(n523), .A2(n522), .ZN(n56) );
  INV_X1 U549 ( .A(n349), .ZN(n348) );
  INV_X1 U550 ( .A(n217), .ZN(n216) );
  INV_X1 U551 ( .A(n218), .ZN(n217) );
  NAND2_X1 U552 ( .A1(n154), .A2(n145), .ZN(n143) );
  OAI21_X1 U553 ( .B1(n256), .B2(n262), .A(n257), .ZN(n255) );
  NOR2_X1 U554 ( .A1(n276), .A2(n271), .ZN(n269) );
  NOR2_X1 U555 ( .A1(n247), .A2(n240), .ZN(n238) );
  AOI21_X1 U556 ( .B1(n522), .B2(n68), .A(n59), .ZN(n57) );
  INV_X1 U557 ( .A(n61), .ZN(n59) );
  NOR2_X1 U558 ( .A1(n94), .A2(n89), .ZN(n85) );
  OAI21_X1 U559 ( .B1(n95), .B2(n89), .A(n90), .ZN(n86) );
  NOR2_X1 U560 ( .A1(n236), .A2(n225), .ZN(n223) );
  OAI21_X1 U561 ( .B1(n233), .B2(n225), .A(n228), .ZN(n224) );
  INV_X1 U562 ( .A(n226), .ZN(n225) );
  INV_X1 U563 ( .A(n262), .ZN(n260) );
  NOR2_X1 U564 ( .A1(n252), .A2(n247), .ZN(n243) );
  OAI21_X1 U565 ( .B1(n253), .B2(n247), .A(n248), .ZN(n244) );
  OAI21_X1 U566 ( .B1(n220), .B2(n228), .A(n221), .ZN(n219) );
  AOI21_X1 U567 ( .B1(n238), .B2(n255), .A(n239), .ZN(n237) );
  AOI21_X1 U568 ( .B1(n299), .B2(n312), .A(n300), .ZN(n298) );
  OAI21_X1 U569 ( .B1(n301), .B2(n307), .A(n302), .ZN(n300) );
  AOI21_X1 U570 ( .B1(n341), .B2(n349), .A(n342), .ZN(n340) );
  NOR2_X1 U571 ( .A1(n346), .A2(n343), .ZN(n341) );
  OAI21_X1 U572 ( .B1(n343), .B2(n347), .A(n344), .ZN(n342) );
  NOR2_X1 U573 ( .A1(n220), .A2(n227), .ZN(n218) );
  OAI21_X1 U574 ( .B1(n313), .B2(n317), .A(n314), .ZN(n312) );
  OAI21_X1 U575 ( .B1(n332), .B2(n338), .A(n333), .ZN(n331) );
  OAI21_X1 U576 ( .B1(n285), .B2(n291), .A(n286), .ZN(n284) );
  OAI21_X1 U577 ( .B1(n350), .B2(n353), .A(n351), .ZN(n349) );
  OAI21_X1 U578 ( .B1(n340), .B2(n320), .A(n321), .ZN(n319) );
  AOI21_X1 U579 ( .B1(n322), .B2(n331), .A(n323), .ZN(n321) );
  NAND2_X1 U580 ( .A1(n330), .A2(n322), .ZN(n320) );
  OAI21_X1 U581 ( .B1(n324), .B2(n328), .A(n325), .ZN(n323) );
  INV_X1 U582 ( .A(n104), .ZN(n102) );
  NOR2_X1 U583 ( .A1(n214), .A2(n535), .ZN(n205) );
  NOR2_X1 U584 ( .A1(n337), .A2(n332), .ZN(n330) );
  NOR2_X1 U585 ( .A1(n327), .A2(n324), .ZN(n322) );
  NOR2_X1 U586 ( .A1(n316), .A2(n313), .ZN(n311) );
  NOR2_X1 U587 ( .A1(n306), .A2(n301), .ZN(n299) );
  OAI21_X1 U588 ( .B1(n135), .B2(n123), .A(n126), .ZN(n122) );
  NOR2_X1 U589 ( .A1(n290), .A2(n285), .ZN(n283) );
  AOI21_X1 U590 ( .B1(n55), .B2(n524), .A(n50), .ZN(n48) );
  INV_X1 U591 ( .A(n52), .ZN(n50) );
  AOI21_X1 U592 ( .B1(n292), .B2(n381), .A(n289), .ZN(n287) );
  INV_X1 U593 ( .A(n291), .ZN(n289) );
  AOI21_X1 U594 ( .B1(n308), .B2(n383), .A(n305), .ZN(n303) );
  INV_X1 U595 ( .A(n307), .ZN(n305) );
  AOI21_X1 U596 ( .B1(n339), .B2(n389), .A(n336), .ZN(n334) );
  INV_X1 U597 ( .A(n338), .ZN(n336) );
  AOI21_X1 U598 ( .B1(n278), .B2(n379), .A(n275), .ZN(n273) );
  INV_X1 U599 ( .A(n277), .ZN(n275) );
  XOR2_X1 U600 ( .A(n329), .B(n35), .Z(SUM[6]) );
  NAND2_X1 U601 ( .A1(n387), .A2(n328), .ZN(n35) );
  INV_X1 U602 ( .A(n529), .ZN(n145) );
  OAI21_X1 U603 ( .B1(n237), .B2(n198), .A(n199), .ZN(n197) );
  OAI21_X1 U604 ( .B1(n318), .B2(n316), .A(n317), .ZN(n315) );
  OAI21_X1 U605 ( .B1(n348), .B2(n346), .A(n347), .ZN(n345) );
  AOI21_X1 U606 ( .B1(n539), .B2(n167), .A(n168), .ZN(n166) );
  INV_X1 U607 ( .A(n170), .ZN(n168) );
  INV_X1 U608 ( .A(n103), .ZN(n361) );
  INV_X1 U609 ( .A(n256), .ZN(n376) );
  INV_X1 U610 ( .A(n533), .ZN(n364) );
  INV_X1 U611 ( .A(n202), .ZN(n370) );
  INV_X1 U612 ( .A(n227), .ZN(n226) );
  INV_X1 U613 ( .A(n552), .ZN(n123) );
  INV_X1 U614 ( .A(n70), .ZN(n68) );
  INV_X1 U615 ( .A(n541), .ZN(n188) );
  INV_X1 U616 ( .A(n535), .ZN(n208) );
  INV_X1 U617 ( .A(n89), .ZN(n88) );
  INV_X1 U618 ( .A(n247), .ZN(n246) );
  INV_X1 U619 ( .A(n538), .ZN(n362) );
  INV_X1 U620 ( .A(n327), .ZN(n387) );
  INV_X1 U621 ( .A(n316), .ZN(n385) );
  INV_X1 U622 ( .A(n346), .ZN(n391) );
  INV_X1 U623 ( .A(n337), .ZN(n389) );
  INV_X1 U624 ( .A(n332), .ZN(n388) );
  INV_X1 U625 ( .A(n285), .ZN(n380) );
  INV_X1 U626 ( .A(n301), .ZN(n382) );
  INV_X1 U627 ( .A(n313), .ZN(n384) );
  INV_X1 U628 ( .A(n343), .ZN(n390) );
  INV_X1 U629 ( .A(n290), .ZN(n381) );
  INV_X1 U630 ( .A(n306), .ZN(n383) );
  INV_X1 U631 ( .A(n220), .ZN(n372) );
  NAND2_X1 U632 ( .A1(n386), .A2(n325), .ZN(n34) );
  INV_X1 U633 ( .A(n324), .ZN(n386) );
  INV_X1 U634 ( .A(n276), .ZN(n379) );
  XOR2_X1 U635 ( .A(n287), .B(n28), .Z(SUM[13]) );
  NAND2_X1 U636 ( .A1(n380), .A2(n286), .ZN(n28) );
  NAND2_X1 U637 ( .A1(n361), .A2(n104), .ZN(n9) );
  XNOR2_X1 U638 ( .A(n278), .B(n27), .ZN(SUM[14]) );
  NAND2_X1 U639 ( .A1(n379), .A2(n277), .ZN(n27) );
  XNOR2_X1 U640 ( .A(n292), .B(n29), .ZN(SUM[12]) );
  NAND2_X1 U641 ( .A1(n381), .A2(n291), .ZN(n29) );
  XOR2_X1 U642 ( .A(n303), .B(n30), .Z(SUM[11]) );
  NAND2_X1 U643 ( .A1(n382), .A2(n302), .ZN(n30) );
  XOR2_X1 U644 ( .A(n40), .B(n353), .Z(SUM[1]) );
  NAND2_X1 U645 ( .A1(n392), .A2(n351), .ZN(n40) );
  XOR2_X1 U646 ( .A(n348), .B(n39), .Z(SUM[2]) );
  NAND2_X1 U647 ( .A1(n391), .A2(n347), .ZN(n39) );
  XNOR2_X1 U648 ( .A(n345), .B(n38), .ZN(SUM[3]) );
  NAND2_X1 U649 ( .A1(n390), .A2(n344), .ZN(n38) );
  XNOR2_X1 U650 ( .A(n339), .B(n37), .ZN(SUM[4]) );
  NAND2_X1 U651 ( .A1(n389), .A2(n338), .ZN(n37) );
  XOR2_X1 U652 ( .A(n334), .B(n36), .Z(SUM[5]) );
  NAND2_X1 U653 ( .A1(n388), .A2(n333), .ZN(n36) );
  XNOR2_X1 U654 ( .A(n308), .B(n31), .ZN(SUM[10]) );
  NAND2_X1 U655 ( .A1(n383), .A2(n307), .ZN(n31) );
  XNOR2_X1 U656 ( .A(n315), .B(n32), .ZN(SUM[9]) );
  NAND2_X1 U657 ( .A1(n384), .A2(n314), .ZN(n32) );
  XOR2_X1 U658 ( .A(n318), .B(n33), .Z(SUM[8]) );
  NAND2_X1 U659 ( .A1(n385), .A2(n317), .ZN(n33) );
  XNOR2_X1 U660 ( .A(n326), .B(n34), .ZN(SUM[7]) );
  OAI21_X1 U661 ( .B1(n329), .B2(n327), .A(n328), .ZN(n326) );
  AND2_X1 U662 ( .A1(n556), .A2(n353), .ZN(SUM[0]) );
  INV_X1 U663 ( .A(n350), .ZN(n392) );
  INV_X1 U664 ( .A(n527), .ZN(n366) );
  INV_X1 U665 ( .A(n534), .ZN(n146) );
  NAND2_X1 U666 ( .A1(n377), .A2(n262), .ZN(n25) );
  INV_X1 U667 ( .A(n261), .ZN(n377) );
  INV_X1 U668 ( .A(n271), .ZN(n378) );
  INV_X1 U669 ( .A(n98), .ZN(n360) );
  NOR2_X1 U670 ( .A1(B[20]), .A2(A[20]), .ZN(n227) );
  NOR2_X1 U671 ( .A1(B[21]), .A2(A[21]), .ZN(n220) );
  OR2_X1 U672 ( .A1(A[0]), .A2(B[0]), .ZN(n556) );
  NOR2_X1 U673 ( .A1(B[22]), .A2(A[22]), .ZN(n209) );
  NOR2_X1 U674 ( .A1(B[24]), .A2(A[24]), .ZN(n189) );
  NOR2_X1 U675 ( .A1(B[26]), .A2(A[26]), .ZN(n169) );
  NOR2_X1 U676 ( .A1(A[35]), .A2(B[35]), .ZN(n82) );
  NOR2_X1 U677 ( .A1(A[18]), .A2(B[18]), .ZN(n247) );
  NAND2_X1 U678 ( .A1(B[30]), .A2(A[30]), .ZN(n126) );
  NAND2_X1 U679 ( .A1(n362), .A2(n115), .ZN(n10) );
  NAND2_X1 U680 ( .A1(n366), .A2(n161), .ZN(n14) );
  NOR2_X1 U681 ( .A1(A[34]), .A2(B[34]), .ZN(n89) );
  NOR2_X1 U682 ( .A1(A[15]), .A2(B[15]), .ZN(n271) );
  NAND2_X1 U683 ( .A1(A[37]), .A2(B[37]), .ZN(n61) );
  NOR2_X1 U684 ( .A1(A[33]), .A2(B[33]), .ZN(n98) );
  NAND2_X1 U685 ( .A1(A[4]), .A2(B[4]), .ZN(n338) );
  NAND2_X1 U686 ( .A1(A[8]), .A2(B[8]), .ZN(n317) );
  NAND2_X1 U687 ( .A1(A[6]), .A2(B[6]), .ZN(n328) );
  XOR2_X1 U688 ( .A(n127), .B(n11), .Z(SUM[30]) );
  NAND2_X1 U689 ( .A1(n552), .A2(n126), .ZN(n11) );
  XOR2_X1 U690 ( .A(n242), .B(n22), .Z(SUM[19]) );
  NAND2_X1 U691 ( .A1(n374), .A2(n241), .ZN(n22) );
  XOR2_X1 U692 ( .A(n258), .B(n24), .Z(SUM[17]) );
  NAND2_X1 U693 ( .A1(n376), .A2(n257), .ZN(n24) );
  XOR2_X1 U694 ( .A(n171), .B(n15), .Z(SUM[26]) );
  NAND2_X1 U695 ( .A1(n167), .A2(n170), .ZN(n15) );
  NAND2_X1 U696 ( .A1(A[7]), .A2(B[7]), .ZN(n325) );
  NAND2_X1 U697 ( .A1(A[12]), .A2(B[12]), .ZN(n291) );
  NAND2_X1 U698 ( .A1(A[10]), .A2(B[10]), .ZN(n307) );
  NAND2_X1 U699 ( .A1(A[2]), .A2(B[2]), .ZN(n347) );
  NAND2_X1 U700 ( .A1(A[34]), .A2(B[34]), .ZN(n90) );
  NAND2_X1 U701 ( .A1(A[38]), .A2(B[38]), .ZN(n52) );
  NAND2_X1 U702 ( .A1(A[0]), .A2(B[0]), .ZN(n353) );
  NAND2_X1 U703 ( .A1(A[18]), .A2(B[18]), .ZN(n248) );
  NAND2_X1 U704 ( .A1(A[16]), .A2(B[16]), .ZN(n262) );
  NAND2_X1 U705 ( .A1(A[14]), .A2(B[14]), .ZN(n277) );
  NAND2_X1 U706 ( .A1(A[36]), .A2(B[36]), .ZN(n70) );
  NAND2_X1 U707 ( .A1(A[33]), .A2(B[33]), .ZN(n99) );
  NAND2_X1 U708 ( .A1(A[5]), .A2(B[5]), .ZN(n333) );
  NAND2_X1 U709 ( .A1(A[13]), .A2(B[13]), .ZN(n286) );
  NAND2_X1 U710 ( .A1(A[11]), .A2(B[11]), .ZN(n302) );
  NAND2_X1 U711 ( .A1(A[3]), .A2(B[3]), .ZN(n344) );
  NAND2_X1 U712 ( .A1(A[9]), .A2(B[9]), .ZN(n314) );
  NAND2_X1 U713 ( .A1(A[1]), .A2(B[1]), .ZN(n351) );
  NAND2_X1 U714 ( .A1(B[22]), .A2(A[22]), .ZN(n210) );
  NAND2_X1 U715 ( .A1(A[39]), .A2(B[39]), .ZN(n43) );
  NAND2_X1 U716 ( .A1(A[15]), .A2(B[15]), .ZN(n272) );
  NAND2_X1 U717 ( .A1(A[21]), .A2(B[21]), .ZN(n221) );
  NAND2_X1 U718 ( .A1(A[19]), .A2(B[19]), .ZN(n241) );
  NAND2_X1 U719 ( .A1(B[25]), .A2(A[25]), .ZN(n183) );
  XOR2_X1 U720 ( .A(n249), .B(n23), .Z(SUM[18]) );
  NAND2_X1 U721 ( .A1(n246), .A2(n248), .ZN(n23) );
  XOR2_X1 U722 ( .A(n222), .B(n20), .Z(SUM[21]) );
  NAND2_X1 U723 ( .A1(n372), .A2(n221), .ZN(n20) );
  XOR2_X1 U724 ( .A(n184), .B(n16), .Z(SUM[25]) );
  NAND2_X1 U725 ( .A1(n368), .A2(n183), .ZN(n16) );
  XOR2_X1 U726 ( .A(n140), .B(n12), .Z(SUM[29]) );
  NAND2_X1 U727 ( .A1(n364), .A2(n139), .ZN(n12) );
  XOR2_X1 U728 ( .A(n191), .B(n17), .Z(SUM[24]) );
  NAND2_X1 U729 ( .A1(n188), .A2(n528), .ZN(n17) );
  XOR2_X1 U730 ( .A(n149), .B(n13), .Z(SUM[28]) );
  NAND2_X1 U731 ( .A1(n145), .A2(n534), .ZN(n13) );
  XOR2_X1 U732 ( .A(n229), .B(n21), .Z(SUM[20]) );
  NAND2_X1 U733 ( .A1(n226), .A2(n228), .ZN(n21) );
  NAND2_X1 U734 ( .A1(n208), .A2(n210), .ZN(n19) );
  NAND2_X1 U735 ( .A1(n370), .A2(n203), .ZN(n18) );
  XOR2_X1 U736 ( .A(n273), .B(n26), .Z(SUM[15]) );
  NAND2_X1 U737 ( .A1(n378), .A2(n272), .ZN(n26) );
  OR2_X1 U738 ( .A1(A[39]), .A2(B[39]), .ZN(n557) );
  AOI21_X1 U739 ( .B1(n200), .B2(n219), .A(n201), .ZN(n199) );
  NAND2_X1 U740 ( .A1(n218), .A2(n200), .ZN(n198) );
  NOR2_X1 U741 ( .A1(n209), .A2(n202), .ZN(n200) );
  NOR2_X1 U742 ( .A1(B[30]), .A2(A[30]), .ZN(n125) );
  XOR2_X1 U743 ( .A(n211), .B(n19), .Z(SUM[22]) );
  OAI21_X1 U744 ( .B1(n215), .B2(n535), .A(n210), .ZN(n206) );
  NOR2_X1 U745 ( .A1(n261), .A2(n256), .ZN(n254) );
  NAND2_X1 U746 ( .A1(A[17]), .A2(B[17]), .ZN(n257) );
  NOR2_X1 U747 ( .A1(A[17]), .A2(B[17]), .ZN(n256) );
  AOI21_X1 U748 ( .B1(n121), .B2(n155), .A(n122), .ZN(n120) );
  AOI21_X1 U749 ( .B1(n155), .B2(n132), .A(n550), .ZN(n131) );
  AOI21_X1 U750 ( .B1(n155), .B2(n145), .A(n146), .ZN(n144) );
  INV_X1 U751 ( .A(n169), .ZN(n167) );
  NOR2_X1 U752 ( .A1(n537), .A2(n169), .ZN(n158) );
  NAND2_X1 U753 ( .A1(B[26]), .A2(A[26]), .ZN(n170) );
  AOI21_X1 U754 ( .B1(n80), .B2(n97), .A(n81), .ZN(n79) );
  NOR2_X1 U755 ( .A1(n89), .A2(n82), .ZN(n80) );
  OAI21_X1 U756 ( .B1(n240), .B2(n248), .A(n241), .ZN(n239) );
  INV_X1 U757 ( .A(n240), .ZN(n374) );
  XOR2_X1 U758 ( .A(n204), .B(n18), .Z(SUM[23]) );
  NOR2_X1 U759 ( .A1(A[19]), .A2(B[19]), .ZN(n240) );
  NAND2_X1 U760 ( .A1(B[27]), .A2(A[27]), .ZN(n161) );
  NOR2_X1 U761 ( .A1(n138), .A2(n147), .ZN(n136) );
  INV_X1 U762 ( .A(n157), .ZN(n155) );
  NOR2_X1 U763 ( .A1(n189), .A2(n536), .ZN(n180) );
  OAI21_X1 U764 ( .B1(n190), .B2(n182), .A(n183), .ZN(n181) );
  XNOR2_X1 U765 ( .A(n263), .B(n25), .ZN(SUM[16]) );
  AOI21_X1 U766 ( .B1(n263), .B2(n254), .A(n255), .ZN(n249) );
  AOI21_X1 U767 ( .B1(n263), .B2(n243), .A(n244), .ZN(n242) );
  AOI21_X1 U768 ( .B1(n263), .B2(n230), .A(n235), .ZN(n229) );
  AOI21_X1 U769 ( .B1(n263), .B2(n223), .A(n224), .ZN(n222) );
  AOI21_X1 U770 ( .B1(n263), .B2(n212), .A(n213), .ZN(n211) );
  AOI21_X1 U771 ( .B1(n263), .B2(n205), .A(n206), .ZN(n204) );
  AOI21_X1 U772 ( .B1(n263), .B2(n192), .A(n193), .ZN(n191) );
  AOI21_X1 U773 ( .B1(n263), .B2(n377), .A(n260), .ZN(n258) );
  OAI21_X1 U774 ( .B1(n271), .B2(n277), .A(n272), .ZN(n270) );
  XOR2_X1 U775 ( .A(n162), .B(n14), .Z(SUM[27]) );
  AOI21_X1 U776 ( .B1(n263), .B2(n163), .A(n164), .ZN(n162) );
  OAI21_X1 U777 ( .B1(n79), .B2(n56), .A(n57), .ZN(n55) );
  INV_X1 U778 ( .A(n79), .ZN(n77) );
  NOR2_X1 U779 ( .A1(A[32]), .A2(B[32]), .ZN(n103) );
  NAND2_X1 U780 ( .A1(A[32]), .A2(B[32]), .ZN(n104) );
  NAND2_X1 U781 ( .A1(A[35]), .A2(B[35]), .ZN(n83) );
  INV_X1 U782 ( .A(n196), .ZN(n194) );
  NAND2_X1 U783 ( .A1(n540), .A2(n167), .ZN(n165) );
  AOI21_X1 U784 ( .B1(n263), .B2(n172), .A(n173), .ZN(n171) );
  NAND2_X1 U785 ( .A1(A[20]), .A2(B[20]), .ZN(n228) );
  AOI21_X1 U786 ( .B1(n263), .B2(n185), .A(n186), .ZN(n184) );
  NAND2_X1 U787 ( .A1(A[23]), .A2(B[23]), .ZN(n203) );
  NOR2_X1 U788 ( .A1(A[23]), .A2(B[23]), .ZN(n202) );
  INV_X1 U789 ( .A(n195), .ZN(n193) );
  INV_X1 U790 ( .A(n197), .ZN(n195) );
  AOI21_X1 U791 ( .B1(n263), .B2(n150), .A(n151), .ZN(n149) );
  AOI21_X1 U792 ( .B1(n158), .B2(n181), .A(n159), .ZN(n157) );
  NAND2_X1 U793 ( .A1(n526), .A2(n180), .ZN(n156) );
  AOI21_X1 U794 ( .B1(n263), .B2(n117), .A(n118), .ZN(n116) );
  NOR2_X1 U795 ( .A1(B[28]), .A2(A[28]), .ZN(n147) );
  NAND2_X1 U796 ( .A1(B[28]), .A2(A[28]), .ZN(n148) );
  AOI21_X1 U797 ( .B1(n263), .B2(n128), .A(n129), .ZN(n127) );
  AOI21_X1 U798 ( .B1(n263), .B2(n141), .A(n142), .ZN(n140) );
  NAND2_X1 U799 ( .A1(B[24]), .A2(A[24]), .ZN(n190) );
  INV_X1 U800 ( .A(n97), .ZN(n95) );
  OAI21_X1 U801 ( .B1(n98), .B2(n104), .A(n99), .ZN(n97) );
  NOR2_X1 U802 ( .A1(n194), .A2(n119), .ZN(n117) );
  NOR2_X1 U803 ( .A1(n194), .A2(n174), .ZN(n172) );
  NOR2_X1 U804 ( .A1(n194), .A2(n165), .ZN(n163) );
  NOR2_X1 U805 ( .A1(n194), .A2(n152), .ZN(n150) );
  NOR2_X1 U806 ( .A1(n194), .A2(n143), .ZN(n141) );
  NOR2_X1 U807 ( .A1(n194), .A2(n130), .ZN(n128) );
  NOR2_X1 U808 ( .A1(n194), .A2(n541), .ZN(n185) );
  OAI21_X1 U809 ( .B1(n202), .B2(n210), .A(n203), .ZN(n201) );
  OAI21_X1 U810 ( .B1(n195), .B2(n119), .A(n120), .ZN(n118) );
  OAI21_X1 U811 ( .B1(n195), .B2(n541), .A(n528), .ZN(n186) );
  OAI21_X1 U812 ( .B1(n195), .B2(n174), .A(n179), .ZN(n173) );
  OAI21_X1 U813 ( .B1(n195), .B2(n152), .A(n153), .ZN(n151) );
  OAI21_X1 U814 ( .B1(n195), .B2(n143), .A(n144), .ZN(n142) );
  OAI21_X1 U815 ( .B1(n195), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U816 ( .B1(n195), .B2(n165), .A(n166), .ZN(n164) );
  INV_X1 U817 ( .A(n532), .ZN(n368) );
  OAI21_X1 U818 ( .B1(n82), .B2(n90), .A(n83), .ZN(n81) );
  NAND2_X1 U819 ( .A1(n96), .A2(n80), .ZN(n78) );
  XOR2_X1 U820 ( .A(n116), .B(n10), .Z(SUM[31]) );
  NOR2_X1 U821 ( .A1(n103), .A2(n98), .ZN(n96) );
  NOR2_X1 U822 ( .A1(n156), .A2(n110), .ZN(n108) );
  NAND2_X1 U823 ( .A1(B[31]), .A2(A[31]), .ZN(n115) );
  AOI21_X1 U824 ( .B1(n197), .B2(n542), .A(n109), .ZN(n107) );
  NAND2_X1 U825 ( .A1(n108), .A2(n196), .ZN(n106) );
  OAI21_X1 U826 ( .B1(n157), .B2(n110), .A(n111), .ZN(n109) );
  OAI21_X1 U827 ( .B1(n160), .B2(n170), .A(n161), .ZN(n159) );
  AOI21_X1 U828 ( .B1(n551), .B2(n137), .A(n113), .ZN(n111) );
  NAND2_X1 U829 ( .A1(n112), .A2(n136), .ZN(n110) );
  NOR2_X1 U830 ( .A1(n125), .A2(n531), .ZN(n112) );
  XNOR2_X1 U831 ( .A(n521), .B(n9), .ZN(SUM[32]) );
  AOI21_X1 U832 ( .B1(n521), .B2(n554), .A(n46), .ZN(n44) );
  AOI21_X1 U833 ( .B1(n521), .B2(n72), .A(n77), .ZN(n71) );
  AOI21_X1 U834 ( .B1(n521), .B2(n96), .A(n93), .ZN(n91) );
  AOI21_X1 U835 ( .B1(n105), .B2(n63), .A(n64), .ZN(n62) );
  AOI21_X1 U836 ( .B1(n105), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U837 ( .B1(n105), .B2(n54), .A(n55), .ZN(n53) );
  AOI21_X1 U838 ( .B1(n105), .B2(n361), .A(n102), .ZN(n100) );
  OAI21_X1 U839 ( .B1(n549), .B2(n148), .A(n139), .ZN(n137) );
  NAND2_X1 U840 ( .A1(B[29]), .A2(A[29]), .ZN(n139) );
  NOR2_X1 U841 ( .A1(B[29]), .A2(A[29]), .ZN(n138) );
  OAI21_X1 U842 ( .B1(n114), .B2(n126), .A(n115), .ZN(n113) );
endmodule


module datapath_DW01_add_15 ( A, B, CI, SUM, CO );
  input [39:0] A;
  input [39:0] B;
  output [39:0] SUM;
  input CI;
  output CO;
  wire   n1, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n43, n44, n46, n48, n50, n52, n53, n54, n55,
         n56, n57, n59, n61, n62, n63, n64, n67, n68, n69, n70, n71, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n88, n89, n90, n91,
         n93, n94, n95, n96, n97, n98, n99, n100, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n179, n180, n181,
         n182, n183, n184, n185, n186, n188, n189, n190, n191, n194, n195,
         n196, n197, n198, n199, n201, n202, n203, n204, n205, n206, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n226, n227, n228, n229, n230, n233,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n246,
         n247, n248, n249, n252, n253, n254, n255, n256, n257, n258, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n275, n276, n277, n278, n279, n280, n283, n284, n285,
         n286, n287, n289, n290, n291, n292, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n353, n358, n360, n361, n362,
         n364, n365, n366, n372, n374, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n561, n562;

  INV_X1 U437 ( .A(n146), .ZN(n520) );
  CLKBUF_X1 U438 ( .A(n161), .Z(n521) );
  NOR2_X2 U439 ( .A1(n236), .A2(n198), .ZN(n196) );
  NOR2_X1 U440 ( .A1(B[25]), .A2(A[25]), .ZN(n522) );
  NAND2_X1 U441 ( .A1(A[22]), .A2(B[22]), .ZN(n210) );
  OR2_X1 U442 ( .A1(A[23]), .A2(B[23]), .ZN(n523) );
  NOR2_X2 U443 ( .A1(A[34]), .A2(B[34]), .ZN(n89) );
  XNOR2_X1 U444 ( .A(n62), .B(n524), .ZN(SUM[37]) );
  AND2_X1 U445 ( .A1(n528), .A2(n61), .ZN(n524) );
  XNOR2_X1 U446 ( .A(n53), .B(n525), .ZN(SUM[38]) );
  AND2_X1 U447 ( .A1(n529), .A2(n52), .ZN(n525) );
  NOR2_X1 U448 ( .A1(A[23]), .A2(B[23]), .ZN(n526) );
  NOR2_X1 U449 ( .A1(n209), .A2(n202), .ZN(n527) );
  NOR2_X1 U450 ( .A1(A[23]), .A2(B[23]), .ZN(n202) );
  NOR2_X1 U451 ( .A1(A[33]), .A2(B[33]), .ZN(n98) );
  BUF_X1 U452 ( .A(n543), .Z(n558) );
  OR2_X1 U453 ( .A1(A[37]), .A2(B[37]), .ZN(n528) );
  OR2_X1 U454 ( .A1(A[38]), .A2(B[38]), .ZN(n529) );
  NOR2_X1 U455 ( .A1(A[20]), .A2(B[20]), .ZN(n227) );
  AND2_X1 U456 ( .A1(n54), .A2(n529), .ZN(n530) );
  NOR2_X1 U457 ( .A1(n156), .A2(n110), .ZN(n531) );
  CLKBUF_X1 U458 ( .A(n147), .Z(n532) );
  BUF_X1 U459 ( .A(n157), .Z(n546) );
  BUF_X2 U460 ( .A(n105), .Z(n552) );
  XNOR2_X1 U461 ( .A(n44), .B(n533), .ZN(SUM[39]) );
  AND2_X1 U462 ( .A1(n561), .A2(n43), .ZN(n533) );
  NOR2_X1 U463 ( .A1(n556), .A2(n169), .ZN(n534) );
  CLKBUF_X1 U464 ( .A(B[25]), .Z(n535) );
  CLKBUF_X1 U465 ( .A(n548), .Z(n536) );
  CLKBUF_X1 U466 ( .A(n556), .Z(n537) );
  NOR2_X1 U467 ( .A1(A[30]), .A2(B[30]), .ZN(n538) );
  CLKBUF_X1 U468 ( .A(n126), .Z(n539) );
  CLKBUF_X1 U469 ( .A(n209), .Z(n540) );
  CLKBUF_X1 U470 ( .A(n181), .Z(n541) );
  NOR2_X1 U471 ( .A1(n548), .A2(n538), .ZN(n542) );
  NOR2_X1 U472 ( .A1(B[29]), .A2(A[29]), .ZN(n543) );
  CLKBUF_X1 U473 ( .A(n538), .Z(n544) );
  CLKBUF_X1 U474 ( .A(n137), .Z(n545) );
  CLKBUF_X1 U475 ( .A(n169), .Z(n547) );
  NOR2_X1 U476 ( .A1(B[31]), .A2(A[31]), .ZN(n548) );
  CLKBUF_X1 U477 ( .A(n180), .Z(n549) );
  CLKBUF_X1 U478 ( .A(n189), .Z(n550) );
  BUF_X1 U479 ( .A(n105), .Z(n1) );
  XNOR2_X1 U480 ( .A(n100), .B(n551), .ZN(SUM[33]) );
  AND2_X1 U481 ( .A1(n360), .A2(n99), .ZN(n551) );
  XNOR2_X1 U482 ( .A(n71), .B(n553), .ZN(SUM[36]) );
  AND2_X1 U483 ( .A1(n67), .A2(n70), .ZN(n553) );
  XNOR2_X1 U484 ( .A(n91), .B(n554), .ZN(SUM[34]) );
  AND2_X1 U485 ( .A1(n88), .A2(n90), .ZN(n554) );
  XNOR2_X1 U486 ( .A(n84), .B(n555), .ZN(SUM[35]) );
  AND2_X1 U487 ( .A1(n358), .A2(n83), .ZN(n555) );
  NOR2_X1 U488 ( .A1(B[27]), .A2(A[27]), .ZN(n556) );
  OR2_X1 U489 ( .A1(n532), .A2(n558), .ZN(n557) );
  OR2_X1 U490 ( .A1(A[25]), .A2(n535), .ZN(n559) );
  NOR2_X1 U491 ( .A1(A[35]), .A2(B[35]), .ZN(n82) );
  NOR2_X1 U492 ( .A1(A[4]), .A2(B[4]), .ZN(n337) );
  NOR2_X1 U493 ( .A1(A[12]), .A2(B[12]), .ZN(n290) );
  NOR2_X1 U494 ( .A1(A[10]), .A2(B[10]), .ZN(n306) );
  NOR2_X1 U495 ( .A1(A[18]), .A2(B[18]), .ZN(n247) );
  NOR2_X1 U496 ( .A1(A[16]), .A2(B[16]), .ZN(n261) );
  NOR2_X1 U497 ( .A1(A[14]), .A2(B[14]), .ZN(n276) );
  NOR2_X1 U498 ( .A1(A[6]), .A2(B[6]), .ZN(n327) );
  NOR2_X1 U499 ( .A1(A[7]), .A2(B[7]), .ZN(n324) );
  NOR2_X1 U500 ( .A1(A[11]), .A2(B[11]), .ZN(n301) );
  NOR2_X1 U501 ( .A1(A[13]), .A2(B[13]), .ZN(n285) );
  NOR2_X1 U502 ( .A1(A[9]), .A2(B[9]), .ZN(n313) );
  NOR2_X1 U503 ( .A1(A[5]), .A2(B[5]), .ZN(n332) );
  NOR2_X1 U504 ( .A1(A[3]), .A2(B[3]), .ZN(n343) );
  NOR2_X1 U505 ( .A1(A[15]), .A2(B[15]), .ZN(n271) );
  NOR2_X1 U506 ( .A1(A[8]), .A2(B[8]), .ZN(n316) );
  NOR2_X1 U507 ( .A1(A[2]), .A2(B[2]), .ZN(n346) );
  NOR2_X1 U508 ( .A1(A[1]), .A2(B[1]), .ZN(n350) );
  AOI21_X1 U509 ( .B1(n263), .B2(n230), .A(n235), .ZN(n229) );
  INV_X1 U510 ( .A(n236), .ZN(n230) );
  INV_X2 U511 ( .A(n264), .ZN(n263) );
  INV_X1 U512 ( .A(n154), .ZN(n152) );
  INV_X1 U513 ( .A(n549), .ZN(n174) );
  INV_X1 U514 ( .A(n156), .ZN(n154) );
  INV_X1 U515 ( .A(n95), .ZN(n93) );
  NAND2_X1 U516 ( .A1(n154), .A2(n132), .ZN(n130) );
  OAI21_X1 U517 ( .B1(n318), .B2(n297), .A(n298), .ZN(n292) );
  AOI21_X1 U518 ( .B1(n263), .B2(n212), .A(n213), .ZN(n211) );
  INV_X1 U519 ( .A(n215), .ZN(n213) );
  INV_X1 U520 ( .A(n214), .ZN(n212) );
  AOI21_X1 U521 ( .B1(n263), .B2(n196), .A(n197), .ZN(n191) );
  AOI21_X1 U522 ( .B1(n263), .B2(n254), .A(n255), .ZN(n249) );
  AOI21_X1 U523 ( .B1(n155), .B2(n132), .A(n545), .ZN(n131) );
  NAND2_X1 U524 ( .A1(n230), .A2(n216), .ZN(n214) );
  INV_X1 U525 ( .A(n557), .ZN(n132) );
  INV_X1 U526 ( .A(n235), .ZN(n233) );
  INV_X1 U527 ( .A(n78), .ZN(n76) );
  INV_X1 U528 ( .A(n297), .ZN(n295) );
  INV_X1 U529 ( .A(n155), .ZN(n153) );
  NAND2_X1 U530 ( .A1(n283), .A2(n269), .ZN(n267) );
  NAND2_X1 U531 ( .A1(n549), .A2(n167), .ZN(n165) );
  AOI21_X1 U532 ( .B1(n339), .B2(n330), .A(n331), .ZN(n329) );
  AOI21_X1 U533 ( .B1(n235), .B2(n216), .A(n219), .ZN(n215) );
  INV_X1 U534 ( .A(n48), .ZN(n46) );
  NAND2_X1 U535 ( .A1(n154), .A2(n365), .ZN(n143) );
  OAI21_X1 U536 ( .B1(n318), .B2(n279), .A(n280), .ZN(n278) );
  NAND2_X1 U537 ( .A1(n295), .A2(n283), .ZN(n279) );
  AOI21_X1 U538 ( .B1(n296), .B2(n283), .A(n284), .ZN(n280) );
  OAI21_X1 U539 ( .B1(n318), .B2(n309), .A(n310), .ZN(n308) );
  INV_X1 U540 ( .A(n312), .ZN(n310) );
  INV_X1 U541 ( .A(n311), .ZN(n309) );
  INV_X1 U542 ( .A(n319), .ZN(n318) );
  NAND2_X1 U543 ( .A1(n254), .A2(n238), .ZN(n236) );
  NAND2_X1 U544 ( .A1(n121), .A2(n154), .ZN(n119) );
  INV_X1 U545 ( .A(n96), .ZN(n94) );
  NAND2_X1 U546 ( .A1(n218), .A2(n527), .ZN(n198) );
  INV_X1 U547 ( .A(n77), .ZN(n75) );
  INV_X1 U548 ( .A(n255), .ZN(n253) );
  INV_X1 U549 ( .A(n254), .ZN(n252) );
  INV_X1 U550 ( .A(n237), .ZN(n235) );
  NOR2_X1 U551 ( .A1(n557), .A2(n544), .ZN(n121) );
  INV_X1 U552 ( .A(n197), .ZN(n195) );
  INV_X1 U553 ( .A(n340), .ZN(n339) );
  NOR2_X1 U554 ( .A1(n78), .A2(n69), .ZN(n63) );
  OAI21_X1 U555 ( .B1(n75), .B2(n69), .A(n70), .ZN(n64) );
  NAND2_X1 U556 ( .A1(n311), .A2(n299), .ZN(n297) );
  INV_X1 U557 ( .A(n298), .ZN(n296) );
  INV_X1 U558 ( .A(n349), .ZN(n348) );
  INV_X1 U559 ( .A(n217), .ZN(n216) );
  INV_X1 U560 ( .A(n218), .ZN(n217) );
  NAND2_X1 U561 ( .A1(n67), .A2(n528), .ZN(n56) );
  AOI21_X1 U562 ( .B1(n263), .B2(n185), .A(n186), .ZN(n184) );
  NOR2_X1 U563 ( .A1(n247), .A2(n240), .ZN(n238) );
  OAI21_X1 U564 ( .B1(n237), .B2(n198), .A(n199), .ZN(n197) );
  INV_X1 U565 ( .A(n52), .ZN(n50) );
  AOI21_X1 U566 ( .B1(n341), .B2(n349), .A(n342), .ZN(n340) );
  NOR2_X1 U567 ( .A1(n346), .A2(n343), .ZN(n341) );
  OAI21_X1 U568 ( .B1(n343), .B2(n347), .A(n344), .ZN(n342) );
  INV_X1 U569 ( .A(n61), .ZN(n59) );
  OAI21_X1 U570 ( .B1(n313), .B2(n317), .A(n314), .ZN(n312) );
  OAI21_X1 U571 ( .B1(n332), .B2(n338), .A(n333), .ZN(n331) );
  OAI21_X1 U572 ( .B1(n285), .B2(n291), .A(n286), .ZN(n284) );
  OAI21_X1 U573 ( .B1(n350), .B2(n353), .A(n351), .ZN(n349) );
  NOR2_X1 U574 ( .A1(n94), .A2(n89), .ZN(n85) );
  OAI21_X1 U575 ( .B1(n95), .B2(n89), .A(n90), .ZN(n86) );
  INV_X1 U576 ( .A(n104), .ZN(n102) );
  OAI21_X1 U577 ( .B1(n220), .B2(n228), .A(n221), .ZN(n219) );
  NOR2_X1 U578 ( .A1(n327), .A2(n324), .ZN(n322) );
  AOI21_X1 U579 ( .B1(n299), .B2(n312), .A(n300), .ZN(n298) );
  OAI21_X1 U580 ( .B1(n301), .B2(n307), .A(n302), .ZN(n300) );
  NOR2_X1 U581 ( .A1(n276), .A2(n271), .ZN(n269) );
  NOR2_X1 U582 ( .A1(n306), .A2(n301), .ZN(n299) );
  NOR2_X1 U583 ( .A1(n337), .A2(n332), .ZN(n330) );
  AOI21_X1 U584 ( .B1(n238), .B2(n255), .A(n239), .ZN(n237) );
  NOR2_X1 U585 ( .A1(n316), .A2(n313), .ZN(n311) );
  NOR2_X1 U586 ( .A1(n290), .A2(n285), .ZN(n283) );
  OAI21_X1 U587 ( .B1(n340), .B2(n320), .A(n321), .ZN(n319) );
  AOI21_X1 U588 ( .B1(n322), .B2(n331), .A(n323), .ZN(n321) );
  NAND2_X1 U589 ( .A1(n330), .A2(n322), .ZN(n320) );
  OAI21_X1 U590 ( .B1(n324), .B2(n328), .A(n325), .ZN(n323) );
  AOI21_X1 U591 ( .B1(n263), .B2(n223), .A(n224), .ZN(n222) );
  OAI21_X1 U592 ( .B1(n233), .B2(n227), .A(n228), .ZN(n224) );
  NOR2_X1 U593 ( .A1(n236), .A2(n227), .ZN(n223) );
  AOI21_X1 U594 ( .B1(n263), .B2(n243), .A(n244), .ZN(n242) );
  NOR2_X1 U595 ( .A1(n252), .A2(n247), .ZN(n243) );
  OAI21_X1 U596 ( .B1(n253), .B2(n247), .A(n248), .ZN(n244) );
  AOI21_X1 U597 ( .B1(n278), .B2(n379), .A(n275), .ZN(n273) );
  INV_X1 U598 ( .A(n277), .ZN(n275) );
  AOI21_X1 U599 ( .B1(n292), .B2(n381), .A(n289), .ZN(n287) );
  INV_X1 U600 ( .A(n291), .ZN(n289) );
  AOI21_X1 U601 ( .B1(n308), .B2(n383), .A(n305), .ZN(n303) );
  INV_X1 U602 ( .A(n307), .ZN(n305) );
  AOI21_X1 U603 ( .B1(n263), .B2(n377), .A(n260), .ZN(n258) );
  INV_X1 U604 ( .A(n262), .ZN(n260) );
  INV_X1 U605 ( .A(n547), .ZN(n167) );
  INV_X1 U606 ( .A(n69), .ZN(n67) );
  INV_X1 U607 ( .A(n540), .ZN(n208) );
  INV_X1 U608 ( .A(n227), .ZN(n226) );
  AOI21_X1 U609 ( .B1(n263), .B2(n205), .A(n206), .ZN(n204) );
  NOR2_X1 U610 ( .A1(n214), .A2(n540), .ZN(n205) );
  OAI21_X1 U611 ( .B1(n318), .B2(n316), .A(n317), .ZN(n315) );
  AOI21_X1 U612 ( .B1(n269), .B2(n284), .A(n270), .ZN(n268) );
  OAI21_X1 U613 ( .B1(n271), .B2(n277), .A(n272), .ZN(n270) );
  INV_X1 U614 ( .A(n550), .ZN(n188) );
  AOI21_X1 U615 ( .B1(n155), .B2(n365), .A(n146), .ZN(n144) );
  INV_X1 U616 ( .A(n148), .ZN(n146) );
  AOI21_X1 U617 ( .B1(n541), .B2(n167), .A(n168), .ZN(n166) );
  INV_X1 U618 ( .A(n170), .ZN(n168) );
  INV_X1 U619 ( .A(n103), .ZN(n361) );
  INV_X1 U620 ( .A(n220), .ZN(n372) );
  INV_X1 U621 ( .A(n537), .ZN(n366) );
  INV_X1 U622 ( .A(n536), .ZN(n362) );
  INV_X1 U623 ( .A(n70), .ZN(n68) );
  INV_X1 U624 ( .A(n247), .ZN(n246) );
  INV_X1 U625 ( .A(n89), .ZN(n88) );
  INV_X1 U626 ( .A(n82), .ZN(n358) );
  INV_X1 U627 ( .A(n98), .ZN(n360) );
  INV_X1 U628 ( .A(n327), .ZN(n387) );
  INV_X1 U629 ( .A(n316), .ZN(n385) );
  INV_X1 U630 ( .A(n346), .ZN(n391) );
  INV_X1 U631 ( .A(n271), .ZN(n378) );
  INV_X1 U632 ( .A(n301), .ZN(n382) );
  INV_X1 U633 ( .A(n285), .ZN(n380) );
  INV_X1 U634 ( .A(n313), .ZN(n384) );
  INV_X1 U635 ( .A(n276), .ZN(n379) );
  INV_X1 U636 ( .A(n290), .ZN(n381) );
  INV_X1 U637 ( .A(n306), .ZN(n383) );
  INV_X1 U638 ( .A(n337), .ZN(n389) );
  NAND2_X1 U639 ( .A1(n386), .A2(n325), .ZN(n34) );
  INV_X1 U640 ( .A(n324), .ZN(n386) );
  NAND2_X1 U641 ( .A1(n390), .A2(n344), .ZN(n38) );
  INV_X1 U642 ( .A(n343), .ZN(n390) );
  INV_X1 U643 ( .A(n261), .ZN(n377) );
  INV_X1 U644 ( .A(n532), .ZN(n365) );
  NAND2_X1 U645 ( .A1(n388), .A2(n333), .ZN(n36) );
  INV_X1 U646 ( .A(n332), .ZN(n388) );
  INV_X1 U647 ( .A(n240), .ZN(n374) );
  INV_X1 U648 ( .A(n350), .ZN(n392) );
  INV_X1 U649 ( .A(n338), .ZN(n336) );
  INV_X1 U650 ( .A(n544), .ZN(n124) );
  INV_X1 U651 ( .A(n256), .ZN(n376) );
  NOR2_X1 U652 ( .A1(A[28]), .A2(B[28]), .ZN(n147) );
  NOR2_X1 U653 ( .A1(B[26]), .A2(A[26]), .ZN(n169) );
  NOR2_X1 U654 ( .A1(B[30]), .A2(A[30]), .ZN(n125) );
  NOR2_X1 U655 ( .A1(A[17]), .A2(B[17]), .ZN(n256) );
  NOR2_X1 U656 ( .A1(B[25]), .A2(A[25]), .ZN(n182) );
  NOR2_X1 U657 ( .A1(A[19]), .A2(B[19]), .ZN(n240) );
  NAND2_X1 U658 ( .A1(A[32]), .A2(B[32]), .ZN(n104) );
  NAND2_X1 U659 ( .A1(B[26]), .A2(A[26]), .ZN(n170) );
  NAND2_X1 U660 ( .A1(A[34]), .A2(B[34]), .ZN(n90) );
  NAND2_X1 U661 ( .A1(n559), .A2(n183), .ZN(n16) );
  NAND2_X1 U662 ( .A1(n362), .A2(n115), .ZN(n10) );
  NAND2_X1 U663 ( .A1(n364), .A2(n139), .ZN(n12) );
  NAND2_X1 U664 ( .A1(n124), .A2(n539), .ZN(n11) );
  NAND2_X1 U665 ( .A1(A[37]), .A2(B[37]), .ZN(n61) );
  NAND2_X1 U666 ( .A1(n361), .A2(n104), .ZN(n9) );
  NAND2_X1 U667 ( .A1(A[6]), .A2(B[6]), .ZN(n328) );
  XOR2_X1 U668 ( .A(n318), .B(n33), .Z(SUM[8]) );
  NAND2_X1 U669 ( .A1(n385), .A2(n317), .ZN(n33) );
  XOR2_X1 U670 ( .A(n329), .B(n35), .Z(SUM[6]) );
  NAND2_X1 U671 ( .A1(n387), .A2(n328), .ZN(n35) );
  XOR2_X1 U672 ( .A(n171), .B(n15), .Z(SUM[26]) );
  NAND2_X1 U673 ( .A1(n167), .A2(n170), .ZN(n15) );
  XNOR2_X1 U674 ( .A(n263), .B(n25), .ZN(SUM[16]) );
  NAND2_X1 U675 ( .A1(n377), .A2(n262), .ZN(n25) );
  NAND2_X1 U676 ( .A1(A[8]), .A2(B[8]), .ZN(n317) );
  NAND2_X1 U677 ( .A1(A[14]), .A2(B[14]), .ZN(n277) );
  NAND2_X1 U678 ( .A1(A[12]), .A2(B[12]), .ZN(n291) );
  NAND2_X1 U679 ( .A1(A[10]), .A2(B[10]), .ZN(n307) );
  NAND2_X1 U680 ( .A1(A[4]), .A2(B[4]), .ZN(n338) );
  NAND2_X1 U681 ( .A1(A[2]), .A2(B[2]), .ZN(n347) );
  XOR2_X1 U682 ( .A(n222), .B(n20), .Z(SUM[21]) );
  NAND2_X1 U683 ( .A1(n372), .A2(n221), .ZN(n20) );
  XOR2_X1 U684 ( .A(n258), .B(n24), .Z(SUM[17]) );
  NAND2_X1 U685 ( .A1(n376), .A2(n257), .ZN(n24) );
  XOR2_X1 U686 ( .A(n249), .B(n23), .Z(SUM[18]) );
  NAND2_X1 U687 ( .A1(n246), .A2(n248), .ZN(n23) );
  XOR2_X1 U688 ( .A(n242), .B(n22), .Z(SUM[19]) );
  NAND2_X1 U689 ( .A1(n374), .A2(n241), .ZN(n22) );
  XOR2_X1 U690 ( .A(n229), .B(n21), .Z(SUM[20]) );
  NAND2_X1 U691 ( .A1(n226), .A2(n228), .ZN(n21) );
  XOR2_X1 U692 ( .A(n211), .B(n19), .Z(SUM[22]) );
  NAND2_X1 U693 ( .A1(n208), .A2(n210), .ZN(n19) );
  XOR2_X1 U694 ( .A(n191), .B(n17), .Z(SUM[24]) );
  NAND2_X1 U695 ( .A1(n188), .A2(n190), .ZN(n17) );
  XOR2_X1 U696 ( .A(n149), .B(n13), .Z(SUM[28]) );
  NAND2_X1 U697 ( .A1(n365), .A2(n520), .ZN(n13) );
  NAND2_X1 U698 ( .A1(n523), .A2(n203), .ZN(n18) );
  XOR2_X1 U699 ( .A(n162), .B(n14), .Z(SUM[27]) );
  NAND2_X1 U700 ( .A1(n366), .A2(n521), .ZN(n14) );
  XOR2_X1 U701 ( .A(n273), .B(n26), .Z(SUM[15]) );
  NAND2_X1 U702 ( .A1(n378), .A2(n272), .ZN(n26) );
  XNOR2_X1 U703 ( .A(n292), .B(n29), .ZN(SUM[12]) );
  NAND2_X1 U704 ( .A1(n381), .A2(n291), .ZN(n29) );
  XNOR2_X1 U705 ( .A(n308), .B(n31), .ZN(SUM[10]) );
  NAND2_X1 U706 ( .A1(n383), .A2(n307), .ZN(n31) );
  XOR2_X1 U707 ( .A(n40), .B(n353), .Z(SUM[1]) );
  NAND2_X1 U708 ( .A1(n392), .A2(n351), .ZN(n40) );
  XOR2_X1 U709 ( .A(n348), .B(n39), .Z(SUM[2]) );
  NAND2_X1 U710 ( .A1(n391), .A2(n347), .ZN(n39) );
  XNOR2_X1 U711 ( .A(n345), .B(n38), .ZN(SUM[3]) );
  OAI21_X1 U712 ( .B1(n348), .B2(n346), .A(n347), .ZN(n345) );
  XNOR2_X1 U713 ( .A(n339), .B(n37), .ZN(SUM[4]) );
  NAND2_X1 U714 ( .A1(n389), .A2(n338), .ZN(n37) );
  XNOR2_X1 U715 ( .A(n315), .B(n32), .ZN(SUM[9]) );
  NAND2_X1 U716 ( .A1(n384), .A2(n314), .ZN(n32) );
  XNOR2_X1 U717 ( .A(n326), .B(n34), .ZN(SUM[7]) );
  OAI21_X1 U718 ( .B1(n329), .B2(n327), .A(n328), .ZN(n326) );
  XOR2_X1 U719 ( .A(n334), .B(n36), .Z(SUM[5]) );
  AOI21_X1 U720 ( .B1(n339), .B2(n389), .A(n336), .ZN(n334) );
  AND2_X1 U721 ( .A1(n562), .A2(n353), .ZN(SUM[0]) );
  NAND2_X1 U722 ( .A1(A[7]), .A2(B[7]), .ZN(n325) );
  NAND2_X1 U723 ( .A1(A[0]), .A2(B[0]), .ZN(n353) );
  NAND2_X1 U724 ( .A1(A[16]), .A2(B[16]), .ZN(n262) );
  NAND2_X1 U725 ( .A1(A[18]), .A2(B[18]), .ZN(n248) );
  NAND2_X1 U726 ( .A1(A[15]), .A2(B[15]), .ZN(n272) );
  XNOR2_X1 U727 ( .A(n278), .B(n27), .ZN(SUM[14]) );
  NAND2_X1 U728 ( .A1(n379), .A2(n277), .ZN(n27) );
  NAND2_X1 U729 ( .A1(A[19]), .A2(B[19]), .ZN(n241) );
  NAND2_X1 U730 ( .A1(A[38]), .A2(B[38]), .ZN(n52) );
  NAND2_X1 U731 ( .A1(A[11]), .A2(B[11]), .ZN(n302) );
  NAND2_X1 U732 ( .A1(A[13]), .A2(B[13]), .ZN(n286) );
  NAND2_X1 U733 ( .A1(A[9]), .A2(B[9]), .ZN(n314) );
  NAND2_X1 U734 ( .A1(A[1]), .A2(B[1]), .ZN(n351) );
  NAND2_X1 U735 ( .A1(A[5]), .A2(B[5]), .ZN(n333) );
  NAND2_X1 U736 ( .A1(A[3]), .A2(B[3]), .ZN(n344) );
  NAND2_X1 U737 ( .A1(A[39]), .A2(B[39]), .ZN(n43) );
  NAND2_X1 U738 ( .A1(B[29]), .A2(A[29]), .ZN(n139) );
  XOR2_X1 U739 ( .A(n287), .B(n28), .Z(SUM[13]) );
  NAND2_X1 U740 ( .A1(n380), .A2(n286), .ZN(n28) );
  XOR2_X1 U741 ( .A(n303), .B(n30), .Z(SUM[11]) );
  NAND2_X1 U742 ( .A1(n382), .A2(n302), .ZN(n30) );
  OR2_X1 U743 ( .A1(A[39]), .A2(B[39]), .ZN(n561) );
  OR2_X1 U744 ( .A1(A[0]), .A2(B[0]), .ZN(n562) );
  NAND2_X1 U745 ( .A1(B[30]), .A2(A[30]), .ZN(n126) );
  INV_X1 U746 ( .A(n541), .ZN(n179) );
  INV_X1 U747 ( .A(n558), .ZN(n364) );
  NOR2_X1 U748 ( .A1(B[29]), .A2(A[29]), .ZN(n138) );
  NOR2_X1 U749 ( .A1(n297), .A2(n267), .ZN(n265) );
  NAND2_X1 U750 ( .A1(A[23]), .A2(B[23]), .ZN(n203) );
  INV_X1 U751 ( .A(n196), .ZN(n194) );
  XOR2_X1 U752 ( .A(n127), .B(n11), .Z(SUM[30]) );
  OAI21_X1 U753 ( .B1(n135), .B2(n544), .A(n539), .ZN(n122) );
  NOR2_X1 U754 ( .A1(n261), .A2(n256), .ZN(n254) );
  OAI21_X1 U755 ( .B1(n256), .B2(n262), .A(n257), .ZN(n255) );
  NAND2_X1 U756 ( .A1(A[17]), .A2(B[17]), .ZN(n257) );
  AOI21_X1 U757 ( .B1(n319), .B2(n265), .A(n266), .ZN(n264) );
  OAI21_X1 U758 ( .B1(n298), .B2(n267), .A(n268), .ZN(n266) );
  NOR2_X1 U759 ( .A1(B[31]), .A2(A[31]), .ZN(n114) );
  INV_X1 U760 ( .A(n545), .ZN(n135) );
  INV_X1 U761 ( .A(n97), .ZN(n95) );
  OAI21_X1 U762 ( .B1(n98), .B2(n104), .A(n99), .ZN(n97) );
  XOR2_X1 U763 ( .A(n204), .B(n18), .Z(SUM[23]) );
  OAI21_X1 U764 ( .B1(n215), .B2(n540), .A(n210), .ZN(n206) );
  OAI21_X1 U765 ( .B1(n240), .B2(n248), .A(n241), .ZN(n239) );
  AOI21_X1 U766 ( .B1(n263), .B2(n117), .A(n118), .ZN(n116) );
  NAND2_X1 U767 ( .A1(A[36]), .A2(B[36]), .ZN(n70) );
  NOR2_X1 U768 ( .A1(A[36]), .A2(B[36]), .ZN(n69) );
  INV_X1 U769 ( .A(n79), .ZN(n77) );
  NOR2_X1 U770 ( .A1(n103), .A2(n98), .ZN(n96) );
  AOI21_X1 U771 ( .B1(n263), .B2(n163), .A(n164), .ZN(n162) );
  AOI21_X1 U772 ( .B1(n527), .B2(n219), .A(n201), .ZN(n199) );
  NAND2_X1 U773 ( .A1(A[20]), .A2(B[20]), .ZN(n228) );
  INV_X1 U774 ( .A(n546), .ZN(n155) );
  AOI21_X1 U775 ( .B1(n80), .B2(n97), .A(n81), .ZN(n79) );
  AOI21_X1 U776 ( .B1(n528), .B2(n68), .A(n59), .ZN(n57) );
  AOI21_X1 U777 ( .B1(n263), .B2(n172), .A(n173), .ZN(n171) );
  NOR2_X1 U778 ( .A1(B[22]), .A2(A[22]), .ZN(n209) );
  AOI21_X1 U779 ( .B1(n263), .B2(n141), .A(n142), .ZN(n140) );
  NAND2_X1 U780 ( .A1(n112), .A2(n136), .ZN(n110) );
  NOR2_X1 U781 ( .A1(n147), .A2(n138), .ZN(n136) );
  NAND2_X1 U782 ( .A1(B[31]), .A2(A[31]), .ZN(n115) );
  AOI21_X1 U783 ( .B1(n263), .B2(n150), .A(n151), .ZN(n149) );
  NAND2_X1 U784 ( .A1(B[25]), .A2(A[25]), .ZN(n183) );
  NOR2_X1 U785 ( .A1(n78), .A2(n56), .ZN(n54) );
  NOR2_X1 U786 ( .A1(n89), .A2(n82), .ZN(n80) );
  AOI21_X1 U787 ( .B1(n108), .B2(n197), .A(n109), .ZN(n107) );
  NOR2_X1 U788 ( .A1(n194), .A2(n130), .ZN(n128) );
  NOR2_X1 U789 ( .A1(n194), .A2(n550), .ZN(n185) );
  NOR2_X1 U790 ( .A1(n194), .A2(n143), .ZN(n141) );
  NOR2_X1 U791 ( .A1(n194), .A2(n119), .ZN(n117) );
  NOR2_X1 U792 ( .A1(n194), .A2(n174), .ZN(n172) );
  NOR2_X1 U793 ( .A1(n194), .A2(n165), .ZN(n163) );
  NOR2_X1 U794 ( .A1(n194), .A2(n152), .ZN(n150) );
  NOR2_X1 U795 ( .A1(n227), .A2(n220), .ZN(n218) );
  NAND2_X1 U796 ( .A1(A[21]), .A2(B[21]), .ZN(n221) );
  NOR2_X1 U797 ( .A1(A[21]), .A2(B[21]), .ZN(n220) );
  AOI21_X1 U798 ( .B1(n263), .B2(n128), .A(n129), .ZN(n127) );
  NAND2_X1 U799 ( .A1(B[28]), .A2(A[28]), .ZN(n148) );
  XOR2_X1 U800 ( .A(n184), .B(n16), .Z(SUM[25]) );
  OAI21_X1 U801 ( .B1(n195), .B2(n550), .A(n190), .ZN(n186) );
  OAI21_X1 U802 ( .B1(n195), .B2(n143), .A(n144), .ZN(n142) );
  OAI21_X1 U803 ( .B1(n195), .B2(n119), .A(n120), .ZN(n118) );
  OAI21_X1 U804 ( .B1(n195), .B2(n174), .A(n179), .ZN(n173) );
  OAI21_X1 U805 ( .B1(n195), .B2(n165), .A(n166), .ZN(n164) );
  OAI21_X1 U806 ( .B1(n195), .B2(n152), .A(n153), .ZN(n151) );
  OAI21_X1 U807 ( .B1(n195), .B2(n130), .A(n131), .ZN(n129) );
  OAI21_X1 U808 ( .B1(n526), .B2(n210), .A(n203), .ZN(n201) );
  NOR2_X1 U809 ( .A1(n156), .A2(n110), .ZN(n108) );
  NOR2_X1 U810 ( .A1(n189), .A2(n182), .ZN(n180) );
  NAND2_X1 U811 ( .A1(B[24]), .A2(A[24]), .ZN(n190) );
  NOR2_X1 U812 ( .A1(A[24]), .A2(B[24]), .ZN(n189) );
  NAND2_X1 U813 ( .A1(n96), .A2(n80), .ZN(n78) );
  NOR2_X1 U814 ( .A1(A[32]), .A2(B[32]), .ZN(n103) );
  AOI21_X1 U815 ( .B1(n55), .B2(n529), .A(n50), .ZN(n48) );
  OAI21_X1 U816 ( .B1(n82), .B2(n90), .A(n83), .ZN(n81) );
  NAND2_X1 U817 ( .A1(A[35]), .A2(B[35]), .ZN(n83) );
  XOR2_X1 U818 ( .A(n140), .B(n12), .Z(SUM[29]) );
  AOI21_X1 U819 ( .B1(n181), .B2(n534), .A(n159), .ZN(n157) );
  NAND2_X1 U820 ( .A1(n180), .A2(n534), .ZN(n156) );
  OAI21_X1 U821 ( .B1(n160), .B2(n170), .A(n161), .ZN(n159) );
  NAND2_X1 U822 ( .A1(B[27]), .A2(A[27]), .ZN(n161) );
  NOR2_X1 U823 ( .A1(B[27]), .A2(A[27]), .ZN(n160) );
  OAI21_X1 U824 ( .B1(n79), .B2(n56), .A(n57), .ZN(n55) );
  NAND2_X1 U825 ( .A1(A[33]), .A2(B[33]), .ZN(n99) );
  XOR2_X1 U826 ( .A(n116), .B(n10), .Z(SUM[31]) );
  AOI21_X1 U827 ( .B1(n121), .B2(n155), .A(n122), .ZN(n120) );
  OAI21_X1 U828 ( .B1(n264), .B2(n106), .A(n107), .ZN(n105) );
  OAI21_X1 U829 ( .B1(n157), .B2(n110), .A(n111), .ZN(n109) );
  OAI21_X1 U830 ( .B1(n522), .B2(n190), .A(n183), .ZN(n181) );
  OAI21_X1 U831 ( .B1(n543), .B2(n148), .A(n139), .ZN(n137) );
  XNOR2_X1 U832 ( .A(n552), .B(n9), .ZN(SUM[32]) );
  AOI21_X1 U833 ( .B1(n552), .B2(n361), .A(n102), .ZN(n100) );
  AOI21_X1 U834 ( .B1(n552), .B2(n76), .A(n77), .ZN(n71) );
  AOI21_X1 U835 ( .B1(n552), .B2(n96), .A(n93), .ZN(n91) );
  AOI21_X1 U836 ( .B1(n1), .B2(n530), .A(n46), .ZN(n44) );
  AOI21_X1 U837 ( .B1(n1), .B2(n63), .A(n64), .ZN(n62) );
  AOI21_X1 U838 ( .B1(n552), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U839 ( .B1(n1), .B2(n54), .A(n55), .ZN(n53) );
  AOI21_X1 U840 ( .B1(n542), .B2(n137), .A(n113), .ZN(n111) );
  NAND2_X1 U841 ( .A1(n531), .A2(n196), .ZN(n106) );
  OAI21_X1 U842 ( .B1(n126), .B2(n114), .A(n115), .ZN(n113) );
  NOR2_X1 U843 ( .A1(n548), .A2(n125), .ZN(n112) );
endmodule


module datapath ( clk, data_in, addr_x, wr_en_x, addr_a1, addr_a2, addr_a3, 
        addr_a4, addr_a5, addr_a6, addr_a7, addr_a8, wr_en_a1, wr_en_a2, 
        wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6, wr_en_a7, wr_en_a8, addr_y, 
        wr_en_y, clear_acc, clc, clc1, data_out );
  input [19:0] data_in;
  input [2:0] addr_x;
  input [2:0] addr_a1;
  input [2:0] addr_a2;
  input [2:0] addr_a3;
  input [2:0] addr_a4;
  input [2:0] addr_a5;
  input [2:0] addr_a6;
  input [2:0] addr_a7;
  input [2:0] addr_a8;
  input [2:0] addr_y;
  output [39:0] data_out;
  input clk, wr_en_x, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5,
         wr_en_a6, wr_en_a7, wr_en_a8, wr_en_y, clear_acc, clc, clc1;
  wire   n27, n28, n29, n30, n31, n32, n33, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n267, n268, n269, n270,
         n271, n272, n273, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n338,
         n339, n340, n341, n343, n344, n345, n349, n350, n351, n352, n355,
         n356, n359, n360, n363, n364, n367, n368, n371, n372, n375, n376,
         n379, n380, n383, n384, n387, n388, n391, n392, n395, n396, n399,
         n400, n403, n404, n407, n408, n411, n412, n415, n416, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n506, n507, n508, n509, n510, n511, n512,
         n513, n515, n516, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, \mul_out1[9] ,
         \mul_out1[8] , \mul_out1[7] , \mul_out1[6] , \mul_out1[5] ,
         \mul_out1[4] , \mul_out1[3] , \mul_out1[39] , \mul_out1[38] ,
         \mul_out1[37] , \mul_out1[36] , \mul_out1[35] , \mul_out1[34] ,
         \mul_out1[33] , \mul_out1[32] , \mul_out1[31] , \mul_out1[30] ,
         \mul_out1[2] , \mul_out1[29] , \mul_out1[28] , \mul_out1[27] ,
         \mul_out1[26] , \mul_out1[25] , \mul_out1[24] , \mul_out1[23] ,
         \mul_out1[22] , \mul_out1[21] , \mul_out1[20] , \mul_out1[1] ,
         \mul_out1[19] , \mul_out1[18] , \mul_out1[17] , \mul_out1[16] ,
         \mul_out1[15] , \mul_out1[14] , \mul_out1[13] , \mul_out1[12] ,
         \mul_out1[11] , \mul_out1[10] , \mul_out1[0] , \mul_out2[9] ,
         \mul_out2[8] , \mul_out2[7] , \mul_out2[6] , \mul_out2[5] ,
         \mul_out2[4] , \mul_out2[3] , \mul_out2[39] , \mul_out2[38] ,
         \mul_out2[37] , \mul_out2[36] , \mul_out2[35] , \mul_out2[34] ,
         \mul_out2[33] , \mul_out2[32] , \mul_out2[31] , \mul_out2[30] ,
         \mul_out2[2] , \mul_out2[29] , \mul_out2[28] , \mul_out2[27] ,
         \mul_out2[26] , \mul_out2[25] , \mul_out2[24] , \mul_out2[23] ,
         \mul_out2[22] , \mul_out2[21] , \mul_out2[20] , \mul_out2[1] ,
         \mul_out2[19] , \mul_out2[18] , \mul_out2[17] , \mul_out2[16] ,
         \mul_out2[15] , \mul_out2[14] , \mul_out2[13] , \mul_out2[12] ,
         \mul_out2[11] , \mul_out2[10] , \mul_out2[0] , \mul_out3[9] ,
         \mul_out3[8] , \mul_out3[7] , \mul_out3[6] , \mul_out3[5] ,
         \mul_out3[4] , \mul_out3[3] , \mul_out3[39] , \mul_out3[38] ,
         \mul_out3[37] , \mul_out3[36] , \mul_out3[35] , \mul_out3[34] ,
         \mul_out3[33] , \mul_out3[32] , \mul_out3[31] , \mul_out3[30] ,
         \mul_out3[2] , \mul_out3[29] , \mul_out3[28] , \mul_out3[27] ,
         \mul_out3[26] , \mul_out3[25] , \mul_out3[24] , \mul_out3[23] ,
         \mul_out3[22] , \mul_out3[21] , \mul_out3[20] , \mul_out3[1] ,
         \mul_out3[19] , \mul_out3[18] , \mul_out3[17] , \mul_out3[16] ,
         \mul_out3[15] , \mul_out3[14] , \mul_out3[13] , \mul_out3[12] ,
         \mul_out3[11] , \mul_out3[10] , \mul_out3[0] , \mul_out4[9] ,
         \mul_out4[8] , \mul_out4[7] , \mul_out4[6] , \mul_out4[5] ,
         \mul_out4[4] , \mul_out4[3] , \mul_out4[39] , \mul_out4[38] ,
         \mul_out4[37] , \mul_out4[36] , \mul_out4[35] , \mul_out4[34] ,
         \mul_out4[33] , \mul_out4[32] , \mul_out4[31] , \mul_out4[30] ,
         \mul_out4[2] , \mul_out4[29] , \mul_out4[28] , \mul_out4[27] ,
         \mul_out4[26] , \mul_out4[25] , \mul_out4[24] , \mul_out4[23] ,
         \mul_out4[22] , \mul_out4[21] , \mul_out4[20] , \mul_out4[1] ,
         \mul_out4[19] , \mul_out4[18] , \mul_out4[17] , \mul_out4[16] ,
         \mul_out4[15] , \mul_out4[14] , \mul_out4[13] , \mul_out4[12] ,
         \mul_out4[11] , \mul_out4[10] , \mul_out4[0] , \mul_out5[9] ,
         \mul_out5[8] , \mul_out5[7] , \mul_out5[6] , \mul_out5[5] ,
         \mul_out5[4] , \mul_out5[3] , \mul_out5[39] , \mul_out5[38] ,
         \mul_out5[37] , \mul_out5[36] , \mul_out5[35] , \mul_out5[34] ,
         \mul_out5[33] , \mul_out5[32] , \mul_out5[31] , \mul_out5[30] ,
         \mul_out5[2] , \mul_out5[29] , \mul_out5[28] , \mul_out5[27] ,
         \mul_out5[26] , \mul_out5[25] , \mul_out5[24] , \mul_out5[23] ,
         \mul_out5[22] , \mul_out5[21] , \mul_out5[20] , \mul_out5[1] ,
         \mul_out5[19] , \mul_out5[18] , \mul_out5[17] , \mul_out5[16] ,
         \mul_out5[15] , \mul_out5[14] , \mul_out5[13] , \mul_out5[12] ,
         \mul_out5[11] , \mul_out5[10] , \mul_out5[0] , \mul_out6[9] ,
         \mul_out6[8] , \mul_out6[7] , \mul_out6[6] , \mul_out6[5] ,
         \mul_out6[4] , \mul_out6[3] , \mul_out6[39] , \mul_out6[38] ,
         \mul_out6[37] , \mul_out6[36] , \mul_out6[35] , \mul_out6[34] ,
         \mul_out6[33] , \mul_out6[32] , \mul_out6[31] , \mul_out6[30] ,
         \mul_out6[2] , \mul_out6[29] , \mul_out6[28] , \mul_out6[27] ,
         \mul_out6[26] , \mul_out6[25] , \mul_out6[24] , \mul_out6[23] ,
         \mul_out6[22] , \mul_out6[21] , \mul_out6[20] , \mul_out6[1] ,
         \mul_out6[19] , \mul_out6[18] , \mul_out6[17] , \mul_out6[16] ,
         \mul_out6[15] , \mul_out6[14] , \mul_out6[13] , \mul_out6[12] ,
         \mul_out6[11] , \mul_out6[10] , \mul_out6[0] , \mul_out7[9] ,
         \mul_out7[8] , \mul_out7[7] , \mul_out7[6] , \mul_out7[5] ,
         \mul_out7[4] , \mul_out7[3] , \mul_out7[39] , \mul_out7[38] ,
         \mul_out7[37] , \mul_out7[36] , \mul_out7[35] , \mul_out7[34] ,
         \mul_out7[33] , \mul_out7[32] , \mul_out7[31] , \mul_out7[30] ,
         \mul_out7[2] , \mul_out7[29] , \mul_out7[28] , \mul_out7[27] ,
         \mul_out7[26] , \mul_out7[25] , \mul_out7[24] , \mul_out7[23] ,
         \mul_out7[22] , \mul_out7[21] , \mul_out7[20] , \mul_out7[1] ,
         \mul_out7[19] , \mul_out7[18] , \mul_out7[17] , \mul_out7[16] ,
         \mul_out7[15] , \mul_out7[14] , \mul_out7[13] , \mul_out7[12] ,
         \mul_out7[11] , \mul_out7[10] , \mul_out7[0] , \mul_out8[9] ,
         \mul_out8[8] , \mul_out8[7] , \mul_out8[6] , \mul_out8[5] ,
         \mul_out8[4] , \mul_out8[3] , \mul_out8[39] , \mul_out8[38] ,
         \mul_out8[37] , \mul_out8[36] , \mul_out8[35] , \mul_out8[34] ,
         \mul_out8[33] , \mul_out8[32] , \mul_out8[31] , \mul_out8[30] ,
         \mul_out8[2] , \mul_out8[29] , \mul_out8[28] , \mul_out8[27] ,
         \mul_out8[26] , \mul_out8[25] , \mul_out8[24] , \mul_out8[23] ,
         \mul_out8[22] , \mul_out8[21] , \mul_out8[20] , \mul_out8[1] ,
         \mul_out8[19] , \mul_out8[18] , \mul_out8[17] , \mul_out8[16] ,
         \mul_out8[15] , \mul_out8[14] , \mul_out8[13] , \mul_out8[12] ,
         \mul_out8[11] , \mul_out8[10] , \mul_out8[0] , n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n342, n346, n347, n348, n353, n354, n357, n358,
         n361, n362, n365, n366, n369, n370, n373, n374, n377, n378, n381,
         n382, n385, n386, n389, n390, n393, n394, n397, n398, n401, n402,
         n405, n406, n409, n410, n413, n414, n417, n418, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n514, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361;
  wire   [19:0] data_out_x;
  wire   [19:0] data_out_a1;
  wire   [19:0] data_out_a2;
  wire   [19:0] data_out_a3;
  wire   [19:0] data_out_a4;
  wire   [19:0] data_out_a5;
  wire   [19:0] data_out_a6;
  wire   [19:0] data_out_a7;
  wire   [19:0] data_out_a8;
  wire   [39:0] f;
  wire   [39:0] f1;
  wire   [39:0] f2;
  wire   [39:0] f3;
  wire   [39:0] f4;
  wire   [39:0] f5;
  wire   [39:0] f6;
  wire   [39:0] f7;
  wire   [39:0] f8;
  wire   [39:0] add_r1;
  wire   [39:0] add_r2;
  wire   [39:0] add_r3;
  wire   [39:0] add_r4;
  wire   [39:0] add_r5;
  wire   [39:0] add_r6;
  wire   [39:0] add_r7;
  wire   [39:0] add_r8;

  DFF_X1 \f1_reg[36]  ( .D(n1195), .CK(clk), .Q(f1[36]), .QN(n1334) );
  DFF_X1 \f1_reg[34]  ( .D(n1193), .CK(clk), .Q(f1[34]), .QN(n1324) );
  DFF_X1 \f1_reg[33]  ( .D(n1192), .CK(clk), .Q(f1[33]), .QN(n1319) );
  DFF_X1 \f1_reg[28]  ( .D(n1187), .CK(clk), .Q(f1[28]), .QN(n1295) );
  DFF_X1 \f1_reg[27]  ( .D(n1186), .CK(clk), .Q(f1[27]), .QN(n1290) );
  DFF_X1 \f1_reg[26]  ( .D(n1185), .CK(clk), .Q(f1[26]), .QN(n1285) );
  DFF_X1 \f1_reg[25]  ( .D(n1184), .CK(clk), .Q(f1[25]), .QN(n1280) );
  DFF_X1 \f1_reg[24]  ( .D(n1183), .CK(clk), .Q(f1[24]), .QN(n1275) );
  DFF_X1 \f2_reg[39]  ( .D(n1158), .CK(clk), .Q(n766), .QN(n49) );
  DFF_X1 \f2_reg[35]  ( .D(n1154), .CK(clk), .Q(n774), .QN(n53) );
  DFF_X1 \f2_reg[34]  ( .D(n1153), .CK(clk), .Q(n776), .QN(n54) );
  DFF_X1 \f2_reg[30]  ( .D(n1149), .CK(clk), .Q(n784), .QN(n58) );
  DFF_X1 \f3_reg[39]  ( .D(n1118), .CK(clk), .Q(n642), .QN(n89) );
  DFF_X1 \f3_reg[37]  ( .D(n1116), .CK(clk), .Q(n646), .QN(n91) );
  DFF_X1 \f3_reg[35]  ( .D(n1114), .CK(clk), .Q(n649), .QN(n93) );
  DFF_X1 \f4_reg[32]  ( .D(n1071), .CK(clk), .Q(f4[32]), .QN(n136) );
  DFF_X1 \f4_reg[31]  ( .D(n1070), .CK(clk), .Q(f4[31]), .QN(n137) );
  DFF_X1 \f4_reg[30]  ( .D(n1069), .CK(clk), .Q(f4[30]), .QN(n138) );
  DFF_X1 \f4_reg[29]  ( .D(n1068), .CK(clk), .Q(f4[29]), .QN(n139) );
  DFF_X1 \f4_reg[28]  ( .D(n1067), .CK(clk), .Q(f4[28]), .QN(n140) );
  DFF_X1 \f5_reg[30]  ( .D(n1029), .CK(clk), .Q(n720), .QN(n178) );
  DFF_X1 \f5_reg[29]  ( .D(n1028), .CK(clk), .Q(n722), .QN(n179) );
  DFF_X1 \f6_reg[39]  ( .D(n998), .CK(clk), .Q(n1355) );
  DFF_X1 \f6_reg[37]  ( .D(n996), .CK(clk), .Q(n1342) );
  DFF_X1 \f6_reg[36]  ( .D(n995), .CK(clk), .Q(n1337) );
  DFF_X1 \f6_reg[35]  ( .D(n994), .CK(clk), .Q(n1332) );
  DFF_X1 \f6_reg[34]  ( .D(n993), .CK(clk), .Q(n1327) );
  DFF_X1 \f6_reg[33]  ( .D(n992), .CK(clk), .Q(n1322) );
  DFF_X1 \f6_reg[32]  ( .D(n991), .CK(clk), .Q(n1317) );
  DFF_X1 \f6_reg[30]  ( .D(n989), .CK(clk), .Q(n1308) );
  DFF_X1 \f6_reg[24]  ( .D(n983), .CK(clk), .Q(n1278) );
  DFF_X1 \f6_reg[23]  ( .D(n982), .CK(clk), .Q(n1273) );
  DFF_X1 \f6_reg[22]  ( .D(n981), .CK(clk), .Q(n1268) );
  DFF_X1 \f7_reg[37]  ( .D(n956), .CK(clk), .Q(n1341) );
  DFF_X1 \f7_reg[34]  ( .D(n953), .CK(clk), .Q(n1326) );
  DFF_X1 \f7_reg[33]  ( .D(n952), .CK(clk), .Q(n1321) );
  DFF_X1 \f7_reg[31]  ( .D(n950), .CK(clk), .Q(n1312) );
  DFF_X1 \f7_reg[30]  ( .D(n949), .CK(clk), .Q(n1307) );
  DFF_X1 \f7_reg[29]  ( .D(n948), .CK(clk), .Q(n1302) );
  DFF_X1 \f7_reg[28]  ( .D(n947), .CK(clk), .Q(n1297) );
  DFF_X1 \f7_reg[27]  ( .D(n946), .CK(clk), .Q(n1292) );
  DFF_X1 \f7_reg[26]  ( .D(n945), .CK(clk), .Q(n1287) );
  DFF_X1 \f7_reg[25]  ( .D(n944), .CK(clk), .Q(n1282) );
  DFF_X1 \f7_reg[24]  ( .D(n943), .CK(clk), .Q(n1277) );
  DFF_X1 \f7_reg[23]  ( .D(n942), .CK(clk), .Q(n1272) );
  DFF_X1 \f7_reg[22]  ( .D(n941), .CK(clk), .Q(n1267) );
  DFF_X1 \f_reg[39]  ( .D(n839), .CK(clk), .Q(f[39]), .QN(n26) );
  DFF_X1 \f8_reg[38]  ( .D(n917), .CK(clk), .Q(f8[38]), .QN(n290) );
  DFF_X1 \f_reg[38]  ( .D(n840), .CK(clk), .Q(f[38]), .QN(n25) );
  DFF_X1 \f_reg[37]  ( .D(n841), .CK(clk), .Q(f[37]), .QN(n24) );
  DFF_X1 \f_reg[36]  ( .D(n842), .CK(clk), .Q(f[36]), .QN(n23) );
  DFF_X1 \f_reg[35]  ( .D(n843), .CK(clk), .Q(f[35]), .QN(n22) );
  DFF_X1 \f_reg[34]  ( .D(n844), .CK(clk), .Q(f[34]), .QN(n21) );
  DFF_X1 \f_reg[33]  ( .D(n845), .CK(clk), .Q(f[33]), .QN(n20) );
  DFF_X1 \f_reg[32]  ( .D(n846), .CK(clk), .Q(f[32]), .QN(n19) );
  DFF_X1 \f_reg[31]  ( .D(n847), .CK(clk), .Q(f[31]), .QN(n18) );
  DFF_X1 \f_reg[30]  ( .D(n848), .CK(clk), .Q(f[30]), .QN(n17) );
  DFF_X1 \f_reg[29]  ( .D(n849), .CK(clk), .Q(f[29]), .QN(n16) );
  DFF_X1 \f_reg[28]  ( .D(n850), .CK(clk), .Q(f[28]), .QN(n15) );
  DFF_X1 \f_reg[27]  ( .D(n851), .CK(clk), .Q(f[27]), .QN(n14) );
  DFF_X1 \f_reg[26]  ( .D(n852), .CK(clk), .Q(f[26]), .QN(n13) );
  DFF_X1 \f_reg[25]  ( .D(n853), .CK(clk), .Q(f[25]), .QN(n12) );
  DFF_X1 \f_reg[24]  ( .D(n854), .CK(clk), .Q(f[24]), .QN(n11) );
  DFF_X1 \f_reg[23]  ( .D(n855), .CK(clk), .Q(f[23]), .QN(n10) );
  DFF_X1 \f_reg[22]  ( .D(n856), .CK(clk), .Q(f[22]), .QN(n9) );
  DFF_X1 \f_reg[21]  ( .D(n857), .CK(clk), .Q(f[21]) );
  DFF_X1 \f_reg[20]  ( .D(n858), .CK(clk), .Q(f[20]) );
  DFF_X1 \f_reg[19]  ( .D(n859), .CK(clk), .Q(f[19]) );
  DFF_X1 \f_reg[18]  ( .D(n860), .CK(clk), .Q(f[18]) );
  DFF_X1 \f_reg[17]  ( .D(n861), .CK(clk), .Q(f[17]) );
  DFF_X1 \f_reg[16]  ( .D(n862), .CK(clk), .Q(f[16]) );
  DFF_X1 \f_reg[15]  ( .D(n863), .CK(clk), .Q(f[15]) );
  DFF_X1 \f_reg[14]  ( .D(n864), .CK(clk), .Q(f[14]), .QN(n34) );
  DFF_X1 \f_reg[13]  ( .D(n865), .CK(clk), .Q(f[13]), .QN(n35) );
  DFF_X1 \f_reg[12]  ( .D(n866), .CK(clk), .Q(f[12]), .QN(n36) );
  DFF_X1 \f_reg[11]  ( .D(n867), .CK(clk), .Q(f[11]), .QN(n37) );
  DFF_X1 \f_reg[10]  ( .D(n868), .CK(clk), .Q(f[10]), .QN(n38) );
  DFF_X1 \f_reg[9]  ( .D(n869), .CK(clk), .Q(f[9]), .QN(n39) );
  DFF_X1 \f_reg[8]  ( .D(n870), .CK(clk), .Q(f[8]), .QN(n40) );
  DFF_X1 \f_reg[7]  ( .D(n871), .CK(clk), .Q(f[7]), .QN(n41) );
  DFF_X1 \f_reg[6]  ( .D(n872), .CK(clk), .Q(f[6]), .QN(n42) );
  DFF_X1 \f_reg[5]  ( .D(n873), .CK(clk), .Q(f[5]), .QN(n43) );
  DFF_X1 \f_reg[4]  ( .D(n874), .CK(clk), .Q(f[4]), .QN(n44) );
  DFF_X1 \f_reg[3]  ( .D(n875), .CK(clk), .Q(f[3]), .QN(n45) );
  DFF_X1 \f_reg[2]  ( .D(n876), .CK(clk), .Q(f[2]), .QN(n46) );
  DFF_X1 \f_reg[1]  ( .D(n877), .CK(clk), .Q(f[1]), .QN(n47) );
  DFF_X1 \f_reg[0]  ( .D(n878), .CK(clk), .Q(f[0]), .QN(n48) );
  memory_WIDTH20_SIZE8_LOGSIZE3_0 mem_x ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_x), .addr(addr_x), .wr_en(wr_en_x) );
  memory_WIDTH20_SIZE8_LOGSIZE3_8 mem_a1 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a1), .addr(addr_a1), .wr_en(wr_en_a1) );
  memory_WIDTH20_SIZE8_LOGSIZE3_7 mem_a2 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a2), .addr(addr_a2), .wr_en(wr_en_a2) );
  memory_WIDTH20_SIZE8_LOGSIZE3_6 mem_a3 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a3), .addr(addr_a3), .wr_en(wr_en_a3) );
  memory_WIDTH20_SIZE8_LOGSIZE3_5 mem_a4 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a4), .addr(addr_a4), .wr_en(wr_en_a4) );
  memory_WIDTH20_SIZE8_LOGSIZE3_4 mem_a5 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a5), .addr(addr_a5), .wr_en(wr_en_a5) );
  memory_WIDTH20_SIZE8_LOGSIZE3_3 mem_a6 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a6), .addr(addr_a6), .wr_en(wr_en_a6) );
  memory_WIDTH20_SIZE8_LOGSIZE3_2 mem_a7 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a7), .addr(addr_a7), .wr_en(wr_en_a7) );
  memory_WIDTH20_SIZE8_LOGSIZE3_1 mem_a8 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a8), .addr(addr_a8), .wr_en(wr_en_a8) );
  memory_WIDTH40_SIZE8_LOGSIZE3 mem_y ( .clk(clk), .data_in(f), .data_out(
        data_out), .addr(addr_y), .wr_en(wr_en_y) );
  datapath_DW_mult_tc_8 mult_84 ( .a(data_out_a1), .b(data_out_x), .product({
        \mul_out1[39] , \mul_out1[38] , \mul_out1[37] , \mul_out1[36] , 
        \mul_out1[35] , \mul_out1[34] , \mul_out1[33] , \mul_out1[32] , 
        \mul_out1[31] , \mul_out1[30] , \mul_out1[29] , \mul_out1[28] , 
        \mul_out1[27] , \mul_out1[26] , \mul_out1[25] , \mul_out1[24] , 
        \mul_out1[23] , \mul_out1[22] , \mul_out1[21] , \mul_out1[20] , 
        \mul_out1[19] , \mul_out1[18] , \mul_out1[17] , \mul_out1[16] , 
        \mul_out1[15] , \mul_out1[14] , \mul_out1[13] , \mul_out1[12] , 
        \mul_out1[11] , \mul_out1[10] , \mul_out1[9] , \mul_out1[8] , 
        \mul_out1[7] , \mul_out1[6] , \mul_out1[5] , \mul_out1[4] , 
        \mul_out1[3] , \mul_out1[2] , \mul_out1[1] , \mul_out1[0] }) );
  datapath_DW_mult_tc_9 mult_86 ( .a(data_out_a2), .b(data_out_x), .product({
        \mul_out2[39] , \mul_out2[38] , \mul_out2[37] , \mul_out2[36] , 
        \mul_out2[35] , \mul_out2[34] , \mul_out2[33] , \mul_out2[32] , 
        \mul_out2[31] , \mul_out2[30] , \mul_out2[29] , \mul_out2[28] , 
        \mul_out2[27] , \mul_out2[26] , \mul_out2[25] , \mul_out2[24] , 
        \mul_out2[23] , \mul_out2[22] , \mul_out2[21] , \mul_out2[20] , 
        \mul_out2[19] , \mul_out2[18] , \mul_out2[17] , \mul_out2[16] , 
        \mul_out2[15] , \mul_out2[14] , \mul_out2[13] , \mul_out2[12] , 
        \mul_out2[11] , \mul_out2[10] , \mul_out2[9] , \mul_out2[8] , 
        \mul_out2[7] , \mul_out2[6] , \mul_out2[5] , \mul_out2[4] , 
        \mul_out2[3] , \mul_out2[2] , \mul_out2[1] , \mul_out2[0] }) );
  datapath_DW_mult_tc_10 mult_88 ( .a(data_out_a3), .b(data_out_x), .product({
        \mul_out3[39] , \mul_out3[38] , \mul_out3[37] , \mul_out3[36] , 
        \mul_out3[35] , \mul_out3[34] , \mul_out3[33] , \mul_out3[32] , 
        \mul_out3[31] , \mul_out3[30] , \mul_out3[29] , \mul_out3[28] , 
        \mul_out3[27] , \mul_out3[26] , \mul_out3[25] , \mul_out3[24] , 
        \mul_out3[23] , \mul_out3[22] , \mul_out3[21] , \mul_out3[20] , 
        \mul_out3[19] , \mul_out3[18] , \mul_out3[17] , \mul_out3[16] , 
        \mul_out3[15] , \mul_out3[14] , \mul_out3[13] , \mul_out3[12] , 
        \mul_out3[11] , \mul_out3[10] , \mul_out3[9] , \mul_out3[8] , 
        \mul_out3[7] , \mul_out3[6] , \mul_out3[5] , \mul_out3[4] , 
        \mul_out3[3] , \mul_out3[2] , \mul_out3[1] , \mul_out3[0] }) );
  datapath_DW_mult_tc_11 mult_90 ( .a(data_out_a4), .b(data_out_x), .product({
        \mul_out4[39] , \mul_out4[38] , \mul_out4[37] , \mul_out4[36] , 
        \mul_out4[35] , \mul_out4[34] , \mul_out4[33] , \mul_out4[32] , 
        \mul_out4[31] , \mul_out4[30] , \mul_out4[29] , \mul_out4[28] , 
        \mul_out4[27] , \mul_out4[26] , \mul_out4[25] , \mul_out4[24] , 
        \mul_out4[23] , \mul_out4[22] , \mul_out4[21] , \mul_out4[20] , 
        \mul_out4[19] , \mul_out4[18] , \mul_out4[17] , \mul_out4[16] , 
        \mul_out4[15] , \mul_out4[14] , \mul_out4[13] , \mul_out4[12] , 
        \mul_out4[11] , \mul_out4[10] , \mul_out4[9] , \mul_out4[8] , 
        \mul_out4[7] , \mul_out4[6] , \mul_out4[5] , \mul_out4[4] , 
        \mul_out4[3] , \mul_out4[2] , \mul_out4[1] , \mul_out4[0] }) );
  datapath_DW_mult_tc_12 mult_92 ( .a(data_out_a5), .b(data_out_x), .product({
        \mul_out5[39] , \mul_out5[38] , \mul_out5[37] , \mul_out5[36] , 
        \mul_out5[35] , \mul_out5[34] , \mul_out5[33] , \mul_out5[32] , 
        \mul_out5[31] , \mul_out5[30] , \mul_out5[29] , \mul_out5[28] , 
        \mul_out5[27] , \mul_out5[26] , \mul_out5[25] , \mul_out5[24] , 
        \mul_out5[23] , \mul_out5[22] , \mul_out5[21] , \mul_out5[20] , 
        \mul_out5[19] , \mul_out5[18] , \mul_out5[17] , \mul_out5[16] , 
        \mul_out5[15] , \mul_out5[14] , \mul_out5[13] , \mul_out5[12] , 
        \mul_out5[11] , \mul_out5[10] , \mul_out5[9] , \mul_out5[8] , 
        \mul_out5[7] , \mul_out5[6] , \mul_out5[5] , \mul_out5[4] , 
        \mul_out5[3] , \mul_out5[2] , \mul_out5[1] , \mul_out5[0] }) );
  datapath_DW_mult_tc_13 mult_94 ( .a(data_out_a6), .b(data_out_x), .product({
        \mul_out6[39] , \mul_out6[38] , \mul_out6[37] , \mul_out6[36] , 
        \mul_out6[35] , \mul_out6[34] , \mul_out6[33] , \mul_out6[32] , 
        \mul_out6[31] , \mul_out6[30] , \mul_out6[29] , \mul_out6[28] , 
        \mul_out6[27] , \mul_out6[26] , \mul_out6[25] , \mul_out6[24] , 
        \mul_out6[23] , \mul_out6[22] , \mul_out6[21] , \mul_out6[20] , 
        \mul_out6[19] , \mul_out6[18] , \mul_out6[17] , \mul_out6[16] , 
        \mul_out6[15] , \mul_out6[14] , \mul_out6[13] , \mul_out6[12] , 
        \mul_out6[11] , \mul_out6[10] , \mul_out6[9] , \mul_out6[8] , 
        \mul_out6[7] , \mul_out6[6] , \mul_out6[5] , \mul_out6[4] , 
        \mul_out6[3] , \mul_out6[2] , \mul_out6[1] , \mul_out6[0] }) );
  datapath_DW_mult_tc_14 mult_96 ( .a(data_out_a7), .b(data_out_x), .product({
        \mul_out7[39] , \mul_out7[38] , \mul_out7[37] , \mul_out7[36] , 
        \mul_out7[35] , \mul_out7[34] , \mul_out7[33] , \mul_out7[32] , 
        \mul_out7[31] , \mul_out7[30] , \mul_out7[29] , \mul_out7[28] , 
        \mul_out7[27] , \mul_out7[26] , \mul_out7[25] , \mul_out7[24] , 
        \mul_out7[23] , \mul_out7[22] , \mul_out7[21] , \mul_out7[20] , 
        \mul_out7[19] , \mul_out7[18] , \mul_out7[17] , \mul_out7[16] , 
        \mul_out7[15] , \mul_out7[14] , \mul_out7[13] , \mul_out7[12] , 
        \mul_out7[11] , \mul_out7[10] , \mul_out7[9] , \mul_out7[8] , 
        \mul_out7[7] , \mul_out7[6] , \mul_out7[5] , \mul_out7[4] , 
        \mul_out7[3] , \mul_out7[2] , \mul_out7[1] , \mul_out7[0] }) );
  datapath_DW_mult_tc_15 mult_98 ( .a(data_out_a8), .b(data_out_x), .product({
        \mul_out8[39] , \mul_out8[38] , \mul_out8[37] , \mul_out8[36] , 
        \mul_out8[35] , \mul_out8[34] , \mul_out8[33] , \mul_out8[32] , 
        \mul_out8[31] , \mul_out8[30] , \mul_out8[29] , \mul_out8[28] , 
        \mul_out8[27] , \mul_out8[26] , \mul_out8[25] , \mul_out8[24] , 
        \mul_out8[23] , \mul_out8[22] , \mul_out8[21] , \mul_out8[20] , 
        \mul_out8[19] , \mul_out8[18] , \mul_out8[17] , \mul_out8[16] , 
        \mul_out8[15] , \mul_out8[14] , \mul_out8[13] , \mul_out8[12] , 
        \mul_out8[11] , \mul_out8[10] , \mul_out8[9] , \mul_out8[8] , 
        \mul_out8[7] , \mul_out8[6] , \mul_out8[5] , \mul_out8[4] , 
        \mul_out8[3] , \mul_out8[2] , \mul_out8[1] , \mul_out8[0] }) );
  datapath_DW01_add_8 add_85 ( .A(f1), .B({\mul_out1[39] , \mul_out1[38] , 
        \mul_out1[37] , \mul_out1[36] , \mul_out1[35] , \mul_out1[34] , 
        \mul_out1[33] , \mul_out1[32] , \mul_out1[31] , \mul_out1[30] , 
        \mul_out1[29] , \mul_out1[28] , \mul_out1[27] , \mul_out1[26] , 
        \mul_out1[25] , \mul_out1[24] , \mul_out1[23] , \mul_out1[22] , 
        \mul_out1[21] , \mul_out1[20] , \mul_out1[19] , \mul_out1[18] , 
        \mul_out1[17] , \mul_out1[16] , \mul_out1[15] , \mul_out1[14] , 
        \mul_out1[13] , \mul_out1[12] , \mul_out1[11] , \mul_out1[10] , 
        \mul_out1[9] , \mul_out1[8] , \mul_out1[7] , \mul_out1[6] , 
        \mul_out1[5] , \mul_out1[4] , \mul_out1[3] , \mul_out1[2] , 
        \mul_out1[1] , \mul_out1[0] }), .CI(1'b0), .SUM(add_r1) );
  datapath_DW01_add_9 add_87 ( .A({n766, n768, n770, n772, n774, n776, n778, 
        n780, n782, n784, n786, n788, n790, n792, n794, n796, n798, n800, n802, 
        n804, n806, n808, n810, f2[16:0]}), .B({\mul_out2[39] , \mul_out2[38] , 
        \mul_out2[37] , \mul_out2[36] , \mul_out2[35] , \mul_out2[34] , 
        \mul_out2[33] , \mul_out2[32] , \mul_out2[31] , \mul_out2[30] , 
        \mul_out2[29] , \mul_out2[28] , \mul_out2[27] , \mul_out2[26] , 
        \mul_out2[25] , \mul_out2[24] , \mul_out2[23] , \mul_out2[22] , 
        \mul_out2[21] , \mul_out2[20] , \mul_out2[19] , \mul_out2[18] , 
        \mul_out2[17] , \mul_out2[16] , \mul_out2[15] , \mul_out2[14] , 
        \mul_out2[13] , \mul_out2[12] , \mul_out2[11] , \mul_out2[10] , 
        \mul_out2[9] , \mul_out2[8] , \mul_out2[7] , \mul_out2[6] , 
        \mul_out2[5] , \mul_out2[4] , \mul_out2[3] , \mul_out2[2] , 
        \mul_out2[1] , \mul_out2[0] }), .CI(1'b0), .SUM(add_r2) );
  datapath_DW01_add_10 add_89 ( .A({n642, n644, n646, n647, n649, n650, n652, 
        n654, n656, n658, n660, n662, n664, n666, n668, n670, n672, n674, n676, 
        n678, n680, n682, n684, f3[16:0]}), .B({\mul_out3[39] , \mul_out3[38] , 
        \mul_out3[37] , \mul_out3[36] , \mul_out3[35] , \mul_out3[34] , 
        \mul_out3[33] , \mul_out3[32] , \mul_out3[31] , \mul_out3[30] , 
        \mul_out3[29] , \mul_out3[28] , \mul_out3[27] , \mul_out3[26] , 
        \mul_out3[25] , \mul_out3[24] , \mul_out3[23] , \mul_out3[22] , 
        \mul_out3[21] , \mul_out3[20] , \mul_out3[19] , \mul_out3[18] , 
        \mul_out3[17] , \mul_out3[16] , \mul_out3[15] , \mul_out3[14] , 
        \mul_out3[13] , \mul_out3[12] , \mul_out3[11] , \mul_out3[10] , 
        \mul_out3[9] , \mul_out3[8] , \mul_out3[7] , \mul_out3[6] , 
        \mul_out3[5] , \mul_out3[4] , \mul_out3[3] , \mul_out3[2] , 
        \mul_out3[1] , \mul_out3[0] }), .CI(1'b0), .SUM(add_r3) );
  datapath_DW01_add_11 add_91 ( .A(f4), .B({\mul_out4[39] , \mul_out4[38] , 
        \mul_out4[37] , \mul_out4[36] , \mul_out4[35] , \mul_out4[34] , 
        \mul_out4[33] , \mul_out4[32] , \mul_out4[31] , \mul_out4[30] , 
        \mul_out4[29] , \mul_out4[28] , \mul_out4[27] , \mul_out4[26] , 
        \mul_out4[25] , \mul_out4[24] , \mul_out4[23] , \mul_out4[22] , 
        \mul_out4[21] , \mul_out4[20] , \mul_out4[19] , \mul_out4[18] , 
        \mul_out4[17] , \mul_out4[16] , \mul_out4[15] , \mul_out4[14] , 
        \mul_out4[13] , \mul_out4[12] , \mul_out4[11] , \mul_out4[10] , 
        \mul_out4[9] , \mul_out4[8] , \mul_out4[7] , \mul_out4[6] , 
        \mul_out4[5] , \mul_out4[4] , \mul_out4[3] , \mul_out4[2] , 
        \mul_out4[1] , \mul_out4[0] }), .CI(1'b0), .SUM(add_r4) );
  datapath_DW01_add_12 add_93 ( .A({n703, n705, n707, n709, n711, n713, n715, 
        f5[32], n718, n720, n722, n724, n726, n728, n730, n732, n734, n736, 
        n738, n740, n742, n744, n746, f5[16], n749, f5[14:0]}), .B({
        \mul_out5[39] , \mul_out5[38] , \mul_out5[37] , \mul_out5[36] , 
        \mul_out5[35] , \mul_out5[34] , \mul_out5[33] , \mul_out5[32] , 
        \mul_out5[31] , \mul_out5[30] , \mul_out5[29] , \mul_out5[28] , 
        \mul_out5[27] , \mul_out5[26] , \mul_out5[25] , \mul_out5[24] , 
        \mul_out5[23] , \mul_out5[22] , \mul_out5[21] , \mul_out5[20] , 
        \mul_out5[19] , \mul_out5[18] , \mul_out5[17] , \mul_out5[16] , 
        \mul_out5[15] , \mul_out5[14] , \mul_out5[13] , \mul_out5[12] , 
        \mul_out5[11] , \mul_out5[10] , \mul_out5[9] , \mul_out5[8] , 
        \mul_out5[7] , \mul_out5[6] , \mul_out5[5] , \mul_out5[4] , 
        \mul_out5[3] , \mul_out5[2] , \mul_out5[1] , \mul_out5[0] }), .CI(1'b0), .SUM(add_r5) );
  datapath_DW01_add_13 add_95 ( .A({n1355, n1347, n1342, n1337, n1332, n1327, 
        n1322, n1317, n1313, n1308, n1303, n1298, n1293, n1288, n1283, n1278, 
        n1273, n1268, n479, n481, n483, n485, n487, f6[16:0]}), .B({
        \mul_out6[39] , \mul_out6[38] , \mul_out6[37] , \mul_out6[36] , 
        \mul_out6[35] , \mul_out6[34] , \mul_out6[33] , \mul_out6[32] , 
        \mul_out6[31] , \mul_out6[30] , \mul_out6[29] , \mul_out6[28] , 
        \mul_out6[27] , \mul_out6[26] , \mul_out6[25] , \mul_out6[24] , 
        \mul_out6[23] , \mul_out6[22] , \mul_out6[21] , \mul_out6[20] , 
        \mul_out6[19] , \mul_out6[18] , \mul_out6[17] , \mul_out6[16] , 
        \mul_out6[15] , \mul_out6[14] , \mul_out6[13] , \mul_out6[12] , 
        \mul_out6[11] , \mul_out6[10] , \mul_out6[9] , \mul_out6[8] , 
        \mul_out6[7] , \mul_out6[6] , \mul_out6[5] , \mul_out6[4] , 
        \mul_out6[3] , \mul_out6[2] , \mul_out6[1] , \mul_out6[0] }), .CI(1'b0), .SUM(add_r6) );
  datapath_DW01_add_14 add_97 ( .A({n1353, n1346, n1341, n1336, n1331, n1326, 
        n1321, f7[32], n1312, n1307, n1302, n1297, n1292, n1287, n1282, n1277, 
        n1272, n1267, n534, n536, n538, n540, n542, f7[16], n545, f7[14:0]}), 
        .B({\mul_out7[39] , \mul_out7[38] , \mul_out7[37] , \mul_out7[36] , 
        \mul_out7[35] , \mul_out7[34] , \mul_out7[33] , \mul_out7[32] , 
        \mul_out7[31] , \mul_out7[30] , \mul_out7[29] , \mul_out7[28] , 
        \mul_out7[27] , \mul_out7[26] , \mul_out7[25] , \mul_out7[24] , 
        \mul_out7[23] , \mul_out7[22] , \mul_out7[21] , \mul_out7[20] , 
        \mul_out7[19] , \mul_out7[18] , \mul_out7[17] , \mul_out7[16] , 
        \mul_out7[15] , \mul_out7[14] , \mul_out7[13] , \mul_out7[12] , 
        \mul_out7[11] , \mul_out7[10] , \mul_out7[9] , \mul_out7[8] , 
        \mul_out7[7] , \mul_out7[6] , \mul_out7[5] , \mul_out7[4] , 
        \mul_out7[3] , \mul_out7[2] , \mul_out7[1] , \mul_out7[0] }), .CI(1'b0), .SUM(add_r7) );
  datapath_DW01_add_15 add_99 ( .A(f8), .B({\mul_out8[39] , \mul_out8[38] , 
        \mul_out8[37] , \mul_out8[36] , \mul_out8[35] , \mul_out8[34] , 
        \mul_out8[33] , \mul_out8[32] , \mul_out8[31] , \mul_out8[30] , 
        \mul_out8[29] , \mul_out8[28] , \mul_out8[27] , \mul_out8[26] , 
        \mul_out8[25] , \mul_out8[24] , \mul_out8[23] , \mul_out8[22] , 
        \mul_out8[21] , \mul_out8[20] , \mul_out8[19] , \mul_out8[18] , 
        \mul_out8[17] , \mul_out8[16] , \mul_out8[15] , \mul_out8[14] , 
        \mul_out8[13] , \mul_out8[12] , \mul_out8[11] , \mul_out8[10] , 
        \mul_out8[9] , \mul_out8[8] , \mul_out8[7] , \mul_out8[6] , 
        \mul_out8[5] , \mul_out8[4] , \mul_out8[3] , \mul_out8[2] , 
        \mul_out8[1] , \mul_out8[0] }), .CI(1'b0), .SUM(add_r8) );
  DFF_X2 \f8_reg[34]  ( .D(n913), .CK(clk), .Q(f8[34]), .QN(n294) );
  DFF_X2 \f8_reg[36]  ( .D(n915), .CK(clk), .Q(f8[36]), .QN(n292) );
  DFF_X1 \f4_reg[2]  ( .D(n1041), .CK(clk), .Q(f4[2]), .QN(n166) );
  DFF_X1 \f4_reg[1]  ( .D(n1040), .CK(clk), .Q(f4[1]), .QN(n167) );
  DFF_X1 \f4_reg[0]  ( .D(n1039), .CK(clk), .Q(f4[0]), .QN(n168) );
  DFF_X1 \f1_reg[0]  ( .D(n1159), .CK(clk), .Q(f1[0]), .QN(n1260) );
  DFF_X1 \f8_reg[3]  ( .D(n882), .CK(clk), .Q(f8[3]), .QN(n325) );
  DFF_X1 \f8_reg[2]  ( .D(n881), .CK(clk), .Q(f8[2]), .QN(n326) );
  DFF_X1 \f8_reg[1]  ( .D(n880), .CK(clk), .Q(f8[1]), .QN(n327) );
  DFF_X1 \f8_reg[0]  ( .D(n879), .CK(clk), .Q(f8[0]), .QN(n328) );
  DFF_X1 \f1_reg[3]  ( .D(n1162), .CK(clk), .Q(f1[3]), .QN(n1245) );
  DFF_X1 \f1_reg[2]  ( .D(n1161), .CK(clk), .Q(f1[2]), .QN(n1250) );
  DFF_X1 \f1_reg[1]  ( .D(n1160), .CK(clk), .Q(f1[1]), .QN(n1255) );
  DFF_X1 \f2_reg[1]  ( .D(n1120), .CK(clk), .Q(f2[1]), .QN(n87) );
  DFF_X1 \f2_reg[0]  ( .D(n1119), .CK(clk), .Q(f2[0]), .QN(n88) );
  DFF_X1 \f7_reg[3]  ( .D(n922), .CK(clk), .Q(f7[3]) );
  DFF_X1 \f7_reg[2]  ( .D(n921), .CK(clk), .Q(f7[2]) );
  DFF_X1 \f7_reg[1]  ( .D(n920), .CK(clk), .Q(f7[1]) );
  DFF_X1 \f7_reg[0]  ( .D(n919), .CK(clk), .Q(f7[0]) );
  DFF_X1 \f5_reg[0]  ( .D(n999), .CK(clk), .Q(f5[0]), .QN(n208) );
  DFF_X1 \f3_reg[2]  ( .D(n1081), .CK(clk), .Q(f3[2]) );
  DFF_X1 \f3_reg[1]  ( .D(n1080), .CK(clk), .Q(f3[1]) );
  DFF_X1 \f3_reg[0]  ( .D(n1079), .CK(clk), .Q(f3[0]) );
  DFF_X1 \f4_reg[3]  ( .D(n1042), .CK(clk), .Q(f4[3]), .QN(n165) );
  DFF_X1 \f2_reg[2]  ( .D(n1121), .CK(clk), .Q(f2[2]), .QN(n86) );
  DFF_X1 \f3_reg[3]  ( .D(n1082), .CK(clk), .Q(f3[3]) );
  DFF_X1 \f6_reg[2]  ( .D(n961), .CK(clk), .Q(f6[2]), .QN(n246) );
  DFF_X1 \f6_reg[1]  ( .D(n960), .CK(clk), .Q(f6[1]), .QN(n247) );
  DFF_X1 \f6_reg[0]  ( .D(n959), .CK(clk), .Q(f6[0]), .QN(n248) );
  DFF_X1 \f5_reg[3]  ( .D(n1002), .CK(clk), .Q(f5[3]), .QN(n205) );
  DFF_X1 \f5_reg[2]  ( .D(n1001), .CK(clk), .Q(f5[2]), .QN(n206) );
  DFF_X1 \f5_reg[1]  ( .D(n1000), .CK(clk), .Q(f5[1]), .QN(n207) );
  DFF_X1 \f6_reg[3]  ( .D(n962), .CK(clk), .Q(f6[3]), .QN(n245) );
  DFF_X1 \f2_reg[3]  ( .D(n1122), .CK(clk), .Q(f2[3]), .QN(n85) );
  DFF_X1 \f8_reg[4]  ( .D(n883), .CK(clk), .Q(f8[4]), .QN(n324) );
  DFF_X1 \f5_reg[4]  ( .D(n1003), .CK(clk), .Q(f5[4]), .QN(n204) );
  DFF_X1 \f7_reg[4]  ( .D(n923), .CK(clk), .Q(f7[4]) );
  DFF_X1 \f1_reg[4]  ( .D(n1163), .CK(clk), .Q(f1[4]), .QN(n1240) );
  DFF_X1 \f4_reg[4]  ( .D(n1043), .CK(clk), .Q(f4[4]), .QN(n164) );
  DFF_X1 \f3_reg[4]  ( .D(n1083), .CK(clk), .Q(f3[4]) );
  DFF_X1 \f6_reg[4]  ( .D(n963), .CK(clk), .Q(f6[4]), .QN(n244) );
  DFF_X1 \f2_reg[4]  ( .D(n1123), .CK(clk), .Q(f2[4]), .QN(n84) );
  DFF_X1 \f8_reg[5]  ( .D(n884), .CK(clk), .Q(f8[5]), .QN(n323) );
  DFF_X1 \f5_reg[5]  ( .D(n1004), .CK(clk), .Q(f5[5]), .QN(n203) );
  DFF_X1 \f1_reg[5]  ( .D(n1164), .CK(clk), .Q(f1[5]), .QN(n1235) );
  DFF_X1 \f4_reg[5]  ( .D(n1044), .CK(clk), .Q(f4[5]), .QN(n163) );
  DFF_X1 \f3_reg[5]  ( .D(n1084), .CK(clk), .Q(f3[5]) );
  DFF_X1 \f6_reg[5]  ( .D(n964), .CK(clk), .Q(f6[5]), .QN(n243) );
  DFF_X1 \f2_reg[5]  ( .D(n1124), .CK(clk), .Q(f2[5]), .QN(n83) );
  DFF_X1 \f7_reg[5]  ( .D(n924), .CK(clk), .Q(f7[5]) );
  DFF_X1 \f1_reg[6]  ( .D(n1165), .CK(clk), .Q(f1[6]), .QN(n1230) );
  DFF_X1 \f6_reg[6]  ( .D(n965), .CK(clk), .Q(f6[6]), .QN(n242) );
  DFF_X1 \f8_reg[6]  ( .D(n885), .CK(clk), .Q(f8[6]), .QN(n322) );
  DFF_X1 \f2_reg[6]  ( .D(n1125), .CK(clk), .Q(f2[6]), .QN(n82) );
  DFF_X1 \f5_reg[6]  ( .D(n1005), .CK(clk), .Q(f5[6]), .QN(n202) );
  DFF_X1 \f4_reg[6]  ( .D(n1045), .CK(clk), .Q(f4[6]), .QN(n162) );
  DFF_X1 \f1_reg[7]  ( .D(n1166), .CK(clk), .Q(f1[7]), .QN(n1225) );
  DFF_X1 \f3_reg[6]  ( .D(n1085), .CK(clk), .Q(f3[6]) );
  DFF_X1 \f7_reg[6]  ( .D(n925), .CK(clk), .Q(f7[6]) );
  DFF_X1 \f8_reg[7]  ( .D(n886), .CK(clk), .Q(f8[7]), .QN(n321) );
  DFF_X1 \f4_reg[7]  ( .D(n1046), .CK(clk), .Q(f4[7]), .QN(n161) );
  DFF_X1 \f6_reg[7]  ( .D(n966), .CK(clk), .Q(f6[7]), .QN(n241) );
  DFF_X1 \f2_reg[7]  ( .D(n1126), .CK(clk), .Q(f2[7]), .QN(n81) );
  DFF_X1 \f5_reg[7]  ( .D(n1006), .CK(clk), .Q(f5[7]), .QN(n201) );
  DFF_X1 \f7_reg[7]  ( .D(n926), .CK(clk), .Q(f7[7]) );
  DFF_X1 \f3_reg[7]  ( .D(n1086), .CK(clk), .Q(f3[7]) );
  DFF_X1 \f1_reg[8]  ( .D(n1167), .CK(clk), .Q(f1[8]), .QN(n1220) );
  DFF_X1 \f8_reg[8]  ( .D(n887), .CK(clk), .Q(f8[8]), .QN(n320) );
  DFF_X1 \f2_reg[8]  ( .D(n1127), .CK(clk), .Q(f2[8]), .QN(n80) );
  DFF_X1 \f6_reg[8]  ( .D(n967), .CK(clk), .Q(f6[8]), .QN(n240) );
  DFF_X1 \f1_reg[9]  ( .D(n1168), .CK(clk), .Q(f1[9]), .QN(n1215) );
  DFF_X1 \f8_reg[9]  ( .D(n888), .CK(clk), .Q(f8[9]), .QN(n319) );
  DFF_X1 \f5_reg[8]  ( .D(n1007), .CK(clk), .Q(f5[8]), .QN(n200) );
  DFF_X1 \f7_reg[8]  ( .D(n927), .CK(clk), .Q(f7[8]) );
  DFF_X1 \f4_reg[8]  ( .D(n1047), .CK(clk), .Q(f4[8]), .QN(n160) );
  DFF_X1 \f1_reg[10]  ( .D(n1169), .CK(clk), .Q(f1[10]), .QN(n1210) );
  DFF_X1 \f5_reg[9]  ( .D(n1008), .CK(clk), .Q(f5[9]), .QN(n199) );
  DFF_X1 \f8_reg[10]  ( .D(n889), .CK(clk), .Q(f8[10]), .QN(n318) );
  DFF_X1 \f2_reg[9]  ( .D(n1128), .CK(clk), .Q(f2[9]), .QN(n79) );
  DFF_X1 \f7_reg[9]  ( .D(n928), .CK(clk), .Q(f7[9]) );
  DFF_X1 \f6_reg[9]  ( .D(n968), .CK(clk), .Q(f6[9]), .QN(n239) );
  DFF_X1 \f2_reg[10]  ( .D(n1129), .CK(clk), .Q(f2[10]), .QN(n78) );
  DFF_X1 \f3_reg[8]  ( .D(n1087), .CK(clk), .Q(f3[8]) );
  DFF_X1 \f4_reg[9]  ( .D(n1048), .CK(clk), .Q(f4[9]), .QN(n159) );
  DFF_X1 \f5_reg[10]  ( .D(n1009), .CK(clk), .Q(f5[10]), .QN(n198) );
  DFF_X1 \f7_reg[10]  ( .D(n929), .CK(clk), .Q(f7[10]) );
  DFF_X1 \f6_reg[10]  ( .D(n969), .CK(clk), .Q(f6[10]), .QN(n238) );
  DFF_X1 \f4_reg[10]  ( .D(n1049), .CK(clk), .Q(f4[10]), .QN(n158) );
  DFF_X1 \f1_reg[11]  ( .D(n1170), .CK(clk), .Q(f1[11]), .QN(n1205) );
  DFF_X1 \f8_reg[11]  ( .D(n890), .CK(clk), .Q(f8[11]), .QN(n317) );
  DFF_X1 \f3_reg[9]  ( .D(n1088), .CK(clk), .Q(f3[9]) );
  DFF_X1 \f3_reg[10]  ( .D(n1089), .CK(clk), .Q(f3[10]) );
  DFF_X1 \f2_reg[11]  ( .D(n1130), .CK(clk), .Q(f2[11]), .QN(n77) );
  DFF_X1 \f7_reg[11]  ( .D(n930), .CK(clk), .Q(f7[11]) );
  DFF_X1 \f6_reg[11]  ( .D(n970), .CK(clk), .Q(f6[11]), .QN(n237) );
  DFF_X1 \f5_reg[11]  ( .D(n1010), .CK(clk), .Q(f5[11]), .QN(n197) );
  DFF_X1 \f4_reg[11]  ( .D(n1050), .CK(clk), .Q(f4[11]), .QN(n157) );
  DFF_X1 \f3_reg[11]  ( .D(n1090), .CK(clk), .Q(f3[11]) );
  DFF_X1 \f1_reg[12]  ( .D(n1171), .CK(clk), .Q(f1[12]), .QN(n1200) );
  DFF_X1 \f8_reg[12]  ( .D(n891), .CK(clk), .Q(f8[12]), .QN(n316) );
  DFF_X1 \f4_reg[12]  ( .D(n1051), .CK(clk), .Q(f4[12]), .QN(n156) );
  DFF_X1 \f7_reg[12]  ( .D(n931), .CK(clk), .Q(f7[12]) );
  DFF_X1 \f2_reg[12]  ( .D(n1131), .CK(clk), .Q(f2[12]), .QN(n76) );
  DFF_X1 \f8_reg[14]  ( .D(n893), .CK(clk), .Q(f8[14]), .QN(n314) );
  DFF_X1 \f2_reg[14]  ( .D(n1133), .CK(clk), .Q(f2[14]), .QN(n74) );
  DFF_X1 \f1_reg[14]  ( .D(n1173), .CK(clk), .Q(f1[14]), .QN(n830) );
  DFF_X1 \f1_reg[13]  ( .D(n1172), .CK(clk), .Q(f1[13]), .QN(n835) );
  DFF_X1 \f8_reg[13]  ( .D(n892), .CK(clk), .Q(f8[13]), .QN(n315) );
  DFF_X1 \f2_reg[13]  ( .D(n1132), .CK(clk), .Q(f2[13]), .QN(n75) );
  DFF_X1 \f6_reg[12]  ( .D(n971), .CK(clk), .Q(f6[12]), .QN(n236) );
  DFF_X1 \f4_reg[13]  ( .D(n1052), .CK(clk), .Q(f4[13]), .QN(n155) );
  DFF_X1 \f5_reg[12]  ( .D(n1011), .CK(clk), .Q(f5[12]), .QN(n196) );
  DFF_X1 \f4_reg[14]  ( .D(n1053), .CK(clk), .Q(f4[14]), .QN(n154) );
  DFF_X1 \f3_reg[12]  ( .D(n1091), .CK(clk), .Q(f3[12]) );
  DFF_X1 \f6_reg[14]  ( .D(n973), .CK(clk), .Q(f6[14]), .QN(n234) );
  DFF_X1 \f7_reg[13]  ( .D(n932), .CK(clk), .Q(f7[13]) );
  DFF_X1 \f2_reg[15]  ( .D(n1134), .CK(clk), .Q(f2[15]), .QN(n73) );
  DFF_X1 \f3_reg[14]  ( .D(n1093), .CK(clk), .Q(f3[14]) );
  DFF_X1 \f7_reg[14]  ( .D(n933), .CK(clk), .Q(f7[14]) );
  DFF_X1 \f8_reg[15]  ( .D(n894), .CK(clk), .Q(f8[15]), .QN(n313) );
  DFF_X1 \f5_reg[14]  ( .D(n1013), .CK(clk), .Q(f5[14]), .QN(n194) );
  DFF_X1 \f3_reg[13]  ( .D(n1092), .CK(clk), .Q(f3[13]) );
  DFF_X1 \f1_reg[15]  ( .D(n1174), .CK(clk), .Q(f1[15]), .QN(n33) );
  DFF_X1 \f4_reg[15]  ( .D(n1054), .CK(clk), .Q(f4[15]), .QN(n153) );
  DFF_X1 \f3_reg[15]  ( .D(n1094), .CK(clk), .Q(f3[15]), .QN(n113) );
  DFF_X1 \f6_reg[13]  ( .D(n972), .CK(clk), .Q(f6[13]), .QN(n235) );
  DFF_X1 \f5_reg[13]  ( .D(n1012), .CK(clk), .Q(f5[13]), .QN(n195) );
  DFF_X1 \f7_reg[15]  ( .D(n934), .CK(clk), .Q(n545), .QN(n273) );
  DFF_X1 \f6_reg[15]  ( .D(n974), .CK(clk), .Q(f6[15]), .QN(n233) );
  DFF_X1 \f5_reg[15]  ( .D(n1014), .CK(clk), .Q(n749), .QN(n193) );
  DFF_X1 \f8_reg[16]  ( .D(n895), .CK(clk), .Q(f8[16]), .QN(n312) );
  DFF_X1 \f6_reg[16]  ( .D(n975), .CK(clk), .Q(f6[16]), .QN(n232) );
  DFF_X1 \f2_reg[16]  ( .D(n1135), .CK(clk), .Q(f2[16]), .QN(n72) );
  DFF_X1 \f8_reg[18]  ( .D(n897), .CK(clk), .Q(f8[18]), .QN(n310) );
  DFF_X1 \f8_reg[17]  ( .D(n896), .CK(clk), .Q(f8[17]), .QN(n311) );
  DFF_X1 \f8_reg[19]  ( .D(n898), .CK(clk), .Q(f8[19]), .QN(n309) );
  DFF_X1 \f3_reg[16]  ( .D(n1095), .CK(clk), .Q(f3[16]), .QN(n112) );
  DFF_X1 \f5_reg[16]  ( .D(n1015), .CK(clk), .Q(f5[16]), .QN(n192) );
  DFF_X1 \f1_reg[16]  ( .D(n1175), .CK(clk), .Q(f1[16]), .QN(n32) );
  DFF_X1 \f6_reg[19]  ( .D(n978), .CK(clk), .Q(n483), .QN(n229) );
  DFF_X1 \f6_reg[18]  ( .D(n977), .CK(clk), .Q(n485), .QN(n230) );
  DFF_X1 \f6_reg[17]  ( .D(n976), .CK(clk), .Q(n487), .QN(n231) );
  DFF_X1 \f8_reg[20]  ( .D(n899), .CK(clk), .Q(f8[20]), .QN(n308) );
  DFF_X1 \f4_reg[16]  ( .D(n1055), .CK(clk), .Q(f4[16]), .QN(n152) );
  DFF_X1 \f7_reg[16]  ( .D(n935), .CK(clk), .Q(f7[16]), .QN(n272) );
  DFF_X1 \f8_reg[21]  ( .D(n900), .CK(clk), .Q(f8[21]), .QN(n307) );
  DFF_X1 \f6_reg[20]  ( .D(n979), .CK(clk), .Q(n481), .QN(n228) );
  DFF_X1 \f2_reg[19]  ( .D(n1138), .CK(clk), .Q(n806), .QN(n69) );
  DFF_X1 \f2_reg[18]  ( .D(n1137), .CK(clk), .Q(n808), .QN(n70) );
  DFF_X1 \f2_reg[17]  ( .D(n1136), .CK(clk), .Q(n810), .QN(n71) );
  DFF_X1 \f2_reg[20]  ( .D(n1139), .CK(clk), .Q(n804), .QN(n68) );
  DFF_X1 \f6_reg[21]  ( .D(n980), .CK(clk), .Q(n479), .QN(n227) );
  DFF_X1 \f8_reg[22]  ( .D(n901), .CK(clk), .Q(f8[22]), .QN(n306) );
  DFF_X1 \f1_reg[21]  ( .D(n1180), .CK(clk), .Q(f1[21]), .QN(n27) );
  DFF_X1 \f1_reg[20]  ( .D(n1179), .CK(clk), .Q(f1[20]), .QN(n28) );
  DFF_X1 \f1_reg[19]  ( .D(n1178), .CK(clk), .Q(f1[19]), .QN(n29) );
  DFF_X1 \f1_reg[18]  ( .D(n1177), .CK(clk), .Q(f1[18]), .QN(n30) );
  DFF_X1 \f1_reg[17]  ( .D(n1176), .CK(clk), .Q(f1[17]), .QN(n31) );
  DFF_X1 \f2_reg[21]  ( .D(n1140), .CK(clk), .Q(n802), .QN(n67) );
  DFF_X1 \f1_reg[22]  ( .D(n1181), .CK(clk), .Q(f1[22]), .QN(n1265) );
  DFF_X1 \f3_reg[19]  ( .D(n1098), .CK(clk), .Q(n680), .QN(n109) );
  DFF_X1 \f3_reg[18]  ( .D(n1097), .CK(clk), .Q(n682), .QN(n110) );
  DFF_X1 \f3_reg[17]  ( .D(n1096), .CK(clk), .Q(n684), .QN(n111) );
  DFF_X1 \f3_reg[22]  ( .D(n1101), .CK(clk), .Q(n674), .QN(n106) );
  DFF_X1 \f3_reg[21]  ( .D(n1100), .CK(clk), .Q(n676), .QN(n107) );
  DFF_X1 \f3_reg[20]  ( .D(n1099), .CK(clk), .Q(n678), .QN(n108) );
  DFF_X1 \f8_reg[23]  ( .D(n902), .CK(clk), .Q(f8[23]), .QN(n305) );
  DFF_X1 \f3_reg[23]  ( .D(n1102), .CK(clk), .Q(n672), .QN(n105) );
  DFF_X1 \f5_reg[21]  ( .D(n1020), .CK(clk), .Q(n738), .QN(n187) );
  DFF_X1 \f5_reg[20]  ( .D(n1019), .CK(clk), .Q(n740), .QN(n188) );
  DFF_X1 \f5_reg[19]  ( .D(n1018), .CK(clk), .Q(n742), .QN(n189) );
  DFF_X1 \f5_reg[18]  ( .D(n1017), .CK(clk), .Q(n744), .QN(n190) );
  DFF_X1 \f5_reg[17]  ( .D(n1016), .CK(clk), .Q(n746), .QN(n191) );
  DFF_X1 \f2_reg[22]  ( .D(n1141), .CK(clk), .Q(n800), .QN(n66) );
  DFF_X1 \f1_reg[23]  ( .D(n1182), .CK(clk), .Q(f1[23]), .QN(n1270) );
  DFF_X1 \f5_reg[22]  ( .D(n1021), .CK(clk), .Q(n736), .QN(n186) );
  DFF_X1 \f4_reg[21]  ( .D(n1060), .CK(clk), .Q(f4[21]), .QN(n147) );
  DFF_X1 \f4_reg[20]  ( .D(n1059), .CK(clk), .Q(f4[20]), .QN(n148) );
  DFF_X1 \f4_reg[19]  ( .D(n1058), .CK(clk), .Q(f4[19]), .QN(n149) );
  DFF_X1 \f4_reg[18]  ( .D(n1057), .CK(clk), .Q(f4[18]), .QN(n150) );
  DFF_X1 \f4_reg[17]  ( .D(n1056), .CK(clk), .Q(f4[17]), .QN(n151) );
  DFF_X1 \f2_reg[23]  ( .D(n1142), .CK(clk), .Q(n798), .QN(n65) );
  DFF_X1 \f5_reg[23]  ( .D(n1022), .CK(clk), .Q(n734), .QN(n185) );
  DFF_X1 \f4_reg[22]  ( .D(n1061), .CK(clk), .Q(f4[22]), .QN(n146) );
  DFF_X1 \f7_reg[21]  ( .D(n940), .CK(clk), .Q(n534), .QN(n267) );
  DFF_X1 \f7_reg[20]  ( .D(n939), .CK(clk), .Q(n536), .QN(n268) );
  DFF_X1 \f7_reg[19]  ( .D(n938), .CK(clk), .Q(n538), .QN(n269) );
  DFF_X1 \f7_reg[18]  ( .D(n937), .CK(clk), .Q(n540), .QN(n270) );
  DFF_X1 \f7_reg[17]  ( .D(n936), .CK(clk), .Q(n542), .QN(n271) );
  DFF_X1 \f8_reg[32]  ( .D(n911), .CK(clk), .Q(f8[32]), .QN(n296) );
  DFF_X1 \f4_reg[23]  ( .D(n1062), .CK(clk), .Q(f4[23]), .QN(n145) );
  DFF_X1 \f4_reg[24]  ( .D(n1063), .CK(clk), .Q(f4[24]), .QN(n144) );
  DFF_X1 \f7_reg[32]  ( .D(n951), .CK(clk), .Q(f7[32]) );
  DFF_X1 \f2_reg[32]  ( .D(n1151), .CK(clk), .Q(n780), .QN(n56) );
  DFF_X1 \f3_reg[32]  ( .D(n1111), .CK(clk), .Q(n654), .QN(n96) );
  DFF_X1 \f3_reg[24]  ( .D(n1103), .CK(clk), .Q(n670), .QN(n104) );
  DFF_X1 \f8_reg[24]  ( .D(n903), .CK(clk), .Q(f8[24]), .QN(n304) );
  DFF_X1 \f5_reg[24]  ( .D(n1023), .CK(clk), .Q(n732), .QN(n184) );
  DFF_X1 \f4_reg[26]  ( .D(n1065), .CK(clk), .Q(f4[26]), .QN(n142) );
  DFF_X1 \f4_reg[27]  ( .D(n1066), .CK(clk), .Q(f4[27]), .QN(n141) );
  DFF_X1 \f4_reg[25]  ( .D(n1064), .CK(clk), .Q(f4[25]), .QN(n143) );
  DFF_X1 \f2_reg[24]  ( .D(n1143), .CK(clk), .Q(n796), .QN(n64) );
  DFF_X1 \f5_reg[31]  ( .D(n1030), .CK(clk), .Q(n718), .QN(n177) );
  DFF_X1 \f3_reg[28]  ( .D(n1107), .CK(clk), .Q(n662), .QN(n100) );
  DFF_X1 \f3_reg[27]  ( .D(n1106), .CK(clk), .Q(n664), .QN(n101) );
  DFF_X1 \f3_reg[26]  ( .D(n1105), .CK(clk), .Q(n666), .QN(n102) );
  DFF_X1 \f3_reg[25]  ( .D(n1104), .CK(clk), .Q(n668), .QN(n103) );
  DFF_X1 \f1_reg[31]  ( .D(n1190), .CK(clk), .Q(f1[31]), .QN(n1310) );
  DFF_X1 \f8_reg[28]  ( .D(n907), .CK(clk), .Q(f8[28]), .QN(n300) );
  DFF_X1 \f8_reg[29]  ( .D(n908), .CK(clk), .Q(f8[29]), .QN(n299) );
  DFF_X1 \f8_reg[30]  ( .D(n909), .CK(clk), .Q(f8[30]), .QN(n298) );
  DFF_X1 \f8_reg[26]  ( .D(n905), .CK(clk), .Q(f8[26]), .QN(n302) );
  DFF_X1 \f8_reg[27]  ( .D(n906), .CK(clk), .Q(f8[27]), .QN(n301) );
  DFF_X1 \f8_reg[25]  ( .D(n904), .CK(clk), .Q(f8[25]), .QN(n303) );
  DFF_X1 \f1_reg[37]  ( .D(n1196), .CK(clk), .Q(f1[37]), .QN(n1339) );
  DFF_X1 \f8_reg[35]  ( .D(n914), .CK(clk), .Q(f8[35]), .QN(n293) );
  DFF_X1 \f4_reg[38]  ( .D(n1077), .CK(clk), .Q(f4[38]), .QN(n130) );
  DFF_X1 \f8_reg[31]  ( .D(n910), .CK(clk), .Q(f8[31]), .QN(n297) );
  DFF_X1 \f8_reg[33]  ( .D(n912), .CK(clk), .Q(f8[33]), .QN(n295) );
  DFF_X1 \f5_reg[36]  ( .D(n1035), .CK(clk), .Q(n709), .QN(n172) );
  DFF_X1 \f5_reg[39]  ( .D(n1038), .CK(clk), .Q(n703), .QN(n169) );
  DFF_X1 \f5_reg[33]  ( .D(n1032), .CK(clk), .Q(n715), .QN(n175) );
  DFF_X1 \f8_reg[39]  ( .D(n918), .CK(clk), .Q(f8[39]), .QN(n289) );
  DFF_X1 \f2_reg[31]  ( .D(n1150), .CK(clk), .Q(n782), .QN(n57) );
  DFF_X1 \f1_reg[32]  ( .D(n1191), .CK(clk), .Q(f1[32]), .QN(n1315) );
  DFF_X1 \f3_reg[33]  ( .D(n1112), .CK(clk), .Q(n652), .QN(n95) );
  DFF_X1 \f3_reg[38]  ( .D(n1117), .CK(clk), .Q(n644), .QN(n90) );
  DFF_X1 \f5_reg[28]  ( .D(n1027), .CK(clk), .Q(n724), .QN(n180) );
  DFF_X1 \f5_reg[27]  ( .D(n1026), .CK(clk), .Q(n726), .QN(n181) );
  DFF_X1 \f5_reg[26]  ( .D(n1025), .CK(clk), .Q(n728), .QN(n182) );
  DFF_X1 \f5_reg[25]  ( .D(n1024), .CK(clk), .Q(n730), .QN(n183) );
  DFF_X1 \f2_reg[28]  ( .D(n1147), .CK(clk), .Q(n788), .QN(n60) );
  DFF_X1 \f2_reg[26]  ( .D(n1145), .CK(clk), .Q(n792), .QN(n62) );
  DFF_X1 \f2_reg[25]  ( .D(n1144), .CK(clk), .Q(n794), .QN(n63) );
  DFF_X1 \f2_reg[27]  ( .D(n1146), .CK(clk), .Q(n790), .QN(n61) );
  DFF_X1 \f4_reg[35]  ( .D(n1074), .CK(clk), .Q(f4[35]), .QN(n133) );
  DFF_X1 \f3_reg[30]  ( .D(n1109), .CK(clk), .Q(n658), .QN(n98) );
  DFF_X1 \f3_reg[29]  ( .D(n1108), .CK(clk), .Q(n660), .QN(n99) );
  DFF_X1 \f4_reg[39]  ( .D(n1078), .CK(clk), .Q(f4[39]), .QN(n129) );
  DFF_X1 \f4_reg[37]  ( .D(n1076), .CK(clk), .Q(f4[37]), .QN(n131) );
  DFF_X1 \f1_reg[39]  ( .D(n1198), .CK(clk), .Q(f1[39]), .QN(n1349) );
  DFF_X1 \f1_reg[35]  ( .D(n1194), .CK(clk), .Q(f1[35]), .QN(n1329) );
  DFF_X1 \f3_reg[36]  ( .D(n1115), .CK(clk), .Q(n647), .QN(n92) );
  DFF_X1 \f3_reg[34]  ( .D(n1113), .CK(clk), .Q(n650), .QN(n94) );
  DFF_X1 \f2_reg[37]  ( .D(n1156), .CK(clk), .Q(n770), .QN(n51) );
  DFF_X1 \f2_reg[36]  ( .D(n1155), .CK(clk), .Q(n772), .QN(n52) );
  DFF_X1 \f2_reg[33]  ( .D(n1152), .CK(clk), .Q(n778), .QN(n55) );
  DFF_X1 \f2_reg[38]  ( .D(n1157), .CK(clk), .Q(n768), .QN(n50) );
  DFF_X1 \f1_reg[29]  ( .D(n1188), .CK(clk), .Q(f1[29]), .QN(n1300) );
  DFF_X1 \f8_reg[37]  ( .D(n916), .CK(clk), .Q(f8[37]), .QN(n291) );
  DFF_X1 \f3_reg[31]  ( .D(n1110), .CK(clk), .Q(n656), .QN(n97) );
  DFF_X1 \f1_reg[38]  ( .D(n1197), .CK(clk), .Q(f1[38]), .QN(n1344) );
  DFF_X1 \f5_reg[32]  ( .D(n1031), .CK(clk), .Q(f5[32]), .QN(n176) );
  DFF_X1 \f5_reg[34]  ( .D(n1033), .CK(clk), .Q(n713), .QN(n174) );
  DFF_X1 \f5_reg[37]  ( .D(n1036), .CK(clk), .Q(n707), .QN(n171) );
  DFF_X1 \f5_reg[35]  ( .D(n1034), .CK(clk), .Q(n711), .QN(n173) );
  DFF_X1 \f5_reg[38]  ( .D(n1037), .CK(clk), .Q(n705), .QN(n170) );
  DFF_X1 \f6_reg[27]  ( .D(n986), .CK(clk), .Q(n1293) );
  DFF_X1 \f6_reg[28]  ( .D(n987), .CK(clk), .Q(n1298) );
  DFF_X1 \f6_reg[26]  ( .D(n985), .CK(clk), .Q(n1288) );
  DFF_X1 \f6_reg[25]  ( .D(n984), .CK(clk), .Q(n1283) );
  DFF_X1 \f6_reg[38]  ( .D(n997), .CK(clk), .Q(n1347) );
  DFF_X1 \f6_reg[29]  ( .D(n988), .CK(clk), .Q(n1303) );
  DFF_X1 \f6_reg[31]  ( .D(n990), .CK(clk), .Q(n1313) );
  DFF_X1 \f7_reg[36]  ( .D(n955), .CK(clk), .Q(n1336) );
  DFF_X1 \f7_reg[39]  ( .D(n958), .CK(clk), .Q(n1353) );
  DFF_X1 \f7_reg[35]  ( .D(n954), .CK(clk), .Q(n1331) );
  DFF_X1 \f7_reg[38]  ( .D(n957), .CK(clk), .Q(n1346) );
  DFF_X2 \f1_reg[30]  ( .D(n1189), .CK(clk), .Q(f1[30]), .QN(n1305) );
  DFF_X1 \f2_reg[29]  ( .D(n1148), .CK(clk), .Q(n786), .QN(n59) );
  DFF_X1 \f4_reg[33]  ( .D(n1072), .CK(clk), .Q(f4[33]), .QN(n135) );
  DFF_X1 \f4_reg[34]  ( .D(n1073), .CK(clk), .Q(f4[34]), .QN(n134) );
  DFF_X1 \f4_reg[36]  ( .D(n1075), .CK(clk), .Q(f4[36]), .QN(n132) );
  OR2_X1 U3 ( .A1(n132), .A2(n286), .ZN(n1) );
  NAND2_X1 U4 ( .A1(n1), .A2(n605), .ZN(n1075) );
  OR2_X1 U5 ( .A1(n1344), .A2(n278), .ZN(n2) );
  NAND2_X1 U6 ( .A1(n2), .A2(n370), .ZN(n1197) );
  OR2_X1 U7 ( .A1(n1349), .A2(n278), .ZN(n3) );
  NAND2_X1 U8 ( .A1(n3), .A2(n369), .ZN(n1198) );
  OR2_X1 U9 ( .A1(n1334), .A2(n279), .ZN(n4) );
  NAND2_X1 U10 ( .A1(n4), .A2(n374), .ZN(n1195) );
  OR2_X1 U11 ( .A1(n292), .A2(n281), .ZN(n5) );
  NAND2_X1 U12 ( .A1(n5), .A2(n565), .ZN(n915) );
  OR2_X1 U13 ( .A1(n294), .A2(n282), .ZN(n6) );
  NAND2_X1 U14 ( .A1(n567), .A2(n6), .ZN(n913) );
  AND3_X1 U15 ( .A1(clc), .A2(n1357), .A3(n366), .ZN(n7) );
  AND2_X1 U16 ( .A1(n278), .A2(n1357), .ZN(n8) );
  AOI22_X1 U17 ( .A1(n828), .A2(n646), .B1(add_r3[37]), .B2(n8), .ZN(n114) );
  INV_X1 U18 ( .A(n114), .ZN(n1116) );
  AOI22_X1 U19 ( .A1(n828), .A2(n649), .B1(add_r3[35]), .B2(n8), .ZN(n115) );
  INV_X1 U20 ( .A(n115), .ZN(n1114) );
  OR2_X1 U21 ( .A1(n293), .A2(n281), .ZN(n116) );
  NAND2_X1 U22 ( .A1(n116), .A2(n566), .ZN(n914) );
  OR2_X1 U23 ( .A1(n1339), .A2(n278), .ZN(n117) );
  NAND2_X1 U24 ( .A1(n117), .A2(n373), .ZN(n1196) );
  OR2_X1 U25 ( .A1(n1310), .A2(n279), .ZN(n118) );
  NAND2_X1 U26 ( .A1(n118), .A2(n385), .ZN(n1190) );
  OR2_X1 U27 ( .A1(n130), .A2(n286), .ZN(n119) );
  NAND2_X1 U28 ( .A1(n119), .A2(n603), .ZN(n1077) );
  OR2_X1 U29 ( .A1(n291), .A2(n281), .ZN(n120) );
  NAND2_X1 U30 ( .A1(n120), .A2(n564), .ZN(n916) );
  OR2_X1 U31 ( .A1(n1324), .A2(n279), .ZN(n121) );
  NAND2_X1 U32 ( .A1(n378), .A2(n121), .ZN(n1193) );
  OR2_X1 U33 ( .A1(n295), .A2(n282), .ZN(n122) );
  NAND2_X1 U34 ( .A1(n122), .A2(n568), .ZN(n912) );
  OR2_X1 U35 ( .A1(n290), .A2(n281), .ZN(n123) );
  NAND2_X1 U36 ( .A1(n123), .A2(n563), .ZN(n917) );
  INV_X1 U37 ( .A(n354), .ZN(n353) );
  BUF_X1 U38 ( .A(n125), .Z(n215) );
  BUF_X1 U39 ( .A(n125), .Z(n216) );
  BUF_X1 U40 ( .A(n125), .Z(n212) );
  BUF_X1 U41 ( .A(n125), .Z(n213) );
  BUF_X1 U42 ( .A(n125), .Z(n214) );
  BUF_X1 U43 ( .A(n126), .Z(n220) );
  BUF_X1 U44 ( .A(n126), .Z(n219) );
  BUF_X1 U45 ( .A(n126), .Z(n217) );
  BUF_X1 U46 ( .A(n126), .Z(n218) );
  BUF_X1 U47 ( .A(n125), .Z(n211) );
  BUF_X1 U48 ( .A(n128), .Z(n256) );
  BUF_X1 U49 ( .A(n128), .Z(n254) );
  BUF_X1 U50 ( .A(n128), .Z(n253) );
  BUF_X1 U51 ( .A(n128), .Z(n252) );
  BUF_X1 U52 ( .A(n128), .Z(n255) );
  BUF_X1 U53 ( .A(n127), .Z(n250) );
  BUF_X1 U54 ( .A(n127), .Z(n249) );
  BUF_X1 U55 ( .A(n126), .Z(n221) );
  BUF_X1 U56 ( .A(n126), .Z(n222) );
  BUF_X1 U57 ( .A(n127), .Z(n223) );
  BUF_X1 U58 ( .A(n128), .Z(n251) );
  BUF_X1 U59 ( .A(n127), .Z(n224) );
  BUF_X1 U60 ( .A(n127), .Z(n225) );
  BUF_X1 U61 ( .A(n127), .Z(n226) );
  BUF_X1 U62 ( .A(n1352), .Z(n346) );
  INV_X1 U63 ( .A(n278), .ZN(n258) );
  BUF_X1 U64 ( .A(n341), .Z(n357) );
  BUF_X1 U65 ( .A(n345), .Z(n347) );
  BUF_X1 U66 ( .A(n344), .Z(n348) );
  BUF_X1 U67 ( .A(n209), .Z(n128) );
  BUF_X1 U68 ( .A(n209), .Z(n127) );
  BUF_X1 U69 ( .A(n210), .Z(n126) );
  BUF_X1 U70 ( .A(n210), .Z(n125) );
  INV_X1 U71 ( .A(n510), .ZN(n1359) );
  BUF_X1 U72 ( .A(n340), .Z(n358) );
  INV_X1 U73 ( .A(n337), .ZN(n342) );
  NOR3_X1 U74 ( .A1(n508), .A2(n509), .A3(n510), .ZN(n506) );
  NAND2_X1 U75 ( .A1(n512), .A2(n511), .ZN(n349) );
  INV_X1 U76 ( .A(n7), .ZN(n335) );
  INV_X1 U77 ( .A(n7), .ZN(n336) );
  NAND2_X1 U78 ( .A1(n506), .A2(n507), .ZN(n343) );
  NAND2_X1 U79 ( .A1(n511), .A2(n1360), .ZN(n510) );
  INV_X1 U80 ( .A(n512), .ZN(n1360) );
  BUF_X1 U81 ( .A(n332), .Z(n278) );
  NAND2_X1 U82 ( .A1(n506), .A2(n1358), .ZN(n345) );
  INV_X1 U83 ( .A(n507), .ZN(n1358) );
  BUF_X1 U84 ( .A(n333), .Z(n277) );
  BUF_X1 U85 ( .A(n333), .Z(n276) );
  NAND2_X1 U86 ( .A1(n1359), .A2(n508), .ZN(n344) );
  AND2_X1 U87 ( .A1(n509), .A2(n1359), .ZN(n341) );
  BUF_X1 U88 ( .A(n1350), .Z(n337) );
  BUF_X1 U89 ( .A(n8), .Z(n209) );
  BUF_X1 U90 ( .A(n8), .Z(n210) );
  NAND2_X1 U91 ( .A1(n512), .A2(n511), .ZN(n124) );
  NAND2_X1 U92 ( .A1(n515), .A2(n1361), .ZN(n350) );
  AND2_X1 U93 ( .A1(n513), .A2(n1361), .ZN(n340) );
  BUF_X1 U94 ( .A(n330), .Z(n284) );
  BUF_X1 U95 ( .A(n330), .Z(n285) );
  BUF_X1 U96 ( .A(n330), .Z(n283) );
  BUF_X1 U97 ( .A(n330), .Z(n282) );
  BUF_X1 U98 ( .A(n330), .Z(n288) );
  BUF_X1 U99 ( .A(n330), .Z(n287) );
  BUF_X1 U100 ( .A(n330), .Z(n286) );
  BUF_X1 U101 ( .A(n330), .Z(n281) );
  BUF_X1 U102 ( .A(n332), .Z(n280) );
  BUF_X1 U103 ( .A(n332), .Z(n279) );
  BUF_X1 U104 ( .A(n330), .Z(n329) );
  NOR3_X1 U105 ( .A1(n513), .A2(n515), .A3(n516), .ZN(n511) );
  NOR3_X1 U106 ( .A1(n361), .A2(addr_y[2]), .A3(n362), .ZN(n508) );
  NOR3_X1 U107 ( .A1(n361), .A2(addr_y[1]), .A3(n365), .ZN(n515) );
  NOR3_X1 U108 ( .A1(n365), .A2(addr_y[0]), .A3(n362), .ZN(n513) );
  NOR2_X1 U109 ( .A1(n365), .A2(addr_y[0]), .ZN(n512) );
  NOR2_X1 U110 ( .A1(n362), .A2(addr_y[0]), .ZN(n509) );
  BUF_X1 U111 ( .A(n334), .Z(n332) );
  BUF_X1 U112 ( .A(n334), .Z(n333) );
  NOR2_X1 U113 ( .A1(n361), .A2(addr_y[1]), .ZN(n507) );
  INV_X1 U114 ( .A(n516), .ZN(n1361) );
  BUF_X1 U115 ( .A(n334), .Z(n330) );
  BUF_X1 U116 ( .A(n334), .Z(n331) );
  NAND2_X1 U117 ( .A1(n351), .A2(n352), .ZN(n840) );
  NAND2_X1 U118 ( .A1(n338), .A2(n339), .ZN(n839) );
  OAI222_X1 U119 ( .A1(n353), .A2(n113), .B1(n344), .B2(n193), .C1(n347), .C2(
        n73), .ZN(n445) );
  OAI222_X1 U120 ( .A1(n353), .A2(n112), .B1(n344), .B2(n192), .C1(n347), .C2(
        n72), .ZN(n441) );
  OAI222_X1 U121 ( .A1(n353), .A2(n111), .B1(n344), .B2(n191), .C1(n347), .C2(
        n71), .ZN(n437) );
  OAI222_X1 U122 ( .A1(n353), .A2(n110), .B1(n344), .B2(n190), .C1(n347), .C2(
        n70), .ZN(n433) );
  OAI222_X1 U123 ( .A1(n353), .A2(n109), .B1(n344), .B2(n189), .C1(n347), .C2(
        n69), .ZN(n429) );
  OAI222_X1 U124 ( .A1(n353), .A2(n108), .B1(n344), .B2(n188), .C1(n347), .C2(
        n68), .ZN(n425) );
  OAI222_X1 U125 ( .A1(n353), .A2(n107), .B1(n344), .B2(n187), .C1(n347), .C2(
        n67), .ZN(n421) );
  INV_X1 U126 ( .A(n828), .ZN(n334) );
  NAND2_X1 U127 ( .A1(clc1), .A2(n1357), .ZN(n516) );
  NAND2_X1 U128 ( .A1(n415), .A2(n416), .ZN(n856) );
  NAND2_X1 U129 ( .A1(n411), .A2(n412), .ZN(n855) );
  NAND2_X1 U130 ( .A1(n407), .A2(n408), .ZN(n854) );
  NAND2_X1 U131 ( .A1(n403), .A2(n404), .ZN(n853) );
  NAND2_X1 U132 ( .A1(n399), .A2(n400), .ZN(n852) );
  NAND2_X1 U133 ( .A1(n395), .A2(n396), .ZN(n851) );
  NAND2_X1 U134 ( .A1(n391), .A2(n392), .ZN(n850) );
  NAND2_X1 U135 ( .A1(n387), .A2(n388), .ZN(n849) );
  NAND2_X1 U136 ( .A1(n383), .A2(n384), .ZN(n848) );
  NAND2_X1 U137 ( .A1(n379), .A2(n380), .ZN(n847) );
  NAND2_X1 U138 ( .A1(n375), .A2(n376), .ZN(n846) );
  NAND2_X1 U139 ( .A1(n371), .A2(n372), .ZN(n845) );
  NAND2_X1 U140 ( .A1(n367), .A2(n368), .ZN(n844) );
  NAND2_X1 U141 ( .A1(n363), .A2(n364), .ZN(n843) );
  NAND2_X1 U142 ( .A1(n359), .A2(n360), .ZN(n842) );
  NAND2_X1 U143 ( .A1(n355), .A2(n356), .ZN(n841) );
  NAND2_X1 U144 ( .A1(n443), .A2(n444), .ZN(n863) );
  AOI221_X1 U145 ( .B1(f1[15]), .B2(n7), .C1(f[15]), .C2(n342), .A(n446), .ZN(
        n443) );
  AOI221_X1 U146 ( .B1(f8[15]), .B2(n340), .C1(f4[15]), .C2(n341), .A(n445), 
        .ZN(n444) );
  OAI22_X1 U147 ( .A1(n124), .A2(n233), .B1(n350), .B2(n273), .ZN(n446) );
  NAND2_X1 U148 ( .A1(n439), .A2(n440), .ZN(n862) );
  AOI221_X1 U149 ( .B1(f1[16]), .B2(n7), .C1(f[16]), .C2(n342), .A(n442), .ZN(
        n439) );
  AOI221_X1 U150 ( .B1(f8[16]), .B2(n340), .C1(f4[16]), .C2(n341), .A(n441), 
        .ZN(n440) );
  OAI22_X1 U151 ( .A1(n349), .A2(n232), .B1(n350), .B2(n272), .ZN(n442) );
  NAND2_X1 U152 ( .A1(n435), .A2(n436), .ZN(n861) );
  AOI221_X1 U153 ( .B1(f1[17]), .B2(n7), .C1(f[17]), .C2(n342), .A(n438), .ZN(
        n435) );
  AOI221_X1 U154 ( .B1(f8[17]), .B2(n340), .C1(f4[17]), .C2(n341), .A(n437), 
        .ZN(n436) );
  OAI22_X1 U155 ( .A1(n124), .A2(n231), .B1(n350), .B2(n271), .ZN(n438) );
  NAND2_X1 U156 ( .A1(n431), .A2(n432), .ZN(n860) );
  AOI221_X1 U157 ( .B1(f1[18]), .B2(n7), .C1(f[18]), .C2(n342), .A(n434), .ZN(
        n431) );
  AOI221_X1 U158 ( .B1(f8[18]), .B2(n340), .C1(f4[18]), .C2(n341), .A(n433), 
        .ZN(n432) );
  OAI22_X1 U159 ( .A1(n349), .A2(n230), .B1(n350), .B2(n270), .ZN(n434) );
  NAND2_X1 U160 ( .A1(n427), .A2(n428), .ZN(n859) );
  AOI221_X1 U161 ( .B1(f1[19]), .B2(n7), .C1(f[19]), .C2(n342), .A(n430), .ZN(
        n427) );
  AOI221_X1 U162 ( .B1(f8[19]), .B2(n340), .C1(f4[19]), .C2(n341), .A(n429), 
        .ZN(n428) );
  OAI22_X1 U163 ( .A1(n124), .A2(n229), .B1(n350), .B2(n269), .ZN(n430) );
  NAND2_X1 U164 ( .A1(n423), .A2(n424), .ZN(n858) );
  AOI221_X1 U165 ( .B1(f1[20]), .B2(n7), .C1(f[20]), .C2(n342), .A(n426), .ZN(
        n423) );
  AOI221_X1 U166 ( .B1(f8[20]), .B2(n340), .C1(f4[20]), .C2(n341), .A(n425), 
        .ZN(n424) );
  OAI22_X1 U167 ( .A1(n349), .A2(n228), .B1(n350), .B2(n268), .ZN(n426) );
  NAND2_X1 U168 ( .A1(n419), .A2(n420), .ZN(n857) );
  AOI221_X1 U169 ( .B1(f1[21]), .B2(n7), .C1(f[21]), .C2(n342), .A(n422), .ZN(
        n419) );
  AOI221_X1 U170 ( .B1(f8[21]), .B2(n340), .C1(f4[21]), .C2(n341), .A(n421), 
        .ZN(n420) );
  OAI22_X1 U171 ( .A1(n124), .A2(n227), .B1(n350), .B2(n267), .ZN(n422) );
  INV_X1 U172 ( .A(n278), .ZN(n257) );
  INV_X1 U173 ( .A(n277), .ZN(n259) );
  INV_X1 U174 ( .A(n277), .ZN(n260) );
  INV_X1 U175 ( .A(n277), .ZN(n261) );
  INV_X1 U176 ( .A(n277), .ZN(n262) );
  INV_X1 U177 ( .A(n277), .ZN(n263) );
  INV_X1 U178 ( .A(n277), .ZN(n264) );
  INV_X1 U179 ( .A(n276), .ZN(n265) );
  INV_X1 U180 ( .A(n276), .ZN(n266) );
  INV_X1 U181 ( .A(n276), .ZN(n274) );
  INV_X1 U182 ( .A(n276), .ZN(n275) );
  INV_X1 U183 ( .A(n343), .ZN(n354) );
  INV_X1 U184 ( .A(addr_y[0]), .ZN(n361) );
  INV_X1 U185 ( .A(addr_y[1]), .ZN(n362) );
  INV_X1 U186 ( .A(addr_y[2]), .ZN(n365) );
  INV_X1 U187 ( .A(clc1), .ZN(n366) );
  INV_X1 U188 ( .A(clear_acc), .ZN(n1357) );
  OAI21_X1 U189 ( .B1(clear_acc), .B2(n366), .A(n335), .ZN(n828) );
  NAND2_X1 U190 ( .A1(add_r1[39]), .A2(n211), .ZN(n369) );
  NAND2_X1 U191 ( .A1(add_r1[38]), .A2(n218), .ZN(n370) );
  NAND2_X1 U192 ( .A1(add_r1[37]), .A2(n218), .ZN(n373) );
  NAND2_X1 U193 ( .A1(add_r1[36]), .A2(n217), .ZN(n374) );
  NAND2_X1 U194 ( .A1(add_r1[35]), .A2(n218), .ZN(n377) );
  OAI21_X1 U195 ( .B1(n1329), .B2(n279), .A(n377), .ZN(n1194) );
  NAND2_X1 U196 ( .A1(add_r1[34]), .A2(n218), .ZN(n378) );
  NAND2_X1 U197 ( .A1(add_r1[33]), .A2(n218), .ZN(n381) );
  OAI21_X1 U198 ( .B1(n1319), .B2(n279), .A(n381), .ZN(n1192) );
  NAND2_X1 U199 ( .A1(add_r1[32]), .A2(n218), .ZN(n382) );
  OAI21_X1 U200 ( .B1(n1315), .B2(n279), .A(n382), .ZN(n1191) );
  NAND2_X1 U201 ( .A1(add_r1[31]), .A2(n219), .ZN(n385) );
  NAND2_X1 U202 ( .A1(add_r1[30]), .A2(n218), .ZN(n386) );
  OAI21_X1 U203 ( .B1(n1305), .B2(n279), .A(n386), .ZN(n1189) );
  NAND2_X1 U204 ( .A1(add_r1[29]), .A2(n219), .ZN(n389) );
  OAI21_X1 U205 ( .B1(n1300), .B2(n280), .A(n389), .ZN(n1188) );
  NAND2_X1 U206 ( .A1(add_r1[28]), .A2(n218), .ZN(n390) );
  OAI21_X1 U207 ( .B1(n1295), .B2(n280), .A(n390), .ZN(n1187) );
  NAND2_X1 U208 ( .A1(add_r1[27]), .A2(n219), .ZN(n393) );
  OAI21_X1 U209 ( .B1(n1290), .B2(n280), .A(n393), .ZN(n1186) );
  NAND2_X1 U210 ( .A1(add_r1[26]), .A2(n218), .ZN(n394) );
  OAI21_X1 U211 ( .B1(n1285), .B2(n280), .A(n394), .ZN(n1185) );
  NAND2_X1 U212 ( .A1(add_r1[25]), .A2(n219), .ZN(n397) );
  OAI21_X1 U213 ( .B1(n1280), .B2(n280), .A(n397), .ZN(n1184) );
  NAND2_X1 U214 ( .A1(add_r1[24]), .A2(n219), .ZN(n398) );
  OAI21_X1 U215 ( .B1(n1275), .B2(n280), .A(n398), .ZN(n1183) );
  NAND2_X1 U216 ( .A1(add_r1[23]), .A2(n219), .ZN(n401) );
  OAI21_X1 U217 ( .B1(n1270), .B2(n280), .A(n401), .ZN(n1182) );
  NAND2_X1 U218 ( .A1(add_r1[22]), .A2(n219), .ZN(n402) );
  OAI21_X1 U219 ( .B1(n1265), .B2(n280), .A(n402), .ZN(n1181) );
  NAND2_X1 U220 ( .A1(add_r1[21]), .A2(n219), .ZN(n405) );
  OAI21_X1 U221 ( .B1(n27), .B2(n331), .A(n405), .ZN(n1180) );
  NAND2_X1 U222 ( .A1(add_r1[20]), .A2(n217), .ZN(n406) );
  OAI21_X1 U223 ( .B1(n28), .B2(n280), .A(n406), .ZN(n1179) );
  NAND2_X1 U224 ( .A1(add_r1[19]), .A2(n218), .ZN(n409) );
  OAI21_X1 U225 ( .B1(n29), .B2(n287), .A(n409), .ZN(n1178) );
  NAND2_X1 U226 ( .A1(add_r1[18]), .A2(n220), .ZN(n410) );
  OAI21_X1 U227 ( .B1(n30), .B2(n280), .A(n410), .ZN(n1177) );
  NAND2_X1 U228 ( .A1(add_r1[17]), .A2(n217), .ZN(n413) );
  OAI21_X1 U229 ( .B1(n31), .B2(n331), .A(n413), .ZN(n1176) );
  NAND2_X1 U230 ( .A1(add_r1[16]), .A2(n220), .ZN(n414) );
  OAI21_X1 U231 ( .B1(n32), .B2(n280), .A(n414), .ZN(n1175) );
  NAND2_X1 U232 ( .A1(add_r1[15]), .A2(n219), .ZN(n417) );
  OAI21_X1 U233 ( .B1(n33), .B2(n331), .A(n417), .ZN(n1174) );
  NAND2_X1 U234 ( .A1(add_r1[13]), .A2(n220), .ZN(n418) );
  OAI21_X1 U235 ( .B1(n835), .B2(n331), .A(n418), .ZN(n1172) );
  NAND2_X1 U236 ( .A1(add_r1[12]), .A2(n218), .ZN(n447) );
  OAI21_X1 U237 ( .B1(n1200), .B2(n331), .A(n447), .ZN(n1171) );
  NAND2_X1 U238 ( .A1(add_r1[11]), .A2(n220), .ZN(n448) );
  OAI21_X1 U239 ( .B1(n1205), .B2(n331), .A(n448), .ZN(n1170) );
  NAND2_X1 U240 ( .A1(add_r1[10]), .A2(n219), .ZN(n449) );
  OAI21_X1 U241 ( .B1(n1210), .B2(n331), .A(n449), .ZN(n1169) );
  NAND2_X1 U242 ( .A1(add_r1[9]), .A2(n220), .ZN(n450) );
  OAI21_X1 U243 ( .B1(n1215), .B2(n331), .A(n450), .ZN(n1168) );
  NAND2_X1 U244 ( .A1(add_r1[8]), .A2(n219), .ZN(n451) );
  OAI21_X1 U245 ( .B1(n1220), .B2(n331), .A(n451), .ZN(n1167) );
  NAND2_X1 U246 ( .A1(add_r1[7]), .A2(n220), .ZN(n452) );
  OAI21_X1 U247 ( .B1(n1225), .B2(n288), .A(n452), .ZN(n1166) );
  NAND2_X1 U248 ( .A1(add_r1[6]), .A2(n218), .ZN(n453) );
  OAI21_X1 U249 ( .B1(n1230), .B2(n331), .A(n453), .ZN(n1165) );
  NAND2_X1 U250 ( .A1(add_r1[5]), .A2(n220), .ZN(n454) );
  OAI21_X1 U251 ( .B1(n1235), .B2(n331), .A(n454), .ZN(n1164) );
  NAND2_X1 U252 ( .A1(add_r1[4]), .A2(n220), .ZN(n455) );
  OAI21_X1 U253 ( .B1(n1240), .B2(n284), .A(n455), .ZN(n1163) );
  NAND2_X1 U254 ( .A1(add_r1[3]), .A2(n220), .ZN(n456) );
  OAI21_X1 U255 ( .B1(n1245), .B2(n329), .A(n456), .ZN(n1162) );
  NAND2_X1 U256 ( .A1(add_r1[2]), .A2(n220), .ZN(n457) );
  OAI21_X1 U257 ( .B1(n1250), .B2(n331), .A(n457), .ZN(n1161) );
  NAND2_X1 U258 ( .A1(add_r1[1]), .A2(n219), .ZN(n458) );
  OAI21_X1 U259 ( .B1(n1255), .B2(n329), .A(n458), .ZN(n1160) );
  NAND2_X1 U260 ( .A1(add_r1[0]), .A2(n220), .ZN(n459) );
  OAI21_X1 U261 ( .B1(n1260), .B2(n281), .A(n459), .ZN(n1159) );
  NAND2_X1 U262 ( .A1(add_r1[14]), .A2(n220), .ZN(n460) );
  OAI21_X1 U263 ( .B1(n830), .B2(n281), .A(n460), .ZN(n1173) );
  AOI22_X1 U264 ( .A1(n257), .A2(n1355), .B1(add_r6[39]), .B2(n222), .ZN(n461)
         );
  INV_X1 U265 ( .A(n461), .ZN(n998) );
  AOI22_X1 U266 ( .A1(n257), .A2(n1347), .B1(add_r6[38]), .B2(n255), .ZN(n462)
         );
  INV_X1 U267 ( .A(n462), .ZN(n997) );
  AOI22_X1 U268 ( .A1(n257), .A2(n1342), .B1(add_r6[37]), .B2(n251), .ZN(n463)
         );
  INV_X1 U269 ( .A(n463), .ZN(n996) );
  AOI22_X1 U270 ( .A1(n257), .A2(n1337), .B1(add_r6[36]), .B2(n251), .ZN(n464)
         );
  INV_X1 U271 ( .A(n464), .ZN(n995) );
  AOI22_X1 U272 ( .A1(n257), .A2(n1332), .B1(add_r6[35]), .B2(n251), .ZN(n465)
         );
  INV_X1 U273 ( .A(n465), .ZN(n994) );
  AOI22_X1 U274 ( .A1(n257), .A2(n1327), .B1(add_r6[34]), .B2(n251), .ZN(n466)
         );
  INV_X1 U275 ( .A(n466), .ZN(n993) );
  AOI22_X1 U276 ( .A1(n257), .A2(n1322), .B1(add_r6[33]), .B2(n251), .ZN(n467)
         );
  INV_X1 U277 ( .A(n467), .ZN(n992) );
  AOI22_X1 U278 ( .A1(n257), .A2(n1317), .B1(add_r6[32]), .B2(n251), .ZN(n468)
         );
  INV_X1 U279 ( .A(n468), .ZN(n991) );
  AOI22_X1 U280 ( .A1(n257), .A2(n1313), .B1(add_r6[31]), .B2(n251), .ZN(n469)
         );
  INV_X1 U281 ( .A(n469), .ZN(n990) );
  AOI22_X1 U282 ( .A1(n257), .A2(n1308), .B1(add_r6[30]), .B2(n252), .ZN(n470)
         );
  INV_X1 U283 ( .A(n470), .ZN(n989) );
  AOI22_X1 U284 ( .A1(n257), .A2(n1303), .B1(add_r6[29]), .B2(n252), .ZN(n471)
         );
  INV_X1 U285 ( .A(n471), .ZN(n988) );
  AOI22_X1 U286 ( .A1(n257), .A2(n1298), .B1(add_r6[28]), .B2(n252), .ZN(n472)
         );
  INV_X1 U287 ( .A(n472), .ZN(n987) );
  AOI22_X1 U288 ( .A1(n258), .A2(n1293), .B1(add_r6[27]), .B2(n252), .ZN(n473)
         );
  INV_X1 U289 ( .A(n473), .ZN(n986) );
  AOI22_X1 U290 ( .A1(n258), .A2(n1288), .B1(add_r6[26]), .B2(n252), .ZN(n474)
         );
  INV_X1 U291 ( .A(n474), .ZN(n985) );
  AOI22_X1 U292 ( .A1(n258), .A2(n1283), .B1(add_r6[25]), .B2(n252), .ZN(n475)
         );
  INV_X1 U293 ( .A(n475), .ZN(n984) );
  AOI22_X1 U294 ( .A1(n258), .A2(n1278), .B1(add_r6[24]), .B2(n252), .ZN(n476)
         );
  INV_X1 U295 ( .A(n476), .ZN(n983) );
  AOI22_X1 U296 ( .A1(n258), .A2(n1273), .B1(add_r6[23]), .B2(n252), .ZN(n477)
         );
  INV_X1 U297 ( .A(n477), .ZN(n982) );
  AOI22_X1 U298 ( .A1(n258), .A2(n1268), .B1(add_r6[22]), .B2(n252), .ZN(n478)
         );
  INV_X1 U299 ( .A(n478), .ZN(n981) );
  AOI22_X1 U300 ( .A1(n258), .A2(n479), .B1(add_r6[21]), .B2(n252), .ZN(n480)
         );
  INV_X1 U301 ( .A(n480), .ZN(n980) );
  AOI22_X1 U302 ( .A1(n258), .A2(n481), .B1(add_r6[20]), .B2(n252), .ZN(n482)
         );
  INV_X1 U303 ( .A(n482), .ZN(n979) );
  AOI22_X1 U304 ( .A1(n258), .A2(n483), .B1(add_r6[19]), .B2(n252), .ZN(n484)
         );
  INV_X1 U305 ( .A(n484), .ZN(n978) );
  AOI22_X1 U306 ( .A1(n258), .A2(n485), .B1(add_r6[18]), .B2(n253), .ZN(n486)
         );
  INV_X1 U307 ( .A(n486), .ZN(n977) );
  AOI22_X1 U308 ( .A1(n258), .A2(n487), .B1(add_r6[17]), .B2(n253), .ZN(n488)
         );
  INV_X1 U309 ( .A(n488), .ZN(n976) );
  AOI22_X1 U310 ( .A1(n258), .A2(f6[16]), .B1(add_r6[16]), .B2(n253), .ZN(n489) );
  INV_X1 U311 ( .A(n489), .ZN(n975) );
  AOI22_X1 U312 ( .A1(n257), .A2(f6[15]), .B1(add_r6[15]), .B2(n253), .ZN(n490) );
  INV_X1 U313 ( .A(n490), .ZN(n974) );
  AOI22_X1 U314 ( .A1(n258), .A2(f6[13]), .B1(add_r6[13]), .B2(n253), .ZN(n491) );
  INV_X1 U315 ( .A(n491), .ZN(n972) );
  AOI22_X1 U316 ( .A1(n265), .A2(f6[12]), .B1(add_r6[12]), .B2(n253), .ZN(n492) );
  INV_X1 U317 ( .A(n492), .ZN(n971) );
  AOI22_X1 U318 ( .A1(n275), .A2(f6[11]), .B1(add_r6[11]), .B2(n253), .ZN(n493) );
  INV_X1 U319 ( .A(n493), .ZN(n970) );
  AOI22_X1 U320 ( .A1(n274), .A2(f6[10]), .B1(add_r6[10]), .B2(n253), .ZN(n494) );
  INV_X1 U321 ( .A(n494), .ZN(n969) );
  AOI22_X1 U322 ( .A1(n266), .A2(f6[9]), .B1(add_r6[9]), .B2(n253), .ZN(n495)
         );
  INV_X1 U323 ( .A(n495), .ZN(n968) );
  AOI22_X1 U324 ( .A1(n265), .A2(f6[8]), .B1(add_r6[8]), .B2(n253), .ZN(n496)
         );
  INV_X1 U325 ( .A(n496), .ZN(n967) );
  AOI22_X1 U326 ( .A1(n265), .A2(f6[7]), .B1(add_r6[7]), .B2(n253), .ZN(n497)
         );
  INV_X1 U327 ( .A(n497), .ZN(n966) );
  AOI22_X1 U328 ( .A1(n257), .A2(f6[6]), .B1(add_r6[6]), .B2(n253), .ZN(n498)
         );
  INV_X1 U329 ( .A(n498), .ZN(n965) );
  AOI22_X1 U330 ( .A1(n258), .A2(f6[5]), .B1(add_r6[5]), .B2(n254), .ZN(n499)
         );
  INV_X1 U331 ( .A(n499), .ZN(n964) );
  AOI22_X1 U332 ( .A1(n257), .A2(f6[4]), .B1(add_r6[4]), .B2(n254), .ZN(n500)
         );
  INV_X1 U333 ( .A(n500), .ZN(n963) );
  AOI22_X1 U334 ( .A1(n258), .A2(f6[3]), .B1(add_r6[3]), .B2(n254), .ZN(n501)
         );
  INV_X1 U335 ( .A(n501), .ZN(n962) );
  AOI22_X1 U336 ( .A1(n259), .A2(f6[2]), .B1(add_r6[2]), .B2(n254), .ZN(n502)
         );
  INV_X1 U337 ( .A(n502), .ZN(n961) );
  AOI22_X1 U338 ( .A1(n259), .A2(f6[1]), .B1(add_r6[1]), .B2(n254), .ZN(n503)
         );
  INV_X1 U339 ( .A(n503), .ZN(n960) );
  AOI22_X1 U340 ( .A1(n259), .A2(f6[0]), .B1(add_r6[0]), .B2(n254), .ZN(n504)
         );
  INV_X1 U341 ( .A(n504), .ZN(n959) );
  AOI22_X1 U342 ( .A1(n259), .A2(f6[14]), .B1(add_r6[14]), .B2(n254), .ZN(n505) );
  INV_X1 U343 ( .A(n505), .ZN(n973) );
  AOI22_X1 U344 ( .A1(n259), .A2(n1353), .B1(add_r7[39]), .B2(n254), .ZN(n514)
         );
  INV_X1 U345 ( .A(n514), .ZN(n958) );
  AOI22_X1 U346 ( .A1(n259), .A2(n1346), .B1(add_r7[38]), .B2(n254), .ZN(n517)
         );
  INV_X1 U347 ( .A(n517), .ZN(n957) );
  AOI22_X1 U348 ( .A1(n259), .A2(n1341), .B1(add_r7[37]), .B2(n254), .ZN(n518)
         );
  INV_X1 U349 ( .A(n518), .ZN(n956) );
  AOI22_X1 U350 ( .A1(n259), .A2(n1336), .B1(add_r7[36]), .B2(n254), .ZN(n519)
         );
  INV_X1 U351 ( .A(n519), .ZN(n955) );
  AOI22_X1 U352 ( .A1(n259), .A2(n1331), .B1(add_r7[35]), .B2(n254), .ZN(n520)
         );
  INV_X1 U353 ( .A(n520), .ZN(n954) );
  AOI22_X1 U354 ( .A1(n259), .A2(n1326), .B1(add_r7[34]), .B2(n255), .ZN(n521)
         );
  INV_X1 U355 ( .A(n521), .ZN(n953) );
  AOI22_X1 U356 ( .A1(n259), .A2(n1321), .B1(add_r7[33]), .B2(n255), .ZN(n522)
         );
  INV_X1 U357 ( .A(n522), .ZN(n952) );
  AOI22_X1 U358 ( .A1(n259), .A2(f7[32]), .B1(add_r7[32]), .B2(n255), .ZN(n523) );
  INV_X1 U359 ( .A(n523), .ZN(n951) );
  AOI22_X1 U360 ( .A1(n260), .A2(n1312), .B1(add_r7[31]), .B2(n255), .ZN(n524)
         );
  INV_X1 U361 ( .A(n524), .ZN(n950) );
  AOI22_X1 U362 ( .A1(n260), .A2(n1307), .B1(add_r7[30]), .B2(n255), .ZN(n525)
         );
  INV_X1 U363 ( .A(n525), .ZN(n949) );
  AOI22_X1 U364 ( .A1(n260), .A2(n1302), .B1(add_r7[29]), .B2(n255), .ZN(n526)
         );
  INV_X1 U365 ( .A(n526), .ZN(n948) );
  AOI22_X1 U366 ( .A1(n260), .A2(n1297), .B1(add_r7[28]), .B2(n255), .ZN(n527)
         );
  INV_X1 U367 ( .A(n527), .ZN(n947) );
  AOI22_X1 U368 ( .A1(n260), .A2(n1292), .B1(add_r7[27]), .B2(n255), .ZN(n528)
         );
  INV_X1 U369 ( .A(n528), .ZN(n946) );
  AOI22_X1 U370 ( .A1(n260), .A2(n1287), .B1(add_r7[26]), .B2(n255), .ZN(n529)
         );
  INV_X1 U371 ( .A(n529), .ZN(n945) );
  AOI22_X1 U372 ( .A1(n260), .A2(n1282), .B1(add_r7[25]), .B2(n255), .ZN(n530)
         );
  INV_X1 U373 ( .A(n530), .ZN(n944) );
  AOI22_X1 U374 ( .A1(n260), .A2(n1277), .B1(add_r7[24]), .B2(n255), .ZN(n531)
         );
  INV_X1 U375 ( .A(n531), .ZN(n943) );
  AOI22_X1 U376 ( .A1(n260), .A2(n1272), .B1(add_r7[23]), .B2(n256), .ZN(n532)
         );
  INV_X1 U377 ( .A(n532), .ZN(n942) );
  AOI22_X1 U378 ( .A1(n260), .A2(n1267), .B1(add_r7[22]), .B2(n256), .ZN(n533)
         );
  INV_X1 U379 ( .A(n533), .ZN(n941) );
  AOI22_X1 U380 ( .A1(n260), .A2(n534), .B1(add_r7[21]), .B2(n256), .ZN(n535)
         );
  INV_X1 U381 ( .A(n535), .ZN(n940) );
  AOI22_X1 U382 ( .A1(n260), .A2(n536), .B1(add_r7[20]), .B2(n256), .ZN(n537)
         );
  INV_X1 U383 ( .A(n537), .ZN(n939) );
  AOI22_X1 U384 ( .A1(n261), .A2(n538), .B1(add_r7[19]), .B2(n256), .ZN(n539)
         );
  INV_X1 U385 ( .A(n539), .ZN(n938) );
  AOI22_X1 U386 ( .A1(n261), .A2(n540), .B1(add_r7[18]), .B2(n256), .ZN(n541)
         );
  INV_X1 U387 ( .A(n541), .ZN(n937) );
  AOI22_X1 U388 ( .A1(n261), .A2(n542), .B1(add_r7[17]), .B2(n256), .ZN(n543)
         );
  INV_X1 U389 ( .A(n543), .ZN(n936) );
  AOI22_X1 U390 ( .A1(n261), .A2(f7[16]), .B1(add_r7[16]), .B2(n256), .ZN(n544) );
  INV_X1 U391 ( .A(n544), .ZN(n935) );
  AOI22_X1 U392 ( .A1(n261), .A2(n545), .B1(add_r7[15]), .B2(n256), .ZN(n546)
         );
  INV_X1 U393 ( .A(n546), .ZN(n934) );
  AOI22_X1 U394 ( .A1(n261), .A2(f7[13]), .B1(add_r7[13]), .B2(n256), .ZN(n547) );
  INV_X1 U395 ( .A(n547), .ZN(n932) );
  AOI22_X1 U396 ( .A1(n261), .A2(f7[12]), .B1(add_r7[12]), .B2(n256), .ZN(n548) );
  INV_X1 U397 ( .A(n548), .ZN(n931) );
  AOI22_X1 U398 ( .A1(n261), .A2(f7[11]), .B1(add_r7[11]), .B2(n256), .ZN(n549) );
  INV_X1 U399 ( .A(n549), .ZN(n930) );
  AOI22_X1 U400 ( .A1(n261), .A2(f7[10]), .B1(add_r7[10]), .B2(n8), .ZN(n550)
         );
  INV_X1 U401 ( .A(n550), .ZN(n929) );
  AOI22_X1 U402 ( .A1(n261), .A2(f7[9]), .B1(add_r7[9]), .B2(n8), .ZN(n551) );
  INV_X1 U403 ( .A(n551), .ZN(n928) );
  AOI22_X1 U404 ( .A1(n261), .A2(f7[8]), .B1(add_r7[8]), .B2(n209), .ZN(n552)
         );
  INV_X1 U405 ( .A(n552), .ZN(n927) );
  AOI22_X1 U406 ( .A1(n261), .A2(f7[7]), .B1(add_r7[7]), .B2(n126), .ZN(n553)
         );
  INV_X1 U407 ( .A(n553), .ZN(n926) );
  AOI22_X1 U408 ( .A1(n262), .A2(f7[6]), .B1(add_r7[6]), .B2(n210), .ZN(n554)
         );
  INV_X1 U409 ( .A(n554), .ZN(n925) );
  AOI22_X1 U410 ( .A1(n262), .A2(f7[5]), .B1(add_r7[5]), .B2(n8), .ZN(n555) );
  INV_X1 U411 ( .A(n555), .ZN(n924) );
  AOI22_X1 U412 ( .A1(n262), .A2(f7[4]), .B1(add_r7[4]), .B2(n8), .ZN(n556) );
  INV_X1 U413 ( .A(n556), .ZN(n923) );
  AOI22_X1 U414 ( .A1(n262), .A2(f7[3]), .B1(add_r7[3]), .B2(n8), .ZN(n557) );
  INV_X1 U415 ( .A(n557), .ZN(n922) );
  AOI22_X1 U416 ( .A1(n262), .A2(f7[2]), .B1(add_r7[2]), .B2(n8), .ZN(n558) );
  INV_X1 U417 ( .A(n558), .ZN(n921) );
  AOI22_X1 U418 ( .A1(n262), .A2(f7[1]), .B1(add_r7[1]), .B2(n8), .ZN(n559) );
  INV_X1 U419 ( .A(n559), .ZN(n920) );
  AOI22_X1 U420 ( .A1(n262), .A2(f7[0]), .B1(add_r7[0]), .B2(n8), .ZN(n560) );
  INV_X1 U421 ( .A(n560), .ZN(n919) );
  AOI22_X1 U422 ( .A1(n262), .A2(f7[14]), .B1(add_r7[14]), .B2(n8), .ZN(n561)
         );
  INV_X1 U423 ( .A(n561), .ZN(n933) );
  NAND2_X1 U424 ( .A1(add_r8[39]), .A2(n217), .ZN(n562) );
  OAI21_X1 U425 ( .B1(n289), .B2(n281), .A(n562), .ZN(n918) );
  NAND2_X1 U426 ( .A1(add_r8[38]), .A2(n217), .ZN(n563) );
  NAND2_X1 U427 ( .A1(add_r8[37]), .A2(n217), .ZN(n564) );
  NAND2_X1 U428 ( .A1(add_r8[36]), .A2(n217), .ZN(n565) );
  NAND2_X1 U429 ( .A1(add_r8[35]), .A2(n217), .ZN(n566) );
  NAND2_X1 U430 ( .A1(add_r8[34]), .A2(n217), .ZN(n567) );
  NAND2_X1 U431 ( .A1(add_r8[33]), .A2(n217), .ZN(n568) );
  NAND2_X1 U432 ( .A1(add_r8[32]), .A2(n217), .ZN(n569) );
  OAI21_X1 U433 ( .B1(n296), .B2(n282), .A(n569), .ZN(n911) );
  NAND2_X1 U434 ( .A1(add_r8[31]), .A2(n216), .ZN(n570) );
  OAI21_X1 U435 ( .B1(n297), .B2(n282), .A(n570), .ZN(n910) );
  NAND2_X1 U436 ( .A1(add_r8[30]), .A2(n216), .ZN(n571) );
  OAI21_X1 U437 ( .B1(n298), .B2(n282), .A(n571), .ZN(n909) );
  NAND2_X1 U438 ( .A1(add_r8[29]), .A2(n216), .ZN(n572) );
  OAI21_X1 U439 ( .B1(n299), .B2(n282), .A(n572), .ZN(n908) );
  NAND2_X1 U440 ( .A1(add_r8[28]), .A2(n216), .ZN(n573) );
  OAI21_X1 U441 ( .B1(n300), .B2(n282), .A(n573), .ZN(n907) );
  NAND2_X1 U442 ( .A1(add_r8[27]), .A2(n216), .ZN(n574) );
  OAI21_X1 U443 ( .B1(n301), .B2(n288), .A(n574), .ZN(n906) );
  NAND2_X1 U444 ( .A1(add_r8[26]), .A2(n216), .ZN(n575) );
  OAI21_X1 U445 ( .B1(n302), .B2(n331), .A(n575), .ZN(n905) );
  NAND2_X1 U446 ( .A1(add_r8[25]), .A2(n216), .ZN(n576) );
  OAI21_X1 U447 ( .B1(n303), .B2(n279), .A(n576), .ZN(n904) );
  NAND2_X1 U448 ( .A1(add_r8[24]), .A2(n216), .ZN(n577) );
  OAI21_X1 U449 ( .B1(n304), .B2(n331), .A(n577), .ZN(n903) );
  NAND2_X1 U450 ( .A1(add_r8[23]), .A2(n216), .ZN(n578) );
  OAI21_X1 U451 ( .B1(n305), .B2(n331), .A(n578), .ZN(n902) );
  NAND2_X1 U452 ( .A1(add_r8[22]), .A2(n216), .ZN(n579) );
  OAI21_X1 U453 ( .B1(n306), .B2(n331), .A(n579), .ZN(n901) );
  NAND2_X1 U454 ( .A1(add_r8[21]), .A2(n216), .ZN(n580) );
  OAI21_X1 U455 ( .B1(n307), .B2(n331), .A(n580), .ZN(n900) );
  NAND2_X1 U456 ( .A1(add_r8[20]), .A2(n216), .ZN(n581) );
  OAI21_X1 U457 ( .B1(n308), .B2(n283), .A(n581), .ZN(n899) );
  NAND2_X1 U458 ( .A1(add_r8[19]), .A2(n215), .ZN(n582) );
  OAI21_X1 U459 ( .B1(n309), .B2(n283), .A(n582), .ZN(n898) );
  NAND2_X1 U460 ( .A1(add_r8[18]), .A2(n215), .ZN(n583) );
  OAI21_X1 U461 ( .B1(n310), .B2(n283), .A(n583), .ZN(n897) );
  NAND2_X1 U462 ( .A1(add_r8[17]), .A2(n215), .ZN(n584) );
  OAI21_X1 U463 ( .B1(n311), .B2(n283), .A(n584), .ZN(n896) );
  NAND2_X1 U464 ( .A1(add_r8[16]), .A2(n215), .ZN(n585) );
  OAI21_X1 U465 ( .B1(n312), .B2(n283), .A(n585), .ZN(n895) );
  NAND2_X1 U466 ( .A1(add_r8[15]), .A2(n215), .ZN(n586) );
  OAI21_X1 U467 ( .B1(n313), .B2(n283), .A(n586), .ZN(n894) );
  NAND2_X1 U468 ( .A1(add_r8[13]), .A2(n215), .ZN(n587) );
  OAI21_X1 U469 ( .B1(n315), .B2(n283), .A(n587), .ZN(n892) );
  NAND2_X1 U470 ( .A1(add_r8[12]), .A2(n215), .ZN(n588) );
  OAI21_X1 U471 ( .B1(n316), .B2(n284), .A(n588), .ZN(n891) );
  NAND2_X1 U472 ( .A1(add_r8[11]), .A2(n215), .ZN(n589) );
  OAI21_X1 U473 ( .B1(n317), .B2(n284), .A(n589), .ZN(n890) );
  NAND2_X1 U474 ( .A1(add_r8[10]), .A2(n215), .ZN(n590) );
  OAI21_X1 U475 ( .B1(n318), .B2(n284), .A(n590), .ZN(n889) );
  NAND2_X1 U476 ( .A1(add_r8[9]), .A2(n215), .ZN(n591) );
  OAI21_X1 U477 ( .B1(n319), .B2(n284), .A(n591), .ZN(n888) );
  NAND2_X1 U478 ( .A1(add_r8[8]), .A2(n215), .ZN(n592) );
  OAI21_X1 U479 ( .B1(n320), .B2(n284), .A(n592), .ZN(n887) );
  NAND2_X1 U480 ( .A1(add_r8[7]), .A2(n215), .ZN(n593) );
  OAI21_X1 U481 ( .B1(n321), .B2(n284), .A(n593), .ZN(n886) );
  NAND2_X1 U482 ( .A1(add_r8[6]), .A2(n214), .ZN(n594) );
  OAI21_X1 U483 ( .B1(n322), .B2(n284), .A(n594), .ZN(n885) );
  NAND2_X1 U484 ( .A1(add_r8[5]), .A2(n214), .ZN(n595) );
  OAI21_X1 U485 ( .B1(n323), .B2(n285), .A(n595), .ZN(n884) );
  NAND2_X1 U486 ( .A1(add_r8[4]), .A2(n214), .ZN(n596) );
  OAI21_X1 U487 ( .B1(n324), .B2(n285), .A(n596), .ZN(n883) );
  NAND2_X1 U488 ( .A1(add_r8[3]), .A2(n214), .ZN(n597) );
  OAI21_X1 U489 ( .B1(n325), .B2(n285), .A(n597), .ZN(n882) );
  NAND2_X1 U490 ( .A1(add_r8[2]), .A2(n214), .ZN(n598) );
  OAI21_X1 U491 ( .B1(n326), .B2(n285), .A(n598), .ZN(n881) );
  NAND2_X1 U492 ( .A1(add_r8[1]), .A2(n214), .ZN(n599) );
  OAI21_X1 U493 ( .B1(n327), .B2(n285), .A(n599), .ZN(n880) );
  NAND2_X1 U494 ( .A1(add_r8[0]), .A2(n214), .ZN(n600) );
  OAI21_X1 U495 ( .B1(n328), .B2(n285), .A(n600), .ZN(n879) );
  NAND2_X1 U496 ( .A1(add_r8[14]), .A2(n214), .ZN(n601) );
  OAI21_X1 U497 ( .B1(n314), .B2(n285), .A(n601), .ZN(n893) );
  NAND2_X1 U498 ( .A1(add_r4[39]), .A2(n214), .ZN(n602) );
  OAI21_X1 U499 ( .B1(n129), .B2(n286), .A(n602), .ZN(n1078) );
  NAND2_X1 U500 ( .A1(add_r4[38]), .A2(n214), .ZN(n603) );
  NAND2_X1 U501 ( .A1(add_r4[37]), .A2(n214), .ZN(n604) );
  OAI21_X1 U502 ( .B1(n131), .B2(n286), .A(n604), .ZN(n1076) );
  NAND2_X1 U503 ( .A1(add_r4[36]), .A2(n214), .ZN(n605) );
  NAND2_X1 U504 ( .A1(add_r4[35]), .A2(n213), .ZN(n606) );
  OAI21_X1 U505 ( .B1(n133), .B2(n286), .A(n606), .ZN(n1074) );
  NAND2_X1 U506 ( .A1(add_r4[34]), .A2(n217), .ZN(n607) );
  OAI21_X1 U507 ( .B1(n134), .B2(n286), .A(n607), .ZN(n1073) );
  NAND2_X1 U508 ( .A1(add_r4[33]), .A2(n213), .ZN(n608) );
  OAI21_X1 U509 ( .B1(n135), .B2(n286), .A(n608), .ZN(n1072) );
  NAND2_X1 U510 ( .A1(add_r4[32]), .A2(n213), .ZN(n609) );
  OAI21_X1 U511 ( .B1(n136), .B2(n287), .A(n609), .ZN(n1071) );
  NAND2_X1 U512 ( .A1(add_r4[31]), .A2(n213), .ZN(n610) );
  OAI21_X1 U513 ( .B1(n137), .B2(n287), .A(n610), .ZN(n1070) );
  NAND2_X1 U514 ( .A1(add_r4[30]), .A2(n213), .ZN(n611) );
  OAI21_X1 U515 ( .B1(n138), .B2(n287), .A(n611), .ZN(n1069) );
  NAND2_X1 U516 ( .A1(add_r4[29]), .A2(n213), .ZN(n612) );
  OAI21_X1 U517 ( .B1(n139), .B2(n287), .A(n612), .ZN(n1068) );
  NAND2_X1 U518 ( .A1(add_r4[28]), .A2(n213), .ZN(n613) );
  OAI21_X1 U519 ( .B1(n140), .B2(n287), .A(n613), .ZN(n1067) );
  NAND2_X1 U520 ( .A1(add_r4[27]), .A2(n213), .ZN(n614) );
  OAI21_X1 U521 ( .B1(n141), .B2(n287), .A(n614), .ZN(n1066) );
  NAND2_X1 U522 ( .A1(add_r4[26]), .A2(n213), .ZN(n615) );
  OAI21_X1 U523 ( .B1(n142), .B2(n287), .A(n615), .ZN(n1065) );
  NAND2_X1 U524 ( .A1(add_r4[25]), .A2(n213), .ZN(n616) );
  OAI21_X1 U525 ( .B1(n143), .B2(n288), .A(n616), .ZN(n1064) );
  NAND2_X1 U526 ( .A1(add_r4[24]), .A2(n213), .ZN(n617) );
  OAI21_X1 U527 ( .B1(n144), .B2(n288), .A(n617), .ZN(n1063) );
  NAND2_X1 U528 ( .A1(add_r4[23]), .A2(n213), .ZN(n618) );
  OAI21_X1 U529 ( .B1(n145), .B2(n288), .A(n618), .ZN(n1062) );
  NAND2_X1 U530 ( .A1(add_r4[22]), .A2(n212), .ZN(n619) );
  OAI21_X1 U531 ( .B1(n146), .B2(n288), .A(n619), .ZN(n1061) );
  NAND2_X1 U532 ( .A1(add_r4[21]), .A2(n212), .ZN(n620) );
  OAI21_X1 U533 ( .B1(n147), .B2(n288), .A(n620), .ZN(n1060) );
  NAND2_X1 U534 ( .A1(add_r4[20]), .A2(n212), .ZN(n621) );
  OAI21_X1 U535 ( .B1(n148), .B2(n288), .A(n621), .ZN(n1059) );
  NAND2_X1 U536 ( .A1(add_r4[19]), .A2(n212), .ZN(n622) );
  OAI21_X1 U537 ( .B1(n149), .B2(n288), .A(n622), .ZN(n1058) );
  NAND2_X1 U538 ( .A1(add_r4[18]), .A2(n212), .ZN(n623) );
  OAI21_X1 U539 ( .B1(n150), .B2(n329), .A(n623), .ZN(n1057) );
  NAND2_X1 U540 ( .A1(add_r4[17]), .A2(n212), .ZN(n624) );
  OAI21_X1 U541 ( .B1(n151), .B2(n329), .A(n624), .ZN(n1056) );
  NAND2_X1 U542 ( .A1(add_r4[16]), .A2(n212), .ZN(n625) );
  OAI21_X1 U543 ( .B1(n152), .B2(n287), .A(n625), .ZN(n1055) );
  NAND2_X1 U544 ( .A1(add_r4[15]), .A2(n212), .ZN(n626) );
  OAI21_X1 U545 ( .B1(n153), .B2(n287), .A(n626), .ZN(n1054) );
  NAND2_X1 U546 ( .A1(add_r4[13]), .A2(n212), .ZN(n627) );
  OAI21_X1 U547 ( .B1(n155), .B2(n288), .A(n627), .ZN(n1052) );
  NAND2_X1 U548 ( .A1(add_r4[12]), .A2(n212), .ZN(n628) );
  OAI21_X1 U549 ( .B1(n156), .B2(n280), .A(n628), .ZN(n1051) );
  NAND2_X1 U550 ( .A1(add_r4[11]), .A2(n212), .ZN(n629) );
  OAI21_X1 U551 ( .B1(n157), .B2(n280), .A(n629), .ZN(n1050) );
  NAND2_X1 U552 ( .A1(add_r4[10]), .A2(n212), .ZN(n630) );
  OAI21_X1 U553 ( .B1(n158), .B2(n329), .A(n630), .ZN(n1049) );
  NAND2_X1 U554 ( .A1(add_r4[9]), .A2(n211), .ZN(n631) );
  OAI21_X1 U555 ( .B1(n159), .B2(n331), .A(n631), .ZN(n1048) );
  NAND2_X1 U556 ( .A1(add_r4[8]), .A2(n211), .ZN(n632) );
  OAI21_X1 U557 ( .B1(n160), .B2(n288), .A(n632), .ZN(n1047) );
  NAND2_X1 U558 ( .A1(add_r4[7]), .A2(n211), .ZN(n633) );
  OAI21_X1 U559 ( .B1(n161), .B2(n287), .A(n633), .ZN(n1046) );
  NAND2_X1 U560 ( .A1(add_r4[6]), .A2(n211), .ZN(n634) );
  OAI21_X1 U561 ( .B1(n162), .B2(n329), .A(n634), .ZN(n1045) );
  NAND2_X1 U562 ( .A1(add_r4[5]), .A2(n211), .ZN(n635) );
  OAI21_X1 U563 ( .B1(n163), .B2(n329), .A(n635), .ZN(n1044) );
  NAND2_X1 U564 ( .A1(add_r4[4]), .A2(n211), .ZN(n636) );
  OAI21_X1 U565 ( .B1(n164), .B2(n288), .A(n636), .ZN(n1043) );
  NAND2_X1 U566 ( .A1(add_r4[3]), .A2(n211), .ZN(n637) );
  OAI21_X1 U567 ( .B1(n165), .B2(n329), .A(n637), .ZN(n1042) );
  NAND2_X1 U568 ( .A1(add_r4[2]), .A2(n211), .ZN(n638) );
  OAI21_X1 U569 ( .B1(n166), .B2(n329), .A(n638), .ZN(n1041) );
  NAND2_X1 U570 ( .A1(add_r4[1]), .A2(n211), .ZN(n639) );
  OAI21_X1 U571 ( .B1(n167), .B2(n329), .A(n639), .ZN(n1040) );
  NAND2_X1 U572 ( .A1(add_r4[0]), .A2(n211), .ZN(n640) );
  OAI21_X1 U573 ( .B1(n168), .B2(n329), .A(n640), .ZN(n1039) );
  NAND2_X1 U574 ( .A1(add_r4[14]), .A2(n211), .ZN(n641) );
  OAI21_X1 U575 ( .B1(n154), .B2(n329), .A(n641), .ZN(n1053) );
  AOI22_X1 U576 ( .A1(n262), .A2(n642), .B1(add_r3[39]), .B2(n8), .ZN(n643) );
  INV_X1 U577 ( .A(n643), .ZN(n1118) );
  AOI22_X1 U578 ( .A1(n262), .A2(n644), .B1(add_r3[38]), .B2(n8), .ZN(n645) );
  INV_X1 U579 ( .A(n645), .ZN(n1117) );
  AOI22_X1 U580 ( .A1(n262), .A2(n647), .B1(add_r3[36]), .B2(n8), .ZN(n648) );
  INV_X1 U581 ( .A(n648), .ZN(n1115) );
  AOI22_X1 U582 ( .A1(n263), .A2(n650), .B1(add_r3[34]), .B2(n210), .ZN(n651)
         );
  INV_X1 U583 ( .A(n651), .ZN(n1113) );
  AOI22_X1 U584 ( .A1(n263), .A2(n652), .B1(add_r3[33]), .B2(n209), .ZN(n653)
         );
  INV_X1 U585 ( .A(n653), .ZN(n1112) );
  AOI22_X1 U586 ( .A1(n263), .A2(n654), .B1(add_r3[32]), .B2(n8), .ZN(n655) );
  INV_X1 U587 ( .A(n655), .ZN(n1111) );
  AOI22_X1 U588 ( .A1(n263), .A2(n656), .B1(add_r3[31]), .B2(n8), .ZN(n657) );
  INV_X1 U589 ( .A(n657), .ZN(n1110) );
  AOI22_X1 U590 ( .A1(n263), .A2(n658), .B1(add_r3[30]), .B2(n210), .ZN(n659)
         );
  INV_X1 U591 ( .A(n659), .ZN(n1109) );
  AOI22_X1 U592 ( .A1(n263), .A2(n660), .B1(add_r3[29]), .B2(n8), .ZN(n661) );
  INV_X1 U593 ( .A(n661), .ZN(n1108) );
  AOI22_X1 U594 ( .A1(n263), .A2(n662), .B1(add_r3[28]), .B2(n125), .ZN(n663)
         );
  INV_X1 U595 ( .A(n663), .ZN(n1107) );
  AOI22_X1 U596 ( .A1(n263), .A2(n664), .B1(add_r3[27]), .B2(n209), .ZN(n665)
         );
  INV_X1 U597 ( .A(n665), .ZN(n1106) );
  AOI22_X1 U598 ( .A1(n263), .A2(n666), .B1(add_r3[26]), .B2(n209), .ZN(n667)
         );
  INV_X1 U599 ( .A(n667), .ZN(n1105) );
  AOI22_X1 U600 ( .A1(n263), .A2(n668), .B1(add_r3[25]), .B2(n125), .ZN(n669)
         );
  INV_X1 U601 ( .A(n669), .ZN(n1104) );
  AOI22_X1 U602 ( .A1(n263), .A2(n670), .B1(add_r3[24]), .B2(n209), .ZN(n671)
         );
  INV_X1 U603 ( .A(n671), .ZN(n1103) );
  AOI22_X1 U604 ( .A1(n264), .A2(n672), .B1(add_r3[23]), .B2(n210), .ZN(n673)
         );
  INV_X1 U605 ( .A(n673), .ZN(n1102) );
  AOI22_X1 U606 ( .A1(n264), .A2(n674), .B1(add_r3[22]), .B2(n8), .ZN(n675) );
  INV_X1 U607 ( .A(n675), .ZN(n1101) );
  AOI22_X1 U608 ( .A1(n264), .A2(n676), .B1(add_r3[21]), .B2(n8), .ZN(n677) );
  INV_X1 U609 ( .A(n677), .ZN(n1100) );
  AOI22_X1 U610 ( .A1(n264), .A2(n678), .B1(add_r3[20]), .B2(n8), .ZN(n679) );
  INV_X1 U611 ( .A(n679), .ZN(n1099) );
  AOI22_X1 U612 ( .A1(n264), .A2(n680), .B1(add_r3[19]), .B2(n222), .ZN(n681)
         );
  INV_X1 U613 ( .A(n681), .ZN(n1098) );
  AOI22_X1 U614 ( .A1(n264), .A2(n682), .B1(add_r3[18]), .B2(n221), .ZN(n683)
         );
  INV_X1 U615 ( .A(n683), .ZN(n1097) );
  AOI22_X1 U616 ( .A1(n264), .A2(n684), .B1(add_r3[17]), .B2(n221), .ZN(n685)
         );
  INV_X1 U617 ( .A(n685), .ZN(n1096) );
  AOI22_X1 U618 ( .A1(n264), .A2(f3[16]), .B1(add_r3[16]), .B2(n222), .ZN(n686) );
  INV_X1 U619 ( .A(n686), .ZN(n1095) );
  AOI22_X1 U620 ( .A1(n264), .A2(f3[15]), .B1(add_r3[15]), .B2(n221), .ZN(n687) );
  INV_X1 U621 ( .A(n687), .ZN(n1094) );
  AOI22_X1 U622 ( .A1(n264), .A2(f3[13]), .B1(add_r3[13]), .B2(n222), .ZN(n688) );
  INV_X1 U623 ( .A(n688), .ZN(n1092) );
  AOI22_X1 U624 ( .A1(n264), .A2(f3[12]), .B1(add_r3[12]), .B2(n221), .ZN(n689) );
  INV_X1 U625 ( .A(n689), .ZN(n1091) );
  AOI22_X1 U626 ( .A1(n264), .A2(f3[11]), .B1(add_r3[11]), .B2(n221), .ZN(n690) );
  INV_X1 U627 ( .A(n690), .ZN(n1090) );
  AOI22_X1 U628 ( .A1(n264), .A2(f3[10]), .B1(add_r3[10]), .B2(n221), .ZN(n691) );
  INV_X1 U629 ( .A(n691), .ZN(n1089) );
  AOI22_X1 U630 ( .A1(n263), .A2(f3[9]), .B1(add_r3[9]), .B2(n222), .ZN(n692)
         );
  INV_X1 U631 ( .A(n692), .ZN(n1088) );
  AOI22_X1 U632 ( .A1(n262), .A2(f3[8]), .B1(add_r3[8]), .B2(n221), .ZN(n693)
         );
  INV_X1 U633 ( .A(n693), .ZN(n1087) );
  AOI22_X1 U634 ( .A1(n261), .A2(f3[7]), .B1(add_r3[7]), .B2(n222), .ZN(n694)
         );
  INV_X1 U635 ( .A(n694), .ZN(n1086) );
  AOI22_X1 U636 ( .A1(n260), .A2(f3[6]), .B1(add_r3[6]), .B2(n221), .ZN(n695)
         );
  INV_X1 U637 ( .A(n695), .ZN(n1085) );
  AOI22_X1 U638 ( .A1(n259), .A2(f3[5]), .B1(add_r3[5]), .B2(n222), .ZN(n696)
         );
  INV_X1 U639 ( .A(n696), .ZN(n1084) );
  AOI22_X1 U640 ( .A1(n264), .A2(f3[4]), .B1(add_r3[4]), .B2(n221), .ZN(n697)
         );
  INV_X1 U641 ( .A(n697), .ZN(n1083) );
  AOI22_X1 U642 ( .A1(n263), .A2(f3[3]), .B1(add_r3[3]), .B2(n222), .ZN(n698)
         );
  INV_X1 U643 ( .A(n698), .ZN(n1082) );
  AOI22_X1 U644 ( .A1(n262), .A2(f3[2]), .B1(add_r3[2]), .B2(n221), .ZN(n699)
         );
  INV_X1 U645 ( .A(n699), .ZN(n1081) );
  AOI22_X1 U646 ( .A1(n261), .A2(f3[1]), .B1(add_r3[1]), .B2(n222), .ZN(n700)
         );
  INV_X1 U647 ( .A(n700), .ZN(n1080) );
  AOI22_X1 U648 ( .A1(n260), .A2(f3[0]), .B1(add_r3[0]), .B2(n221), .ZN(n701)
         );
  INV_X1 U649 ( .A(n701), .ZN(n1079) );
  AOI22_X1 U650 ( .A1(n259), .A2(f3[14]), .B1(add_r3[14]), .B2(n222), .ZN(n702) );
  INV_X1 U651 ( .A(n702), .ZN(n1093) );
  AOI22_X1 U652 ( .A1(n265), .A2(n703), .B1(add_r5[39]), .B2(n226), .ZN(n704)
         );
  INV_X1 U653 ( .A(n704), .ZN(n1038) );
  AOI22_X1 U654 ( .A1(n265), .A2(n705), .B1(add_r5[38]), .B2(n226), .ZN(n706)
         );
  INV_X1 U655 ( .A(n706), .ZN(n1037) );
  AOI22_X1 U656 ( .A1(n265), .A2(n707), .B1(add_r5[37]), .B2(n226), .ZN(n708)
         );
  INV_X1 U657 ( .A(n708), .ZN(n1036) );
  AOI22_X1 U658 ( .A1(n265), .A2(n709), .B1(add_r5[36]), .B2(n226), .ZN(n710)
         );
  INV_X1 U659 ( .A(n710), .ZN(n1035) );
  AOI22_X1 U660 ( .A1(n265), .A2(n711), .B1(add_r5[35]), .B2(n226), .ZN(n712)
         );
  INV_X1 U661 ( .A(n712), .ZN(n1034) );
  AOI22_X1 U662 ( .A1(n265), .A2(n713), .B1(add_r5[34]), .B2(n223), .ZN(n714)
         );
  INV_X1 U663 ( .A(n714), .ZN(n1033) );
  AOI22_X1 U664 ( .A1(n265), .A2(n715), .B1(add_r5[33]), .B2(n226), .ZN(n716)
         );
  INV_X1 U665 ( .A(n716), .ZN(n1032) );
  AOI22_X1 U666 ( .A1(n265), .A2(f5[32]), .B1(add_r5[32]), .B2(n226), .ZN(n717) );
  INV_X1 U667 ( .A(n717), .ZN(n1031) );
  AOI22_X1 U668 ( .A1(n265), .A2(n718), .B1(add_r5[31]), .B2(n226), .ZN(n719)
         );
  INV_X1 U669 ( .A(n719), .ZN(n1030) );
  AOI22_X1 U670 ( .A1(n265), .A2(n720), .B1(add_r5[30]), .B2(n226), .ZN(n721)
         );
  INV_X1 U671 ( .A(n721), .ZN(n1029) );
  AOI22_X1 U672 ( .A1(n265), .A2(n722), .B1(add_r5[29]), .B2(n249), .ZN(n723)
         );
  INV_X1 U673 ( .A(n723), .ZN(n1028) );
  AOI22_X1 U674 ( .A1(n265), .A2(n724), .B1(add_r5[28]), .B2(n249), .ZN(n725)
         );
  INV_X1 U675 ( .A(n725), .ZN(n1027) );
  AOI22_X1 U676 ( .A1(n266), .A2(n726), .B1(add_r5[27]), .B2(n249), .ZN(n727)
         );
  INV_X1 U677 ( .A(n727), .ZN(n1026) );
  AOI22_X1 U678 ( .A1(n266), .A2(n728), .B1(add_r5[26]), .B2(n249), .ZN(n729)
         );
  INV_X1 U679 ( .A(n729), .ZN(n1025) );
  AOI22_X1 U680 ( .A1(n266), .A2(n730), .B1(add_r5[25]), .B2(n249), .ZN(n731)
         );
  INV_X1 U681 ( .A(n731), .ZN(n1024) );
  AOI22_X1 U682 ( .A1(n266), .A2(n732), .B1(add_r5[24]), .B2(n249), .ZN(n733)
         );
  INV_X1 U683 ( .A(n733), .ZN(n1023) );
  AOI22_X1 U684 ( .A1(n266), .A2(n734), .B1(add_r5[23]), .B2(n249), .ZN(n735)
         );
  INV_X1 U685 ( .A(n735), .ZN(n1022) );
  AOI22_X1 U686 ( .A1(n266), .A2(n736), .B1(add_r5[22]), .B2(n249), .ZN(n737)
         );
  INV_X1 U687 ( .A(n737), .ZN(n1021) );
  AOI22_X1 U688 ( .A1(n266), .A2(n738), .B1(add_r5[21]), .B2(n249), .ZN(n739)
         );
  INV_X1 U689 ( .A(n739), .ZN(n1020) );
  AOI22_X1 U690 ( .A1(n266), .A2(n740), .B1(add_r5[20]), .B2(n249), .ZN(n741)
         );
  INV_X1 U691 ( .A(n741), .ZN(n1019) );
  AOI22_X1 U692 ( .A1(n266), .A2(n742), .B1(add_r5[19]), .B2(n249), .ZN(n743)
         );
  INV_X1 U693 ( .A(n743), .ZN(n1018) );
  AOI22_X1 U694 ( .A1(n266), .A2(n744), .B1(add_r5[18]), .B2(n249), .ZN(n745)
         );
  INV_X1 U695 ( .A(n745), .ZN(n1017) );
  AOI22_X1 U696 ( .A1(n266), .A2(n746), .B1(add_r5[17]), .B2(n250), .ZN(n747)
         );
  INV_X1 U697 ( .A(n747), .ZN(n1016) );
  AOI22_X1 U698 ( .A1(n266), .A2(f5[16]), .B1(add_r5[16]), .B2(n250), .ZN(n748) );
  INV_X1 U699 ( .A(n748), .ZN(n1015) );
  AOI22_X1 U700 ( .A1(n274), .A2(n749), .B1(add_r5[15]), .B2(n250), .ZN(n750)
         );
  INV_X1 U701 ( .A(n750), .ZN(n1014) );
  AOI22_X1 U702 ( .A1(n274), .A2(f5[13]), .B1(add_r5[13]), .B2(n250), .ZN(n751) );
  INV_X1 U703 ( .A(n751), .ZN(n1012) );
  AOI22_X1 U704 ( .A1(n274), .A2(f5[12]), .B1(add_r5[12]), .B2(n250), .ZN(n752) );
  INV_X1 U705 ( .A(n752), .ZN(n1011) );
  AOI22_X1 U706 ( .A1(n274), .A2(f5[11]), .B1(add_r5[11]), .B2(n250), .ZN(n753) );
  INV_X1 U707 ( .A(n753), .ZN(n1010) );
  AOI22_X1 U708 ( .A1(n274), .A2(f5[10]), .B1(add_r5[10]), .B2(n250), .ZN(n754) );
  INV_X1 U709 ( .A(n754), .ZN(n1009) );
  AOI22_X1 U710 ( .A1(n274), .A2(f5[9]), .B1(add_r5[9]), .B2(n250), .ZN(n755)
         );
  INV_X1 U711 ( .A(n755), .ZN(n1008) );
  AOI22_X1 U712 ( .A1(n274), .A2(f5[8]), .B1(add_r5[8]), .B2(n250), .ZN(n756)
         );
  INV_X1 U713 ( .A(n756), .ZN(n1007) );
  AOI22_X1 U714 ( .A1(n274), .A2(f5[7]), .B1(add_r5[7]), .B2(n250), .ZN(n757)
         );
  INV_X1 U715 ( .A(n757), .ZN(n1006) );
  AOI22_X1 U716 ( .A1(n274), .A2(f5[6]), .B1(add_r5[6]), .B2(n250), .ZN(n758)
         );
  INV_X1 U717 ( .A(n758), .ZN(n1005) );
  AOI22_X1 U718 ( .A1(n274), .A2(f5[5]), .B1(add_r5[5]), .B2(n250), .ZN(n759)
         );
  INV_X1 U719 ( .A(n759), .ZN(n1004) );
  AOI22_X1 U720 ( .A1(n274), .A2(f5[4]), .B1(add_r5[4]), .B2(n251), .ZN(n760)
         );
  INV_X1 U721 ( .A(n760), .ZN(n1003) );
  AOI22_X1 U722 ( .A1(n274), .A2(f5[3]), .B1(add_r5[3]), .B2(n251), .ZN(n761)
         );
  INV_X1 U723 ( .A(n761), .ZN(n1002) );
  AOI22_X1 U724 ( .A1(n275), .A2(f5[2]), .B1(add_r5[2]), .B2(n251), .ZN(n762)
         );
  INV_X1 U725 ( .A(n762), .ZN(n1001) );
  AOI22_X1 U726 ( .A1(n275), .A2(f5[1]), .B1(add_r5[1]), .B2(n251), .ZN(n763)
         );
  INV_X1 U727 ( .A(n763), .ZN(n1000) );
  AOI22_X1 U728 ( .A1(n275), .A2(f5[0]), .B1(add_r5[0]), .B2(n221), .ZN(n764)
         );
  INV_X1 U729 ( .A(n764), .ZN(n999) );
  AOI22_X1 U730 ( .A1(n275), .A2(f5[14]), .B1(add_r5[14]), .B2(n226), .ZN(n765) );
  INV_X1 U731 ( .A(n765), .ZN(n1013) );
  AOI22_X1 U732 ( .A1(n275), .A2(n766), .B1(add_r2[39]), .B2(n226), .ZN(n767)
         );
  INV_X1 U733 ( .A(n767), .ZN(n1158) );
  AOI22_X1 U734 ( .A1(n275), .A2(n768), .B1(add_r2[38]), .B2(n226), .ZN(n769)
         );
  INV_X1 U735 ( .A(n769), .ZN(n1157) );
  AOI22_X1 U736 ( .A1(n275), .A2(n770), .B1(add_r2[37]), .B2(n225), .ZN(n771)
         );
  INV_X1 U737 ( .A(n771), .ZN(n1156) );
  AOI22_X1 U738 ( .A1(n275), .A2(n772), .B1(add_r2[36]), .B2(n225), .ZN(n773)
         );
  INV_X1 U739 ( .A(n773), .ZN(n1155) );
  AOI22_X1 U740 ( .A1(n275), .A2(n774), .B1(add_r2[35]), .B2(n225), .ZN(n775)
         );
  INV_X1 U741 ( .A(n775), .ZN(n1154) );
  AOI22_X1 U742 ( .A1(n275), .A2(n776), .B1(add_r2[34]), .B2(n225), .ZN(n777)
         );
  INV_X1 U743 ( .A(n777), .ZN(n1153) );
  AOI22_X1 U744 ( .A1(n275), .A2(n778), .B1(add_r2[33]), .B2(n225), .ZN(n779)
         );
  INV_X1 U745 ( .A(n779), .ZN(n1152) );
  AOI22_X1 U746 ( .A1(n275), .A2(n780), .B1(add_r2[32]), .B2(n225), .ZN(n781)
         );
  INV_X1 U747 ( .A(n781), .ZN(n1151) );
  AOI22_X1 U748 ( .A1(n266), .A2(n782), .B1(add_r2[31]), .B2(n225), .ZN(n783)
         );
  INV_X1 U749 ( .A(n783), .ZN(n1150) );
  AOI22_X1 U750 ( .A1(n265), .A2(n784), .B1(add_r2[30]), .B2(n225), .ZN(n785)
         );
  INV_X1 U751 ( .A(n785), .ZN(n1149) );
  AOI22_X1 U752 ( .A1(n257), .A2(n786), .B1(add_r2[29]), .B2(n225), .ZN(n787)
         );
  INV_X1 U753 ( .A(n787), .ZN(n1148) );
  AOI22_X1 U754 ( .A1(n258), .A2(n788), .B1(add_r2[28]), .B2(n225), .ZN(n789)
         );
  INV_X1 U755 ( .A(n789), .ZN(n1147) );
  AOI22_X1 U756 ( .A1(n264), .A2(n790), .B1(add_r2[27]), .B2(n225), .ZN(n791)
         );
  INV_X1 U757 ( .A(n791), .ZN(n1146) );
  AOI22_X1 U758 ( .A1(n263), .A2(n792), .B1(add_r2[26]), .B2(n225), .ZN(n793)
         );
  INV_X1 U759 ( .A(n793), .ZN(n1145) );
  AOI22_X1 U760 ( .A1(n262), .A2(n794), .B1(add_r2[25]), .B2(n224), .ZN(n795)
         );
  INV_X1 U761 ( .A(n795), .ZN(n1144) );
  AOI22_X1 U762 ( .A1(n261), .A2(n796), .B1(add_r2[24]), .B2(n224), .ZN(n797)
         );
  INV_X1 U763 ( .A(n797), .ZN(n1143) );
  AOI22_X1 U764 ( .A1(n260), .A2(n798), .B1(add_r2[23]), .B2(n224), .ZN(n799)
         );
  INV_X1 U765 ( .A(n799), .ZN(n1142) );
  AOI22_X1 U766 ( .A1(n259), .A2(n800), .B1(add_r2[22]), .B2(n224), .ZN(n801)
         );
  INV_X1 U767 ( .A(n801), .ZN(n1141) );
  AOI22_X1 U768 ( .A1(n275), .A2(n802), .B1(add_r2[21]), .B2(n224), .ZN(n803)
         );
  INV_X1 U769 ( .A(n803), .ZN(n1140) );
  AOI22_X1 U770 ( .A1(n274), .A2(n804), .B1(add_r2[20]), .B2(n224), .ZN(n805)
         );
  INV_X1 U771 ( .A(n805), .ZN(n1139) );
  AOI22_X1 U772 ( .A1(n274), .A2(n806), .B1(add_r2[19]), .B2(n224), .ZN(n807)
         );
  INV_X1 U773 ( .A(n807), .ZN(n1138) );
  AOI22_X1 U774 ( .A1(n266), .A2(n808), .B1(add_r2[18]), .B2(n224), .ZN(n809)
         );
  INV_X1 U775 ( .A(n809), .ZN(n1137) );
  AOI22_X1 U776 ( .A1(n265), .A2(n810), .B1(add_r2[17]), .B2(n224), .ZN(n811)
         );
  INV_X1 U777 ( .A(n811), .ZN(n1136) );
  AOI22_X1 U778 ( .A1(n264), .A2(f2[16]), .B1(add_r2[16]), .B2(n224), .ZN(n812) );
  INV_X1 U779 ( .A(n812), .ZN(n1135) );
  AOI22_X1 U780 ( .A1(n263), .A2(f2[15]), .B1(add_r2[15]), .B2(n224), .ZN(n813) );
  INV_X1 U781 ( .A(n813), .ZN(n1134) );
  AOI22_X1 U782 ( .A1(n262), .A2(f2[13]), .B1(add_r2[13]), .B2(n224), .ZN(n814) );
  INV_X1 U783 ( .A(n814), .ZN(n1132) );
  AOI22_X1 U784 ( .A1(n261), .A2(f2[12]), .B1(add_r2[12]), .B2(n223), .ZN(n815) );
  INV_X1 U785 ( .A(n815), .ZN(n1131) );
  AOI22_X1 U786 ( .A1(n260), .A2(f2[11]), .B1(add_r2[11]), .B2(n223), .ZN(n816) );
  INV_X1 U787 ( .A(n816), .ZN(n1130) );
  AOI22_X1 U788 ( .A1(n259), .A2(f2[10]), .B1(add_r2[10]), .B2(n223), .ZN(n817) );
  INV_X1 U789 ( .A(n817), .ZN(n1129) );
  AOI22_X1 U790 ( .A1(n275), .A2(f2[9]), .B1(add_r2[9]), .B2(n223), .ZN(n818)
         );
  INV_X1 U791 ( .A(n818), .ZN(n1128) );
  AOI22_X1 U792 ( .A1(n275), .A2(f2[8]), .B1(add_r2[8]), .B2(n223), .ZN(n819)
         );
  INV_X1 U793 ( .A(n819), .ZN(n1127) );
  AOI22_X1 U794 ( .A1(n274), .A2(f2[7]), .B1(add_r2[7]), .B2(n223), .ZN(n820)
         );
  INV_X1 U795 ( .A(n820), .ZN(n1126) );
  AOI22_X1 U796 ( .A1(n263), .A2(f2[6]), .B1(add_r2[6]), .B2(n223), .ZN(n821)
         );
  INV_X1 U797 ( .A(n821), .ZN(n1125) );
  AOI22_X1 U798 ( .A1(n262), .A2(f2[5]), .B1(add_r2[5]), .B2(n223), .ZN(n822)
         );
  INV_X1 U799 ( .A(n822), .ZN(n1124) );
  AOI22_X1 U800 ( .A1(n266), .A2(f2[4]), .B1(add_r2[4]), .B2(n223), .ZN(n823)
         );
  INV_X1 U801 ( .A(n823), .ZN(n1123) );
  AOI22_X1 U802 ( .A1(n275), .A2(f2[3]), .B1(add_r2[3]), .B2(n223), .ZN(n824)
         );
  INV_X1 U803 ( .A(n824), .ZN(n1122) );
  AOI22_X1 U804 ( .A1(n274), .A2(f2[2]), .B1(add_r2[2]), .B2(n223), .ZN(n825)
         );
  INV_X1 U805 ( .A(n825), .ZN(n1121) );
  AOI22_X1 U806 ( .A1(n266), .A2(f2[1]), .B1(add_r2[1]), .B2(n222), .ZN(n826)
         );
  INV_X1 U807 ( .A(n826), .ZN(n1120) );
  AOI22_X1 U808 ( .A1(n265), .A2(f2[0]), .B1(add_r2[0]), .B2(n222), .ZN(n827)
         );
  INV_X1 U809 ( .A(n827), .ZN(n1119) );
  AOI22_X1 U810 ( .A1(n266), .A2(f2[14]), .B1(add_r2[14]), .B2(n251), .ZN(n829) );
  INV_X1 U811 ( .A(n829), .ZN(n1133) );
  INV_X1 U812 ( .A(n350), .ZN(n1352) );
  NAND2_X1 U813 ( .A1(n336), .A2(n516), .ZN(n1350) );
  OAI222_X1 U814 ( .A1(n337), .A2(n34), .B1(n336), .B2(n830), .C1(n124), .C2(
        n234), .ZN(n831) );
  AOI221_X1 U815 ( .B1(f7[14]), .B2(n346), .C1(f8[14]), .C2(n340), .A(n831), 
        .ZN(n834) );
  OAI22_X1 U816 ( .A1(n345), .A2(n74), .B1(n348), .B2(n194), .ZN(n832) );
  AOI221_X1 U817 ( .B1(f4[14]), .B2(n341), .C1(f3[14]), .C2(n354), .A(n832), 
        .ZN(n833) );
  NAND2_X1 U818 ( .A1(n834), .A2(n833), .ZN(n864) );
  OAI222_X1 U819 ( .A1(n1350), .A2(n35), .B1(n336), .B2(n835), .C1(n124), .C2(
        n235), .ZN(n836) );
  AOI221_X1 U820 ( .B1(f7[13]), .B2(n1352), .C1(f8[13]), .C2(n340), .A(n836), 
        .ZN(n1199) );
  OAI22_X1 U821 ( .A1(n347), .A2(n75), .B1(n344), .B2(n195), .ZN(n837) );
  AOI221_X1 U822 ( .B1(f4[13]), .B2(n341), .C1(f3[13]), .C2(n354), .A(n837), 
        .ZN(n838) );
  NAND2_X1 U823 ( .A1(n1199), .A2(n838), .ZN(n865) );
  OAI222_X1 U824 ( .A1(n1350), .A2(n36), .B1(n336), .B2(n1200), .C1(n349), 
        .C2(n236), .ZN(n1201) );
  AOI221_X1 U825 ( .B1(f7[12]), .B2(n1352), .C1(f8[12]), .C2(n340), .A(n1201), 
        .ZN(n1204) );
  OAI22_X1 U826 ( .A1(n347), .A2(n76), .B1(n344), .B2(n196), .ZN(n1202) );
  AOI221_X1 U827 ( .B1(f4[12]), .B2(n341), .C1(f3[12]), .C2(n354), .A(n1202), 
        .ZN(n1203) );
  NAND2_X1 U828 ( .A1(n1204), .A2(n1203), .ZN(n866) );
  OAI222_X1 U829 ( .A1(n1350), .A2(n37), .B1(n336), .B2(n1205), .C1(n124), 
        .C2(n237), .ZN(n1206) );
  AOI221_X1 U830 ( .B1(f7[11]), .B2(n1352), .C1(f8[11]), .C2(n340), .A(n1206), 
        .ZN(n1209) );
  OAI22_X1 U831 ( .A1(n347), .A2(n77), .B1(n344), .B2(n197), .ZN(n1207) );
  AOI221_X1 U832 ( .B1(f4[11]), .B2(n341), .C1(f3[11]), .C2(n354), .A(n1207), 
        .ZN(n1208) );
  NAND2_X1 U833 ( .A1(n1209), .A2(n1208), .ZN(n867) );
  OAI222_X1 U834 ( .A1(n1350), .A2(n38), .B1(n336), .B2(n1210), .C1(n349), 
        .C2(n238), .ZN(n1211) );
  AOI221_X1 U835 ( .B1(f7[10]), .B2(n1352), .C1(f8[10]), .C2(n340), .A(n1211), 
        .ZN(n1214) );
  OAI22_X1 U836 ( .A1(n347), .A2(n78), .B1(n344), .B2(n198), .ZN(n1212) );
  AOI221_X1 U837 ( .B1(f4[10]), .B2(n357), .C1(f3[10]), .C2(n354), .A(n1212), 
        .ZN(n1213) );
  NAND2_X1 U838 ( .A1(n1214), .A2(n1213), .ZN(n868) );
  OAI222_X1 U839 ( .A1(n1350), .A2(n39), .B1(n336), .B2(n1215), .C1(n124), 
        .C2(n239), .ZN(n1216) );
  AOI221_X1 U840 ( .B1(f7[9]), .B2(n1352), .C1(f8[9]), .C2(n340), .A(n1216), 
        .ZN(n1219) );
  OAI22_X1 U841 ( .A1(n347), .A2(n79), .B1(n344), .B2(n199), .ZN(n1217) );
  AOI221_X1 U842 ( .B1(f4[9]), .B2(n357), .C1(f3[9]), .C2(n354), .A(n1217), 
        .ZN(n1218) );
  NAND2_X1 U843 ( .A1(n1219), .A2(n1218), .ZN(n869) );
  OAI222_X1 U844 ( .A1(n1350), .A2(n40), .B1(n336), .B2(n1220), .C1(n349), 
        .C2(n240), .ZN(n1221) );
  AOI221_X1 U845 ( .B1(f7[8]), .B2(n1352), .C1(f8[8]), .C2(n340), .A(n1221), 
        .ZN(n1224) );
  OAI22_X1 U846 ( .A1(n347), .A2(n80), .B1(n344), .B2(n200), .ZN(n1222) );
  AOI221_X1 U847 ( .B1(f4[8]), .B2(n357), .C1(f3[8]), .C2(n354), .A(n1222), 
        .ZN(n1223) );
  NAND2_X1 U848 ( .A1(n1224), .A2(n1223), .ZN(n870) );
  OAI222_X1 U849 ( .A1(n1350), .A2(n41), .B1(n336), .B2(n1225), .C1(n124), 
        .C2(n241), .ZN(n1226) );
  AOI221_X1 U850 ( .B1(f7[7]), .B2(n1352), .C1(f8[7]), .C2(n340), .A(n1226), 
        .ZN(n1229) );
  OAI22_X1 U851 ( .A1(n347), .A2(n81), .B1(n344), .B2(n201), .ZN(n1227) );
  AOI221_X1 U852 ( .B1(f4[7]), .B2(n357), .C1(f3[7]), .C2(n354), .A(n1227), 
        .ZN(n1228) );
  NAND2_X1 U853 ( .A1(n1229), .A2(n1228), .ZN(n871) );
  OAI222_X1 U854 ( .A1(n1350), .A2(n42), .B1(n336), .B2(n1230), .C1(n349), 
        .C2(n242), .ZN(n1231) );
  AOI221_X1 U855 ( .B1(f7[6]), .B2(n1352), .C1(f8[6]), .C2(n358), .A(n1231), 
        .ZN(n1234) );
  OAI22_X1 U856 ( .A1(n347), .A2(n82), .B1(n344), .B2(n202), .ZN(n1232) );
  AOI221_X1 U857 ( .B1(f4[6]), .B2(n357), .C1(f3[6]), .C2(n354), .A(n1232), 
        .ZN(n1233) );
  NAND2_X1 U858 ( .A1(n1234), .A2(n1233), .ZN(n872) );
  OAI222_X1 U859 ( .A1(n337), .A2(n43), .B1(n336), .B2(n1235), .C1(n124), .C2(
        n243), .ZN(n1236) );
  AOI221_X1 U860 ( .B1(f7[5]), .B2(n1352), .C1(f8[5]), .C2(n358), .A(n1236), 
        .ZN(n1239) );
  OAI22_X1 U861 ( .A1(n345), .A2(n83), .B1(n348), .B2(n203), .ZN(n1237) );
  AOI221_X1 U862 ( .B1(f4[5]), .B2(n357), .C1(f3[5]), .C2(n354), .A(n1237), 
        .ZN(n1238) );
  NAND2_X1 U863 ( .A1(n1239), .A2(n1238), .ZN(n873) );
  OAI222_X1 U864 ( .A1(n337), .A2(n44), .B1(n336), .B2(n1240), .C1(n349), .C2(
        n244), .ZN(n1241) );
  AOI221_X1 U865 ( .B1(f7[4]), .B2(n1352), .C1(f8[4]), .C2(n358), .A(n1241), 
        .ZN(n1244) );
  OAI22_X1 U866 ( .A1(n345), .A2(n84), .B1(n348), .B2(n204), .ZN(n1242) );
  AOI221_X1 U867 ( .B1(f4[4]), .B2(n357), .C1(f3[4]), .C2(n354), .A(n1242), 
        .ZN(n1243) );
  NAND2_X1 U868 ( .A1(n1244), .A2(n1243), .ZN(n874) );
  OAI222_X1 U869 ( .A1(n337), .A2(n45), .B1(n336), .B2(n1245), .C1(n124), .C2(
        n245), .ZN(n1246) );
  AOI221_X1 U870 ( .B1(f7[3]), .B2(n1352), .C1(f8[3]), .C2(n358), .A(n1246), 
        .ZN(n1249) );
  OAI22_X1 U871 ( .A1(n345), .A2(n85), .B1(n348), .B2(n205), .ZN(n1247) );
  AOI221_X1 U872 ( .B1(f4[3]), .B2(n357), .C1(f3[3]), .C2(n354), .A(n1247), 
        .ZN(n1248) );
  NAND2_X1 U873 ( .A1(n1249), .A2(n1248), .ZN(n875) );
  OAI222_X1 U874 ( .A1(n337), .A2(n46), .B1(n336), .B2(n1250), .C1(n349), .C2(
        n246), .ZN(n1251) );
  AOI221_X1 U875 ( .B1(f7[2]), .B2(n1352), .C1(f8[2]), .C2(n358), .A(n1251), 
        .ZN(n1254) );
  OAI22_X1 U876 ( .A1(n345), .A2(n86), .B1(n348), .B2(n206), .ZN(n1252) );
  AOI221_X1 U877 ( .B1(f4[2]), .B2(n357), .C1(f3[2]), .C2(n354), .A(n1252), 
        .ZN(n1253) );
  NAND2_X1 U878 ( .A1(n1254), .A2(n1253), .ZN(n876) );
  OAI222_X1 U879 ( .A1(n1350), .A2(n47), .B1(n336), .B2(n1255), .C1(n124), 
        .C2(n247), .ZN(n1256) );
  AOI221_X1 U880 ( .B1(f7[1]), .B2(n1352), .C1(f8[1]), .C2(n358), .A(n1256), 
        .ZN(n1259) );
  OAI22_X1 U881 ( .A1(n345), .A2(n87), .B1(n348), .B2(n207), .ZN(n1257) );
  AOI221_X1 U882 ( .B1(f4[1]), .B2(n357), .C1(f3[1]), .C2(n354), .A(n1257), 
        .ZN(n1258) );
  NAND2_X1 U883 ( .A1(n1259), .A2(n1258), .ZN(n877) );
  OAI222_X1 U884 ( .A1(n1350), .A2(n48), .B1(n336), .B2(n1260), .C1(n349), 
        .C2(n248), .ZN(n1261) );
  AOI221_X1 U885 ( .B1(f7[0]), .B2(n1352), .C1(f8[0]), .C2(n358), .A(n1261), 
        .ZN(n1264) );
  OAI22_X1 U886 ( .A1(n345), .A2(n88), .B1(n348), .B2(n208), .ZN(n1262) );
  AOI221_X1 U887 ( .B1(f4[0]), .B2(n357), .C1(f3[0]), .C2(n354), .A(n1262), 
        .ZN(n1263) );
  NAND2_X1 U888 ( .A1(n1264), .A2(n1263), .ZN(n878) );
  INV_X1 U889 ( .A(n349), .ZN(n1354) );
  OAI22_X1 U890 ( .A1(n1350), .A2(n9), .B1(n336), .B2(n1265), .ZN(n1266) );
  AOI221_X1 U891 ( .B1(n1268), .B2(n1354), .C1(n1267), .C2(n1352), .A(n1266), 
        .ZN(n415) );
  OAI222_X1 U892 ( .A1(n348), .A2(n186), .B1(n343), .B2(n106), .C1(n345), .C2(
        n66), .ZN(n1269) );
  AOI221_X1 U893 ( .B1(f4[22]), .B2(n357), .C1(f8[22]), .C2(n358), .A(n1269), 
        .ZN(n416) );
  OAI22_X1 U894 ( .A1(n1350), .A2(n10), .B1(n336), .B2(n1270), .ZN(n1271) );
  AOI221_X1 U895 ( .B1(n1273), .B2(n1354), .C1(n1272), .C2(n1352), .A(n1271), 
        .ZN(n411) );
  OAI222_X1 U896 ( .A1(n348), .A2(n185), .B1(n343), .B2(n105), .C1(n345), .C2(
        n65), .ZN(n1274) );
  AOI221_X1 U897 ( .B1(f4[23]), .B2(n357), .C1(f8[23]), .C2(n358), .A(n1274), 
        .ZN(n412) );
  OAI22_X1 U898 ( .A1(n1350), .A2(n11), .B1(n336), .B2(n1275), .ZN(n1276) );
  AOI221_X1 U899 ( .B1(n1278), .B2(n1354), .C1(n1277), .C2(n1352), .A(n1276), 
        .ZN(n407) );
  OAI222_X1 U900 ( .A1(n348), .A2(n184), .B1(n343), .B2(n104), .C1(n345), .C2(
        n64), .ZN(n1279) );
  AOI221_X1 U901 ( .B1(f4[24]), .B2(n357), .C1(f8[24]), .C2(n358), .A(n1279), 
        .ZN(n408) );
  OAI22_X1 U902 ( .A1(n1350), .A2(n12), .B1(n336), .B2(n1280), .ZN(n1281) );
  AOI221_X1 U903 ( .B1(n1283), .B2(n1354), .C1(n1282), .C2(n1352), .A(n1281), 
        .ZN(n403) );
  OAI222_X1 U904 ( .A1(n348), .A2(n183), .B1(n343), .B2(n103), .C1(n345), .C2(
        n63), .ZN(n1284) );
  AOI221_X1 U905 ( .B1(f4[25]), .B2(n357), .C1(f8[25]), .C2(n358), .A(n1284), 
        .ZN(n404) );
  OAI22_X1 U906 ( .A1(n1350), .A2(n13), .B1(n336), .B2(n1285), .ZN(n1286) );
  AOI221_X1 U907 ( .B1(n1288), .B2(n1354), .C1(n1287), .C2(n1352), .A(n1286), 
        .ZN(n399) );
  OAI222_X1 U908 ( .A1(n348), .A2(n182), .B1(n343), .B2(n102), .C1(n345), .C2(
        n62), .ZN(n1289) );
  AOI221_X1 U909 ( .B1(f4[26]), .B2(n357), .C1(f8[26]), .C2(n358), .A(n1289), 
        .ZN(n400) );
  OAI22_X1 U910 ( .A1(n1350), .A2(n14), .B1(n336), .B2(n1290), .ZN(n1291) );
  AOI221_X1 U911 ( .B1(n1293), .B2(n1354), .C1(n1292), .C2(n1352), .A(n1291), 
        .ZN(n395) );
  OAI222_X1 U912 ( .A1(n348), .A2(n181), .B1(n343), .B2(n101), .C1(n345), .C2(
        n61), .ZN(n1294) );
  AOI221_X1 U913 ( .B1(f4[27]), .B2(n357), .C1(f8[27]), .C2(n358), .A(n1294), 
        .ZN(n396) );
  OAI22_X1 U914 ( .A1(n337), .A2(n15), .B1(n335), .B2(n1295), .ZN(n1296) );
  AOI221_X1 U915 ( .B1(n1298), .B2(n1354), .C1(n1297), .C2(n346), .A(n1296), 
        .ZN(n391) );
  OAI222_X1 U916 ( .A1(n348), .A2(n180), .B1(n343), .B2(n100), .C1(n345), .C2(
        n60), .ZN(n1299) );
  AOI221_X1 U917 ( .B1(f4[28]), .B2(n357), .C1(f8[28]), .C2(n358), .A(n1299), 
        .ZN(n392) );
  OAI22_X1 U918 ( .A1(n337), .A2(n16), .B1(n335), .B2(n1300), .ZN(n1301) );
  AOI221_X1 U919 ( .B1(n1303), .B2(n1354), .C1(n1302), .C2(n346), .A(n1301), 
        .ZN(n387) );
  OAI222_X1 U920 ( .A1(n348), .A2(n179), .B1(n343), .B2(n99), .C1(n345), .C2(
        n59), .ZN(n1304) );
  AOI221_X1 U921 ( .B1(f4[29]), .B2(n357), .C1(f8[29]), .C2(n358), .A(n1304), 
        .ZN(n388) );
  OAI22_X1 U922 ( .A1(n337), .A2(n17), .B1(n335), .B2(n1305), .ZN(n1306) );
  AOI221_X1 U923 ( .B1(n1308), .B2(n1354), .C1(n1307), .C2(n346), .A(n1306), 
        .ZN(n383) );
  OAI222_X1 U924 ( .A1(n348), .A2(n178), .B1(n343), .B2(n98), .C1(n345), .C2(
        n58), .ZN(n1309) );
  AOI221_X1 U925 ( .B1(f4[30]), .B2(n357), .C1(f8[30]), .C2(n358), .A(n1309), 
        .ZN(n384) );
  OAI22_X1 U926 ( .A1(n337), .A2(n18), .B1(n335), .B2(n1310), .ZN(n1311) );
  AOI221_X1 U927 ( .B1(n1313), .B2(n1354), .C1(n1312), .C2(n346), .A(n1311), 
        .ZN(n379) );
  OAI222_X1 U928 ( .A1(n348), .A2(n177), .B1(n343), .B2(n97), .C1(n345), .C2(
        n57), .ZN(n1314) );
  AOI221_X1 U929 ( .B1(f4[31]), .B2(n357), .C1(f8[31]), .C2(n358), .A(n1314), 
        .ZN(n380) );
  OAI22_X1 U930 ( .A1(n337), .A2(n19), .B1(n335), .B2(n1315), .ZN(n1316) );
  AOI221_X1 U931 ( .B1(n1317), .B2(n1354), .C1(f7[32]), .C2(n346), .A(n1316), 
        .ZN(n375) );
  OAI222_X1 U932 ( .A1(n348), .A2(n176), .B1(n353), .B2(n96), .C1(n345), .C2(
        n56), .ZN(n1318) );
  AOI221_X1 U933 ( .B1(f4[32]), .B2(n341), .C1(f8[32]), .C2(n358), .A(n1318), 
        .ZN(n376) );
  OAI22_X1 U934 ( .A1(n337), .A2(n20), .B1(n335), .B2(n1319), .ZN(n1320) );
  AOI221_X1 U935 ( .B1(n1322), .B2(n1354), .C1(n1321), .C2(n346), .A(n1320), 
        .ZN(n371) );
  OAI222_X1 U936 ( .A1(n348), .A2(n175), .B1(n353), .B2(n95), .C1(n345), .C2(
        n55), .ZN(n1323) );
  AOI221_X1 U937 ( .B1(f4[33]), .B2(n357), .C1(f8[33]), .C2(n340), .A(n1323), 
        .ZN(n372) );
  OAI22_X1 U938 ( .A1(n337), .A2(n21), .B1(n335), .B2(n1324), .ZN(n1325) );
  AOI221_X1 U939 ( .B1(n1327), .B2(n1354), .C1(n1326), .C2(n346), .A(n1325), 
        .ZN(n367) );
  OAI222_X1 U940 ( .A1(n348), .A2(n174), .B1(n353), .B2(n94), .C1(n345), .C2(
        n54), .ZN(n1328) );
  AOI221_X1 U941 ( .B1(f4[34]), .B2(n341), .C1(f8[34]), .C2(n340), .A(n1328), 
        .ZN(n368) );
  OAI22_X1 U942 ( .A1(n337), .A2(n22), .B1(n335), .B2(n1329), .ZN(n1330) );
  AOI221_X1 U943 ( .B1(n1332), .B2(n1354), .C1(n1331), .C2(n346), .A(n1330), 
        .ZN(n363) );
  OAI222_X1 U944 ( .A1(n344), .A2(n173), .B1(n353), .B2(n93), .C1(n347), .C2(
        n53), .ZN(n1333) );
  AOI221_X1 U945 ( .B1(f4[35]), .B2(n341), .C1(f8[35]), .C2(n340), .A(n1333), 
        .ZN(n364) );
  OAI22_X1 U946 ( .A1(n337), .A2(n23), .B1(n335), .B2(n1334), .ZN(n1335) );
  AOI221_X1 U947 ( .B1(n1337), .B2(n1354), .C1(n1336), .C2(n346), .A(n1335), 
        .ZN(n359) );
  OAI222_X1 U948 ( .A1(n344), .A2(n172), .B1(n353), .B2(n92), .C1(n347), .C2(
        n52), .ZN(n1338) );
  AOI221_X1 U949 ( .B1(f4[36]), .B2(n341), .C1(f8[36]), .C2(n340), .A(n1338), 
        .ZN(n360) );
  OAI22_X1 U950 ( .A1(n337), .A2(n24), .B1(n335), .B2(n1339), .ZN(n1340) );
  AOI221_X1 U951 ( .B1(n1342), .B2(n1354), .C1(n1341), .C2(n346), .A(n1340), 
        .ZN(n355) );
  OAI222_X1 U952 ( .A1(n344), .A2(n171), .B1(n353), .B2(n91), .C1(n347), .C2(
        n51), .ZN(n1343) );
  AOI221_X1 U953 ( .B1(f4[37]), .B2(n341), .C1(f8[37]), .C2(n340), .A(n1343), 
        .ZN(n356) );
  OAI22_X1 U954 ( .A1(n337), .A2(n25), .B1(n335), .B2(n1344), .ZN(n1345) );
  AOI221_X1 U955 ( .B1(n1347), .B2(n1354), .C1(n1346), .C2(n346), .A(n1345), 
        .ZN(n351) );
  OAI222_X1 U956 ( .A1(n344), .A2(n170), .B1(n353), .B2(n90), .C1(n347), .C2(
        n50), .ZN(n1348) );
  AOI221_X1 U957 ( .B1(f4[38]), .B2(n341), .C1(f8[38]), .C2(n340), .A(n1348), 
        .ZN(n352) );
  OAI22_X1 U958 ( .A1(n337), .A2(n26), .B1(n336), .B2(n1349), .ZN(n1351) );
  AOI221_X1 U959 ( .B1(n1355), .B2(n1354), .C1(n1353), .C2(n346), .A(n1351), 
        .ZN(n338) );
  OAI222_X1 U960 ( .A1(n344), .A2(n169), .B1(n353), .B2(n89), .C1(n347), .C2(
        n49), .ZN(n1356) );
  AOI221_X1 U961 ( .B1(f4[39]), .B2(n341), .C1(f8[39]), .C2(n340), .A(n1356), 
        .ZN(n339) );
endmodule


module ctrlpath ( clk, reset, start, addr_x, wr_en_x, addr_a1, addr_a2, 
        addr_a3, addr_a4, addr_a5, addr_a6, addr_a7, addr_a8, wr_en_a1, 
        wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6, wr_en_a7, wr_en_a8, 
        clear_acc, clc, clc1, addr_y, wr_en_y, done, loadMatrix, loadVector );
  output [2:0] addr_x;
  output [2:0] addr_a1;
  output [2:0] addr_a2;
  output [2:0] addr_a3;
  output [2:0] addr_a4;
  output [2:0] addr_a5;
  output [2:0] addr_a6;
  output [2:0] addr_a7;
  output [2:0] addr_a8;
  output [2:0] addr_y;
  input clk, reset, start, loadMatrix, loadVector;
  output wr_en_x, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6,
         wr_en_a7, wr_en_a8, clear_acc, clc, clc1, wr_en_y, done;
  wire   N32, N33, N34, N35, N37, N45, N46, N56, N57, N67, N68, N78, N79, N89,
         N90, N100, N101, N111, N112, N122, N123, N131, N132, N133, N141, N142,
         N143, N146, N147, N148, n76, n79, n80, n81, n83, n84, n85, n86, n87,
         n88, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n111, n112, n113, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39;
  wire   [4:0] state;

  DFF_X1 \state_reg[3]  ( .D(N35), .CK(clk), .Q(state[3]) );
  DFF_X1 done_reg ( .D(N37), .CK(clk), .Q(done) );
  DFF_X1 \addr_x_reg[0]  ( .D(N131), .CK(clk), .Q(addr_x[0]) );
  DFF_X1 \addr_x_reg[1]  ( .D(N132), .CK(clk), .Q(addr_x[1]) );
  DFF_X1 clear_acc_reg ( .D(N146), .CK(clk), .Q(clear_acc) );
  DFF_X1 clc_reg ( .D(N147), .CK(clk), .Q(clc) );
  DFF_X1 clc1_reg ( .D(N148), .CK(clk), .Q(clc1) );
  NAND3_X1 U201 ( .A1(n127), .A2(n97), .A3(addr_a5[0]), .ZN(n129) );
  NAND3_X1 U202 ( .A1(n133), .A2(n121), .A3(n134), .ZN(n132) );
  NAND3_X1 U203 ( .A1(n137), .A2(n94), .A3(addr_a4[0]), .ZN(n139) );
  NAND3_X1 U204 ( .A1(n120), .A2(n119), .A3(n142), .ZN(n141) );
  NAND3_X1 U205 ( .A1(n145), .A2(n91), .A3(addr_a3[0]), .ZN(n147) );
  NAND3_X1 U206 ( .A1(n142), .A2(n120), .A3(n27), .ZN(n149) );
  NAND3_X1 U207 ( .A1(n153), .A2(n87), .A3(addr_a2[0]), .ZN(n155) );
  NAND3_X1 U208 ( .A1(n119), .A2(n118), .A3(n142), .ZN(n157) );
  NAND3_X1 U209 ( .A1(n162), .A2(n84), .A3(addr_a1[0]), .ZN(n164) );
  NAND3_X1 U210 ( .A1(n133), .A2(n167), .A3(n134), .ZN(n166) );
  NAND3_X1 U211 ( .A1(n178), .A2(n179), .A3(n31), .ZN(n175) );
  NAND3_X1 U212 ( .A1(addr_a8[1]), .A2(addr_a8[0]), .A3(addr_a8[2]), .ZN(n170)
         );
  NAND3_X1 U213 ( .A1(addr_a7[1]), .A2(addr_a7[0]), .A3(addr_a7[2]), .ZN(n195)
         );
  NAND3_X1 U214 ( .A1(addr_y[0]), .A2(n112), .A3(n216), .ZN(n218) );
  NAND3_X1 U215 ( .A1(n219), .A2(n30), .A3(addr_y[0]), .ZN(n220) );
  NAND3_X1 U216 ( .A1(addr_x[0]), .A2(n224), .A3(addr_x[1]), .ZN(n223) );
  NAND3_X1 U217 ( .A1(n228), .A2(n106), .A3(addr_a8[0]), .ZN(n230) );
  NAND3_X1 U218 ( .A1(n233), .A2(n172), .A3(n134), .ZN(n232) );
  NAND3_X1 U219 ( .A1(n236), .A2(n103), .A3(addr_a7[0]), .ZN(n238) );
  NAND3_X1 U220 ( .A1(n233), .A2(n173), .A3(n134), .ZN(n240) );
  NAND3_X1 U221 ( .A1(n123), .A2(n100), .A3(addr_a6[0]), .ZN(n244) );
  NAND3_X1 U222 ( .A1(n22), .A2(n158), .A3(n28), .ZN(n245) );
  NAND3_X1 U223 ( .A1(n119), .A2(n118), .A3(n120), .ZN(n246) );
  NAND3_X1 U224 ( .A1(addr_x[1]), .A2(addr_x[0]), .A3(addr_x[2]), .ZN(n205) );
  DFF_X1 \state_reg[4]  ( .D(n21), .CK(clk), .Q(state[4]), .QN(n76) );
  DFF_X1 \state_reg[2]  ( .D(N34), .CK(clk), .Q(state[2]), .QN(n79) );
  DFF_X1 \addr_y_reg[0]  ( .D(N141), .CK(clk), .Q(addr_y[0]), .QN(n113) );
  DFF_X1 \addr_y_reg[1]  ( .D(N142), .CK(clk), .Q(addr_y[1]), .QN(n112) );
  DFF_X1 \state_reg[1]  ( .D(N33), .CK(clk), .Q(state[1]), .QN(n80) );
  DFF_X1 \addr_y_reg[2]  ( .D(N143), .CK(clk), .Q(addr_y[2]), .QN(n111) );
  DFF_X1 \state_reg[0]  ( .D(N32), .CK(clk), .Q(state[0]), .QN(n81) );
  DFF_X1 \addr_x_reg[2]  ( .D(N133), .CK(clk), .Q(addr_x[2]), .QN(n108) );
  DFF_X1 \addr_a8_reg[0]  ( .D(n8), .CK(clk), .Q(addr_a8[0]), .QN(n107) );
  DFF_X1 \addr_a7_reg[0]  ( .D(n6), .CK(clk), .Q(addr_a7[0]), .QN(n104) );
  DFF_X1 \addr_a6_reg[0]  ( .D(n5), .CK(clk), .Q(addr_a6[0]), .QN(n101) );
  DFF_X1 \addr_a5_reg[0]  ( .D(n19), .CK(clk), .Q(addr_a5[0]), .QN(n98) );
  DFF_X1 \addr_a4_reg[0]  ( .D(n17), .CK(clk), .Q(addr_a4[0]), .QN(n95) );
  DFF_X1 \addr_a3_reg[0]  ( .D(n15), .CK(clk), .Q(addr_a3[0]), .QN(n92) );
  DFF_X1 \addr_a2_reg[0]  ( .D(n13), .CK(clk), .Q(addr_a2[0]), .QN(n88) );
  DFF_X1 \addr_a1_reg[0]  ( .D(n11), .CK(clk), .Q(addr_a1[0]), .QN(n85) );
  DFF_X1 \addr_a8_reg[1]  ( .D(N122), .CK(clk), .Q(addr_a8[1]), .QN(n106) );
  DFF_X1 \addr_a7_reg[1]  ( .D(N111), .CK(clk), .Q(addr_a7[1]), .QN(n103) );
  DFF_X1 \addr_a6_reg[1]  ( .D(N100), .CK(clk), .Q(addr_a6[1]), .QN(n100) );
  DFF_X1 \addr_a5_reg[1]  ( .D(N89), .CK(clk), .Q(addr_a5[1]), .QN(n97) );
  DFF_X1 \addr_a4_reg[1]  ( .D(N78), .CK(clk), .Q(addr_a4[1]), .QN(n94) );
  DFF_X1 \addr_a3_reg[1]  ( .D(N67), .CK(clk), .Q(addr_a3[1]), .QN(n91) );
  DFF_X1 \addr_a2_reg[1]  ( .D(N56), .CK(clk), .Q(addr_a2[1]), .QN(n87) );
  DFF_X1 \addr_a1_reg[1]  ( .D(N45), .CK(clk), .Q(addr_a1[1]), .QN(n84) );
  DFF_X1 \addr_a8_reg[2]  ( .D(N123), .CK(clk), .Q(addr_a8[2]), .QN(n105) );
  DFF_X1 \addr_a7_reg[2]  ( .D(N112), .CK(clk), .Q(addr_a7[2]), .QN(n102) );
  DFF_X1 \addr_a6_reg[2]  ( .D(N101), .CK(clk), .Q(addr_a6[2]), .QN(n99) );
  DFF_X1 \addr_a5_reg[2]  ( .D(N90), .CK(clk), .Q(addr_a5[2]), .QN(n96) );
  DFF_X1 \addr_a4_reg[2]  ( .D(N79), .CK(clk), .Q(addr_a4[2]), .QN(n93) );
  DFF_X1 \addr_a3_reg[2]  ( .D(N68), .CK(clk), .Q(addr_a3[2]), .QN(n90) );
  DFF_X1 \addr_a2_reg[2]  ( .D(N57), .CK(clk), .Q(addr_a2[2]), .QN(n86) );
  DFF_X1 \addr_a1_reg[2]  ( .D(N46), .CK(clk), .Q(addr_a1[2]), .QN(n83) );
  INV_X1 U3 ( .A(n248), .ZN(n22) );
  INV_X1 U4 ( .A(n224), .ZN(n10) );
  INV_X1 U5 ( .A(n246), .ZN(n28) );
  NAND2_X1 U6 ( .A1(n233), .A2(n133), .ZN(n248) );
  NAND2_X1 U7 ( .A1(n131), .A2(n245), .ZN(n123) );
  NAND2_X1 U8 ( .A1(n131), .A2(n149), .ZN(n145) );
  INV_X1 U9 ( .A(n150), .ZN(n27) );
  NAND2_X1 U10 ( .A1(n131), .A2(n157), .ZN(n153) );
  NAND2_X1 U11 ( .A1(n131), .A2(n141), .ZN(n137) );
  NAND2_X1 U12 ( .A1(n131), .A2(n132), .ZN(n127) );
  NAND2_X1 U13 ( .A1(n131), .A2(n166), .ZN(n162) );
  NOR2_X1 U14 ( .A1(n32), .A2(n23), .ZN(n133) );
  OAI21_X1 U15 ( .B1(n37), .B2(n117), .A(n131), .ZN(n224) );
  NAND2_X1 U16 ( .A1(n202), .A2(n116), .ZN(N148) );
  AND2_X1 U17 ( .A1(n207), .A2(n180), .ZN(n191) );
  NAND2_X1 U18 ( .A1(n117), .A2(n180), .ZN(N146) );
  AND2_X1 U19 ( .A1(n121), .A2(n167), .ZN(n233) );
  AND4_X1 U20 ( .A1(n247), .A2(n178), .A3(n210), .A4(n26), .ZN(n158) );
  INV_X1 U21 ( .A(N148), .ZN(n26) );
  INV_X1 U22 ( .A(n210), .ZN(n29) );
  OR2_X1 U23 ( .A1(n189), .A2(N37), .ZN(n188) );
  OAI211_X2 U24 ( .C1(n205), .C2(n210), .A(n116), .B(n178), .ZN(n124) );
  AOI21_X1 U25 ( .B1(n251), .B2(n33), .A(n189), .ZN(n178) );
  NAND4_X1 U26 ( .A1(n202), .A2(n159), .A3(n247), .A4(n249), .ZN(n131) );
  NOR3_X1 U27 ( .A1(n124), .A2(n248), .A3(n246), .ZN(n249) );
  NAND2_X1 U28 ( .A1(n222), .A2(n252), .ZN(n116) );
  NAND2_X1 U29 ( .A1(n254), .A2(n251), .ZN(n117) );
  OAI21_X1 U30 ( .B1(n119), .B2(n36), .A(n118), .ZN(n150) );
  INV_X1 U31 ( .A(n194), .ZN(n36) );
  NAND2_X1 U32 ( .A1(n254), .A2(n252), .ZN(n121) );
  NAND2_X1 U33 ( .A1(n131), .A2(n232), .ZN(n228) );
  NAND2_X1 U34 ( .A1(n131), .A2(n240), .ZN(n236) );
  NAND2_X1 U35 ( .A1(n250), .A2(n252), .ZN(n119) );
  NAND2_X1 U36 ( .A1(n255), .A2(n254), .ZN(n210) );
  NAND2_X1 U37 ( .A1(n255), .A2(n250), .ZN(n167) );
  NAND2_X1 U38 ( .A1(n250), .A2(n251), .ZN(n118) );
  NAND2_X1 U39 ( .A1(n251), .A2(n222), .ZN(n209) );
  NAND2_X1 U40 ( .A1(n221), .A2(n250), .ZN(n120) );
  NAND2_X1 U41 ( .A1(n33), .A2(n221), .ZN(n202) );
  INV_X1 U42 ( .A(n212), .ZN(n33) );
  NAND2_X1 U43 ( .A1(n33), .A2(n252), .ZN(n180) );
  NAND2_X1 U44 ( .A1(n255), .A2(n222), .ZN(n208) );
  INV_X1 U45 ( .A(n172), .ZN(n32) );
  NAND2_X1 U46 ( .A1(n221), .A2(n254), .ZN(n207) );
  AND3_X1 U47 ( .A1(n158), .A2(n159), .A3(n28), .ZN(n134) );
  AND4_X1 U48 ( .A1(n207), .A2(n25), .A3(n209), .A4(n256), .ZN(n247) );
  AND2_X1 U49 ( .A1(n208), .A2(n31), .ZN(n256) );
  INV_X1 U50 ( .A(N146), .ZN(n25) );
  AND3_X1 U51 ( .A1(n158), .A2(n159), .A3(n22), .ZN(n142) );
  AND2_X1 U52 ( .A1(n221), .A2(n222), .ZN(n189) );
  INV_X1 U53 ( .A(n173), .ZN(n23) );
  OAI221_X1 U54 ( .B1(n169), .B2(n167), .C1(n121), .C2(n35), .A(n28), .ZN(n177) );
  INV_X1 U55 ( .A(n184), .ZN(n35) );
  OAI22_X1 U56 ( .A1(n117), .A2(n205), .B1(n173), .B2(n170), .ZN(n176) );
  OAI22_X1 U57 ( .A1(n37), .A2(n117), .B1(n172), .B2(n195), .ZN(n192) );
  OAI22_X1 U58 ( .A1(n190), .A2(n116), .B1(n184), .B2(n121), .ZN(n204) );
  OAI21_X1 U59 ( .B1(n190), .B2(n208), .A(n209), .ZN(n183) );
  INV_X1 U60 ( .A(n205), .ZN(n37) );
  INV_X1 U61 ( .A(n216), .ZN(n30) );
  NOR2_X1 U62 ( .A1(n2), .A2(n116), .ZN(N37) );
  INV_X1 U63 ( .A(n190), .ZN(n2) );
  INV_X1 U64 ( .A(n222), .ZN(n34) );
  INV_X1 U65 ( .A(n193), .ZN(n3) );
  INV_X1 U66 ( .A(n168), .ZN(n21) );
  AOI221_X1 U67 ( .B1(n169), .B2(wr_en_a5), .C1(n170), .C2(wr_en_a8), .A(n171), 
        .ZN(n168) );
  OR2_X1 U68 ( .A1(wr_en_a7), .A2(wr_en_a6), .ZN(n171) );
  NOR3_X1 U69 ( .A1(state[0]), .A2(state[4]), .A3(n80), .ZN(n251) );
  NOR2_X1 U70 ( .A1(state[3]), .A2(state[2]), .ZN(n254) );
  NOR3_X1 U71 ( .A1(n81), .A2(state[4]), .A3(n80), .ZN(n255) );
  AOI211_X1 U72 ( .C1(n205), .C2(n29), .A(n183), .B(n206), .ZN(n193) );
  OAI22_X1 U73 ( .A1(n39), .A2(n191), .B1(n167), .B2(n169), .ZN(n206) );
  INV_X1 U74 ( .A(start), .ZN(n39) );
  NOR2_X1 U75 ( .A1(n79), .A2(state[3]), .ZN(n222) );
  NOR2_X1 U76 ( .A1(n211), .A2(state[0]), .ZN(n221) );
  NOR2_X1 U77 ( .A1(n81), .A2(n211), .ZN(n252) );
  NAND4_X1 U78 ( .A1(state[4]), .A2(n254), .A3(state[0]), .A4(n80), .ZN(n172)
         );
  AOI21_X1 U79 ( .B1(n101), .B2(n123), .A(n124), .ZN(n243) );
  AOI21_X1 U80 ( .B1(n92), .B2(n145), .A(n124), .ZN(n146) );
  AOI21_X1 U81 ( .B1(n88), .B2(n153), .A(n124), .ZN(n154) );
  AOI21_X1 U82 ( .B1(n95), .B2(n137), .A(n124), .ZN(n138) );
  AOI21_X1 U83 ( .B1(n98), .B2(n127), .A(n124), .ZN(n128) );
  AOI21_X1 U84 ( .B1(n85), .B2(n162), .A(n124), .ZN(n163) );
  AOI21_X1 U85 ( .B1(n107), .B2(n228), .A(n124), .ZN(n229) );
  AOI21_X1 U86 ( .B1(n104), .B2(n236), .A(n124), .ZN(n237) );
  NOR2_X1 U87 ( .A1(n173), .A2(reset), .ZN(wr_en_a8) );
  NOR2_X1 U88 ( .A1(n167), .A2(reset), .ZN(wr_en_a5) );
  NOR2_X1 U89 ( .A1(n172), .A2(reset), .ZN(wr_en_a7) );
  NAND2_X1 U90 ( .A1(n253), .A2(n80), .ZN(n159) );
  NOR2_X1 U91 ( .A1(n159), .A2(reset), .ZN(wr_en_a6) );
  NOR2_X1 U92 ( .A1(reset), .A2(n117), .ZN(wr_en_x) );
  NOR2_X1 U93 ( .A1(reset), .A2(n116), .ZN(wr_en_y) );
  NOR2_X1 U94 ( .A1(reset), .A2(n121), .ZN(wr_en_a1) );
  OAI211_X1 U95 ( .C1(loadVector), .C2(n180), .A(n24), .B(n193), .ZN(n203) );
  INV_X1 U96 ( .A(n176), .ZN(n24) );
  NOR2_X1 U97 ( .A1(reset), .A2(n118), .ZN(wr_en_a4) );
  NOR2_X1 U98 ( .A1(reset), .A2(n120), .ZN(wr_en_a2) );
  NOR2_X1 U99 ( .A1(reset), .A2(n119), .ZN(wr_en_a3) );
  AND2_X1 U100 ( .A1(state[3]), .A2(state[2]), .ZN(n250) );
  NAND2_X1 U101 ( .A1(n76), .A2(n80), .ZN(n211) );
  NAND2_X1 U102 ( .A1(n253), .A2(state[1]), .ZN(n173) );
  AOI21_X1 U103 ( .B1(n196), .B2(n197), .A(reset), .ZN(N32) );
  NOR4_X1 U104 ( .A1(n198), .A2(n199), .A3(n200), .A4(n201), .ZN(n197) );
  AOI211_X1 U105 ( .C1(n32), .C2(n195), .A(n203), .B(n204), .ZN(n196) );
  NOR4_X1 U106 ( .A1(n118), .A2(n95), .A3(n94), .A4(n93), .ZN(n201) );
  OAI21_X1 U107 ( .B1(n243), .B2(n100), .A(n244), .ZN(N100) );
  OAI21_X1 U108 ( .B1(n237), .B2(n103), .A(n238), .ZN(N111) );
  OAI21_X1 U109 ( .B1(n229), .B2(n106), .A(n230), .ZN(N122) );
  OAI21_X1 U110 ( .B1(n146), .B2(n91), .A(n147), .ZN(N67) );
  OAI21_X1 U111 ( .B1(n154), .B2(n87), .A(n155), .ZN(N56) );
  OAI21_X1 U112 ( .B1(n138), .B2(n94), .A(n139), .ZN(N78) );
  OAI21_X1 U113 ( .B1(n163), .B2(n84), .A(n164), .ZN(N45) );
  OAI21_X1 U114 ( .B1(n128), .B2(n97), .A(n129), .ZN(N89) );
  AND3_X1 U115 ( .A1(n254), .A2(n81), .A3(state[4]), .ZN(n253) );
  NAND2_X1 U116 ( .A1(state[3]), .A2(n79), .ZN(n212) );
  OAI21_X1 U117 ( .B1(n241), .B2(n99), .A(n242), .ZN(N101) );
  NAND4_X1 U118 ( .A1(addr_a6[1]), .A2(addr_a6[0]), .A3(n123), .A4(n99), .ZN(
        n242) );
  AOI21_X1 U119 ( .B1(n123), .B2(n100), .A(n4), .ZN(n241) );
  INV_X1 U120 ( .A(n243), .ZN(n4) );
  OAI21_X1 U121 ( .B1(n151), .B2(n86), .A(n152), .ZN(N57) );
  NAND4_X1 U122 ( .A1(addr_a2[1]), .A2(addr_a2[0]), .A3(n153), .A4(n86), .ZN(
        n152) );
  AOI21_X1 U123 ( .B1(n153), .B2(n87), .A(n14), .ZN(n151) );
  INV_X1 U124 ( .A(n154), .ZN(n14) );
  OAI21_X1 U125 ( .B1(n135), .B2(n93), .A(n136), .ZN(N79) );
  NAND4_X1 U126 ( .A1(addr_a4[1]), .A2(addr_a4[0]), .A3(n137), .A4(n93), .ZN(
        n136) );
  AOI21_X1 U127 ( .B1(n137), .B2(n94), .A(n18), .ZN(n135) );
  INV_X1 U128 ( .A(n138), .ZN(n18) );
  OAI21_X1 U129 ( .B1(n143), .B2(n90), .A(n144), .ZN(N68) );
  NAND4_X1 U130 ( .A1(addr_a3[1]), .A2(addr_a3[0]), .A3(n145), .A4(n90), .ZN(
        n144) );
  AOI21_X1 U131 ( .B1(n145), .B2(n91), .A(n16), .ZN(n143) );
  INV_X1 U132 ( .A(n146), .ZN(n16) );
  OAI21_X1 U133 ( .B1(n125), .B2(n96), .A(n126), .ZN(N90) );
  NAND4_X1 U134 ( .A1(addr_a5[1]), .A2(addr_a5[0]), .A3(n127), .A4(n96), .ZN(
        n126) );
  AOI21_X1 U135 ( .B1(n127), .B2(n97), .A(n20), .ZN(n125) );
  INV_X1 U136 ( .A(n128), .ZN(n20) );
  OAI21_X1 U137 ( .B1(n160), .B2(n83), .A(n161), .ZN(N46) );
  NAND4_X1 U138 ( .A1(addr_a1[1]), .A2(addr_a1[0]), .A3(n162), .A4(n83), .ZN(
        n161) );
  AOI21_X1 U139 ( .B1(n162), .B2(n84), .A(n12), .ZN(n160) );
  INV_X1 U140 ( .A(n163), .ZN(n12) );
  OAI21_X1 U141 ( .B1(n226), .B2(n105), .A(n227), .ZN(N123) );
  NAND4_X1 U142 ( .A1(addr_a8[1]), .A2(addr_a8[0]), .A3(n228), .A4(n105), .ZN(
        n227) );
  AOI21_X1 U143 ( .B1(n228), .B2(n106), .A(n9), .ZN(n226) );
  INV_X1 U144 ( .A(n229), .ZN(n9) );
  OAI21_X1 U145 ( .B1(n234), .B2(n102), .A(n235), .ZN(N112) );
  NAND4_X1 U146 ( .A1(addr_a7[1]), .A2(addr_a7[0]), .A3(n236), .A4(n102), .ZN(
        n235) );
  AOI21_X1 U147 ( .B1(n236), .B2(n103), .A(n7), .ZN(n234) );
  INV_X1 U148 ( .A(n237), .ZN(n7) );
  OAI21_X1 U149 ( .B1(n10), .B2(n108), .A(n223), .ZN(N133) );
  NOR2_X1 U150 ( .A1(addr_x[0]), .A2(n10), .ZN(N131) );
  NOR2_X1 U151 ( .A1(n10), .A2(n225), .ZN(N132) );
  XNOR2_X1 U152 ( .A(addr_x[1]), .B(addr_x[0]), .ZN(n225) );
  INV_X1 U153 ( .A(n257), .ZN(n31) );
  OAI21_X1 U154 ( .B1(n254), .B2(n76), .A(n258), .ZN(n257) );
  OAI211_X1 U155 ( .C1(n33), .C2(state[4]), .A(state[0]), .B(state[1]), .ZN(
        n258) );
  INV_X1 U156 ( .A(n122), .ZN(n5) );
  AOI22_X1 U157 ( .A1(n101), .A2(n123), .B1(n124), .B2(addr_a6[0]), .ZN(n122)
         );
  INV_X1 U158 ( .A(n148), .ZN(n15) );
  AOI22_X1 U159 ( .A1(n92), .A2(n145), .B1(n124), .B2(addr_a3[0]), .ZN(n148)
         );
  INV_X1 U160 ( .A(n156), .ZN(n13) );
  AOI22_X1 U161 ( .A1(n88), .A2(n153), .B1(n124), .B2(addr_a2[0]), .ZN(n156)
         );
  INV_X1 U162 ( .A(n140), .ZN(n17) );
  AOI22_X1 U163 ( .A1(n95), .A2(n137), .B1(n124), .B2(addr_a4[0]), .ZN(n140)
         );
  INV_X1 U164 ( .A(n130), .ZN(n19) );
  AOI22_X1 U165 ( .A1(n98), .A2(n127), .B1(n124), .B2(addr_a5[0]), .ZN(n130)
         );
  INV_X1 U166 ( .A(n165), .ZN(n11) );
  AOI22_X1 U167 ( .A1(n85), .A2(n162), .B1(n124), .B2(addr_a1[0]), .ZN(n165)
         );
  INV_X1 U168 ( .A(n231), .ZN(n8) );
  AOI22_X1 U169 ( .A1(n107), .A2(n228), .B1(n124), .B2(addr_a8[0]), .ZN(n231)
         );
  INV_X1 U170 ( .A(n239), .ZN(n6) );
  AOI22_X1 U171 ( .A1(n104), .A2(n236), .B1(n124), .B2(addr_a7[0]), .ZN(n239)
         );
  AOI211_X1 U172 ( .C1(n80), .C2(n81), .A(state[4]), .B(n34), .ZN(n216) );
  NOR3_X1 U173 ( .A1(n97), .A2(n98), .A3(n96), .ZN(n169) );
  NOR3_X1 U174 ( .A1(n112), .A2(n113), .A3(n111), .ZN(n190) );
  NOR4_X1 U175 ( .A1(n159), .A2(n101), .A3(n100), .A4(n99), .ZN(n200) );
  NOR4_X1 U176 ( .A1(n120), .A2(n88), .A3(n87), .A4(n86), .ZN(n199) );
  NOR3_X1 U177 ( .A1(n84), .A2(n85), .A3(n83), .ZN(n184) );
  NOR3_X1 U178 ( .A1(n91), .A2(n92), .A3(n90), .ZN(n194) );
  OAI221_X1 U179 ( .B1(n191), .B2(n38), .C1(n194), .C2(n119), .A(n202), .ZN(
        n198) );
  INV_X1 U180 ( .A(loadMatrix), .ZN(n38) );
  AOI22_X1 U181 ( .A1(n113), .A2(n216), .B1(n30), .B2(n219), .ZN(n217) );
  OAI22_X1 U182 ( .A1(n211), .A2(n34), .B1(n212), .B2(n213), .ZN(N147) );
  NAND2_X1 U183 ( .A1(n81), .A2(n76), .ZN(n213) );
  AOI21_X1 U184 ( .B1(n181), .B2(n182), .A(reset), .ZN(N34) );
  AOI21_X1 U185 ( .B1(n29), .B2(n37), .A(N148), .ZN(n182) );
  NOR2_X1 U186 ( .A1(n177), .A2(n183), .ZN(n181) );
  AOI21_X1 U187 ( .B1(n185), .B2(n186), .A(reset), .ZN(N33) );
  AOI221_X1 U188 ( .B1(n187), .B2(loadVector), .C1(n23), .C2(n170), .A(n188), 
        .ZN(n186) );
  NOR3_X1 U189 ( .A1(n192), .A2(n150), .A3(n3), .ZN(n185) );
  NOR2_X1 U190 ( .A1(loadMatrix), .A2(n191), .ZN(n187) );
  NAND2_X1 U191 ( .A1(n221), .A2(n79), .ZN(n219) );
  OAI21_X1 U192 ( .B1(n217), .B2(n112), .A(n218), .ZN(N142) );
  OAI21_X1 U193 ( .B1(n214), .B2(n111), .A(n215), .ZN(N143) );
  NAND4_X1 U194 ( .A1(n216), .A2(addr_y[1]), .A3(addr_y[0]), .A4(n111), .ZN(
        n215) );
  AOI21_X1 U195 ( .B1(n216), .B2(n112), .A(n1), .ZN(n214) );
  INV_X1 U196 ( .A(n217), .ZN(n1) );
  OAI21_X1 U197 ( .B1(addr_y[0]), .B2(n30), .A(n220), .ZN(N141) );
  NOR2_X1 U198 ( .A1(reset), .A2(n174), .ZN(N35) );
  NOR3_X1 U199 ( .A1(n175), .A2(n176), .A3(n177), .ZN(n174) );
  OR4_X1 U200 ( .A1(n180), .A2(loadMatrix), .A3(loadVector), .A4(start), .ZN(
        n179) );
endmodule


module mvm_8_8_20_1 ( clk, reset, loadMatrix, loadVector, start, done, data_in, 
        data_out );
  input [19:0] data_in;
  output [39:0] data_out;
  input clk, reset, loadMatrix, loadVector, start;
  output done;
  wire   wr_en_x, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6,
         wr_en_a7, wr_en_a8, wr_en_y, clear_acc, clc, clc1;
  wire   [2:0] addr_x;
  wire   [2:0] addr_a1;
  wire   [2:0] addr_a2;
  wire   [2:0] addr_a3;
  wire   [2:0] addr_a4;
  wire   [2:0] addr_a5;
  wire   [2:0] addr_a6;
  wire   [2:0] addr_a7;
  wire   [2:0] addr_a8;
  wire   [2:0] addr_y;

  datapath d ( .clk(clk), .data_in(data_in), .addr_x(addr_x), .wr_en_x(wr_en_x), .addr_a1(addr_a1), .addr_a2(addr_a2), .addr_a3(addr_a3), .addr_a4(addr_a4), 
        .addr_a5(addr_a5), .addr_a6(addr_a6), .addr_a7(addr_a7), .addr_a8(
        addr_a8), .wr_en_a1(wr_en_a1), .wr_en_a2(wr_en_a2), .wr_en_a3(wr_en_a3), .wr_en_a4(wr_en_a4), .wr_en_a5(wr_en_a5), .wr_en_a6(wr_en_a6), .wr_en_a7(
        wr_en_a7), .wr_en_a8(wr_en_a8), .addr_y(addr_y), .wr_en_y(wr_en_y), 
        .clear_acc(clear_acc), .clc(clc), .clc1(clc1), .data_out(data_out) );
  ctrlpath c ( .clk(clk), .reset(reset), .start(start), .addr_x(addr_x), 
        .wr_en_x(wr_en_x), .addr_a1(addr_a1), .addr_a2(addr_a2), .addr_a3(
        addr_a3), .addr_a4(addr_a4), .addr_a5(addr_a5), .addr_a6(addr_a6), 
        .addr_a7(addr_a7), .addr_a8(addr_a8), .wr_en_a1(wr_en_a1), .wr_en_a2(
        wr_en_a2), .wr_en_a3(wr_en_a3), .wr_en_a4(wr_en_a4), .wr_en_a5(
        wr_en_a5), .wr_en_a6(wr_en_a6), .wr_en_a7(wr_en_a7), .wr_en_a8(
        wr_en_a8), .clear_acc(clear_acc), .clc(clc), .clc1(clc1), .addr_y(
        addr_y), .wr_en_y(wr_en_y), .done(done), .loadMatrix(loadMatrix), 
        .loadVector(loadVector) );
endmodule

