
module memory_WIDTH8_SIZE16_LOGSIZE4_0 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N16), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n293), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n292), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n291), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n290), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n289), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n288), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n287), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n286), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n285), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n284), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n283), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n282), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n281), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n280), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n279), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n278), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n277), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n276), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n275), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n274), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n273), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n272), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n271), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n270), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n269), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n268), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n267), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n266), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n265), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n264), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n263), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n262), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n261), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n260), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n259), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n258), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n257), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n256), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n255), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n254), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n253), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n252), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n251), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n250), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n249), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n248), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n247), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n246), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n245), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n244), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n243), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n242), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n241), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n240), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n239), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n238), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n237), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n236), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n235), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n234), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n233), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n232), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n231), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n230), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n229), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n228), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n227), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n226), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n225), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n224), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n223), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n222), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n221), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n220), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n219), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n218), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n217), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n216), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n215), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n214), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n213), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n212), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n211), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n210), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n209), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n208), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n207), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n206), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n205), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n204), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n203), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n202), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n201), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n200), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n199), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n198), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n197), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n196), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n195), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n194), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n193), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n192), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n191), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n190), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n189), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n188), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n187), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n186), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n185), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n184), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n183), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n182), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n181), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n180), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n179), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n178), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n177), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n176), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n175), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n174), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n173), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n172), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n171), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n170), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n169), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n168), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n167), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n166), .CK(clk), .Q(\mem[0][0] ) );
  SDFF_X1 \data_out_reg[2]  ( .D(n324), .SI(n317), .SE(N13), .CK(clk), .Q(
        data_out[2]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n296), .SI(n7), .SE(N13), .CK(clk), .Q(
        data_out[0]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n310), .SI(n303), .SE(N13), .CK(clk), .Q(
        data_out[1]) );
  BUF_X1 U3 ( .A(N10), .Z(n397) );
  BUF_X1 U4 ( .A(N10), .Z(n398) );
  BUF_X1 U5 ( .A(N11), .Z(n395) );
  NAND2_X1 U6 ( .A1(n42), .A2(n22), .ZN(n33) );
  NAND2_X1 U7 ( .A1(n42), .A2(n32), .ZN(n43) );
  NAND2_X1 U8 ( .A1(n21), .A2(n22), .ZN(n12) );
  NAND2_X1 U9 ( .A1(n32), .A2(n21), .ZN(n23) );
  NAND2_X1 U10 ( .A1(n100), .A2(n21), .ZN(n91) );
  NAND2_X1 U11 ( .A1(n110), .A2(n21), .ZN(n101) );
  NAND2_X1 U12 ( .A1(n100), .A2(n42), .ZN(n111) );
  NAND2_X1 U13 ( .A1(n110), .A2(n42), .ZN(n120) );
  NAND2_X1 U14 ( .A1(n61), .A2(n22), .ZN(n52) );
  NAND2_X1 U15 ( .A1(n61), .A2(n32), .ZN(n62) );
  NAND2_X1 U16 ( .A1(n80), .A2(n22), .ZN(n71) );
  NAND2_X1 U17 ( .A1(n80), .A2(n32), .ZN(n82) );
  NAND2_X1 U18 ( .A1(n100), .A2(n61), .ZN(n129) );
  NAND2_X1 U19 ( .A1(n110), .A2(n61), .ZN(n138) );
  NAND2_X1 U20 ( .A1(n100), .A2(n80), .ZN(n147) );
  NAND2_X1 U21 ( .A1(n110), .A2(n80), .ZN(n157) );
  AND2_X1 U22 ( .A1(n156), .A2(N10), .ZN(n110) );
  AND2_X1 U23 ( .A1(n156), .A2(n399), .ZN(n100) );
  AND2_X1 U24 ( .A1(N10), .A2(n81), .ZN(n32) );
  AND2_X1 U25 ( .A1(n81), .A2(n399), .ZN(n22) );
  OAI21_X1 U26 ( .B1(n12), .B2(n409), .A(n13), .ZN(n166) );
  NAND2_X1 U27 ( .A1(\mem[0][0] ), .A2(n12), .ZN(n13) );
  OAI21_X1 U28 ( .B1(n12), .B2(n408), .A(n14), .ZN(n167) );
  NAND2_X1 U29 ( .A1(\mem[0][1] ), .A2(n12), .ZN(n14) );
  OAI21_X1 U30 ( .B1(n12), .B2(n407), .A(n15), .ZN(n168) );
  NAND2_X1 U31 ( .A1(\mem[0][2] ), .A2(n12), .ZN(n15) );
  OAI21_X1 U32 ( .B1(n12), .B2(n406), .A(n16), .ZN(n169) );
  NAND2_X1 U33 ( .A1(\mem[0][3] ), .A2(n12), .ZN(n16) );
  OAI21_X1 U34 ( .B1(n12), .B2(n405), .A(n17), .ZN(n170) );
  NAND2_X1 U35 ( .A1(\mem[0][4] ), .A2(n12), .ZN(n17) );
  OAI21_X1 U36 ( .B1(n12), .B2(n404), .A(n18), .ZN(n171) );
  NAND2_X1 U37 ( .A1(\mem[0][5] ), .A2(n12), .ZN(n18) );
  OAI21_X1 U38 ( .B1(n12), .B2(n403), .A(n19), .ZN(n172) );
  NAND2_X1 U39 ( .A1(\mem[0][6] ), .A2(n12), .ZN(n19) );
  OAI21_X1 U40 ( .B1(n12), .B2(n402), .A(n20), .ZN(n173) );
  NAND2_X1 U41 ( .A1(\mem[0][7] ), .A2(n12), .ZN(n20) );
  OAI21_X1 U42 ( .B1(n409), .B2(n33), .A(n34), .ZN(n182) );
  NAND2_X1 U43 ( .A1(\mem[2][0] ), .A2(n33), .ZN(n34) );
  OAI21_X1 U44 ( .B1(n408), .B2(n33), .A(n35), .ZN(n183) );
  NAND2_X1 U45 ( .A1(\mem[2][1] ), .A2(n33), .ZN(n35) );
  OAI21_X1 U46 ( .B1(n407), .B2(n33), .A(n36), .ZN(n184) );
  NAND2_X1 U47 ( .A1(\mem[2][2] ), .A2(n33), .ZN(n36) );
  OAI21_X1 U48 ( .B1(n406), .B2(n33), .A(n37), .ZN(n185) );
  NAND2_X1 U49 ( .A1(\mem[2][3] ), .A2(n33), .ZN(n37) );
  OAI21_X1 U50 ( .B1(n405), .B2(n33), .A(n38), .ZN(n186) );
  NAND2_X1 U51 ( .A1(\mem[2][4] ), .A2(n33), .ZN(n38) );
  OAI21_X1 U52 ( .B1(n404), .B2(n33), .A(n39), .ZN(n187) );
  NAND2_X1 U53 ( .A1(\mem[2][5] ), .A2(n33), .ZN(n39) );
  OAI21_X1 U54 ( .B1(n403), .B2(n33), .A(n40), .ZN(n188) );
  NAND2_X1 U55 ( .A1(\mem[2][6] ), .A2(n33), .ZN(n40) );
  OAI21_X1 U56 ( .B1(n402), .B2(n33), .A(n41), .ZN(n189) );
  NAND2_X1 U57 ( .A1(\mem[2][7] ), .A2(n33), .ZN(n41) );
  OAI21_X1 U58 ( .B1(n409), .B2(n43), .A(n44), .ZN(n190) );
  NAND2_X1 U59 ( .A1(\mem[3][0] ), .A2(n43), .ZN(n44) );
  OAI21_X1 U60 ( .B1(n408), .B2(n43), .A(n45), .ZN(n191) );
  NAND2_X1 U61 ( .A1(\mem[3][1] ), .A2(n43), .ZN(n45) );
  OAI21_X1 U62 ( .B1(n407), .B2(n43), .A(n46), .ZN(n192) );
  NAND2_X1 U63 ( .A1(\mem[3][2] ), .A2(n43), .ZN(n46) );
  OAI21_X1 U64 ( .B1(n406), .B2(n43), .A(n47), .ZN(n193) );
  NAND2_X1 U65 ( .A1(\mem[3][3] ), .A2(n43), .ZN(n47) );
  OAI21_X1 U66 ( .B1(n405), .B2(n43), .A(n48), .ZN(n194) );
  NAND2_X1 U67 ( .A1(\mem[3][4] ), .A2(n43), .ZN(n48) );
  OAI21_X1 U68 ( .B1(n404), .B2(n43), .A(n49), .ZN(n195) );
  NAND2_X1 U69 ( .A1(\mem[3][5] ), .A2(n43), .ZN(n49) );
  OAI21_X1 U70 ( .B1(n403), .B2(n43), .A(n50), .ZN(n196) );
  NAND2_X1 U71 ( .A1(\mem[3][6] ), .A2(n43), .ZN(n50) );
  OAI21_X1 U72 ( .B1(n402), .B2(n43), .A(n51), .ZN(n197) );
  NAND2_X1 U73 ( .A1(\mem[3][7] ), .A2(n43), .ZN(n51) );
  NOR2_X1 U74 ( .A1(n401), .A2(N13), .ZN(n81) );
  INV_X1 U75 ( .A(wr_en), .ZN(n401) );
  OAI21_X1 U76 ( .B1(n409), .B2(n23), .A(n24), .ZN(n174) );
  NAND2_X1 U77 ( .A1(\mem[1][0] ), .A2(n23), .ZN(n24) );
  OAI21_X1 U78 ( .B1(n408), .B2(n23), .A(n25), .ZN(n175) );
  NAND2_X1 U79 ( .A1(\mem[1][1] ), .A2(n23), .ZN(n25) );
  OAI21_X1 U80 ( .B1(n407), .B2(n23), .A(n26), .ZN(n176) );
  NAND2_X1 U81 ( .A1(\mem[1][2] ), .A2(n23), .ZN(n26) );
  OAI21_X1 U82 ( .B1(n406), .B2(n23), .A(n27), .ZN(n177) );
  NAND2_X1 U83 ( .A1(\mem[1][3] ), .A2(n23), .ZN(n27) );
  OAI21_X1 U84 ( .B1(n405), .B2(n23), .A(n28), .ZN(n178) );
  NAND2_X1 U85 ( .A1(\mem[1][4] ), .A2(n23), .ZN(n28) );
  OAI21_X1 U86 ( .B1(n404), .B2(n23), .A(n29), .ZN(n179) );
  NAND2_X1 U87 ( .A1(\mem[1][5] ), .A2(n23), .ZN(n29) );
  OAI21_X1 U88 ( .B1(n403), .B2(n23), .A(n30), .ZN(n180) );
  NAND2_X1 U89 ( .A1(\mem[1][6] ), .A2(n23), .ZN(n30) );
  OAI21_X1 U90 ( .B1(n402), .B2(n23), .A(n31), .ZN(n181) );
  NAND2_X1 U91 ( .A1(\mem[1][7] ), .A2(n23), .ZN(n31) );
  OAI21_X1 U92 ( .B1(n409), .B2(n52), .A(n53), .ZN(n198) );
  NAND2_X1 U93 ( .A1(\mem[4][0] ), .A2(n52), .ZN(n53) );
  OAI21_X1 U94 ( .B1(n408), .B2(n52), .A(n54), .ZN(n199) );
  NAND2_X1 U95 ( .A1(\mem[4][1] ), .A2(n52), .ZN(n54) );
  OAI21_X1 U96 ( .B1(n407), .B2(n52), .A(n55), .ZN(n200) );
  NAND2_X1 U97 ( .A1(\mem[4][2] ), .A2(n52), .ZN(n55) );
  OAI21_X1 U98 ( .B1(n406), .B2(n52), .A(n56), .ZN(n201) );
  NAND2_X1 U99 ( .A1(\mem[4][3] ), .A2(n52), .ZN(n56) );
  OAI21_X1 U100 ( .B1(n405), .B2(n52), .A(n57), .ZN(n202) );
  NAND2_X1 U101 ( .A1(\mem[4][4] ), .A2(n52), .ZN(n57) );
  OAI21_X1 U102 ( .B1(n404), .B2(n52), .A(n58), .ZN(n203) );
  NAND2_X1 U103 ( .A1(\mem[4][5] ), .A2(n52), .ZN(n58) );
  OAI21_X1 U104 ( .B1(n403), .B2(n52), .A(n59), .ZN(n204) );
  NAND2_X1 U105 ( .A1(\mem[4][6] ), .A2(n52), .ZN(n59) );
  OAI21_X1 U106 ( .B1(n402), .B2(n52), .A(n60), .ZN(n205) );
  NAND2_X1 U107 ( .A1(\mem[4][7] ), .A2(n52), .ZN(n60) );
  OAI21_X1 U108 ( .B1(n409), .B2(n62), .A(n63), .ZN(n206) );
  NAND2_X1 U109 ( .A1(\mem[5][0] ), .A2(n62), .ZN(n63) );
  OAI21_X1 U110 ( .B1(n408), .B2(n62), .A(n64), .ZN(n207) );
  NAND2_X1 U111 ( .A1(\mem[5][1] ), .A2(n62), .ZN(n64) );
  OAI21_X1 U112 ( .B1(n407), .B2(n62), .A(n65), .ZN(n208) );
  NAND2_X1 U113 ( .A1(\mem[5][2] ), .A2(n62), .ZN(n65) );
  OAI21_X1 U114 ( .B1(n406), .B2(n62), .A(n66), .ZN(n209) );
  NAND2_X1 U115 ( .A1(\mem[5][3] ), .A2(n62), .ZN(n66) );
  OAI21_X1 U116 ( .B1(n405), .B2(n62), .A(n67), .ZN(n210) );
  NAND2_X1 U117 ( .A1(\mem[5][4] ), .A2(n62), .ZN(n67) );
  OAI21_X1 U118 ( .B1(n404), .B2(n62), .A(n68), .ZN(n211) );
  NAND2_X1 U119 ( .A1(\mem[5][5] ), .A2(n62), .ZN(n68) );
  OAI21_X1 U120 ( .B1(n403), .B2(n62), .A(n69), .ZN(n212) );
  NAND2_X1 U121 ( .A1(\mem[5][6] ), .A2(n62), .ZN(n69) );
  OAI21_X1 U122 ( .B1(n402), .B2(n62), .A(n70), .ZN(n213) );
  NAND2_X1 U123 ( .A1(\mem[5][7] ), .A2(n62), .ZN(n70) );
  OAI21_X1 U124 ( .B1(n409), .B2(n71), .A(n72), .ZN(n214) );
  NAND2_X1 U125 ( .A1(\mem[6][0] ), .A2(n71), .ZN(n72) );
  OAI21_X1 U126 ( .B1(n408), .B2(n71), .A(n73), .ZN(n215) );
  NAND2_X1 U127 ( .A1(\mem[6][1] ), .A2(n71), .ZN(n73) );
  OAI21_X1 U128 ( .B1(n407), .B2(n71), .A(n74), .ZN(n216) );
  NAND2_X1 U129 ( .A1(\mem[6][2] ), .A2(n71), .ZN(n74) );
  OAI21_X1 U130 ( .B1(n406), .B2(n71), .A(n75), .ZN(n217) );
  NAND2_X1 U131 ( .A1(\mem[6][3] ), .A2(n71), .ZN(n75) );
  OAI21_X1 U132 ( .B1(n405), .B2(n71), .A(n76), .ZN(n218) );
  NAND2_X1 U133 ( .A1(\mem[6][4] ), .A2(n71), .ZN(n76) );
  OAI21_X1 U134 ( .B1(n404), .B2(n71), .A(n77), .ZN(n219) );
  NAND2_X1 U135 ( .A1(\mem[6][5] ), .A2(n71), .ZN(n77) );
  OAI21_X1 U136 ( .B1(n403), .B2(n71), .A(n78), .ZN(n220) );
  NAND2_X1 U137 ( .A1(\mem[6][6] ), .A2(n71), .ZN(n78) );
  OAI21_X1 U138 ( .B1(n402), .B2(n71), .A(n79), .ZN(n221) );
  NAND2_X1 U139 ( .A1(\mem[6][7] ), .A2(n71), .ZN(n79) );
  OAI21_X1 U140 ( .B1(n409), .B2(n82), .A(n83), .ZN(n222) );
  NAND2_X1 U141 ( .A1(\mem[7][0] ), .A2(n82), .ZN(n83) );
  OAI21_X1 U142 ( .B1(n408), .B2(n82), .A(n84), .ZN(n223) );
  NAND2_X1 U143 ( .A1(\mem[7][1] ), .A2(n82), .ZN(n84) );
  OAI21_X1 U144 ( .B1(n407), .B2(n82), .A(n85), .ZN(n224) );
  NAND2_X1 U145 ( .A1(\mem[7][2] ), .A2(n82), .ZN(n85) );
  OAI21_X1 U146 ( .B1(n406), .B2(n82), .A(n86), .ZN(n225) );
  NAND2_X1 U147 ( .A1(\mem[7][3] ), .A2(n82), .ZN(n86) );
  OAI21_X1 U148 ( .B1(n405), .B2(n82), .A(n87), .ZN(n226) );
  NAND2_X1 U149 ( .A1(\mem[7][4] ), .A2(n82), .ZN(n87) );
  OAI21_X1 U150 ( .B1(n404), .B2(n82), .A(n88), .ZN(n227) );
  NAND2_X1 U151 ( .A1(\mem[7][5] ), .A2(n82), .ZN(n88) );
  OAI21_X1 U152 ( .B1(n403), .B2(n82), .A(n89), .ZN(n228) );
  NAND2_X1 U153 ( .A1(\mem[7][6] ), .A2(n82), .ZN(n89) );
  OAI21_X1 U154 ( .B1(n402), .B2(n82), .A(n90), .ZN(n229) );
  NAND2_X1 U155 ( .A1(\mem[7][7] ), .A2(n82), .ZN(n90) );
  OAI21_X1 U156 ( .B1(n409), .B2(n91), .A(n92), .ZN(n230) );
  NAND2_X1 U157 ( .A1(\mem[8][0] ), .A2(n91), .ZN(n92) );
  OAI21_X1 U158 ( .B1(n408), .B2(n91), .A(n93), .ZN(n231) );
  NAND2_X1 U159 ( .A1(\mem[8][1] ), .A2(n91), .ZN(n93) );
  OAI21_X1 U160 ( .B1(n407), .B2(n91), .A(n94), .ZN(n232) );
  NAND2_X1 U161 ( .A1(\mem[8][2] ), .A2(n91), .ZN(n94) );
  OAI21_X1 U162 ( .B1(n406), .B2(n91), .A(n95), .ZN(n233) );
  NAND2_X1 U163 ( .A1(\mem[8][3] ), .A2(n91), .ZN(n95) );
  OAI21_X1 U164 ( .B1(n405), .B2(n91), .A(n96), .ZN(n234) );
  NAND2_X1 U165 ( .A1(\mem[8][4] ), .A2(n91), .ZN(n96) );
  OAI21_X1 U166 ( .B1(n404), .B2(n91), .A(n97), .ZN(n235) );
  NAND2_X1 U167 ( .A1(\mem[8][5] ), .A2(n91), .ZN(n97) );
  OAI21_X1 U168 ( .B1(n403), .B2(n91), .A(n98), .ZN(n236) );
  NAND2_X1 U169 ( .A1(\mem[8][6] ), .A2(n91), .ZN(n98) );
  OAI21_X1 U170 ( .B1(n402), .B2(n91), .A(n99), .ZN(n237) );
  NAND2_X1 U171 ( .A1(\mem[8][7] ), .A2(n91), .ZN(n99) );
  OAI21_X1 U172 ( .B1(n409), .B2(n101), .A(n102), .ZN(n238) );
  NAND2_X1 U173 ( .A1(\mem[9][0] ), .A2(n101), .ZN(n102) );
  OAI21_X1 U174 ( .B1(n408), .B2(n101), .A(n103), .ZN(n239) );
  NAND2_X1 U175 ( .A1(\mem[9][1] ), .A2(n101), .ZN(n103) );
  OAI21_X1 U176 ( .B1(n407), .B2(n101), .A(n104), .ZN(n240) );
  NAND2_X1 U177 ( .A1(\mem[9][2] ), .A2(n101), .ZN(n104) );
  OAI21_X1 U178 ( .B1(n406), .B2(n101), .A(n105), .ZN(n241) );
  NAND2_X1 U179 ( .A1(\mem[9][3] ), .A2(n101), .ZN(n105) );
  OAI21_X1 U180 ( .B1(n405), .B2(n101), .A(n106), .ZN(n242) );
  NAND2_X1 U181 ( .A1(\mem[9][4] ), .A2(n101), .ZN(n106) );
  OAI21_X1 U182 ( .B1(n404), .B2(n101), .A(n107), .ZN(n243) );
  NAND2_X1 U183 ( .A1(\mem[9][5] ), .A2(n101), .ZN(n107) );
  OAI21_X1 U184 ( .B1(n403), .B2(n101), .A(n108), .ZN(n244) );
  NAND2_X1 U185 ( .A1(\mem[9][6] ), .A2(n101), .ZN(n108) );
  OAI21_X1 U186 ( .B1(n402), .B2(n101), .A(n109), .ZN(n245) );
  NAND2_X1 U187 ( .A1(\mem[9][7] ), .A2(n101), .ZN(n109) );
  OAI21_X1 U188 ( .B1(n409), .B2(n111), .A(n112), .ZN(n246) );
  NAND2_X1 U189 ( .A1(\mem[10][0] ), .A2(n111), .ZN(n112) );
  OAI21_X1 U190 ( .B1(n408), .B2(n111), .A(n113), .ZN(n247) );
  NAND2_X1 U191 ( .A1(\mem[10][1] ), .A2(n111), .ZN(n113) );
  OAI21_X1 U192 ( .B1(n407), .B2(n111), .A(n114), .ZN(n248) );
  NAND2_X1 U193 ( .A1(\mem[10][2] ), .A2(n111), .ZN(n114) );
  OAI21_X1 U194 ( .B1(n406), .B2(n111), .A(n115), .ZN(n249) );
  NAND2_X1 U195 ( .A1(\mem[10][3] ), .A2(n111), .ZN(n115) );
  OAI21_X1 U196 ( .B1(n405), .B2(n111), .A(n116), .ZN(n250) );
  NAND2_X1 U197 ( .A1(\mem[10][4] ), .A2(n111), .ZN(n116) );
  OAI21_X1 U198 ( .B1(n404), .B2(n111), .A(n117), .ZN(n251) );
  NAND2_X1 U199 ( .A1(\mem[10][5] ), .A2(n111), .ZN(n117) );
  OAI21_X1 U200 ( .B1(n403), .B2(n111), .A(n118), .ZN(n252) );
  NAND2_X1 U201 ( .A1(\mem[10][6] ), .A2(n111), .ZN(n118) );
  OAI21_X1 U202 ( .B1(n402), .B2(n111), .A(n119), .ZN(n253) );
  NAND2_X1 U203 ( .A1(\mem[10][7] ), .A2(n111), .ZN(n119) );
  OAI21_X1 U204 ( .B1(n409), .B2(n120), .A(n121), .ZN(n254) );
  NAND2_X1 U205 ( .A1(\mem[11][0] ), .A2(n120), .ZN(n121) );
  OAI21_X1 U206 ( .B1(n408), .B2(n120), .A(n122), .ZN(n255) );
  NAND2_X1 U207 ( .A1(\mem[11][1] ), .A2(n120), .ZN(n122) );
  OAI21_X1 U208 ( .B1(n407), .B2(n120), .A(n123), .ZN(n256) );
  NAND2_X1 U209 ( .A1(\mem[11][2] ), .A2(n120), .ZN(n123) );
  OAI21_X1 U210 ( .B1(n406), .B2(n120), .A(n124), .ZN(n257) );
  NAND2_X1 U211 ( .A1(\mem[11][3] ), .A2(n120), .ZN(n124) );
  OAI21_X1 U212 ( .B1(n405), .B2(n120), .A(n125), .ZN(n258) );
  NAND2_X1 U213 ( .A1(\mem[11][4] ), .A2(n120), .ZN(n125) );
  OAI21_X1 U214 ( .B1(n404), .B2(n120), .A(n126), .ZN(n259) );
  NAND2_X1 U215 ( .A1(\mem[11][5] ), .A2(n120), .ZN(n126) );
  OAI21_X1 U216 ( .B1(n403), .B2(n120), .A(n127), .ZN(n260) );
  NAND2_X1 U217 ( .A1(\mem[11][6] ), .A2(n120), .ZN(n127) );
  OAI21_X1 U218 ( .B1(n402), .B2(n120), .A(n128), .ZN(n261) );
  NAND2_X1 U219 ( .A1(\mem[11][7] ), .A2(n120), .ZN(n128) );
  OAI21_X1 U220 ( .B1(n409), .B2(n129), .A(n130), .ZN(n262) );
  NAND2_X1 U221 ( .A1(\mem[12][0] ), .A2(n129), .ZN(n130) );
  OAI21_X1 U222 ( .B1(n408), .B2(n129), .A(n131), .ZN(n263) );
  NAND2_X1 U223 ( .A1(\mem[12][1] ), .A2(n129), .ZN(n131) );
  OAI21_X1 U224 ( .B1(n407), .B2(n129), .A(n132), .ZN(n264) );
  NAND2_X1 U225 ( .A1(\mem[12][2] ), .A2(n129), .ZN(n132) );
  OAI21_X1 U226 ( .B1(n406), .B2(n129), .A(n133), .ZN(n265) );
  NAND2_X1 U227 ( .A1(\mem[12][3] ), .A2(n129), .ZN(n133) );
  OAI21_X1 U228 ( .B1(n405), .B2(n129), .A(n134), .ZN(n266) );
  NAND2_X1 U229 ( .A1(\mem[12][4] ), .A2(n129), .ZN(n134) );
  OAI21_X1 U230 ( .B1(n404), .B2(n129), .A(n135), .ZN(n267) );
  NAND2_X1 U231 ( .A1(\mem[12][5] ), .A2(n129), .ZN(n135) );
  OAI21_X1 U232 ( .B1(n403), .B2(n129), .A(n136), .ZN(n268) );
  NAND2_X1 U233 ( .A1(\mem[12][6] ), .A2(n129), .ZN(n136) );
  OAI21_X1 U234 ( .B1(n402), .B2(n129), .A(n137), .ZN(n269) );
  NAND2_X1 U235 ( .A1(\mem[12][7] ), .A2(n129), .ZN(n137) );
  OAI21_X1 U236 ( .B1(n409), .B2(n138), .A(n139), .ZN(n270) );
  NAND2_X1 U237 ( .A1(\mem[13][0] ), .A2(n138), .ZN(n139) );
  OAI21_X1 U238 ( .B1(n408), .B2(n138), .A(n140), .ZN(n271) );
  NAND2_X1 U239 ( .A1(\mem[13][1] ), .A2(n138), .ZN(n140) );
  OAI21_X1 U240 ( .B1(n407), .B2(n138), .A(n141), .ZN(n272) );
  NAND2_X1 U241 ( .A1(\mem[13][2] ), .A2(n138), .ZN(n141) );
  OAI21_X1 U242 ( .B1(n406), .B2(n138), .A(n142), .ZN(n273) );
  NAND2_X1 U243 ( .A1(\mem[13][3] ), .A2(n138), .ZN(n142) );
  OAI21_X1 U244 ( .B1(n405), .B2(n138), .A(n143), .ZN(n274) );
  NAND2_X1 U245 ( .A1(\mem[13][4] ), .A2(n138), .ZN(n143) );
  OAI21_X1 U246 ( .B1(n404), .B2(n138), .A(n144), .ZN(n275) );
  NAND2_X1 U247 ( .A1(\mem[13][5] ), .A2(n138), .ZN(n144) );
  OAI21_X1 U248 ( .B1(n403), .B2(n138), .A(n145), .ZN(n276) );
  NAND2_X1 U249 ( .A1(\mem[13][6] ), .A2(n138), .ZN(n145) );
  OAI21_X1 U250 ( .B1(n402), .B2(n138), .A(n146), .ZN(n277) );
  NAND2_X1 U251 ( .A1(\mem[13][7] ), .A2(n138), .ZN(n146) );
  OAI21_X1 U252 ( .B1(n409), .B2(n147), .A(n148), .ZN(n278) );
  NAND2_X1 U253 ( .A1(\mem[14][0] ), .A2(n147), .ZN(n148) );
  OAI21_X1 U254 ( .B1(n408), .B2(n147), .A(n149), .ZN(n279) );
  NAND2_X1 U255 ( .A1(\mem[14][1] ), .A2(n147), .ZN(n149) );
  OAI21_X1 U256 ( .B1(n407), .B2(n147), .A(n150), .ZN(n280) );
  NAND2_X1 U257 ( .A1(\mem[14][2] ), .A2(n147), .ZN(n150) );
  OAI21_X1 U258 ( .B1(n406), .B2(n147), .A(n151), .ZN(n281) );
  NAND2_X1 U259 ( .A1(\mem[14][3] ), .A2(n147), .ZN(n151) );
  OAI21_X1 U260 ( .B1(n405), .B2(n147), .A(n152), .ZN(n282) );
  NAND2_X1 U261 ( .A1(\mem[14][4] ), .A2(n147), .ZN(n152) );
  OAI21_X1 U262 ( .B1(n404), .B2(n147), .A(n153), .ZN(n283) );
  NAND2_X1 U263 ( .A1(\mem[14][5] ), .A2(n147), .ZN(n153) );
  OAI21_X1 U264 ( .B1(n403), .B2(n147), .A(n154), .ZN(n284) );
  NAND2_X1 U265 ( .A1(\mem[14][6] ), .A2(n147), .ZN(n154) );
  OAI21_X1 U266 ( .B1(n402), .B2(n147), .A(n155), .ZN(n285) );
  NAND2_X1 U267 ( .A1(\mem[14][7] ), .A2(n147), .ZN(n155) );
  OAI21_X1 U268 ( .B1(n409), .B2(n157), .A(n158), .ZN(n286) );
  NAND2_X1 U269 ( .A1(\mem[15][0] ), .A2(n157), .ZN(n158) );
  OAI21_X1 U270 ( .B1(n408), .B2(n157), .A(n159), .ZN(n287) );
  NAND2_X1 U271 ( .A1(\mem[15][1] ), .A2(n157), .ZN(n159) );
  OAI21_X1 U272 ( .B1(n407), .B2(n157), .A(n160), .ZN(n288) );
  NAND2_X1 U273 ( .A1(\mem[15][2] ), .A2(n157), .ZN(n160) );
  OAI21_X1 U274 ( .B1(n406), .B2(n157), .A(n161), .ZN(n289) );
  NAND2_X1 U275 ( .A1(\mem[15][3] ), .A2(n157), .ZN(n161) );
  OAI21_X1 U276 ( .B1(n405), .B2(n157), .A(n162), .ZN(n290) );
  NAND2_X1 U277 ( .A1(\mem[15][4] ), .A2(n157), .ZN(n162) );
  OAI21_X1 U278 ( .B1(n404), .B2(n157), .A(n163), .ZN(n291) );
  NAND2_X1 U279 ( .A1(\mem[15][5] ), .A2(n157), .ZN(n163) );
  OAI21_X1 U280 ( .B1(n403), .B2(n157), .A(n164), .ZN(n292) );
  NAND2_X1 U281 ( .A1(\mem[15][6] ), .A2(n157), .ZN(n164) );
  OAI21_X1 U282 ( .B1(n402), .B2(n157), .A(n165), .ZN(n293) );
  NAND2_X1 U283 ( .A1(\mem[15][7] ), .A2(n157), .ZN(n165) );
  AND2_X1 U284 ( .A1(N13), .A2(wr_en), .ZN(n156) );
  NOR2_X1 U285 ( .A1(N11), .A2(N12), .ZN(n21) );
  NOR2_X1 U286 ( .A1(n400), .A2(N12), .ZN(n42) );
  AND2_X1 U287 ( .A1(N12), .A2(n400), .ZN(n61) );
  AND2_X1 U288 ( .A1(N12), .A2(N11), .ZN(n80) );
  INV_X1 U289 ( .A(data_in[0]), .ZN(n409) );
  INV_X1 U290 ( .A(data_in[1]), .ZN(n408) );
  INV_X1 U291 ( .A(data_in[2]), .ZN(n407) );
  INV_X1 U292 ( .A(data_in[3]), .ZN(n406) );
  INV_X1 U293 ( .A(data_in[4]), .ZN(n405) );
  INV_X1 U294 ( .A(data_in[5]), .ZN(n404) );
  INV_X1 U295 ( .A(data_in[6]), .ZN(n403) );
  INV_X1 U296 ( .A(data_in[7]), .ZN(n402) );
  MUX2_X1 U297 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n396), .Z(n1) );
  MUX2_X1 U298 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n396), .Z(n2) );
  MUX2_X1 U299 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U300 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n396), .Z(n4) );
  MUX2_X1 U301 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n396), .Z(n5) );
  MUX2_X1 U302 ( .A(n5), .B(n4), .S(N11), .Z(n6) );
  MUX2_X1 U303 ( .A(n6), .B(n3), .S(N12), .Z(n7) );
  MUX2_X1 U304 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n397), .Z(n8) );
  MUX2_X1 U305 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n396), .Z(n9) );
  MUX2_X1 U306 ( .A(n9), .B(n8), .S(N11), .Z(n10) );
  MUX2_X1 U307 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n398), .Z(n11) );
  MUX2_X1 U308 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n397), .Z(n294) );
  MUX2_X1 U309 ( .A(n294), .B(n11), .S(N11), .Z(n295) );
  MUX2_X1 U310 ( .A(n295), .B(n10), .S(N12), .Z(n296) );
  MUX2_X1 U311 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n397), .Z(n297) );
  MUX2_X1 U312 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n396), .Z(n298) );
  MUX2_X1 U313 ( .A(n298), .B(n297), .S(N11), .Z(n299) );
  MUX2_X1 U314 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(N10), .Z(n300) );
  MUX2_X1 U315 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n398), .Z(n301) );
  MUX2_X1 U316 ( .A(n301), .B(n300), .S(N11), .Z(n302) );
  MUX2_X1 U317 ( .A(n302), .B(n299), .S(N12), .Z(n303) );
  MUX2_X1 U318 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n396), .Z(n304) );
  MUX2_X1 U319 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n398), .Z(n305) );
  MUX2_X1 U320 ( .A(n305), .B(n304), .S(N11), .Z(n306) );
  MUX2_X1 U321 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n397), .Z(n307) );
  MUX2_X1 U322 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n396), .Z(n308) );
  MUX2_X1 U323 ( .A(n308), .B(n307), .S(N11), .Z(n309) );
  MUX2_X1 U324 ( .A(n309), .B(n306), .S(N12), .Z(n310) );
  MUX2_X1 U325 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(N10), .Z(n311) );
  MUX2_X1 U326 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(N10), .Z(n312) );
  MUX2_X1 U327 ( .A(n312), .B(n311), .S(n395), .Z(n313) );
  MUX2_X1 U328 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(N10), .Z(n314) );
  MUX2_X1 U329 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(N10), .Z(n315) );
  MUX2_X1 U330 ( .A(n315), .B(n314), .S(n395), .Z(n316) );
  MUX2_X1 U331 ( .A(n316), .B(n313), .S(N12), .Z(n317) );
  MUX2_X1 U332 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(N10), .Z(n318) );
  MUX2_X1 U333 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(N10), .Z(n319) );
  MUX2_X1 U334 ( .A(n319), .B(n318), .S(n395), .Z(n320) );
  MUX2_X1 U335 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(N10), .Z(n321) );
  MUX2_X1 U336 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(N10), .Z(n322) );
  MUX2_X1 U337 ( .A(n322), .B(n321), .S(n395), .Z(n323) );
  MUX2_X1 U338 ( .A(n323), .B(n320), .S(N12), .Z(n324) );
  MUX2_X1 U339 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n397), .Z(n325) );
  MUX2_X1 U340 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n398), .Z(n326) );
  MUX2_X1 U341 ( .A(n326), .B(n325), .S(n395), .Z(n327) );
  MUX2_X1 U342 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n398), .Z(n328) );
  MUX2_X1 U343 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n329) );
  MUX2_X1 U344 ( .A(n329), .B(n328), .S(n395), .Z(n330) );
  MUX2_X1 U345 ( .A(n330), .B(n327), .S(N12), .Z(n331) );
  MUX2_X1 U346 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n396), .Z(n332) );
  MUX2_X1 U347 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n333) );
  MUX2_X1 U348 ( .A(n333), .B(n332), .S(n395), .Z(n334) );
  MUX2_X1 U349 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n396), .Z(n335) );
  MUX2_X1 U350 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n336) );
  MUX2_X1 U351 ( .A(n336), .B(n335), .S(n395), .Z(n337) );
  MUX2_X1 U352 ( .A(n337), .B(n334), .S(N12), .Z(n338) );
  MUX2_X1 U353 ( .A(n338), .B(n331), .S(N13), .Z(N18) );
  MUX2_X1 U354 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n396), .Z(n339) );
  MUX2_X1 U355 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n396), .Z(n340) );
  MUX2_X1 U356 ( .A(n340), .B(n339), .S(n395), .Z(n341) );
  MUX2_X1 U357 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n396), .Z(n342) );
  MUX2_X1 U358 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(N10), .Z(n343) );
  MUX2_X1 U359 ( .A(n343), .B(n342), .S(n395), .Z(n344) );
  MUX2_X1 U360 ( .A(n344), .B(n341), .S(N12), .Z(n345) );
  MUX2_X1 U361 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n396), .Z(n346) );
  MUX2_X1 U362 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(N10), .Z(n347) );
  MUX2_X1 U363 ( .A(n347), .B(n346), .S(n395), .Z(n348) );
  MUX2_X1 U364 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n396), .Z(n349) );
  MUX2_X1 U365 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n350) );
  MUX2_X1 U366 ( .A(n350), .B(n349), .S(n395), .Z(n351) );
  MUX2_X1 U367 ( .A(n351), .B(n348), .S(N12), .Z(n352) );
  MUX2_X1 U368 ( .A(n352), .B(n345), .S(N13), .Z(N17) );
  MUX2_X1 U369 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n397), .Z(n353) );
  MUX2_X1 U370 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n397), .Z(n354) );
  MUX2_X1 U371 ( .A(n354), .B(n353), .S(N11), .Z(n355) );
  MUX2_X1 U372 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n397), .Z(n356) );
  MUX2_X1 U373 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n397), .Z(n357) );
  MUX2_X1 U374 ( .A(n357), .B(n356), .S(N11), .Z(n358) );
  MUX2_X1 U375 ( .A(n358), .B(n355), .S(N12), .Z(n359) );
  MUX2_X1 U376 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n397), .Z(n360) );
  MUX2_X1 U377 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n397), .Z(n361) );
  MUX2_X1 U378 ( .A(n361), .B(n360), .S(N11), .Z(n362) );
  MUX2_X1 U379 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n397), .Z(n363) );
  MUX2_X1 U380 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n397), .Z(n364) );
  MUX2_X1 U381 ( .A(n364), .B(n363), .S(n395), .Z(n365) );
  MUX2_X1 U382 ( .A(n365), .B(n362), .S(N12), .Z(n366) );
  MUX2_X1 U383 ( .A(n366), .B(n359), .S(N13), .Z(N16) );
  MUX2_X1 U384 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n397), .Z(n367) );
  MUX2_X1 U385 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n397), .Z(n368) );
  MUX2_X1 U386 ( .A(n368), .B(n367), .S(N11), .Z(n369) );
  MUX2_X1 U387 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n397), .Z(n370) );
  MUX2_X1 U388 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n397), .Z(n371) );
  MUX2_X1 U389 ( .A(n371), .B(n370), .S(N11), .Z(n372) );
  MUX2_X1 U390 ( .A(n372), .B(n369), .S(N12), .Z(n373) );
  MUX2_X1 U391 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n398), .Z(n374) );
  MUX2_X1 U392 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n398), .Z(n375) );
  MUX2_X1 U393 ( .A(n375), .B(n374), .S(N11), .Z(n376) );
  MUX2_X1 U394 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n398), .Z(n377) );
  MUX2_X1 U395 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n398), .Z(n378) );
  MUX2_X1 U396 ( .A(n378), .B(n377), .S(n395), .Z(n379) );
  MUX2_X1 U397 ( .A(n379), .B(n376), .S(N12), .Z(n380) );
  MUX2_X1 U398 ( .A(n380), .B(n373), .S(N13), .Z(N15) );
  MUX2_X1 U399 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n398), .Z(n381) );
  MUX2_X1 U400 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n398), .Z(n382) );
  MUX2_X1 U401 ( .A(n382), .B(n381), .S(N11), .Z(n383) );
  MUX2_X1 U402 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n398), .Z(n384) );
  MUX2_X1 U403 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n398), .Z(n385) );
  MUX2_X1 U404 ( .A(n385), .B(n384), .S(N11), .Z(n386) );
  MUX2_X1 U405 ( .A(n386), .B(n383), .S(N12), .Z(n387) );
  MUX2_X1 U406 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n398), .Z(n388) );
  MUX2_X1 U407 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n398), .Z(n389) );
  MUX2_X1 U408 ( .A(n389), .B(n388), .S(N11), .Z(n390) );
  MUX2_X1 U409 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n398), .Z(n391) );
  MUX2_X1 U410 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n398), .Z(n392) );
  MUX2_X1 U411 ( .A(n392), .B(n391), .S(n395), .Z(n393) );
  MUX2_X1 U412 ( .A(n393), .B(n390), .S(N12), .Z(n394) );
  MUX2_X1 U413 ( .A(n394), .B(n387), .S(N13), .Z(N14) );
  CLKBUF_X1 U414 ( .A(N10), .Z(n396) );
  INV_X1 U415 ( .A(N10), .ZN(n399) );
  INV_X1 U416 ( .A(N11), .ZN(n400) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_16 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, N19, N20, N21, n2, n4, n6, n7, n8, n9, n10, n11,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n415), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n416), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n417), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n418), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n419), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n420), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n421), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n422), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n423), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n424), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n425), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n426), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n427), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n428), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n429), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n430), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n431), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n432), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n433), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n434), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n435), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n436), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n437), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n438), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n439), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n440), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n441), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n442), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n443), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n444), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n445), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n446), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n447), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n448), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n449), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n450), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n451), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n452), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n453), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n454), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n455), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n456), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n457), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n458), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n459), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n460), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n461), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n462), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n463), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n464), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n465), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n466), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n467), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n468), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n469), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n470), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n471), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n472), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n473), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n474), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n475), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n476), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n477), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n478), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n479), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n480), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n481), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n482), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n483), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n484), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n485), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n486), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n487), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n488), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n489), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n490), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n491), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n492), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n493), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n494), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n495), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n496), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n497), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n498), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n499), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n500), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n501), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n502), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n503), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n504), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n505), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n506), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n507), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n508), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n509), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n510), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n511), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n512), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n513), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n514), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n515), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n516), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n517), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n518), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n519), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n520), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n521), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n522), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n523), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n524), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n525), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n526), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n527), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n528), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n529), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n530), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n531), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n532), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n533), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n534), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n535), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n536), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n537), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n538), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n539), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n540), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n541), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n542), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[1]  ( .D(N20), .CK(clk), .QN(n4) );
  DFF_X1 \data_out_reg[5]  ( .D(N16), .CK(clk), .QN(n2) );
  INV_X2 U3 ( .A(n2), .ZN(data_out[5]) );
  INV_X2 U4 ( .A(n4), .ZN(data_out[1]) );
  BUF_X1 U5 ( .A(N10), .Z(n401) );
  BUF_X1 U6 ( .A(N10), .Z(n402) );
  BUF_X1 U7 ( .A(N10), .Z(n403) );
  BUF_X1 U8 ( .A(N11), .Z(n400) );
  NAND2_X1 U9 ( .A1(n666), .A2(n686), .ZN(n675) );
  NAND2_X1 U10 ( .A1(n666), .A2(n676), .ZN(n665) );
  NAND2_X1 U11 ( .A1(n687), .A2(n686), .ZN(n696) );
  NAND2_X1 U12 ( .A1(n676), .A2(n687), .ZN(n685) );
  NAND2_X1 U13 ( .A1(n608), .A2(n687), .ZN(n617) );
  NAND2_X1 U14 ( .A1(n598), .A2(n687), .ZN(n607) );
  NAND2_X1 U15 ( .A1(n608), .A2(n666), .ZN(n597) );
  NAND2_X1 U16 ( .A1(n598), .A2(n666), .ZN(n588) );
  NAND2_X1 U17 ( .A1(n647), .A2(n686), .ZN(n656) );
  NAND2_X1 U18 ( .A1(n647), .A2(n676), .ZN(n646) );
  NAND2_X1 U19 ( .A1(n628), .A2(n686), .ZN(n637) );
  NAND2_X1 U20 ( .A1(n628), .A2(n676), .ZN(n626) );
  NAND2_X1 U21 ( .A1(n608), .A2(n647), .ZN(n579) );
  NAND2_X1 U22 ( .A1(n598), .A2(n647), .ZN(n570) );
  NAND2_X1 U23 ( .A1(n608), .A2(n628), .ZN(n561) );
  NAND2_X1 U24 ( .A1(n598), .A2(n628), .ZN(n551) );
  AND2_X1 U25 ( .A1(n552), .A2(N10), .ZN(n598) );
  AND2_X1 U26 ( .A1(n552), .A2(n404), .ZN(n608) );
  AND2_X1 U27 ( .A1(N10), .A2(n627), .ZN(n676) );
  AND2_X1 U28 ( .A1(n627), .A2(n404), .ZN(n686) );
  OAI21_X1 U29 ( .B1(n696), .B2(n414), .A(n695), .ZN(n542) );
  NAND2_X1 U30 ( .A1(\mem[0][0] ), .A2(n696), .ZN(n695) );
  OAI21_X1 U31 ( .B1(n696), .B2(n413), .A(n694), .ZN(n541) );
  NAND2_X1 U32 ( .A1(\mem[0][1] ), .A2(n696), .ZN(n694) );
  OAI21_X1 U33 ( .B1(n696), .B2(n412), .A(n693), .ZN(n540) );
  NAND2_X1 U34 ( .A1(\mem[0][2] ), .A2(n696), .ZN(n693) );
  OAI21_X1 U35 ( .B1(n696), .B2(n411), .A(n692), .ZN(n539) );
  NAND2_X1 U36 ( .A1(\mem[0][3] ), .A2(n696), .ZN(n692) );
  OAI21_X1 U37 ( .B1(n696), .B2(n410), .A(n691), .ZN(n538) );
  NAND2_X1 U38 ( .A1(\mem[0][4] ), .A2(n696), .ZN(n691) );
  OAI21_X1 U39 ( .B1(n696), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U40 ( .A1(\mem[0][5] ), .A2(n696), .ZN(n690) );
  OAI21_X1 U41 ( .B1(n696), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U42 ( .A1(\mem[0][6] ), .A2(n696), .ZN(n689) );
  OAI21_X1 U43 ( .B1(n696), .B2(n407), .A(n688), .ZN(n535) );
  NAND2_X1 U44 ( .A1(\mem[0][7] ), .A2(n696), .ZN(n688) );
  OAI21_X1 U45 ( .B1(n414), .B2(n675), .A(n674), .ZN(n526) );
  NAND2_X1 U46 ( .A1(\mem[2][0] ), .A2(n675), .ZN(n674) );
  OAI21_X1 U47 ( .B1(n413), .B2(n675), .A(n673), .ZN(n525) );
  NAND2_X1 U48 ( .A1(\mem[2][1] ), .A2(n675), .ZN(n673) );
  OAI21_X1 U49 ( .B1(n412), .B2(n675), .A(n672), .ZN(n524) );
  NAND2_X1 U50 ( .A1(\mem[2][2] ), .A2(n675), .ZN(n672) );
  OAI21_X1 U51 ( .B1(n411), .B2(n675), .A(n671), .ZN(n523) );
  NAND2_X1 U52 ( .A1(\mem[2][3] ), .A2(n675), .ZN(n671) );
  OAI21_X1 U53 ( .B1(n410), .B2(n675), .A(n670), .ZN(n522) );
  NAND2_X1 U54 ( .A1(\mem[2][4] ), .A2(n675), .ZN(n670) );
  OAI21_X1 U55 ( .B1(n409), .B2(n675), .A(n669), .ZN(n521) );
  NAND2_X1 U56 ( .A1(\mem[2][5] ), .A2(n675), .ZN(n669) );
  OAI21_X1 U57 ( .B1(n408), .B2(n675), .A(n668), .ZN(n520) );
  NAND2_X1 U58 ( .A1(\mem[2][6] ), .A2(n675), .ZN(n668) );
  OAI21_X1 U59 ( .B1(n407), .B2(n675), .A(n667), .ZN(n519) );
  NAND2_X1 U60 ( .A1(\mem[2][7] ), .A2(n675), .ZN(n667) );
  OAI21_X1 U61 ( .B1(n414), .B2(n665), .A(n664), .ZN(n518) );
  NAND2_X1 U62 ( .A1(\mem[3][0] ), .A2(n665), .ZN(n664) );
  OAI21_X1 U63 ( .B1(n413), .B2(n665), .A(n663), .ZN(n517) );
  NAND2_X1 U64 ( .A1(\mem[3][1] ), .A2(n665), .ZN(n663) );
  OAI21_X1 U65 ( .B1(n412), .B2(n665), .A(n662), .ZN(n516) );
  NAND2_X1 U66 ( .A1(\mem[3][2] ), .A2(n665), .ZN(n662) );
  OAI21_X1 U67 ( .B1(n411), .B2(n665), .A(n661), .ZN(n515) );
  NAND2_X1 U68 ( .A1(\mem[3][3] ), .A2(n665), .ZN(n661) );
  OAI21_X1 U69 ( .B1(n410), .B2(n665), .A(n660), .ZN(n514) );
  NAND2_X1 U70 ( .A1(\mem[3][4] ), .A2(n665), .ZN(n660) );
  OAI21_X1 U71 ( .B1(n409), .B2(n665), .A(n659), .ZN(n513) );
  NAND2_X1 U72 ( .A1(\mem[3][5] ), .A2(n665), .ZN(n659) );
  OAI21_X1 U73 ( .B1(n408), .B2(n665), .A(n658), .ZN(n512) );
  NAND2_X1 U74 ( .A1(\mem[3][6] ), .A2(n665), .ZN(n658) );
  OAI21_X1 U75 ( .B1(n407), .B2(n665), .A(n657), .ZN(n511) );
  NAND2_X1 U76 ( .A1(\mem[3][7] ), .A2(n665), .ZN(n657) );
  NOR2_X1 U77 ( .A1(n406), .A2(N13), .ZN(n627) );
  INV_X1 U78 ( .A(wr_en), .ZN(n406) );
  OAI21_X1 U79 ( .B1(n414), .B2(n685), .A(n684), .ZN(n534) );
  NAND2_X1 U80 ( .A1(\mem[1][0] ), .A2(n685), .ZN(n684) );
  OAI21_X1 U81 ( .B1(n413), .B2(n685), .A(n683), .ZN(n533) );
  NAND2_X1 U82 ( .A1(\mem[1][1] ), .A2(n685), .ZN(n683) );
  OAI21_X1 U83 ( .B1(n412), .B2(n685), .A(n682), .ZN(n532) );
  NAND2_X1 U84 ( .A1(\mem[1][2] ), .A2(n685), .ZN(n682) );
  OAI21_X1 U85 ( .B1(n411), .B2(n685), .A(n681), .ZN(n531) );
  NAND2_X1 U86 ( .A1(\mem[1][3] ), .A2(n685), .ZN(n681) );
  OAI21_X1 U87 ( .B1(n410), .B2(n685), .A(n680), .ZN(n530) );
  NAND2_X1 U88 ( .A1(\mem[1][4] ), .A2(n685), .ZN(n680) );
  OAI21_X1 U89 ( .B1(n409), .B2(n685), .A(n679), .ZN(n529) );
  NAND2_X1 U90 ( .A1(\mem[1][5] ), .A2(n685), .ZN(n679) );
  OAI21_X1 U91 ( .B1(n408), .B2(n685), .A(n678), .ZN(n528) );
  NAND2_X1 U92 ( .A1(\mem[1][6] ), .A2(n685), .ZN(n678) );
  OAI21_X1 U93 ( .B1(n407), .B2(n685), .A(n677), .ZN(n527) );
  NAND2_X1 U94 ( .A1(\mem[1][7] ), .A2(n685), .ZN(n677) );
  OAI21_X1 U95 ( .B1(n414), .B2(n656), .A(n655), .ZN(n510) );
  NAND2_X1 U96 ( .A1(\mem[4][0] ), .A2(n656), .ZN(n655) );
  OAI21_X1 U97 ( .B1(n413), .B2(n656), .A(n654), .ZN(n509) );
  NAND2_X1 U98 ( .A1(\mem[4][1] ), .A2(n656), .ZN(n654) );
  OAI21_X1 U99 ( .B1(n412), .B2(n656), .A(n653), .ZN(n508) );
  NAND2_X1 U100 ( .A1(\mem[4][2] ), .A2(n656), .ZN(n653) );
  OAI21_X1 U101 ( .B1(n411), .B2(n656), .A(n652), .ZN(n507) );
  NAND2_X1 U102 ( .A1(\mem[4][3] ), .A2(n656), .ZN(n652) );
  OAI21_X1 U103 ( .B1(n410), .B2(n656), .A(n651), .ZN(n506) );
  NAND2_X1 U104 ( .A1(\mem[4][4] ), .A2(n656), .ZN(n651) );
  OAI21_X1 U105 ( .B1(n409), .B2(n656), .A(n650), .ZN(n505) );
  NAND2_X1 U106 ( .A1(\mem[4][5] ), .A2(n656), .ZN(n650) );
  OAI21_X1 U107 ( .B1(n408), .B2(n656), .A(n649), .ZN(n504) );
  NAND2_X1 U108 ( .A1(\mem[4][6] ), .A2(n656), .ZN(n649) );
  OAI21_X1 U109 ( .B1(n407), .B2(n656), .A(n648), .ZN(n503) );
  NAND2_X1 U110 ( .A1(\mem[4][7] ), .A2(n656), .ZN(n648) );
  OAI21_X1 U111 ( .B1(n414), .B2(n646), .A(n645), .ZN(n502) );
  NAND2_X1 U112 ( .A1(\mem[5][0] ), .A2(n646), .ZN(n645) );
  OAI21_X1 U113 ( .B1(n413), .B2(n646), .A(n644), .ZN(n501) );
  NAND2_X1 U114 ( .A1(\mem[5][1] ), .A2(n646), .ZN(n644) );
  OAI21_X1 U115 ( .B1(n412), .B2(n646), .A(n643), .ZN(n500) );
  NAND2_X1 U116 ( .A1(\mem[5][2] ), .A2(n646), .ZN(n643) );
  OAI21_X1 U117 ( .B1(n411), .B2(n646), .A(n642), .ZN(n499) );
  NAND2_X1 U118 ( .A1(\mem[5][3] ), .A2(n646), .ZN(n642) );
  OAI21_X1 U119 ( .B1(n410), .B2(n646), .A(n641), .ZN(n498) );
  NAND2_X1 U120 ( .A1(\mem[5][4] ), .A2(n646), .ZN(n641) );
  OAI21_X1 U121 ( .B1(n409), .B2(n646), .A(n640), .ZN(n497) );
  NAND2_X1 U122 ( .A1(\mem[5][5] ), .A2(n646), .ZN(n640) );
  OAI21_X1 U123 ( .B1(n408), .B2(n646), .A(n639), .ZN(n496) );
  NAND2_X1 U124 ( .A1(\mem[5][6] ), .A2(n646), .ZN(n639) );
  OAI21_X1 U125 ( .B1(n407), .B2(n646), .A(n638), .ZN(n495) );
  NAND2_X1 U126 ( .A1(\mem[5][7] ), .A2(n646), .ZN(n638) );
  OAI21_X1 U127 ( .B1(n414), .B2(n637), .A(n636), .ZN(n494) );
  NAND2_X1 U128 ( .A1(\mem[6][0] ), .A2(n637), .ZN(n636) );
  OAI21_X1 U129 ( .B1(n413), .B2(n637), .A(n635), .ZN(n493) );
  NAND2_X1 U130 ( .A1(\mem[6][1] ), .A2(n637), .ZN(n635) );
  OAI21_X1 U131 ( .B1(n412), .B2(n637), .A(n634), .ZN(n492) );
  NAND2_X1 U132 ( .A1(\mem[6][2] ), .A2(n637), .ZN(n634) );
  OAI21_X1 U133 ( .B1(n411), .B2(n637), .A(n633), .ZN(n491) );
  NAND2_X1 U134 ( .A1(\mem[6][3] ), .A2(n637), .ZN(n633) );
  OAI21_X1 U135 ( .B1(n410), .B2(n637), .A(n632), .ZN(n490) );
  NAND2_X1 U136 ( .A1(\mem[6][4] ), .A2(n637), .ZN(n632) );
  OAI21_X1 U137 ( .B1(n409), .B2(n637), .A(n631), .ZN(n489) );
  NAND2_X1 U138 ( .A1(\mem[6][5] ), .A2(n637), .ZN(n631) );
  OAI21_X1 U139 ( .B1(n408), .B2(n637), .A(n630), .ZN(n488) );
  NAND2_X1 U140 ( .A1(\mem[6][6] ), .A2(n637), .ZN(n630) );
  OAI21_X1 U141 ( .B1(n407), .B2(n637), .A(n629), .ZN(n487) );
  NAND2_X1 U142 ( .A1(\mem[6][7] ), .A2(n637), .ZN(n629) );
  OAI21_X1 U143 ( .B1(n414), .B2(n626), .A(n625), .ZN(n486) );
  NAND2_X1 U144 ( .A1(\mem[7][0] ), .A2(n626), .ZN(n625) );
  OAI21_X1 U145 ( .B1(n413), .B2(n626), .A(n624), .ZN(n485) );
  NAND2_X1 U146 ( .A1(\mem[7][1] ), .A2(n626), .ZN(n624) );
  OAI21_X1 U147 ( .B1(n412), .B2(n626), .A(n623), .ZN(n484) );
  NAND2_X1 U148 ( .A1(\mem[7][2] ), .A2(n626), .ZN(n623) );
  OAI21_X1 U149 ( .B1(n411), .B2(n626), .A(n622), .ZN(n483) );
  NAND2_X1 U150 ( .A1(\mem[7][3] ), .A2(n626), .ZN(n622) );
  OAI21_X1 U151 ( .B1(n410), .B2(n626), .A(n621), .ZN(n482) );
  NAND2_X1 U152 ( .A1(\mem[7][4] ), .A2(n626), .ZN(n621) );
  OAI21_X1 U153 ( .B1(n409), .B2(n626), .A(n620), .ZN(n481) );
  NAND2_X1 U154 ( .A1(\mem[7][5] ), .A2(n626), .ZN(n620) );
  OAI21_X1 U155 ( .B1(n408), .B2(n626), .A(n619), .ZN(n480) );
  NAND2_X1 U156 ( .A1(\mem[7][6] ), .A2(n626), .ZN(n619) );
  OAI21_X1 U157 ( .B1(n407), .B2(n626), .A(n618), .ZN(n479) );
  NAND2_X1 U158 ( .A1(\mem[7][7] ), .A2(n626), .ZN(n618) );
  OAI21_X1 U159 ( .B1(n414), .B2(n617), .A(n616), .ZN(n478) );
  NAND2_X1 U160 ( .A1(\mem[8][0] ), .A2(n617), .ZN(n616) );
  OAI21_X1 U161 ( .B1(n413), .B2(n617), .A(n615), .ZN(n477) );
  NAND2_X1 U162 ( .A1(\mem[8][1] ), .A2(n617), .ZN(n615) );
  OAI21_X1 U163 ( .B1(n412), .B2(n617), .A(n614), .ZN(n476) );
  NAND2_X1 U164 ( .A1(\mem[8][2] ), .A2(n617), .ZN(n614) );
  OAI21_X1 U165 ( .B1(n411), .B2(n617), .A(n613), .ZN(n475) );
  NAND2_X1 U166 ( .A1(\mem[8][3] ), .A2(n617), .ZN(n613) );
  OAI21_X1 U167 ( .B1(n410), .B2(n617), .A(n612), .ZN(n474) );
  NAND2_X1 U168 ( .A1(\mem[8][4] ), .A2(n617), .ZN(n612) );
  OAI21_X1 U169 ( .B1(n409), .B2(n617), .A(n611), .ZN(n473) );
  NAND2_X1 U170 ( .A1(\mem[8][5] ), .A2(n617), .ZN(n611) );
  OAI21_X1 U171 ( .B1(n408), .B2(n617), .A(n610), .ZN(n472) );
  NAND2_X1 U172 ( .A1(\mem[8][6] ), .A2(n617), .ZN(n610) );
  OAI21_X1 U173 ( .B1(n407), .B2(n617), .A(n609), .ZN(n471) );
  NAND2_X1 U174 ( .A1(\mem[8][7] ), .A2(n617), .ZN(n609) );
  OAI21_X1 U175 ( .B1(n414), .B2(n607), .A(n606), .ZN(n470) );
  NAND2_X1 U176 ( .A1(\mem[9][0] ), .A2(n607), .ZN(n606) );
  OAI21_X1 U177 ( .B1(n413), .B2(n607), .A(n605), .ZN(n469) );
  NAND2_X1 U178 ( .A1(\mem[9][1] ), .A2(n607), .ZN(n605) );
  OAI21_X1 U179 ( .B1(n412), .B2(n607), .A(n604), .ZN(n468) );
  NAND2_X1 U180 ( .A1(\mem[9][2] ), .A2(n607), .ZN(n604) );
  OAI21_X1 U181 ( .B1(n411), .B2(n607), .A(n603), .ZN(n467) );
  NAND2_X1 U182 ( .A1(\mem[9][3] ), .A2(n607), .ZN(n603) );
  OAI21_X1 U183 ( .B1(n410), .B2(n607), .A(n602), .ZN(n466) );
  NAND2_X1 U184 ( .A1(\mem[9][4] ), .A2(n607), .ZN(n602) );
  OAI21_X1 U185 ( .B1(n409), .B2(n607), .A(n601), .ZN(n465) );
  NAND2_X1 U186 ( .A1(\mem[9][5] ), .A2(n607), .ZN(n601) );
  OAI21_X1 U187 ( .B1(n408), .B2(n607), .A(n600), .ZN(n464) );
  NAND2_X1 U188 ( .A1(\mem[9][6] ), .A2(n607), .ZN(n600) );
  OAI21_X1 U189 ( .B1(n407), .B2(n607), .A(n599), .ZN(n463) );
  NAND2_X1 U190 ( .A1(\mem[9][7] ), .A2(n607), .ZN(n599) );
  OAI21_X1 U191 ( .B1(n414), .B2(n597), .A(n596), .ZN(n462) );
  NAND2_X1 U192 ( .A1(\mem[10][0] ), .A2(n597), .ZN(n596) );
  OAI21_X1 U193 ( .B1(n413), .B2(n597), .A(n595), .ZN(n461) );
  NAND2_X1 U194 ( .A1(\mem[10][1] ), .A2(n597), .ZN(n595) );
  OAI21_X1 U195 ( .B1(n412), .B2(n597), .A(n594), .ZN(n460) );
  NAND2_X1 U196 ( .A1(\mem[10][2] ), .A2(n597), .ZN(n594) );
  OAI21_X1 U197 ( .B1(n411), .B2(n597), .A(n593), .ZN(n459) );
  NAND2_X1 U198 ( .A1(\mem[10][3] ), .A2(n597), .ZN(n593) );
  OAI21_X1 U199 ( .B1(n410), .B2(n597), .A(n592), .ZN(n458) );
  NAND2_X1 U200 ( .A1(\mem[10][4] ), .A2(n597), .ZN(n592) );
  OAI21_X1 U201 ( .B1(n409), .B2(n597), .A(n591), .ZN(n457) );
  NAND2_X1 U202 ( .A1(\mem[10][5] ), .A2(n597), .ZN(n591) );
  OAI21_X1 U203 ( .B1(n408), .B2(n597), .A(n590), .ZN(n456) );
  NAND2_X1 U204 ( .A1(\mem[10][6] ), .A2(n597), .ZN(n590) );
  OAI21_X1 U205 ( .B1(n407), .B2(n597), .A(n589), .ZN(n455) );
  NAND2_X1 U206 ( .A1(\mem[10][7] ), .A2(n597), .ZN(n589) );
  OAI21_X1 U207 ( .B1(n414), .B2(n588), .A(n587), .ZN(n454) );
  NAND2_X1 U208 ( .A1(\mem[11][0] ), .A2(n588), .ZN(n587) );
  OAI21_X1 U209 ( .B1(n413), .B2(n588), .A(n586), .ZN(n453) );
  NAND2_X1 U210 ( .A1(\mem[11][1] ), .A2(n588), .ZN(n586) );
  OAI21_X1 U211 ( .B1(n412), .B2(n588), .A(n585), .ZN(n452) );
  NAND2_X1 U212 ( .A1(\mem[11][2] ), .A2(n588), .ZN(n585) );
  OAI21_X1 U213 ( .B1(n411), .B2(n588), .A(n584), .ZN(n451) );
  NAND2_X1 U214 ( .A1(\mem[11][3] ), .A2(n588), .ZN(n584) );
  OAI21_X1 U215 ( .B1(n410), .B2(n588), .A(n583), .ZN(n450) );
  NAND2_X1 U216 ( .A1(\mem[11][4] ), .A2(n588), .ZN(n583) );
  OAI21_X1 U217 ( .B1(n409), .B2(n588), .A(n582), .ZN(n449) );
  NAND2_X1 U218 ( .A1(\mem[11][5] ), .A2(n588), .ZN(n582) );
  OAI21_X1 U219 ( .B1(n408), .B2(n588), .A(n581), .ZN(n448) );
  NAND2_X1 U220 ( .A1(\mem[11][6] ), .A2(n588), .ZN(n581) );
  OAI21_X1 U221 ( .B1(n407), .B2(n588), .A(n580), .ZN(n447) );
  NAND2_X1 U222 ( .A1(\mem[11][7] ), .A2(n588), .ZN(n580) );
  OAI21_X1 U223 ( .B1(n414), .B2(n579), .A(n578), .ZN(n446) );
  NAND2_X1 U224 ( .A1(\mem[12][0] ), .A2(n579), .ZN(n578) );
  OAI21_X1 U225 ( .B1(n413), .B2(n579), .A(n577), .ZN(n445) );
  NAND2_X1 U226 ( .A1(\mem[12][1] ), .A2(n579), .ZN(n577) );
  OAI21_X1 U227 ( .B1(n412), .B2(n579), .A(n576), .ZN(n444) );
  NAND2_X1 U228 ( .A1(\mem[12][2] ), .A2(n579), .ZN(n576) );
  OAI21_X1 U229 ( .B1(n411), .B2(n579), .A(n575), .ZN(n443) );
  NAND2_X1 U230 ( .A1(\mem[12][3] ), .A2(n579), .ZN(n575) );
  OAI21_X1 U231 ( .B1(n410), .B2(n579), .A(n574), .ZN(n442) );
  NAND2_X1 U232 ( .A1(\mem[12][4] ), .A2(n579), .ZN(n574) );
  OAI21_X1 U233 ( .B1(n409), .B2(n579), .A(n573), .ZN(n441) );
  NAND2_X1 U234 ( .A1(\mem[12][5] ), .A2(n579), .ZN(n573) );
  OAI21_X1 U235 ( .B1(n408), .B2(n579), .A(n572), .ZN(n440) );
  NAND2_X1 U236 ( .A1(\mem[12][6] ), .A2(n579), .ZN(n572) );
  OAI21_X1 U237 ( .B1(n407), .B2(n579), .A(n571), .ZN(n439) );
  NAND2_X1 U238 ( .A1(\mem[12][7] ), .A2(n579), .ZN(n571) );
  OAI21_X1 U239 ( .B1(n414), .B2(n570), .A(n569), .ZN(n438) );
  NAND2_X1 U240 ( .A1(\mem[13][0] ), .A2(n570), .ZN(n569) );
  OAI21_X1 U241 ( .B1(n413), .B2(n570), .A(n568), .ZN(n437) );
  NAND2_X1 U242 ( .A1(\mem[13][1] ), .A2(n570), .ZN(n568) );
  OAI21_X1 U243 ( .B1(n412), .B2(n570), .A(n567), .ZN(n436) );
  NAND2_X1 U244 ( .A1(\mem[13][2] ), .A2(n570), .ZN(n567) );
  OAI21_X1 U245 ( .B1(n411), .B2(n570), .A(n566), .ZN(n435) );
  NAND2_X1 U246 ( .A1(\mem[13][3] ), .A2(n570), .ZN(n566) );
  OAI21_X1 U247 ( .B1(n410), .B2(n570), .A(n565), .ZN(n434) );
  NAND2_X1 U248 ( .A1(\mem[13][4] ), .A2(n570), .ZN(n565) );
  OAI21_X1 U249 ( .B1(n409), .B2(n570), .A(n564), .ZN(n433) );
  NAND2_X1 U250 ( .A1(\mem[13][5] ), .A2(n570), .ZN(n564) );
  OAI21_X1 U251 ( .B1(n408), .B2(n570), .A(n563), .ZN(n432) );
  NAND2_X1 U252 ( .A1(\mem[13][6] ), .A2(n570), .ZN(n563) );
  OAI21_X1 U253 ( .B1(n407), .B2(n570), .A(n562), .ZN(n431) );
  NAND2_X1 U254 ( .A1(\mem[13][7] ), .A2(n570), .ZN(n562) );
  OAI21_X1 U255 ( .B1(n414), .B2(n561), .A(n560), .ZN(n430) );
  NAND2_X1 U256 ( .A1(\mem[14][0] ), .A2(n561), .ZN(n560) );
  OAI21_X1 U257 ( .B1(n413), .B2(n561), .A(n559), .ZN(n429) );
  NAND2_X1 U258 ( .A1(\mem[14][1] ), .A2(n561), .ZN(n559) );
  OAI21_X1 U259 ( .B1(n412), .B2(n561), .A(n558), .ZN(n428) );
  NAND2_X1 U260 ( .A1(\mem[14][2] ), .A2(n561), .ZN(n558) );
  OAI21_X1 U261 ( .B1(n411), .B2(n561), .A(n557), .ZN(n427) );
  NAND2_X1 U262 ( .A1(\mem[14][3] ), .A2(n561), .ZN(n557) );
  OAI21_X1 U263 ( .B1(n410), .B2(n561), .A(n556), .ZN(n426) );
  NAND2_X1 U264 ( .A1(\mem[14][4] ), .A2(n561), .ZN(n556) );
  OAI21_X1 U265 ( .B1(n409), .B2(n561), .A(n555), .ZN(n425) );
  NAND2_X1 U266 ( .A1(\mem[14][5] ), .A2(n561), .ZN(n555) );
  OAI21_X1 U267 ( .B1(n408), .B2(n561), .A(n554), .ZN(n424) );
  NAND2_X1 U268 ( .A1(\mem[14][6] ), .A2(n561), .ZN(n554) );
  OAI21_X1 U269 ( .B1(n407), .B2(n561), .A(n553), .ZN(n423) );
  NAND2_X1 U270 ( .A1(\mem[14][7] ), .A2(n561), .ZN(n553) );
  OAI21_X1 U271 ( .B1(n414), .B2(n551), .A(n550), .ZN(n422) );
  NAND2_X1 U272 ( .A1(\mem[15][0] ), .A2(n551), .ZN(n550) );
  OAI21_X1 U273 ( .B1(n413), .B2(n551), .A(n549), .ZN(n421) );
  NAND2_X1 U274 ( .A1(\mem[15][1] ), .A2(n551), .ZN(n549) );
  OAI21_X1 U275 ( .B1(n412), .B2(n551), .A(n548), .ZN(n420) );
  NAND2_X1 U276 ( .A1(\mem[15][2] ), .A2(n551), .ZN(n548) );
  OAI21_X1 U277 ( .B1(n411), .B2(n551), .A(n547), .ZN(n419) );
  NAND2_X1 U278 ( .A1(\mem[15][3] ), .A2(n551), .ZN(n547) );
  OAI21_X1 U279 ( .B1(n410), .B2(n551), .A(n546), .ZN(n418) );
  NAND2_X1 U280 ( .A1(\mem[15][4] ), .A2(n551), .ZN(n546) );
  OAI21_X1 U281 ( .B1(n409), .B2(n551), .A(n545), .ZN(n417) );
  NAND2_X1 U282 ( .A1(\mem[15][5] ), .A2(n551), .ZN(n545) );
  OAI21_X1 U283 ( .B1(n408), .B2(n551), .A(n544), .ZN(n416) );
  NAND2_X1 U284 ( .A1(\mem[15][6] ), .A2(n551), .ZN(n544) );
  OAI21_X1 U285 ( .B1(n407), .B2(n551), .A(n543), .ZN(n415) );
  NAND2_X1 U286 ( .A1(\mem[15][7] ), .A2(n551), .ZN(n543) );
  AND2_X1 U287 ( .A1(N13), .A2(wr_en), .ZN(n552) );
  NOR2_X1 U288 ( .A1(N11), .A2(N12), .ZN(n687) );
  NOR2_X1 U289 ( .A1(n405), .A2(N12), .ZN(n666) );
  AND2_X1 U290 ( .A1(N12), .A2(n405), .ZN(n647) );
  AND2_X1 U291 ( .A1(N12), .A2(N11), .ZN(n628) );
  INV_X1 U292 ( .A(data_in[0]), .ZN(n414) );
  INV_X1 U293 ( .A(data_in[1]), .ZN(n413) );
  INV_X1 U294 ( .A(data_in[2]), .ZN(n412) );
  INV_X1 U295 ( .A(data_in[3]), .ZN(n411) );
  INV_X1 U296 ( .A(data_in[4]), .ZN(n410) );
  INV_X1 U297 ( .A(data_in[5]), .ZN(n409) );
  INV_X1 U298 ( .A(data_in[6]), .ZN(n408) );
  INV_X1 U299 ( .A(data_in[7]), .ZN(n407) );
  MUX2_X1 U300 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(N10), .Z(n6) );
  MUX2_X1 U301 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(N10), .Z(n7) );
  MUX2_X1 U302 ( .A(n7), .B(n6), .S(N11), .Z(n8) );
  MUX2_X1 U303 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(N10), .Z(n9) );
  MUX2_X1 U304 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n10) );
  MUX2_X1 U305 ( .A(n10), .B(n9), .S(N11), .Z(n11) );
  MUX2_X1 U306 ( .A(n11), .B(n8), .S(N12), .Z(n294) );
  MUX2_X1 U307 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n401), .Z(n295) );
  MUX2_X1 U308 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n401), .Z(n296) );
  MUX2_X1 U309 ( .A(n296), .B(n295), .S(N11), .Z(n297) );
  MUX2_X1 U310 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n401), .Z(n298) );
  MUX2_X1 U311 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n401), .Z(n299) );
  MUX2_X1 U312 ( .A(n299), .B(n298), .S(n400), .Z(n300) );
  MUX2_X1 U313 ( .A(n300), .B(n297), .S(N12), .Z(n301) );
  MUX2_X1 U314 ( .A(n301), .B(n294), .S(N13), .Z(N21) );
  MUX2_X1 U315 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n401), .Z(n302) );
  MUX2_X1 U316 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n401), .Z(n303) );
  MUX2_X1 U317 ( .A(n303), .B(n302), .S(N11), .Z(n304) );
  MUX2_X1 U318 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n401), .Z(n305) );
  MUX2_X1 U319 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n401), .Z(n306) );
  MUX2_X1 U320 ( .A(n306), .B(n305), .S(N11), .Z(n307) );
  MUX2_X1 U321 ( .A(n307), .B(n304), .S(N12), .Z(n308) );
  MUX2_X1 U322 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n401), .Z(n309) );
  MUX2_X1 U323 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n401), .Z(n310) );
  MUX2_X1 U324 ( .A(n310), .B(n309), .S(N11), .Z(n311) );
  MUX2_X1 U325 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n401), .Z(n312) );
  MUX2_X1 U326 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n401), .Z(n313) );
  MUX2_X1 U327 ( .A(n313), .B(n312), .S(n400), .Z(n314) );
  MUX2_X1 U328 ( .A(n314), .B(n311), .S(N12), .Z(n315) );
  MUX2_X1 U329 ( .A(n315), .B(n308), .S(N13), .Z(N20) );
  MUX2_X1 U330 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n402), .Z(n316) );
  MUX2_X1 U331 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n402), .Z(n317) );
  MUX2_X1 U332 ( .A(n317), .B(n316), .S(N11), .Z(n318) );
  MUX2_X1 U333 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n402), .Z(n319) );
  MUX2_X1 U334 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n402), .Z(n320) );
  MUX2_X1 U335 ( .A(n320), .B(n319), .S(N11), .Z(n321) );
  MUX2_X1 U336 ( .A(n321), .B(n318), .S(N12), .Z(n322) );
  MUX2_X1 U337 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n402), .Z(n323) );
  MUX2_X1 U338 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n402), .Z(n324) );
  MUX2_X1 U339 ( .A(n324), .B(n323), .S(N11), .Z(n325) );
  MUX2_X1 U340 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n402), .Z(n326) );
  MUX2_X1 U341 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n402), .Z(n327) );
  MUX2_X1 U342 ( .A(n327), .B(n326), .S(N11), .Z(n328) );
  MUX2_X1 U343 ( .A(n328), .B(n325), .S(N12), .Z(n329) );
  MUX2_X1 U344 ( .A(n329), .B(n322), .S(N13), .Z(N19) );
  MUX2_X1 U345 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n402), .Z(n330) );
  MUX2_X1 U346 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n402), .Z(n331) );
  MUX2_X1 U347 ( .A(n331), .B(n330), .S(N11), .Z(n332) );
  MUX2_X1 U348 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n402), .Z(n333) );
  MUX2_X1 U349 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n402), .Z(n334) );
  MUX2_X1 U350 ( .A(n334), .B(n333), .S(N11), .Z(n335) );
  MUX2_X1 U351 ( .A(n335), .B(n332), .S(N12), .Z(n336) );
  MUX2_X1 U352 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n403), .Z(n337) );
  MUX2_X1 U353 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n403), .Z(n338) );
  MUX2_X1 U354 ( .A(n338), .B(n337), .S(N11), .Z(n339) );
  MUX2_X1 U355 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n403), .Z(n340) );
  MUX2_X1 U356 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n403), .Z(n341) );
  MUX2_X1 U357 ( .A(n341), .B(n340), .S(N11), .Z(n342) );
  MUX2_X1 U358 ( .A(n342), .B(n339), .S(N12), .Z(n343) );
  MUX2_X1 U359 ( .A(n343), .B(n336), .S(N13), .Z(N18) );
  MUX2_X1 U360 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n403), .Z(n344) );
  MUX2_X1 U361 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n403), .Z(n345) );
  MUX2_X1 U362 ( .A(n345), .B(n344), .S(N11), .Z(n346) );
  MUX2_X1 U363 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n403), .Z(n347) );
  MUX2_X1 U364 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n403), .Z(n348) );
  MUX2_X1 U365 ( .A(n348), .B(n347), .S(N11), .Z(n349) );
  MUX2_X1 U366 ( .A(n349), .B(n346), .S(N12), .Z(n350) );
  MUX2_X1 U367 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n403), .Z(n351) );
  MUX2_X1 U368 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n403), .Z(n352) );
  MUX2_X1 U369 ( .A(n352), .B(n351), .S(N11), .Z(n353) );
  MUX2_X1 U370 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n403), .Z(n354) );
  MUX2_X1 U371 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n403), .Z(n355) );
  MUX2_X1 U372 ( .A(n355), .B(n354), .S(N11), .Z(n356) );
  MUX2_X1 U373 ( .A(n356), .B(n353), .S(N12), .Z(n357) );
  MUX2_X1 U374 ( .A(n357), .B(n350), .S(N13), .Z(N17) );
  MUX2_X1 U375 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(N10), .Z(n358) );
  MUX2_X1 U376 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n402), .Z(n359) );
  MUX2_X1 U377 ( .A(n359), .B(n358), .S(n400), .Z(n360) );
  MUX2_X1 U378 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n403), .Z(n361) );
  MUX2_X1 U379 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n403), .Z(n362) );
  MUX2_X1 U380 ( .A(n362), .B(n361), .S(n400), .Z(n363) );
  MUX2_X1 U381 ( .A(n363), .B(n360), .S(N12), .Z(n364) );
  MUX2_X1 U382 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n402), .Z(n365) );
  MUX2_X1 U383 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n402), .Z(n366) );
  MUX2_X1 U384 ( .A(n366), .B(n365), .S(n400), .Z(n367) );
  MUX2_X1 U385 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n401), .Z(n368) );
  MUX2_X1 U386 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n402), .Z(n369) );
  MUX2_X1 U387 ( .A(n369), .B(n368), .S(n400), .Z(n370) );
  MUX2_X1 U388 ( .A(n370), .B(n367), .S(N12), .Z(n371) );
  MUX2_X1 U389 ( .A(n371), .B(n364), .S(N13), .Z(N16) );
  MUX2_X1 U390 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n401), .Z(n372) );
  MUX2_X1 U391 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n403), .Z(n373) );
  MUX2_X1 U392 ( .A(n373), .B(n372), .S(n400), .Z(n374) );
  MUX2_X1 U393 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n401), .Z(n375) );
  MUX2_X1 U394 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n401), .Z(n376) );
  MUX2_X1 U395 ( .A(n376), .B(n375), .S(n400), .Z(n377) );
  MUX2_X1 U396 ( .A(n377), .B(n374), .S(N12), .Z(n378) );
  MUX2_X1 U397 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n379) );
  MUX2_X1 U398 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n380) );
  MUX2_X1 U399 ( .A(n380), .B(n379), .S(n400), .Z(n381) );
  MUX2_X1 U400 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n382) );
  MUX2_X1 U401 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n383) );
  MUX2_X1 U402 ( .A(n383), .B(n382), .S(n400), .Z(n384) );
  MUX2_X1 U403 ( .A(n384), .B(n381), .S(N12), .Z(n385) );
  MUX2_X1 U404 ( .A(n385), .B(n378), .S(N13), .Z(N15) );
  MUX2_X1 U405 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(N10), .Z(n386) );
  MUX2_X1 U406 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n387) );
  MUX2_X1 U407 ( .A(n387), .B(n386), .S(n400), .Z(n388) );
  MUX2_X1 U408 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(N10), .Z(n389) );
  MUX2_X1 U409 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n390) );
  MUX2_X1 U410 ( .A(n390), .B(n389), .S(n400), .Z(n391) );
  MUX2_X1 U411 ( .A(n391), .B(n388), .S(N12), .Z(n392) );
  MUX2_X1 U412 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n393) );
  MUX2_X1 U413 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n394) );
  MUX2_X1 U414 ( .A(n394), .B(n393), .S(n400), .Z(n395) );
  MUX2_X1 U415 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n396) );
  MUX2_X1 U416 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n403), .Z(n397) );
  MUX2_X1 U417 ( .A(n397), .B(n396), .S(n400), .Z(n398) );
  MUX2_X1 U418 ( .A(n398), .B(n395), .S(N12), .Z(n399) );
  MUX2_X1 U419 ( .A(n399), .B(n392), .S(N13), .Z(N14) );
  INV_X1 U420 ( .A(N10), .ZN(n404) );
  INV_X1 U421 ( .A(N11), .ZN(n405) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_15 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, N19, N20, N21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n412), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n413), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n414), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n415), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n416), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n417), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n418), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n419), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n420), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n421), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n422), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n423), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n424), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n425), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n426), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n427), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n428), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n429), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n430), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n431), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n432), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n433), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n434), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n435), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n436), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n437), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n438), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n439), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n440), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n441), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n442), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n443), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n444), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n445), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n446), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n447), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n448), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n449), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n450), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n451), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n452), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n453), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n454), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n455), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n456), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n457), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n458), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n459), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n460), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n461), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n462), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n463), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n464), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n465), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n466), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n467), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n468), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n469), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n470), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n471), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n472), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n473), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n474), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n475), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n476), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n477), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n478), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n479), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n480), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n481), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n482), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n483), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n484), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n485), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n486), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n487), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n488), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n489), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n490), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n491), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n492), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n493), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n494), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n495), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n496), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n497), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n498), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n499), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n500), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n501), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n502), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n503), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n504), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n505), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n506), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n507), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n508), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n509), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n510), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n511), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n512), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n513), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n514), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n515), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n516), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n517), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n518), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n519), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n520), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n521), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n522), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n523), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n524), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n525), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n526), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n527), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n528), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n529), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n530), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n531), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n532), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n533), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n534), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n535), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n536), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n537), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n538), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n539), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N20), .CK(clk), .QN(n399) );
  DFF_X1 \data_out_reg[5]  ( .D(N16), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(N10), .Z(n396) );
  BUF_X1 U4 ( .A(N10), .Z(n397) );
  BUF_X1 U5 ( .A(N10), .Z(n398) );
  BUF_X1 U6 ( .A(N11), .Z(n395) );
  NAND2_X1 U7 ( .A1(n663), .A2(n683), .ZN(n672) );
  NAND2_X1 U8 ( .A1(n663), .A2(n673), .ZN(n662) );
  NAND2_X1 U9 ( .A1(n684), .A2(n683), .ZN(n693) );
  NAND2_X1 U10 ( .A1(n673), .A2(n684), .ZN(n682) );
  NAND2_X1 U11 ( .A1(n605), .A2(n684), .ZN(n614) );
  NAND2_X1 U12 ( .A1(n595), .A2(n684), .ZN(n604) );
  NAND2_X1 U13 ( .A1(n605), .A2(n663), .ZN(n594) );
  NAND2_X1 U14 ( .A1(n595), .A2(n663), .ZN(n585) );
  NAND2_X1 U15 ( .A1(n644), .A2(n683), .ZN(n653) );
  NAND2_X1 U16 ( .A1(n644), .A2(n673), .ZN(n643) );
  NAND2_X1 U17 ( .A1(n625), .A2(n683), .ZN(n634) );
  NAND2_X1 U18 ( .A1(n625), .A2(n673), .ZN(n623) );
  NAND2_X1 U19 ( .A1(n605), .A2(n644), .ZN(n576) );
  NAND2_X1 U20 ( .A1(n595), .A2(n644), .ZN(n567) );
  NAND2_X1 U21 ( .A1(n605), .A2(n625), .ZN(n558) );
  NAND2_X1 U22 ( .A1(n595), .A2(n625), .ZN(n548) );
  AND2_X1 U23 ( .A1(n549), .A2(N10), .ZN(n595) );
  AND2_X1 U24 ( .A1(n549), .A2(n401), .ZN(n605) );
  AND2_X1 U25 ( .A1(N10), .A2(n624), .ZN(n673) );
  AND2_X1 U26 ( .A1(n624), .A2(n401), .ZN(n683) );
  OAI21_X1 U27 ( .B1(n693), .B2(n411), .A(n692), .ZN(n539) );
  NAND2_X1 U28 ( .A1(\mem[0][0] ), .A2(n693), .ZN(n692) );
  OAI21_X1 U29 ( .B1(n693), .B2(n410), .A(n691), .ZN(n538) );
  NAND2_X1 U30 ( .A1(\mem[0][1] ), .A2(n693), .ZN(n691) );
  OAI21_X1 U31 ( .B1(n693), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U32 ( .A1(\mem[0][2] ), .A2(n693), .ZN(n690) );
  OAI21_X1 U33 ( .B1(n693), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U34 ( .A1(\mem[0][3] ), .A2(n693), .ZN(n689) );
  OAI21_X1 U35 ( .B1(n693), .B2(n407), .A(n688), .ZN(n535) );
  NAND2_X1 U36 ( .A1(\mem[0][4] ), .A2(n693), .ZN(n688) );
  OAI21_X1 U37 ( .B1(n693), .B2(n406), .A(n687), .ZN(n534) );
  NAND2_X1 U38 ( .A1(\mem[0][5] ), .A2(n693), .ZN(n687) );
  OAI21_X1 U39 ( .B1(n693), .B2(n405), .A(n686), .ZN(n533) );
  NAND2_X1 U40 ( .A1(\mem[0][6] ), .A2(n693), .ZN(n686) );
  OAI21_X1 U41 ( .B1(n693), .B2(n404), .A(n685), .ZN(n532) );
  NAND2_X1 U42 ( .A1(\mem[0][7] ), .A2(n693), .ZN(n685) );
  OAI21_X1 U43 ( .B1(n411), .B2(n672), .A(n671), .ZN(n523) );
  NAND2_X1 U44 ( .A1(\mem[2][0] ), .A2(n672), .ZN(n671) );
  OAI21_X1 U45 ( .B1(n410), .B2(n672), .A(n670), .ZN(n522) );
  NAND2_X1 U46 ( .A1(\mem[2][1] ), .A2(n672), .ZN(n670) );
  OAI21_X1 U47 ( .B1(n409), .B2(n672), .A(n669), .ZN(n521) );
  NAND2_X1 U48 ( .A1(\mem[2][2] ), .A2(n672), .ZN(n669) );
  OAI21_X1 U49 ( .B1(n408), .B2(n672), .A(n668), .ZN(n520) );
  NAND2_X1 U50 ( .A1(\mem[2][3] ), .A2(n672), .ZN(n668) );
  OAI21_X1 U51 ( .B1(n407), .B2(n672), .A(n667), .ZN(n519) );
  NAND2_X1 U52 ( .A1(\mem[2][4] ), .A2(n672), .ZN(n667) );
  OAI21_X1 U53 ( .B1(n406), .B2(n672), .A(n666), .ZN(n518) );
  NAND2_X1 U54 ( .A1(\mem[2][5] ), .A2(n672), .ZN(n666) );
  OAI21_X1 U55 ( .B1(n405), .B2(n672), .A(n665), .ZN(n517) );
  NAND2_X1 U56 ( .A1(\mem[2][6] ), .A2(n672), .ZN(n665) );
  OAI21_X1 U57 ( .B1(n404), .B2(n672), .A(n664), .ZN(n516) );
  NAND2_X1 U58 ( .A1(\mem[2][7] ), .A2(n672), .ZN(n664) );
  OAI21_X1 U59 ( .B1(n411), .B2(n662), .A(n661), .ZN(n515) );
  NAND2_X1 U60 ( .A1(\mem[3][0] ), .A2(n662), .ZN(n661) );
  OAI21_X1 U61 ( .B1(n410), .B2(n662), .A(n660), .ZN(n514) );
  NAND2_X1 U62 ( .A1(\mem[3][1] ), .A2(n662), .ZN(n660) );
  OAI21_X1 U63 ( .B1(n409), .B2(n662), .A(n659), .ZN(n513) );
  NAND2_X1 U64 ( .A1(\mem[3][2] ), .A2(n662), .ZN(n659) );
  OAI21_X1 U65 ( .B1(n408), .B2(n662), .A(n658), .ZN(n512) );
  NAND2_X1 U66 ( .A1(\mem[3][3] ), .A2(n662), .ZN(n658) );
  OAI21_X1 U67 ( .B1(n407), .B2(n662), .A(n657), .ZN(n511) );
  NAND2_X1 U68 ( .A1(\mem[3][4] ), .A2(n662), .ZN(n657) );
  OAI21_X1 U69 ( .B1(n406), .B2(n662), .A(n656), .ZN(n510) );
  NAND2_X1 U70 ( .A1(\mem[3][5] ), .A2(n662), .ZN(n656) );
  OAI21_X1 U71 ( .B1(n405), .B2(n662), .A(n655), .ZN(n509) );
  NAND2_X1 U72 ( .A1(\mem[3][6] ), .A2(n662), .ZN(n655) );
  OAI21_X1 U73 ( .B1(n404), .B2(n662), .A(n654), .ZN(n508) );
  NAND2_X1 U74 ( .A1(\mem[3][7] ), .A2(n662), .ZN(n654) );
  NOR2_X1 U75 ( .A1(n403), .A2(N13), .ZN(n624) );
  INV_X1 U76 ( .A(wr_en), .ZN(n403) );
  OAI21_X1 U77 ( .B1(n411), .B2(n682), .A(n681), .ZN(n531) );
  NAND2_X1 U78 ( .A1(\mem[1][0] ), .A2(n682), .ZN(n681) );
  OAI21_X1 U79 ( .B1(n410), .B2(n682), .A(n680), .ZN(n530) );
  NAND2_X1 U80 ( .A1(\mem[1][1] ), .A2(n682), .ZN(n680) );
  OAI21_X1 U81 ( .B1(n409), .B2(n682), .A(n679), .ZN(n529) );
  NAND2_X1 U82 ( .A1(\mem[1][2] ), .A2(n682), .ZN(n679) );
  OAI21_X1 U83 ( .B1(n408), .B2(n682), .A(n678), .ZN(n528) );
  NAND2_X1 U84 ( .A1(\mem[1][3] ), .A2(n682), .ZN(n678) );
  OAI21_X1 U85 ( .B1(n407), .B2(n682), .A(n677), .ZN(n527) );
  NAND2_X1 U86 ( .A1(\mem[1][4] ), .A2(n682), .ZN(n677) );
  OAI21_X1 U87 ( .B1(n406), .B2(n682), .A(n676), .ZN(n526) );
  NAND2_X1 U88 ( .A1(\mem[1][5] ), .A2(n682), .ZN(n676) );
  OAI21_X1 U89 ( .B1(n405), .B2(n682), .A(n675), .ZN(n525) );
  NAND2_X1 U90 ( .A1(\mem[1][6] ), .A2(n682), .ZN(n675) );
  OAI21_X1 U91 ( .B1(n404), .B2(n682), .A(n674), .ZN(n524) );
  NAND2_X1 U92 ( .A1(\mem[1][7] ), .A2(n682), .ZN(n674) );
  OAI21_X1 U93 ( .B1(n411), .B2(n653), .A(n652), .ZN(n507) );
  NAND2_X1 U94 ( .A1(\mem[4][0] ), .A2(n653), .ZN(n652) );
  OAI21_X1 U95 ( .B1(n410), .B2(n653), .A(n651), .ZN(n506) );
  NAND2_X1 U96 ( .A1(\mem[4][1] ), .A2(n653), .ZN(n651) );
  OAI21_X1 U97 ( .B1(n409), .B2(n653), .A(n650), .ZN(n505) );
  NAND2_X1 U98 ( .A1(\mem[4][2] ), .A2(n653), .ZN(n650) );
  OAI21_X1 U99 ( .B1(n408), .B2(n653), .A(n649), .ZN(n504) );
  NAND2_X1 U100 ( .A1(\mem[4][3] ), .A2(n653), .ZN(n649) );
  OAI21_X1 U101 ( .B1(n407), .B2(n653), .A(n648), .ZN(n503) );
  NAND2_X1 U102 ( .A1(\mem[4][4] ), .A2(n653), .ZN(n648) );
  OAI21_X1 U103 ( .B1(n406), .B2(n653), .A(n647), .ZN(n502) );
  NAND2_X1 U104 ( .A1(\mem[4][5] ), .A2(n653), .ZN(n647) );
  OAI21_X1 U105 ( .B1(n405), .B2(n653), .A(n646), .ZN(n501) );
  NAND2_X1 U106 ( .A1(\mem[4][6] ), .A2(n653), .ZN(n646) );
  OAI21_X1 U107 ( .B1(n404), .B2(n653), .A(n645), .ZN(n500) );
  NAND2_X1 U108 ( .A1(\mem[4][7] ), .A2(n653), .ZN(n645) );
  OAI21_X1 U109 ( .B1(n411), .B2(n643), .A(n642), .ZN(n499) );
  NAND2_X1 U110 ( .A1(\mem[5][0] ), .A2(n643), .ZN(n642) );
  OAI21_X1 U111 ( .B1(n410), .B2(n643), .A(n641), .ZN(n498) );
  NAND2_X1 U112 ( .A1(\mem[5][1] ), .A2(n643), .ZN(n641) );
  OAI21_X1 U113 ( .B1(n409), .B2(n643), .A(n640), .ZN(n497) );
  NAND2_X1 U114 ( .A1(\mem[5][2] ), .A2(n643), .ZN(n640) );
  OAI21_X1 U115 ( .B1(n408), .B2(n643), .A(n639), .ZN(n496) );
  NAND2_X1 U116 ( .A1(\mem[5][3] ), .A2(n643), .ZN(n639) );
  OAI21_X1 U117 ( .B1(n407), .B2(n643), .A(n638), .ZN(n495) );
  NAND2_X1 U118 ( .A1(\mem[5][4] ), .A2(n643), .ZN(n638) );
  OAI21_X1 U119 ( .B1(n406), .B2(n643), .A(n637), .ZN(n494) );
  NAND2_X1 U120 ( .A1(\mem[5][5] ), .A2(n643), .ZN(n637) );
  OAI21_X1 U121 ( .B1(n405), .B2(n643), .A(n636), .ZN(n493) );
  NAND2_X1 U122 ( .A1(\mem[5][6] ), .A2(n643), .ZN(n636) );
  OAI21_X1 U123 ( .B1(n404), .B2(n643), .A(n635), .ZN(n492) );
  NAND2_X1 U124 ( .A1(\mem[5][7] ), .A2(n643), .ZN(n635) );
  OAI21_X1 U125 ( .B1(n411), .B2(n634), .A(n633), .ZN(n491) );
  NAND2_X1 U126 ( .A1(\mem[6][0] ), .A2(n634), .ZN(n633) );
  OAI21_X1 U127 ( .B1(n410), .B2(n634), .A(n632), .ZN(n490) );
  NAND2_X1 U128 ( .A1(\mem[6][1] ), .A2(n634), .ZN(n632) );
  OAI21_X1 U129 ( .B1(n409), .B2(n634), .A(n631), .ZN(n489) );
  NAND2_X1 U130 ( .A1(\mem[6][2] ), .A2(n634), .ZN(n631) );
  OAI21_X1 U131 ( .B1(n408), .B2(n634), .A(n630), .ZN(n488) );
  NAND2_X1 U132 ( .A1(\mem[6][3] ), .A2(n634), .ZN(n630) );
  OAI21_X1 U133 ( .B1(n407), .B2(n634), .A(n629), .ZN(n487) );
  NAND2_X1 U134 ( .A1(\mem[6][4] ), .A2(n634), .ZN(n629) );
  OAI21_X1 U135 ( .B1(n406), .B2(n634), .A(n628), .ZN(n486) );
  NAND2_X1 U136 ( .A1(\mem[6][5] ), .A2(n634), .ZN(n628) );
  OAI21_X1 U137 ( .B1(n405), .B2(n634), .A(n627), .ZN(n485) );
  NAND2_X1 U138 ( .A1(\mem[6][6] ), .A2(n634), .ZN(n627) );
  OAI21_X1 U139 ( .B1(n404), .B2(n634), .A(n626), .ZN(n484) );
  NAND2_X1 U140 ( .A1(\mem[6][7] ), .A2(n634), .ZN(n626) );
  OAI21_X1 U141 ( .B1(n411), .B2(n623), .A(n622), .ZN(n483) );
  NAND2_X1 U142 ( .A1(\mem[7][0] ), .A2(n623), .ZN(n622) );
  OAI21_X1 U143 ( .B1(n410), .B2(n623), .A(n621), .ZN(n482) );
  NAND2_X1 U144 ( .A1(\mem[7][1] ), .A2(n623), .ZN(n621) );
  OAI21_X1 U145 ( .B1(n409), .B2(n623), .A(n620), .ZN(n481) );
  NAND2_X1 U146 ( .A1(\mem[7][2] ), .A2(n623), .ZN(n620) );
  OAI21_X1 U147 ( .B1(n408), .B2(n623), .A(n619), .ZN(n480) );
  NAND2_X1 U148 ( .A1(\mem[7][3] ), .A2(n623), .ZN(n619) );
  OAI21_X1 U149 ( .B1(n407), .B2(n623), .A(n618), .ZN(n479) );
  NAND2_X1 U150 ( .A1(\mem[7][4] ), .A2(n623), .ZN(n618) );
  OAI21_X1 U151 ( .B1(n406), .B2(n623), .A(n617), .ZN(n478) );
  NAND2_X1 U152 ( .A1(\mem[7][5] ), .A2(n623), .ZN(n617) );
  OAI21_X1 U153 ( .B1(n405), .B2(n623), .A(n616), .ZN(n477) );
  NAND2_X1 U154 ( .A1(\mem[7][6] ), .A2(n623), .ZN(n616) );
  OAI21_X1 U155 ( .B1(n404), .B2(n623), .A(n615), .ZN(n476) );
  NAND2_X1 U156 ( .A1(\mem[7][7] ), .A2(n623), .ZN(n615) );
  OAI21_X1 U157 ( .B1(n411), .B2(n614), .A(n613), .ZN(n475) );
  NAND2_X1 U158 ( .A1(\mem[8][0] ), .A2(n614), .ZN(n613) );
  OAI21_X1 U159 ( .B1(n410), .B2(n614), .A(n612), .ZN(n474) );
  NAND2_X1 U160 ( .A1(\mem[8][1] ), .A2(n614), .ZN(n612) );
  OAI21_X1 U161 ( .B1(n409), .B2(n614), .A(n611), .ZN(n473) );
  NAND2_X1 U162 ( .A1(\mem[8][2] ), .A2(n614), .ZN(n611) );
  OAI21_X1 U163 ( .B1(n408), .B2(n614), .A(n610), .ZN(n472) );
  NAND2_X1 U164 ( .A1(\mem[8][3] ), .A2(n614), .ZN(n610) );
  OAI21_X1 U165 ( .B1(n407), .B2(n614), .A(n609), .ZN(n471) );
  NAND2_X1 U166 ( .A1(\mem[8][4] ), .A2(n614), .ZN(n609) );
  OAI21_X1 U167 ( .B1(n406), .B2(n614), .A(n608), .ZN(n470) );
  NAND2_X1 U168 ( .A1(\mem[8][5] ), .A2(n614), .ZN(n608) );
  OAI21_X1 U169 ( .B1(n405), .B2(n614), .A(n607), .ZN(n469) );
  NAND2_X1 U170 ( .A1(\mem[8][6] ), .A2(n614), .ZN(n607) );
  OAI21_X1 U171 ( .B1(n404), .B2(n614), .A(n606), .ZN(n468) );
  NAND2_X1 U172 ( .A1(\mem[8][7] ), .A2(n614), .ZN(n606) );
  OAI21_X1 U173 ( .B1(n411), .B2(n604), .A(n603), .ZN(n467) );
  NAND2_X1 U174 ( .A1(\mem[9][0] ), .A2(n604), .ZN(n603) );
  OAI21_X1 U175 ( .B1(n410), .B2(n604), .A(n602), .ZN(n466) );
  NAND2_X1 U176 ( .A1(\mem[9][1] ), .A2(n604), .ZN(n602) );
  OAI21_X1 U177 ( .B1(n409), .B2(n604), .A(n601), .ZN(n465) );
  NAND2_X1 U178 ( .A1(\mem[9][2] ), .A2(n604), .ZN(n601) );
  OAI21_X1 U179 ( .B1(n408), .B2(n604), .A(n600), .ZN(n464) );
  NAND2_X1 U180 ( .A1(\mem[9][3] ), .A2(n604), .ZN(n600) );
  OAI21_X1 U181 ( .B1(n407), .B2(n604), .A(n599), .ZN(n463) );
  NAND2_X1 U182 ( .A1(\mem[9][4] ), .A2(n604), .ZN(n599) );
  OAI21_X1 U183 ( .B1(n406), .B2(n604), .A(n598), .ZN(n462) );
  NAND2_X1 U184 ( .A1(\mem[9][5] ), .A2(n604), .ZN(n598) );
  OAI21_X1 U185 ( .B1(n405), .B2(n604), .A(n597), .ZN(n461) );
  NAND2_X1 U186 ( .A1(\mem[9][6] ), .A2(n604), .ZN(n597) );
  OAI21_X1 U187 ( .B1(n404), .B2(n604), .A(n596), .ZN(n460) );
  NAND2_X1 U188 ( .A1(\mem[9][7] ), .A2(n604), .ZN(n596) );
  OAI21_X1 U189 ( .B1(n411), .B2(n594), .A(n593), .ZN(n459) );
  NAND2_X1 U190 ( .A1(\mem[10][0] ), .A2(n594), .ZN(n593) );
  OAI21_X1 U191 ( .B1(n410), .B2(n594), .A(n592), .ZN(n458) );
  NAND2_X1 U192 ( .A1(\mem[10][1] ), .A2(n594), .ZN(n592) );
  OAI21_X1 U193 ( .B1(n409), .B2(n594), .A(n591), .ZN(n457) );
  NAND2_X1 U194 ( .A1(\mem[10][2] ), .A2(n594), .ZN(n591) );
  OAI21_X1 U195 ( .B1(n408), .B2(n594), .A(n590), .ZN(n456) );
  NAND2_X1 U196 ( .A1(\mem[10][3] ), .A2(n594), .ZN(n590) );
  OAI21_X1 U197 ( .B1(n407), .B2(n594), .A(n589), .ZN(n455) );
  NAND2_X1 U198 ( .A1(\mem[10][4] ), .A2(n594), .ZN(n589) );
  OAI21_X1 U199 ( .B1(n406), .B2(n594), .A(n588), .ZN(n454) );
  NAND2_X1 U200 ( .A1(\mem[10][5] ), .A2(n594), .ZN(n588) );
  OAI21_X1 U201 ( .B1(n405), .B2(n594), .A(n587), .ZN(n453) );
  NAND2_X1 U202 ( .A1(\mem[10][6] ), .A2(n594), .ZN(n587) );
  OAI21_X1 U203 ( .B1(n404), .B2(n594), .A(n586), .ZN(n452) );
  NAND2_X1 U204 ( .A1(\mem[10][7] ), .A2(n594), .ZN(n586) );
  OAI21_X1 U205 ( .B1(n411), .B2(n585), .A(n584), .ZN(n451) );
  NAND2_X1 U206 ( .A1(\mem[11][0] ), .A2(n585), .ZN(n584) );
  OAI21_X1 U207 ( .B1(n410), .B2(n585), .A(n583), .ZN(n450) );
  NAND2_X1 U208 ( .A1(\mem[11][1] ), .A2(n585), .ZN(n583) );
  OAI21_X1 U209 ( .B1(n409), .B2(n585), .A(n582), .ZN(n449) );
  NAND2_X1 U210 ( .A1(\mem[11][2] ), .A2(n585), .ZN(n582) );
  OAI21_X1 U211 ( .B1(n408), .B2(n585), .A(n581), .ZN(n448) );
  NAND2_X1 U212 ( .A1(\mem[11][3] ), .A2(n585), .ZN(n581) );
  OAI21_X1 U213 ( .B1(n407), .B2(n585), .A(n580), .ZN(n447) );
  NAND2_X1 U214 ( .A1(\mem[11][4] ), .A2(n585), .ZN(n580) );
  OAI21_X1 U215 ( .B1(n406), .B2(n585), .A(n579), .ZN(n446) );
  NAND2_X1 U216 ( .A1(\mem[11][5] ), .A2(n585), .ZN(n579) );
  OAI21_X1 U217 ( .B1(n405), .B2(n585), .A(n578), .ZN(n445) );
  NAND2_X1 U218 ( .A1(\mem[11][6] ), .A2(n585), .ZN(n578) );
  OAI21_X1 U219 ( .B1(n404), .B2(n585), .A(n577), .ZN(n444) );
  NAND2_X1 U220 ( .A1(\mem[11][7] ), .A2(n585), .ZN(n577) );
  OAI21_X1 U221 ( .B1(n411), .B2(n576), .A(n575), .ZN(n443) );
  NAND2_X1 U222 ( .A1(\mem[12][0] ), .A2(n576), .ZN(n575) );
  OAI21_X1 U223 ( .B1(n410), .B2(n576), .A(n574), .ZN(n442) );
  NAND2_X1 U224 ( .A1(\mem[12][1] ), .A2(n576), .ZN(n574) );
  OAI21_X1 U225 ( .B1(n409), .B2(n576), .A(n573), .ZN(n441) );
  NAND2_X1 U226 ( .A1(\mem[12][2] ), .A2(n576), .ZN(n573) );
  OAI21_X1 U227 ( .B1(n408), .B2(n576), .A(n572), .ZN(n440) );
  NAND2_X1 U228 ( .A1(\mem[12][3] ), .A2(n576), .ZN(n572) );
  OAI21_X1 U229 ( .B1(n407), .B2(n576), .A(n571), .ZN(n439) );
  NAND2_X1 U230 ( .A1(\mem[12][4] ), .A2(n576), .ZN(n571) );
  OAI21_X1 U231 ( .B1(n406), .B2(n576), .A(n570), .ZN(n438) );
  NAND2_X1 U232 ( .A1(\mem[12][5] ), .A2(n576), .ZN(n570) );
  OAI21_X1 U233 ( .B1(n405), .B2(n576), .A(n569), .ZN(n437) );
  NAND2_X1 U234 ( .A1(\mem[12][6] ), .A2(n576), .ZN(n569) );
  OAI21_X1 U235 ( .B1(n404), .B2(n576), .A(n568), .ZN(n436) );
  NAND2_X1 U236 ( .A1(\mem[12][7] ), .A2(n576), .ZN(n568) );
  OAI21_X1 U237 ( .B1(n411), .B2(n567), .A(n566), .ZN(n435) );
  NAND2_X1 U238 ( .A1(\mem[13][0] ), .A2(n567), .ZN(n566) );
  OAI21_X1 U239 ( .B1(n410), .B2(n567), .A(n565), .ZN(n434) );
  NAND2_X1 U240 ( .A1(\mem[13][1] ), .A2(n567), .ZN(n565) );
  OAI21_X1 U241 ( .B1(n409), .B2(n567), .A(n564), .ZN(n433) );
  NAND2_X1 U242 ( .A1(\mem[13][2] ), .A2(n567), .ZN(n564) );
  OAI21_X1 U243 ( .B1(n408), .B2(n567), .A(n563), .ZN(n432) );
  NAND2_X1 U244 ( .A1(\mem[13][3] ), .A2(n567), .ZN(n563) );
  OAI21_X1 U245 ( .B1(n407), .B2(n567), .A(n562), .ZN(n431) );
  NAND2_X1 U246 ( .A1(\mem[13][4] ), .A2(n567), .ZN(n562) );
  OAI21_X1 U247 ( .B1(n406), .B2(n567), .A(n561), .ZN(n430) );
  NAND2_X1 U248 ( .A1(\mem[13][5] ), .A2(n567), .ZN(n561) );
  OAI21_X1 U249 ( .B1(n405), .B2(n567), .A(n560), .ZN(n429) );
  NAND2_X1 U250 ( .A1(\mem[13][6] ), .A2(n567), .ZN(n560) );
  OAI21_X1 U251 ( .B1(n404), .B2(n567), .A(n559), .ZN(n428) );
  NAND2_X1 U252 ( .A1(\mem[13][7] ), .A2(n567), .ZN(n559) );
  OAI21_X1 U253 ( .B1(n411), .B2(n558), .A(n557), .ZN(n427) );
  NAND2_X1 U254 ( .A1(\mem[14][0] ), .A2(n558), .ZN(n557) );
  OAI21_X1 U255 ( .B1(n410), .B2(n558), .A(n556), .ZN(n426) );
  NAND2_X1 U256 ( .A1(\mem[14][1] ), .A2(n558), .ZN(n556) );
  OAI21_X1 U257 ( .B1(n409), .B2(n558), .A(n555), .ZN(n425) );
  NAND2_X1 U258 ( .A1(\mem[14][2] ), .A2(n558), .ZN(n555) );
  OAI21_X1 U259 ( .B1(n408), .B2(n558), .A(n554), .ZN(n424) );
  NAND2_X1 U260 ( .A1(\mem[14][3] ), .A2(n558), .ZN(n554) );
  OAI21_X1 U261 ( .B1(n407), .B2(n558), .A(n553), .ZN(n423) );
  NAND2_X1 U262 ( .A1(\mem[14][4] ), .A2(n558), .ZN(n553) );
  OAI21_X1 U263 ( .B1(n406), .B2(n558), .A(n552), .ZN(n422) );
  NAND2_X1 U264 ( .A1(\mem[14][5] ), .A2(n558), .ZN(n552) );
  OAI21_X1 U265 ( .B1(n405), .B2(n558), .A(n551), .ZN(n421) );
  NAND2_X1 U266 ( .A1(\mem[14][6] ), .A2(n558), .ZN(n551) );
  OAI21_X1 U267 ( .B1(n404), .B2(n558), .A(n550), .ZN(n420) );
  NAND2_X1 U268 ( .A1(\mem[14][7] ), .A2(n558), .ZN(n550) );
  OAI21_X1 U269 ( .B1(n411), .B2(n548), .A(n547), .ZN(n419) );
  NAND2_X1 U270 ( .A1(\mem[15][0] ), .A2(n548), .ZN(n547) );
  OAI21_X1 U271 ( .B1(n410), .B2(n548), .A(n546), .ZN(n418) );
  NAND2_X1 U272 ( .A1(\mem[15][1] ), .A2(n548), .ZN(n546) );
  OAI21_X1 U273 ( .B1(n409), .B2(n548), .A(n545), .ZN(n417) );
  NAND2_X1 U274 ( .A1(\mem[15][2] ), .A2(n548), .ZN(n545) );
  OAI21_X1 U275 ( .B1(n408), .B2(n548), .A(n544), .ZN(n416) );
  NAND2_X1 U276 ( .A1(\mem[15][3] ), .A2(n548), .ZN(n544) );
  OAI21_X1 U277 ( .B1(n407), .B2(n548), .A(n543), .ZN(n415) );
  NAND2_X1 U278 ( .A1(\mem[15][4] ), .A2(n548), .ZN(n543) );
  OAI21_X1 U279 ( .B1(n406), .B2(n548), .A(n542), .ZN(n414) );
  NAND2_X1 U280 ( .A1(\mem[15][5] ), .A2(n548), .ZN(n542) );
  OAI21_X1 U281 ( .B1(n405), .B2(n548), .A(n541), .ZN(n413) );
  NAND2_X1 U282 ( .A1(\mem[15][6] ), .A2(n548), .ZN(n541) );
  OAI21_X1 U283 ( .B1(n404), .B2(n548), .A(n540), .ZN(n412) );
  NAND2_X1 U284 ( .A1(\mem[15][7] ), .A2(n548), .ZN(n540) );
  AND2_X1 U285 ( .A1(N13), .A2(wr_en), .ZN(n549) );
  NOR2_X1 U286 ( .A1(N11), .A2(N12), .ZN(n684) );
  NOR2_X1 U287 ( .A1(n402), .A2(N12), .ZN(n663) );
  AND2_X1 U288 ( .A1(N12), .A2(n402), .ZN(n644) );
  AND2_X1 U289 ( .A1(N12), .A2(N11), .ZN(n625) );
  INV_X1 U290 ( .A(data_in[0]), .ZN(n411) );
  INV_X1 U291 ( .A(data_in[1]), .ZN(n410) );
  INV_X1 U292 ( .A(data_in[2]), .ZN(n409) );
  INV_X1 U293 ( .A(data_in[3]), .ZN(n408) );
  INV_X1 U294 ( .A(data_in[4]), .ZN(n407) );
  INV_X1 U295 ( .A(data_in[5]), .ZN(n406) );
  INV_X1 U296 ( .A(data_in[6]), .ZN(n405) );
  INV_X1 U297 ( .A(data_in[7]), .ZN(n404) );
  MUX2_X1 U298 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n398), .Z(n1) );
  MUX2_X1 U299 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n396), .Z(n2) );
  MUX2_X1 U300 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U301 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n398), .Z(n4) );
  MUX2_X1 U302 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n397), .Z(n5) );
  MUX2_X1 U303 ( .A(n5), .B(n4), .S(N11), .Z(n6) );
  MUX2_X1 U304 ( .A(n6), .B(n3), .S(N12), .Z(n7) );
  MUX2_X1 U305 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n397), .Z(n8) );
  MUX2_X1 U306 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(N10), .Z(n9) );
  MUX2_X1 U307 ( .A(n9), .B(n8), .S(N11), .Z(n10) );
  MUX2_X1 U308 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(N10), .Z(n11) );
  MUX2_X1 U309 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n294) );
  MUX2_X1 U310 ( .A(n294), .B(n11), .S(n395), .Z(n295) );
  MUX2_X1 U311 ( .A(n295), .B(n10), .S(N12), .Z(n296) );
  MUX2_X1 U312 ( .A(n296), .B(n7), .S(N13), .Z(N21) );
  MUX2_X1 U313 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n396), .Z(n297) );
  MUX2_X1 U314 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(N10), .Z(n298) );
  MUX2_X1 U315 ( .A(n298), .B(n297), .S(N11), .Z(n299) );
  MUX2_X1 U316 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(N10), .Z(n300) );
  MUX2_X1 U317 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(N10), .Z(n301) );
  MUX2_X1 U318 ( .A(n301), .B(n300), .S(n395), .Z(n302) );
  MUX2_X1 U319 ( .A(n302), .B(n299), .S(N12), .Z(n303) );
  MUX2_X1 U320 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n398), .Z(n304) );
  MUX2_X1 U321 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(N10), .Z(n305) );
  MUX2_X1 U322 ( .A(n305), .B(n304), .S(N11), .Z(n306) );
  MUX2_X1 U323 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(N10), .Z(n307) );
  MUX2_X1 U324 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(N10), .Z(n308) );
  MUX2_X1 U325 ( .A(n308), .B(n307), .S(n395), .Z(n309) );
  MUX2_X1 U326 ( .A(n309), .B(n306), .S(N12), .Z(n310) );
  MUX2_X1 U327 ( .A(n310), .B(n303), .S(N13), .Z(N20) );
  MUX2_X1 U328 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(N10), .Z(n311) );
  MUX2_X1 U329 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n397), .Z(n312) );
  MUX2_X1 U330 ( .A(n312), .B(n311), .S(N11), .Z(n313) );
  MUX2_X1 U331 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n396), .Z(n314) );
  MUX2_X1 U332 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(N10), .Z(n315) );
  MUX2_X1 U333 ( .A(n315), .B(n314), .S(N11), .Z(n316) );
  MUX2_X1 U334 ( .A(n316), .B(n313), .S(N12), .Z(n317) );
  MUX2_X1 U335 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n396), .Z(n318) );
  MUX2_X1 U336 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(N10), .Z(n319) );
  MUX2_X1 U337 ( .A(n319), .B(n318), .S(N11), .Z(n320) );
  MUX2_X1 U338 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(N10), .Z(n321) );
  MUX2_X1 U339 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(N10), .Z(n322) );
  MUX2_X1 U340 ( .A(n322), .B(n321), .S(N11), .Z(n323) );
  MUX2_X1 U341 ( .A(n323), .B(n320), .S(N12), .Z(n324) );
  MUX2_X1 U342 ( .A(n324), .B(n317), .S(N13), .Z(N19) );
  MUX2_X1 U343 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n397), .Z(n325) );
  MUX2_X1 U344 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n398), .Z(n326) );
  MUX2_X1 U345 ( .A(n326), .B(n325), .S(N11), .Z(n327) );
  MUX2_X1 U346 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n397), .Z(n328) );
  MUX2_X1 U347 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n329) );
  MUX2_X1 U348 ( .A(n329), .B(n328), .S(N11), .Z(n330) );
  MUX2_X1 U349 ( .A(n330), .B(n327), .S(N12), .Z(n331) );
  MUX2_X1 U350 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n396), .Z(n332) );
  MUX2_X1 U351 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n396), .Z(n333) );
  MUX2_X1 U352 ( .A(n333), .B(n332), .S(N11), .Z(n334) );
  MUX2_X1 U353 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n396), .Z(n335) );
  MUX2_X1 U354 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n396), .Z(n336) );
  MUX2_X1 U355 ( .A(n336), .B(n335), .S(N11), .Z(n337) );
  MUX2_X1 U356 ( .A(n337), .B(n334), .S(N12), .Z(n338) );
  MUX2_X1 U357 ( .A(n338), .B(n331), .S(N13), .Z(N18) );
  MUX2_X1 U358 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n396), .Z(n339) );
  MUX2_X1 U359 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n396), .Z(n340) );
  MUX2_X1 U360 ( .A(n340), .B(n339), .S(N11), .Z(n341) );
  MUX2_X1 U361 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n396), .Z(n342) );
  MUX2_X1 U362 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n396), .Z(n343) );
  MUX2_X1 U363 ( .A(n343), .B(n342), .S(N11), .Z(n344) );
  MUX2_X1 U364 ( .A(n344), .B(n341), .S(N12), .Z(n345) );
  MUX2_X1 U365 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n396), .Z(n346) );
  MUX2_X1 U366 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n396), .Z(n347) );
  MUX2_X1 U367 ( .A(n347), .B(n346), .S(N11), .Z(n348) );
  MUX2_X1 U368 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n396), .Z(n349) );
  MUX2_X1 U369 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n396), .Z(n350) );
  MUX2_X1 U370 ( .A(n350), .B(n349), .S(N11), .Z(n351) );
  MUX2_X1 U371 ( .A(n351), .B(n348), .S(N12), .Z(n352) );
  MUX2_X1 U372 ( .A(n352), .B(n345), .S(N13), .Z(N17) );
  MUX2_X1 U373 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n397), .Z(n353) );
  MUX2_X1 U374 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n397), .Z(n354) );
  MUX2_X1 U375 ( .A(n354), .B(n353), .S(n395), .Z(n355) );
  MUX2_X1 U376 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n397), .Z(n356) );
  MUX2_X1 U377 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n397), .Z(n357) );
  MUX2_X1 U378 ( .A(n357), .B(n356), .S(n395), .Z(n358) );
  MUX2_X1 U379 ( .A(n358), .B(n355), .S(N12), .Z(n359) );
  MUX2_X1 U380 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n397), .Z(n360) );
  MUX2_X1 U381 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n397), .Z(n361) );
  MUX2_X1 U382 ( .A(n361), .B(n360), .S(n395), .Z(n362) );
  MUX2_X1 U383 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n397), .Z(n363) );
  MUX2_X1 U384 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n397), .Z(n364) );
  MUX2_X1 U385 ( .A(n364), .B(n363), .S(n395), .Z(n365) );
  MUX2_X1 U386 ( .A(n365), .B(n362), .S(N12), .Z(n366) );
  MUX2_X1 U387 ( .A(n366), .B(n359), .S(N13), .Z(N16) );
  MUX2_X1 U388 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n397), .Z(n367) );
  MUX2_X1 U389 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n397), .Z(n368) );
  MUX2_X1 U390 ( .A(n368), .B(n367), .S(n395), .Z(n369) );
  MUX2_X1 U391 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n397), .Z(n370) );
  MUX2_X1 U392 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n397), .Z(n371) );
  MUX2_X1 U393 ( .A(n371), .B(n370), .S(n395), .Z(n372) );
  MUX2_X1 U394 ( .A(n372), .B(n369), .S(N12), .Z(n373) );
  MUX2_X1 U395 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n398), .Z(n374) );
  MUX2_X1 U396 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n398), .Z(n375) );
  MUX2_X1 U397 ( .A(n375), .B(n374), .S(n395), .Z(n376) );
  MUX2_X1 U398 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n398), .Z(n377) );
  MUX2_X1 U399 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n398), .Z(n378) );
  MUX2_X1 U400 ( .A(n378), .B(n377), .S(n395), .Z(n379) );
  MUX2_X1 U401 ( .A(n379), .B(n376), .S(N12), .Z(n380) );
  MUX2_X1 U402 ( .A(n380), .B(n373), .S(N13), .Z(N15) );
  MUX2_X1 U403 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n398), .Z(n381) );
  MUX2_X1 U404 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n398), .Z(n382) );
  MUX2_X1 U405 ( .A(n382), .B(n381), .S(n395), .Z(n383) );
  MUX2_X1 U406 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n398), .Z(n384) );
  MUX2_X1 U407 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n398), .Z(n385) );
  MUX2_X1 U408 ( .A(n385), .B(n384), .S(n395), .Z(n386) );
  MUX2_X1 U409 ( .A(n386), .B(n383), .S(N12), .Z(n387) );
  MUX2_X1 U410 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n398), .Z(n388) );
  MUX2_X1 U411 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n398), .Z(n389) );
  MUX2_X1 U412 ( .A(n389), .B(n388), .S(n395), .Z(n390) );
  MUX2_X1 U413 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n398), .Z(n391) );
  MUX2_X1 U414 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n398), .Z(n392) );
  MUX2_X1 U415 ( .A(n392), .B(n391), .S(n395), .Z(n393) );
  MUX2_X1 U416 ( .A(n393), .B(n390), .S(N12), .Z(n394) );
  MUX2_X1 U417 ( .A(n394), .B(n387), .S(N13), .Z(N14) );
  INV_X2 U418 ( .A(n399), .ZN(data_out[1]) );
  INV_X1 U419 ( .A(N10), .ZN(n401) );
  INV_X1 U420 ( .A(N11), .ZN(n402) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_14 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, N19, N20, N21, n1, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N20), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n412), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n413), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n414), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n415), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n416), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n417), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n418), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n419), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n420), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n421), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n422), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n423), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n424), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n425), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n426), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n427), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n428), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n429), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n430), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n431), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n432), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n433), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n434), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n435), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n436), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n437), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n438), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n439), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n440), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n441), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n442), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n443), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n444), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n445), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n446), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n447), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n448), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n449), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n450), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n451), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n452), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n453), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n454), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n455), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n456), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n457), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n458), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n459), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n460), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n461), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n462), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n463), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n464), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n465), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n466), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n467), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n468), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n469), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n470), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n471), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n472), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n473), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n474), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n475), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n476), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n477), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n478), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n479), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n480), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n481), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n482), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n483), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n484), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n485), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n486), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n487), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n488), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n489), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n490), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n491), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n492), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n493), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n494), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n495), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n496), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n497), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n498), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n499), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n500), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n501), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n502), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n503), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n504), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n505), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n506), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n507), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n508), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n509), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n510), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n511), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n512), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n513), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n514), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n515), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n516), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n517), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n518), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n519), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n520), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n521), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n522), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n523), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n524), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n525), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n526), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n527), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n528), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n529), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n530), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n531), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n532), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n533), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n534), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n535), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n536), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n537), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n538), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n539), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .QN(n1) );
  DFF_X2 \data_out_reg[5]  ( .D(N16), .CK(clk), .Q(data_out[5]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(N10), .Z(n398) );
  BUF_X1 U5 ( .A(N10), .Z(n399) );
  BUF_X1 U6 ( .A(N10), .Z(n400) );
  BUF_X1 U7 ( .A(N11), .Z(n397) );
  NAND2_X1 U8 ( .A1(n663), .A2(n683), .ZN(n672) );
  NAND2_X1 U9 ( .A1(n663), .A2(n673), .ZN(n662) );
  NAND2_X1 U10 ( .A1(n684), .A2(n683), .ZN(n693) );
  NAND2_X1 U11 ( .A1(n673), .A2(n684), .ZN(n682) );
  NAND2_X1 U12 ( .A1(n605), .A2(n684), .ZN(n614) );
  NAND2_X1 U13 ( .A1(n595), .A2(n684), .ZN(n604) );
  NAND2_X1 U14 ( .A1(n605), .A2(n663), .ZN(n594) );
  NAND2_X1 U15 ( .A1(n595), .A2(n663), .ZN(n585) );
  NAND2_X1 U16 ( .A1(n644), .A2(n683), .ZN(n653) );
  NAND2_X1 U17 ( .A1(n644), .A2(n673), .ZN(n643) );
  NAND2_X1 U18 ( .A1(n625), .A2(n683), .ZN(n634) );
  NAND2_X1 U19 ( .A1(n625), .A2(n673), .ZN(n623) );
  NAND2_X1 U20 ( .A1(n605), .A2(n644), .ZN(n576) );
  NAND2_X1 U21 ( .A1(n595), .A2(n644), .ZN(n567) );
  NAND2_X1 U22 ( .A1(n605), .A2(n625), .ZN(n558) );
  NAND2_X1 U23 ( .A1(n595), .A2(n625), .ZN(n548) );
  AND2_X1 U24 ( .A1(n549), .A2(N10), .ZN(n595) );
  AND2_X1 U25 ( .A1(n549), .A2(n401), .ZN(n605) );
  AND2_X1 U26 ( .A1(N10), .A2(n624), .ZN(n673) );
  AND2_X1 U27 ( .A1(n624), .A2(n401), .ZN(n683) );
  OAI21_X1 U28 ( .B1(n693), .B2(n411), .A(n692), .ZN(n539) );
  NAND2_X1 U29 ( .A1(\mem[0][0] ), .A2(n693), .ZN(n692) );
  OAI21_X1 U30 ( .B1(n693), .B2(n410), .A(n691), .ZN(n538) );
  NAND2_X1 U31 ( .A1(\mem[0][1] ), .A2(n693), .ZN(n691) );
  OAI21_X1 U32 ( .B1(n693), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U33 ( .A1(\mem[0][2] ), .A2(n693), .ZN(n690) );
  OAI21_X1 U34 ( .B1(n693), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U35 ( .A1(\mem[0][3] ), .A2(n693), .ZN(n689) );
  OAI21_X1 U36 ( .B1(n693), .B2(n407), .A(n688), .ZN(n535) );
  NAND2_X1 U37 ( .A1(\mem[0][4] ), .A2(n693), .ZN(n688) );
  OAI21_X1 U38 ( .B1(n693), .B2(n406), .A(n687), .ZN(n534) );
  NAND2_X1 U39 ( .A1(\mem[0][5] ), .A2(n693), .ZN(n687) );
  OAI21_X1 U40 ( .B1(n693), .B2(n405), .A(n686), .ZN(n533) );
  NAND2_X1 U41 ( .A1(\mem[0][6] ), .A2(n693), .ZN(n686) );
  OAI21_X1 U42 ( .B1(n693), .B2(n404), .A(n685), .ZN(n532) );
  NAND2_X1 U43 ( .A1(\mem[0][7] ), .A2(n693), .ZN(n685) );
  OAI21_X1 U44 ( .B1(n411), .B2(n672), .A(n671), .ZN(n523) );
  NAND2_X1 U45 ( .A1(\mem[2][0] ), .A2(n672), .ZN(n671) );
  OAI21_X1 U46 ( .B1(n410), .B2(n672), .A(n670), .ZN(n522) );
  NAND2_X1 U47 ( .A1(\mem[2][1] ), .A2(n672), .ZN(n670) );
  OAI21_X1 U48 ( .B1(n409), .B2(n672), .A(n669), .ZN(n521) );
  NAND2_X1 U49 ( .A1(\mem[2][2] ), .A2(n672), .ZN(n669) );
  OAI21_X1 U50 ( .B1(n408), .B2(n672), .A(n668), .ZN(n520) );
  NAND2_X1 U51 ( .A1(\mem[2][3] ), .A2(n672), .ZN(n668) );
  OAI21_X1 U52 ( .B1(n407), .B2(n672), .A(n667), .ZN(n519) );
  NAND2_X1 U53 ( .A1(\mem[2][4] ), .A2(n672), .ZN(n667) );
  OAI21_X1 U54 ( .B1(n406), .B2(n672), .A(n666), .ZN(n518) );
  NAND2_X1 U55 ( .A1(\mem[2][5] ), .A2(n672), .ZN(n666) );
  OAI21_X1 U56 ( .B1(n405), .B2(n672), .A(n665), .ZN(n517) );
  NAND2_X1 U57 ( .A1(\mem[2][6] ), .A2(n672), .ZN(n665) );
  OAI21_X1 U58 ( .B1(n404), .B2(n672), .A(n664), .ZN(n516) );
  NAND2_X1 U59 ( .A1(\mem[2][7] ), .A2(n672), .ZN(n664) );
  OAI21_X1 U60 ( .B1(n411), .B2(n662), .A(n661), .ZN(n515) );
  NAND2_X1 U61 ( .A1(\mem[3][0] ), .A2(n662), .ZN(n661) );
  OAI21_X1 U62 ( .B1(n410), .B2(n662), .A(n660), .ZN(n514) );
  NAND2_X1 U63 ( .A1(\mem[3][1] ), .A2(n662), .ZN(n660) );
  OAI21_X1 U64 ( .B1(n409), .B2(n662), .A(n659), .ZN(n513) );
  NAND2_X1 U65 ( .A1(\mem[3][2] ), .A2(n662), .ZN(n659) );
  OAI21_X1 U66 ( .B1(n408), .B2(n662), .A(n658), .ZN(n512) );
  NAND2_X1 U67 ( .A1(\mem[3][3] ), .A2(n662), .ZN(n658) );
  OAI21_X1 U68 ( .B1(n407), .B2(n662), .A(n657), .ZN(n511) );
  NAND2_X1 U69 ( .A1(\mem[3][4] ), .A2(n662), .ZN(n657) );
  OAI21_X1 U70 ( .B1(n406), .B2(n662), .A(n656), .ZN(n510) );
  NAND2_X1 U71 ( .A1(\mem[3][5] ), .A2(n662), .ZN(n656) );
  OAI21_X1 U72 ( .B1(n405), .B2(n662), .A(n655), .ZN(n509) );
  NAND2_X1 U73 ( .A1(\mem[3][6] ), .A2(n662), .ZN(n655) );
  OAI21_X1 U74 ( .B1(n404), .B2(n662), .A(n654), .ZN(n508) );
  NAND2_X1 U75 ( .A1(\mem[3][7] ), .A2(n662), .ZN(n654) );
  NOR2_X1 U76 ( .A1(n403), .A2(N13), .ZN(n624) );
  INV_X1 U77 ( .A(wr_en), .ZN(n403) );
  OAI21_X1 U78 ( .B1(n411), .B2(n682), .A(n681), .ZN(n531) );
  NAND2_X1 U79 ( .A1(\mem[1][0] ), .A2(n682), .ZN(n681) );
  OAI21_X1 U80 ( .B1(n410), .B2(n682), .A(n680), .ZN(n530) );
  NAND2_X1 U81 ( .A1(\mem[1][1] ), .A2(n682), .ZN(n680) );
  OAI21_X1 U82 ( .B1(n409), .B2(n682), .A(n679), .ZN(n529) );
  NAND2_X1 U83 ( .A1(\mem[1][2] ), .A2(n682), .ZN(n679) );
  OAI21_X1 U84 ( .B1(n408), .B2(n682), .A(n678), .ZN(n528) );
  NAND2_X1 U85 ( .A1(\mem[1][3] ), .A2(n682), .ZN(n678) );
  OAI21_X1 U86 ( .B1(n407), .B2(n682), .A(n677), .ZN(n527) );
  NAND2_X1 U87 ( .A1(\mem[1][4] ), .A2(n682), .ZN(n677) );
  OAI21_X1 U88 ( .B1(n406), .B2(n682), .A(n676), .ZN(n526) );
  NAND2_X1 U89 ( .A1(\mem[1][5] ), .A2(n682), .ZN(n676) );
  OAI21_X1 U90 ( .B1(n405), .B2(n682), .A(n675), .ZN(n525) );
  NAND2_X1 U91 ( .A1(\mem[1][6] ), .A2(n682), .ZN(n675) );
  OAI21_X1 U92 ( .B1(n404), .B2(n682), .A(n674), .ZN(n524) );
  NAND2_X1 U93 ( .A1(\mem[1][7] ), .A2(n682), .ZN(n674) );
  OAI21_X1 U94 ( .B1(n411), .B2(n653), .A(n652), .ZN(n507) );
  NAND2_X1 U95 ( .A1(\mem[4][0] ), .A2(n653), .ZN(n652) );
  OAI21_X1 U96 ( .B1(n410), .B2(n653), .A(n651), .ZN(n506) );
  NAND2_X1 U97 ( .A1(\mem[4][1] ), .A2(n653), .ZN(n651) );
  OAI21_X1 U98 ( .B1(n409), .B2(n653), .A(n650), .ZN(n505) );
  NAND2_X1 U99 ( .A1(\mem[4][2] ), .A2(n653), .ZN(n650) );
  OAI21_X1 U100 ( .B1(n408), .B2(n653), .A(n649), .ZN(n504) );
  NAND2_X1 U101 ( .A1(\mem[4][3] ), .A2(n653), .ZN(n649) );
  OAI21_X1 U102 ( .B1(n407), .B2(n653), .A(n648), .ZN(n503) );
  NAND2_X1 U103 ( .A1(\mem[4][4] ), .A2(n653), .ZN(n648) );
  OAI21_X1 U104 ( .B1(n406), .B2(n653), .A(n647), .ZN(n502) );
  NAND2_X1 U105 ( .A1(\mem[4][5] ), .A2(n653), .ZN(n647) );
  OAI21_X1 U106 ( .B1(n405), .B2(n653), .A(n646), .ZN(n501) );
  NAND2_X1 U107 ( .A1(\mem[4][6] ), .A2(n653), .ZN(n646) );
  OAI21_X1 U108 ( .B1(n404), .B2(n653), .A(n645), .ZN(n500) );
  NAND2_X1 U109 ( .A1(\mem[4][7] ), .A2(n653), .ZN(n645) );
  OAI21_X1 U110 ( .B1(n411), .B2(n643), .A(n642), .ZN(n499) );
  NAND2_X1 U111 ( .A1(\mem[5][0] ), .A2(n643), .ZN(n642) );
  OAI21_X1 U112 ( .B1(n410), .B2(n643), .A(n641), .ZN(n498) );
  NAND2_X1 U113 ( .A1(\mem[5][1] ), .A2(n643), .ZN(n641) );
  OAI21_X1 U114 ( .B1(n409), .B2(n643), .A(n640), .ZN(n497) );
  NAND2_X1 U115 ( .A1(\mem[5][2] ), .A2(n643), .ZN(n640) );
  OAI21_X1 U116 ( .B1(n408), .B2(n643), .A(n639), .ZN(n496) );
  NAND2_X1 U117 ( .A1(\mem[5][3] ), .A2(n643), .ZN(n639) );
  OAI21_X1 U118 ( .B1(n407), .B2(n643), .A(n638), .ZN(n495) );
  NAND2_X1 U119 ( .A1(\mem[5][4] ), .A2(n643), .ZN(n638) );
  OAI21_X1 U120 ( .B1(n406), .B2(n643), .A(n637), .ZN(n494) );
  NAND2_X1 U121 ( .A1(\mem[5][5] ), .A2(n643), .ZN(n637) );
  OAI21_X1 U122 ( .B1(n405), .B2(n643), .A(n636), .ZN(n493) );
  NAND2_X1 U123 ( .A1(\mem[5][6] ), .A2(n643), .ZN(n636) );
  OAI21_X1 U124 ( .B1(n404), .B2(n643), .A(n635), .ZN(n492) );
  NAND2_X1 U125 ( .A1(\mem[5][7] ), .A2(n643), .ZN(n635) );
  OAI21_X1 U126 ( .B1(n411), .B2(n634), .A(n633), .ZN(n491) );
  NAND2_X1 U127 ( .A1(\mem[6][0] ), .A2(n634), .ZN(n633) );
  OAI21_X1 U128 ( .B1(n410), .B2(n634), .A(n632), .ZN(n490) );
  NAND2_X1 U129 ( .A1(\mem[6][1] ), .A2(n634), .ZN(n632) );
  OAI21_X1 U130 ( .B1(n409), .B2(n634), .A(n631), .ZN(n489) );
  NAND2_X1 U131 ( .A1(\mem[6][2] ), .A2(n634), .ZN(n631) );
  OAI21_X1 U132 ( .B1(n408), .B2(n634), .A(n630), .ZN(n488) );
  NAND2_X1 U133 ( .A1(\mem[6][3] ), .A2(n634), .ZN(n630) );
  OAI21_X1 U134 ( .B1(n407), .B2(n634), .A(n629), .ZN(n487) );
  NAND2_X1 U135 ( .A1(\mem[6][4] ), .A2(n634), .ZN(n629) );
  OAI21_X1 U136 ( .B1(n406), .B2(n634), .A(n628), .ZN(n486) );
  NAND2_X1 U137 ( .A1(\mem[6][5] ), .A2(n634), .ZN(n628) );
  OAI21_X1 U138 ( .B1(n405), .B2(n634), .A(n627), .ZN(n485) );
  NAND2_X1 U139 ( .A1(\mem[6][6] ), .A2(n634), .ZN(n627) );
  OAI21_X1 U140 ( .B1(n404), .B2(n634), .A(n626), .ZN(n484) );
  NAND2_X1 U141 ( .A1(\mem[6][7] ), .A2(n634), .ZN(n626) );
  OAI21_X1 U142 ( .B1(n411), .B2(n623), .A(n622), .ZN(n483) );
  NAND2_X1 U143 ( .A1(\mem[7][0] ), .A2(n623), .ZN(n622) );
  OAI21_X1 U144 ( .B1(n410), .B2(n623), .A(n621), .ZN(n482) );
  NAND2_X1 U145 ( .A1(\mem[7][1] ), .A2(n623), .ZN(n621) );
  OAI21_X1 U146 ( .B1(n409), .B2(n623), .A(n620), .ZN(n481) );
  NAND2_X1 U147 ( .A1(\mem[7][2] ), .A2(n623), .ZN(n620) );
  OAI21_X1 U148 ( .B1(n408), .B2(n623), .A(n619), .ZN(n480) );
  NAND2_X1 U149 ( .A1(\mem[7][3] ), .A2(n623), .ZN(n619) );
  OAI21_X1 U150 ( .B1(n407), .B2(n623), .A(n618), .ZN(n479) );
  NAND2_X1 U151 ( .A1(\mem[7][4] ), .A2(n623), .ZN(n618) );
  OAI21_X1 U152 ( .B1(n406), .B2(n623), .A(n617), .ZN(n478) );
  NAND2_X1 U153 ( .A1(\mem[7][5] ), .A2(n623), .ZN(n617) );
  OAI21_X1 U154 ( .B1(n405), .B2(n623), .A(n616), .ZN(n477) );
  NAND2_X1 U155 ( .A1(\mem[7][6] ), .A2(n623), .ZN(n616) );
  OAI21_X1 U156 ( .B1(n404), .B2(n623), .A(n615), .ZN(n476) );
  NAND2_X1 U157 ( .A1(\mem[7][7] ), .A2(n623), .ZN(n615) );
  OAI21_X1 U158 ( .B1(n411), .B2(n614), .A(n613), .ZN(n475) );
  NAND2_X1 U159 ( .A1(\mem[8][0] ), .A2(n614), .ZN(n613) );
  OAI21_X1 U160 ( .B1(n410), .B2(n614), .A(n612), .ZN(n474) );
  NAND2_X1 U161 ( .A1(\mem[8][1] ), .A2(n614), .ZN(n612) );
  OAI21_X1 U162 ( .B1(n409), .B2(n614), .A(n611), .ZN(n473) );
  NAND2_X1 U163 ( .A1(\mem[8][2] ), .A2(n614), .ZN(n611) );
  OAI21_X1 U164 ( .B1(n408), .B2(n614), .A(n610), .ZN(n472) );
  NAND2_X1 U165 ( .A1(\mem[8][3] ), .A2(n614), .ZN(n610) );
  OAI21_X1 U166 ( .B1(n407), .B2(n614), .A(n609), .ZN(n471) );
  NAND2_X1 U167 ( .A1(\mem[8][4] ), .A2(n614), .ZN(n609) );
  OAI21_X1 U168 ( .B1(n406), .B2(n614), .A(n608), .ZN(n470) );
  NAND2_X1 U169 ( .A1(\mem[8][5] ), .A2(n614), .ZN(n608) );
  OAI21_X1 U170 ( .B1(n405), .B2(n614), .A(n607), .ZN(n469) );
  NAND2_X1 U171 ( .A1(\mem[8][6] ), .A2(n614), .ZN(n607) );
  OAI21_X1 U172 ( .B1(n404), .B2(n614), .A(n606), .ZN(n468) );
  NAND2_X1 U173 ( .A1(\mem[8][7] ), .A2(n614), .ZN(n606) );
  OAI21_X1 U174 ( .B1(n411), .B2(n604), .A(n603), .ZN(n467) );
  NAND2_X1 U175 ( .A1(\mem[9][0] ), .A2(n604), .ZN(n603) );
  OAI21_X1 U176 ( .B1(n410), .B2(n604), .A(n602), .ZN(n466) );
  NAND2_X1 U177 ( .A1(\mem[9][1] ), .A2(n604), .ZN(n602) );
  OAI21_X1 U178 ( .B1(n409), .B2(n604), .A(n601), .ZN(n465) );
  NAND2_X1 U179 ( .A1(\mem[9][2] ), .A2(n604), .ZN(n601) );
  OAI21_X1 U180 ( .B1(n408), .B2(n604), .A(n600), .ZN(n464) );
  NAND2_X1 U181 ( .A1(\mem[9][3] ), .A2(n604), .ZN(n600) );
  OAI21_X1 U182 ( .B1(n407), .B2(n604), .A(n599), .ZN(n463) );
  NAND2_X1 U183 ( .A1(\mem[9][4] ), .A2(n604), .ZN(n599) );
  OAI21_X1 U184 ( .B1(n406), .B2(n604), .A(n598), .ZN(n462) );
  NAND2_X1 U185 ( .A1(\mem[9][5] ), .A2(n604), .ZN(n598) );
  OAI21_X1 U186 ( .B1(n405), .B2(n604), .A(n597), .ZN(n461) );
  NAND2_X1 U187 ( .A1(\mem[9][6] ), .A2(n604), .ZN(n597) );
  OAI21_X1 U188 ( .B1(n404), .B2(n604), .A(n596), .ZN(n460) );
  NAND2_X1 U189 ( .A1(\mem[9][7] ), .A2(n604), .ZN(n596) );
  OAI21_X1 U190 ( .B1(n411), .B2(n594), .A(n593), .ZN(n459) );
  NAND2_X1 U191 ( .A1(\mem[10][0] ), .A2(n594), .ZN(n593) );
  OAI21_X1 U192 ( .B1(n410), .B2(n594), .A(n592), .ZN(n458) );
  NAND2_X1 U193 ( .A1(\mem[10][1] ), .A2(n594), .ZN(n592) );
  OAI21_X1 U194 ( .B1(n409), .B2(n594), .A(n591), .ZN(n457) );
  NAND2_X1 U195 ( .A1(\mem[10][2] ), .A2(n594), .ZN(n591) );
  OAI21_X1 U196 ( .B1(n408), .B2(n594), .A(n590), .ZN(n456) );
  NAND2_X1 U197 ( .A1(\mem[10][3] ), .A2(n594), .ZN(n590) );
  OAI21_X1 U198 ( .B1(n407), .B2(n594), .A(n589), .ZN(n455) );
  NAND2_X1 U199 ( .A1(\mem[10][4] ), .A2(n594), .ZN(n589) );
  OAI21_X1 U200 ( .B1(n406), .B2(n594), .A(n588), .ZN(n454) );
  NAND2_X1 U201 ( .A1(\mem[10][5] ), .A2(n594), .ZN(n588) );
  OAI21_X1 U202 ( .B1(n405), .B2(n594), .A(n587), .ZN(n453) );
  NAND2_X1 U203 ( .A1(\mem[10][6] ), .A2(n594), .ZN(n587) );
  OAI21_X1 U204 ( .B1(n404), .B2(n594), .A(n586), .ZN(n452) );
  NAND2_X1 U205 ( .A1(\mem[10][7] ), .A2(n594), .ZN(n586) );
  OAI21_X1 U206 ( .B1(n411), .B2(n585), .A(n584), .ZN(n451) );
  NAND2_X1 U207 ( .A1(\mem[11][0] ), .A2(n585), .ZN(n584) );
  OAI21_X1 U208 ( .B1(n410), .B2(n585), .A(n583), .ZN(n450) );
  NAND2_X1 U209 ( .A1(\mem[11][1] ), .A2(n585), .ZN(n583) );
  OAI21_X1 U210 ( .B1(n409), .B2(n585), .A(n582), .ZN(n449) );
  NAND2_X1 U211 ( .A1(\mem[11][2] ), .A2(n585), .ZN(n582) );
  OAI21_X1 U212 ( .B1(n408), .B2(n585), .A(n581), .ZN(n448) );
  NAND2_X1 U213 ( .A1(\mem[11][3] ), .A2(n585), .ZN(n581) );
  OAI21_X1 U214 ( .B1(n407), .B2(n585), .A(n580), .ZN(n447) );
  NAND2_X1 U215 ( .A1(\mem[11][4] ), .A2(n585), .ZN(n580) );
  OAI21_X1 U216 ( .B1(n406), .B2(n585), .A(n579), .ZN(n446) );
  NAND2_X1 U217 ( .A1(\mem[11][5] ), .A2(n585), .ZN(n579) );
  OAI21_X1 U218 ( .B1(n405), .B2(n585), .A(n578), .ZN(n445) );
  NAND2_X1 U219 ( .A1(\mem[11][6] ), .A2(n585), .ZN(n578) );
  OAI21_X1 U220 ( .B1(n404), .B2(n585), .A(n577), .ZN(n444) );
  NAND2_X1 U221 ( .A1(\mem[11][7] ), .A2(n585), .ZN(n577) );
  OAI21_X1 U222 ( .B1(n411), .B2(n576), .A(n575), .ZN(n443) );
  NAND2_X1 U223 ( .A1(\mem[12][0] ), .A2(n576), .ZN(n575) );
  OAI21_X1 U224 ( .B1(n410), .B2(n576), .A(n574), .ZN(n442) );
  NAND2_X1 U225 ( .A1(\mem[12][1] ), .A2(n576), .ZN(n574) );
  OAI21_X1 U226 ( .B1(n409), .B2(n576), .A(n573), .ZN(n441) );
  NAND2_X1 U227 ( .A1(\mem[12][2] ), .A2(n576), .ZN(n573) );
  OAI21_X1 U228 ( .B1(n408), .B2(n576), .A(n572), .ZN(n440) );
  NAND2_X1 U229 ( .A1(\mem[12][3] ), .A2(n576), .ZN(n572) );
  OAI21_X1 U230 ( .B1(n407), .B2(n576), .A(n571), .ZN(n439) );
  NAND2_X1 U231 ( .A1(\mem[12][4] ), .A2(n576), .ZN(n571) );
  OAI21_X1 U232 ( .B1(n406), .B2(n576), .A(n570), .ZN(n438) );
  NAND2_X1 U233 ( .A1(\mem[12][5] ), .A2(n576), .ZN(n570) );
  OAI21_X1 U234 ( .B1(n405), .B2(n576), .A(n569), .ZN(n437) );
  NAND2_X1 U235 ( .A1(\mem[12][6] ), .A2(n576), .ZN(n569) );
  OAI21_X1 U236 ( .B1(n404), .B2(n576), .A(n568), .ZN(n436) );
  NAND2_X1 U237 ( .A1(\mem[12][7] ), .A2(n576), .ZN(n568) );
  OAI21_X1 U238 ( .B1(n411), .B2(n567), .A(n566), .ZN(n435) );
  NAND2_X1 U239 ( .A1(\mem[13][0] ), .A2(n567), .ZN(n566) );
  OAI21_X1 U240 ( .B1(n410), .B2(n567), .A(n565), .ZN(n434) );
  NAND2_X1 U241 ( .A1(\mem[13][1] ), .A2(n567), .ZN(n565) );
  OAI21_X1 U242 ( .B1(n409), .B2(n567), .A(n564), .ZN(n433) );
  NAND2_X1 U243 ( .A1(\mem[13][2] ), .A2(n567), .ZN(n564) );
  OAI21_X1 U244 ( .B1(n408), .B2(n567), .A(n563), .ZN(n432) );
  NAND2_X1 U245 ( .A1(\mem[13][3] ), .A2(n567), .ZN(n563) );
  OAI21_X1 U246 ( .B1(n407), .B2(n567), .A(n562), .ZN(n431) );
  NAND2_X1 U247 ( .A1(\mem[13][4] ), .A2(n567), .ZN(n562) );
  OAI21_X1 U248 ( .B1(n406), .B2(n567), .A(n561), .ZN(n430) );
  NAND2_X1 U249 ( .A1(\mem[13][5] ), .A2(n567), .ZN(n561) );
  OAI21_X1 U250 ( .B1(n405), .B2(n567), .A(n560), .ZN(n429) );
  NAND2_X1 U251 ( .A1(\mem[13][6] ), .A2(n567), .ZN(n560) );
  OAI21_X1 U252 ( .B1(n404), .B2(n567), .A(n559), .ZN(n428) );
  NAND2_X1 U253 ( .A1(\mem[13][7] ), .A2(n567), .ZN(n559) );
  OAI21_X1 U254 ( .B1(n411), .B2(n558), .A(n557), .ZN(n427) );
  NAND2_X1 U255 ( .A1(\mem[14][0] ), .A2(n558), .ZN(n557) );
  OAI21_X1 U256 ( .B1(n410), .B2(n558), .A(n556), .ZN(n426) );
  NAND2_X1 U257 ( .A1(\mem[14][1] ), .A2(n558), .ZN(n556) );
  OAI21_X1 U258 ( .B1(n409), .B2(n558), .A(n555), .ZN(n425) );
  NAND2_X1 U259 ( .A1(\mem[14][2] ), .A2(n558), .ZN(n555) );
  OAI21_X1 U260 ( .B1(n408), .B2(n558), .A(n554), .ZN(n424) );
  NAND2_X1 U261 ( .A1(\mem[14][3] ), .A2(n558), .ZN(n554) );
  OAI21_X1 U262 ( .B1(n407), .B2(n558), .A(n553), .ZN(n423) );
  NAND2_X1 U263 ( .A1(\mem[14][4] ), .A2(n558), .ZN(n553) );
  OAI21_X1 U264 ( .B1(n406), .B2(n558), .A(n552), .ZN(n422) );
  NAND2_X1 U265 ( .A1(\mem[14][5] ), .A2(n558), .ZN(n552) );
  OAI21_X1 U266 ( .B1(n405), .B2(n558), .A(n551), .ZN(n421) );
  NAND2_X1 U267 ( .A1(\mem[14][6] ), .A2(n558), .ZN(n551) );
  OAI21_X1 U268 ( .B1(n404), .B2(n558), .A(n550), .ZN(n420) );
  NAND2_X1 U269 ( .A1(\mem[14][7] ), .A2(n558), .ZN(n550) );
  OAI21_X1 U270 ( .B1(n411), .B2(n548), .A(n547), .ZN(n419) );
  NAND2_X1 U271 ( .A1(\mem[15][0] ), .A2(n548), .ZN(n547) );
  OAI21_X1 U272 ( .B1(n410), .B2(n548), .A(n546), .ZN(n418) );
  NAND2_X1 U273 ( .A1(\mem[15][1] ), .A2(n548), .ZN(n546) );
  OAI21_X1 U274 ( .B1(n409), .B2(n548), .A(n545), .ZN(n417) );
  NAND2_X1 U275 ( .A1(\mem[15][2] ), .A2(n548), .ZN(n545) );
  OAI21_X1 U276 ( .B1(n408), .B2(n548), .A(n544), .ZN(n416) );
  NAND2_X1 U277 ( .A1(\mem[15][3] ), .A2(n548), .ZN(n544) );
  OAI21_X1 U278 ( .B1(n407), .B2(n548), .A(n543), .ZN(n415) );
  NAND2_X1 U279 ( .A1(\mem[15][4] ), .A2(n548), .ZN(n543) );
  OAI21_X1 U280 ( .B1(n406), .B2(n548), .A(n542), .ZN(n414) );
  NAND2_X1 U281 ( .A1(\mem[15][5] ), .A2(n548), .ZN(n542) );
  OAI21_X1 U282 ( .B1(n405), .B2(n548), .A(n541), .ZN(n413) );
  NAND2_X1 U283 ( .A1(\mem[15][6] ), .A2(n548), .ZN(n541) );
  OAI21_X1 U284 ( .B1(n404), .B2(n548), .A(n540), .ZN(n412) );
  NAND2_X1 U285 ( .A1(\mem[15][7] ), .A2(n548), .ZN(n540) );
  AND2_X1 U286 ( .A1(N13), .A2(wr_en), .ZN(n549) );
  NOR2_X1 U287 ( .A1(N11), .A2(N12), .ZN(n684) );
  NOR2_X1 U288 ( .A1(n402), .A2(N12), .ZN(n663) );
  AND2_X1 U289 ( .A1(N12), .A2(n402), .ZN(n644) );
  AND2_X1 U290 ( .A1(N12), .A2(N11), .ZN(n625) );
  INV_X1 U291 ( .A(data_in[0]), .ZN(n411) );
  INV_X1 U292 ( .A(data_in[1]), .ZN(n410) );
  INV_X1 U293 ( .A(data_in[2]), .ZN(n409) );
  INV_X1 U294 ( .A(data_in[3]), .ZN(n408) );
  INV_X1 U295 ( .A(data_in[4]), .ZN(n407) );
  INV_X1 U296 ( .A(data_in[5]), .ZN(n406) );
  INV_X1 U297 ( .A(data_in[6]), .ZN(n405) );
  INV_X1 U298 ( .A(data_in[7]), .ZN(n404) );
  MUX2_X1 U299 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n400), .Z(n3) );
  MUX2_X1 U300 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(N10), .Z(n4) );
  MUX2_X1 U301 ( .A(n4), .B(n3), .S(n397), .Z(n5) );
  MUX2_X1 U302 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n399), .Z(n6) );
  MUX2_X1 U303 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n398), .Z(n7) );
  MUX2_X1 U304 ( .A(n7), .B(n6), .S(N11), .Z(n8) );
  MUX2_X1 U305 ( .A(n8), .B(n5), .S(N12), .Z(n9) );
  MUX2_X1 U306 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n398), .Z(n10) );
  MUX2_X1 U307 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n398), .Z(n11) );
  MUX2_X1 U308 ( .A(n11), .B(n10), .S(N11), .Z(n294) );
  MUX2_X1 U309 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n398), .Z(n295) );
  MUX2_X1 U310 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n398), .Z(n296) );
  MUX2_X1 U311 ( .A(n296), .B(n295), .S(N11), .Z(n297) );
  MUX2_X1 U312 ( .A(n297), .B(n294), .S(N12), .Z(n298) );
  MUX2_X1 U313 ( .A(n298), .B(n9), .S(N13), .Z(N21) );
  MUX2_X1 U314 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n398), .Z(n299) );
  MUX2_X1 U315 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n398), .Z(n300) );
  MUX2_X1 U316 ( .A(n300), .B(n299), .S(N11), .Z(n301) );
  MUX2_X1 U317 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n398), .Z(n302) );
  MUX2_X1 U318 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n398), .Z(n303) );
  MUX2_X1 U319 ( .A(n303), .B(n302), .S(N11), .Z(n304) );
  MUX2_X1 U320 ( .A(n304), .B(n301), .S(N12), .Z(n305) );
  MUX2_X1 U321 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n398), .Z(n306) );
  MUX2_X1 U322 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n398), .Z(n307) );
  MUX2_X1 U323 ( .A(n307), .B(n306), .S(N11), .Z(n308) );
  MUX2_X1 U324 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n398), .Z(n309) );
  MUX2_X1 U325 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n398), .Z(n310) );
  MUX2_X1 U326 ( .A(n310), .B(n309), .S(N11), .Z(n311) );
  MUX2_X1 U327 ( .A(n311), .B(n308), .S(N12), .Z(n312) );
  MUX2_X1 U328 ( .A(n312), .B(n305), .S(N13), .Z(N20) );
  MUX2_X1 U329 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n399), .Z(n313) );
  MUX2_X1 U330 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n399), .Z(n314) );
  MUX2_X1 U331 ( .A(n314), .B(n313), .S(n397), .Z(n315) );
  MUX2_X1 U332 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n399), .Z(n316) );
  MUX2_X1 U333 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n399), .Z(n317) );
  MUX2_X1 U334 ( .A(n317), .B(n316), .S(n397), .Z(n318) );
  MUX2_X1 U335 ( .A(n318), .B(n315), .S(N12), .Z(n319) );
  MUX2_X1 U336 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n399), .Z(n320) );
  MUX2_X1 U337 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n399), .Z(n321) );
  MUX2_X1 U338 ( .A(n321), .B(n320), .S(n397), .Z(n322) );
  MUX2_X1 U339 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n399), .Z(n323) );
  MUX2_X1 U340 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n399), .Z(n324) );
  MUX2_X1 U341 ( .A(n324), .B(n323), .S(n397), .Z(n325) );
  MUX2_X1 U342 ( .A(n325), .B(n322), .S(N12), .Z(n326) );
  MUX2_X1 U343 ( .A(n326), .B(n319), .S(N13), .Z(N19) );
  MUX2_X1 U344 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n399), .Z(n327) );
  MUX2_X1 U345 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n399), .Z(n328) );
  MUX2_X1 U346 ( .A(n328), .B(n327), .S(n397), .Z(n329) );
  MUX2_X1 U347 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n399), .Z(n330) );
  MUX2_X1 U348 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n399), .Z(n331) );
  MUX2_X1 U349 ( .A(n331), .B(n330), .S(n397), .Z(n332) );
  MUX2_X1 U350 ( .A(n332), .B(n329), .S(N12), .Z(n333) );
  MUX2_X1 U351 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n400), .Z(n334) );
  MUX2_X1 U352 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n400), .Z(n335) );
  MUX2_X1 U353 ( .A(n335), .B(n334), .S(n397), .Z(n336) );
  MUX2_X1 U354 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n400), .Z(n337) );
  MUX2_X1 U355 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n400), .Z(n338) );
  MUX2_X1 U356 ( .A(n338), .B(n337), .S(n397), .Z(n339) );
  MUX2_X1 U357 ( .A(n339), .B(n336), .S(N12), .Z(n340) );
  MUX2_X1 U358 ( .A(n340), .B(n333), .S(N13), .Z(N18) );
  MUX2_X1 U359 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n400), .Z(n341) );
  MUX2_X1 U360 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n400), .Z(n342) );
  MUX2_X1 U361 ( .A(n342), .B(n341), .S(n397), .Z(n343) );
  MUX2_X1 U362 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n400), .Z(n344) );
  MUX2_X1 U363 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n400), .Z(n345) );
  MUX2_X1 U364 ( .A(n345), .B(n344), .S(n397), .Z(n346) );
  MUX2_X1 U365 ( .A(n346), .B(n343), .S(N12), .Z(n347) );
  MUX2_X1 U366 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n400), .Z(n348) );
  MUX2_X1 U367 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n400), .Z(n349) );
  MUX2_X1 U368 ( .A(n349), .B(n348), .S(n397), .Z(n350) );
  MUX2_X1 U369 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n400), .Z(n351) );
  MUX2_X1 U370 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n400), .Z(n352) );
  MUX2_X1 U371 ( .A(n352), .B(n351), .S(n397), .Z(n353) );
  MUX2_X1 U372 ( .A(n353), .B(n350), .S(N12), .Z(n354) );
  MUX2_X1 U373 ( .A(n354), .B(n347), .S(N13), .Z(N17) );
  MUX2_X1 U374 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(N10), .Z(n355) );
  MUX2_X1 U375 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(N10), .Z(n356) );
  MUX2_X1 U376 ( .A(n356), .B(n355), .S(N11), .Z(n357) );
  MUX2_X1 U377 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(N10), .Z(n358) );
  MUX2_X1 U378 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n399), .Z(n359) );
  MUX2_X1 U379 ( .A(n359), .B(n358), .S(N11), .Z(n360) );
  MUX2_X1 U380 ( .A(n360), .B(n357), .S(N12), .Z(n361) );
  MUX2_X1 U381 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(N10), .Z(n362) );
  MUX2_X1 U382 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n400), .Z(n363) );
  MUX2_X1 U383 ( .A(n363), .B(n362), .S(N11), .Z(n364) );
  MUX2_X1 U384 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n398), .Z(n365) );
  MUX2_X1 U385 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n399), .Z(n366) );
  MUX2_X1 U386 ( .A(n366), .B(n365), .S(N11), .Z(n367) );
  MUX2_X1 U387 ( .A(n367), .B(n364), .S(N12), .Z(n368) );
  MUX2_X1 U388 ( .A(n368), .B(n361), .S(N13), .Z(N16) );
  MUX2_X1 U389 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n400), .Z(n369) );
  MUX2_X1 U390 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n400), .Z(n370) );
  MUX2_X1 U391 ( .A(n370), .B(n369), .S(N11), .Z(n371) );
  MUX2_X1 U392 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n399), .Z(n372) );
  MUX2_X1 U393 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n398), .Z(n373) );
  MUX2_X1 U394 ( .A(n373), .B(n372), .S(N11), .Z(n374) );
  MUX2_X1 U395 ( .A(n374), .B(n371), .S(N12), .Z(n375) );
  MUX2_X1 U396 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n376) );
  MUX2_X1 U397 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n377) );
  MUX2_X1 U398 ( .A(n377), .B(n376), .S(N11), .Z(n378) );
  MUX2_X1 U399 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n379) );
  MUX2_X1 U400 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n380) );
  MUX2_X1 U401 ( .A(n380), .B(n379), .S(N11), .Z(n381) );
  MUX2_X1 U402 ( .A(n381), .B(n378), .S(N12), .Z(n382) );
  MUX2_X1 U403 ( .A(n382), .B(n375), .S(N13), .Z(N15) );
  MUX2_X1 U404 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n398), .Z(n383) );
  MUX2_X1 U405 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n384) );
  MUX2_X1 U406 ( .A(n384), .B(n383), .S(N11), .Z(n385) );
  MUX2_X1 U407 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(N10), .Z(n386) );
  MUX2_X1 U408 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n387) );
  MUX2_X1 U409 ( .A(n387), .B(n386), .S(N11), .Z(n388) );
  MUX2_X1 U410 ( .A(n388), .B(n385), .S(N12), .Z(n389) );
  MUX2_X1 U411 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n390) );
  MUX2_X1 U412 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n391) );
  MUX2_X1 U413 ( .A(n391), .B(n390), .S(N11), .Z(n392) );
  MUX2_X1 U414 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n393) );
  MUX2_X1 U415 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n394) );
  MUX2_X1 U416 ( .A(n394), .B(n393), .S(n397), .Z(n395) );
  MUX2_X1 U417 ( .A(n395), .B(n392), .S(N12), .Z(n396) );
  MUX2_X1 U418 ( .A(n396), .B(n389), .S(N13), .Z(N14) );
  INV_X1 U419 ( .A(N10), .ZN(n401) );
  INV_X1 U420 ( .A(N11), .ZN(n402) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_13 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, N19, N20, N21, n2, n4, n5, n6, n7, n8, n9, n10,
         n11, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N16), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n413), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n414), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n415), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n416), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n417), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n418), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n419), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n420), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n421), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n422), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n423), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n424), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n425), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n426), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n427), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n428), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n429), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n430), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n431), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n432), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n433), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n434), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n435), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n436), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n437), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n438), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n439), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n440), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n441), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n442), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n443), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n444), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n445), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n446), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n447), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n448), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n449), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n450), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n451), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n452), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n453), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n454), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n455), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n456), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n457), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n458), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n459), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n460), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n461), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n462), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n463), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n464), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n465), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n466), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n467), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n468), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n469), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n470), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n471), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n472), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n473), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n474), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n475), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n476), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n477), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n478), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n479), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n480), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n481), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n482), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n483), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n484), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n485), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n486), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n487), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n488), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n489), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n490), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n491), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n492), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n493), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n494), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n495), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n496), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n497), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n498), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n499), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n500), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n501), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n502), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n503), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n504), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n505), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n506), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n507), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n508), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n509), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n510), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n511), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n512), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n513), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n514), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n515), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n516), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n517), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n518), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n519), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n520), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n521), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n522), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n523), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n524), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n525), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n526), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n527), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n528), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n529), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n530), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n531), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n532), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n533), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n534), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n535), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n536), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n537), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n538), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n539), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n540), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N20), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .QN(n2) );
  INV_X2 U3 ( .A(n2), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(N10), .Z(n399) );
  BUF_X1 U5 ( .A(N10), .Z(n400) );
  BUF_X1 U6 ( .A(N10), .Z(n401) );
  BUF_X1 U7 ( .A(N11), .Z(n398) );
  NAND2_X1 U8 ( .A1(n664), .A2(n684), .ZN(n673) );
  NAND2_X1 U9 ( .A1(n664), .A2(n674), .ZN(n663) );
  NAND2_X1 U10 ( .A1(n685), .A2(n684), .ZN(n694) );
  NAND2_X1 U11 ( .A1(n674), .A2(n685), .ZN(n683) );
  NAND2_X1 U12 ( .A1(n606), .A2(n685), .ZN(n615) );
  NAND2_X1 U13 ( .A1(n596), .A2(n685), .ZN(n605) );
  NAND2_X1 U14 ( .A1(n606), .A2(n664), .ZN(n595) );
  NAND2_X1 U15 ( .A1(n596), .A2(n664), .ZN(n586) );
  NAND2_X1 U16 ( .A1(n645), .A2(n684), .ZN(n654) );
  NAND2_X1 U17 ( .A1(n645), .A2(n674), .ZN(n644) );
  NAND2_X1 U18 ( .A1(n626), .A2(n684), .ZN(n635) );
  NAND2_X1 U19 ( .A1(n626), .A2(n674), .ZN(n624) );
  NAND2_X1 U20 ( .A1(n606), .A2(n645), .ZN(n577) );
  NAND2_X1 U21 ( .A1(n596), .A2(n645), .ZN(n568) );
  NAND2_X1 U22 ( .A1(n606), .A2(n626), .ZN(n559) );
  NAND2_X1 U23 ( .A1(n596), .A2(n626), .ZN(n549) );
  AND2_X1 U24 ( .A1(n550), .A2(N10), .ZN(n596) );
  AND2_X1 U25 ( .A1(n550), .A2(n402), .ZN(n606) );
  AND2_X1 U26 ( .A1(N10), .A2(n625), .ZN(n674) );
  AND2_X1 U27 ( .A1(n625), .A2(n402), .ZN(n684) );
  OAI21_X1 U28 ( .B1(n694), .B2(n412), .A(n693), .ZN(n540) );
  NAND2_X1 U29 ( .A1(\mem[0][0] ), .A2(n694), .ZN(n693) );
  OAI21_X1 U30 ( .B1(n694), .B2(n411), .A(n692), .ZN(n539) );
  NAND2_X1 U31 ( .A1(\mem[0][1] ), .A2(n694), .ZN(n692) );
  OAI21_X1 U32 ( .B1(n694), .B2(n410), .A(n691), .ZN(n538) );
  NAND2_X1 U33 ( .A1(\mem[0][2] ), .A2(n694), .ZN(n691) );
  OAI21_X1 U34 ( .B1(n694), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U35 ( .A1(\mem[0][3] ), .A2(n694), .ZN(n690) );
  OAI21_X1 U36 ( .B1(n694), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U37 ( .A1(\mem[0][4] ), .A2(n694), .ZN(n689) );
  OAI21_X1 U38 ( .B1(n694), .B2(n407), .A(n688), .ZN(n535) );
  NAND2_X1 U39 ( .A1(\mem[0][5] ), .A2(n694), .ZN(n688) );
  OAI21_X1 U40 ( .B1(n694), .B2(n406), .A(n687), .ZN(n534) );
  NAND2_X1 U41 ( .A1(\mem[0][6] ), .A2(n694), .ZN(n687) );
  OAI21_X1 U42 ( .B1(n694), .B2(n405), .A(n686), .ZN(n533) );
  NAND2_X1 U43 ( .A1(\mem[0][7] ), .A2(n694), .ZN(n686) );
  OAI21_X1 U44 ( .B1(n412), .B2(n673), .A(n672), .ZN(n524) );
  NAND2_X1 U45 ( .A1(\mem[2][0] ), .A2(n673), .ZN(n672) );
  OAI21_X1 U46 ( .B1(n411), .B2(n673), .A(n671), .ZN(n523) );
  NAND2_X1 U47 ( .A1(\mem[2][1] ), .A2(n673), .ZN(n671) );
  OAI21_X1 U48 ( .B1(n410), .B2(n673), .A(n670), .ZN(n522) );
  NAND2_X1 U49 ( .A1(\mem[2][2] ), .A2(n673), .ZN(n670) );
  OAI21_X1 U50 ( .B1(n409), .B2(n673), .A(n669), .ZN(n521) );
  NAND2_X1 U51 ( .A1(\mem[2][3] ), .A2(n673), .ZN(n669) );
  OAI21_X1 U52 ( .B1(n408), .B2(n673), .A(n668), .ZN(n520) );
  NAND2_X1 U53 ( .A1(\mem[2][4] ), .A2(n673), .ZN(n668) );
  OAI21_X1 U54 ( .B1(n407), .B2(n673), .A(n667), .ZN(n519) );
  NAND2_X1 U55 ( .A1(\mem[2][5] ), .A2(n673), .ZN(n667) );
  OAI21_X1 U56 ( .B1(n406), .B2(n673), .A(n666), .ZN(n518) );
  NAND2_X1 U57 ( .A1(\mem[2][6] ), .A2(n673), .ZN(n666) );
  OAI21_X1 U58 ( .B1(n405), .B2(n673), .A(n665), .ZN(n517) );
  NAND2_X1 U59 ( .A1(\mem[2][7] ), .A2(n673), .ZN(n665) );
  OAI21_X1 U60 ( .B1(n412), .B2(n663), .A(n662), .ZN(n516) );
  NAND2_X1 U61 ( .A1(\mem[3][0] ), .A2(n663), .ZN(n662) );
  OAI21_X1 U62 ( .B1(n411), .B2(n663), .A(n661), .ZN(n515) );
  NAND2_X1 U63 ( .A1(\mem[3][1] ), .A2(n663), .ZN(n661) );
  OAI21_X1 U64 ( .B1(n410), .B2(n663), .A(n660), .ZN(n514) );
  NAND2_X1 U65 ( .A1(\mem[3][2] ), .A2(n663), .ZN(n660) );
  OAI21_X1 U66 ( .B1(n409), .B2(n663), .A(n659), .ZN(n513) );
  NAND2_X1 U67 ( .A1(\mem[3][3] ), .A2(n663), .ZN(n659) );
  OAI21_X1 U68 ( .B1(n408), .B2(n663), .A(n658), .ZN(n512) );
  NAND2_X1 U69 ( .A1(\mem[3][4] ), .A2(n663), .ZN(n658) );
  OAI21_X1 U70 ( .B1(n407), .B2(n663), .A(n657), .ZN(n511) );
  NAND2_X1 U71 ( .A1(\mem[3][5] ), .A2(n663), .ZN(n657) );
  OAI21_X1 U72 ( .B1(n406), .B2(n663), .A(n656), .ZN(n510) );
  NAND2_X1 U73 ( .A1(\mem[3][6] ), .A2(n663), .ZN(n656) );
  OAI21_X1 U74 ( .B1(n405), .B2(n663), .A(n655), .ZN(n509) );
  NAND2_X1 U75 ( .A1(\mem[3][7] ), .A2(n663), .ZN(n655) );
  NOR2_X1 U76 ( .A1(n404), .A2(N13), .ZN(n625) );
  INV_X1 U77 ( .A(wr_en), .ZN(n404) );
  OAI21_X1 U78 ( .B1(n412), .B2(n683), .A(n682), .ZN(n532) );
  NAND2_X1 U79 ( .A1(\mem[1][0] ), .A2(n683), .ZN(n682) );
  OAI21_X1 U80 ( .B1(n411), .B2(n683), .A(n681), .ZN(n531) );
  NAND2_X1 U81 ( .A1(\mem[1][1] ), .A2(n683), .ZN(n681) );
  OAI21_X1 U82 ( .B1(n410), .B2(n683), .A(n680), .ZN(n530) );
  NAND2_X1 U83 ( .A1(\mem[1][2] ), .A2(n683), .ZN(n680) );
  OAI21_X1 U84 ( .B1(n409), .B2(n683), .A(n679), .ZN(n529) );
  NAND2_X1 U85 ( .A1(\mem[1][3] ), .A2(n683), .ZN(n679) );
  OAI21_X1 U86 ( .B1(n408), .B2(n683), .A(n678), .ZN(n528) );
  NAND2_X1 U87 ( .A1(\mem[1][4] ), .A2(n683), .ZN(n678) );
  OAI21_X1 U88 ( .B1(n407), .B2(n683), .A(n677), .ZN(n527) );
  NAND2_X1 U89 ( .A1(\mem[1][5] ), .A2(n683), .ZN(n677) );
  OAI21_X1 U90 ( .B1(n406), .B2(n683), .A(n676), .ZN(n526) );
  NAND2_X1 U91 ( .A1(\mem[1][6] ), .A2(n683), .ZN(n676) );
  OAI21_X1 U92 ( .B1(n405), .B2(n683), .A(n675), .ZN(n525) );
  NAND2_X1 U93 ( .A1(\mem[1][7] ), .A2(n683), .ZN(n675) );
  OAI21_X1 U94 ( .B1(n412), .B2(n654), .A(n653), .ZN(n508) );
  NAND2_X1 U95 ( .A1(\mem[4][0] ), .A2(n654), .ZN(n653) );
  OAI21_X1 U96 ( .B1(n411), .B2(n654), .A(n652), .ZN(n507) );
  NAND2_X1 U97 ( .A1(\mem[4][1] ), .A2(n654), .ZN(n652) );
  OAI21_X1 U98 ( .B1(n410), .B2(n654), .A(n651), .ZN(n506) );
  NAND2_X1 U99 ( .A1(\mem[4][2] ), .A2(n654), .ZN(n651) );
  OAI21_X1 U100 ( .B1(n409), .B2(n654), .A(n650), .ZN(n505) );
  NAND2_X1 U101 ( .A1(\mem[4][3] ), .A2(n654), .ZN(n650) );
  OAI21_X1 U102 ( .B1(n408), .B2(n654), .A(n649), .ZN(n504) );
  NAND2_X1 U103 ( .A1(\mem[4][4] ), .A2(n654), .ZN(n649) );
  OAI21_X1 U104 ( .B1(n407), .B2(n654), .A(n648), .ZN(n503) );
  NAND2_X1 U105 ( .A1(\mem[4][5] ), .A2(n654), .ZN(n648) );
  OAI21_X1 U106 ( .B1(n406), .B2(n654), .A(n647), .ZN(n502) );
  NAND2_X1 U107 ( .A1(\mem[4][6] ), .A2(n654), .ZN(n647) );
  OAI21_X1 U108 ( .B1(n405), .B2(n654), .A(n646), .ZN(n501) );
  NAND2_X1 U109 ( .A1(\mem[4][7] ), .A2(n654), .ZN(n646) );
  OAI21_X1 U110 ( .B1(n412), .B2(n644), .A(n643), .ZN(n500) );
  NAND2_X1 U111 ( .A1(\mem[5][0] ), .A2(n644), .ZN(n643) );
  OAI21_X1 U112 ( .B1(n411), .B2(n644), .A(n642), .ZN(n499) );
  NAND2_X1 U113 ( .A1(\mem[5][1] ), .A2(n644), .ZN(n642) );
  OAI21_X1 U114 ( .B1(n410), .B2(n644), .A(n641), .ZN(n498) );
  NAND2_X1 U115 ( .A1(\mem[5][2] ), .A2(n644), .ZN(n641) );
  OAI21_X1 U116 ( .B1(n409), .B2(n644), .A(n640), .ZN(n497) );
  NAND2_X1 U117 ( .A1(\mem[5][3] ), .A2(n644), .ZN(n640) );
  OAI21_X1 U118 ( .B1(n408), .B2(n644), .A(n639), .ZN(n496) );
  NAND2_X1 U119 ( .A1(\mem[5][4] ), .A2(n644), .ZN(n639) );
  OAI21_X1 U120 ( .B1(n407), .B2(n644), .A(n638), .ZN(n495) );
  NAND2_X1 U121 ( .A1(\mem[5][5] ), .A2(n644), .ZN(n638) );
  OAI21_X1 U122 ( .B1(n406), .B2(n644), .A(n637), .ZN(n494) );
  NAND2_X1 U123 ( .A1(\mem[5][6] ), .A2(n644), .ZN(n637) );
  OAI21_X1 U124 ( .B1(n405), .B2(n644), .A(n636), .ZN(n493) );
  NAND2_X1 U125 ( .A1(\mem[5][7] ), .A2(n644), .ZN(n636) );
  OAI21_X1 U126 ( .B1(n412), .B2(n635), .A(n634), .ZN(n492) );
  NAND2_X1 U127 ( .A1(\mem[6][0] ), .A2(n635), .ZN(n634) );
  OAI21_X1 U128 ( .B1(n411), .B2(n635), .A(n633), .ZN(n491) );
  NAND2_X1 U129 ( .A1(\mem[6][1] ), .A2(n635), .ZN(n633) );
  OAI21_X1 U130 ( .B1(n410), .B2(n635), .A(n632), .ZN(n490) );
  NAND2_X1 U131 ( .A1(\mem[6][2] ), .A2(n635), .ZN(n632) );
  OAI21_X1 U132 ( .B1(n409), .B2(n635), .A(n631), .ZN(n489) );
  NAND2_X1 U133 ( .A1(\mem[6][3] ), .A2(n635), .ZN(n631) );
  OAI21_X1 U134 ( .B1(n408), .B2(n635), .A(n630), .ZN(n488) );
  NAND2_X1 U135 ( .A1(\mem[6][4] ), .A2(n635), .ZN(n630) );
  OAI21_X1 U136 ( .B1(n407), .B2(n635), .A(n629), .ZN(n487) );
  NAND2_X1 U137 ( .A1(\mem[6][5] ), .A2(n635), .ZN(n629) );
  OAI21_X1 U138 ( .B1(n406), .B2(n635), .A(n628), .ZN(n486) );
  NAND2_X1 U139 ( .A1(\mem[6][6] ), .A2(n635), .ZN(n628) );
  OAI21_X1 U140 ( .B1(n405), .B2(n635), .A(n627), .ZN(n485) );
  NAND2_X1 U141 ( .A1(\mem[6][7] ), .A2(n635), .ZN(n627) );
  OAI21_X1 U142 ( .B1(n412), .B2(n624), .A(n623), .ZN(n484) );
  NAND2_X1 U143 ( .A1(\mem[7][0] ), .A2(n624), .ZN(n623) );
  OAI21_X1 U144 ( .B1(n411), .B2(n624), .A(n622), .ZN(n483) );
  NAND2_X1 U145 ( .A1(\mem[7][1] ), .A2(n624), .ZN(n622) );
  OAI21_X1 U146 ( .B1(n410), .B2(n624), .A(n621), .ZN(n482) );
  NAND2_X1 U147 ( .A1(\mem[7][2] ), .A2(n624), .ZN(n621) );
  OAI21_X1 U148 ( .B1(n409), .B2(n624), .A(n620), .ZN(n481) );
  NAND2_X1 U149 ( .A1(\mem[7][3] ), .A2(n624), .ZN(n620) );
  OAI21_X1 U150 ( .B1(n408), .B2(n624), .A(n619), .ZN(n480) );
  NAND2_X1 U151 ( .A1(\mem[7][4] ), .A2(n624), .ZN(n619) );
  OAI21_X1 U152 ( .B1(n407), .B2(n624), .A(n618), .ZN(n479) );
  NAND2_X1 U153 ( .A1(\mem[7][5] ), .A2(n624), .ZN(n618) );
  OAI21_X1 U154 ( .B1(n406), .B2(n624), .A(n617), .ZN(n478) );
  NAND2_X1 U155 ( .A1(\mem[7][6] ), .A2(n624), .ZN(n617) );
  OAI21_X1 U156 ( .B1(n405), .B2(n624), .A(n616), .ZN(n477) );
  NAND2_X1 U157 ( .A1(\mem[7][7] ), .A2(n624), .ZN(n616) );
  OAI21_X1 U158 ( .B1(n412), .B2(n615), .A(n614), .ZN(n476) );
  NAND2_X1 U159 ( .A1(\mem[8][0] ), .A2(n615), .ZN(n614) );
  OAI21_X1 U160 ( .B1(n411), .B2(n615), .A(n613), .ZN(n475) );
  NAND2_X1 U161 ( .A1(\mem[8][1] ), .A2(n615), .ZN(n613) );
  OAI21_X1 U162 ( .B1(n410), .B2(n615), .A(n612), .ZN(n474) );
  NAND2_X1 U163 ( .A1(\mem[8][2] ), .A2(n615), .ZN(n612) );
  OAI21_X1 U164 ( .B1(n409), .B2(n615), .A(n611), .ZN(n473) );
  NAND2_X1 U165 ( .A1(\mem[8][3] ), .A2(n615), .ZN(n611) );
  OAI21_X1 U166 ( .B1(n408), .B2(n615), .A(n610), .ZN(n472) );
  NAND2_X1 U167 ( .A1(\mem[8][4] ), .A2(n615), .ZN(n610) );
  OAI21_X1 U168 ( .B1(n407), .B2(n615), .A(n609), .ZN(n471) );
  NAND2_X1 U169 ( .A1(\mem[8][5] ), .A2(n615), .ZN(n609) );
  OAI21_X1 U170 ( .B1(n406), .B2(n615), .A(n608), .ZN(n470) );
  NAND2_X1 U171 ( .A1(\mem[8][6] ), .A2(n615), .ZN(n608) );
  OAI21_X1 U172 ( .B1(n405), .B2(n615), .A(n607), .ZN(n469) );
  NAND2_X1 U173 ( .A1(\mem[8][7] ), .A2(n615), .ZN(n607) );
  OAI21_X1 U174 ( .B1(n412), .B2(n605), .A(n604), .ZN(n468) );
  NAND2_X1 U175 ( .A1(\mem[9][0] ), .A2(n605), .ZN(n604) );
  OAI21_X1 U176 ( .B1(n411), .B2(n605), .A(n603), .ZN(n467) );
  NAND2_X1 U177 ( .A1(\mem[9][1] ), .A2(n605), .ZN(n603) );
  OAI21_X1 U178 ( .B1(n410), .B2(n605), .A(n602), .ZN(n466) );
  NAND2_X1 U179 ( .A1(\mem[9][2] ), .A2(n605), .ZN(n602) );
  OAI21_X1 U180 ( .B1(n409), .B2(n605), .A(n601), .ZN(n465) );
  NAND2_X1 U181 ( .A1(\mem[9][3] ), .A2(n605), .ZN(n601) );
  OAI21_X1 U182 ( .B1(n408), .B2(n605), .A(n600), .ZN(n464) );
  NAND2_X1 U183 ( .A1(\mem[9][4] ), .A2(n605), .ZN(n600) );
  OAI21_X1 U184 ( .B1(n407), .B2(n605), .A(n599), .ZN(n463) );
  NAND2_X1 U185 ( .A1(\mem[9][5] ), .A2(n605), .ZN(n599) );
  OAI21_X1 U186 ( .B1(n406), .B2(n605), .A(n598), .ZN(n462) );
  NAND2_X1 U187 ( .A1(\mem[9][6] ), .A2(n605), .ZN(n598) );
  OAI21_X1 U188 ( .B1(n405), .B2(n605), .A(n597), .ZN(n461) );
  NAND2_X1 U189 ( .A1(\mem[9][7] ), .A2(n605), .ZN(n597) );
  OAI21_X1 U190 ( .B1(n412), .B2(n595), .A(n594), .ZN(n460) );
  NAND2_X1 U191 ( .A1(\mem[10][0] ), .A2(n595), .ZN(n594) );
  OAI21_X1 U192 ( .B1(n411), .B2(n595), .A(n593), .ZN(n459) );
  NAND2_X1 U193 ( .A1(\mem[10][1] ), .A2(n595), .ZN(n593) );
  OAI21_X1 U194 ( .B1(n410), .B2(n595), .A(n592), .ZN(n458) );
  NAND2_X1 U195 ( .A1(\mem[10][2] ), .A2(n595), .ZN(n592) );
  OAI21_X1 U196 ( .B1(n409), .B2(n595), .A(n591), .ZN(n457) );
  NAND2_X1 U197 ( .A1(\mem[10][3] ), .A2(n595), .ZN(n591) );
  OAI21_X1 U198 ( .B1(n408), .B2(n595), .A(n590), .ZN(n456) );
  NAND2_X1 U199 ( .A1(\mem[10][4] ), .A2(n595), .ZN(n590) );
  OAI21_X1 U200 ( .B1(n407), .B2(n595), .A(n589), .ZN(n455) );
  NAND2_X1 U201 ( .A1(\mem[10][5] ), .A2(n595), .ZN(n589) );
  OAI21_X1 U202 ( .B1(n406), .B2(n595), .A(n588), .ZN(n454) );
  NAND2_X1 U203 ( .A1(\mem[10][6] ), .A2(n595), .ZN(n588) );
  OAI21_X1 U204 ( .B1(n405), .B2(n595), .A(n587), .ZN(n453) );
  NAND2_X1 U205 ( .A1(\mem[10][7] ), .A2(n595), .ZN(n587) );
  OAI21_X1 U206 ( .B1(n412), .B2(n586), .A(n585), .ZN(n452) );
  NAND2_X1 U207 ( .A1(\mem[11][0] ), .A2(n586), .ZN(n585) );
  OAI21_X1 U208 ( .B1(n411), .B2(n586), .A(n584), .ZN(n451) );
  NAND2_X1 U209 ( .A1(\mem[11][1] ), .A2(n586), .ZN(n584) );
  OAI21_X1 U210 ( .B1(n410), .B2(n586), .A(n583), .ZN(n450) );
  NAND2_X1 U211 ( .A1(\mem[11][2] ), .A2(n586), .ZN(n583) );
  OAI21_X1 U212 ( .B1(n409), .B2(n586), .A(n582), .ZN(n449) );
  NAND2_X1 U213 ( .A1(\mem[11][3] ), .A2(n586), .ZN(n582) );
  OAI21_X1 U214 ( .B1(n408), .B2(n586), .A(n581), .ZN(n448) );
  NAND2_X1 U215 ( .A1(\mem[11][4] ), .A2(n586), .ZN(n581) );
  OAI21_X1 U216 ( .B1(n407), .B2(n586), .A(n580), .ZN(n447) );
  NAND2_X1 U217 ( .A1(\mem[11][5] ), .A2(n586), .ZN(n580) );
  OAI21_X1 U218 ( .B1(n406), .B2(n586), .A(n579), .ZN(n446) );
  NAND2_X1 U219 ( .A1(\mem[11][6] ), .A2(n586), .ZN(n579) );
  OAI21_X1 U220 ( .B1(n405), .B2(n586), .A(n578), .ZN(n445) );
  NAND2_X1 U221 ( .A1(\mem[11][7] ), .A2(n586), .ZN(n578) );
  OAI21_X1 U222 ( .B1(n412), .B2(n577), .A(n576), .ZN(n444) );
  NAND2_X1 U223 ( .A1(\mem[12][0] ), .A2(n577), .ZN(n576) );
  OAI21_X1 U224 ( .B1(n411), .B2(n577), .A(n575), .ZN(n443) );
  NAND2_X1 U225 ( .A1(\mem[12][1] ), .A2(n577), .ZN(n575) );
  OAI21_X1 U226 ( .B1(n410), .B2(n577), .A(n574), .ZN(n442) );
  NAND2_X1 U227 ( .A1(\mem[12][2] ), .A2(n577), .ZN(n574) );
  OAI21_X1 U228 ( .B1(n409), .B2(n577), .A(n573), .ZN(n441) );
  NAND2_X1 U229 ( .A1(\mem[12][3] ), .A2(n577), .ZN(n573) );
  OAI21_X1 U230 ( .B1(n408), .B2(n577), .A(n572), .ZN(n440) );
  NAND2_X1 U231 ( .A1(\mem[12][4] ), .A2(n577), .ZN(n572) );
  OAI21_X1 U232 ( .B1(n407), .B2(n577), .A(n571), .ZN(n439) );
  NAND2_X1 U233 ( .A1(\mem[12][5] ), .A2(n577), .ZN(n571) );
  OAI21_X1 U234 ( .B1(n406), .B2(n577), .A(n570), .ZN(n438) );
  NAND2_X1 U235 ( .A1(\mem[12][6] ), .A2(n577), .ZN(n570) );
  OAI21_X1 U236 ( .B1(n405), .B2(n577), .A(n569), .ZN(n437) );
  NAND2_X1 U237 ( .A1(\mem[12][7] ), .A2(n577), .ZN(n569) );
  OAI21_X1 U238 ( .B1(n412), .B2(n568), .A(n567), .ZN(n436) );
  NAND2_X1 U239 ( .A1(\mem[13][0] ), .A2(n568), .ZN(n567) );
  OAI21_X1 U240 ( .B1(n411), .B2(n568), .A(n566), .ZN(n435) );
  NAND2_X1 U241 ( .A1(\mem[13][1] ), .A2(n568), .ZN(n566) );
  OAI21_X1 U242 ( .B1(n410), .B2(n568), .A(n565), .ZN(n434) );
  NAND2_X1 U243 ( .A1(\mem[13][2] ), .A2(n568), .ZN(n565) );
  OAI21_X1 U244 ( .B1(n409), .B2(n568), .A(n564), .ZN(n433) );
  NAND2_X1 U245 ( .A1(\mem[13][3] ), .A2(n568), .ZN(n564) );
  OAI21_X1 U246 ( .B1(n408), .B2(n568), .A(n563), .ZN(n432) );
  NAND2_X1 U247 ( .A1(\mem[13][4] ), .A2(n568), .ZN(n563) );
  OAI21_X1 U248 ( .B1(n407), .B2(n568), .A(n562), .ZN(n431) );
  NAND2_X1 U249 ( .A1(\mem[13][5] ), .A2(n568), .ZN(n562) );
  OAI21_X1 U250 ( .B1(n406), .B2(n568), .A(n561), .ZN(n430) );
  NAND2_X1 U251 ( .A1(\mem[13][6] ), .A2(n568), .ZN(n561) );
  OAI21_X1 U252 ( .B1(n405), .B2(n568), .A(n560), .ZN(n429) );
  NAND2_X1 U253 ( .A1(\mem[13][7] ), .A2(n568), .ZN(n560) );
  OAI21_X1 U254 ( .B1(n412), .B2(n559), .A(n558), .ZN(n428) );
  NAND2_X1 U255 ( .A1(\mem[14][0] ), .A2(n559), .ZN(n558) );
  OAI21_X1 U256 ( .B1(n411), .B2(n559), .A(n557), .ZN(n427) );
  NAND2_X1 U257 ( .A1(\mem[14][1] ), .A2(n559), .ZN(n557) );
  OAI21_X1 U258 ( .B1(n410), .B2(n559), .A(n556), .ZN(n426) );
  NAND2_X1 U259 ( .A1(\mem[14][2] ), .A2(n559), .ZN(n556) );
  OAI21_X1 U260 ( .B1(n409), .B2(n559), .A(n555), .ZN(n425) );
  NAND2_X1 U261 ( .A1(\mem[14][3] ), .A2(n559), .ZN(n555) );
  OAI21_X1 U262 ( .B1(n408), .B2(n559), .A(n554), .ZN(n424) );
  NAND2_X1 U263 ( .A1(\mem[14][4] ), .A2(n559), .ZN(n554) );
  OAI21_X1 U264 ( .B1(n407), .B2(n559), .A(n553), .ZN(n423) );
  NAND2_X1 U265 ( .A1(\mem[14][5] ), .A2(n559), .ZN(n553) );
  OAI21_X1 U266 ( .B1(n406), .B2(n559), .A(n552), .ZN(n422) );
  NAND2_X1 U267 ( .A1(\mem[14][6] ), .A2(n559), .ZN(n552) );
  OAI21_X1 U268 ( .B1(n405), .B2(n559), .A(n551), .ZN(n421) );
  NAND2_X1 U269 ( .A1(\mem[14][7] ), .A2(n559), .ZN(n551) );
  OAI21_X1 U270 ( .B1(n412), .B2(n549), .A(n548), .ZN(n420) );
  NAND2_X1 U271 ( .A1(\mem[15][0] ), .A2(n549), .ZN(n548) );
  OAI21_X1 U272 ( .B1(n411), .B2(n549), .A(n547), .ZN(n419) );
  NAND2_X1 U273 ( .A1(\mem[15][1] ), .A2(n549), .ZN(n547) );
  OAI21_X1 U274 ( .B1(n410), .B2(n549), .A(n546), .ZN(n418) );
  NAND2_X1 U275 ( .A1(\mem[15][2] ), .A2(n549), .ZN(n546) );
  OAI21_X1 U276 ( .B1(n409), .B2(n549), .A(n545), .ZN(n417) );
  NAND2_X1 U277 ( .A1(\mem[15][3] ), .A2(n549), .ZN(n545) );
  OAI21_X1 U278 ( .B1(n408), .B2(n549), .A(n544), .ZN(n416) );
  NAND2_X1 U279 ( .A1(\mem[15][4] ), .A2(n549), .ZN(n544) );
  OAI21_X1 U280 ( .B1(n407), .B2(n549), .A(n543), .ZN(n415) );
  NAND2_X1 U281 ( .A1(\mem[15][5] ), .A2(n549), .ZN(n543) );
  OAI21_X1 U282 ( .B1(n406), .B2(n549), .A(n542), .ZN(n414) );
  NAND2_X1 U283 ( .A1(\mem[15][6] ), .A2(n549), .ZN(n542) );
  OAI21_X1 U284 ( .B1(n405), .B2(n549), .A(n541), .ZN(n413) );
  NAND2_X1 U285 ( .A1(\mem[15][7] ), .A2(n549), .ZN(n541) );
  AND2_X1 U286 ( .A1(N13), .A2(wr_en), .ZN(n550) );
  NOR2_X1 U287 ( .A1(N11), .A2(N12), .ZN(n685) );
  NOR2_X1 U288 ( .A1(n403), .A2(N12), .ZN(n664) );
  AND2_X1 U289 ( .A1(N12), .A2(n403), .ZN(n645) );
  AND2_X1 U290 ( .A1(N12), .A2(N11), .ZN(n626) );
  INV_X1 U291 ( .A(data_in[0]), .ZN(n412) );
  INV_X1 U292 ( .A(data_in[1]), .ZN(n411) );
  INV_X1 U293 ( .A(data_in[2]), .ZN(n410) );
  INV_X1 U294 ( .A(data_in[3]), .ZN(n409) );
  INV_X1 U295 ( .A(data_in[4]), .ZN(n408) );
  INV_X1 U296 ( .A(data_in[5]), .ZN(n407) );
  INV_X1 U297 ( .A(data_in[6]), .ZN(n406) );
  INV_X1 U298 ( .A(data_in[7]), .ZN(n405) );
  MUX2_X1 U299 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(N10), .Z(n4) );
  MUX2_X1 U300 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(N10), .Z(n5) );
  MUX2_X1 U301 ( .A(n5), .B(n4), .S(N11), .Z(n6) );
  MUX2_X1 U302 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(N10), .Z(n7) );
  MUX2_X1 U303 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n8) );
  MUX2_X1 U304 ( .A(n8), .B(n7), .S(N11), .Z(n9) );
  MUX2_X1 U305 ( .A(n9), .B(n6), .S(N12), .Z(n10) );
  MUX2_X1 U306 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n399), .Z(n11) );
  MUX2_X1 U307 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n399), .Z(n294) );
  MUX2_X1 U308 ( .A(n294), .B(n11), .S(N11), .Z(n295) );
  MUX2_X1 U309 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n399), .Z(n296) );
  MUX2_X1 U310 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n399), .Z(n297) );
  MUX2_X1 U311 ( .A(n297), .B(n296), .S(N11), .Z(n298) );
  MUX2_X1 U312 ( .A(n298), .B(n295), .S(N12), .Z(n299) );
  MUX2_X1 U313 ( .A(n299), .B(n10), .S(N13), .Z(N21) );
  MUX2_X1 U314 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n399), .Z(n300) );
  MUX2_X1 U315 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n399), .Z(n301) );
  MUX2_X1 U316 ( .A(n301), .B(n300), .S(N11), .Z(n302) );
  MUX2_X1 U317 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n399), .Z(n303) );
  MUX2_X1 U318 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n399), .Z(n304) );
  MUX2_X1 U319 ( .A(n304), .B(n303), .S(N11), .Z(n305) );
  MUX2_X1 U320 ( .A(n305), .B(n302), .S(N12), .Z(n306) );
  MUX2_X1 U321 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n399), .Z(n307) );
  MUX2_X1 U322 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n399), .Z(n308) );
  MUX2_X1 U323 ( .A(n308), .B(n307), .S(N11), .Z(n309) );
  MUX2_X1 U324 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n399), .Z(n310) );
  MUX2_X1 U325 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n399), .Z(n311) );
  MUX2_X1 U326 ( .A(n311), .B(n310), .S(N11), .Z(n312) );
  MUX2_X1 U327 ( .A(n312), .B(n309), .S(N12), .Z(n313) );
  MUX2_X1 U328 ( .A(n313), .B(n306), .S(N13), .Z(N20) );
  MUX2_X1 U329 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n400), .Z(n314) );
  MUX2_X1 U330 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n400), .Z(n315) );
  MUX2_X1 U331 ( .A(n315), .B(n314), .S(n398), .Z(n316) );
  MUX2_X1 U332 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n400), .Z(n317) );
  MUX2_X1 U333 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n400), .Z(n318) );
  MUX2_X1 U334 ( .A(n318), .B(n317), .S(n398), .Z(n319) );
  MUX2_X1 U335 ( .A(n319), .B(n316), .S(N12), .Z(n320) );
  MUX2_X1 U336 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n400), .Z(n321) );
  MUX2_X1 U337 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n400), .Z(n322) );
  MUX2_X1 U338 ( .A(n322), .B(n321), .S(n398), .Z(n323) );
  MUX2_X1 U339 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n400), .Z(n324) );
  MUX2_X1 U340 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n400), .Z(n325) );
  MUX2_X1 U341 ( .A(n325), .B(n324), .S(n398), .Z(n326) );
  MUX2_X1 U342 ( .A(n326), .B(n323), .S(N12), .Z(n327) );
  MUX2_X1 U343 ( .A(n327), .B(n320), .S(N13), .Z(N19) );
  MUX2_X1 U344 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n400), .Z(n328) );
  MUX2_X1 U345 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n400), .Z(n329) );
  MUX2_X1 U346 ( .A(n329), .B(n328), .S(n398), .Z(n330) );
  MUX2_X1 U347 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n400), .Z(n331) );
  MUX2_X1 U348 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n400), .Z(n332) );
  MUX2_X1 U349 ( .A(n332), .B(n331), .S(n398), .Z(n333) );
  MUX2_X1 U350 ( .A(n333), .B(n330), .S(N12), .Z(n334) );
  MUX2_X1 U351 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n401), .Z(n335) );
  MUX2_X1 U352 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n401), .Z(n336) );
  MUX2_X1 U353 ( .A(n336), .B(n335), .S(n398), .Z(n337) );
  MUX2_X1 U354 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n401), .Z(n338) );
  MUX2_X1 U355 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n401), .Z(n339) );
  MUX2_X1 U356 ( .A(n339), .B(n338), .S(n398), .Z(n340) );
  MUX2_X1 U357 ( .A(n340), .B(n337), .S(N12), .Z(n341) );
  MUX2_X1 U358 ( .A(n341), .B(n334), .S(N13), .Z(N18) );
  MUX2_X1 U359 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n401), .Z(n342) );
  MUX2_X1 U360 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n401), .Z(n343) );
  MUX2_X1 U361 ( .A(n343), .B(n342), .S(n398), .Z(n344) );
  MUX2_X1 U362 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n401), .Z(n345) );
  MUX2_X1 U363 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n401), .Z(n346) );
  MUX2_X1 U364 ( .A(n346), .B(n345), .S(n398), .Z(n347) );
  MUX2_X1 U365 ( .A(n347), .B(n344), .S(N12), .Z(n348) );
  MUX2_X1 U366 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n401), .Z(n349) );
  MUX2_X1 U367 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n401), .Z(n350) );
  MUX2_X1 U368 ( .A(n350), .B(n349), .S(n398), .Z(n351) );
  MUX2_X1 U369 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n401), .Z(n352) );
  MUX2_X1 U370 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n401), .Z(n353) );
  MUX2_X1 U371 ( .A(n353), .B(n352), .S(n398), .Z(n354) );
  MUX2_X1 U372 ( .A(n354), .B(n351), .S(N12), .Z(n355) );
  MUX2_X1 U373 ( .A(n355), .B(n348), .S(N13), .Z(N17) );
  MUX2_X1 U374 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n399), .Z(n356) );
  MUX2_X1 U375 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n400), .Z(n357) );
  MUX2_X1 U376 ( .A(n357), .B(n356), .S(N11), .Z(n358) );
  MUX2_X1 U377 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n400), .Z(n359) );
  MUX2_X1 U378 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n399), .Z(n360) );
  MUX2_X1 U379 ( .A(n360), .B(n359), .S(N11), .Z(n361) );
  MUX2_X1 U380 ( .A(n361), .B(n358), .S(N12), .Z(n362) );
  MUX2_X1 U381 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n399), .Z(n363) );
  MUX2_X1 U382 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n401), .Z(n364) );
  MUX2_X1 U383 ( .A(n364), .B(n363), .S(N11), .Z(n365) );
  MUX2_X1 U384 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n399), .Z(n366) );
  MUX2_X1 U385 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n400), .Z(n367) );
  MUX2_X1 U386 ( .A(n367), .B(n366), .S(n398), .Z(n368) );
  MUX2_X1 U387 ( .A(n368), .B(n365), .S(N12), .Z(n369) );
  MUX2_X1 U388 ( .A(n369), .B(n362), .S(N13), .Z(N16) );
  MUX2_X1 U389 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(N10), .Z(n370) );
  MUX2_X1 U390 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n401), .Z(n371) );
  MUX2_X1 U391 ( .A(n371), .B(n370), .S(N11), .Z(n372) );
  MUX2_X1 U392 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n401), .Z(n373) );
  MUX2_X1 U393 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n400), .Z(n374) );
  MUX2_X1 U394 ( .A(n374), .B(n373), .S(N11), .Z(n375) );
  MUX2_X1 U395 ( .A(n375), .B(n372), .S(N12), .Z(n376) );
  MUX2_X1 U396 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n377) );
  MUX2_X1 U397 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n378) );
  MUX2_X1 U398 ( .A(n378), .B(n377), .S(N11), .Z(n379) );
  MUX2_X1 U399 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n380) );
  MUX2_X1 U400 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n400), .Z(n381) );
  MUX2_X1 U401 ( .A(n381), .B(n380), .S(n398), .Z(n382) );
  MUX2_X1 U402 ( .A(n382), .B(n379), .S(N12), .Z(n383) );
  MUX2_X1 U403 ( .A(n383), .B(n376), .S(N13), .Z(N15) );
  MUX2_X1 U404 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(N10), .Z(n384) );
  MUX2_X1 U405 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n385) );
  MUX2_X1 U406 ( .A(n385), .B(n384), .S(N11), .Z(n386) );
  MUX2_X1 U407 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(N10), .Z(n387) );
  MUX2_X1 U408 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n388) );
  MUX2_X1 U409 ( .A(n388), .B(n387), .S(N11), .Z(n389) );
  MUX2_X1 U410 ( .A(n389), .B(n386), .S(N12), .Z(n390) );
  MUX2_X1 U411 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n391) );
  MUX2_X1 U412 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n392) );
  MUX2_X1 U413 ( .A(n392), .B(n391), .S(N11), .Z(n393) );
  MUX2_X1 U414 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n394) );
  MUX2_X1 U415 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n401), .Z(n395) );
  MUX2_X1 U416 ( .A(n395), .B(n394), .S(n398), .Z(n396) );
  MUX2_X1 U417 ( .A(n396), .B(n393), .S(N12), .Z(n397) );
  MUX2_X1 U418 ( .A(n397), .B(n390), .S(N13), .Z(N14) );
  INV_X1 U419 ( .A(N10), .ZN(n402) );
  INV_X1 U420 ( .A(N11), .ZN(n403) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_12 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, N19, N20, N21, n2, n4, n6, n7, n8, n9, n10, n11,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n415), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n416), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n417), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n418), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n419), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n420), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n421), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n422), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n423), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n424), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n425), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n426), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n427), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n428), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n429), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n430), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n431), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n432), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n433), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n434), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n435), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n436), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n437), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n438), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n439), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n440), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n441), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n442), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n443), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n444), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n445), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n446), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n447), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n448), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n449), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n450), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n451), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n452), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n453), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n454), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n455), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n456), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n457), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n458), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n459), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n460), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n461), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n462), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n463), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n464), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n465), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n466), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n467), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n468), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n469), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n470), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n471), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n472), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n473), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n474), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n475), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n476), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n477), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n478), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n479), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n480), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n481), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n482), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n483), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n484), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n485), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n486), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n487), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n488), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n489), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n490), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n491), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n492), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n493), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n494), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n495), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n496), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n497), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n498), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n499), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n500), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n501), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n502), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n503), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n504), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n505), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n506), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n507), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n508), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n509), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n510), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n511), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n512), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n513), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n514), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n515), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n516), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n517), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n518), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n519), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n520), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n521), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n522), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n523), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n524), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n525), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n526), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n527), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n528), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n529), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n530), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n531), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n532), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n533), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n534), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n535), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n536), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n537), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n538), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n539), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n540), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n541), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n542), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N20), .CK(clk), .QN(n4) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[5]  ( .D(N16), .CK(clk), .QN(n2) );
  INV_X2 U3 ( .A(n2), .ZN(data_out[5]) );
  INV_X2 U4 ( .A(n4), .ZN(data_out[1]) );
  BUF_X1 U5 ( .A(N10), .Z(n401) );
  BUF_X1 U6 ( .A(N10), .Z(n402) );
  BUF_X1 U7 ( .A(N10), .Z(n403) );
  BUF_X1 U8 ( .A(N11), .Z(n400) );
  NAND2_X1 U9 ( .A1(n666), .A2(n686), .ZN(n675) );
  NAND2_X1 U10 ( .A1(n666), .A2(n676), .ZN(n665) );
  NAND2_X1 U11 ( .A1(n687), .A2(n686), .ZN(n696) );
  NAND2_X1 U12 ( .A1(n676), .A2(n687), .ZN(n685) );
  NAND2_X1 U13 ( .A1(n608), .A2(n687), .ZN(n617) );
  NAND2_X1 U14 ( .A1(n598), .A2(n687), .ZN(n607) );
  NAND2_X1 U15 ( .A1(n608), .A2(n666), .ZN(n597) );
  NAND2_X1 U16 ( .A1(n598), .A2(n666), .ZN(n588) );
  NAND2_X1 U17 ( .A1(n647), .A2(n686), .ZN(n656) );
  NAND2_X1 U18 ( .A1(n647), .A2(n676), .ZN(n646) );
  NAND2_X1 U19 ( .A1(n628), .A2(n686), .ZN(n637) );
  NAND2_X1 U20 ( .A1(n628), .A2(n676), .ZN(n626) );
  NAND2_X1 U21 ( .A1(n608), .A2(n647), .ZN(n579) );
  NAND2_X1 U22 ( .A1(n598), .A2(n647), .ZN(n570) );
  NAND2_X1 U23 ( .A1(n608), .A2(n628), .ZN(n561) );
  NAND2_X1 U24 ( .A1(n598), .A2(n628), .ZN(n551) );
  AND2_X1 U25 ( .A1(n552), .A2(N10), .ZN(n598) );
  AND2_X1 U26 ( .A1(n552), .A2(n404), .ZN(n608) );
  AND2_X1 U27 ( .A1(N10), .A2(n627), .ZN(n676) );
  AND2_X1 U28 ( .A1(n627), .A2(n404), .ZN(n686) );
  OAI21_X1 U29 ( .B1(n696), .B2(n414), .A(n695), .ZN(n542) );
  NAND2_X1 U30 ( .A1(\mem[0][0] ), .A2(n696), .ZN(n695) );
  OAI21_X1 U31 ( .B1(n696), .B2(n413), .A(n694), .ZN(n541) );
  NAND2_X1 U32 ( .A1(\mem[0][1] ), .A2(n696), .ZN(n694) );
  OAI21_X1 U33 ( .B1(n696), .B2(n412), .A(n693), .ZN(n540) );
  NAND2_X1 U34 ( .A1(\mem[0][2] ), .A2(n696), .ZN(n693) );
  OAI21_X1 U35 ( .B1(n696), .B2(n411), .A(n692), .ZN(n539) );
  NAND2_X1 U36 ( .A1(\mem[0][3] ), .A2(n696), .ZN(n692) );
  OAI21_X1 U37 ( .B1(n696), .B2(n410), .A(n691), .ZN(n538) );
  NAND2_X1 U38 ( .A1(\mem[0][4] ), .A2(n696), .ZN(n691) );
  OAI21_X1 U39 ( .B1(n696), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U40 ( .A1(\mem[0][5] ), .A2(n696), .ZN(n690) );
  OAI21_X1 U41 ( .B1(n696), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U42 ( .A1(\mem[0][6] ), .A2(n696), .ZN(n689) );
  OAI21_X1 U43 ( .B1(n696), .B2(n407), .A(n688), .ZN(n535) );
  NAND2_X1 U44 ( .A1(\mem[0][7] ), .A2(n696), .ZN(n688) );
  OAI21_X1 U45 ( .B1(n414), .B2(n675), .A(n674), .ZN(n526) );
  NAND2_X1 U46 ( .A1(\mem[2][0] ), .A2(n675), .ZN(n674) );
  OAI21_X1 U47 ( .B1(n413), .B2(n675), .A(n673), .ZN(n525) );
  NAND2_X1 U48 ( .A1(\mem[2][1] ), .A2(n675), .ZN(n673) );
  OAI21_X1 U49 ( .B1(n412), .B2(n675), .A(n672), .ZN(n524) );
  NAND2_X1 U50 ( .A1(\mem[2][2] ), .A2(n675), .ZN(n672) );
  OAI21_X1 U51 ( .B1(n411), .B2(n675), .A(n671), .ZN(n523) );
  NAND2_X1 U52 ( .A1(\mem[2][3] ), .A2(n675), .ZN(n671) );
  OAI21_X1 U53 ( .B1(n410), .B2(n675), .A(n670), .ZN(n522) );
  NAND2_X1 U54 ( .A1(\mem[2][4] ), .A2(n675), .ZN(n670) );
  OAI21_X1 U55 ( .B1(n409), .B2(n675), .A(n669), .ZN(n521) );
  NAND2_X1 U56 ( .A1(\mem[2][5] ), .A2(n675), .ZN(n669) );
  OAI21_X1 U57 ( .B1(n408), .B2(n675), .A(n668), .ZN(n520) );
  NAND2_X1 U58 ( .A1(\mem[2][6] ), .A2(n675), .ZN(n668) );
  OAI21_X1 U59 ( .B1(n407), .B2(n675), .A(n667), .ZN(n519) );
  NAND2_X1 U60 ( .A1(\mem[2][7] ), .A2(n675), .ZN(n667) );
  OAI21_X1 U61 ( .B1(n414), .B2(n665), .A(n664), .ZN(n518) );
  NAND2_X1 U62 ( .A1(\mem[3][0] ), .A2(n665), .ZN(n664) );
  OAI21_X1 U63 ( .B1(n413), .B2(n665), .A(n663), .ZN(n517) );
  NAND2_X1 U64 ( .A1(\mem[3][1] ), .A2(n665), .ZN(n663) );
  OAI21_X1 U65 ( .B1(n412), .B2(n665), .A(n662), .ZN(n516) );
  NAND2_X1 U66 ( .A1(\mem[3][2] ), .A2(n665), .ZN(n662) );
  OAI21_X1 U67 ( .B1(n411), .B2(n665), .A(n661), .ZN(n515) );
  NAND2_X1 U68 ( .A1(\mem[3][3] ), .A2(n665), .ZN(n661) );
  OAI21_X1 U69 ( .B1(n410), .B2(n665), .A(n660), .ZN(n514) );
  NAND2_X1 U70 ( .A1(\mem[3][4] ), .A2(n665), .ZN(n660) );
  OAI21_X1 U71 ( .B1(n409), .B2(n665), .A(n659), .ZN(n513) );
  NAND2_X1 U72 ( .A1(\mem[3][5] ), .A2(n665), .ZN(n659) );
  OAI21_X1 U73 ( .B1(n408), .B2(n665), .A(n658), .ZN(n512) );
  NAND2_X1 U74 ( .A1(\mem[3][6] ), .A2(n665), .ZN(n658) );
  OAI21_X1 U75 ( .B1(n407), .B2(n665), .A(n657), .ZN(n511) );
  NAND2_X1 U76 ( .A1(\mem[3][7] ), .A2(n665), .ZN(n657) );
  NOR2_X1 U77 ( .A1(n406), .A2(N13), .ZN(n627) );
  INV_X1 U78 ( .A(wr_en), .ZN(n406) );
  OAI21_X1 U79 ( .B1(n414), .B2(n685), .A(n684), .ZN(n534) );
  NAND2_X1 U80 ( .A1(\mem[1][0] ), .A2(n685), .ZN(n684) );
  OAI21_X1 U81 ( .B1(n413), .B2(n685), .A(n683), .ZN(n533) );
  NAND2_X1 U82 ( .A1(\mem[1][1] ), .A2(n685), .ZN(n683) );
  OAI21_X1 U83 ( .B1(n412), .B2(n685), .A(n682), .ZN(n532) );
  NAND2_X1 U84 ( .A1(\mem[1][2] ), .A2(n685), .ZN(n682) );
  OAI21_X1 U85 ( .B1(n411), .B2(n685), .A(n681), .ZN(n531) );
  NAND2_X1 U86 ( .A1(\mem[1][3] ), .A2(n685), .ZN(n681) );
  OAI21_X1 U87 ( .B1(n410), .B2(n685), .A(n680), .ZN(n530) );
  NAND2_X1 U88 ( .A1(\mem[1][4] ), .A2(n685), .ZN(n680) );
  OAI21_X1 U89 ( .B1(n409), .B2(n685), .A(n679), .ZN(n529) );
  NAND2_X1 U90 ( .A1(\mem[1][5] ), .A2(n685), .ZN(n679) );
  OAI21_X1 U91 ( .B1(n408), .B2(n685), .A(n678), .ZN(n528) );
  NAND2_X1 U92 ( .A1(\mem[1][6] ), .A2(n685), .ZN(n678) );
  OAI21_X1 U93 ( .B1(n407), .B2(n685), .A(n677), .ZN(n527) );
  NAND2_X1 U94 ( .A1(\mem[1][7] ), .A2(n685), .ZN(n677) );
  OAI21_X1 U95 ( .B1(n414), .B2(n656), .A(n655), .ZN(n510) );
  NAND2_X1 U96 ( .A1(\mem[4][0] ), .A2(n656), .ZN(n655) );
  OAI21_X1 U97 ( .B1(n413), .B2(n656), .A(n654), .ZN(n509) );
  NAND2_X1 U98 ( .A1(\mem[4][1] ), .A2(n656), .ZN(n654) );
  OAI21_X1 U99 ( .B1(n412), .B2(n656), .A(n653), .ZN(n508) );
  NAND2_X1 U100 ( .A1(\mem[4][2] ), .A2(n656), .ZN(n653) );
  OAI21_X1 U101 ( .B1(n411), .B2(n656), .A(n652), .ZN(n507) );
  NAND2_X1 U102 ( .A1(\mem[4][3] ), .A2(n656), .ZN(n652) );
  OAI21_X1 U103 ( .B1(n410), .B2(n656), .A(n651), .ZN(n506) );
  NAND2_X1 U104 ( .A1(\mem[4][4] ), .A2(n656), .ZN(n651) );
  OAI21_X1 U105 ( .B1(n409), .B2(n656), .A(n650), .ZN(n505) );
  NAND2_X1 U106 ( .A1(\mem[4][5] ), .A2(n656), .ZN(n650) );
  OAI21_X1 U107 ( .B1(n408), .B2(n656), .A(n649), .ZN(n504) );
  NAND2_X1 U108 ( .A1(\mem[4][6] ), .A2(n656), .ZN(n649) );
  OAI21_X1 U109 ( .B1(n407), .B2(n656), .A(n648), .ZN(n503) );
  NAND2_X1 U110 ( .A1(\mem[4][7] ), .A2(n656), .ZN(n648) );
  OAI21_X1 U111 ( .B1(n414), .B2(n646), .A(n645), .ZN(n502) );
  NAND2_X1 U112 ( .A1(\mem[5][0] ), .A2(n646), .ZN(n645) );
  OAI21_X1 U113 ( .B1(n413), .B2(n646), .A(n644), .ZN(n501) );
  NAND2_X1 U114 ( .A1(\mem[5][1] ), .A2(n646), .ZN(n644) );
  OAI21_X1 U115 ( .B1(n412), .B2(n646), .A(n643), .ZN(n500) );
  NAND2_X1 U116 ( .A1(\mem[5][2] ), .A2(n646), .ZN(n643) );
  OAI21_X1 U117 ( .B1(n411), .B2(n646), .A(n642), .ZN(n499) );
  NAND2_X1 U118 ( .A1(\mem[5][3] ), .A2(n646), .ZN(n642) );
  OAI21_X1 U119 ( .B1(n410), .B2(n646), .A(n641), .ZN(n498) );
  NAND2_X1 U120 ( .A1(\mem[5][4] ), .A2(n646), .ZN(n641) );
  OAI21_X1 U121 ( .B1(n409), .B2(n646), .A(n640), .ZN(n497) );
  NAND2_X1 U122 ( .A1(\mem[5][5] ), .A2(n646), .ZN(n640) );
  OAI21_X1 U123 ( .B1(n408), .B2(n646), .A(n639), .ZN(n496) );
  NAND2_X1 U124 ( .A1(\mem[5][6] ), .A2(n646), .ZN(n639) );
  OAI21_X1 U125 ( .B1(n407), .B2(n646), .A(n638), .ZN(n495) );
  NAND2_X1 U126 ( .A1(\mem[5][7] ), .A2(n646), .ZN(n638) );
  OAI21_X1 U127 ( .B1(n414), .B2(n637), .A(n636), .ZN(n494) );
  NAND2_X1 U128 ( .A1(\mem[6][0] ), .A2(n637), .ZN(n636) );
  OAI21_X1 U129 ( .B1(n413), .B2(n637), .A(n635), .ZN(n493) );
  NAND2_X1 U130 ( .A1(\mem[6][1] ), .A2(n637), .ZN(n635) );
  OAI21_X1 U131 ( .B1(n412), .B2(n637), .A(n634), .ZN(n492) );
  NAND2_X1 U132 ( .A1(\mem[6][2] ), .A2(n637), .ZN(n634) );
  OAI21_X1 U133 ( .B1(n411), .B2(n637), .A(n633), .ZN(n491) );
  NAND2_X1 U134 ( .A1(\mem[6][3] ), .A2(n637), .ZN(n633) );
  OAI21_X1 U135 ( .B1(n410), .B2(n637), .A(n632), .ZN(n490) );
  NAND2_X1 U136 ( .A1(\mem[6][4] ), .A2(n637), .ZN(n632) );
  OAI21_X1 U137 ( .B1(n409), .B2(n637), .A(n631), .ZN(n489) );
  NAND2_X1 U138 ( .A1(\mem[6][5] ), .A2(n637), .ZN(n631) );
  OAI21_X1 U139 ( .B1(n408), .B2(n637), .A(n630), .ZN(n488) );
  NAND2_X1 U140 ( .A1(\mem[6][6] ), .A2(n637), .ZN(n630) );
  OAI21_X1 U141 ( .B1(n407), .B2(n637), .A(n629), .ZN(n487) );
  NAND2_X1 U142 ( .A1(\mem[6][7] ), .A2(n637), .ZN(n629) );
  OAI21_X1 U143 ( .B1(n414), .B2(n626), .A(n625), .ZN(n486) );
  NAND2_X1 U144 ( .A1(\mem[7][0] ), .A2(n626), .ZN(n625) );
  OAI21_X1 U145 ( .B1(n413), .B2(n626), .A(n624), .ZN(n485) );
  NAND2_X1 U146 ( .A1(\mem[7][1] ), .A2(n626), .ZN(n624) );
  OAI21_X1 U147 ( .B1(n412), .B2(n626), .A(n623), .ZN(n484) );
  NAND2_X1 U148 ( .A1(\mem[7][2] ), .A2(n626), .ZN(n623) );
  OAI21_X1 U149 ( .B1(n411), .B2(n626), .A(n622), .ZN(n483) );
  NAND2_X1 U150 ( .A1(\mem[7][3] ), .A2(n626), .ZN(n622) );
  OAI21_X1 U151 ( .B1(n410), .B2(n626), .A(n621), .ZN(n482) );
  NAND2_X1 U152 ( .A1(\mem[7][4] ), .A2(n626), .ZN(n621) );
  OAI21_X1 U153 ( .B1(n409), .B2(n626), .A(n620), .ZN(n481) );
  NAND2_X1 U154 ( .A1(\mem[7][5] ), .A2(n626), .ZN(n620) );
  OAI21_X1 U155 ( .B1(n408), .B2(n626), .A(n619), .ZN(n480) );
  NAND2_X1 U156 ( .A1(\mem[7][6] ), .A2(n626), .ZN(n619) );
  OAI21_X1 U157 ( .B1(n407), .B2(n626), .A(n618), .ZN(n479) );
  NAND2_X1 U158 ( .A1(\mem[7][7] ), .A2(n626), .ZN(n618) );
  OAI21_X1 U159 ( .B1(n414), .B2(n617), .A(n616), .ZN(n478) );
  NAND2_X1 U160 ( .A1(\mem[8][0] ), .A2(n617), .ZN(n616) );
  OAI21_X1 U161 ( .B1(n413), .B2(n617), .A(n615), .ZN(n477) );
  NAND2_X1 U162 ( .A1(\mem[8][1] ), .A2(n617), .ZN(n615) );
  OAI21_X1 U163 ( .B1(n412), .B2(n617), .A(n614), .ZN(n476) );
  NAND2_X1 U164 ( .A1(\mem[8][2] ), .A2(n617), .ZN(n614) );
  OAI21_X1 U165 ( .B1(n411), .B2(n617), .A(n613), .ZN(n475) );
  NAND2_X1 U166 ( .A1(\mem[8][3] ), .A2(n617), .ZN(n613) );
  OAI21_X1 U167 ( .B1(n410), .B2(n617), .A(n612), .ZN(n474) );
  NAND2_X1 U168 ( .A1(\mem[8][4] ), .A2(n617), .ZN(n612) );
  OAI21_X1 U169 ( .B1(n409), .B2(n617), .A(n611), .ZN(n473) );
  NAND2_X1 U170 ( .A1(\mem[8][5] ), .A2(n617), .ZN(n611) );
  OAI21_X1 U171 ( .B1(n408), .B2(n617), .A(n610), .ZN(n472) );
  NAND2_X1 U172 ( .A1(\mem[8][6] ), .A2(n617), .ZN(n610) );
  OAI21_X1 U173 ( .B1(n407), .B2(n617), .A(n609), .ZN(n471) );
  NAND2_X1 U174 ( .A1(\mem[8][7] ), .A2(n617), .ZN(n609) );
  OAI21_X1 U175 ( .B1(n414), .B2(n607), .A(n606), .ZN(n470) );
  NAND2_X1 U176 ( .A1(\mem[9][0] ), .A2(n607), .ZN(n606) );
  OAI21_X1 U177 ( .B1(n413), .B2(n607), .A(n605), .ZN(n469) );
  NAND2_X1 U178 ( .A1(\mem[9][1] ), .A2(n607), .ZN(n605) );
  OAI21_X1 U179 ( .B1(n412), .B2(n607), .A(n604), .ZN(n468) );
  NAND2_X1 U180 ( .A1(\mem[9][2] ), .A2(n607), .ZN(n604) );
  OAI21_X1 U181 ( .B1(n411), .B2(n607), .A(n603), .ZN(n467) );
  NAND2_X1 U182 ( .A1(\mem[9][3] ), .A2(n607), .ZN(n603) );
  OAI21_X1 U183 ( .B1(n410), .B2(n607), .A(n602), .ZN(n466) );
  NAND2_X1 U184 ( .A1(\mem[9][4] ), .A2(n607), .ZN(n602) );
  OAI21_X1 U185 ( .B1(n409), .B2(n607), .A(n601), .ZN(n465) );
  NAND2_X1 U186 ( .A1(\mem[9][5] ), .A2(n607), .ZN(n601) );
  OAI21_X1 U187 ( .B1(n408), .B2(n607), .A(n600), .ZN(n464) );
  NAND2_X1 U188 ( .A1(\mem[9][6] ), .A2(n607), .ZN(n600) );
  OAI21_X1 U189 ( .B1(n407), .B2(n607), .A(n599), .ZN(n463) );
  NAND2_X1 U190 ( .A1(\mem[9][7] ), .A2(n607), .ZN(n599) );
  OAI21_X1 U191 ( .B1(n414), .B2(n597), .A(n596), .ZN(n462) );
  NAND2_X1 U192 ( .A1(\mem[10][0] ), .A2(n597), .ZN(n596) );
  OAI21_X1 U193 ( .B1(n413), .B2(n597), .A(n595), .ZN(n461) );
  NAND2_X1 U194 ( .A1(\mem[10][1] ), .A2(n597), .ZN(n595) );
  OAI21_X1 U195 ( .B1(n412), .B2(n597), .A(n594), .ZN(n460) );
  NAND2_X1 U196 ( .A1(\mem[10][2] ), .A2(n597), .ZN(n594) );
  OAI21_X1 U197 ( .B1(n411), .B2(n597), .A(n593), .ZN(n459) );
  NAND2_X1 U198 ( .A1(\mem[10][3] ), .A2(n597), .ZN(n593) );
  OAI21_X1 U199 ( .B1(n410), .B2(n597), .A(n592), .ZN(n458) );
  NAND2_X1 U200 ( .A1(\mem[10][4] ), .A2(n597), .ZN(n592) );
  OAI21_X1 U201 ( .B1(n409), .B2(n597), .A(n591), .ZN(n457) );
  NAND2_X1 U202 ( .A1(\mem[10][5] ), .A2(n597), .ZN(n591) );
  OAI21_X1 U203 ( .B1(n408), .B2(n597), .A(n590), .ZN(n456) );
  NAND2_X1 U204 ( .A1(\mem[10][6] ), .A2(n597), .ZN(n590) );
  OAI21_X1 U205 ( .B1(n407), .B2(n597), .A(n589), .ZN(n455) );
  NAND2_X1 U206 ( .A1(\mem[10][7] ), .A2(n597), .ZN(n589) );
  OAI21_X1 U207 ( .B1(n414), .B2(n588), .A(n587), .ZN(n454) );
  NAND2_X1 U208 ( .A1(\mem[11][0] ), .A2(n588), .ZN(n587) );
  OAI21_X1 U209 ( .B1(n413), .B2(n588), .A(n586), .ZN(n453) );
  NAND2_X1 U210 ( .A1(\mem[11][1] ), .A2(n588), .ZN(n586) );
  OAI21_X1 U211 ( .B1(n412), .B2(n588), .A(n585), .ZN(n452) );
  NAND2_X1 U212 ( .A1(\mem[11][2] ), .A2(n588), .ZN(n585) );
  OAI21_X1 U213 ( .B1(n411), .B2(n588), .A(n584), .ZN(n451) );
  NAND2_X1 U214 ( .A1(\mem[11][3] ), .A2(n588), .ZN(n584) );
  OAI21_X1 U215 ( .B1(n410), .B2(n588), .A(n583), .ZN(n450) );
  NAND2_X1 U216 ( .A1(\mem[11][4] ), .A2(n588), .ZN(n583) );
  OAI21_X1 U217 ( .B1(n409), .B2(n588), .A(n582), .ZN(n449) );
  NAND2_X1 U218 ( .A1(\mem[11][5] ), .A2(n588), .ZN(n582) );
  OAI21_X1 U219 ( .B1(n408), .B2(n588), .A(n581), .ZN(n448) );
  NAND2_X1 U220 ( .A1(\mem[11][6] ), .A2(n588), .ZN(n581) );
  OAI21_X1 U221 ( .B1(n407), .B2(n588), .A(n580), .ZN(n447) );
  NAND2_X1 U222 ( .A1(\mem[11][7] ), .A2(n588), .ZN(n580) );
  OAI21_X1 U223 ( .B1(n414), .B2(n579), .A(n578), .ZN(n446) );
  NAND2_X1 U224 ( .A1(\mem[12][0] ), .A2(n579), .ZN(n578) );
  OAI21_X1 U225 ( .B1(n413), .B2(n579), .A(n577), .ZN(n445) );
  NAND2_X1 U226 ( .A1(\mem[12][1] ), .A2(n579), .ZN(n577) );
  OAI21_X1 U227 ( .B1(n412), .B2(n579), .A(n576), .ZN(n444) );
  NAND2_X1 U228 ( .A1(\mem[12][2] ), .A2(n579), .ZN(n576) );
  OAI21_X1 U229 ( .B1(n411), .B2(n579), .A(n575), .ZN(n443) );
  NAND2_X1 U230 ( .A1(\mem[12][3] ), .A2(n579), .ZN(n575) );
  OAI21_X1 U231 ( .B1(n410), .B2(n579), .A(n574), .ZN(n442) );
  NAND2_X1 U232 ( .A1(\mem[12][4] ), .A2(n579), .ZN(n574) );
  OAI21_X1 U233 ( .B1(n409), .B2(n579), .A(n573), .ZN(n441) );
  NAND2_X1 U234 ( .A1(\mem[12][5] ), .A2(n579), .ZN(n573) );
  OAI21_X1 U235 ( .B1(n408), .B2(n579), .A(n572), .ZN(n440) );
  NAND2_X1 U236 ( .A1(\mem[12][6] ), .A2(n579), .ZN(n572) );
  OAI21_X1 U237 ( .B1(n407), .B2(n579), .A(n571), .ZN(n439) );
  NAND2_X1 U238 ( .A1(\mem[12][7] ), .A2(n579), .ZN(n571) );
  OAI21_X1 U239 ( .B1(n414), .B2(n570), .A(n569), .ZN(n438) );
  NAND2_X1 U240 ( .A1(\mem[13][0] ), .A2(n570), .ZN(n569) );
  OAI21_X1 U241 ( .B1(n413), .B2(n570), .A(n568), .ZN(n437) );
  NAND2_X1 U242 ( .A1(\mem[13][1] ), .A2(n570), .ZN(n568) );
  OAI21_X1 U243 ( .B1(n412), .B2(n570), .A(n567), .ZN(n436) );
  NAND2_X1 U244 ( .A1(\mem[13][2] ), .A2(n570), .ZN(n567) );
  OAI21_X1 U245 ( .B1(n411), .B2(n570), .A(n566), .ZN(n435) );
  NAND2_X1 U246 ( .A1(\mem[13][3] ), .A2(n570), .ZN(n566) );
  OAI21_X1 U247 ( .B1(n410), .B2(n570), .A(n565), .ZN(n434) );
  NAND2_X1 U248 ( .A1(\mem[13][4] ), .A2(n570), .ZN(n565) );
  OAI21_X1 U249 ( .B1(n409), .B2(n570), .A(n564), .ZN(n433) );
  NAND2_X1 U250 ( .A1(\mem[13][5] ), .A2(n570), .ZN(n564) );
  OAI21_X1 U251 ( .B1(n408), .B2(n570), .A(n563), .ZN(n432) );
  NAND2_X1 U252 ( .A1(\mem[13][6] ), .A2(n570), .ZN(n563) );
  OAI21_X1 U253 ( .B1(n407), .B2(n570), .A(n562), .ZN(n431) );
  NAND2_X1 U254 ( .A1(\mem[13][7] ), .A2(n570), .ZN(n562) );
  OAI21_X1 U255 ( .B1(n414), .B2(n561), .A(n560), .ZN(n430) );
  NAND2_X1 U256 ( .A1(\mem[14][0] ), .A2(n561), .ZN(n560) );
  OAI21_X1 U257 ( .B1(n413), .B2(n561), .A(n559), .ZN(n429) );
  NAND2_X1 U258 ( .A1(\mem[14][1] ), .A2(n561), .ZN(n559) );
  OAI21_X1 U259 ( .B1(n412), .B2(n561), .A(n558), .ZN(n428) );
  NAND2_X1 U260 ( .A1(\mem[14][2] ), .A2(n561), .ZN(n558) );
  OAI21_X1 U261 ( .B1(n411), .B2(n561), .A(n557), .ZN(n427) );
  NAND2_X1 U262 ( .A1(\mem[14][3] ), .A2(n561), .ZN(n557) );
  OAI21_X1 U263 ( .B1(n410), .B2(n561), .A(n556), .ZN(n426) );
  NAND2_X1 U264 ( .A1(\mem[14][4] ), .A2(n561), .ZN(n556) );
  OAI21_X1 U265 ( .B1(n409), .B2(n561), .A(n555), .ZN(n425) );
  NAND2_X1 U266 ( .A1(\mem[14][5] ), .A2(n561), .ZN(n555) );
  OAI21_X1 U267 ( .B1(n408), .B2(n561), .A(n554), .ZN(n424) );
  NAND2_X1 U268 ( .A1(\mem[14][6] ), .A2(n561), .ZN(n554) );
  OAI21_X1 U269 ( .B1(n407), .B2(n561), .A(n553), .ZN(n423) );
  NAND2_X1 U270 ( .A1(\mem[14][7] ), .A2(n561), .ZN(n553) );
  OAI21_X1 U271 ( .B1(n414), .B2(n551), .A(n550), .ZN(n422) );
  NAND2_X1 U272 ( .A1(\mem[15][0] ), .A2(n551), .ZN(n550) );
  OAI21_X1 U273 ( .B1(n413), .B2(n551), .A(n549), .ZN(n421) );
  NAND2_X1 U274 ( .A1(\mem[15][1] ), .A2(n551), .ZN(n549) );
  OAI21_X1 U275 ( .B1(n412), .B2(n551), .A(n548), .ZN(n420) );
  NAND2_X1 U276 ( .A1(\mem[15][2] ), .A2(n551), .ZN(n548) );
  OAI21_X1 U277 ( .B1(n411), .B2(n551), .A(n547), .ZN(n419) );
  NAND2_X1 U278 ( .A1(\mem[15][3] ), .A2(n551), .ZN(n547) );
  OAI21_X1 U279 ( .B1(n410), .B2(n551), .A(n546), .ZN(n418) );
  NAND2_X1 U280 ( .A1(\mem[15][4] ), .A2(n551), .ZN(n546) );
  OAI21_X1 U281 ( .B1(n409), .B2(n551), .A(n545), .ZN(n417) );
  NAND2_X1 U282 ( .A1(\mem[15][5] ), .A2(n551), .ZN(n545) );
  OAI21_X1 U283 ( .B1(n408), .B2(n551), .A(n544), .ZN(n416) );
  NAND2_X1 U284 ( .A1(\mem[15][6] ), .A2(n551), .ZN(n544) );
  OAI21_X1 U285 ( .B1(n407), .B2(n551), .A(n543), .ZN(n415) );
  NAND2_X1 U286 ( .A1(\mem[15][7] ), .A2(n551), .ZN(n543) );
  AND2_X1 U287 ( .A1(N13), .A2(wr_en), .ZN(n552) );
  NOR2_X1 U288 ( .A1(N11), .A2(N12), .ZN(n687) );
  NOR2_X1 U289 ( .A1(n405), .A2(N12), .ZN(n666) );
  AND2_X1 U290 ( .A1(N12), .A2(n405), .ZN(n647) );
  AND2_X1 U291 ( .A1(N12), .A2(N11), .ZN(n628) );
  INV_X1 U292 ( .A(data_in[0]), .ZN(n414) );
  INV_X1 U293 ( .A(data_in[1]), .ZN(n413) );
  INV_X1 U294 ( .A(data_in[2]), .ZN(n412) );
  INV_X1 U295 ( .A(data_in[3]), .ZN(n411) );
  INV_X1 U296 ( .A(data_in[4]), .ZN(n410) );
  INV_X1 U297 ( .A(data_in[5]), .ZN(n409) );
  INV_X1 U298 ( .A(data_in[6]), .ZN(n408) );
  INV_X1 U299 ( .A(data_in[7]), .ZN(n407) );
  MUX2_X1 U300 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(N10), .Z(n6) );
  MUX2_X1 U301 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n401), .Z(n7) );
  MUX2_X1 U302 ( .A(n7), .B(n6), .S(N11), .Z(n8) );
  MUX2_X1 U303 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(N10), .Z(n9) );
  MUX2_X1 U304 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n401), .Z(n10) );
  MUX2_X1 U305 ( .A(n10), .B(n9), .S(N11), .Z(n11) );
  MUX2_X1 U306 ( .A(n11), .B(n8), .S(N12), .Z(n294) );
  MUX2_X1 U307 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(N10), .Z(n295) );
  MUX2_X1 U308 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(N10), .Z(n296) );
  MUX2_X1 U309 ( .A(n296), .B(n295), .S(N11), .Z(n297) );
  MUX2_X1 U310 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(N10), .Z(n298) );
  MUX2_X1 U311 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n299) );
  MUX2_X1 U312 ( .A(n299), .B(n298), .S(N11), .Z(n300) );
  MUX2_X1 U313 ( .A(n300), .B(n297), .S(N12), .Z(n301) );
  MUX2_X1 U314 ( .A(n301), .B(n294), .S(N13), .Z(N21) );
  MUX2_X1 U315 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n402), .Z(n302) );
  MUX2_X1 U316 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(N10), .Z(n303) );
  MUX2_X1 U317 ( .A(n303), .B(n302), .S(N11), .Z(n304) );
  MUX2_X1 U318 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n403), .Z(n305) );
  MUX2_X1 U319 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(N10), .Z(n306) );
  MUX2_X1 U320 ( .A(n306), .B(n305), .S(N11), .Z(n307) );
  MUX2_X1 U321 ( .A(n307), .B(n304), .S(N12), .Z(n308) );
  MUX2_X1 U322 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(N10), .Z(n309) );
  MUX2_X1 U323 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(N10), .Z(n310) );
  MUX2_X1 U324 ( .A(n310), .B(n309), .S(N11), .Z(n311) );
  MUX2_X1 U325 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(N10), .Z(n312) );
  MUX2_X1 U326 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(N10), .Z(n313) );
  MUX2_X1 U327 ( .A(n313), .B(n312), .S(N11), .Z(n314) );
  MUX2_X1 U328 ( .A(n314), .B(n311), .S(N12), .Z(n315) );
  MUX2_X1 U329 ( .A(n315), .B(n308), .S(N13), .Z(N20) );
  MUX2_X1 U330 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n402), .Z(n316) );
  MUX2_X1 U331 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n402), .Z(n317) );
  MUX2_X1 U332 ( .A(n317), .B(n316), .S(n400), .Z(n318) );
  MUX2_X1 U333 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n403), .Z(n319) );
  MUX2_X1 U334 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(N10), .Z(n320) );
  MUX2_X1 U335 ( .A(n320), .B(n319), .S(n400), .Z(n321) );
  MUX2_X1 U336 ( .A(n321), .B(n318), .S(N12), .Z(n322) );
  MUX2_X1 U337 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n402), .Z(n323) );
  MUX2_X1 U338 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(N10), .Z(n324) );
  MUX2_X1 U339 ( .A(n324), .B(n323), .S(n400), .Z(n325) );
  MUX2_X1 U340 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n401), .Z(n326) );
  MUX2_X1 U341 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(N10), .Z(n327) );
  MUX2_X1 U342 ( .A(n327), .B(n326), .S(n400), .Z(n328) );
  MUX2_X1 U343 ( .A(n328), .B(n325), .S(N12), .Z(n329) );
  MUX2_X1 U344 ( .A(n329), .B(n322), .S(N13), .Z(N19) );
  MUX2_X1 U345 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n403), .Z(n330) );
  MUX2_X1 U346 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n403), .Z(n331) );
  MUX2_X1 U347 ( .A(n331), .B(n330), .S(n400), .Z(n332) );
  MUX2_X1 U348 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n401), .Z(n333) );
  MUX2_X1 U349 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n334) );
  MUX2_X1 U350 ( .A(n334), .B(n333), .S(n400), .Z(n335) );
  MUX2_X1 U351 ( .A(n335), .B(n332), .S(N12), .Z(n336) );
  MUX2_X1 U352 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n401), .Z(n337) );
  MUX2_X1 U353 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n401), .Z(n338) );
  MUX2_X1 U354 ( .A(n338), .B(n337), .S(n400), .Z(n339) );
  MUX2_X1 U355 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n401), .Z(n340) );
  MUX2_X1 U356 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n401), .Z(n341) );
  MUX2_X1 U357 ( .A(n341), .B(n340), .S(n400), .Z(n342) );
  MUX2_X1 U358 ( .A(n342), .B(n339), .S(N12), .Z(n343) );
  MUX2_X1 U359 ( .A(n343), .B(n336), .S(N13), .Z(N18) );
  MUX2_X1 U360 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n401), .Z(n344) );
  MUX2_X1 U361 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n401), .Z(n345) );
  MUX2_X1 U362 ( .A(n345), .B(n344), .S(n400), .Z(n346) );
  MUX2_X1 U363 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n401), .Z(n347) );
  MUX2_X1 U364 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n401), .Z(n348) );
  MUX2_X1 U365 ( .A(n348), .B(n347), .S(n400), .Z(n349) );
  MUX2_X1 U366 ( .A(n349), .B(n346), .S(N12), .Z(n350) );
  MUX2_X1 U367 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n401), .Z(n351) );
  MUX2_X1 U368 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n401), .Z(n352) );
  MUX2_X1 U369 ( .A(n352), .B(n351), .S(n400), .Z(n353) );
  MUX2_X1 U370 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n401), .Z(n354) );
  MUX2_X1 U371 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n401), .Z(n355) );
  MUX2_X1 U372 ( .A(n355), .B(n354), .S(n400), .Z(n356) );
  MUX2_X1 U373 ( .A(n356), .B(n353), .S(N12), .Z(n357) );
  MUX2_X1 U374 ( .A(n357), .B(n350), .S(N13), .Z(N17) );
  MUX2_X1 U375 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n402), .Z(n358) );
  MUX2_X1 U376 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n402), .Z(n359) );
  MUX2_X1 U377 ( .A(n359), .B(n358), .S(N11), .Z(n360) );
  MUX2_X1 U378 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n402), .Z(n361) );
  MUX2_X1 U379 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n402), .Z(n362) );
  MUX2_X1 U380 ( .A(n362), .B(n361), .S(N11), .Z(n363) );
  MUX2_X1 U381 ( .A(n363), .B(n360), .S(N12), .Z(n364) );
  MUX2_X1 U382 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n402), .Z(n365) );
  MUX2_X1 U383 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n402), .Z(n366) );
  MUX2_X1 U384 ( .A(n366), .B(n365), .S(N11), .Z(n367) );
  MUX2_X1 U385 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n402), .Z(n368) );
  MUX2_X1 U386 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n402), .Z(n369) );
  MUX2_X1 U387 ( .A(n369), .B(n368), .S(N11), .Z(n370) );
  MUX2_X1 U388 ( .A(n370), .B(n367), .S(N12), .Z(n371) );
  MUX2_X1 U389 ( .A(n371), .B(n364), .S(N13), .Z(N16) );
  MUX2_X1 U390 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n402), .Z(n372) );
  MUX2_X1 U391 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n402), .Z(n373) );
  MUX2_X1 U392 ( .A(n373), .B(n372), .S(N11), .Z(n374) );
  MUX2_X1 U393 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n402), .Z(n375) );
  MUX2_X1 U394 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n402), .Z(n376) );
  MUX2_X1 U395 ( .A(n376), .B(n375), .S(N11), .Z(n377) );
  MUX2_X1 U396 ( .A(n377), .B(n374), .S(N12), .Z(n378) );
  MUX2_X1 U397 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n403), .Z(n379) );
  MUX2_X1 U398 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n403), .Z(n380) );
  MUX2_X1 U399 ( .A(n380), .B(n379), .S(N11), .Z(n381) );
  MUX2_X1 U400 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n403), .Z(n382) );
  MUX2_X1 U401 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n403), .Z(n383) );
  MUX2_X1 U402 ( .A(n383), .B(n382), .S(n400), .Z(n384) );
  MUX2_X1 U403 ( .A(n384), .B(n381), .S(N12), .Z(n385) );
  MUX2_X1 U404 ( .A(n385), .B(n378), .S(N13), .Z(N15) );
  MUX2_X1 U405 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n403), .Z(n386) );
  MUX2_X1 U406 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n403), .Z(n387) );
  MUX2_X1 U407 ( .A(n387), .B(n386), .S(N11), .Z(n388) );
  MUX2_X1 U408 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n403), .Z(n389) );
  MUX2_X1 U409 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n403), .Z(n390) );
  MUX2_X1 U410 ( .A(n390), .B(n389), .S(N11), .Z(n391) );
  MUX2_X1 U411 ( .A(n391), .B(n388), .S(N12), .Z(n392) );
  MUX2_X1 U412 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n403), .Z(n393) );
  MUX2_X1 U413 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n403), .Z(n394) );
  MUX2_X1 U414 ( .A(n394), .B(n393), .S(N11), .Z(n395) );
  MUX2_X1 U415 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n403), .Z(n396) );
  MUX2_X1 U416 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n403), .Z(n397) );
  MUX2_X1 U417 ( .A(n397), .B(n396), .S(n400), .Z(n398) );
  MUX2_X1 U418 ( .A(n398), .B(n395), .S(N12), .Z(n399) );
  MUX2_X1 U419 ( .A(n399), .B(n392), .S(N13), .Z(N14) );
  INV_X1 U420 ( .A(N10), .ZN(n404) );
  INV_X1 U421 ( .A(N11), .ZN(n405) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_11 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, N19, N21, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n411), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n412), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n413), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n414), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n415), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n416), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n417), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n418), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n419), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n420), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n421), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n422), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n423), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n424), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n425), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n426), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n427), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n428), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n429), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n430), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n431), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n432), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n433), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n434), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n435), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n436), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n437), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n438), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n439), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n440), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n441), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n442), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n443), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n444), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n445), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n446), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n447), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n448), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n449), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n450), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n451), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n452), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n453), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n454), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n455), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n456), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n457), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n458), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n459), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n460), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n461), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n462), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n463), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n464), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n465), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n466), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n467), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n468), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n469), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n470), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n471), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n472), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n473), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n474), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n475), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n476), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n477), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n478), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n479), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n480), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n481), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n482), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n483), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n484), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n485), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n486), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n487), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n488), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n489), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n490), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n491), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n492), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n493), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n494), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n495), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n496), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n497), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n498), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n499), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n500), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n501), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n502), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n503), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n504), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n505), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n506), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n507), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n508), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n509), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n510), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n511), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n512), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n513), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n514), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n515), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n516), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n517), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n518), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n519), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n520), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n521), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n522), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n523), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n524), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n525), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n526), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n527), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n528), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n529), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n530), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n531), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n532), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n533), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n534), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n535), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n536), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n537), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n538), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .Q(data_out[3]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n311), .SI(n304), .SE(N13), .CK(clk), .Q(
        data_out[1]) );
  DFF_X1 \data_out_reg[5]  ( .D(N16), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(N10), .Z(n398) );
  BUF_X1 U4 ( .A(N10), .Z(n399) );
  BUF_X1 U5 ( .A(N11), .Z(n396) );
  NAND2_X1 U6 ( .A1(n662), .A2(n682), .ZN(n671) );
  NAND2_X1 U7 ( .A1(n662), .A2(n672), .ZN(n661) );
  NAND2_X1 U8 ( .A1(n683), .A2(n682), .ZN(n692) );
  NAND2_X1 U9 ( .A1(n672), .A2(n683), .ZN(n681) );
  NAND2_X1 U10 ( .A1(n604), .A2(n683), .ZN(n613) );
  NAND2_X1 U11 ( .A1(n594), .A2(n683), .ZN(n603) );
  NAND2_X1 U12 ( .A1(n604), .A2(n662), .ZN(n593) );
  NAND2_X1 U13 ( .A1(n594), .A2(n662), .ZN(n584) );
  NAND2_X1 U14 ( .A1(n643), .A2(n682), .ZN(n652) );
  NAND2_X1 U15 ( .A1(n643), .A2(n672), .ZN(n642) );
  NAND2_X1 U16 ( .A1(n624), .A2(n682), .ZN(n633) );
  NAND2_X1 U17 ( .A1(n624), .A2(n672), .ZN(n622) );
  NAND2_X1 U18 ( .A1(n604), .A2(n643), .ZN(n575) );
  NAND2_X1 U19 ( .A1(n594), .A2(n643), .ZN(n566) );
  NAND2_X1 U20 ( .A1(n604), .A2(n624), .ZN(n557) );
  NAND2_X1 U21 ( .A1(n594), .A2(n624), .ZN(n547) );
  AND2_X1 U22 ( .A1(n548), .A2(N10), .ZN(n594) );
  AND2_X1 U23 ( .A1(n548), .A2(n400), .ZN(n604) );
  AND2_X1 U24 ( .A1(N10), .A2(n623), .ZN(n672) );
  AND2_X1 U25 ( .A1(n623), .A2(n400), .ZN(n682) );
  OAI21_X1 U26 ( .B1(n692), .B2(n410), .A(n691), .ZN(n538) );
  NAND2_X1 U27 ( .A1(\mem[0][0] ), .A2(n692), .ZN(n691) );
  OAI21_X1 U28 ( .B1(n692), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U29 ( .A1(\mem[0][1] ), .A2(n692), .ZN(n690) );
  OAI21_X1 U30 ( .B1(n692), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U31 ( .A1(\mem[0][2] ), .A2(n692), .ZN(n689) );
  OAI21_X1 U32 ( .B1(n692), .B2(n407), .A(n688), .ZN(n535) );
  NAND2_X1 U33 ( .A1(\mem[0][3] ), .A2(n692), .ZN(n688) );
  OAI21_X1 U34 ( .B1(n692), .B2(n406), .A(n687), .ZN(n534) );
  NAND2_X1 U35 ( .A1(\mem[0][4] ), .A2(n692), .ZN(n687) );
  OAI21_X1 U36 ( .B1(n692), .B2(n405), .A(n686), .ZN(n533) );
  NAND2_X1 U37 ( .A1(\mem[0][5] ), .A2(n692), .ZN(n686) );
  OAI21_X1 U38 ( .B1(n692), .B2(n404), .A(n685), .ZN(n532) );
  NAND2_X1 U39 ( .A1(\mem[0][6] ), .A2(n692), .ZN(n685) );
  OAI21_X1 U40 ( .B1(n692), .B2(n403), .A(n684), .ZN(n531) );
  NAND2_X1 U41 ( .A1(\mem[0][7] ), .A2(n692), .ZN(n684) );
  OAI21_X1 U42 ( .B1(n410), .B2(n671), .A(n670), .ZN(n522) );
  NAND2_X1 U43 ( .A1(\mem[2][0] ), .A2(n671), .ZN(n670) );
  OAI21_X1 U44 ( .B1(n409), .B2(n671), .A(n669), .ZN(n521) );
  NAND2_X1 U45 ( .A1(\mem[2][1] ), .A2(n671), .ZN(n669) );
  OAI21_X1 U46 ( .B1(n408), .B2(n671), .A(n668), .ZN(n520) );
  NAND2_X1 U47 ( .A1(\mem[2][2] ), .A2(n671), .ZN(n668) );
  OAI21_X1 U48 ( .B1(n407), .B2(n671), .A(n667), .ZN(n519) );
  NAND2_X1 U49 ( .A1(\mem[2][3] ), .A2(n671), .ZN(n667) );
  OAI21_X1 U50 ( .B1(n406), .B2(n671), .A(n666), .ZN(n518) );
  NAND2_X1 U51 ( .A1(\mem[2][4] ), .A2(n671), .ZN(n666) );
  OAI21_X1 U52 ( .B1(n405), .B2(n671), .A(n665), .ZN(n517) );
  NAND2_X1 U53 ( .A1(\mem[2][5] ), .A2(n671), .ZN(n665) );
  OAI21_X1 U54 ( .B1(n404), .B2(n671), .A(n664), .ZN(n516) );
  NAND2_X1 U55 ( .A1(\mem[2][6] ), .A2(n671), .ZN(n664) );
  OAI21_X1 U56 ( .B1(n403), .B2(n671), .A(n663), .ZN(n515) );
  NAND2_X1 U57 ( .A1(\mem[2][7] ), .A2(n671), .ZN(n663) );
  OAI21_X1 U58 ( .B1(n410), .B2(n661), .A(n660), .ZN(n514) );
  NAND2_X1 U59 ( .A1(\mem[3][0] ), .A2(n661), .ZN(n660) );
  OAI21_X1 U60 ( .B1(n409), .B2(n661), .A(n659), .ZN(n513) );
  NAND2_X1 U61 ( .A1(\mem[3][1] ), .A2(n661), .ZN(n659) );
  OAI21_X1 U62 ( .B1(n408), .B2(n661), .A(n658), .ZN(n512) );
  NAND2_X1 U63 ( .A1(\mem[3][2] ), .A2(n661), .ZN(n658) );
  OAI21_X1 U64 ( .B1(n407), .B2(n661), .A(n657), .ZN(n511) );
  NAND2_X1 U65 ( .A1(\mem[3][3] ), .A2(n661), .ZN(n657) );
  OAI21_X1 U66 ( .B1(n406), .B2(n661), .A(n656), .ZN(n510) );
  NAND2_X1 U67 ( .A1(\mem[3][4] ), .A2(n661), .ZN(n656) );
  OAI21_X1 U68 ( .B1(n405), .B2(n661), .A(n655), .ZN(n509) );
  NAND2_X1 U69 ( .A1(\mem[3][5] ), .A2(n661), .ZN(n655) );
  OAI21_X1 U70 ( .B1(n404), .B2(n661), .A(n654), .ZN(n508) );
  NAND2_X1 U71 ( .A1(\mem[3][6] ), .A2(n661), .ZN(n654) );
  OAI21_X1 U72 ( .B1(n403), .B2(n661), .A(n653), .ZN(n507) );
  NAND2_X1 U73 ( .A1(\mem[3][7] ), .A2(n661), .ZN(n653) );
  NOR2_X1 U74 ( .A1(n402), .A2(N13), .ZN(n623) );
  INV_X1 U75 ( .A(wr_en), .ZN(n402) );
  OAI21_X1 U76 ( .B1(n410), .B2(n681), .A(n680), .ZN(n530) );
  NAND2_X1 U77 ( .A1(\mem[1][0] ), .A2(n681), .ZN(n680) );
  OAI21_X1 U78 ( .B1(n409), .B2(n681), .A(n679), .ZN(n529) );
  NAND2_X1 U79 ( .A1(\mem[1][1] ), .A2(n681), .ZN(n679) );
  OAI21_X1 U80 ( .B1(n408), .B2(n681), .A(n678), .ZN(n528) );
  NAND2_X1 U81 ( .A1(\mem[1][2] ), .A2(n681), .ZN(n678) );
  OAI21_X1 U82 ( .B1(n407), .B2(n681), .A(n677), .ZN(n527) );
  NAND2_X1 U83 ( .A1(\mem[1][3] ), .A2(n681), .ZN(n677) );
  OAI21_X1 U84 ( .B1(n406), .B2(n681), .A(n676), .ZN(n526) );
  NAND2_X1 U85 ( .A1(\mem[1][4] ), .A2(n681), .ZN(n676) );
  OAI21_X1 U86 ( .B1(n405), .B2(n681), .A(n675), .ZN(n525) );
  NAND2_X1 U87 ( .A1(\mem[1][5] ), .A2(n681), .ZN(n675) );
  OAI21_X1 U88 ( .B1(n404), .B2(n681), .A(n674), .ZN(n524) );
  NAND2_X1 U89 ( .A1(\mem[1][6] ), .A2(n681), .ZN(n674) );
  OAI21_X1 U90 ( .B1(n403), .B2(n681), .A(n673), .ZN(n523) );
  NAND2_X1 U91 ( .A1(\mem[1][7] ), .A2(n681), .ZN(n673) );
  OAI21_X1 U92 ( .B1(n410), .B2(n652), .A(n651), .ZN(n506) );
  NAND2_X1 U93 ( .A1(\mem[4][0] ), .A2(n652), .ZN(n651) );
  OAI21_X1 U94 ( .B1(n409), .B2(n652), .A(n650), .ZN(n505) );
  NAND2_X1 U95 ( .A1(\mem[4][1] ), .A2(n652), .ZN(n650) );
  OAI21_X1 U96 ( .B1(n408), .B2(n652), .A(n649), .ZN(n504) );
  NAND2_X1 U97 ( .A1(\mem[4][2] ), .A2(n652), .ZN(n649) );
  OAI21_X1 U98 ( .B1(n407), .B2(n652), .A(n648), .ZN(n503) );
  NAND2_X1 U99 ( .A1(\mem[4][3] ), .A2(n652), .ZN(n648) );
  OAI21_X1 U100 ( .B1(n406), .B2(n652), .A(n647), .ZN(n502) );
  NAND2_X1 U101 ( .A1(\mem[4][4] ), .A2(n652), .ZN(n647) );
  OAI21_X1 U102 ( .B1(n405), .B2(n652), .A(n646), .ZN(n501) );
  NAND2_X1 U103 ( .A1(\mem[4][5] ), .A2(n652), .ZN(n646) );
  OAI21_X1 U104 ( .B1(n404), .B2(n652), .A(n645), .ZN(n500) );
  NAND2_X1 U105 ( .A1(\mem[4][6] ), .A2(n652), .ZN(n645) );
  OAI21_X1 U106 ( .B1(n403), .B2(n652), .A(n644), .ZN(n499) );
  NAND2_X1 U107 ( .A1(\mem[4][7] ), .A2(n652), .ZN(n644) );
  OAI21_X1 U108 ( .B1(n410), .B2(n642), .A(n641), .ZN(n498) );
  NAND2_X1 U109 ( .A1(\mem[5][0] ), .A2(n642), .ZN(n641) );
  OAI21_X1 U110 ( .B1(n409), .B2(n642), .A(n640), .ZN(n497) );
  NAND2_X1 U111 ( .A1(\mem[5][1] ), .A2(n642), .ZN(n640) );
  OAI21_X1 U112 ( .B1(n408), .B2(n642), .A(n639), .ZN(n496) );
  NAND2_X1 U113 ( .A1(\mem[5][2] ), .A2(n642), .ZN(n639) );
  OAI21_X1 U114 ( .B1(n407), .B2(n642), .A(n638), .ZN(n495) );
  NAND2_X1 U115 ( .A1(\mem[5][3] ), .A2(n642), .ZN(n638) );
  OAI21_X1 U116 ( .B1(n406), .B2(n642), .A(n637), .ZN(n494) );
  NAND2_X1 U117 ( .A1(\mem[5][4] ), .A2(n642), .ZN(n637) );
  OAI21_X1 U118 ( .B1(n405), .B2(n642), .A(n636), .ZN(n493) );
  NAND2_X1 U119 ( .A1(\mem[5][5] ), .A2(n642), .ZN(n636) );
  OAI21_X1 U120 ( .B1(n404), .B2(n642), .A(n635), .ZN(n492) );
  NAND2_X1 U121 ( .A1(\mem[5][6] ), .A2(n642), .ZN(n635) );
  OAI21_X1 U122 ( .B1(n403), .B2(n642), .A(n634), .ZN(n491) );
  NAND2_X1 U123 ( .A1(\mem[5][7] ), .A2(n642), .ZN(n634) );
  OAI21_X1 U124 ( .B1(n410), .B2(n633), .A(n632), .ZN(n490) );
  NAND2_X1 U125 ( .A1(\mem[6][0] ), .A2(n633), .ZN(n632) );
  OAI21_X1 U126 ( .B1(n409), .B2(n633), .A(n631), .ZN(n489) );
  NAND2_X1 U127 ( .A1(\mem[6][1] ), .A2(n633), .ZN(n631) );
  OAI21_X1 U128 ( .B1(n408), .B2(n633), .A(n630), .ZN(n488) );
  NAND2_X1 U129 ( .A1(\mem[6][2] ), .A2(n633), .ZN(n630) );
  OAI21_X1 U130 ( .B1(n407), .B2(n633), .A(n629), .ZN(n487) );
  NAND2_X1 U131 ( .A1(\mem[6][3] ), .A2(n633), .ZN(n629) );
  OAI21_X1 U132 ( .B1(n406), .B2(n633), .A(n628), .ZN(n486) );
  NAND2_X1 U133 ( .A1(\mem[6][4] ), .A2(n633), .ZN(n628) );
  OAI21_X1 U134 ( .B1(n405), .B2(n633), .A(n627), .ZN(n485) );
  NAND2_X1 U135 ( .A1(\mem[6][5] ), .A2(n633), .ZN(n627) );
  OAI21_X1 U136 ( .B1(n404), .B2(n633), .A(n626), .ZN(n484) );
  NAND2_X1 U137 ( .A1(\mem[6][6] ), .A2(n633), .ZN(n626) );
  OAI21_X1 U138 ( .B1(n403), .B2(n633), .A(n625), .ZN(n483) );
  NAND2_X1 U139 ( .A1(\mem[6][7] ), .A2(n633), .ZN(n625) );
  OAI21_X1 U140 ( .B1(n410), .B2(n622), .A(n621), .ZN(n482) );
  NAND2_X1 U141 ( .A1(\mem[7][0] ), .A2(n622), .ZN(n621) );
  OAI21_X1 U142 ( .B1(n409), .B2(n622), .A(n620), .ZN(n481) );
  NAND2_X1 U143 ( .A1(\mem[7][1] ), .A2(n622), .ZN(n620) );
  OAI21_X1 U144 ( .B1(n408), .B2(n622), .A(n619), .ZN(n480) );
  NAND2_X1 U145 ( .A1(\mem[7][2] ), .A2(n622), .ZN(n619) );
  OAI21_X1 U146 ( .B1(n407), .B2(n622), .A(n618), .ZN(n479) );
  NAND2_X1 U147 ( .A1(\mem[7][3] ), .A2(n622), .ZN(n618) );
  OAI21_X1 U148 ( .B1(n406), .B2(n622), .A(n617), .ZN(n478) );
  NAND2_X1 U149 ( .A1(\mem[7][4] ), .A2(n622), .ZN(n617) );
  OAI21_X1 U150 ( .B1(n405), .B2(n622), .A(n616), .ZN(n477) );
  NAND2_X1 U151 ( .A1(\mem[7][5] ), .A2(n622), .ZN(n616) );
  OAI21_X1 U152 ( .B1(n404), .B2(n622), .A(n615), .ZN(n476) );
  NAND2_X1 U153 ( .A1(\mem[7][6] ), .A2(n622), .ZN(n615) );
  OAI21_X1 U154 ( .B1(n403), .B2(n622), .A(n614), .ZN(n475) );
  NAND2_X1 U155 ( .A1(\mem[7][7] ), .A2(n622), .ZN(n614) );
  OAI21_X1 U156 ( .B1(n410), .B2(n613), .A(n612), .ZN(n474) );
  NAND2_X1 U157 ( .A1(\mem[8][0] ), .A2(n613), .ZN(n612) );
  OAI21_X1 U158 ( .B1(n409), .B2(n613), .A(n611), .ZN(n473) );
  NAND2_X1 U159 ( .A1(\mem[8][1] ), .A2(n613), .ZN(n611) );
  OAI21_X1 U160 ( .B1(n408), .B2(n613), .A(n610), .ZN(n472) );
  NAND2_X1 U161 ( .A1(\mem[8][2] ), .A2(n613), .ZN(n610) );
  OAI21_X1 U162 ( .B1(n407), .B2(n613), .A(n609), .ZN(n471) );
  NAND2_X1 U163 ( .A1(\mem[8][3] ), .A2(n613), .ZN(n609) );
  OAI21_X1 U164 ( .B1(n406), .B2(n613), .A(n608), .ZN(n470) );
  NAND2_X1 U165 ( .A1(\mem[8][4] ), .A2(n613), .ZN(n608) );
  OAI21_X1 U166 ( .B1(n405), .B2(n613), .A(n607), .ZN(n469) );
  NAND2_X1 U167 ( .A1(\mem[8][5] ), .A2(n613), .ZN(n607) );
  OAI21_X1 U168 ( .B1(n404), .B2(n613), .A(n606), .ZN(n468) );
  NAND2_X1 U169 ( .A1(\mem[8][6] ), .A2(n613), .ZN(n606) );
  OAI21_X1 U170 ( .B1(n403), .B2(n613), .A(n605), .ZN(n467) );
  NAND2_X1 U171 ( .A1(\mem[8][7] ), .A2(n613), .ZN(n605) );
  OAI21_X1 U172 ( .B1(n410), .B2(n603), .A(n602), .ZN(n466) );
  NAND2_X1 U173 ( .A1(\mem[9][0] ), .A2(n603), .ZN(n602) );
  OAI21_X1 U174 ( .B1(n409), .B2(n603), .A(n601), .ZN(n465) );
  NAND2_X1 U175 ( .A1(\mem[9][1] ), .A2(n603), .ZN(n601) );
  OAI21_X1 U176 ( .B1(n408), .B2(n603), .A(n600), .ZN(n464) );
  NAND2_X1 U177 ( .A1(\mem[9][2] ), .A2(n603), .ZN(n600) );
  OAI21_X1 U178 ( .B1(n407), .B2(n603), .A(n599), .ZN(n463) );
  NAND2_X1 U179 ( .A1(\mem[9][3] ), .A2(n603), .ZN(n599) );
  OAI21_X1 U180 ( .B1(n406), .B2(n603), .A(n598), .ZN(n462) );
  NAND2_X1 U181 ( .A1(\mem[9][4] ), .A2(n603), .ZN(n598) );
  OAI21_X1 U182 ( .B1(n405), .B2(n603), .A(n597), .ZN(n461) );
  NAND2_X1 U183 ( .A1(\mem[9][5] ), .A2(n603), .ZN(n597) );
  OAI21_X1 U184 ( .B1(n404), .B2(n603), .A(n596), .ZN(n460) );
  NAND2_X1 U185 ( .A1(\mem[9][6] ), .A2(n603), .ZN(n596) );
  OAI21_X1 U186 ( .B1(n403), .B2(n603), .A(n595), .ZN(n459) );
  NAND2_X1 U187 ( .A1(\mem[9][7] ), .A2(n603), .ZN(n595) );
  OAI21_X1 U188 ( .B1(n410), .B2(n593), .A(n592), .ZN(n458) );
  NAND2_X1 U189 ( .A1(\mem[10][0] ), .A2(n593), .ZN(n592) );
  OAI21_X1 U190 ( .B1(n409), .B2(n593), .A(n591), .ZN(n457) );
  NAND2_X1 U191 ( .A1(\mem[10][1] ), .A2(n593), .ZN(n591) );
  OAI21_X1 U192 ( .B1(n408), .B2(n593), .A(n590), .ZN(n456) );
  NAND2_X1 U193 ( .A1(\mem[10][2] ), .A2(n593), .ZN(n590) );
  OAI21_X1 U194 ( .B1(n407), .B2(n593), .A(n589), .ZN(n455) );
  NAND2_X1 U195 ( .A1(\mem[10][3] ), .A2(n593), .ZN(n589) );
  OAI21_X1 U196 ( .B1(n406), .B2(n593), .A(n588), .ZN(n454) );
  NAND2_X1 U197 ( .A1(\mem[10][4] ), .A2(n593), .ZN(n588) );
  OAI21_X1 U198 ( .B1(n405), .B2(n593), .A(n587), .ZN(n453) );
  NAND2_X1 U199 ( .A1(\mem[10][5] ), .A2(n593), .ZN(n587) );
  OAI21_X1 U200 ( .B1(n404), .B2(n593), .A(n586), .ZN(n452) );
  NAND2_X1 U201 ( .A1(\mem[10][6] ), .A2(n593), .ZN(n586) );
  OAI21_X1 U202 ( .B1(n403), .B2(n593), .A(n585), .ZN(n451) );
  NAND2_X1 U203 ( .A1(\mem[10][7] ), .A2(n593), .ZN(n585) );
  OAI21_X1 U204 ( .B1(n410), .B2(n584), .A(n583), .ZN(n450) );
  NAND2_X1 U205 ( .A1(\mem[11][0] ), .A2(n584), .ZN(n583) );
  OAI21_X1 U206 ( .B1(n409), .B2(n584), .A(n582), .ZN(n449) );
  NAND2_X1 U207 ( .A1(\mem[11][1] ), .A2(n584), .ZN(n582) );
  OAI21_X1 U208 ( .B1(n408), .B2(n584), .A(n581), .ZN(n448) );
  NAND2_X1 U209 ( .A1(\mem[11][2] ), .A2(n584), .ZN(n581) );
  OAI21_X1 U210 ( .B1(n407), .B2(n584), .A(n580), .ZN(n447) );
  NAND2_X1 U211 ( .A1(\mem[11][3] ), .A2(n584), .ZN(n580) );
  OAI21_X1 U212 ( .B1(n406), .B2(n584), .A(n579), .ZN(n446) );
  NAND2_X1 U213 ( .A1(\mem[11][4] ), .A2(n584), .ZN(n579) );
  OAI21_X1 U214 ( .B1(n405), .B2(n584), .A(n578), .ZN(n445) );
  NAND2_X1 U215 ( .A1(\mem[11][5] ), .A2(n584), .ZN(n578) );
  OAI21_X1 U216 ( .B1(n404), .B2(n584), .A(n577), .ZN(n444) );
  NAND2_X1 U217 ( .A1(\mem[11][6] ), .A2(n584), .ZN(n577) );
  OAI21_X1 U218 ( .B1(n403), .B2(n584), .A(n576), .ZN(n443) );
  NAND2_X1 U219 ( .A1(\mem[11][7] ), .A2(n584), .ZN(n576) );
  OAI21_X1 U220 ( .B1(n410), .B2(n575), .A(n574), .ZN(n442) );
  NAND2_X1 U221 ( .A1(\mem[12][0] ), .A2(n575), .ZN(n574) );
  OAI21_X1 U222 ( .B1(n409), .B2(n575), .A(n573), .ZN(n441) );
  NAND2_X1 U223 ( .A1(\mem[12][1] ), .A2(n575), .ZN(n573) );
  OAI21_X1 U224 ( .B1(n408), .B2(n575), .A(n572), .ZN(n440) );
  NAND2_X1 U225 ( .A1(\mem[12][2] ), .A2(n575), .ZN(n572) );
  OAI21_X1 U226 ( .B1(n407), .B2(n575), .A(n571), .ZN(n439) );
  NAND2_X1 U227 ( .A1(\mem[12][3] ), .A2(n575), .ZN(n571) );
  OAI21_X1 U228 ( .B1(n406), .B2(n575), .A(n570), .ZN(n438) );
  NAND2_X1 U229 ( .A1(\mem[12][4] ), .A2(n575), .ZN(n570) );
  OAI21_X1 U230 ( .B1(n405), .B2(n575), .A(n569), .ZN(n437) );
  NAND2_X1 U231 ( .A1(\mem[12][5] ), .A2(n575), .ZN(n569) );
  OAI21_X1 U232 ( .B1(n404), .B2(n575), .A(n568), .ZN(n436) );
  NAND2_X1 U233 ( .A1(\mem[12][6] ), .A2(n575), .ZN(n568) );
  OAI21_X1 U234 ( .B1(n403), .B2(n575), .A(n567), .ZN(n435) );
  NAND2_X1 U235 ( .A1(\mem[12][7] ), .A2(n575), .ZN(n567) );
  OAI21_X1 U236 ( .B1(n410), .B2(n566), .A(n565), .ZN(n434) );
  NAND2_X1 U237 ( .A1(\mem[13][0] ), .A2(n566), .ZN(n565) );
  OAI21_X1 U238 ( .B1(n409), .B2(n566), .A(n564), .ZN(n433) );
  NAND2_X1 U239 ( .A1(\mem[13][1] ), .A2(n566), .ZN(n564) );
  OAI21_X1 U240 ( .B1(n408), .B2(n566), .A(n563), .ZN(n432) );
  NAND2_X1 U241 ( .A1(\mem[13][2] ), .A2(n566), .ZN(n563) );
  OAI21_X1 U242 ( .B1(n407), .B2(n566), .A(n562), .ZN(n431) );
  NAND2_X1 U243 ( .A1(\mem[13][3] ), .A2(n566), .ZN(n562) );
  OAI21_X1 U244 ( .B1(n406), .B2(n566), .A(n561), .ZN(n430) );
  NAND2_X1 U245 ( .A1(\mem[13][4] ), .A2(n566), .ZN(n561) );
  OAI21_X1 U246 ( .B1(n405), .B2(n566), .A(n560), .ZN(n429) );
  NAND2_X1 U247 ( .A1(\mem[13][5] ), .A2(n566), .ZN(n560) );
  OAI21_X1 U248 ( .B1(n404), .B2(n566), .A(n559), .ZN(n428) );
  NAND2_X1 U249 ( .A1(\mem[13][6] ), .A2(n566), .ZN(n559) );
  OAI21_X1 U250 ( .B1(n403), .B2(n566), .A(n558), .ZN(n427) );
  NAND2_X1 U251 ( .A1(\mem[13][7] ), .A2(n566), .ZN(n558) );
  OAI21_X1 U252 ( .B1(n410), .B2(n557), .A(n556), .ZN(n426) );
  NAND2_X1 U253 ( .A1(\mem[14][0] ), .A2(n557), .ZN(n556) );
  OAI21_X1 U254 ( .B1(n409), .B2(n557), .A(n555), .ZN(n425) );
  NAND2_X1 U255 ( .A1(\mem[14][1] ), .A2(n557), .ZN(n555) );
  OAI21_X1 U256 ( .B1(n408), .B2(n557), .A(n554), .ZN(n424) );
  NAND2_X1 U257 ( .A1(\mem[14][2] ), .A2(n557), .ZN(n554) );
  OAI21_X1 U258 ( .B1(n407), .B2(n557), .A(n553), .ZN(n423) );
  NAND2_X1 U259 ( .A1(\mem[14][3] ), .A2(n557), .ZN(n553) );
  OAI21_X1 U260 ( .B1(n406), .B2(n557), .A(n552), .ZN(n422) );
  NAND2_X1 U261 ( .A1(\mem[14][4] ), .A2(n557), .ZN(n552) );
  OAI21_X1 U262 ( .B1(n405), .B2(n557), .A(n551), .ZN(n421) );
  NAND2_X1 U263 ( .A1(\mem[14][5] ), .A2(n557), .ZN(n551) );
  OAI21_X1 U264 ( .B1(n404), .B2(n557), .A(n550), .ZN(n420) );
  NAND2_X1 U265 ( .A1(\mem[14][6] ), .A2(n557), .ZN(n550) );
  OAI21_X1 U266 ( .B1(n403), .B2(n557), .A(n549), .ZN(n419) );
  NAND2_X1 U267 ( .A1(\mem[14][7] ), .A2(n557), .ZN(n549) );
  OAI21_X1 U268 ( .B1(n410), .B2(n547), .A(n546), .ZN(n418) );
  NAND2_X1 U269 ( .A1(\mem[15][0] ), .A2(n547), .ZN(n546) );
  OAI21_X1 U270 ( .B1(n409), .B2(n547), .A(n545), .ZN(n417) );
  NAND2_X1 U271 ( .A1(\mem[15][1] ), .A2(n547), .ZN(n545) );
  OAI21_X1 U272 ( .B1(n408), .B2(n547), .A(n544), .ZN(n416) );
  NAND2_X1 U273 ( .A1(\mem[15][2] ), .A2(n547), .ZN(n544) );
  OAI21_X1 U274 ( .B1(n407), .B2(n547), .A(n543), .ZN(n415) );
  NAND2_X1 U275 ( .A1(\mem[15][3] ), .A2(n547), .ZN(n543) );
  OAI21_X1 U276 ( .B1(n406), .B2(n547), .A(n542), .ZN(n414) );
  NAND2_X1 U277 ( .A1(\mem[15][4] ), .A2(n547), .ZN(n542) );
  OAI21_X1 U278 ( .B1(n405), .B2(n547), .A(n541), .ZN(n413) );
  NAND2_X1 U279 ( .A1(\mem[15][5] ), .A2(n547), .ZN(n541) );
  OAI21_X1 U280 ( .B1(n404), .B2(n547), .A(n540), .ZN(n412) );
  NAND2_X1 U281 ( .A1(\mem[15][6] ), .A2(n547), .ZN(n540) );
  OAI21_X1 U282 ( .B1(n403), .B2(n547), .A(n539), .ZN(n411) );
  NAND2_X1 U283 ( .A1(\mem[15][7] ), .A2(n547), .ZN(n539) );
  AND2_X1 U284 ( .A1(N13), .A2(wr_en), .ZN(n548) );
  NOR2_X1 U285 ( .A1(N11), .A2(N12), .ZN(n683) );
  NOR2_X1 U286 ( .A1(n401), .A2(N12), .ZN(n662) );
  AND2_X1 U287 ( .A1(N12), .A2(n401), .ZN(n643) );
  AND2_X1 U288 ( .A1(N12), .A2(N11), .ZN(n624) );
  INV_X1 U289 ( .A(data_in[0]), .ZN(n410) );
  INV_X1 U290 ( .A(data_in[1]), .ZN(n409) );
  INV_X1 U291 ( .A(data_in[2]), .ZN(n408) );
  INV_X1 U292 ( .A(data_in[3]), .ZN(n407) );
  INV_X1 U293 ( .A(data_in[4]), .ZN(n406) );
  INV_X1 U294 ( .A(data_in[5]), .ZN(n405) );
  INV_X1 U295 ( .A(data_in[6]), .ZN(n404) );
  INV_X1 U296 ( .A(data_in[7]), .ZN(n403) );
  MUX2_X1 U297 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n397), .Z(n2) );
  MUX2_X1 U298 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n397), .Z(n3) );
  MUX2_X1 U299 ( .A(n3), .B(n2), .S(N11), .Z(n4) );
  MUX2_X1 U300 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n397), .Z(n5) );
  MUX2_X1 U301 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n397), .Z(n6) );
  MUX2_X1 U302 ( .A(n6), .B(n5), .S(N11), .Z(n7) );
  MUX2_X1 U303 ( .A(n7), .B(n4), .S(N12), .Z(n8) );
  MUX2_X1 U304 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n398), .Z(n9) );
  MUX2_X1 U305 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n398), .Z(n10) );
  MUX2_X1 U306 ( .A(n10), .B(n9), .S(N11), .Z(n11) );
  MUX2_X1 U307 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n398), .Z(n294) );
  MUX2_X1 U308 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n398), .Z(n295) );
  MUX2_X1 U309 ( .A(n295), .B(n294), .S(N11), .Z(n296) );
  MUX2_X1 U310 ( .A(n296), .B(n11), .S(N12), .Z(n297) );
  MUX2_X1 U311 ( .A(n297), .B(n8), .S(N13), .Z(N21) );
  MUX2_X1 U312 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n398), .Z(n298) );
  MUX2_X1 U313 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n398), .Z(n299) );
  MUX2_X1 U314 ( .A(n299), .B(n298), .S(N11), .Z(n300) );
  MUX2_X1 U315 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n398), .Z(n301) );
  MUX2_X1 U316 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n398), .Z(n302) );
  MUX2_X1 U317 ( .A(n302), .B(n301), .S(N11), .Z(n303) );
  MUX2_X1 U318 ( .A(n303), .B(n300), .S(N12), .Z(n304) );
  MUX2_X1 U319 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n398), .Z(n305) );
  MUX2_X1 U320 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n398), .Z(n306) );
  MUX2_X1 U321 ( .A(n306), .B(n305), .S(N11), .Z(n307) );
  MUX2_X1 U322 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n398), .Z(n308) );
  MUX2_X1 U323 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n398), .Z(n309) );
  MUX2_X1 U324 ( .A(n309), .B(n308), .S(N11), .Z(n310) );
  MUX2_X1 U325 ( .A(n310), .B(n307), .S(N12), .Z(n311) );
  MUX2_X1 U326 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n399), .Z(n312) );
  MUX2_X1 U327 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n399), .Z(n313) );
  MUX2_X1 U328 ( .A(n313), .B(n312), .S(n396), .Z(n314) );
  MUX2_X1 U329 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n399), .Z(n315) );
  MUX2_X1 U330 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n399), .Z(n316) );
  MUX2_X1 U331 ( .A(n316), .B(n315), .S(n396), .Z(n317) );
  MUX2_X1 U332 ( .A(n317), .B(n314), .S(N12), .Z(n318) );
  MUX2_X1 U333 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n399), .Z(n319) );
  MUX2_X1 U334 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n399), .Z(n320) );
  MUX2_X1 U335 ( .A(n320), .B(n319), .S(n396), .Z(n321) );
  MUX2_X1 U336 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n399), .Z(n322) );
  MUX2_X1 U337 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n399), .Z(n323) );
  MUX2_X1 U338 ( .A(n323), .B(n322), .S(n396), .Z(n324) );
  MUX2_X1 U339 ( .A(n324), .B(n321), .S(N12), .Z(n325) );
  MUX2_X1 U340 ( .A(n325), .B(n318), .S(N13), .Z(N19) );
  MUX2_X1 U341 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n399), .Z(n326) );
  MUX2_X1 U342 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n399), .Z(n327) );
  MUX2_X1 U343 ( .A(n327), .B(n326), .S(n396), .Z(n328) );
  MUX2_X1 U344 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n399), .Z(n329) );
  MUX2_X1 U345 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n399), .Z(n330) );
  MUX2_X1 U346 ( .A(n330), .B(n329), .S(n396), .Z(n331) );
  MUX2_X1 U347 ( .A(n331), .B(n328), .S(N12), .Z(n332) );
  MUX2_X1 U348 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(N10), .Z(n333) );
  MUX2_X1 U349 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n399), .Z(n334) );
  MUX2_X1 U350 ( .A(n334), .B(n333), .S(n396), .Z(n335) );
  MUX2_X1 U351 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n397), .Z(n336) );
  MUX2_X1 U352 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n399), .Z(n337) );
  MUX2_X1 U353 ( .A(n337), .B(n336), .S(n396), .Z(n338) );
  MUX2_X1 U354 ( .A(n338), .B(n335), .S(N12), .Z(n339) );
  MUX2_X1 U355 ( .A(n339), .B(n332), .S(N13), .Z(N18) );
  MUX2_X1 U356 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n399), .Z(n340) );
  MUX2_X1 U357 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n399), .Z(n341) );
  MUX2_X1 U358 ( .A(n341), .B(n340), .S(n396), .Z(n342) );
  MUX2_X1 U359 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n398), .Z(n343) );
  MUX2_X1 U360 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n398), .Z(n344) );
  MUX2_X1 U361 ( .A(n344), .B(n343), .S(n396), .Z(n345) );
  MUX2_X1 U362 ( .A(n345), .B(n342), .S(N12), .Z(n346) );
  MUX2_X1 U363 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n397), .Z(n347) );
  MUX2_X1 U364 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n397), .Z(n348) );
  MUX2_X1 U365 ( .A(n348), .B(n347), .S(n396), .Z(n349) );
  MUX2_X1 U366 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n398), .Z(n350) );
  MUX2_X1 U367 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n397), .Z(n351) );
  MUX2_X1 U368 ( .A(n351), .B(n350), .S(n396), .Z(n352) );
  MUX2_X1 U369 ( .A(n352), .B(n349), .S(N12), .Z(n353) );
  MUX2_X1 U370 ( .A(n353), .B(n346), .S(N13), .Z(N17) );
  MUX2_X1 U371 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n398), .Z(n354) );
  MUX2_X1 U372 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(N10), .Z(n355) );
  MUX2_X1 U373 ( .A(n355), .B(n354), .S(N11), .Z(n356) );
  MUX2_X1 U374 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n398), .Z(n357) );
  MUX2_X1 U375 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(N10), .Z(n358) );
  MUX2_X1 U376 ( .A(n358), .B(n357), .S(N11), .Z(n359) );
  MUX2_X1 U377 ( .A(n359), .B(n356), .S(N12), .Z(n360) );
  MUX2_X1 U378 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(N10), .Z(n361) );
  MUX2_X1 U379 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(N10), .Z(n362) );
  MUX2_X1 U380 ( .A(n362), .B(n361), .S(N11), .Z(n363) );
  MUX2_X1 U381 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n364) );
  MUX2_X1 U382 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(N10), .Z(n365) );
  MUX2_X1 U383 ( .A(n365), .B(n364), .S(n396), .Z(n366) );
  MUX2_X1 U384 ( .A(n366), .B(n363), .S(N12), .Z(n367) );
  MUX2_X1 U385 ( .A(n367), .B(n360), .S(N13), .Z(N16) );
  MUX2_X1 U386 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n399), .Z(n368) );
  MUX2_X1 U387 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(N10), .Z(n369) );
  MUX2_X1 U388 ( .A(n369), .B(n368), .S(N11), .Z(n370) );
  MUX2_X1 U389 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(N10), .Z(n371) );
  MUX2_X1 U390 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n372) );
  MUX2_X1 U391 ( .A(n372), .B(n371), .S(N11), .Z(n373) );
  MUX2_X1 U392 ( .A(n373), .B(n370), .S(N12), .Z(n374) );
  MUX2_X1 U393 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n397), .Z(n375) );
  MUX2_X1 U394 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n397), .Z(n376) );
  MUX2_X1 U395 ( .A(n376), .B(n375), .S(N11), .Z(n377) );
  MUX2_X1 U396 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n378) );
  MUX2_X1 U397 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n379) );
  MUX2_X1 U398 ( .A(n379), .B(n378), .S(n396), .Z(n380) );
  MUX2_X1 U399 ( .A(n380), .B(n377), .S(N12), .Z(n381) );
  MUX2_X1 U400 ( .A(n381), .B(n374), .S(N13), .Z(N15) );
  MUX2_X1 U401 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n397), .Z(n382) );
  MUX2_X1 U402 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n397), .Z(n383) );
  MUX2_X1 U403 ( .A(n383), .B(n382), .S(N11), .Z(n384) );
  MUX2_X1 U404 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n397), .Z(n385) );
  MUX2_X1 U405 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n397), .Z(n386) );
  MUX2_X1 U406 ( .A(n386), .B(n385), .S(N11), .Z(n387) );
  MUX2_X1 U407 ( .A(n387), .B(n384), .S(N12), .Z(n388) );
  MUX2_X1 U408 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n397), .Z(n389) );
  MUX2_X1 U409 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n390) );
  MUX2_X1 U410 ( .A(n390), .B(n389), .S(N11), .Z(n391) );
  MUX2_X1 U411 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n392) );
  MUX2_X1 U412 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n393) );
  MUX2_X1 U413 ( .A(n393), .B(n392), .S(n396), .Z(n394) );
  MUX2_X1 U414 ( .A(n394), .B(n391), .S(N12), .Z(n395) );
  MUX2_X1 U415 ( .A(n395), .B(n388), .S(N13), .Z(N14) );
  CLKBUF_X1 U416 ( .A(N10), .Z(n397) );
  INV_X1 U417 ( .A(N10), .ZN(n400) );
  INV_X1 U418 ( .A(N11), .ZN(n401) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_10 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N19, N20, N21, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n411), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n412), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n413), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n414), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n415), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n416), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n417), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n418), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n419), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n420), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n421), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n422), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n423), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n424), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n425), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n426), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n427), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n428), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n429), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n430), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n431), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n432), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n433), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n434), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n435), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n436), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n437), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n438), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n439), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n440), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n441), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n442), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n443), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n444), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n445), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n446), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n447), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n448), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n449), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n450), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n451), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n452), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n453), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n454), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n455), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n456), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n457), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n458), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n459), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n460), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n461), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n462), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n463), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n464), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n465), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n466), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n467), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n468), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n469), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n470), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n471), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n472), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n473), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n474), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n475), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n476), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n477), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n478), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n479), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n480), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n481), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n482), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n483), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n484), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n485), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n486), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n487), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n488), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n489), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n490), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n491), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n492), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n493), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n494), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n495), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n496), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n497), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n498), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n499), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n500), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n501), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n502), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n503), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n504), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n505), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n506), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n507), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n508), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n509), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n510), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n511), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n512), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n513), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n514), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n515), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n516), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n517), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n518), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n519), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n520), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n521), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n522), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n523), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n524), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n525), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n526), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n527), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n528), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n529), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n530), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n531), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n532), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n533), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n534), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n535), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n536), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n537), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n538), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N20), .CK(clk), .Q(data_out[1]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n339), .SI(n332), .SE(N13), .CK(clk), .Q(
        data_out[3]) );
  DFF_X1 \data_out_reg[5]  ( .D(N16), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(N10), .Z(n397) );
  BUF_X1 U4 ( .A(N10), .Z(n398) );
  BUF_X1 U5 ( .A(N10), .Z(n399) );
  BUF_X1 U6 ( .A(N11), .Z(n396) );
  NAND2_X1 U7 ( .A1(n662), .A2(n682), .ZN(n671) );
  NAND2_X1 U8 ( .A1(n662), .A2(n672), .ZN(n661) );
  NAND2_X1 U9 ( .A1(n683), .A2(n682), .ZN(n692) );
  NAND2_X1 U10 ( .A1(n672), .A2(n683), .ZN(n681) );
  NAND2_X1 U11 ( .A1(n604), .A2(n683), .ZN(n613) );
  NAND2_X1 U12 ( .A1(n594), .A2(n683), .ZN(n603) );
  NAND2_X1 U13 ( .A1(n604), .A2(n662), .ZN(n593) );
  NAND2_X1 U14 ( .A1(n594), .A2(n662), .ZN(n584) );
  NAND2_X1 U15 ( .A1(n643), .A2(n682), .ZN(n652) );
  NAND2_X1 U16 ( .A1(n643), .A2(n672), .ZN(n642) );
  NAND2_X1 U17 ( .A1(n624), .A2(n682), .ZN(n633) );
  NAND2_X1 U18 ( .A1(n624), .A2(n672), .ZN(n622) );
  NAND2_X1 U19 ( .A1(n604), .A2(n643), .ZN(n575) );
  NAND2_X1 U20 ( .A1(n594), .A2(n643), .ZN(n566) );
  NAND2_X1 U21 ( .A1(n604), .A2(n624), .ZN(n557) );
  NAND2_X1 U22 ( .A1(n594), .A2(n624), .ZN(n547) );
  AND2_X1 U23 ( .A1(n548), .A2(N10), .ZN(n594) );
  AND2_X1 U24 ( .A1(n548), .A2(n400), .ZN(n604) );
  AND2_X1 U25 ( .A1(N10), .A2(n623), .ZN(n672) );
  AND2_X1 U26 ( .A1(n623), .A2(n400), .ZN(n682) );
  OAI21_X1 U27 ( .B1(n692), .B2(n410), .A(n691), .ZN(n538) );
  NAND2_X1 U28 ( .A1(\mem[0][0] ), .A2(n692), .ZN(n691) );
  OAI21_X1 U29 ( .B1(n692), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U30 ( .A1(\mem[0][1] ), .A2(n692), .ZN(n690) );
  OAI21_X1 U31 ( .B1(n692), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U32 ( .A1(\mem[0][2] ), .A2(n692), .ZN(n689) );
  OAI21_X1 U33 ( .B1(n692), .B2(n407), .A(n688), .ZN(n535) );
  NAND2_X1 U34 ( .A1(\mem[0][3] ), .A2(n692), .ZN(n688) );
  OAI21_X1 U35 ( .B1(n692), .B2(n406), .A(n687), .ZN(n534) );
  NAND2_X1 U36 ( .A1(\mem[0][4] ), .A2(n692), .ZN(n687) );
  OAI21_X1 U37 ( .B1(n692), .B2(n405), .A(n686), .ZN(n533) );
  NAND2_X1 U38 ( .A1(\mem[0][5] ), .A2(n692), .ZN(n686) );
  OAI21_X1 U39 ( .B1(n692), .B2(n404), .A(n685), .ZN(n532) );
  NAND2_X1 U40 ( .A1(\mem[0][6] ), .A2(n692), .ZN(n685) );
  OAI21_X1 U41 ( .B1(n692), .B2(n403), .A(n684), .ZN(n531) );
  NAND2_X1 U42 ( .A1(\mem[0][7] ), .A2(n692), .ZN(n684) );
  OAI21_X1 U43 ( .B1(n410), .B2(n671), .A(n670), .ZN(n522) );
  NAND2_X1 U44 ( .A1(\mem[2][0] ), .A2(n671), .ZN(n670) );
  OAI21_X1 U45 ( .B1(n409), .B2(n671), .A(n669), .ZN(n521) );
  NAND2_X1 U46 ( .A1(\mem[2][1] ), .A2(n671), .ZN(n669) );
  OAI21_X1 U47 ( .B1(n408), .B2(n671), .A(n668), .ZN(n520) );
  NAND2_X1 U48 ( .A1(\mem[2][2] ), .A2(n671), .ZN(n668) );
  OAI21_X1 U49 ( .B1(n407), .B2(n671), .A(n667), .ZN(n519) );
  NAND2_X1 U50 ( .A1(\mem[2][3] ), .A2(n671), .ZN(n667) );
  OAI21_X1 U51 ( .B1(n406), .B2(n671), .A(n666), .ZN(n518) );
  NAND2_X1 U52 ( .A1(\mem[2][4] ), .A2(n671), .ZN(n666) );
  OAI21_X1 U53 ( .B1(n405), .B2(n671), .A(n665), .ZN(n517) );
  NAND2_X1 U54 ( .A1(\mem[2][5] ), .A2(n671), .ZN(n665) );
  OAI21_X1 U55 ( .B1(n404), .B2(n671), .A(n664), .ZN(n516) );
  NAND2_X1 U56 ( .A1(\mem[2][6] ), .A2(n671), .ZN(n664) );
  OAI21_X1 U57 ( .B1(n403), .B2(n671), .A(n663), .ZN(n515) );
  NAND2_X1 U58 ( .A1(\mem[2][7] ), .A2(n671), .ZN(n663) );
  OAI21_X1 U59 ( .B1(n410), .B2(n661), .A(n660), .ZN(n514) );
  NAND2_X1 U60 ( .A1(\mem[3][0] ), .A2(n661), .ZN(n660) );
  OAI21_X1 U61 ( .B1(n409), .B2(n661), .A(n659), .ZN(n513) );
  NAND2_X1 U62 ( .A1(\mem[3][1] ), .A2(n661), .ZN(n659) );
  OAI21_X1 U63 ( .B1(n408), .B2(n661), .A(n658), .ZN(n512) );
  NAND2_X1 U64 ( .A1(\mem[3][2] ), .A2(n661), .ZN(n658) );
  OAI21_X1 U65 ( .B1(n407), .B2(n661), .A(n657), .ZN(n511) );
  NAND2_X1 U66 ( .A1(\mem[3][3] ), .A2(n661), .ZN(n657) );
  OAI21_X1 U67 ( .B1(n406), .B2(n661), .A(n656), .ZN(n510) );
  NAND2_X1 U68 ( .A1(\mem[3][4] ), .A2(n661), .ZN(n656) );
  OAI21_X1 U69 ( .B1(n405), .B2(n661), .A(n655), .ZN(n509) );
  NAND2_X1 U70 ( .A1(\mem[3][5] ), .A2(n661), .ZN(n655) );
  OAI21_X1 U71 ( .B1(n404), .B2(n661), .A(n654), .ZN(n508) );
  NAND2_X1 U72 ( .A1(\mem[3][6] ), .A2(n661), .ZN(n654) );
  OAI21_X1 U73 ( .B1(n403), .B2(n661), .A(n653), .ZN(n507) );
  NAND2_X1 U74 ( .A1(\mem[3][7] ), .A2(n661), .ZN(n653) );
  NOR2_X1 U75 ( .A1(n402), .A2(N13), .ZN(n623) );
  INV_X1 U76 ( .A(wr_en), .ZN(n402) );
  OAI21_X1 U77 ( .B1(n410), .B2(n681), .A(n680), .ZN(n530) );
  NAND2_X1 U78 ( .A1(\mem[1][0] ), .A2(n681), .ZN(n680) );
  OAI21_X1 U79 ( .B1(n409), .B2(n681), .A(n679), .ZN(n529) );
  NAND2_X1 U80 ( .A1(\mem[1][1] ), .A2(n681), .ZN(n679) );
  OAI21_X1 U81 ( .B1(n408), .B2(n681), .A(n678), .ZN(n528) );
  NAND2_X1 U82 ( .A1(\mem[1][2] ), .A2(n681), .ZN(n678) );
  OAI21_X1 U83 ( .B1(n407), .B2(n681), .A(n677), .ZN(n527) );
  NAND2_X1 U84 ( .A1(\mem[1][3] ), .A2(n681), .ZN(n677) );
  OAI21_X1 U85 ( .B1(n406), .B2(n681), .A(n676), .ZN(n526) );
  NAND2_X1 U86 ( .A1(\mem[1][4] ), .A2(n681), .ZN(n676) );
  OAI21_X1 U87 ( .B1(n405), .B2(n681), .A(n675), .ZN(n525) );
  NAND2_X1 U88 ( .A1(\mem[1][5] ), .A2(n681), .ZN(n675) );
  OAI21_X1 U89 ( .B1(n404), .B2(n681), .A(n674), .ZN(n524) );
  NAND2_X1 U90 ( .A1(\mem[1][6] ), .A2(n681), .ZN(n674) );
  OAI21_X1 U91 ( .B1(n403), .B2(n681), .A(n673), .ZN(n523) );
  NAND2_X1 U92 ( .A1(\mem[1][7] ), .A2(n681), .ZN(n673) );
  OAI21_X1 U93 ( .B1(n410), .B2(n652), .A(n651), .ZN(n506) );
  NAND2_X1 U94 ( .A1(\mem[4][0] ), .A2(n652), .ZN(n651) );
  OAI21_X1 U95 ( .B1(n409), .B2(n652), .A(n650), .ZN(n505) );
  NAND2_X1 U96 ( .A1(\mem[4][1] ), .A2(n652), .ZN(n650) );
  OAI21_X1 U97 ( .B1(n408), .B2(n652), .A(n649), .ZN(n504) );
  NAND2_X1 U98 ( .A1(\mem[4][2] ), .A2(n652), .ZN(n649) );
  OAI21_X1 U99 ( .B1(n407), .B2(n652), .A(n648), .ZN(n503) );
  NAND2_X1 U100 ( .A1(\mem[4][3] ), .A2(n652), .ZN(n648) );
  OAI21_X1 U101 ( .B1(n406), .B2(n652), .A(n647), .ZN(n502) );
  NAND2_X1 U102 ( .A1(\mem[4][4] ), .A2(n652), .ZN(n647) );
  OAI21_X1 U103 ( .B1(n405), .B2(n652), .A(n646), .ZN(n501) );
  NAND2_X1 U104 ( .A1(\mem[4][5] ), .A2(n652), .ZN(n646) );
  OAI21_X1 U105 ( .B1(n404), .B2(n652), .A(n645), .ZN(n500) );
  NAND2_X1 U106 ( .A1(\mem[4][6] ), .A2(n652), .ZN(n645) );
  OAI21_X1 U107 ( .B1(n403), .B2(n652), .A(n644), .ZN(n499) );
  NAND2_X1 U108 ( .A1(\mem[4][7] ), .A2(n652), .ZN(n644) );
  OAI21_X1 U109 ( .B1(n410), .B2(n642), .A(n641), .ZN(n498) );
  NAND2_X1 U110 ( .A1(\mem[5][0] ), .A2(n642), .ZN(n641) );
  OAI21_X1 U111 ( .B1(n409), .B2(n642), .A(n640), .ZN(n497) );
  NAND2_X1 U112 ( .A1(\mem[5][1] ), .A2(n642), .ZN(n640) );
  OAI21_X1 U113 ( .B1(n408), .B2(n642), .A(n639), .ZN(n496) );
  NAND2_X1 U114 ( .A1(\mem[5][2] ), .A2(n642), .ZN(n639) );
  OAI21_X1 U115 ( .B1(n407), .B2(n642), .A(n638), .ZN(n495) );
  NAND2_X1 U116 ( .A1(\mem[5][3] ), .A2(n642), .ZN(n638) );
  OAI21_X1 U117 ( .B1(n406), .B2(n642), .A(n637), .ZN(n494) );
  NAND2_X1 U118 ( .A1(\mem[5][4] ), .A2(n642), .ZN(n637) );
  OAI21_X1 U119 ( .B1(n405), .B2(n642), .A(n636), .ZN(n493) );
  NAND2_X1 U120 ( .A1(\mem[5][5] ), .A2(n642), .ZN(n636) );
  OAI21_X1 U121 ( .B1(n404), .B2(n642), .A(n635), .ZN(n492) );
  NAND2_X1 U122 ( .A1(\mem[5][6] ), .A2(n642), .ZN(n635) );
  OAI21_X1 U123 ( .B1(n403), .B2(n642), .A(n634), .ZN(n491) );
  NAND2_X1 U124 ( .A1(\mem[5][7] ), .A2(n642), .ZN(n634) );
  OAI21_X1 U125 ( .B1(n410), .B2(n633), .A(n632), .ZN(n490) );
  NAND2_X1 U126 ( .A1(\mem[6][0] ), .A2(n633), .ZN(n632) );
  OAI21_X1 U127 ( .B1(n409), .B2(n633), .A(n631), .ZN(n489) );
  NAND2_X1 U128 ( .A1(\mem[6][1] ), .A2(n633), .ZN(n631) );
  OAI21_X1 U129 ( .B1(n408), .B2(n633), .A(n630), .ZN(n488) );
  NAND2_X1 U130 ( .A1(\mem[6][2] ), .A2(n633), .ZN(n630) );
  OAI21_X1 U131 ( .B1(n407), .B2(n633), .A(n629), .ZN(n487) );
  NAND2_X1 U132 ( .A1(\mem[6][3] ), .A2(n633), .ZN(n629) );
  OAI21_X1 U133 ( .B1(n406), .B2(n633), .A(n628), .ZN(n486) );
  NAND2_X1 U134 ( .A1(\mem[6][4] ), .A2(n633), .ZN(n628) );
  OAI21_X1 U135 ( .B1(n405), .B2(n633), .A(n627), .ZN(n485) );
  NAND2_X1 U136 ( .A1(\mem[6][5] ), .A2(n633), .ZN(n627) );
  OAI21_X1 U137 ( .B1(n404), .B2(n633), .A(n626), .ZN(n484) );
  NAND2_X1 U138 ( .A1(\mem[6][6] ), .A2(n633), .ZN(n626) );
  OAI21_X1 U139 ( .B1(n403), .B2(n633), .A(n625), .ZN(n483) );
  NAND2_X1 U140 ( .A1(\mem[6][7] ), .A2(n633), .ZN(n625) );
  OAI21_X1 U141 ( .B1(n410), .B2(n622), .A(n621), .ZN(n482) );
  NAND2_X1 U142 ( .A1(\mem[7][0] ), .A2(n622), .ZN(n621) );
  OAI21_X1 U143 ( .B1(n409), .B2(n622), .A(n620), .ZN(n481) );
  NAND2_X1 U144 ( .A1(\mem[7][1] ), .A2(n622), .ZN(n620) );
  OAI21_X1 U145 ( .B1(n408), .B2(n622), .A(n619), .ZN(n480) );
  NAND2_X1 U146 ( .A1(\mem[7][2] ), .A2(n622), .ZN(n619) );
  OAI21_X1 U147 ( .B1(n407), .B2(n622), .A(n618), .ZN(n479) );
  NAND2_X1 U148 ( .A1(\mem[7][3] ), .A2(n622), .ZN(n618) );
  OAI21_X1 U149 ( .B1(n406), .B2(n622), .A(n617), .ZN(n478) );
  NAND2_X1 U150 ( .A1(\mem[7][4] ), .A2(n622), .ZN(n617) );
  OAI21_X1 U151 ( .B1(n405), .B2(n622), .A(n616), .ZN(n477) );
  NAND2_X1 U152 ( .A1(\mem[7][5] ), .A2(n622), .ZN(n616) );
  OAI21_X1 U153 ( .B1(n404), .B2(n622), .A(n615), .ZN(n476) );
  NAND2_X1 U154 ( .A1(\mem[7][6] ), .A2(n622), .ZN(n615) );
  OAI21_X1 U155 ( .B1(n403), .B2(n622), .A(n614), .ZN(n475) );
  NAND2_X1 U156 ( .A1(\mem[7][7] ), .A2(n622), .ZN(n614) );
  OAI21_X1 U157 ( .B1(n410), .B2(n613), .A(n612), .ZN(n474) );
  NAND2_X1 U158 ( .A1(\mem[8][0] ), .A2(n613), .ZN(n612) );
  OAI21_X1 U159 ( .B1(n409), .B2(n613), .A(n611), .ZN(n473) );
  NAND2_X1 U160 ( .A1(\mem[8][1] ), .A2(n613), .ZN(n611) );
  OAI21_X1 U161 ( .B1(n408), .B2(n613), .A(n610), .ZN(n472) );
  NAND2_X1 U162 ( .A1(\mem[8][2] ), .A2(n613), .ZN(n610) );
  OAI21_X1 U163 ( .B1(n407), .B2(n613), .A(n609), .ZN(n471) );
  NAND2_X1 U164 ( .A1(\mem[8][3] ), .A2(n613), .ZN(n609) );
  OAI21_X1 U165 ( .B1(n406), .B2(n613), .A(n608), .ZN(n470) );
  NAND2_X1 U166 ( .A1(\mem[8][4] ), .A2(n613), .ZN(n608) );
  OAI21_X1 U167 ( .B1(n405), .B2(n613), .A(n607), .ZN(n469) );
  NAND2_X1 U168 ( .A1(\mem[8][5] ), .A2(n613), .ZN(n607) );
  OAI21_X1 U169 ( .B1(n404), .B2(n613), .A(n606), .ZN(n468) );
  NAND2_X1 U170 ( .A1(\mem[8][6] ), .A2(n613), .ZN(n606) );
  OAI21_X1 U171 ( .B1(n403), .B2(n613), .A(n605), .ZN(n467) );
  NAND2_X1 U172 ( .A1(\mem[8][7] ), .A2(n613), .ZN(n605) );
  OAI21_X1 U173 ( .B1(n410), .B2(n603), .A(n602), .ZN(n466) );
  NAND2_X1 U174 ( .A1(\mem[9][0] ), .A2(n603), .ZN(n602) );
  OAI21_X1 U175 ( .B1(n409), .B2(n603), .A(n601), .ZN(n465) );
  NAND2_X1 U176 ( .A1(\mem[9][1] ), .A2(n603), .ZN(n601) );
  OAI21_X1 U177 ( .B1(n408), .B2(n603), .A(n600), .ZN(n464) );
  NAND2_X1 U178 ( .A1(\mem[9][2] ), .A2(n603), .ZN(n600) );
  OAI21_X1 U179 ( .B1(n407), .B2(n603), .A(n599), .ZN(n463) );
  NAND2_X1 U180 ( .A1(\mem[9][3] ), .A2(n603), .ZN(n599) );
  OAI21_X1 U181 ( .B1(n406), .B2(n603), .A(n598), .ZN(n462) );
  NAND2_X1 U182 ( .A1(\mem[9][4] ), .A2(n603), .ZN(n598) );
  OAI21_X1 U183 ( .B1(n405), .B2(n603), .A(n597), .ZN(n461) );
  NAND2_X1 U184 ( .A1(\mem[9][5] ), .A2(n603), .ZN(n597) );
  OAI21_X1 U185 ( .B1(n404), .B2(n603), .A(n596), .ZN(n460) );
  NAND2_X1 U186 ( .A1(\mem[9][6] ), .A2(n603), .ZN(n596) );
  OAI21_X1 U187 ( .B1(n403), .B2(n603), .A(n595), .ZN(n459) );
  NAND2_X1 U188 ( .A1(\mem[9][7] ), .A2(n603), .ZN(n595) );
  OAI21_X1 U189 ( .B1(n410), .B2(n593), .A(n592), .ZN(n458) );
  NAND2_X1 U190 ( .A1(\mem[10][0] ), .A2(n593), .ZN(n592) );
  OAI21_X1 U191 ( .B1(n409), .B2(n593), .A(n591), .ZN(n457) );
  NAND2_X1 U192 ( .A1(\mem[10][1] ), .A2(n593), .ZN(n591) );
  OAI21_X1 U193 ( .B1(n408), .B2(n593), .A(n590), .ZN(n456) );
  NAND2_X1 U194 ( .A1(\mem[10][2] ), .A2(n593), .ZN(n590) );
  OAI21_X1 U195 ( .B1(n407), .B2(n593), .A(n589), .ZN(n455) );
  NAND2_X1 U196 ( .A1(\mem[10][3] ), .A2(n593), .ZN(n589) );
  OAI21_X1 U197 ( .B1(n406), .B2(n593), .A(n588), .ZN(n454) );
  NAND2_X1 U198 ( .A1(\mem[10][4] ), .A2(n593), .ZN(n588) );
  OAI21_X1 U199 ( .B1(n405), .B2(n593), .A(n587), .ZN(n453) );
  NAND2_X1 U200 ( .A1(\mem[10][5] ), .A2(n593), .ZN(n587) );
  OAI21_X1 U201 ( .B1(n404), .B2(n593), .A(n586), .ZN(n452) );
  NAND2_X1 U202 ( .A1(\mem[10][6] ), .A2(n593), .ZN(n586) );
  OAI21_X1 U203 ( .B1(n403), .B2(n593), .A(n585), .ZN(n451) );
  NAND2_X1 U204 ( .A1(\mem[10][7] ), .A2(n593), .ZN(n585) );
  OAI21_X1 U205 ( .B1(n410), .B2(n584), .A(n583), .ZN(n450) );
  NAND2_X1 U206 ( .A1(\mem[11][0] ), .A2(n584), .ZN(n583) );
  OAI21_X1 U207 ( .B1(n409), .B2(n584), .A(n582), .ZN(n449) );
  NAND2_X1 U208 ( .A1(\mem[11][1] ), .A2(n584), .ZN(n582) );
  OAI21_X1 U209 ( .B1(n408), .B2(n584), .A(n581), .ZN(n448) );
  NAND2_X1 U210 ( .A1(\mem[11][2] ), .A2(n584), .ZN(n581) );
  OAI21_X1 U211 ( .B1(n407), .B2(n584), .A(n580), .ZN(n447) );
  NAND2_X1 U212 ( .A1(\mem[11][3] ), .A2(n584), .ZN(n580) );
  OAI21_X1 U213 ( .B1(n406), .B2(n584), .A(n579), .ZN(n446) );
  NAND2_X1 U214 ( .A1(\mem[11][4] ), .A2(n584), .ZN(n579) );
  OAI21_X1 U215 ( .B1(n405), .B2(n584), .A(n578), .ZN(n445) );
  NAND2_X1 U216 ( .A1(\mem[11][5] ), .A2(n584), .ZN(n578) );
  OAI21_X1 U217 ( .B1(n404), .B2(n584), .A(n577), .ZN(n444) );
  NAND2_X1 U218 ( .A1(\mem[11][6] ), .A2(n584), .ZN(n577) );
  OAI21_X1 U219 ( .B1(n403), .B2(n584), .A(n576), .ZN(n443) );
  NAND2_X1 U220 ( .A1(\mem[11][7] ), .A2(n584), .ZN(n576) );
  OAI21_X1 U221 ( .B1(n410), .B2(n575), .A(n574), .ZN(n442) );
  NAND2_X1 U222 ( .A1(\mem[12][0] ), .A2(n575), .ZN(n574) );
  OAI21_X1 U223 ( .B1(n409), .B2(n575), .A(n573), .ZN(n441) );
  NAND2_X1 U224 ( .A1(\mem[12][1] ), .A2(n575), .ZN(n573) );
  OAI21_X1 U225 ( .B1(n408), .B2(n575), .A(n572), .ZN(n440) );
  NAND2_X1 U226 ( .A1(\mem[12][2] ), .A2(n575), .ZN(n572) );
  OAI21_X1 U227 ( .B1(n407), .B2(n575), .A(n571), .ZN(n439) );
  NAND2_X1 U228 ( .A1(\mem[12][3] ), .A2(n575), .ZN(n571) );
  OAI21_X1 U229 ( .B1(n406), .B2(n575), .A(n570), .ZN(n438) );
  NAND2_X1 U230 ( .A1(\mem[12][4] ), .A2(n575), .ZN(n570) );
  OAI21_X1 U231 ( .B1(n405), .B2(n575), .A(n569), .ZN(n437) );
  NAND2_X1 U232 ( .A1(\mem[12][5] ), .A2(n575), .ZN(n569) );
  OAI21_X1 U233 ( .B1(n404), .B2(n575), .A(n568), .ZN(n436) );
  NAND2_X1 U234 ( .A1(\mem[12][6] ), .A2(n575), .ZN(n568) );
  OAI21_X1 U235 ( .B1(n403), .B2(n575), .A(n567), .ZN(n435) );
  NAND2_X1 U236 ( .A1(\mem[12][7] ), .A2(n575), .ZN(n567) );
  OAI21_X1 U237 ( .B1(n410), .B2(n566), .A(n565), .ZN(n434) );
  NAND2_X1 U238 ( .A1(\mem[13][0] ), .A2(n566), .ZN(n565) );
  OAI21_X1 U239 ( .B1(n409), .B2(n566), .A(n564), .ZN(n433) );
  NAND2_X1 U240 ( .A1(\mem[13][1] ), .A2(n566), .ZN(n564) );
  OAI21_X1 U241 ( .B1(n408), .B2(n566), .A(n563), .ZN(n432) );
  NAND2_X1 U242 ( .A1(\mem[13][2] ), .A2(n566), .ZN(n563) );
  OAI21_X1 U243 ( .B1(n407), .B2(n566), .A(n562), .ZN(n431) );
  NAND2_X1 U244 ( .A1(\mem[13][3] ), .A2(n566), .ZN(n562) );
  OAI21_X1 U245 ( .B1(n406), .B2(n566), .A(n561), .ZN(n430) );
  NAND2_X1 U246 ( .A1(\mem[13][4] ), .A2(n566), .ZN(n561) );
  OAI21_X1 U247 ( .B1(n405), .B2(n566), .A(n560), .ZN(n429) );
  NAND2_X1 U248 ( .A1(\mem[13][5] ), .A2(n566), .ZN(n560) );
  OAI21_X1 U249 ( .B1(n404), .B2(n566), .A(n559), .ZN(n428) );
  NAND2_X1 U250 ( .A1(\mem[13][6] ), .A2(n566), .ZN(n559) );
  OAI21_X1 U251 ( .B1(n403), .B2(n566), .A(n558), .ZN(n427) );
  NAND2_X1 U252 ( .A1(\mem[13][7] ), .A2(n566), .ZN(n558) );
  OAI21_X1 U253 ( .B1(n410), .B2(n557), .A(n556), .ZN(n426) );
  NAND2_X1 U254 ( .A1(\mem[14][0] ), .A2(n557), .ZN(n556) );
  OAI21_X1 U255 ( .B1(n409), .B2(n557), .A(n555), .ZN(n425) );
  NAND2_X1 U256 ( .A1(\mem[14][1] ), .A2(n557), .ZN(n555) );
  OAI21_X1 U257 ( .B1(n408), .B2(n557), .A(n554), .ZN(n424) );
  NAND2_X1 U258 ( .A1(\mem[14][2] ), .A2(n557), .ZN(n554) );
  OAI21_X1 U259 ( .B1(n407), .B2(n557), .A(n553), .ZN(n423) );
  NAND2_X1 U260 ( .A1(\mem[14][3] ), .A2(n557), .ZN(n553) );
  OAI21_X1 U261 ( .B1(n406), .B2(n557), .A(n552), .ZN(n422) );
  NAND2_X1 U262 ( .A1(\mem[14][4] ), .A2(n557), .ZN(n552) );
  OAI21_X1 U263 ( .B1(n405), .B2(n557), .A(n551), .ZN(n421) );
  NAND2_X1 U264 ( .A1(\mem[14][5] ), .A2(n557), .ZN(n551) );
  OAI21_X1 U265 ( .B1(n404), .B2(n557), .A(n550), .ZN(n420) );
  NAND2_X1 U266 ( .A1(\mem[14][6] ), .A2(n557), .ZN(n550) );
  OAI21_X1 U267 ( .B1(n403), .B2(n557), .A(n549), .ZN(n419) );
  NAND2_X1 U268 ( .A1(\mem[14][7] ), .A2(n557), .ZN(n549) );
  OAI21_X1 U269 ( .B1(n410), .B2(n547), .A(n546), .ZN(n418) );
  NAND2_X1 U270 ( .A1(\mem[15][0] ), .A2(n547), .ZN(n546) );
  OAI21_X1 U271 ( .B1(n409), .B2(n547), .A(n545), .ZN(n417) );
  NAND2_X1 U272 ( .A1(\mem[15][1] ), .A2(n547), .ZN(n545) );
  OAI21_X1 U273 ( .B1(n408), .B2(n547), .A(n544), .ZN(n416) );
  NAND2_X1 U274 ( .A1(\mem[15][2] ), .A2(n547), .ZN(n544) );
  OAI21_X1 U275 ( .B1(n407), .B2(n547), .A(n543), .ZN(n415) );
  NAND2_X1 U276 ( .A1(\mem[15][3] ), .A2(n547), .ZN(n543) );
  OAI21_X1 U277 ( .B1(n406), .B2(n547), .A(n542), .ZN(n414) );
  NAND2_X1 U278 ( .A1(\mem[15][4] ), .A2(n547), .ZN(n542) );
  OAI21_X1 U279 ( .B1(n405), .B2(n547), .A(n541), .ZN(n413) );
  NAND2_X1 U280 ( .A1(\mem[15][5] ), .A2(n547), .ZN(n541) );
  OAI21_X1 U281 ( .B1(n404), .B2(n547), .A(n540), .ZN(n412) );
  NAND2_X1 U282 ( .A1(\mem[15][6] ), .A2(n547), .ZN(n540) );
  OAI21_X1 U283 ( .B1(n403), .B2(n547), .A(n539), .ZN(n411) );
  NAND2_X1 U284 ( .A1(\mem[15][7] ), .A2(n547), .ZN(n539) );
  AND2_X1 U285 ( .A1(N13), .A2(wr_en), .ZN(n548) );
  NOR2_X1 U286 ( .A1(N11), .A2(N12), .ZN(n683) );
  NOR2_X1 U287 ( .A1(n401), .A2(N12), .ZN(n662) );
  AND2_X1 U288 ( .A1(N12), .A2(n401), .ZN(n643) );
  AND2_X1 U289 ( .A1(N12), .A2(N11), .ZN(n624) );
  INV_X1 U290 ( .A(data_in[0]), .ZN(n410) );
  INV_X1 U291 ( .A(data_in[1]), .ZN(n409) );
  INV_X1 U292 ( .A(data_in[2]), .ZN(n408) );
  INV_X1 U293 ( .A(data_in[3]), .ZN(n407) );
  INV_X1 U294 ( .A(data_in[4]), .ZN(n406) );
  INV_X1 U295 ( .A(data_in[5]), .ZN(n405) );
  INV_X1 U296 ( .A(data_in[6]), .ZN(n404) );
  INV_X1 U297 ( .A(data_in[7]), .ZN(n403) );
  MUX2_X1 U298 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(N10), .Z(n2) );
  MUX2_X1 U299 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(N10), .Z(n3) );
  MUX2_X1 U300 ( .A(n3), .B(n2), .S(N11), .Z(n4) );
  MUX2_X1 U301 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(N10), .Z(n5) );
  MUX2_X1 U302 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n6) );
  MUX2_X1 U303 ( .A(n6), .B(n5), .S(N11), .Z(n7) );
  MUX2_X1 U304 ( .A(n7), .B(n4), .S(N12), .Z(n8) );
  MUX2_X1 U305 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n397), .Z(n9) );
  MUX2_X1 U306 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n397), .Z(n10) );
  MUX2_X1 U307 ( .A(n10), .B(n9), .S(N11), .Z(n11) );
  MUX2_X1 U308 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n397), .Z(n294) );
  MUX2_X1 U309 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n397), .Z(n295) );
  MUX2_X1 U310 ( .A(n295), .B(n294), .S(N11), .Z(n296) );
  MUX2_X1 U311 ( .A(n296), .B(n11), .S(N12), .Z(n297) );
  MUX2_X1 U312 ( .A(n297), .B(n8), .S(N13), .Z(N21) );
  MUX2_X1 U313 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n397), .Z(n298) );
  MUX2_X1 U314 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n397), .Z(n299) );
  MUX2_X1 U315 ( .A(n299), .B(n298), .S(N11), .Z(n300) );
  MUX2_X1 U316 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n397), .Z(n301) );
  MUX2_X1 U317 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n397), .Z(n302) );
  MUX2_X1 U318 ( .A(n302), .B(n301), .S(N11), .Z(n303) );
  MUX2_X1 U319 ( .A(n303), .B(n300), .S(N12), .Z(n304) );
  MUX2_X1 U320 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n397), .Z(n305) );
  MUX2_X1 U321 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n397), .Z(n306) );
  MUX2_X1 U322 ( .A(n306), .B(n305), .S(N11), .Z(n307) );
  MUX2_X1 U323 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n397), .Z(n308) );
  MUX2_X1 U324 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n397), .Z(n309) );
  MUX2_X1 U325 ( .A(n309), .B(n308), .S(N11), .Z(n310) );
  MUX2_X1 U326 ( .A(n310), .B(n307), .S(N12), .Z(n311) );
  MUX2_X1 U327 ( .A(n311), .B(n304), .S(N13), .Z(N20) );
  MUX2_X1 U328 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n398), .Z(n312) );
  MUX2_X1 U329 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n398), .Z(n313) );
  MUX2_X1 U330 ( .A(n313), .B(n312), .S(n396), .Z(n314) );
  MUX2_X1 U331 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n398), .Z(n315) );
  MUX2_X1 U332 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n398), .Z(n316) );
  MUX2_X1 U333 ( .A(n316), .B(n315), .S(n396), .Z(n317) );
  MUX2_X1 U334 ( .A(n317), .B(n314), .S(N12), .Z(n318) );
  MUX2_X1 U335 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n398), .Z(n319) );
  MUX2_X1 U336 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n398), .Z(n320) );
  MUX2_X1 U337 ( .A(n320), .B(n319), .S(n396), .Z(n321) );
  MUX2_X1 U338 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n398), .Z(n322) );
  MUX2_X1 U339 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n398), .Z(n323) );
  MUX2_X1 U340 ( .A(n323), .B(n322), .S(n396), .Z(n324) );
  MUX2_X1 U341 ( .A(n324), .B(n321), .S(N12), .Z(n325) );
  MUX2_X1 U342 ( .A(n325), .B(n318), .S(N13), .Z(N19) );
  MUX2_X1 U343 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n398), .Z(n326) );
  MUX2_X1 U344 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n398), .Z(n327) );
  MUX2_X1 U345 ( .A(n327), .B(n326), .S(n396), .Z(n328) );
  MUX2_X1 U346 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n398), .Z(n329) );
  MUX2_X1 U347 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n398), .Z(n330) );
  MUX2_X1 U348 ( .A(n330), .B(n329), .S(n396), .Z(n331) );
  MUX2_X1 U349 ( .A(n331), .B(n328), .S(N12), .Z(n332) );
  MUX2_X1 U350 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n399), .Z(n333) );
  MUX2_X1 U351 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n399), .Z(n334) );
  MUX2_X1 U352 ( .A(n334), .B(n333), .S(n396), .Z(n335) );
  MUX2_X1 U353 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n399), .Z(n336) );
  MUX2_X1 U354 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n399), .Z(n337) );
  MUX2_X1 U355 ( .A(n337), .B(n336), .S(n396), .Z(n338) );
  MUX2_X1 U356 ( .A(n338), .B(n335), .S(N12), .Z(n339) );
  MUX2_X1 U357 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n399), .Z(n340) );
  MUX2_X1 U358 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n399), .Z(n341) );
  MUX2_X1 U359 ( .A(n341), .B(n340), .S(n396), .Z(n342) );
  MUX2_X1 U360 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n399), .Z(n343) );
  MUX2_X1 U361 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n399), .Z(n344) );
  MUX2_X1 U362 ( .A(n344), .B(n343), .S(n396), .Z(n345) );
  MUX2_X1 U363 ( .A(n345), .B(n342), .S(N12), .Z(n346) );
  MUX2_X1 U364 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n399), .Z(n347) );
  MUX2_X1 U365 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n399), .Z(n348) );
  MUX2_X1 U366 ( .A(n348), .B(n347), .S(n396), .Z(n349) );
  MUX2_X1 U367 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n399), .Z(n350) );
  MUX2_X1 U368 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n399), .Z(n351) );
  MUX2_X1 U369 ( .A(n351), .B(n350), .S(n396), .Z(n352) );
  MUX2_X1 U370 ( .A(n352), .B(n349), .S(N12), .Z(n353) );
  MUX2_X1 U371 ( .A(n353), .B(n346), .S(N13), .Z(N17) );
  MUX2_X1 U372 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n397), .Z(n354) );
  MUX2_X1 U373 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n399), .Z(n355) );
  MUX2_X1 U374 ( .A(n355), .B(n354), .S(N11), .Z(n356) );
  MUX2_X1 U375 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(N10), .Z(n357) );
  MUX2_X1 U376 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n399), .Z(n358) );
  MUX2_X1 U377 ( .A(n358), .B(n357), .S(N11), .Z(n359) );
  MUX2_X1 U378 ( .A(n359), .B(n356), .S(N12), .Z(n360) );
  MUX2_X1 U379 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n397), .Z(n361) );
  MUX2_X1 U380 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n397), .Z(n362) );
  MUX2_X1 U381 ( .A(n362), .B(n361), .S(N11), .Z(n363) );
  MUX2_X1 U382 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n397), .Z(n364) );
  MUX2_X1 U383 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n399), .Z(n365) );
  MUX2_X1 U384 ( .A(n365), .B(n364), .S(N11), .Z(n366) );
  MUX2_X1 U385 ( .A(n366), .B(n363), .S(N12), .Z(n367) );
  MUX2_X1 U386 ( .A(n367), .B(n360), .S(N13), .Z(N16) );
  MUX2_X1 U387 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n399), .Z(n368) );
  MUX2_X1 U388 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n398), .Z(n369) );
  MUX2_X1 U389 ( .A(n369), .B(n368), .S(N11), .Z(n370) );
  MUX2_X1 U390 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n398), .Z(n371) );
  MUX2_X1 U391 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n398), .Z(n372) );
  MUX2_X1 U392 ( .A(n372), .B(n371), .S(N11), .Z(n373) );
  MUX2_X1 U393 ( .A(n373), .B(n370), .S(N12), .Z(n374) );
  MUX2_X1 U394 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n375) );
  MUX2_X1 U395 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n376) );
  MUX2_X1 U396 ( .A(n376), .B(n375), .S(N11), .Z(n377) );
  MUX2_X1 U397 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n378) );
  MUX2_X1 U398 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n379) );
  MUX2_X1 U399 ( .A(n379), .B(n378), .S(n396), .Z(n380) );
  MUX2_X1 U400 ( .A(n380), .B(n377), .S(N12), .Z(n381) );
  MUX2_X1 U401 ( .A(n381), .B(n374), .S(N13), .Z(N15) );
  MUX2_X1 U402 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(N10), .Z(n382) );
  MUX2_X1 U403 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n383) );
  MUX2_X1 U404 ( .A(n383), .B(n382), .S(N11), .Z(n384) );
  MUX2_X1 U405 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(N10), .Z(n385) );
  MUX2_X1 U406 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n386) );
  MUX2_X1 U407 ( .A(n386), .B(n385), .S(N11), .Z(n387) );
  MUX2_X1 U408 ( .A(n387), .B(n384), .S(N12), .Z(n388) );
  MUX2_X1 U409 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n389) );
  MUX2_X1 U410 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n390) );
  MUX2_X1 U411 ( .A(n390), .B(n389), .S(N11), .Z(n391) );
  MUX2_X1 U412 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n392) );
  MUX2_X1 U413 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n398), .Z(n393) );
  MUX2_X1 U414 ( .A(n393), .B(n392), .S(n396), .Z(n394) );
  MUX2_X1 U415 ( .A(n394), .B(n391), .S(N12), .Z(n395) );
  MUX2_X1 U416 ( .A(n395), .B(n388), .S(N13), .Z(N14) );
  INV_X1 U417 ( .A(N10), .ZN(n400) );
  INV_X1 U418 ( .A(N11), .ZN(n401) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_9 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, N19, N20, N21, n1, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N16), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n412), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n413), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n414), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n415), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n416), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n417), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n418), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n419), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n420), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n421), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n422), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n423), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n424), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n425), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n426), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n427), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n428), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n429), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n430), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n431), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n432), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n433), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n434), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n435), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n436), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n437), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n438), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n439), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n440), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n441), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n442), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n443), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n444), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n445), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n446), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n447), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n448), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n449), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n450), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n451), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n452), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n453), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n454), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n455), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n456), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n457), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n458), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n459), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n460), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n461), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n462), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n463), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n464), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n465), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n466), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n467), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n468), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n469), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n470), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n471), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n472), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n473), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n474), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n475), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n476), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n477), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n478), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n479), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n480), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n481), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n482), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n483), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n484), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n485), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n486), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n487), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n488), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n489), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n490), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n491), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n492), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n493), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n494), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n495), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n496), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n497), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n498), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n499), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n500), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n501), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n502), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n503), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n504), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n505), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n506), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n507), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n508), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n509), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n510), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n511), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n512), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n513), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n514), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n515), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n516), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n517), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n518), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n519), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n520), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n521), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n522), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n523), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n524), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n525), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n526), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n527), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n528), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n529), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n530), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n531), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n532), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n533), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n534), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n535), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n536), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n537), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n538), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n539), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N20), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .QN(n1) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(N10), .Z(n398) );
  BUF_X1 U5 ( .A(N10), .Z(n399) );
  BUF_X1 U6 ( .A(N10), .Z(n400) );
  BUF_X1 U7 ( .A(N11), .Z(n397) );
  NAND2_X1 U8 ( .A1(n663), .A2(n683), .ZN(n672) );
  NAND2_X1 U9 ( .A1(n663), .A2(n673), .ZN(n662) );
  NAND2_X1 U10 ( .A1(n684), .A2(n683), .ZN(n693) );
  NAND2_X1 U11 ( .A1(n673), .A2(n684), .ZN(n682) );
  NAND2_X1 U12 ( .A1(n605), .A2(n684), .ZN(n614) );
  NAND2_X1 U13 ( .A1(n595), .A2(n684), .ZN(n604) );
  NAND2_X1 U14 ( .A1(n605), .A2(n663), .ZN(n594) );
  NAND2_X1 U15 ( .A1(n595), .A2(n663), .ZN(n585) );
  NAND2_X1 U16 ( .A1(n644), .A2(n683), .ZN(n653) );
  NAND2_X1 U17 ( .A1(n644), .A2(n673), .ZN(n643) );
  NAND2_X1 U18 ( .A1(n625), .A2(n683), .ZN(n634) );
  NAND2_X1 U19 ( .A1(n625), .A2(n673), .ZN(n623) );
  NAND2_X1 U20 ( .A1(n605), .A2(n644), .ZN(n576) );
  NAND2_X1 U21 ( .A1(n595), .A2(n644), .ZN(n567) );
  NAND2_X1 U22 ( .A1(n605), .A2(n625), .ZN(n558) );
  NAND2_X1 U23 ( .A1(n595), .A2(n625), .ZN(n548) );
  AND2_X1 U24 ( .A1(n549), .A2(N10), .ZN(n595) );
  AND2_X1 U25 ( .A1(n549), .A2(n401), .ZN(n605) );
  AND2_X1 U26 ( .A1(N10), .A2(n624), .ZN(n673) );
  AND2_X1 U27 ( .A1(n624), .A2(n401), .ZN(n683) );
  OAI21_X1 U28 ( .B1(n693), .B2(n411), .A(n692), .ZN(n539) );
  NAND2_X1 U29 ( .A1(\mem[0][0] ), .A2(n693), .ZN(n692) );
  OAI21_X1 U30 ( .B1(n693), .B2(n410), .A(n691), .ZN(n538) );
  NAND2_X1 U31 ( .A1(\mem[0][1] ), .A2(n693), .ZN(n691) );
  OAI21_X1 U32 ( .B1(n693), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U33 ( .A1(\mem[0][2] ), .A2(n693), .ZN(n690) );
  OAI21_X1 U34 ( .B1(n693), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U35 ( .A1(\mem[0][3] ), .A2(n693), .ZN(n689) );
  OAI21_X1 U36 ( .B1(n693), .B2(n407), .A(n688), .ZN(n535) );
  NAND2_X1 U37 ( .A1(\mem[0][4] ), .A2(n693), .ZN(n688) );
  OAI21_X1 U38 ( .B1(n693), .B2(n406), .A(n687), .ZN(n534) );
  NAND2_X1 U39 ( .A1(\mem[0][5] ), .A2(n693), .ZN(n687) );
  OAI21_X1 U40 ( .B1(n693), .B2(n405), .A(n686), .ZN(n533) );
  NAND2_X1 U41 ( .A1(\mem[0][6] ), .A2(n693), .ZN(n686) );
  OAI21_X1 U42 ( .B1(n693), .B2(n404), .A(n685), .ZN(n532) );
  NAND2_X1 U43 ( .A1(\mem[0][7] ), .A2(n693), .ZN(n685) );
  OAI21_X1 U44 ( .B1(n411), .B2(n672), .A(n671), .ZN(n523) );
  NAND2_X1 U45 ( .A1(\mem[2][0] ), .A2(n672), .ZN(n671) );
  OAI21_X1 U46 ( .B1(n410), .B2(n672), .A(n670), .ZN(n522) );
  NAND2_X1 U47 ( .A1(\mem[2][1] ), .A2(n672), .ZN(n670) );
  OAI21_X1 U48 ( .B1(n409), .B2(n672), .A(n669), .ZN(n521) );
  NAND2_X1 U49 ( .A1(\mem[2][2] ), .A2(n672), .ZN(n669) );
  OAI21_X1 U50 ( .B1(n408), .B2(n672), .A(n668), .ZN(n520) );
  NAND2_X1 U51 ( .A1(\mem[2][3] ), .A2(n672), .ZN(n668) );
  OAI21_X1 U52 ( .B1(n407), .B2(n672), .A(n667), .ZN(n519) );
  NAND2_X1 U53 ( .A1(\mem[2][4] ), .A2(n672), .ZN(n667) );
  OAI21_X1 U54 ( .B1(n406), .B2(n672), .A(n666), .ZN(n518) );
  NAND2_X1 U55 ( .A1(\mem[2][5] ), .A2(n672), .ZN(n666) );
  OAI21_X1 U56 ( .B1(n405), .B2(n672), .A(n665), .ZN(n517) );
  NAND2_X1 U57 ( .A1(\mem[2][6] ), .A2(n672), .ZN(n665) );
  OAI21_X1 U58 ( .B1(n404), .B2(n672), .A(n664), .ZN(n516) );
  NAND2_X1 U59 ( .A1(\mem[2][7] ), .A2(n672), .ZN(n664) );
  OAI21_X1 U60 ( .B1(n411), .B2(n662), .A(n661), .ZN(n515) );
  NAND2_X1 U61 ( .A1(\mem[3][0] ), .A2(n662), .ZN(n661) );
  OAI21_X1 U62 ( .B1(n410), .B2(n662), .A(n660), .ZN(n514) );
  NAND2_X1 U63 ( .A1(\mem[3][1] ), .A2(n662), .ZN(n660) );
  OAI21_X1 U64 ( .B1(n409), .B2(n662), .A(n659), .ZN(n513) );
  NAND2_X1 U65 ( .A1(\mem[3][2] ), .A2(n662), .ZN(n659) );
  OAI21_X1 U66 ( .B1(n408), .B2(n662), .A(n658), .ZN(n512) );
  NAND2_X1 U67 ( .A1(\mem[3][3] ), .A2(n662), .ZN(n658) );
  OAI21_X1 U68 ( .B1(n407), .B2(n662), .A(n657), .ZN(n511) );
  NAND2_X1 U69 ( .A1(\mem[3][4] ), .A2(n662), .ZN(n657) );
  OAI21_X1 U70 ( .B1(n406), .B2(n662), .A(n656), .ZN(n510) );
  NAND2_X1 U71 ( .A1(\mem[3][5] ), .A2(n662), .ZN(n656) );
  OAI21_X1 U72 ( .B1(n405), .B2(n662), .A(n655), .ZN(n509) );
  NAND2_X1 U73 ( .A1(\mem[3][6] ), .A2(n662), .ZN(n655) );
  OAI21_X1 U74 ( .B1(n404), .B2(n662), .A(n654), .ZN(n508) );
  NAND2_X1 U75 ( .A1(\mem[3][7] ), .A2(n662), .ZN(n654) );
  NOR2_X1 U76 ( .A1(n403), .A2(N13), .ZN(n624) );
  INV_X1 U77 ( .A(wr_en), .ZN(n403) );
  OAI21_X1 U78 ( .B1(n411), .B2(n682), .A(n681), .ZN(n531) );
  NAND2_X1 U79 ( .A1(\mem[1][0] ), .A2(n682), .ZN(n681) );
  OAI21_X1 U80 ( .B1(n410), .B2(n682), .A(n680), .ZN(n530) );
  NAND2_X1 U81 ( .A1(\mem[1][1] ), .A2(n682), .ZN(n680) );
  OAI21_X1 U82 ( .B1(n409), .B2(n682), .A(n679), .ZN(n529) );
  NAND2_X1 U83 ( .A1(\mem[1][2] ), .A2(n682), .ZN(n679) );
  OAI21_X1 U84 ( .B1(n408), .B2(n682), .A(n678), .ZN(n528) );
  NAND2_X1 U85 ( .A1(\mem[1][3] ), .A2(n682), .ZN(n678) );
  OAI21_X1 U86 ( .B1(n407), .B2(n682), .A(n677), .ZN(n527) );
  NAND2_X1 U87 ( .A1(\mem[1][4] ), .A2(n682), .ZN(n677) );
  OAI21_X1 U88 ( .B1(n406), .B2(n682), .A(n676), .ZN(n526) );
  NAND2_X1 U89 ( .A1(\mem[1][5] ), .A2(n682), .ZN(n676) );
  OAI21_X1 U90 ( .B1(n405), .B2(n682), .A(n675), .ZN(n525) );
  NAND2_X1 U91 ( .A1(\mem[1][6] ), .A2(n682), .ZN(n675) );
  OAI21_X1 U92 ( .B1(n404), .B2(n682), .A(n674), .ZN(n524) );
  NAND2_X1 U93 ( .A1(\mem[1][7] ), .A2(n682), .ZN(n674) );
  OAI21_X1 U94 ( .B1(n411), .B2(n653), .A(n652), .ZN(n507) );
  NAND2_X1 U95 ( .A1(\mem[4][0] ), .A2(n653), .ZN(n652) );
  OAI21_X1 U96 ( .B1(n410), .B2(n653), .A(n651), .ZN(n506) );
  NAND2_X1 U97 ( .A1(\mem[4][1] ), .A2(n653), .ZN(n651) );
  OAI21_X1 U98 ( .B1(n409), .B2(n653), .A(n650), .ZN(n505) );
  NAND2_X1 U99 ( .A1(\mem[4][2] ), .A2(n653), .ZN(n650) );
  OAI21_X1 U100 ( .B1(n408), .B2(n653), .A(n649), .ZN(n504) );
  NAND2_X1 U101 ( .A1(\mem[4][3] ), .A2(n653), .ZN(n649) );
  OAI21_X1 U102 ( .B1(n407), .B2(n653), .A(n648), .ZN(n503) );
  NAND2_X1 U103 ( .A1(\mem[4][4] ), .A2(n653), .ZN(n648) );
  OAI21_X1 U104 ( .B1(n406), .B2(n653), .A(n647), .ZN(n502) );
  NAND2_X1 U105 ( .A1(\mem[4][5] ), .A2(n653), .ZN(n647) );
  OAI21_X1 U106 ( .B1(n405), .B2(n653), .A(n646), .ZN(n501) );
  NAND2_X1 U107 ( .A1(\mem[4][6] ), .A2(n653), .ZN(n646) );
  OAI21_X1 U108 ( .B1(n404), .B2(n653), .A(n645), .ZN(n500) );
  NAND2_X1 U109 ( .A1(\mem[4][7] ), .A2(n653), .ZN(n645) );
  OAI21_X1 U110 ( .B1(n411), .B2(n643), .A(n642), .ZN(n499) );
  NAND2_X1 U111 ( .A1(\mem[5][0] ), .A2(n643), .ZN(n642) );
  OAI21_X1 U112 ( .B1(n410), .B2(n643), .A(n641), .ZN(n498) );
  NAND2_X1 U113 ( .A1(\mem[5][1] ), .A2(n643), .ZN(n641) );
  OAI21_X1 U114 ( .B1(n409), .B2(n643), .A(n640), .ZN(n497) );
  NAND2_X1 U115 ( .A1(\mem[5][2] ), .A2(n643), .ZN(n640) );
  OAI21_X1 U116 ( .B1(n408), .B2(n643), .A(n639), .ZN(n496) );
  NAND2_X1 U117 ( .A1(\mem[5][3] ), .A2(n643), .ZN(n639) );
  OAI21_X1 U118 ( .B1(n407), .B2(n643), .A(n638), .ZN(n495) );
  NAND2_X1 U119 ( .A1(\mem[5][4] ), .A2(n643), .ZN(n638) );
  OAI21_X1 U120 ( .B1(n406), .B2(n643), .A(n637), .ZN(n494) );
  NAND2_X1 U121 ( .A1(\mem[5][5] ), .A2(n643), .ZN(n637) );
  OAI21_X1 U122 ( .B1(n405), .B2(n643), .A(n636), .ZN(n493) );
  NAND2_X1 U123 ( .A1(\mem[5][6] ), .A2(n643), .ZN(n636) );
  OAI21_X1 U124 ( .B1(n404), .B2(n643), .A(n635), .ZN(n492) );
  NAND2_X1 U125 ( .A1(\mem[5][7] ), .A2(n643), .ZN(n635) );
  OAI21_X1 U126 ( .B1(n411), .B2(n634), .A(n633), .ZN(n491) );
  NAND2_X1 U127 ( .A1(\mem[6][0] ), .A2(n634), .ZN(n633) );
  OAI21_X1 U128 ( .B1(n410), .B2(n634), .A(n632), .ZN(n490) );
  NAND2_X1 U129 ( .A1(\mem[6][1] ), .A2(n634), .ZN(n632) );
  OAI21_X1 U130 ( .B1(n409), .B2(n634), .A(n631), .ZN(n489) );
  NAND2_X1 U131 ( .A1(\mem[6][2] ), .A2(n634), .ZN(n631) );
  OAI21_X1 U132 ( .B1(n408), .B2(n634), .A(n630), .ZN(n488) );
  NAND2_X1 U133 ( .A1(\mem[6][3] ), .A2(n634), .ZN(n630) );
  OAI21_X1 U134 ( .B1(n407), .B2(n634), .A(n629), .ZN(n487) );
  NAND2_X1 U135 ( .A1(\mem[6][4] ), .A2(n634), .ZN(n629) );
  OAI21_X1 U136 ( .B1(n406), .B2(n634), .A(n628), .ZN(n486) );
  NAND2_X1 U137 ( .A1(\mem[6][5] ), .A2(n634), .ZN(n628) );
  OAI21_X1 U138 ( .B1(n405), .B2(n634), .A(n627), .ZN(n485) );
  NAND2_X1 U139 ( .A1(\mem[6][6] ), .A2(n634), .ZN(n627) );
  OAI21_X1 U140 ( .B1(n404), .B2(n634), .A(n626), .ZN(n484) );
  NAND2_X1 U141 ( .A1(\mem[6][7] ), .A2(n634), .ZN(n626) );
  OAI21_X1 U142 ( .B1(n411), .B2(n623), .A(n622), .ZN(n483) );
  NAND2_X1 U143 ( .A1(\mem[7][0] ), .A2(n623), .ZN(n622) );
  OAI21_X1 U144 ( .B1(n410), .B2(n623), .A(n621), .ZN(n482) );
  NAND2_X1 U145 ( .A1(\mem[7][1] ), .A2(n623), .ZN(n621) );
  OAI21_X1 U146 ( .B1(n409), .B2(n623), .A(n620), .ZN(n481) );
  NAND2_X1 U147 ( .A1(\mem[7][2] ), .A2(n623), .ZN(n620) );
  OAI21_X1 U148 ( .B1(n408), .B2(n623), .A(n619), .ZN(n480) );
  NAND2_X1 U149 ( .A1(\mem[7][3] ), .A2(n623), .ZN(n619) );
  OAI21_X1 U150 ( .B1(n407), .B2(n623), .A(n618), .ZN(n479) );
  NAND2_X1 U151 ( .A1(\mem[7][4] ), .A2(n623), .ZN(n618) );
  OAI21_X1 U152 ( .B1(n406), .B2(n623), .A(n617), .ZN(n478) );
  NAND2_X1 U153 ( .A1(\mem[7][5] ), .A2(n623), .ZN(n617) );
  OAI21_X1 U154 ( .B1(n405), .B2(n623), .A(n616), .ZN(n477) );
  NAND2_X1 U155 ( .A1(\mem[7][6] ), .A2(n623), .ZN(n616) );
  OAI21_X1 U156 ( .B1(n404), .B2(n623), .A(n615), .ZN(n476) );
  NAND2_X1 U157 ( .A1(\mem[7][7] ), .A2(n623), .ZN(n615) );
  OAI21_X1 U158 ( .B1(n411), .B2(n614), .A(n613), .ZN(n475) );
  NAND2_X1 U159 ( .A1(\mem[8][0] ), .A2(n614), .ZN(n613) );
  OAI21_X1 U160 ( .B1(n410), .B2(n614), .A(n612), .ZN(n474) );
  NAND2_X1 U161 ( .A1(\mem[8][1] ), .A2(n614), .ZN(n612) );
  OAI21_X1 U162 ( .B1(n409), .B2(n614), .A(n611), .ZN(n473) );
  NAND2_X1 U163 ( .A1(\mem[8][2] ), .A2(n614), .ZN(n611) );
  OAI21_X1 U164 ( .B1(n408), .B2(n614), .A(n610), .ZN(n472) );
  NAND2_X1 U165 ( .A1(\mem[8][3] ), .A2(n614), .ZN(n610) );
  OAI21_X1 U166 ( .B1(n407), .B2(n614), .A(n609), .ZN(n471) );
  NAND2_X1 U167 ( .A1(\mem[8][4] ), .A2(n614), .ZN(n609) );
  OAI21_X1 U168 ( .B1(n406), .B2(n614), .A(n608), .ZN(n470) );
  NAND2_X1 U169 ( .A1(\mem[8][5] ), .A2(n614), .ZN(n608) );
  OAI21_X1 U170 ( .B1(n405), .B2(n614), .A(n607), .ZN(n469) );
  NAND2_X1 U171 ( .A1(\mem[8][6] ), .A2(n614), .ZN(n607) );
  OAI21_X1 U172 ( .B1(n404), .B2(n614), .A(n606), .ZN(n468) );
  NAND2_X1 U173 ( .A1(\mem[8][7] ), .A2(n614), .ZN(n606) );
  OAI21_X1 U174 ( .B1(n411), .B2(n604), .A(n603), .ZN(n467) );
  NAND2_X1 U175 ( .A1(\mem[9][0] ), .A2(n604), .ZN(n603) );
  OAI21_X1 U176 ( .B1(n410), .B2(n604), .A(n602), .ZN(n466) );
  NAND2_X1 U177 ( .A1(\mem[9][1] ), .A2(n604), .ZN(n602) );
  OAI21_X1 U178 ( .B1(n409), .B2(n604), .A(n601), .ZN(n465) );
  NAND2_X1 U179 ( .A1(\mem[9][2] ), .A2(n604), .ZN(n601) );
  OAI21_X1 U180 ( .B1(n408), .B2(n604), .A(n600), .ZN(n464) );
  NAND2_X1 U181 ( .A1(\mem[9][3] ), .A2(n604), .ZN(n600) );
  OAI21_X1 U182 ( .B1(n407), .B2(n604), .A(n599), .ZN(n463) );
  NAND2_X1 U183 ( .A1(\mem[9][4] ), .A2(n604), .ZN(n599) );
  OAI21_X1 U184 ( .B1(n406), .B2(n604), .A(n598), .ZN(n462) );
  NAND2_X1 U185 ( .A1(\mem[9][5] ), .A2(n604), .ZN(n598) );
  OAI21_X1 U186 ( .B1(n405), .B2(n604), .A(n597), .ZN(n461) );
  NAND2_X1 U187 ( .A1(\mem[9][6] ), .A2(n604), .ZN(n597) );
  OAI21_X1 U188 ( .B1(n404), .B2(n604), .A(n596), .ZN(n460) );
  NAND2_X1 U189 ( .A1(\mem[9][7] ), .A2(n604), .ZN(n596) );
  OAI21_X1 U190 ( .B1(n411), .B2(n594), .A(n593), .ZN(n459) );
  NAND2_X1 U191 ( .A1(\mem[10][0] ), .A2(n594), .ZN(n593) );
  OAI21_X1 U192 ( .B1(n410), .B2(n594), .A(n592), .ZN(n458) );
  NAND2_X1 U193 ( .A1(\mem[10][1] ), .A2(n594), .ZN(n592) );
  OAI21_X1 U194 ( .B1(n409), .B2(n594), .A(n591), .ZN(n457) );
  NAND2_X1 U195 ( .A1(\mem[10][2] ), .A2(n594), .ZN(n591) );
  OAI21_X1 U196 ( .B1(n408), .B2(n594), .A(n590), .ZN(n456) );
  NAND2_X1 U197 ( .A1(\mem[10][3] ), .A2(n594), .ZN(n590) );
  OAI21_X1 U198 ( .B1(n407), .B2(n594), .A(n589), .ZN(n455) );
  NAND2_X1 U199 ( .A1(\mem[10][4] ), .A2(n594), .ZN(n589) );
  OAI21_X1 U200 ( .B1(n406), .B2(n594), .A(n588), .ZN(n454) );
  NAND2_X1 U201 ( .A1(\mem[10][5] ), .A2(n594), .ZN(n588) );
  OAI21_X1 U202 ( .B1(n405), .B2(n594), .A(n587), .ZN(n453) );
  NAND2_X1 U203 ( .A1(\mem[10][6] ), .A2(n594), .ZN(n587) );
  OAI21_X1 U204 ( .B1(n404), .B2(n594), .A(n586), .ZN(n452) );
  NAND2_X1 U205 ( .A1(\mem[10][7] ), .A2(n594), .ZN(n586) );
  OAI21_X1 U206 ( .B1(n411), .B2(n585), .A(n584), .ZN(n451) );
  NAND2_X1 U207 ( .A1(\mem[11][0] ), .A2(n585), .ZN(n584) );
  OAI21_X1 U208 ( .B1(n410), .B2(n585), .A(n583), .ZN(n450) );
  NAND2_X1 U209 ( .A1(\mem[11][1] ), .A2(n585), .ZN(n583) );
  OAI21_X1 U210 ( .B1(n409), .B2(n585), .A(n582), .ZN(n449) );
  NAND2_X1 U211 ( .A1(\mem[11][2] ), .A2(n585), .ZN(n582) );
  OAI21_X1 U212 ( .B1(n408), .B2(n585), .A(n581), .ZN(n448) );
  NAND2_X1 U213 ( .A1(\mem[11][3] ), .A2(n585), .ZN(n581) );
  OAI21_X1 U214 ( .B1(n407), .B2(n585), .A(n580), .ZN(n447) );
  NAND2_X1 U215 ( .A1(\mem[11][4] ), .A2(n585), .ZN(n580) );
  OAI21_X1 U216 ( .B1(n406), .B2(n585), .A(n579), .ZN(n446) );
  NAND2_X1 U217 ( .A1(\mem[11][5] ), .A2(n585), .ZN(n579) );
  OAI21_X1 U218 ( .B1(n405), .B2(n585), .A(n578), .ZN(n445) );
  NAND2_X1 U219 ( .A1(\mem[11][6] ), .A2(n585), .ZN(n578) );
  OAI21_X1 U220 ( .B1(n404), .B2(n585), .A(n577), .ZN(n444) );
  NAND2_X1 U221 ( .A1(\mem[11][7] ), .A2(n585), .ZN(n577) );
  OAI21_X1 U222 ( .B1(n411), .B2(n576), .A(n575), .ZN(n443) );
  NAND2_X1 U223 ( .A1(\mem[12][0] ), .A2(n576), .ZN(n575) );
  OAI21_X1 U224 ( .B1(n410), .B2(n576), .A(n574), .ZN(n442) );
  NAND2_X1 U225 ( .A1(\mem[12][1] ), .A2(n576), .ZN(n574) );
  OAI21_X1 U226 ( .B1(n409), .B2(n576), .A(n573), .ZN(n441) );
  NAND2_X1 U227 ( .A1(\mem[12][2] ), .A2(n576), .ZN(n573) );
  OAI21_X1 U228 ( .B1(n408), .B2(n576), .A(n572), .ZN(n440) );
  NAND2_X1 U229 ( .A1(\mem[12][3] ), .A2(n576), .ZN(n572) );
  OAI21_X1 U230 ( .B1(n407), .B2(n576), .A(n571), .ZN(n439) );
  NAND2_X1 U231 ( .A1(\mem[12][4] ), .A2(n576), .ZN(n571) );
  OAI21_X1 U232 ( .B1(n406), .B2(n576), .A(n570), .ZN(n438) );
  NAND2_X1 U233 ( .A1(\mem[12][5] ), .A2(n576), .ZN(n570) );
  OAI21_X1 U234 ( .B1(n405), .B2(n576), .A(n569), .ZN(n437) );
  NAND2_X1 U235 ( .A1(\mem[12][6] ), .A2(n576), .ZN(n569) );
  OAI21_X1 U236 ( .B1(n404), .B2(n576), .A(n568), .ZN(n436) );
  NAND2_X1 U237 ( .A1(\mem[12][7] ), .A2(n576), .ZN(n568) );
  OAI21_X1 U238 ( .B1(n411), .B2(n567), .A(n566), .ZN(n435) );
  NAND2_X1 U239 ( .A1(\mem[13][0] ), .A2(n567), .ZN(n566) );
  OAI21_X1 U240 ( .B1(n410), .B2(n567), .A(n565), .ZN(n434) );
  NAND2_X1 U241 ( .A1(\mem[13][1] ), .A2(n567), .ZN(n565) );
  OAI21_X1 U242 ( .B1(n409), .B2(n567), .A(n564), .ZN(n433) );
  NAND2_X1 U243 ( .A1(\mem[13][2] ), .A2(n567), .ZN(n564) );
  OAI21_X1 U244 ( .B1(n408), .B2(n567), .A(n563), .ZN(n432) );
  NAND2_X1 U245 ( .A1(\mem[13][3] ), .A2(n567), .ZN(n563) );
  OAI21_X1 U246 ( .B1(n407), .B2(n567), .A(n562), .ZN(n431) );
  NAND2_X1 U247 ( .A1(\mem[13][4] ), .A2(n567), .ZN(n562) );
  OAI21_X1 U248 ( .B1(n406), .B2(n567), .A(n561), .ZN(n430) );
  NAND2_X1 U249 ( .A1(\mem[13][5] ), .A2(n567), .ZN(n561) );
  OAI21_X1 U250 ( .B1(n405), .B2(n567), .A(n560), .ZN(n429) );
  NAND2_X1 U251 ( .A1(\mem[13][6] ), .A2(n567), .ZN(n560) );
  OAI21_X1 U252 ( .B1(n404), .B2(n567), .A(n559), .ZN(n428) );
  NAND2_X1 U253 ( .A1(\mem[13][7] ), .A2(n567), .ZN(n559) );
  OAI21_X1 U254 ( .B1(n411), .B2(n558), .A(n557), .ZN(n427) );
  NAND2_X1 U255 ( .A1(\mem[14][0] ), .A2(n558), .ZN(n557) );
  OAI21_X1 U256 ( .B1(n410), .B2(n558), .A(n556), .ZN(n426) );
  NAND2_X1 U257 ( .A1(\mem[14][1] ), .A2(n558), .ZN(n556) );
  OAI21_X1 U258 ( .B1(n409), .B2(n558), .A(n555), .ZN(n425) );
  NAND2_X1 U259 ( .A1(\mem[14][2] ), .A2(n558), .ZN(n555) );
  OAI21_X1 U260 ( .B1(n408), .B2(n558), .A(n554), .ZN(n424) );
  NAND2_X1 U261 ( .A1(\mem[14][3] ), .A2(n558), .ZN(n554) );
  OAI21_X1 U262 ( .B1(n407), .B2(n558), .A(n553), .ZN(n423) );
  NAND2_X1 U263 ( .A1(\mem[14][4] ), .A2(n558), .ZN(n553) );
  OAI21_X1 U264 ( .B1(n406), .B2(n558), .A(n552), .ZN(n422) );
  NAND2_X1 U265 ( .A1(\mem[14][5] ), .A2(n558), .ZN(n552) );
  OAI21_X1 U266 ( .B1(n405), .B2(n558), .A(n551), .ZN(n421) );
  NAND2_X1 U267 ( .A1(\mem[14][6] ), .A2(n558), .ZN(n551) );
  OAI21_X1 U268 ( .B1(n404), .B2(n558), .A(n550), .ZN(n420) );
  NAND2_X1 U269 ( .A1(\mem[14][7] ), .A2(n558), .ZN(n550) );
  OAI21_X1 U270 ( .B1(n411), .B2(n548), .A(n547), .ZN(n419) );
  NAND2_X1 U271 ( .A1(\mem[15][0] ), .A2(n548), .ZN(n547) );
  OAI21_X1 U272 ( .B1(n410), .B2(n548), .A(n546), .ZN(n418) );
  NAND2_X1 U273 ( .A1(\mem[15][1] ), .A2(n548), .ZN(n546) );
  OAI21_X1 U274 ( .B1(n409), .B2(n548), .A(n545), .ZN(n417) );
  NAND2_X1 U275 ( .A1(\mem[15][2] ), .A2(n548), .ZN(n545) );
  OAI21_X1 U276 ( .B1(n408), .B2(n548), .A(n544), .ZN(n416) );
  NAND2_X1 U277 ( .A1(\mem[15][3] ), .A2(n548), .ZN(n544) );
  OAI21_X1 U278 ( .B1(n407), .B2(n548), .A(n543), .ZN(n415) );
  NAND2_X1 U279 ( .A1(\mem[15][4] ), .A2(n548), .ZN(n543) );
  OAI21_X1 U280 ( .B1(n406), .B2(n548), .A(n542), .ZN(n414) );
  NAND2_X1 U281 ( .A1(\mem[15][5] ), .A2(n548), .ZN(n542) );
  OAI21_X1 U282 ( .B1(n405), .B2(n548), .A(n541), .ZN(n413) );
  NAND2_X1 U283 ( .A1(\mem[15][6] ), .A2(n548), .ZN(n541) );
  OAI21_X1 U284 ( .B1(n404), .B2(n548), .A(n540), .ZN(n412) );
  NAND2_X1 U285 ( .A1(\mem[15][7] ), .A2(n548), .ZN(n540) );
  AND2_X1 U286 ( .A1(N13), .A2(wr_en), .ZN(n549) );
  NOR2_X1 U287 ( .A1(N11), .A2(N12), .ZN(n684) );
  NOR2_X1 U288 ( .A1(n402), .A2(N12), .ZN(n663) );
  AND2_X1 U289 ( .A1(N12), .A2(n402), .ZN(n644) );
  AND2_X1 U290 ( .A1(N12), .A2(N11), .ZN(n625) );
  INV_X1 U291 ( .A(data_in[0]), .ZN(n411) );
  INV_X1 U292 ( .A(data_in[1]), .ZN(n410) );
  INV_X1 U293 ( .A(data_in[2]), .ZN(n409) );
  INV_X1 U294 ( .A(data_in[3]), .ZN(n408) );
  INV_X1 U295 ( .A(data_in[4]), .ZN(n407) );
  INV_X1 U296 ( .A(data_in[5]), .ZN(n406) );
  INV_X1 U297 ( .A(data_in[6]), .ZN(n405) );
  INV_X1 U298 ( .A(data_in[7]), .ZN(n404) );
  MUX2_X1 U299 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(N10), .Z(n3) );
  MUX2_X1 U300 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(N10), .Z(n4) );
  MUX2_X1 U301 ( .A(n4), .B(n3), .S(N11), .Z(n5) );
  MUX2_X1 U302 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(N10), .Z(n6) );
  MUX2_X1 U303 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n7) );
  MUX2_X1 U304 ( .A(n7), .B(n6), .S(N11), .Z(n8) );
  MUX2_X1 U305 ( .A(n8), .B(n5), .S(N12), .Z(n9) );
  MUX2_X1 U306 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n398), .Z(n10) );
  MUX2_X1 U307 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n398), .Z(n11) );
  MUX2_X1 U308 ( .A(n11), .B(n10), .S(N11), .Z(n294) );
  MUX2_X1 U309 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n398), .Z(n295) );
  MUX2_X1 U310 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n398), .Z(n296) );
  MUX2_X1 U311 ( .A(n296), .B(n295), .S(N11), .Z(n297) );
  MUX2_X1 U312 ( .A(n297), .B(n294), .S(N12), .Z(n298) );
  MUX2_X1 U313 ( .A(n298), .B(n9), .S(N13), .Z(N21) );
  MUX2_X1 U314 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n398), .Z(n299) );
  MUX2_X1 U315 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n398), .Z(n300) );
  MUX2_X1 U316 ( .A(n300), .B(n299), .S(N11), .Z(n301) );
  MUX2_X1 U317 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n398), .Z(n302) );
  MUX2_X1 U318 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n398), .Z(n303) );
  MUX2_X1 U319 ( .A(n303), .B(n302), .S(N11), .Z(n304) );
  MUX2_X1 U320 ( .A(n304), .B(n301), .S(N12), .Z(n305) );
  MUX2_X1 U321 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n398), .Z(n306) );
  MUX2_X1 U322 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n398), .Z(n307) );
  MUX2_X1 U323 ( .A(n307), .B(n306), .S(N11), .Z(n308) );
  MUX2_X1 U324 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n398), .Z(n309) );
  MUX2_X1 U325 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n398), .Z(n310) );
  MUX2_X1 U326 ( .A(n310), .B(n309), .S(N11), .Z(n311) );
  MUX2_X1 U327 ( .A(n311), .B(n308), .S(N12), .Z(n312) );
  MUX2_X1 U328 ( .A(n312), .B(n305), .S(N13), .Z(N20) );
  MUX2_X1 U329 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n399), .Z(n313) );
  MUX2_X1 U330 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n399), .Z(n314) );
  MUX2_X1 U331 ( .A(n314), .B(n313), .S(n397), .Z(n315) );
  MUX2_X1 U332 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n399), .Z(n316) );
  MUX2_X1 U333 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n399), .Z(n317) );
  MUX2_X1 U334 ( .A(n317), .B(n316), .S(n397), .Z(n318) );
  MUX2_X1 U335 ( .A(n318), .B(n315), .S(N12), .Z(n319) );
  MUX2_X1 U336 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n399), .Z(n320) );
  MUX2_X1 U337 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n399), .Z(n321) );
  MUX2_X1 U338 ( .A(n321), .B(n320), .S(n397), .Z(n322) );
  MUX2_X1 U339 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n399), .Z(n323) );
  MUX2_X1 U340 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n399), .Z(n324) );
  MUX2_X1 U341 ( .A(n324), .B(n323), .S(n397), .Z(n325) );
  MUX2_X1 U342 ( .A(n325), .B(n322), .S(N12), .Z(n326) );
  MUX2_X1 U343 ( .A(n326), .B(n319), .S(N13), .Z(N19) );
  MUX2_X1 U344 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n399), .Z(n327) );
  MUX2_X1 U345 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n399), .Z(n328) );
  MUX2_X1 U346 ( .A(n328), .B(n327), .S(n397), .Z(n329) );
  MUX2_X1 U347 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n399), .Z(n330) );
  MUX2_X1 U348 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n399), .Z(n331) );
  MUX2_X1 U349 ( .A(n331), .B(n330), .S(n397), .Z(n332) );
  MUX2_X1 U350 ( .A(n332), .B(n329), .S(N12), .Z(n333) );
  MUX2_X1 U351 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n400), .Z(n334) );
  MUX2_X1 U352 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n400), .Z(n335) );
  MUX2_X1 U353 ( .A(n335), .B(n334), .S(n397), .Z(n336) );
  MUX2_X1 U354 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n400), .Z(n337) );
  MUX2_X1 U355 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n400), .Z(n338) );
  MUX2_X1 U356 ( .A(n338), .B(n337), .S(n397), .Z(n339) );
  MUX2_X1 U357 ( .A(n339), .B(n336), .S(N12), .Z(n340) );
  MUX2_X1 U358 ( .A(n340), .B(n333), .S(N13), .Z(N18) );
  MUX2_X1 U359 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n400), .Z(n341) );
  MUX2_X1 U360 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n400), .Z(n342) );
  MUX2_X1 U361 ( .A(n342), .B(n341), .S(n397), .Z(n343) );
  MUX2_X1 U362 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n400), .Z(n344) );
  MUX2_X1 U363 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n400), .Z(n345) );
  MUX2_X1 U364 ( .A(n345), .B(n344), .S(n397), .Z(n346) );
  MUX2_X1 U365 ( .A(n346), .B(n343), .S(N12), .Z(n347) );
  MUX2_X1 U366 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n400), .Z(n348) );
  MUX2_X1 U367 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n400), .Z(n349) );
  MUX2_X1 U368 ( .A(n349), .B(n348), .S(n397), .Z(n350) );
  MUX2_X1 U369 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n400), .Z(n351) );
  MUX2_X1 U370 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n400), .Z(n352) );
  MUX2_X1 U371 ( .A(n352), .B(n351), .S(n397), .Z(n353) );
  MUX2_X1 U372 ( .A(n353), .B(n350), .S(N12), .Z(n354) );
  MUX2_X1 U373 ( .A(n354), .B(n347), .S(N13), .Z(N17) );
  MUX2_X1 U374 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n398), .Z(n355) );
  MUX2_X1 U375 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n400), .Z(n356) );
  MUX2_X1 U376 ( .A(n356), .B(n355), .S(N11), .Z(n357) );
  MUX2_X1 U377 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(N10), .Z(n358) );
  MUX2_X1 U378 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n400), .Z(n359) );
  MUX2_X1 U379 ( .A(n359), .B(n358), .S(N11), .Z(n360) );
  MUX2_X1 U380 ( .A(n360), .B(n357), .S(N12), .Z(n361) );
  MUX2_X1 U381 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n398), .Z(n362) );
  MUX2_X1 U382 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n398), .Z(n363) );
  MUX2_X1 U383 ( .A(n363), .B(n362), .S(N11), .Z(n364) );
  MUX2_X1 U384 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n398), .Z(n365) );
  MUX2_X1 U385 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n400), .Z(n366) );
  MUX2_X1 U386 ( .A(n366), .B(n365), .S(N11), .Z(n367) );
  MUX2_X1 U387 ( .A(n367), .B(n364), .S(N12), .Z(n368) );
  MUX2_X1 U388 ( .A(n368), .B(n361), .S(N13), .Z(N16) );
  MUX2_X1 U389 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n400), .Z(n369) );
  MUX2_X1 U390 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n399), .Z(n370) );
  MUX2_X1 U391 ( .A(n370), .B(n369), .S(N11), .Z(n371) );
  MUX2_X1 U392 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n399), .Z(n372) );
  MUX2_X1 U393 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n399), .Z(n373) );
  MUX2_X1 U394 ( .A(n373), .B(n372), .S(N11), .Z(n374) );
  MUX2_X1 U395 ( .A(n374), .B(n371), .S(N12), .Z(n375) );
  MUX2_X1 U396 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n376) );
  MUX2_X1 U397 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n377) );
  MUX2_X1 U398 ( .A(n377), .B(n376), .S(N11), .Z(n378) );
  MUX2_X1 U399 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n379) );
  MUX2_X1 U400 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n380) );
  MUX2_X1 U401 ( .A(n380), .B(n379), .S(n397), .Z(n381) );
  MUX2_X1 U402 ( .A(n381), .B(n378), .S(N12), .Z(n382) );
  MUX2_X1 U403 ( .A(n382), .B(n375), .S(N13), .Z(N15) );
  MUX2_X1 U404 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(N10), .Z(n383) );
  MUX2_X1 U405 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n384) );
  MUX2_X1 U406 ( .A(n384), .B(n383), .S(N11), .Z(n385) );
  MUX2_X1 U407 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(N10), .Z(n386) );
  MUX2_X1 U408 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n387) );
  MUX2_X1 U409 ( .A(n387), .B(n386), .S(N11), .Z(n388) );
  MUX2_X1 U410 ( .A(n388), .B(n385), .S(N12), .Z(n389) );
  MUX2_X1 U411 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n390) );
  MUX2_X1 U412 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n391) );
  MUX2_X1 U413 ( .A(n391), .B(n390), .S(N11), .Z(n392) );
  MUX2_X1 U414 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n393) );
  MUX2_X1 U415 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n399), .Z(n394) );
  MUX2_X1 U416 ( .A(n394), .B(n393), .S(n397), .Z(n395) );
  MUX2_X1 U417 ( .A(n395), .B(n392), .S(N12), .Z(n396) );
  MUX2_X1 U418 ( .A(n396), .B(n389), .S(N13), .Z(N14) );
  INV_X1 U419 ( .A(N10), .ZN(n401) );
  INV_X1 U420 ( .A(N11), .ZN(n402) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_8 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, N19, N20, N21, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N16), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n410), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n411), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n412), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n413), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n414), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n415), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n416), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n417), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n418), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n419), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n420), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n421), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n422), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n423), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n424), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n425), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n426), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n427), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n428), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n429), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n430), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n431), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n432), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n433), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n434), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n435), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n436), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n437), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n438), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n439), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n440), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n441), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n442), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n443), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n444), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n445), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n446), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n447), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n448), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n449), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n450), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n451), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n452), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n453), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n454), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n455), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n456), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n457), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n458), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n459), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n460), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n461), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n462), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n463), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n464), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n465), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n466), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n467), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n468), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n469), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n470), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n471), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n472), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n473), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n474), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n475), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n476), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n477), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n478), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n479), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n480), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n481), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n482), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n483), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n484), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n485), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n486), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n487), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n488), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n489), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n490), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n491), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n492), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n493), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n494), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n495), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n496), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n497), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n498), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n499), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n500), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n501), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n502), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n503), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n504), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n505), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n506), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n507), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n508), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n509), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n510), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n511), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n512), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n513), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n514), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n515), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n516), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n517), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n518), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n519), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n520), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n521), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n522), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n523), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n524), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n525), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n526), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n527), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n528), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n529), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n530), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n531), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n532), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n533), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n534), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n535), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n536), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n537), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[1]  ( .D(N20), .CK(clk), .Q(data_out[1]) );
  BUF_X1 U3 ( .A(N10), .Z(n396) );
  BUF_X1 U4 ( .A(N10), .Z(n397) );
  BUF_X1 U5 ( .A(N10), .Z(n398) );
  BUF_X1 U6 ( .A(N11), .Z(n395) );
  NAND2_X1 U7 ( .A1(n661), .A2(n681), .ZN(n670) );
  NAND2_X1 U8 ( .A1(n661), .A2(n671), .ZN(n660) );
  NAND2_X1 U9 ( .A1(n682), .A2(n681), .ZN(n691) );
  NAND2_X1 U10 ( .A1(n671), .A2(n682), .ZN(n680) );
  NAND2_X1 U11 ( .A1(n603), .A2(n682), .ZN(n612) );
  NAND2_X1 U12 ( .A1(n593), .A2(n682), .ZN(n602) );
  NAND2_X1 U13 ( .A1(n603), .A2(n661), .ZN(n592) );
  NAND2_X1 U14 ( .A1(n593), .A2(n661), .ZN(n583) );
  NAND2_X1 U15 ( .A1(n642), .A2(n681), .ZN(n651) );
  NAND2_X1 U16 ( .A1(n642), .A2(n671), .ZN(n641) );
  NAND2_X1 U17 ( .A1(n623), .A2(n681), .ZN(n632) );
  NAND2_X1 U18 ( .A1(n623), .A2(n671), .ZN(n621) );
  NAND2_X1 U19 ( .A1(n603), .A2(n642), .ZN(n574) );
  NAND2_X1 U20 ( .A1(n593), .A2(n642), .ZN(n565) );
  NAND2_X1 U21 ( .A1(n603), .A2(n623), .ZN(n556) );
  NAND2_X1 U22 ( .A1(n593), .A2(n623), .ZN(n546) );
  AND2_X1 U23 ( .A1(n547), .A2(N10), .ZN(n593) );
  AND2_X1 U24 ( .A1(n547), .A2(n399), .ZN(n603) );
  AND2_X1 U25 ( .A1(N10), .A2(n622), .ZN(n671) );
  AND2_X1 U26 ( .A1(n622), .A2(n399), .ZN(n681) );
  OAI21_X1 U27 ( .B1(n691), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U28 ( .A1(\mem[0][0] ), .A2(n691), .ZN(n690) );
  OAI21_X1 U29 ( .B1(n691), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U30 ( .A1(\mem[0][1] ), .A2(n691), .ZN(n689) );
  OAI21_X1 U31 ( .B1(n691), .B2(n407), .A(n688), .ZN(n535) );
  NAND2_X1 U32 ( .A1(\mem[0][2] ), .A2(n691), .ZN(n688) );
  OAI21_X1 U33 ( .B1(n691), .B2(n406), .A(n687), .ZN(n534) );
  NAND2_X1 U34 ( .A1(\mem[0][3] ), .A2(n691), .ZN(n687) );
  OAI21_X1 U35 ( .B1(n691), .B2(n405), .A(n686), .ZN(n533) );
  NAND2_X1 U36 ( .A1(\mem[0][4] ), .A2(n691), .ZN(n686) );
  OAI21_X1 U37 ( .B1(n691), .B2(n404), .A(n685), .ZN(n532) );
  NAND2_X1 U38 ( .A1(\mem[0][5] ), .A2(n691), .ZN(n685) );
  OAI21_X1 U39 ( .B1(n691), .B2(n403), .A(n684), .ZN(n531) );
  NAND2_X1 U40 ( .A1(\mem[0][6] ), .A2(n691), .ZN(n684) );
  OAI21_X1 U41 ( .B1(n691), .B2(n402), .A(n683), .ZN(n530) );
  NAND2_X1 U42 ( .A1(\mem[0][7] ), .A2(n691), .ZN(n683) );
  OAI21_X1 U43 ( .B1(n409), .B2(n670), .A(n669), .ZN(n521) );
  NAND2_X1 U44 ( .A1(\mem[2][0] ), .A2(n670), .ZN(n669) );
  OAI21_X1 U45 ( .B1(n408), .B2(n670), .A(n668), .ZN(n520) );
  NAND2_X1 U46 ( .A1(\mem[2][1] ), .A2(n670), .ZN(n668) );
  OAI21_X1 U47 ( .B1(n407), .B2(n670), .A(n667), .ZN(n519) );
  NAND2_X1 U48 ( .A1(\mem[2][2] ), .A2(n670), .ZN(n667) );
  OAI21_X1 U49 ( .B1(n406), .B2(n670), .A(n666), .ZN(n518) );
  NAND2_X1 U50 ( .A1(\mem[2][3] ), .A2(n670), .ZN(n666) );
  OAI21_X1 U51 ( .B1(n405), .B2(n670), .A(n665), .ZN(n517) );
  NAND2_X1 U52 ( .A1(\mem[2][4] ), .A2(n670), .ZN(n665) );
  OAI21_X1 U53 ( .B1(n404), .B2(n670), .A(n664), .ZN(n516) );
  NAND2_X1 U54 ( .A1(\mem[2][5] ), .A2(n670), .ZN(n664) );
  OAI21_X1 U55 ( .B1(n403), .B2(n670), .A(n663), .ZN(n515) );
  NAND2_X1 U56 ( .A1(\mem[2][6] ), .A2(n670), .ZN(n663) );
  OAI21_X1 U57 ( .B1(n402), .B2(n670), .A(n662), .ZN(n514) );
  NAND2_X1 U58 ( .A1(\mem[2][7] ), .A2(n670), .ZN(n662) );
  OAI21_X1 U59 ( .B1(n409), .B2(n660), .A(n659), .ZN(n513) );
  NAND2_X1 U60 ( .A1(\mem[3][0] ), .A2(n660), .ZN(n659) );
  OAI21_X1 U61 ( .B1(n408), .B2(n660), .A(n658), .ZN(n512) );
  NAND2_X1 U62 ( .A1(\mem[3][1] ), .A2(n660), .ZN(n658) );
  OAI21_X1 U63 ( .B1(n407), .B2(n660), .A(n657), .ZN(n511) );
  NAND2_X1 U64 ( .A1(\mem[3][2] ), .A2(n660), .ZN(n657) );
  OAI21_X1 U65 ( .B1(n406), .B2(n660), .A(n656), .ZN(n510) );
  NAND2_X1 U66 ( .A1(\mem[3][3] ), .A2(n660), .ZN(n656) );
  OAI21_X1 U67 ( .B1(n405), .B2(n660), .A(n655), .ZN(n509) );
  NAND2_X1 U68 ( .A1(\mem[3][4] ), .A2(n660), .ZN(n655) );
  OAI21_X1 U69 ( .B1(n404), .B2(n660), .A(n654), .ZN(n508) );
  NAND2_X1 U70 ( .A1(\mem[3][5] ), .A2(n660), .ZN(n654) );
  OAI21_X1 U71 ( .B1(n403), .B2(n660), .A(n653), .ZN(n507) );
  NAND2_X1 U72 ( .A1(\mem[3][6] ), .A2(n660), .ZN(n653) );
  OAI21_X1 U73 ( .B1(n402), .B2(n660), .A(n652), .ZN(n506) );
  NAND2_X1 U74 ( .A1(\mem[3][7] ), .A2(n660), .ZN(n652) );
  NOR2_X1 U75 ( .A1(n401), .A2(N13), .ZN(n622) );
  INV_X1 U76 ( .A(wr_en), .ZN(n401) );
  OAI21_X1 U77 ( .B1(n409), .B2(n680), .A(n679), .ZN(n529) );
  NAND2_X1 U78 ( .A1(\mem[1][0] ), .A2(n680), .ZN(n679) );
  OAI21_X1 U79 ( .B1(n408), .B2(n680), .A(n678), .ZN(n528) );
  NAND2_X1 U80 ( .A1(\mem[1][1] ), .A2(n680), .ZN(n678) );
  OAI21_X1 U81 ( .B1(n407), .B2(n680), .A(n677), .ZN(n527) );
  NAND2_X1 U82 ( .A1(\mem[1][2] ), .A2(n680), .ZN(n677) );
  OAI21_X1 U83 ( .B1(n406), .B2(n680), .A(n676), .ZN(n526) );
  NAND2_X1 U84 ( .A1(\mem[1][3] ), .A2(n680), .ZN(n676) );
  OAI21_X1 U85 ( .B1(n405), .B2(n680), .A(n675), .ZN(n525) );
  NAND2_X1 U86 ( .A1(\mem[1][4] ), .A2(n680), .ZN(n675) );
  OAI21_X1 U87 ( .B1(n404), .B2(n680), .A(n674), .ZN(n524) );
  NAND2_X1 U88 ( .A1(\mem[1][5] ), .A2(n680), .ZN(n674) );
  OAI21_X1 U89 ( .B1(n403), .B2(n680), .A(n673), .ZN(n523) );
  NAND2_X1 U90 ( .A1(\mem[1][6] ), .A2(n680), .ZN(n673) );
  OAI21_X1 U91 ( .B1(n402), .B2(n680), .A(n672), .ZN(n522) );
  NAND2_X1 U92 ( .A1(\mem[1][7] ), .A2(n680), .ZN(n672) );
  OAI21_X1 U93 ( .B1(n409), .B2(n651), .A(n650), .ZN(n505) );
  NAND2_X1 U94 ( .A1(\mem[4][0] ), .A2(n651), .ZN(n650) );
  OAI21_X1 U95 ( .B1(n408), .B2(n651), .A(n649), .ZN(n504) );
  NAND2_X1 U96 ( .A1(\mem[4][1] ), .A2(n651), .ZN(n649) );
  OAI21_X1 U97 ( .B1(n407), .B2(n651), .A(n648), .ZN(n503) );
  NAND2_X1 U98 ( .A1(\mem[4][2] ), .A2(n651), .ZN(n648) );
  OAI21_X1 U99 ( .B1(n406), .B2(n651), .A(n647), .ZN(n502) );
  NAND2_X1 U100 ( .A1(\mem[4][3] ), .A2(n651), .ZN(n647) );
  OAI21_X1 U101 ( .B1(n405), .B2(n651), .A(n646), .ZN(n501) );
  NAND2_X1 U102 ( .A1(\mem[4][4] ), .A2(n651), .ZN(n646) );
  OAI21_X1 U103 ( .B1(n404), .B2(n651), .A(n645), .ZN(n500) );
  NAND2_X1 U104 ( .A1(\mem[4][5] ), .A2(n651), .ZN(n645) );
  OAI21_X1 U105 ( .B1(n403), .B2(n651), .A(n644), .ZN(n499) );
  NAND2_X1 U106 ( .A1(\mem[4][6] ), .A2(n651), .ZN(n644) );
  OAI21_X1 U107 ( .B1(n402), .B2(n651), .A(n643), .ZN(n498) );
  NAND2_X1 U108 ( .A1(\mem[4][7] ), .A2(n651), .ZN(n643) );
  OAI21_X1 U109 ( .B1(n409), .B2(n641), .A(n640), .ZN(n497) );
  NAND2_X1 U110 ( .A1(\mem[5][0] ), .A2(n641), .ZN(n640) );
  OAI21_X1 U111 ( .B1(n408), .B2(n641), .A(n639), .ZN(n496) );
  NAND2_X1 U112 ( .A1(\mem[5][1] ), .A2(n641), .ZN(n639) );
  OAI21_X1 U113 ( .B1(n407), .B2(n641), .A(n638), .ZN(n495) );
  NAND2_X1 U114 ( .A1(\mem[5][2] ), .A2(n641), .ZN(n638) );
  OAI21_X1 U115 ( .B1(n406), .B2(n641), .A(n637), .ZN(n494) );
  NAND2_X1 U116 ( .A1(\mem[5][3] ), .A2(n641), .ZN(n637) );
  OAI21_X1 U117 ( .B1(n405), .B2(n641), .A(n636), .ZN(n493) );
  NAND2_X1 U118 ( .A1(\mem[5][4] ), .A2(n641), .ZN(n636) );
  OAI21_X1 U119 ( .B1(n404), .B2(n641), .A(n635), .ZN(n492) );
  NAND2_X1 U120 ( .A1(\mem[5][5] ), .A2(n641), .ZN(n635) );
  OAI21_X1 U121 ( .B1(n403), .B2(n641), .A(n634), .ZN(n491) );
  NAND2_X1 U122 ( .A1(\mem[5][6] ), .A2(n641), .ZN(n634) );
  OAI21_X1 U123 ( .B1(n402), .B2(n641), .A(n633), .ZN(n490) );
  NAND2_X1 U124 ( .A1(\mem[5][7] ), .A2(n641), .ZN(n633) );
  OAI21_X1 U125 ( .B1(n409), .B2(n632), .A(n631), .ZN(n489) );
  NAND2_X1 U126 ( .A1(\mem[6][0] ), .A2(n632), .ZN(n631) );
  OAI21_X1 U127 ( .B1(n408), .B2(n632), .A(n630), .ZN(n488) );
  NAND2_X1 U128 ( .A1(\mem[6][1] ), .A2(n632), .ZN(n630) );
  OAI21_X1 U129 ( .B1(n407), .B2(n632), .A(n629), .ZN(n487) );
  NAND2_X1 U130 ( .A1(\mem[6][2] ), .A2(n632), .ZN(n629) );
  OAI21_X1 U131 ( .B1(n406), .B2(n632), .A(n628), .ZN(n486) );
  NAND2_X1 U132 ( .A1(\mem[6][3] ), .A2(n632), .ZN(n628) );
  OAI21_X1 U133 ( .B1(n405), .B2(n632), .A(n627), .ZN(n485) );
  NAND2_X1 U134 ( .A1(\mem[6][4] ), .A2(n632), .ZN(n627) );
  OAI21_X1 U135 ( .B1(n404), .B2(n632), .A(n626), .ZN(n484) );
  NAND2_X1 U136 ( .A1(\mem[6][5] ), .A2(n632), .ZN(n626) );
  OAI21_X1 U137 ( .B1(n403), .B2(n632), .A(n625), .ZN(n483) );
  NAND2_X1 U138 ( .A1(\mem[6][6] ), .A2(n632), .ZN(n625) );
  OAI21_X1 U139 ( .B1(n402), .B2(n632), .A(n624), .ZN(n482) );
  NAND2_X1 U140 ( .A1(\mem[6][7] ), .A2(n632), .ZN(n624) );
  OAI21_X1 U141 ( .B1(n409), .B2(n621), .A(n620), .ZN(n481) );
  NAND2_X1 U142 ( .A1(\mem[7][0] ), .A2(n621), .ZN(n620) );
  OAI21_X1 U143 ( .B1(n408), .B2(n621), .A(n619), .ZN(n480) );
  NAND2_X1 U144 ( .A1(\mem[7][1] ), .A2(n621), .ZN(n619) );
  OAI21_X1 U145 ( .B1(n407), .B2(n621), .A(n618), .ZN(n479) );
  NAND2_X1 U146 ( .A1(\mem[7][2] ), .A2(n621), .ZN(n618) );
  OAI21_X1 U147 ( .B1(n406), .B2(n621), .A(n617), .ZN(n478) );
  NAND2_X1 U148 ( .A1(\mem[7][3] ), .A2(n621), .ZN(n617) );
  OAI21_X1 U149 ( .B1(n405), .B2(n621), .A(n616), .ZN(n477) );
  NAND2_X1 U150 ( .A1(\mem[7][4] ), .A2(n621), .ZN(n616) );
  OAI21_X1 U151 ( .B1(n404), .B2(n621), .A(n615), .ZN(n476) );
  NAND2_X1 U152 ( .A1(\mem[7][5] ), .A2(n621), .ZN(n615) );
  OAI21_X1 U153 ( .B1(n403), .B2(n621), .A(n614), .ZN(n475) );
  NAND2_X1 U154 ( .A1(\mem[7][6] ), .A2(n621), .ZN(n614) );
  OAI21_X1 U155 ( .B1(n402), .B2(n621), .A(n613), .ZN(n474) );
  NAND2_X1 U156 ( .A1(\mem[7][7] ), .A2(n621), .ZN(n613) );
  OAI21_X1 U157 ( .B1(n409), .B2(n612), .A(n611), .ZN(n473) );
  NAND2_X1 U158 ( .A1(\mem[8][0] ), .A2(n612), .ZN(n611) );
  OAI21_X1 U159 ( .B1(n408), .B2(n612), .A(n610), .ZN(n472) );
  NAND2_X1 U160 ( .A1(\mem[8][1] ), .A2(n612), .ZN(n610) );
  OAI21_X1 U161 ( .B1(n407), .B2(n612), .A(n609), .ZN(n471) );
  NAND2_X1 U162 ( .A1(\mem[8][2] ), .A2(n612), .ZN(n609) );
  OAI21_X1 U163 ( .B1(n406), .B2(n612), .A(n608), .ZN(n470) );
  NAND2_X1 U164 ( .A1(\mem[8][3] ), .A2(n612), .ZN(n608) );
  OAI21_X1 U165 ( .B1(n405), .B2(n612), .A(n607), .ZN(n469) );
  NAND2_X1 U166 ( .A1(\mem[8][4] ), .A2(n612), .ZN(n607) );
  OAI21_X1 U167 ( .B1(n404), .B2(n612), .A(n606), .ZN(n468) );
  NAND2_X1 U168 ( .A1(\mem[8][5] ), .A2(n612), .ZN(n606) );
  OAI21_X1 U169 ( .B1(n403), .B2(n612), .A(n605), .ZN(n467) );
  NAND2_X1 U170 ( .A1(\mem[8][6] ), .A2(n612), .ZN(n605) );
  OAI21_X1 U171 ( .B1(n402), .B2(n612), .A(n604), .ZN(n466) );
  NAND2_X1 U172 ( .A1(\mem[8][7] ), .A2(n612), .ZN(n604) );
  OAI21_X1 U173 ( .B1(n409), .B2(n602), .A(n601), .ZN(n465) );
  NAND2_X1 U174 ( .A1(\mem[9][0] ), .A2(n602), .ZN(n601) );
  OAI21_X1 U175 ( .B1(n408), .B2(n602), .A(n600), .ZN(n464) );
  NAND2_X1 U176 ( .A1(\mem[9][1] ), .A2(n602), .ZN(n600) );
  OAI21_X1 U177 ( .B1(n407), .B2(n602), .A(n599), .ZN(n463) );
  NAND2_X1 U178 ( .A1(\mem[9][2] ), .A2(n602), .ZN(n599) );
  OAI21_X1 U179 ( .B1(n406), .B2(n602), .A(n598), .ZN(n462) );
  NAND2_X1 U180 ( .A1(\mem[9][3] ), .A2(n602), .ZN(n598) );
  OAI21_X1 U181 ( .B1(n405), .B2(n602), .A(n597), .ZN(n461) );
  NAND2_X1 U182 ( .A1(\mem[9][4] ), .A2(n602), .ZN(n597) );
  OAI21_X1 U183 ( .B1(n404), .B2(n602), .A(n596), .ZN(n460) );
  NAND2_X1 U184 ( .A1(\mem[9][5] ), .A2(n602), .ZN(n596) );
  OAI21_X1 U185 ( .B1(n403), .B2(n602), .A(n595), .ZN(n459) );
  NAND2_X1 U186 ( .A1(\mem[9][6] ), .A2(n602), .ZN(n595) );
  OAI21_X1 U187 ( .B1(n402), .B2(n602), .A(n594), .ZN(n458) );
  NAND2_X1 U188 ( .A1(\mem[9][7] ), .A2(n602), .ZN(n594) );
  OAI21_X1 U189 ( .B1(n409), .B2(n592), .A(n591), .ZN(n457) );
  NAND2_X1 U190 ( .A1(\mem[10][0] ), .A2(n592), .ZN(n591) );
  OAI21_X1 U191 ( .B1(n408), .B2(n592), .A(n590), .ZN(n456) );
  NAND2_X1 U192 ( .A1(\mem[10][1] ), .A2(n592), .ZN(n590) );
  OAI21_X1 U193 ( .B1(n407), .B2(n592), .A(n589), .ZN(n455) );
  NAND2_X1 U194 ( .A1(\mem[10][2] ), .A2(n592), .ZN(n589) );
  OAI21_X1 U195 ( .B1(n406), .B2(n592), .A(n588), .ZN(n454) );
  NAND2_X1 U196 ( .A1(\mem[10][3] ), .A2(n592), .ZN(n588) );
  OAI21_X1 U197 ( .B1(n405), .B2(n592), .A(n587), .ZN(n453) );
  NAND2_X1 U198 ( .A1(\mem[10][4] ), .A2(n592), .ZN(n587) );
  OAI21_X1 U199 ( .B1(n404), .B2(n592), .A(n586), .ZN(n452) );
  NAND2_X1 U200 ( .A1(\mem[10][5] ), .A2(n592), .ZN(n586) );
  OAI21_X1 U201 ( .B1(n403), .B2(n592), .A(n585), .ZN(n451) );
  NAND2_X1 U202 ( .A1(\mem[10][6] ), .A2(n592), .ZN(n585) );
  OAI21_X1 U203 ( .B1(n402), .B2(n592), .A(n584), .ZN(n450) );
  NAND2_X1 U204 ( .A1(\mem[10][7] ), .A2(n592), .ZN(n584) );
  OAI21_X1 U205 ( .B1(n409), .B2(n583), .A(n582), .ZN(n449) );
  NAND2_X1 U206 ( .A1(\mem[11][0] ), .A2(n583), .ZN(n582) );
  OAI21_X1 U207 ( .B1(n408), .B2(n583), .A(n581), .ZN(n448) );
  NAND2_X1 U208 ( .A1(\mem[11][1] ), .A2(n583), .ZN(n581) );
  OAI21_X1 U209 ( .B1(n407), .B2(n583), .A(n580), .ZN(n447) );
  NAND2_X1 U210 ( .A1(\mem[11][2] ), .A2(n583), .ZN(n580) );
  OAI21_X1 U211 ( .B1(n406), .B2(n583), .A(n579), .ZN(n446) );
  NAND2_X1 U212 ( .A1(\mem[11][3] ), .A2(n583), .ZN(n579) );
  OAI21_X1 U213 ( .B1(n405), .B2(n583), .A(n578), .ZN(n445) );
  NAND2_X1 U214 ( .A1(\mem[11][4] ), .A2(n583), .ZN(n578) );
  OAI21_X1 U215 ( .B1(n404), .B2(n583), .A(n577), .ZN(n444) );
  NAND2_X1 U216 ( .A1(\mem[11][5] ), .A2(n583), .ZN(n577) );
  OAI21_X1 U217 ( .B1(n403), .B2(n583), .A(n576), .ZN(n443) );
  NAND2_X1 U218 ( .A1(\mem[11][6] ), .A2(n583), .ZN(n576) );
  OAI21_X1 U219 ( .B1(n402), .B2(n583), .A(n575), .ZN(n442) );
  NAND2_X1 U220 ( .A1(\mem[11][7] ), .A2(n583), .ZN(n575) );
  OAI21_X1 U221 ( .B1(n409), .B2(n574), .A(n573), .ZN(n441) );
  NAND2_X1 U222 ( .A1(\mem[12][0] ), .A2(n574), .ZN(n573) );
  OAI21_X1 U223 ( .B1(n408), .B2(n574), .A(n572), .ZN(n440) );
  NAND2_X1 U224 ( .A1(\mem[12][1] ), .A2(n574), .ZN(n572) );
  OAI21_X1 U225 ( .B1(n407), .B2(n574), .A(n571), .ZN(n439) );
  NAND2_X1 U226 ( .A1(\mem[12][2] ), .A2(n574), .ZN(n571) );
  OAI21_X1 U227 ( .B1(n406), .B2(n574), .A(n570), .ZN(n438) );
  NAND2_X1 U228 ( .A1(\mem[12][3] ), .A2(n574), .ZN(n570) );
  OAI21_X1 U229 ( .B1(n405), .B2(n574), .A(n569), .ZN(n437) );
  NAND2_X1 U230 ( .A1(\mem[12][4] ), .A2(n574), .ZN(n569) );
  OAI21_X1 U231 ( .B1(n404), .B2(n574), .A(n568), .ZN(n436) );
  NAND2_X1 U232 ( .A1(\mem[12][5] ), .A2(n574), .ZN(n568) );
  OAI21_X1 U233 ( .B1(n403), .B2(n574), .A(n567), .ZN(n435) );
  NAND2_X1 U234 ( .A1(\mem[12][6] ), .A2(n574), .ZN(n567) );
  OAI21_X1 U235 ( .B1(n402), .B2(n574), .A(n566), .ZN(n434) );
  NAND2_X1 U236 ( .A1(\mem[12][7] ), .A2(n574), .ZN(n566) );
  OAI21_X1 U237 ( .B1(n409), .B2(n565), .A(n564), .ZN(n433) );
  NAND2_X1 U238 ( .A1(\mem[13][0] ), .A2(n565), .ZN(n564) );
  OAI21_X1 U239 ( .B1(n408), .B2(n565), .A(n563), .ZN(n432) );
  NAND2_X1 U240 ( .A1(\mem[13][1] ), .A2(n565), .ZN(n563) );
  OAI21_X1 U241 ( .B1(n407), .B2(n565), .A(n562), .ZN(n431) );
  NAND2_X1 U242 ( .A1(\mem[13][2] ), .A2(n565), .ZN(n562) );
  OAI21_X1 U243 ( .B1(n406), .B2(n565), .A(n561), .ZN(n430) );
  NAND2_X1 U244 ( .A1(\mem[13][3] ), .A2(n565), .ZN(n561) );
  OAI21_X1 U245 ( .B1(n405), .B2(n565), .A(n560), .ZN(n429) );
  NAND2_X1 U246 ( .A1(\mem[13][4] ), .A2(n565), .ZN(n560) );
  OAI21_X1 U247 ( .B1(n404), .B2(n565), .A(n559), .ZN(n428) );
  NAND2_X1 U248 ( .A1(\mem[13][5] ), .A2(n565), .ZN(n559) );
  OAI21_X1 U249 ( .B1(n403), .B2(n565), .A(n558), .ZN(n427) );
  NAND2_X1 U250 ( .A1(\mem[13][6] ), .A2(n565), .ZN(n558) );
  OAI21_X1 U251 ( .B1(n402), .B2(n565), .A(n557), .ZN(n426) );
  NAND2_X1 U252 ( .A1(\mem[13][7] ), .A2(n565), .ZN(n557) );
  OAI21_X1 U253 ( .B1(n409), .B2(n556), .A(n555), .ZN(n425) );
  NAND2_X1 U254 ( .A1(\mem[14][0] ), .A2(n556), .ZN(n555) );
  OAI21_X1 U255 ( .B1(n408), .B2(n556), .A(n554), .ZN(n424) );
  NAND2_X1 U256 ( .A1(\mem[14][1] ), .A2(n556), .ZN(n554) );
  OAI21_X1 U257 ( .B1(n407), .B2(n556), .A(n553), .ZN(n423) );
  NAND2_X1 U258 ( .A1(\mem[14][2] ), .A2(n556), .ZN(n553) );
  OAI21_X1 U259 ( .B1(n406), .B2(n556), .A(n552), .ZN(n422) );
  NAND2_X1 U260 ( .A1(\mem[14][3] ), .A2(n556), .ZN(n552) );
  OAI21_X1 U261 ( .B1(n405), .B2(n556), .A(n551), .ZN(n421) );
  NAND2_X1 U262 ( .A1(\mem[14][4] ), .A2(n556), .ZN(n551) );
  OAI21_X1 U263 ( .B1(n404), .B2(n556), .A(n550), .ZN(n420) );
  NAND2_X1 U264 ( .A1(\mem[14][5] ), .A2(n556), .ZN(n550) );
  OAI21_X1 U265 ( .B1(n403), .B2(n556), .A(n549), .ZN(n419) );
  NAND2_X1 U266 ( .A1(\mem[14][6] ), .A2(n556), .ZN(n549) );
  OAI21_X1 U267 ( .B1(n402), .B2(n556), .A(n548), .ZN(n418) );
  NAND2_X1 U268 ( .A1(\mem[14][7] ), .A2(n556), .ZN(n548) );
  OAI21_X1 U269 ( .B1(n409), .B2(n546), .A(n545), .ZN(n417) );
  NAND2_X1 U270 ( .A1(\mem[15][0] ), .A2(n546), .ZN(n545) );
  OAI21_X1 U271 ( .B1(n408), .B2(n546), .A(n544), .ZN(n416) );
  NAND2_X1 U272 ( .A1(\mem[15][1] ), .A2(n546), .ZN(n544) );
  OAI21_X1 U273 ( .B1(n407), .B2(n546), .A(n543), .ZN(n415) );
  NAND2_X1 U274 ( .A1(\mem[15][2] ), .A2(n546), .ZN(n543) );
  OAI21_X1 U275 ( .B1(n406), .B2(n546), .A(n542), .ZN(n414) );
  NAND2_X1 U276 ( .A1(\mem[15][3] ), .A2(n546), .ZN(n542) );
  OAI21_X1 U277 ( .B1(n405), .B2(n546), .A(n541), .ZN(n413) );
  NAND2_X1 U278 ( .A1(\mem[15][4] ), .A2(n546), .ZN(n541) );
  OAI21_X1 U279 ( .B1(n404), .B2(n546), .A(n540), .ZN(n412) );
  NAND2_X1 U280 ( .A1(\mem[15][5] ), .A2(n546), .ZN(n540) );
  OAI21_X1 U281 ( .B1(n403), .B2(n546), .A(n539), .ZN(n411) );
  NAND2_X1 U282 ( .A1(\mem[15][6] ), .A2(n546), .ZN(n539) );
  OAI21_X1 U283 ( .B1(n402), .B2(n546), .A(n538), .ZN(n410) );
  NAND2_X1 U284 ( .A1(\mem[15][7] ), .A2(n546), .ZN(n538) );
  AND2_X1 U285 ( .A1(N13), .A2(wr_en), .ZN(n547) );
  NOR2_X1 U286 ( .A1(N11), .A2(N12), .ZN(n682) );
  NOR2_X1 U287 ( .A1(n400), .A2(N12), .ZN(n661) );
  AND2_X1 U288 ( .A1(N12), .A2(n400), .ZN(n642) );
  AND2_X1 U289 ( .A1(N12), .A2(N11), .ZN(n623) );
  INV_X1 U290 ( .A(data_in[0]), .ZN(n409) );
  INV_X1 U291 ( .A(data_in[1]), .ZN(n408) );
  INV_X1 U292 ( .A(data_in[2]), .ZN(n407) );
  INV_X1 U293 ( .A(data_in[3]), .ZN(n406) );
  INV_X1 U294 ( .A(data_in[4]), .ZN(n405) );
  INV_X1 U295 ( .A(data_in[5]), .ZN(n404) );
  INV_X1 U296 ( .A(data_in[6]), .ZN(n403) );
  INV_X1 U297 ( .A(data_in[7]), .ZN(n402) );
  MUX2_X1 U298 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n397), .Z(n1) );
  MUX2_X1 U299 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n397), .Z(n2) );
  MUX2_X1 U300 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U301 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n398), .Z(n4) );
  MUX2_X1 U302 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n5) );
  MUX2_X1 U303 ( .A(n5), .B(n4), .S(N11), .Z(n6) );
  MUX2_X1 U304 ( .A(n6), .B(n3), .S(N12), .Z(n7) );
  MUX2_X1 U305 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n396), .Z(n8) );
  MUX2_X1 U306 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n396), .Z(n9) );
  MUX2_X1 U307 ( .A(n9), .B(n8), .S(N11), .Z(n10) );
  MUX2_X1 U308 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n396), .Z(n11) );
  MUX2_X1 U309 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n396), .Z(n294) );
  MUX2_X1 U310 ( .A(n294), .B(n11), .S(N11), .Z(n295) );
  MUX2_X1 U311 ( .A(n295), .B(n10), .S(N12), .Z(n296) );
  MUX2_X1 U312 ( .A(n296), .B(n7), .S(N13), .Z(N21) );
  MUX2_X1 U313 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n396), .Z(n297) );
  MUX2_X1 U314 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n396), .Z(n298) );
  MUX2_X1 U315 ( .A(n298), .B(n297), .S(N11), .Z(n299) );
  MUX2_X1 U316 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n396), .Z(n300) );
  MUX2_X1 U317 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n396), .Z(n301) );
  MUX2_X1 U318 ( .A(n301), .B(n300), .S(N11), .Z(n302) );
  MUX2_X1 U319 ( .A(n302), .B(n299), .S(N12), .Z(n303) );
  MUX2_X1 U320 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n396), .Z(n304) );
  MUX2_X1 U321 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n396), .Z(n305) );
  MUX2_X1 U322 ( .A(n305), .B(n304), .S(N11), .Z(n306) );
  MUX2_X1 U323 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n396), .Z(n307) );
  MUX2_X1 U324 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n396), .Z(n308) );
  MUX2_X1 U325 ( .A(n308), .B(n307), .S(N11), .Z(n309) );
  MUX2_X1 U326 ( .A(n309), .B(n306), .S(N12), .Z(n310) );
  MUX2_X1 U327 ( .A(n310), .B(n303), .S(N13), .Z(N20) );
  MUX2_X1 U328 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n397), .Z(n311) );
  MUX2_X1 U329 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n397), .Z(n312) );
  MUX2_X1 U330 ( .A(n312), .B(n311), .S(n395), .Z(n313) );
  MUX2_X1 U331 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n397), .Z(n314) );
  MUX2_X1 U332 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n397), .Z(n315) );
  MUX2_X1 U333 ( .A(n315), .B(n314), .S(n395), .Z(n316) );
  MUX2_X1 U334 ( .A(n316), .B(n313), .S(N12), .Z(n317) );
  MUX2_X1 U335 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n397), .Z(n318) );
  MUX2_X1 U336 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n397), .Z(n319) );
  MUX2_X1 U337 ( .A(n319), .B(n318), .S(n395), .Z(n320) );
  MUX2_X1 U338 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n397), .Z(n321) );
  MUX2_X1 U339 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n397), .Z(n322) );
  MUX2_X1 U340 ( .A(n322), .B(n321), .S(n395), .Z(n323) );
  MUX2_X1 U341 ( .A(n323), .B(n320), .S(N12), .Z(n324) );
  MUX2_X1 U342 ( .A(n324), .B(n317), .S(N13), .Z(N19) );
  MUX2_X1 U343 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n397), .Z(n325) );
  MUX2_X1 U344 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n397), .Z(n326) );
  MUX2_X1 U345 ( .A(n326), .B(n325), .S(n395), .Z(n327) );
  MUX2_X1 U346 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n397), .Z(n328) );
  MUX2_X1 U347 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n397), .Z(n329) );
  MUX2_X1 U348 ( .A(n329), .B(n328), .S(n395), .Z(n330) );
  MUX2_X1 U349 ( .A(n330), .B(n327), .S(N12), .Z(n331) );
  MUX2_X1 U350 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n398), .Z(n332) );
  MUX2_X1 U351 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n398), .Z(n333) );
  MUX2_X1 U352 ( .A(n333), .B(n332), .S(n395), .Z(n334) );
  MUX2_X1 U353 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n398), .Z(n335) );
  MUX2_X1 U354 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n398), .Z(n336) );
  MUX2_X1 U355 ( .A(n336), .B(n335), .S(n395), .Z(n337) );
  MUX2_X1 U356 ( .A(n337), .B(n334), .S(N12), .Z(n338) );
  MUX2_X1 U357 ( .A(n338), .B(n331), .S(N13), .Z(N18) );
  MUX2_X1 U358 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n398), .Z(n339) );
  MUX2_X1 U359 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n398), .Z(n340) );
  MUX2_X1 U360 ( .A(n340), .B(n339), .S(n395), .Z(n341) );
  MUX2_X1 U361 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n398), .Z(n342) );
  MUX2_X1 U362 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n398), .Z(n343) );
  MUX2_X1 U363 ( .A(n343), .B(n342), .S(n395), .Z(n344) );
  MUX2_X1 U364 ( .A(n344), .B(n341), .S(N12), .Z(n345) );
  MUX2_X1 U365 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n398), .Z(n346) );
  MUX2_X1 U366 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n398), .Z(n347) );
  MUX2_X1 U367 ( .A(n347), .B(n346), .S(n395), .Z(n348) );
  MUX2_X1 U368 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n398), .Z(n349) );
  MUX2_X1 U369 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n398), .Z(n350) );
  MUX2_X1 U370 ( .A(n350), .B(n349), .S(n395), .Z(n351) );
  MUX2_X1 U371 ( .A(n351), .B(n348), .S(N12), .Z(n352) );
  MUX2_X1 U372 ( .A(n352), .B(n345), .S(N13), .Z(N17) );
  MUX2_X1 U373 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n397), .Z(n353) );
  MUX2_X1 U374 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(N10), .Z(n354) );
  MUX2_X1 U375 ( .A(n354), .B(n353), .S(N11), .Z(n355) );
  MUX2_X1 U376 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(N10), .Z(n356) );
  MUX2_X1 U377 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n396), .Z(n357) );
  MUX2_X1 U378 ( .A(n357), .B(n356), .S(N11), .Z(n358) );
  MUX2_X1 U379 ( .A(n358), .B(n355), .S(N12), .Z(n359) );
  MUX2_X1 U380 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(N10), .Z(n360) );
  MUX2_X1 U381 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n398), .Z(n361) );
  MUX2_X1 U382 ( .A(n361), .B(n360), .S(N11), .Z(n362) );
  MUX2_X1 U383 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n398), .Z(n363) );
  MUX2_X1 U384 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n396), .Z(n364) );
  MUX2_X1 U385 ( .A(n364), .B(n363), .S(N11), .Z(n365) );
  MUX2_X1 U386 ( .A(n365), .B(n362), .S(N12), .Z(n366) );
  MUX2_X1 U387 ( .A(n366), .B(n359), .S(N13), .Z(N16) );
  MUX2_X1 U388 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n398), .Z(n367) );
  MUX2_X1 U389 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n396), .Z(n368) );
  MUX2_X1 U390 ( .A(n368), .B(n367), .S(N11), .Z(n369) );
  MUX2_X1 U391 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(N10), .Z(n370) );
  MUX2_X1 U392 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n397), .Z(n371) );
  MUX2_X1 U393 ( .A(n371), .B(n370), .S(N11), .Z(n372) );
  MUX2_X1 U394 ( .A(n372), .B(n369), .S(N12), .Z(n373) );
  MUX2_X1 U395 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n374) );
  MUX2_X1 U396 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n375) );
  MUX2_X1 U397 ( .A(n375), .B(n374), .S(N11), .Z(n376) );
  MUX2_X1 U398 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n377) );
  MUX2_X1 U399 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n378) );
  MUX2_X1 U400 ( .A(n378), .B(n377), .S(n395), .Z(n379) );
  MUX2_X1 U401 ( .A(n379), .B(n376), .S(N12), .Z(n380) );
  MUX2_X1 U402 ( .A(n380), .B(n373), .S(N13), .Z(N15) );
  MUX2_X1 U403 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n396), .Z(n381) );
  MUX2_X1 U404 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n382) );
  MUX2_X1 U405 ( .A(n382), .B(n381), .S(N11), .Z(n383) );
  MUX2_X1 U406 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(N10), .Z(n384) );
  MUX2_X1 U407 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n385) );
  MUX2_X1 U408 ( .A(n385), .B(n384), .S(N11), .Z(n386) );
  MUX2_X1 U409 ( .A(n386), .B(n383), .S(N12), .Z(n387) );
  MUX2_X1 U410 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n388) );
  MUX2_X1 U411 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n389) );
  MUX2_X1 U412 ( .A(n389), .B(n388), .S(N11), .Z(n390) );
  MUX2_X1 U413 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n391) );
  MUX2_X1 U414 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n392) );
  MUX2_X1 U415 ( .A(n392), .B(n391), .S(n395), .Z(n393) );
  MUX2_X1 U416 ( .A(n393), .B(n390), .S(N12), .Z(n394) );
  MUX2_X1 U417 ( .A(n394), .B(n387), .S(N13), .Z(N14) );
  INV_X1 U418 ( .A(N10), .ZN(n399) );
  INV_X1 U419 ( .A(N11), .ZN(n400) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_7 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, N19, N20, N21, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N20), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n411), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n412), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n413), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n414), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n415), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n416), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n417), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n418), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n419), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n420), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n421), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n422), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n423), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n424), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n425), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n426), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n427), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n428), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n429), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n430), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n431), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n432), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n433), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n434), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n435), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n436), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n437), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n438), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n439), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n440), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n441), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n442), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n443), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n444), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n445), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n446), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n447), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n448), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n449), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n450), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n451), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n452), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n453), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n454), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n455), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n456), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n457), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n458), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n459), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n460), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n461), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n462), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n463), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n464), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n465), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n466), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n467), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n468), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n469), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n470), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n471), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n472), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n473), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n474), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n475), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n476), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n477), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n478), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n479), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n480), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n481), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n482), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n483), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n484), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n485), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n486), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n487), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n488), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n489), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n490), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n491), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n492), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n493), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n494), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n495), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n496), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n497), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n498), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n499), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n500), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n501), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n502), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n503), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n504), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n505), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n506), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n507), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n508), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n509), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n510), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n511), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n512), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n513), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n514), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n515), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n516), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n517), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n518), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n519), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n520), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n521), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n522), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n523), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n524), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n525), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n526), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n527), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n528), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n529), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n530), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n531), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n532), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n533), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n534), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n535), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n536), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n537), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n538), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .Q(data_out[3]) );
  DFF_X2 \data_out_reg[5]  ( .D(N16), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(N10), .Z(n398) );
  BUF_X1 U4 ( .A(N10), .Z(n399) );
  BUF_X1 U5 ( .A(N11), .Z(n396) );
  NAND2_X1 U6 ( .A1(n662), .A2(n682), .ZN(n671) );
  NAND2_X1 U7 ( .A1(n662), .A2(n672), .ZN(n661) );
  NAND2_X1 U8 ( .A1(n683), .A2(n682), .ZN(n692) );
  NAND2_X1 U9 ( .A1(n672), .A2(n683), .ZN(n681) );
  NAND2_X1 U10 ( .A1(n604), .A2(n683), .ZN(n613) );
  NAND2_X1 U11 ( .A1(n594), .A2(n683), .ZN(n603) );
  NAND2_X1 U12 ( .A1(n604), .A2(n662), .ZN(n593) );
  NAND2_X1 U13 ( .A1(n594), .A2(n662), .ZN(n584) );
  NAND2_X1 U14 ( .A1(n643), .A2(n682), .ZN(n652) );
  NAND2_X1 U15 ( .A1(n643), .A2(n672), .ZN(n642) );
  NAND2_X1 U16 ( .A1(n624), .A2(n682), .ZN(n633) );
  NAND2_X1 U17 ( .A1(n624), .A2(n672), .ZN(n622) );
  NAND2_X1 U18 ( .A1(n604), .A2(n643), .ZN(n575) );
  NAND2_X1 U19 ( .A1(n594), .A2(n643), .ZN(n566) );
  NAND2_X1 U20 ( .A1(n604), .A2(n624), .ZN(n557) );
  NAND2_X1 U21 ( .A1(n594), .A2(n624), .ZN(n547) );
  AND2_X1 U22 ( .A1(n548), .A2(N10), .ZN(n594) );
  AND2_X1 U23 ( .A1(n548), .A2(n400), .ZN(n604) );
  AND2_X1 U24 ( .A1(N10), .A2(n623), .ZN(n672) );
  AND2_X1 U25 ( .A1(n623), .A2(n400), .ZN(n682) );
  OAI21_X1 U26 ( .B1(n692), .B2(n410), .A(n691), .ZN(n538) );
  NAND2_X1 U27 ( .A1(\mem[0][0] ), .A2(n692), .ZN(n691) );
  OAI21_X1 U28 ( .B1(n692), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U29 ( .A1(\mem[0][1] ), .A2(n692), .ZN(n690) );
  OAI21_X1 U30 ( .B1(n692), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U31 ( .A1(\mem[0][2] ), .A2(n692), .ZN(n689) );
  OAI21_X1 U32 ( .B1(n692), .B2(n407), .A(n688), .ZN(n535) );
  NAND2_X1 U33 ( .A1(\mem[0][3] ), .A2(n692), .ZN(n688) );
  OAI21_X1 U34 ( .B1(n692), .B2(n406), .A(n687), .ZN(n534) );
  NAND2_X1 U35 ( .A1(\mem[0][4] ), .A2(n692), .ZN(n687) );
  OAI21_X1 U36 ( .B1(n692), .B2(n405), .A(n686), .ZN(n533) );
  NAND2_X1 U37 ( .A1(\mem[0][5] ), .A2(n692), .ZN(n686) );
  OAI21_X1 U38 ( .B1(n692), .B2(n404), .A(n685), .ZN(n532) );
  NAND2_X1 U39 ( .A1(\mem[0][6] ), .A2(n692), .ZN(n685) );
  OAI21_X1 U40 ( .B1(n692), .B2(n403), .A(n684), .ZN(n531) );
  NAND2_X1 U41 ( .A1(\mem[0][7] ), .A2(n692), .ZN(n684) );
  OAI21_X1 U42 ( .B1(n410), .B2(n671), .A(n670), .ZN(n522) );
  NAND2_X1 U43 ( .A1(\mem[2][0] ), .A2(n671), .ZN(n670) );
  OAI21_X1 U44 ( .B1(n409), .B2(n671), .A(n669), .ZN(n521) );
  NAND2_X1 U45 ( .A1(\mem[2][1] ), .A2(n671), .ZN(n669) );
  OAI21_X1 U46 ( .B1(n408), .B2(n671), .A(n668), .ZN(n520) );
  NAND2_X1 U47 ( .A1(\mem[2][2] ), .A2(n671), .ZN(n668) );
  OAI21_X1 U48 ( .B1(n407), .B2(n671), .A(n667), .ZN(n519) );
  NAND2_X1 U49 ( .A1(\mem[2][3] ), .A2(n671), .ZN(n667) );
  OAI21_X1 U50 ( .B1(n406), .B2(n671), .A(n666), .ZN(n518) );
  NAND2_X1 U51 ( .A1(\mem[2][4] ), .A2(n671), .ZN(n666) );
  OAI21_X1 U52 ( .B1(n405), .B2(n671), .A(n665), .ZN(n517) );
  NAND2_X1 U53 ( .A1(\mem[2][5] ), .A2(n671), .ZN(n665) );
  OAI21_X1 U54 ( .B1(n404), .B2(n671), .A(n664), .ZN(n516) );
  NAND2_X1 U55 ( .A1(\mem[2][6] ), .A2(n671), .ZN(n664) );
  OAI21_X1 U56 ( .B1(n403), .B2(n671), .A(n663), .ZN(n515) );
  NAND2_X1 U57 ( .A1(\mem[2][7] ), .A2(n671), .ZN(n663) );
  OAI21_X1 U58 ( .B1(n410), .B2(n661), .A(n660), .ZN(n514) );
  NAND2_X1 U59 ( .A1(\mem[3][0] ), .A2(n661), .ZN(n660) );
  OAI21_X1 U60 ( .B1(n409), .B2(n661), .A(n659), .ZN(n513) );
  NAND2_X1 U61 ( .A1(\mem[3][1] ), .A2(n661), .ZN(n659) );
  OAI21_X1 U62 ( .B1(n408), .B2(n661), .A(n658), .ZN(n512) );
  NAND2_X1 U63 ( .A1(\mem[3][2] ), .A2(n661), .ZN(n658) );
  OAI21_X1 U64 ( .B1(n407), .B2(n661), .A(n657), .ZN(n511) );
  NAND2_X1 U65 ( .A1(\mem[3][3] ), .A2(n661), .ZN(n657) );
  OAI21_X1 U66 ( .B1(n406), .B2(n661), .A(n656), .ZN(n510) );
  NAND2_X1 U67 ( .A1(\mem[3][4] ), .A2(n661), .ZN(n656) );
  OAI21_X1 U68 ( .B1(n405), .B2(n661), .A(n655), .ZN(n509) );
  NAND2_X1 U69 ( .A1(\mem[3][5] ), .A2(n661), .ZN(n655) );
  OAI21_X1 U70 ( .B1(n404), .B2(n661), .A(n654), .ZN(n508) );
  NAND2_X1 U71 ( .A1(\mem[3][6] ), .A2(n661), .ZN(n654) );
  OAI21_X1 U72 ( .B1(n403), .B2(n661), .A(n653), .ZN(n507) );
  NAND2_X1 U73 ( .A1(\mem[3][7] ), .A2(n661), .ZN(n653) );
  NOR2_X1 U74 ( .A1(n402), .A2(N13), .ZN(n623) );
  INV_X1 U75 ( .A(wr_en), .ZN(n402) );
  OAI21_X1 U76 ( .B1(n410), .B2(n681), .A(n680), .ZN(n530) );
  NAND2_X1 U77 ( .A1(\mem[1][0] ), .A2(n681), .ZN(n680) );
  OAI21_X1 U78 ( .B1(n409), .B2(n681), .A(n679), .ZN(n529) );
  NAND2_X1 U79 ( .A1(\mem[1][1] ), .A2(n681), .ZN(n679) );
  OAI21_X1 U80 ( .B1(n408), .B2(n681), .A(n678), .ZN(n528) );
  NAND2_X1 U81 ( .A1(\mem[1][2] ), .A2(n681), .ZN(n678) );
  OAI21_X1 U82 ( .B1(n407), .B2(n681), .A(n677), .ZN(n527) );
  NAND2_X1 U83 ( .A1(\mem[1][3] ), .A2(n681), .ZN(n677) );
  OAI21_X1 U84 ( .B1(n406), .B2(n681), .A(n676), .ZN(n526) );
  NAND2_X1 U85 ( .A1(\mem[1][4] ), .A2(n681), .ZN(n676) );
  OAI21_X1 U86 ( .B1(n405), .B2(n681), .A(n675), .ZN(n525) );
  NAND2_X1 U87 ( .A1(\mem[1][5] ), .A2(n681), .ZN(n675) );
  OAI21_X1 U88 ( .B1(n404), .B2(n681), .A(n674), .ZN(n524) );
  NAND2_X1 U89 ( .A1(\mem[1][6] ), .A2(n681), .ZN(n674) );
  OAI21_X1 U90 ( .B1(n403), .B2(n681), .A(n673), .ZN(n523) );
  NAND2_X1 U91 ( .A1(\mem[1][7] ), .A2(n681), .ZN(n673) );
  OAI21_X1 U92 ( .B1(n410), .B2(n652), .A(n651), .ZN(n506) );
  NAND2_X1 U93 ( .A1(\mem[4][0] ), .A2(n652), .ZN(n651) );
  OAI21_X1 U94 ( .B1(n409), .B2(n652), .A(n650), .ZN(n505) );
  NAND2_X1 U95 ( .A1(\mem[4][1] ), .A2(n652), .ZN(n650) );
  OAI21_X1 U96 ( .B1(n408), .B2(n652), .A(n649), .ZN(n504) );
  NAND2_X1 U97 ( .A1(\mem[4][2] ), .A2(n652), .ZN(n649) );
  OAI21_X1 U98 ( .B1(n407), .B2(n652), .A(n648), .ZN(n503) );
  NAND2_X1 U99 ( .A1(\mem[4][3] ), .A2(n652), .ZN(n648) );
  OAI21_X1 U100 ( .B1(n406), .B2(n652), .A(n647), .ZN(n502) );
  NAND2_X1 U101 ( .A1(\mem[4][4] ), .A2(n652), .ZN(n647) );
  OAI21_X1 U102 ( .B1(n405), .B2(n652), .A(n646), .ZN(n501) );
  NAND2_X1 U103 ( .A1(\mem[4][5] ), .A2(n652), .ZN(n646) );
  OAI21_X1 U104 ( .B1(n404), .B2(n652), .A(n645), .ZN(n500) );
  NAND2_X1 U105 ( .A1(\mem[4][6] ), .A2(n652), .ZN(n645) );
  OAI21_X1 U106 ( .B1(n403), .B2(n652), .A(n644), .ZN(n499) );
  NAND2_X1 U107 ( .A1(\mem[4][7] ), .A2(n652), .ZN(n644) );
  OAI21_X1 U108 ( .B1(n410), .B2(n642), .A(n641), .ZN(n498) );
  NAND2_X1 U109 ( .A1(\mem[5][0] ), .A2(n642), .ZN(n641) );
  OAI21_X1 U110 ( .B1(n409), .B2(n642), .A(n640), .ZN(n497) );
  NAND2_X1 U111 ( .A1(\mem[5][1] ), .A2(n642), .ZN(n640) );
  OAI21_X1 U112 ( .B1(n408), .B2(n642), .A(n639), .ZN(n496) );
  NAND2_X1 U113 ( .A1(\mem[5][2] ), .A2(n642), .ZN(n639) );
  OAI21_X1 U114 ( .B1(n407), .B2(n642), .A(n638), .ZN(n495) );
  NAND2_X1 U115 ( .A1(\mem[5][3] ), .A2(n642), .ZN(n638) );
  OAI21_X1 U116 ( .B1(n406), .B2(n642), .A(n637), .ZN(n494) );
  NAND2_X1 U117 ( .A1(\mem[5][4] ), .A2(n642), .ZN(n637) );
  OAI21_X1 U118 ( .B1(n405), .B2(n642), .A(n636), .ZN(n493) );
  NAND2_X1 U119 ( .A1(\mem[5][5] ), .A2(n642), .ZN(n636) );
  OAI21_X1 U120 ( .B1(n404), .B2(n642), .A(n635), .ZN(n492) );
  NAND2_X1 U121 ( .A1(\mem[5][6] ), .A2(n642), .ZN(n635) );
  OAI21_X1 U122 ( .B1(n403), .B2(n642), .A(n634), .ZN(n491) );
  NAND2_X1 U123 ( .A1(\mem[5][7] ), .A2(n642), .ZN(n634) );
  OAI21_X1 U124 ( .B1(n410), .B2(n633), .A(n632), .ZN(n490) );
  NAND2_X1 U125 ( .A1(\mem[6][0] ), .A2(n633), .ZN(n632) );
  OAI21_X1 U126 ( .B1(n409), .B2(n633), .A(n631), .ZN(n489) );
  NAND2_X1 U127 ( .A1(\mem[6][1] ), .A2(n633), .ZN(n631) );
  OAI21_X1 U128 ( .B1(n408), .B2(n633), .A(n630), .ZN(n488) );
  NAND2_X1 U129 ( .A1(\mem[6][2] ), .A2(n633), .ZN(n630) );
  OAI21_X1 U130 ( .B1(n407), .B2(n633), .A(n629), .ZN(n487) );
  NAND2_X1 U131 ( .A1(\mem[6][3] ), .A2(n633), .ZN(n629) );
  OAI21_X1 U132 ( .B1(n406), .B2(n633), .A(n628), .ZN(n486) );
  NAND2_X1 U133 ( .A1(\mem[6][4] ), .A2(n633), .ZN(n628) );
  OAI21_X1 U134 ( .B1(n405), .B2(n633), .A(n627), .ZN(n485) );
  NAND2_X1 U135 ( .A1(\mem[6][5] ), .A2(n633), .ZN(n627) );
  OAI21_X1 U136 ( .B1(n404), .B2(n633), .A(n626), .ZN(n484) );
  NAND2_X1 U137 ( .A1(\mem[6][6] ), .A2(n633), .ZN(n626) );
  OAI21_X1 U138 ( .B1(n403), .B2(n633), .A(n625), .ZN(n483) );
  NAND2_X1 U139 ( .A1(\mem[6][7] ), .A2(n633), .ZN(n625) );
  OAI21_X1 U140 ( .B1(n410), .B2(n622), .A(n621), .ZN(n482) );
  NAND2_X1 U141 ( .A1(\mem[7][0] ), .A2(n622), .ZN(n621) );
  OAI21_X1 U142 ( .B1(n409), .B2(n622), .A(n620), .ZN(n481) );
  NAND2_X1 U143 ( .A1(\mem[7][1] ), .A2(n622), .ZN(n620) );
  OAI21_X1 U144 ( .B1(n408), .B2(n622), .A(n619), .ZN(n480) );
  NAND2_X1 U145 ( .A1(\mem[7][2] ), .A2(n622), .ZN(n619) );
  OAI21_X1 U146 ( .B1(n407), .B2(n622), .A(n618), .ZN(n479) );
  NAND2_X1 U147 ( .A1(\mem[7][3] ), .A2(n622), .ZN(n618) );
  OAI21_X1 U148 ( .B1(n406), .B2(n622), .A(n617), .ZN(n478) );
  NAND2_X1 U149 ( .A1(\mem[7][4] ), .A2(n622), .ZN(n617) );
  OAI21_X1 U150 ( .B1(n405), .B2(n622), .A(n616), .ZN(n477) );
  NAND2_X1 U151 ( .A1(\mem[7][5] ), .A2(n622), .ZN(n616) );
  OAI21_X1 U152 ( .B1(n404), .B2(n622), .A(n615), .ZN(n476) );
  NAND2_X1 U153 ( .A1(\mem[7][6] ), .A2(n622), .ZN(n615) );
  OAI21_X1 U154 ( .B1(n403), .B2(n622), .A(n614), .ZN(n475) );
  NAND2_X1 U155 ( .A1(\mem[7][7] ), .A2(n622), .ZN(n614) );
  OAI21_X1 U156 ( .B1(n410), .B2(n613), .A(n612), .ZN(n474) );
  NAND2_X1 U157 ( .A1(\mem[8][0] ), .A2(n613), .ZN(n612) );
  OAI21_X1 U158 ( .B1(n409), .B2(n613), .A(n611), .ZN(n473) );
  NAND2_X1 U159 ( .A1(\mem[8][1] ), .A2(n613), .ZN(n611) );
  OAI21_X1 U160 ( .B1(n408), .B2(n613), .A(n610), .ZN(n472) );
  NAND2_X1 U161 ( .A1(\mem[8][2] ), .A2(n613), .ZN(n610) );
  OAI21_X1 U162 ( .B1(n407), .B2(n613), .A(n609), .ZN(n471) );
  NAND2_X1 U163 ( .A1(\mem[8][3] ), .A2(n613), .ZN(n609) );
  OAI21_X1 U164 ( .B1(n406), .B2(n613), .A(n608), .ZN(n470) );
  NAND2_X1 U165 ( .A1(\mem[8][4] ), .A2(n613), .ZN(n608) );
  OAI21_X1 U166 ( .B1(n405), .B2(n613), .A(n607), .ZN(n469) );
  NAND2_X1 U167 ( .A1(\mem[8][5] ), .A2(n613), .ZN(n607) );
  OAI21_X1 U168 ( .B1(n404), .B2(n613), .A(n606), .ZN(n468) );
  NAND2_X1 U169 ( .A1(\mem[8][6] ), .A2(n613), .ZN(n606) );
  OAI21_X1 U170 ( .B1(n403), .B2(n613), .A(n605), .ZN(n467) );
  NAND2_X1 U171 ( .A1(\mem[8][7] ), .A2(n613), .ZN(n605) );
  OAI21_X1 U172 ( .B1(n410), .B2(n603), .A(n602), .ZN(n466) );
  NAND2_X1 U173 ( .A1(\mem[9][0] ), .A2(n603), .ZN(n602) );
  OAI21_X1 U174 ( .B1(n409), .B2(n603), .A(n601), .ZN(n465) );
  NAND2_X1 U175 ( .A1(\mem[9][1] ), .A2(n603), .ZN(n601) );
  OAI21_X1 U176 ( .B1(n408), .B2(n603), .A(n600), .ZN(n464) );
  NAND2_X1 U177 ( .A1(\mem[9][2] ), .A2(n603), .ZN(n600) );
  OAI21_X1 U178 ( .B1(n407), .B2(n603), .A(n599), .ZN(n463) );
  NAND2_X1 U179 ( .A1(\mem[9][3] ), .A2(n603), .ZN(n599) );
  OAI21_X1 U180 ( .B1(n406), .B2(n603), .A(n598), .ZN(n462) );
  NAND2_X1 U181 ( .A1(\mem[9][4] ), .A2(n603), .ZN(n598) );
  OAI21_X1 U182 ( .B1(n405), .B2(n603), .A(n597), .ZN(n461) );
  NAND2_X1 U183 ( .A1(\mem[9][5] ), .A2(n603), .ZN(n597) );
  OAI21_X1 U184 ( .B1(n404), .B2(n603), .A(n596), .ZN(n460) );
  NAND2_X1 U185 ( .A1(\mem[9][6] ), .A2(n603), .ZN(n596) );
  OAI21_X1 U186 ( .B1(n403), .B2(n603), .A(n595), .ZN(n459) );
  NAND2_X1 U187 ( .A1(\mem[9][7] ), .A2(n603), .ZN(n595) );
  OAI21_X1 U188 ( .B1(n410), .B2(n593), .A(n592), .ZN(n458) );
  NAND2_X1 U189 ( .A1(\mem[10][0] ), .A2(n593), .ZN(n592) );
  OAI21_X1 U190 ( .B1(n409), .B2(n593), .A(n591), .ZN(n457) );
  NAND2_X1 U191 ( .A1(\mem[10][1] ), .A2(n593), .ZN(n591) );
  OAI21_X1 U192 ( .B1(n408), .B2(n593), .A(n590), .ZN(n456) );
  NAND2_X1 U193 ( .A1(\mem[10][2] ), .A2(n593), .ZN(n590) );
  OAI21_X1 U194 ( .B1(n407), .B2(n593), .A(n589), .ZN(n455) );
  NAND2_X1 U195 ( .A1(\mem[10][3] ), .A2(n593), .ZN(n589) );
  OAI21_X1 U196 ( .B1(n406), .B2(n593), .A(n588), .ZN(n454) );
  NAND2_X1 U197 ( .A1(\mem[10][4] ), .A2(n593), .ZN(n588) );
  OAI21_X1 U198 ( .B1(n405), .B2(n593), .A(n587), .ZN(n453) );
  NAND2_X1 U199 ( .A1(\mem[10][5] ), .A2(n593), .ZN(n587) );
  OAI21_X1 U200 ( .B1(n404), .B2(n593), .A(n586), .ZN(n452) );
  NAND2_X1 U201 ( .A1(\mem[10][6] ), .A2(n593), .ZN(n586) );
  OAI21_X1 U202 ( .B1(n403), .B2(n593), .A(n585), .ZN(n451) );
  NAND2_X1 U203 ( .A1(\mem[10][7] ), .A2(n593), .ZN(n585) );
  OAI21_X1 U204 ( .B1(n410), .B2(n584), .A(n583), .ZN(n450) );
  NAND2_X1 U205 ( .A1(\mem[11][0] ), .A2(n584), .ZN(n583) );
  OAI21_X1 U206 ( .B1(n409), .B2(n584), .A(n582), .ZN(n449) );
  NAND2_X1 U207 ( .A1(\mem[11][1] ), .A2(n584), .ZN(n582) );
  OAI21_X1 U208 ( .B1(n408), .B2(n584), .A(n581), .ZN(n448) );
  NAND2_X1 U209 ( .A1(\mem[11][2] ), .A2(n584), .ZN(n581) );
  OAI21_X1 U210 ( .B1(n407), .B2(n584), .A(n580), .ZN(n447) );
  NAND2_X1 U211 ( .A1(\mem[11][3] ), .A2(n584), .ZN(n580) );
  OAI21_X1 U212 ( .B1(n406), .B2(n584), .A(n579), .ZN(n446) );
  NAND2_X1 U213 ( .A1(\mem[11][4] ), .A2(n584), .ZN(n579) );
  OAI21_X1 U214 ( .B1(n405), .B2(n584), .A(n578), .ZN(n445) );
  NAND2_X1 U215 ( .A1(\mem[11][5] ), .A2(n584), .ZN(n578) );
  OAI21_X1 U216 ( .B1(n404), .B2(n584), .A(n577), .ZN(n444) );
  NAND2_X1 U217 ( .A1(\mem[11][6] ), .A2(n584), .ZN(n577) );
  OAI21_X1 U218 ( .B1(n403), .B2(n584), .A(n576), .ZN(n443) );
  NAND2_X1 U219 ( .A1(\mem[11][7] ), .A2(n584), .ZN(n576) );
  OAI21_X1 U220 ( .B1(n410), .B2(n575), .A(n574), .ZN(n442) );
  NAND2_X1 U221 ( .A1(\mem[12][0] ), .A2(n575), .ZN(n574) );
  OAI21_X1 U222 ( .B1(n409), .B2(n575), .A(n573), .ZN(n441) );
  NAND2_X1 U223 ( .A1(\mem[12][1] ), .A2(n575), .ZN(n573) );
  OAI21_X1 U224 ( .B1(n408), .B2(n575), .A(n572), .ZN(n440) );
  NAND2_X1 U225 ( .A1(\mem[12][2] ), .A2(n575), .ZN(n572) );
  OAI21_X1 U226 ( .B1(n407), .B2(n575), .A(n571), .ZN(n439) );
  NAND2_X1 U227 ( .A1(\mem[12][3] ), .A2(n575), .ZN(n571) );
  OAI21_X1 U228 ( .B1(n406), .B2(n575), .A(n570), .ZN(n438) );
  NAND2_X1 U229 ( .A1(\mem[12][4] ), .A2(n575), .ZN(n570) );
  OAI21_X1 U230 ( .B1(n405), .B2(n575), .A(n569), .ZN(n437) );
  NAND2_X1 U231 ( .A1(\mem[12][5] ), .A2(n575), .ZN(n569) );
  OAI21_X1 U232 ( .B1(n404), .B2(n575), .A(n568), .ZN(n436) );
  NAND2_X1 U233 ( .A1(\mem[12][6] ), .A2(n575), .ZN(n568) );
  OAI21_X1 U234 ( .B1(n403), .B2(n575), .A(n567), .ZN(n435) );
  NAND2_X1 U235 ( .A1(\mem[12][7] ), .A2(n575), .ZN(n567) );
  OAI21_X1 U236 ( .B1(n410), .B2(n566), .A(n565), .ZN(n434) );
  NAND2_X1 U237 ( .A1(\mem[13][0] ), .A2(n566), .ZN(n565) );
  OAI21_X1 U238 ( .B1(n409), .B2(n566), .A(n564), .ZN(n433) );
  NAND2_X1 U239 ( .A1(\mem[13][1] ), .A2(n566), .ZN(n564) );
  OAI21_X1 U240 ( .B1(n408), .B2(n566), .A(n563), .ZN(n432) );
  NAND2_X1 U241 ( .A1(\mem[13][2] ), .A2(n566), .ZN(n563) );
  OAI21_X1 U242 ( .B1(n407), .B2(n566), .A(n562), .ZN(n431) );
  NAND2_X1 U243 ( .A1(\mem[13][3] ), .A2(n566), .ZN(n562) );
  OAI21_X1 U244 ( .B1(n406), .B2(n566), .A(n561), .ZN(n430) );
  NAND2_X1 U245 ( .A1(\mem[13][4] ), .A2(n566), .ZN(n561) );
  OAI21_X1 U246 ( .B1(n405), .B2(n566), .A(n560), .ZN(n429) );
  NAND2_X1 U247 ( .A1(\mem[13][5] ), .A2(n566), .ZN(n560) );
  OAI21_X1 U248 ( .B1(n404), .B2(n566), .A(n559), .ZN(n428) );
  NAND2_X1 U249 ( .A1(\mem[13][6] ), .A2(n566), .ZN(n559) );
  OAI21_X1 U250 ( .B1(n403), .B2(n566), .A(n558), .ZN(n427) );
  NAND2_X1 U251 ( .A1(\mem[13][7] ), .A2(n566), .ZN(n558) );
  OAI21_X1 U252 ( .B1(n410), .B2(n557), .A(n556), .ZN(n426) );
  NAND2_X1 U253 ( .A1(\mem[14][0] ), .A2(n557), .ZN(n556) );
  OAI21_X1 U254 ( .B1(n409), .B2(n557), .A(n555), .ZN(n425) );
  NAND2_X1 U255 ( .A1(\mem[14][1] ), .A2(n557), .ZN(n555) );
  OAI21_X1 U256 ( .B1(n408), .B2(n557), .A(n554), .ZN(n424) );
  NAND2_X1 U257 ( .A1(\mem[14][2] ), .A2(n557), .ZN(n554) );
  OAI21_X1 U258 ( .B1(n407), .B2(n557), .A(n553), .ZN(n423) );
  NAND2_X1 U259 ( .A1(\mem[14][3] ), .A2(n557), .ZN(n553) );
  OAI21_X1 U260 ( .B1(n406), .B2(n557), .A(n552), .ZN(n422) );
  NAND2_X1 U261 ( .A1(\mem[14][4] ), .A2(n557), .ZN(n552) );
  OAI21_X1 U262 ( .B1(n405), .B2(n557), .A(n551), .ZN(n421) );
  NAND2_X1 U263 ( .A1(\mem[14][5] ), .A2(n557), .ZN(n551) );
  OAI21_X1 U264 ( .B1(n404), .B2(n557), .A(n550), .ZN(n420) );
  NAND2_X1 U265 ( .A1(\mem[14][6] ), .A2(n557), .ZN(n550) );
  OAI21_X1 U266 ( .B1(n403), .B2(n557), .A(n549), .ZN(n419) );
  NAND2_X1 U267 ( .A1(\mem[14][7] ), .A2(n557), .ZN(n549) );
  OAI21_X1 U268 ( .B1(n410), .B2(n547), .A(n546), .ZN(n418) );
  NAND2_X1 U269 ( .A1(\mem[15][0] ), .A2(n547), .ZN(n546) );
  OAI21_X1 U270 ( .B1(n409), .B2(n547), .A(n545), .ZN(n417) );
  NAND2_X1 U271 ( .A1(\mem[15][1] ), .A2(n547), .ZN(n545) );
  OAI21_X1 U272 ( .B1(n408), .B2(n547), .A(n544), .ZN(n416) );
  NAND2_X1 U273 ( .A1(\mem[15][2] ), .A2(n547), .ZN(n544) );
  OAI21_X1 U274 ( .B1(n407), .B2(n547), .A(n543), .ZN(n415) );
  NAND2_X1 U275 ( .A1(\mem[15][3] ), .A2(n547), .ZN(n543) );
  OAI21_X1 U276 ( .B1(n406), .B2(n547), .A(n542), .ZN(n414) );
  NAND2_X1 U277 ( .A1(\mem[15][4] ), .A2(n547), .ZN(n542) );
  OAI21_X1 U278 ( .B1(n405), .B2(n547), .A(n541), .ZN(n413) );
  NAND2_X1 U279 ( .A1(\mem[15][5] ), .A2(n547), .ZN(n541) );
  OAI21_X1 U280 ( .B1(n404), .B2(n547), .A(n540), .ZN(n412) );
  NAND2_X1 U281 ( .A1(\mem[15][6] ), .A2(n547), .ZN(n540) );
  OAI21_X1 U282 ( .B1(n403), .B2(n547), .A(n539), .ZN(n411) );
  NAND2_X1 U283 ( .A1(\mem[15][7] ), .A2(n547), .ZN(n539) );
  AND2_X1 U284 ( .A1(N13), .A2(wr_en), .ZN(n548) );
  NOR2_X1 U285 ( .A1(N11), .A2(N12), .ZN(n683) );
  NOR2_X1 U286 ( .A1(n401), .A2(N12), .ZN(n662) );
  AND2_X1 U287 ( .A1(N12), .A2(n401), .ZN(n643) );
  AND2_X1 U288 ( .A1(N12), .A2(N11), .ZN(n624) );
  INV_X1 U289 ( .A(data_in[0]), .ZN(n410) );
  INV_X1 U290 ( .A(data_in[1]), .ZN(n409) );
  INV_X1 U291 ( .A(data_in[2]), .ZN(n408) );
  INV_X1 U292 ( .A(data_in[3]), .ZN(n407) );
  INV_X1 U293 ( .A(data_in[4]), .ZN(n406) );
  INV_X1 U294 ( .A(data_in[5]), .ZN(n405) );
  INV_X1 U295 ( .A(data_in[6]), .ZN(n404) );
  INV_X1 U296 ( .A(data_in[7]), .ZN(n403) );
  MUX2_X1 U297 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n397), .Z(n2) );
  MUX2_X1 U298 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n397), .Z(n3) );
  MUX2_X1 U299 ( .A(n3), .B(n2), .S(N11), .Z(n4) );
  MUX2_X1 U300 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n397), .Z(n5) );
  MUX2_X1 U301 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n397), .Z(n6) );
  MUX2_X1 U302 ( .A(n6), .B(n5), .S(N11), .Z(n7) );
  MUX2_X1 U303 ( .A(n7), .B(n4), .S(N12), .Z(n8) );
  MUX2_X1 U304 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n398), .Z(n9) );
  MUX2_X1 U305 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n398), .Z(n10) );
  MUX2_X1 U306 ( .A(n10), .B(n9), .S(N11), .Z(n11) );
  MUX2_X1 U307 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n398), .Z(n294) );
  MUX2_X1 U308 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n398), .Z(n295) );
  MUX2_X1 U309 ( .A(n295), .B(n294), .S(N11), .Z(n296) );
  MUX2_X1 U310 ( .A(n296), .B(n11), .S(N12), .Z(n297) );
  MUX2_X1 U311 ( .A(n297), .B(n8), .S(N13), .Z(N21) );
  MUX2_X1 U312 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n398), .Z(n298) );
  MUX2_X1 U313 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n398), .Z(n299) );
  MUX2_X1 U314 ( .A(n299), .B(n298), .S(N11), .Z(n300) );
  MUX2_X1 U315 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n398), .Z(n301) );
  MUX2_X1 U316 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n398), .Z(n302) );
  MUX2_X1 U317 ( .A(n302), .B(n301), .S(N11), .Z(n303) );
  MUX2_X1 U318 ( .A(n303), .B(n300), .S(N12), .Z(n304) );
  MUX2_X1 U319 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n398), .Z(n305) );
  MUX2_X1 U320 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n398), .Z(n306) );
  MUX2_X1 U321 ( .A(n306), .B(n305), .S(N11), .Z(n307) );
  MUX2_X1 U322 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n398), .Z(n308) );
  MUX2_X1 U323 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n398), .Z(n309) );
  MUX2_X1 U324 ( .A(n309), .B(n308), .S(N11), .Z(n310) );
  MUX2_X1 U325 ( .A(n310), .B(n307), .S(N12), .Z(n311) );
  MUX2_X1 U326 ( .A(n311), .B(n304), .S(N13), .Z(N20) );
  MUX2_X1 U327 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n399), .Z(n312) );
  MUX2_X1 U328 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n399), .Z(n313) );
  MUX2_X1 U329 ( .A(n313), .B(n312), .S(n396), .Z(n314) );
  MUX2_X1 U330 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n399), .Z(n315) );
  MUX2_X1 U331 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n399), .Z(n316) );
  MUX2_X1 U332 ( .A(n316), .B(n315), .S(n396), .Z(n317) );
  MUX2_X1 U333 ( .A(n317), .B(n314), .S(N12), .Z(n318) );
  MUX2_X1 U334 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n399), .Z(n319) );
  MUX2_X1 U335 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n399), .Z(n320) );
  MUX2_X1 U336 ( .A(n320), .B(n319), .S(n396), .Z(n321) );
  MUX2_X1 U337 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n399), .Z(n322) );
  MUX2_X1 U338 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n399), .Z(n323) );
  MUX2_X1 U339 ( .A(n323), .B(n322), .S(n396), .Z(n324) );
  MUX2_X1 U340 ( .A(n324), .B(n321), .S(N12), .Z(n325) );
  MUX2_X1 U341 ( .A(n325), .B(n318), .S(N13), .Z(N19) );
  MUX2_X1 U342 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n399), .Z(n326) );
  MUX2_X1 U343 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n399), .Z(n327) );
  MUX2_X1 U344 ( .A(n327), .B(n326), .S(n396), .Z(n328) );
  MUX2_X1 U345 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n399), .Z(n329) );
  MUX2_X1 U346 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n399), .Z(n330) );
  MUX2_X1 U347 ( .A(n330), .B(n329), .S(n396), .Z(n331) );
  MUX2_X1 U348 ( .A(n331), .B(n328), .S(N12), .Z(n332) );
  MUX2_X1 U349 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n398), .Z(n333) );
  MUX2_X1 U350 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n398), .Z(n334) );
  MUX2_X1 U351 ( .A(n334), .B(n333), .S(n396), .Z(n335) );
  MUX2_X1 U352 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n336) );
  MUX2_X1 U353 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n398), .Z(n337) );
  MUX2_X1 U354 ( .A(n337), .B(n336), .S(n396), .Z(n338) );
  MUX2_X1 U355 ( .A(n338), .B(n335), .S(N12), .Z(n339) );
  MUX2_X1 U356 ( .A(n339), .B(n332), .S(N13), .Z(N18) );
  MUX2_X1 U357 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n399), .Z(n340) );
  MUX2_X1 U358 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(N10), .Z(n341) );
  MUX2_X1 U359 ( .A(n341), .B(n340), .S(n396), .Z(n342) );
  MUX2_X1 U360 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n398), .Z(n343) );
  MUX2_X1 U361 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n399), .Z(n344) );
  MUX2_X1 U362 ( .A(n344), .B(n343), .S(n396), .Z(n345) );
  MUX2_X1 U363 ( .A(n345), .B(n342), .S(N12), .Z(n346) );
  MUX2_X1 U364 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n399), .Z(n347) );
  MUX2_X1 U365 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n397), .Z(n348) );
  MUX2_X1 U366 ( .A(n348), .B(n347), .S(n396), .Z(n349) );
  MUX2_X1 U367 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n397), .Z(n350) );
  MUX2_X1 U368 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n397), .Z(n351) );
  MUX2_X1 U369 ( .A(n351), .B(n350), .S(n396), .Z(n352) );
  MUX2_X1 U370 ( .A(n352), .B(n349), .S(N12), .Z(n353) );
  MUX2_X1 U371 ( .A(n353), .B(n346), .S(N13), .Z(N17) );
  MUX2_X1 U372 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n397), .Z(n354) );
  MUX2_X1 U373 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(N10), .Z(n355) );
  MUX2_X1 U374 ( .A(n355), .B(n354), .S(N11), .Z(n356) );
  MUX2_X1 U375 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(N10), .Z(n357) );
  MUX2_X1 U376 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(N10), .Z(n358) );
  MUX2_X1 U377 ( .A(n358), .B(n357), .S(N11), .Z(n359) );
  MUX2_X1 U378 ( .A(n359), .B(n356), .S(N12), .Z(n360) );
  MUX2_X1 U379 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(N10), .Z(n361) );
  MUX2_X1 U380 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(N10), .Z(n362) );
  MUX2_X1 U381 ( .A(n362), .B(n361), .S(N11), .Z(n363) );
  MUX2_X1 U382 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n364) );
  MUX2_X1 U383 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(N10), .Z(n365) );
  MUX2_X1 U384 ( .A(n365), .B(n364), .S(N11), .Z(n366) );
  MUX2_X1 U385 ( .A(n366), .B(n363), .S(N12), .Z(n367) );
  MUX2_X1 U386 ( .A(n367), .B(n360), .S(N13), .Z(N16) );
  MUX2_X1 U387 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(N10), .Z(n368) );
  MUX2_X1 U388 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(N10), .Z(n369) );
  MUX2_X1 U389 ( .A(n369), .B(n368), .S(N11), .Z(n370) );
  MUX2_X1 U390 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(N10), .Z(n371) );
  MUX2_X1 U391 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n372) );
  MUX2_X1 U392 ( .A(n372), .B(n371), .S(N11), .Z(n373) );
  MUX2_X1 U393 ( .A(n373), .B(n370), .S(N12), .Z(n374) );
  MUX2_X1 U394 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n397), .Z(n375) );
  MUX2_X1 U395 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n397), .Z(n376) );
  MUX2_X1 U396 ( .A(n376), .B(n375), .S(N11), .Z(n377) );
  MUX2_X1 U397 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n399), .Z(n378) );
  MUX2_X1 U398 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n379) );
  MUX2_X1 U399 ( .A(n379), .B(n378), .S(n396), .Z(n380) );
  MUX2_X1 U400 ( .A(n380), .B(n377), .S(N12), .Z(n381) );
  MUX2_X1 U401 ( .A(n381), .B(n374), .S(N13), .Z(N15) );
  MUX2_X1 U402 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n397), .Z(n382) );
  MUX2_X1 U403 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n397), .Z(n383) );
  MUX2_X1 U404 ( .A(n383), .B(n382), .S(N11), .Z(n384) );
  MUX2_X1 U405 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n397), .Z(n385) );
  MUX2_X1 U406 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n398), .Z(n386) );
  MUX2_X1 U407 ( .A(n386), .B(n385), .S(n396), .Z(n387) );
  MUX2_X1 U408 ( .A(n387), .B(n384), .S(N12), .Z(n388) );
  MUX2_X1 U409 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n397), .Z(n389) );
  MUX2_X1 U410 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n397), .Z(n390) );
  MUX2_X1 U411 ( .A(n390), .B(n389), .S(N11), .Z(n391) );
  MUX2_X1 U412 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n399), .Z(n392) );
  MUX2_X1 U413 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n393) );
  MUX2_X1 U414 ( .A(n393), .B(n392), .S(n396), .Z(n394) );
  MUX2_X1 U415 ( .A(n394), .B(n391), .S(N12), .Z(n395) );
  MUX2_X1 U416 ( .A(n395), .B(n388), .S(N13), .Z(N14) );
  CLKBUF_X1 U417 ( .A(N10), .Z(n397) );
  INV_X1 U418 ( .A(N10), .ZN(n400) );
  INV_X1 U419 ( .A(N11), .ZN(n401) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_6 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, N19, N20, N21, n1, n3, n5, n6, n7, n8, n9, n10,
         n11, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n414), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n415), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n416), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n417), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n418), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n419), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n420), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n421), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n422), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n423), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n424), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n425), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n426), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n427), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n428), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n429), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n430), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n431), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n432), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n433), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n434), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n435), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n436), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n437), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n438), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n439), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n440), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n441), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n442), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n443), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n444), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n445), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n446), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n447), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n448), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n449), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n450), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n451), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n452), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n453), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n454), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n455), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n456), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n457), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n458), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n459), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n460), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n461), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n462), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n463), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n464), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n465), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n466), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n467), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n468), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n469), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n470), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n471), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n472), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n473), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n474), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n475), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n476), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n477), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n478), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n479), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n480), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n481), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n482), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n483), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n484), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n485), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n486), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n487), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n488), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n489), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n490), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n491), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n492), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n493), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n494), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n495), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n496), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n497), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n498), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n499), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n500), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n501), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n502), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n503), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n504), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n505), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n506), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n507), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n508), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n509), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n510), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n511), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n512), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n513), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n514), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n515), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n516), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n517), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n518), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n519), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n520), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n521), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n522), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n523), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n524), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n525), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n526), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n527), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n528), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n529), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n530), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n531), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n532), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n533), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n534), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n535), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n536), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n537), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n538), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n539), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n540), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n541), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N20), .CK(clk), .QN(n3) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .QN(n1) );
  DFF_X2 \data_out_reg[5]  ( .D(N16), .CK(clk), .Q(data_out[5]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  INV_X2 U4 ( .A(n3), .ZN(data_out[1]) );
  BUF_X1 U5 ( .A(N10), .Z(n400) );
  BUF_X1 U6 ( .A(N10), .Z(n401) );
  BUF_X1 U7 ( .A(N10), .Z(n402) );
  BUF_X1 U8 ( .A(N11), .Z(n399) );
  NAND2_X1 U9 ( .A1(n665), .A2(n685), .ZN(n674) );
  NAND2_X1 U10 ( .A1(n665), .A2(n675), .ZN(n664) );
  NAND2_X1 U11 ( .A1(n686), .A2(n685), .ZN(n695) );
  NAND2_X1 U12 ( .A1(n675), .A2(n686), .ZN(n684) );
  NAND2_X1 U13 ( .A1(n607), .A2(n686), .ZN(n616) );
  NAND2_X1 U14 ( .A1(n597), .A2(n686), .ZN(n606) );
  NAND2_X1 U15 ( .A1(n607), .A2(n665), .ZN(n596) );
  NAND2_X1 U16 ( .A1(n597), .A2(n665), .ZN(n587) );
  NAND2_X1 U17 ( .A1(n646), .A2(n685), .ZN(n655) );
  NAND2_X1 U18 ( .A1(n646), .A2(n675), .ZN(n645) );
  NAND2_X1 U19 ( .A1(n627), .A2(n685), .ZN(n636) );
  NAND2_X1 U20 ( .A1(n627), .A2(n675), .ZN(n625) );
  NAND2_X1 U21 ( .A1(n607), .A2(n646), .ZN(n578) );
  NAND2_X1 U22 ( .A1(n597), .A2(n646), .ZN(n569) );
  NAND2_X1 U23 ( .A1(n607), .A2(n627), .ZN(n560) );
  NAND2_X1 U24 ( .A1(n597), .A2(n627), .ZN(n550) );
  AND2_X1 U25 ( .A1(n551), .A2(N10), .ZN(n597) );
  AND2_X1 U26 ( .A1(n551), .A2(n403), .ZN(n607) );
  AND2_X1 U27 ( .A1(N10), .A2(n626), .ZN(n675) );
  AND2_X1 U28 ( .A1(n626), .A2(n403), .ZN(n685) );
  OAI21_X1 U29 ( .B1(n695), .B2(n413), .A(n694), .ZN(n541) );
  NAND2_X1 U30 ( .A1(\mem[0][0] ), .A2(n695), .ZN(n694) );
  OAI21_X1 U31 ( .B1(n695), .B2(n412), .A(n693), .ZN(n540) );
  NAND2_X1 U32 ( .A1(\mem[0][1] ), .A2(n695), .ZN(n693) );
  OAI21_X1 U33 ( .B1(n695), .B2(n411), .A(n692), .ZN(n539) );
  NAND2_X1 U34 ( .A1(\mem[0][2] ), .A2(n695), .ZN(n692) );
  OAI21_X1 U35 ( .B1(n695), .B2(n410), .A(n691), .ZN(n538) );
  NAND2_X1 U36 ( .A1(\mem[0][3] ), .A2(n695), .ZN(n691) );
  OAI21_X1 U37 ( .B1(n695), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U38 ( .A1(\mem[0][4] ), .A2(n695), .ZN(n690) );
  OAI21_X1 U39 ( .B1(n695), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U40 ( .A1(\mem[0][5] ), .A2(n695), .ZN(n689) );
  OAI21_X1 U41 ( .B1(n695), .B2(n407), .A(n688), .ZN(n535) );
  NAND2_X1 U42 ( .A1(\mem[0][6] ), .A2(n695), .ZN(n688) );
  OAI21_X1 U43 ( .B1(n695), .B2(n406), .A(n687), .ZN(n534) );
  NAND2_X1 U44 ( .A1(\mem[0][7] ), .A2(n695), .ZN(n687) );
  OAI21_X1 U45 ( .B1(n413), .B2(n674), .A(n673), .ZN(n525) );
  NAND2_X1 U46 ( .A1(\mem[2][0] ), .A2(n674), .ZN(n673) );
  OAI21_X1 U47 ( .B1(n412), .B2(n674), .A(n672), .ZN(n524) );
  NAND2_X1 U48 ( .A1(\mem[2][1] ), .A2(n674), .ZN(n672) );
  OAI21_X1 U49 ( .B1(n411), .B2(n674), .A(n671), .ZN(n523) );
  NAND2_X1 U50 ( .A1(\mem[2][2] ), .A2(n674), .ZN(n671) );
  OAI21_X1 U51 ( .B1(n410), .B2(n674), .A(n670), .ZN(n522) );
  NAND2_X1 U52 ( .A1(\mem[2][3] ), .A2(n674), .ZN(n670) );
  OAI21_X1 U53 ( .B1(n409), .B2(n674), .A(n669), .ZN(n521) );
  NAND2_X1 U54 ( .A1(\mem[2][4] ), .A2(n674), .ZN(n669) );
  OAI21_X1 U55 ( .B1(n408), .B2(n674), .A(n668), .ZN(n520) );
  NAND2_X1 U56 ( .A1(\mem[2][5] ), .A2(n674), .ZN(n668) );
  OAI21_X1 U57 ( .B1(n407), .B2(n674), .A(n667), .ZN(n519) );
  NAND2_X1 U58 ( .A1(\mem[2][6] ), .A2(n674), .ZN(n667) );
  OAI21_X1 U59 ( .B1(n406), .B2(n674), .A(n666), .ZN(n518) );
  NAND2_X1 U60 ( .A1(\mem[2][7] ), .A2(n674), .ZN(n666) );
  OAI21_X1 U61 ( .B1(n413), .B2(n664), .A(n663), .ZN(n517) );
  NAND2_X1 U62 ( .A1(\mem[3][0] ), .A2(n664), .ZN(n663) );
  OAI21_X1 U63 ( .B1(n412), .B2(n664), .A(n662), .ZN(n516) );
  NAND2_X1 U64 ( .A1(\mem[3][1] ), .A2(n664), .ZN(n662) );
  OAI21_X1 U65 ( .B1(n411), .B2(n664), .A(n661), .ZN(n515) );
  NAND2_X1 U66 ( .A1(\mem[3][2] ), .A2(n664), .ZN(n661) );
  OAI21_X1 U67 ( .B1(n410), .B2(n664), .A(n660), .ZN(n514) );
  NAND2_X1 U68 ( .A1(\mem[3][3] ), .A2(n664), .ZN(n660) );
  OAI21_X1 U69 ( .B1(n409), .B2(n664), .A(n659), .ZN(n513) );
  NAND2_X1 U70 ( .A1(\mem[3][4] ), .A2(n664), .ZN(n659) );
  OAI21_X1 U71 ( .B1(n408), .B2(n664), .A(n658), .ZN(n512) );
  NAND2_X1 U72 ( .A1(\mem[3][5] ), .A2(n664), .ZN(n658) );
  OAI21_X1 U73 ( .B1(n407), .B2(n664), .A(n657), .ZN(n511) );
  NAND2_X1 U74 ( .A1(\mem[3][6] ), .A2(n664), .ZN(n657) );
  OAI21_X1 U75 ( .B1(n406), .B2(n664), .A(n656), .ZN(n510) );
  NAND2_X1 U76 ( .A1(\mem[3][7] ), .A2(n664), .ZN(n656) );
  NOR2_X1 U77 ( .A1(n405), .A2(N13), .ZN(n626) );
  INV_X1 U78 ( .A(wr_en), .ZN(n405) );
  OAI21_X1 U79 ( .B1(n413), .B2(n684), .A(n683), .ZN(n533) );
  NAND2_X1 U80 ( .A1(\mem[1][0] ), .A2(n684), .ZN(n683) );
  OAI21_X1 U81 ( .B1(n412), .B2(n684), .A(n682), .ZN(n532) );
  NAND2_X1 U82 ( .A1(\mem[1][1] ), .A2(n684), .ZN(n682) );
  OAI21_X1 U83 ( .B1(n411), .B2(n684), .A(n681), .ZN(n531) );
  NAND2_X1 U84 ( .A1(\mem[1][2] ), .A2(n684), .ZN(n681) );
  OAI21_X1 U85 ( .B1(n410), .B2(n684), .A(n680), .ZN(n530) );
  NAND2_X1 U86 ( .A1(\mem[1][3] ), .A2(n684), .ZN(n680) );
  OAI21_X1 U87 ( .B1(n409), .B2(n684), .A(n679), .ZN(n529) );
  NAND2_X1 U88 ( .A1(\mem[1][4] ), .A2(n684), .ZN(n679) );
  OAI21_X1 U89 ( .B1(n408), .B2(n684), .A(n678), .ZN(n528) );
  NAND2_X1 U90 ( .A1(\mem[1][5] ), .A2(n684), .ZN(n678) );
  OAI21_X1 U91 ( .B1(n407), .B2(n684), .A(n677), .ZN(n527) );
  NAND2_X1 U92 ( .A1(\mem[1][6] ), .A2(n684), .ZN(n677) );
  OAI21_X1 U93 ( .B1(n406), .B2(n684), .A(n676), .ZN(n526) );
  NAND2_X1 U94 ( .A1(\mem[1][7] ), .A2(n684), .ZN(n676) );
  OAI21_X1 U95 ( .B1(n413), .B2(n655), .A(n654), .ZN(n509) );
  NAND2_X1 U96 ( .A1(\mem[4][0] ), .A2(n655), .ZN(n654) );
  OAI21_X1 U97 ( .B1(n412), .B2(n655), .A(n653), .ZN(n508) );
  NAND2_X1 U98 ( .A1(\mem[4][1] ), .A2(n655), .ZN(n653) );
  OAI21_X1 U99 ( .B1(n411), .B2(n655), .A(n652), .ZN(n507) );
  NAND2_X1 U100 ( .A1(\mem[4][2] ), .A2(n655), .ZN(n652) );
  OAI21_X1 U101 ( .B1(n410), .B2(n655), .A(n651), .ZN(n506) );
  NAND2_X1 U102 ( .A1(\mem[4][3] ), .A2(n655), .ZN(n651) );
  OAI21_X1 U103 ( .B1(n409), .B2(n655), .A(n650), .ZN(n505) );
  NAND2_X1 U104 ( .A1(\mem[4][4] ), .A2(n655), .ZN(n650) );
  OAI21_X1 U105 ( .B1(n408), .B2(n655), .A(n649), .ZN(n504) );
  NAND2_X1 U106 ( .A1(\mem[4][5] ), .A2(n655), .ZN(n649) );
  OAI21_X1 U107 ( .B1(n407), .B2(n655), .A(n648), .ZN(n503) );
  NAND2_X1 U108 ( .A1(\mem[4][6] ), .A2(n655), .ZN(n648) );
  OAI21_X1 U109 ( .B1(n406), .B2(n655), .A(n647), .ZN(n502) );
  NAND2_X1 U110 ( .A1(\mem[4][7] ), .A2(n655), .ZN(n647) );
  OAI21_X1 U111 ( .B1(n413), .B2(n645), .A(n644), .ZN(n501) );
  NAND2_X1 U112 ( .A1(\mem[5][0] ), .A2(n645), .ZN(n644) );
  OAI21_X1 U113 ( .B1(n412), .B2(n645), .A(n643), .ZN(n500) );
  NAND2_X1 U114 ( .A1(\mem[5][1] ), .A2(n645), .ZN(n643) );
  OAI21_X1 U115 ( .B1(n411), .B2(n645), .A(n642), .ZN(n499) );
  NAND2_X1 U116 ( .A1(\mem[5][2] ), .A2(n645), .ZN(n642) );
  OAI21_X1 U117 ( .B1(n410), .B2(n645), .A(n641), .ZN(n498) );
  NAND2_X1 U118 ( .A1(\mem[5][3] ), .A2(n645), .ZN(n641) );
  OAI21_X1 U119 ( .B1(n409), .B2(n645), .A(n640), .ZN(n497) );
  NAND2_X1 U120 ( .A1(\mem[5][4] ), .A2(n645), .ZN(n640) );
  OAI21_X1 U121 ( .B1(n408), .B2(n645), .A(n639), .ZN(n496) );
  NAND2_X1 U122 ( .A1(\mem[5][5] ), .A2(n645), .ZN(n639) );
  OAI21_X1 U123 ( .B1(n407), .B2(n645), .A(n638), .ZN(n495) );
  NAND2_X1 U124 ( .A1(\mem[5][6] ), .A2(n645), .ZN(n638) );
  OAI21_X1 U125 ( .B1(n406), .B2(n645), .A(n637), .ZN(n494) );
  NAND2_X1 U126 ( .A1(\mem[5][7] ), .A2(n645), .ZN(n637) );
  OAI21_X1 U127 ( .B1(n413), .B2(n636), .A(n635), .ZN(n493) );
  NAND2_X1 U128 ( .A1(\mem[6][0] ), .A2(n636), .ZN(n635) );
  OAI21_X1 U129 ( .B1(n412), .B2(n636), .A(n634), .ZN(n492) );
  NAND2_X1 U130 ( .A1(\mem[6][1] ), .A2(n636), .ZN(n634) );
  OAI21_X1 U131 ( .B1(n411), .B2(n636), .A(n633), .ZN(n491) );
  NAND2_X1 U132 ( .A1(\mem[6][2] ), .A2(n636), .ZN(n633) );
  OAI21_X1 U133 ( .B1(n410), .B2(n636), .A(n632), .ZN(n490) );
  NAND2_X1 U134 ( .A1(\mem[6][3] ), .A2(n636), .ZN(n632) );
  OAI21_X1 U135 ( .B1(n409), .B2(n636), .A(n631), .ZN(n489) );
  NAND2_X1 U136 ( .A1(\mem[6][4] ), .A2(n636), .ZN(n631) );
  OAI21_X1 U137 ( .B1(n408), .B2(n636), .A(n630), .ZN(n488) );
  NAND2_X1 U138 ( .A1(\mem[6][5] ), .A2(n636), .ZN(n630) );
  OAI21_X1 U139 ( .B1(n407), .B2(n636), .A(n629), .ZN(n487) );
  NAND2_X1 U140 ( .A1(\mem[6][6] ), .A2(n636), .ZN(n629) );
  OAI21_X1 U141 ( .B1(n406), .B2(n636), .A(n628), .ZN(n486) );
  NAND2_X1 U142 ( .A1(\mem[6][7] ), .A2(n636), .ZN(n628) );
  OAI21_X1 U143 ( .B1(n413), .B2(n625), .A(n624), .ZN(n485) );
  NAND2_X1 U144 ( .A1(\mem[7][0] ), .A2(n625), .ZN(n624) );
  OAI21_X1 U145 ( .B1(n412), .B2(n625), .A(n623), .ZN(n484) );
  NAND2_X1 U146 ( .A1(\mem[7][1] ), .A2(n625), .ZN(n623) );
  OAI21_X1 U147 ( .B1(n411), .B2(n625), .A(n622), .ZN(n483) );
  NAND2_X1 U148 ( .A1(\mem[7][2] ), .A2(n625), .ZN(n622) );
  OAI21_X1 U149 ( .B1(n410), .B2(n625), .A(n621), .ZN(n482) );
  NAND2_X1 U150 ( .A1(\mem[7][3] ), .A2(n625), .ZN(n621) );
  OAI21_X1 U151 ( .B1(n409), .B2(n625), .A(n620), .ZN(n481) );
  NAND2_X1 U152 ( .A1(\mem[7][4] ), .A2(n625), .ZN(n620) );
  OAI21_X1 U153 ( .B1(n408), .B2(n625), .A(n619), .ZN(n480) );
  NAND2_X1 U154 ( .A1(\mem[7][5] ), .A2(n625), .ZN(n619) );
  OAI21_X1 U155 ( .B1(n407), .B2(n625), .A(n618), .ZN(n479) );
  NAND2_X1 U156 ( .A1(\mem[7][6] ), .A2(n625), .ZN(n618) );
  OAI21_X1 U157 ( .B1(n406), .B2(n625), .A(n617), .ZN(n478) );
  NAND2_X1 U158 ( .A1(\mem[7][7] ), .A2(n625), .ZN(n617) );
  OAI21_X1 U159 ( .B1(n413), .B2(n616), .A(n615), .ZN(n477) );
  NAND2_X1 U160 ( .A1(\mem[8][0] ), .A2(n616), .ZN(n615) );
  OAI21_X1 U161 ( .B1(n412), .B2(n616), .A(n614), .ZN(n476) );
  NAND2_X1 U162 ( .A1(\mem[8][1] ), .A2(n616), .ZN(n614) );
  OAI21_X1 U163 ( .B1(n411), .B2(n616), .A(n613), .ZN(n475) );
  NAND2_X1 U164 ( .A1(\mem[8][2] ), .A2(n616), .ZN(n613) );
  OAI21_X1 U165 ( .B1(n410), .B2(n616), .A(n612), .ZN(n474) );
  NAND2_X1 U166 ( .A1(\mem[8][3] ), .A2(n616), .ZN(n612) );
  OAI21_X1 U167 ( .B1(n409), .B2(n616), .A(n611), .ZN(n473) );
  NAND2_X1 U168 ( .A1(\mem[8][4] ), .A2(n616), .ZN(n611) );
  OAI21_X1 U169 ( .B1(n408), .B2(n616), .A(n610), .ZN(n472) );
  NAND2_X1 U170 ( .A1(\mem[8][5] ), .A2(n616), .ZN(n610) );
  OAI21_X1 U171 ( .B1(n407), .B2(n616), .A(n609), .ZN(n471) );
  NAND2_X1 U172 ( .A1(\mem[8][6] ), .A2(n616), .ZN(n609) );
  OAI21_X1 U173 ( .B1(n406), .B2(n616), .A(n608), .ZN(n470) );
  NAND2_X1 U174 ( .A1(\mem[8][7] ), .A2(n616), .ZN(n608) );
  OAI21_X1 U175 ( .B1(n413), .B2(n606), .A(n605), .ZN(n469) );
  NAND2_X1 U176 ( .A1(\mem[9][0] ), .A2(n606), .ZN(n605) );
  OAI21_X1 U177 ( .B1(n412), .B2(n606), .A(n604), .ZN(n468) );
  NAND2_X1 U178 ( .A1(\mem[9][1] ), .A2(n606), .ZN(n604) );
  OAI21_X1 U179 ( .B1(n411), .B2(n606), .A(n603), .ZN(n467) );
  NAND2_X1 U180 ( .A1(\mem[9][2] ), .A2(n606), .ZN(n603) );
  OAI21_X1 U181 ( .B1(n410), .B2(n606), .A(n602), .ZN(n466) );
  NAND2_X1 U182 ( .A1(\mem[9][3] ), .A2(n606), .ZN(n602) );
  OAI21_X1 U183 ( .B1(n409), .B2(n606), .A(n601), .ZN(n465) );
  NAND2_X1 U184 ( .A1(\mem[9][4] ), .A2(n606), .ZN(n601) );
  OAI21_X1 U185 ( .B1(n408), .B2(n606), .A(n600), .ZN(n464) );
  NAND2_X1 U186 ( .A1(\mem[9][5] ), .A2(n606), .ZN(n600) );
  OAI21_X1 U187 ( .B1(n407), .B2(n606), .A(n599), .ZN(n463) );
  NAND2_X1 U188 ( .A1(\mem[9][6] ), .A2(n606), .ZN(n599) );
  OAI21_X1 U189 ( .B1(n406), .B2(n606), .A(n598), .ZN(n462) );
  NAND2_X1 U190 ( .A1(\mem[9][7] ), .A2(n606), .ZN(n598) );
  OAI21_X1 U191 ( .B1(n413), .B2(n596), .A(n595), .ZN(n461) );
  NAND2_X1 U192 ( .A1(\mem[10][0] ), .A2(n596), .ZN(n595) );
  OAI21_X1 U193 ( .B1(n412), .B2(n596), .A(n594), .ZN(n460) );
  NAND2_X1 U194 ( .A1(\mem[10][1] ), .A2(n596), .ZN(n594) );
  OAI21_X1 U195 ( .B1(n411), .B2(n596), .A(n593), .ZN(n459) );
  NAND2_X1 U196 ( .A1(\mem[10][2] ), .A2(n596), .ZN(n593) );
  OAI21_X1 U197 ( .B1(n410), .B2(n596), .A(n592), .ZN(n458) );
  NAND2_X1 U198 ( .A1(\mem[10][3] ), .A2(n596), .ZN(n592) );
  OAI21_X1 U199 ( .B1(n409), .B2(n596), .A(n591), .ZN(n457) );
  NAND2_X1 U200 ( .A1(\mem[10][4] ), .A2(n596), .ZN(n591) );
  OAI21_X1 U201 ( .B1(n408), .B2(n596), .A(n590), .ZN(n456) );
  NAND2_X1 U202 ( .A1(\mem[10][5] ), .A2(n596), .ZN(n590) );
  OAI21_X1 U203 ( .B1(n407), .B2(n596), .A(n589), .ZN(n455) );
  NAND2_X1 U204 ( .A1(\mem[10][6] ), .A2(n596), .ZN(n589) );
  OAI21_X1 U205 ( .B1(n406), .B2(n596), .A(n588), .ZN(n454) );
  NAND2_X1 U206 ( .A1(\mem[10][7] ), .A2(n596), .ZN(n588) );
  OAI21_X1 U207 ( .B1(n413), .B2(n587), .A(n586), .ZN(n453) );
  NAND2_X1 U208 ( .A1(\mem[11][0] ), .A2(n587), .ZN(n586) );
  OAI21_X1 U209 ( .B1(n412), .B2(n587), .A(n585), .ZN(n452) );
  NAND2_X1 U210 ( .A1(\mem[11][1] ), .A2(n587), .ZN(n585) );
  OAI21_X1 U211 ( .B1(n411), .B2(n587), .A(n584), .ZN(n451) );
  NAND2_X1 U212 ( .A1(\mem[11][2] ), .A2(n587), .ZN(n584) );
  OAI21_X1 U213 ( .B1(n410), .B2(n587), .A(n583), .ZN(n450) );
  NAND2_X1 U214 ( .A1(\mem[11][3] ), .A2(n587), .ZN(n583) );
  OAI21_X1 U215 ( .B1(n409), .B2(n587), .A(n582), .ZN(n449) );
  NAND2_X1 U216 ( .A1(\mem[11][4] ), .A2(n587), .ZN(n582) );
  OAI21_X1 U217 ( .B1(n408), .B2(n587), .A(n581), .ZN(n448) );
  NAND2_X1 U218 ( .A1(\mem[11][5] ), .A2(n587), .ZN(n581) );
  OAI21_X1 U219 ( .B1(n407), .B2(n587), .A(n580), .ZN(n447) );
  NAND2_X1 U220 ( .A1(\mem[11][6] ), .A2(n587), .ZN(n580) );
  OAI21_X1 U221 ( .B1(n406), .B2(n587), .A(n579), .ZN(n446) );
  NAND2_X1 U222 ( .A1(\mem[11][7] ), .A2(n587), .ZN(n579) );
  OAI21_X1 U223 ( .B1(n413), .B2(n578), .A(n577), .ZN(n445) );
  NAND2_X1 U224 ( .A1(\mem[12][0] ), .A2(n578), .ZN(n577) );
  OAI21_X1 U225 ( .B1(n412), .B2(n578), .A(n576), .ZN(n444) );
  NAND2_X1 U226 ( .A1(\mem[12][1] ), .A2(n578), .ZN(n576) );
  OAI21_X1 U227 ( .B1(n411), .B2(n578), .A(n575), .ZN(n443) );
  NAND2_X1 U228 ( .A1(\mem[12][2] ), .A2(n578), .ZN(n575) );
  OAI21_X1 U229 ( .B1(n410), .B2(n578), .A(n574), .ZN(n442) );
  NAND2_X1 U230 ( .A1(\mem[12][3] ), .A2(n578), .ZN(n574) );
  OAI21_X1 U231 ( .B1(n409), .B2(n578), .A(n573), .ZN(n441) );
  NAND2_X1 U232 ( .A1(\mem[12][4] ), .A2(n578), .ZN(n573) );
  OAI21_X1 U233 ( .B1(n408), .B2(n578), .A(n572), .ZN(n440) );
  NAND2_X1 U234 ( .A1(\mem[12][5] ), .A2(n578), .ZN(n572) );
  OAI21_X1 U235 ( .B1(n407), .B2(n578), .A(n571), .ZN(n439) );
  NAND2_X1 U236 ( .A1(\mem[12][6] ), .A2(n578), .ZN(n571) );
  OAI21_X1 U237 ( .B1(n406), .B2(n578), .A(n570), .ZN(n438) );
  NAND2_X1 U238 ( .A1(\mem[12][7] ), .A2(n578), .ZN(n570) );
  OAI21_X1 U239 ( .B1(n413), .B2(n569), .A(n568), .ZN(n437) );
  NAND2_X1 U240 ( .A1(\mem[13][0] ), .A2(n569), .ZN(n568) );
  OAI21_X1 U241 ( .B1(n412), .B2(n569), .A(n567), .ZN(n436) );
  NAND2_X1 U242 ( .A1(\mem[13][1] ), .A2(n569), .ZN(n567) );
  OAI21_X1 U243 ( .B1(n411), .B2(n569), .A(n566), .ZN(n435) );
  NAND2_X1 U244 ( .A1(\mem[13][2] ), .A2(n569), .ZN(n566) );
  OAI21_X1 U245 ( .B1(n410), .B2(n569), .A(n565), .ZN(n434) );
  NAND2_X1 U246 ( .A1(\mem[13][3] ), .A2(n569), .ZN(n565) );
  OAI21_X1 U247 ( .B1(n409), .B2(n569), .A(n564), .ZN(n433) );
  NAND2_X1 U248 ( .A1(\mem[13][4] ), .A2(n569), .ZN(n564) );
  OAI21_X1 U249 ( .B1(n408), .B2(n569), .A(n563), .ZN(n432) );
  NAND2_X1 U250 ( .A1(\mem[13][5] ), .A2(n569), .ZN(n563) );
  OAI21_X1 U251 ( .B1(n407), .B2(n569), .A(n562), .ZN(n431) );
  NAND2_X1 U252 ( .A1(\mem[13][6] ), .A2(n569), .ZN(n562) );
  OAI21_X1 U253 ( .B1(n406), .B2(n569), .A(n561), .ZN(n430) );
  NAND2_X1 U254 ( .A1(\mem[13][7] ), .A2(n569), .ZN(n561) );
  OAI21_X1 U255 ( .B1(n413), .B2(n560), .A(n559), .ZN(n429) );
  NAND2_X1 U256 ( .A1(\mem[14][0] ), .A2(n560), .ZN(n559) );
  OAI21_X1 U257 ( .B1(n412), .B2(n560), .A(n558), .ZN(n428) );
  NAND2_X1 U258 ( .A1(\mem[14][1] ), .A2(n560), .ZN(n558) );
  OAI21_X1 U259 ( .B1(n411), .B2(n560), .A(n557), .ZN(n427) );
  NAND2_X1 U260 ( .A1(\mem[14][2] ), .A2(n560), .ZN(n557) );
  OAI21_X1 U261 ( .B1(n410), .B2(n560), .A(n556), .ZN(n426) );
  NAND2_X1 U262 ( .A1(\mem[14][3] ), .A2(n560), .ZN(n556) );
  OAI21_X1 U263 ( .B1(n409), .B2(n560), .A(n555), .ZN(n425) );
  NAND2_X1 U264 ( .A1(\mem[14][4] ), .A2(n560), .ZN(n555) );
  OAI21_X1 U265 ( .B1(n408), .B2(n560), .A(n554), .ZN(n424) );
  NAND2_X1 U266 ( .A1(\mem[14][5] ), .A2(n560), .ZN(n554) );
  OAI21_X1 U267 ( .B1(n407), .B2(n560), .A(n553), .ZN(n423) );
  NAND2_X1 U268 ( .A1(\mem[14][6] ), .A2(n560), .ZN(n553) );
  OAI21_X1 U269 ( .B1(n406), .B2(n560), .A(n552), .ZN(n422) );
  NAND2_X1 U270 ( .A1(\mem[14][7] ), .A2(n560), .ZN(n552) );
  OAI21_X1 U271 ( .B1(n413), .B2(n550), .A(n549), .ZN(n421) );
  NAND2_X1 U272 ( .A1(\mem[15][0] ), .A2(n550), .ZN(n549) );
  OAI21_X1 U273 ( .B1(n412), .B2(n550), .A(n548), .ZN(n420) );
  NAND2_X1 U274 ( .A1(\mem[15][1] ), .A2(n550), .ZN(n548) );
  OAI21_X1 U275 ( .B1(n411), .B2(n550), .A(n547), .ZN(n419) );
  NAND2_X1 U276 ( .A1(\mem[15][2] ), .A2(n550), .ZN(n547) );
  OAI21_X1 U277 ( .B1(n410), .B2(n550), .A(n546), .ZN(n418) );
  NAND2_X1 U278 ( .A1(\mem[15][3] ), .A2(n550), .ZN(n546) );
  OAI21_X1 U279 ( .B1(n409), .B2(n550), .A(n545), .ZN(n417) );
  NAND2_X1 U280 ( .A1(\mem[15][4] ), .A2(n550), .ZN(n545) );
  OAI21_X1 U281 ( .B1(n408), .B2(n550), .A(n544), .ZN(n416) );
  NAND2_X1 U282 ( .A1(\mem[15][5] ), .A2(n550), .ZN(n544) );
  OAI21_X1 U283 ( .B1(n407), .B2(n550), .A(n543), .ZN(n415) );
  NAND2_X1 U284 ( .A1(\mem[15][6] ), .A2(n550), .ZN(n543) );
  OAI21_X1 U285 ( .B1(n406), .B2(n550), .A(n542), .ZN(n414) );
  NAND2_X1 U286 ( .A1(\mem[15][7] ), .A2(n550), .ZN(n542) );
  AND2_X1 U287 ( .A1(N13), .A2(wr_en), .ZN(n551) );
  NOR2_X1 U288 ( .A1(N11), .A2(N12), .ZN(n686) );
  NOR2_X1 U289 ( .A1(n404), .A2(N12), .ZN(n665) );
  AND2_X1 U290 ( .A1(N12), .A2(n404), .ZN(n646) );
  AND2_X1 U291 ( .A1(N12), .A2(N11), .ZN(n627) );
  INV_X1 U292 ( .A(data_in[0]), .ZN(n413) );
  INV_X1 U293 ( .A(data_in[1]), .ZN(n412) );
  INV_X1 U294 ( .A(data_in[2]), .ZN(n411) );
  INV_X1 U295 ( .A(data_in[3]), .ZN(n410) );
  INV_X1 U296 ( .A(data_in[4]), .ZN(n409) );
  INV_X1 U297 ( .A(data_in[5]), .ZN(n408) );
  INV_X1 U298 ( .A(data_in[6]), .ZN(n407) );
  INV_X1 U299 ( .A(data_in[7]), .ZN(n406) );
  MUX2_X1 U300 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(N10), .Z(n5) );
  MUX2_X1 U301 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n401), .Z(n6) );
  MUX2_X1 U302 ( .A(n6), .B(n5), .S(n399), .Z(n7) );
  MUX2_X1 U303 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n400), .Z(n8) );
  MUX2_X1 U304 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n401), .Z(n9) );
  MUX2_X1 U305 ( .A(n9), .B(n8), .S(N11), .Z(n10) );
  MUX2_X1 U306 ( .A(n10), .B(n7), .S(N12), .Z(n11) );
  MUX2_X1 U307 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(N10), .Z(n294) );
  MUX2_X1 U308 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(N10), .Z(n295) );
  MUX2_X1 U309 ( .A(n295), .B(n294), .S(N11), .Z(n296) );
  MUX2_X1 U310 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(N10), .Z(n297) );
  MUX2_X1 U311 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n298) );
  MUX2_X1 U312 ( .A(n298), .B(n297), .S(N11), .Z(n299) );
  MUX2_X1 U313 ( .A(n299), .B(n296), .S(N12), .Z(n300) );
  MUX2_X1 U314 ( .A(n300), .B(n11), .S(N13), .Z(N21) );
  MUX2_X1 U315 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n401), .Z(n301) );
  MUX2_X1 U316 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(N10), .Z(n302) );
  MUX2_X1 U317 ( .A(n302), .B(n301), .S(N11), .Z(n303) );
  MUX2_X1 U318 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n402), .Z(n304) );
  MUX2_X1 U319 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(N10), .Z(n305) );
  MUX2_X1 U320 ( .A(n305), .B(n304), .S(N11), .Z(n306) );
  MUX2_X1 U321 ( .A(n306), .B(n303), .S(N12), .Z(n307) );
  MUX2_X1 U322 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(N10), .Z(n308) );
  MUX2_X1 U323 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(N10), .Z(n309) );
  MUX2_X1 U324 ( .A(n309), .B(n308), .S(N11), .Z(n310) );
  MUX2_X1 U325 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(N10), .Z(n311) );
  MUX2_X1 U326 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(N10), .Z(n312) );
  MUX2_X1 U327 ( .A(n312), .B(n311), .S(N11), .Z(n313) );
  MUX2_X1 U328 ( .A(n313), .B(n310), .S(N12), .Z(n314) );
  MUX2_X1 U329 ( .A(n314), .B(n307), .S(N13), .Z(N20) );
  MUX2_X1 U330 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(N10), .Z(n315) );
  MUX2_X1 U331 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n402), .Z(n316) );
  MUX2_X1 U332 ( .A(n316), .B(n315), .S(n399), .Z(n317) );
  MUX2_X1 U333 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n400), .Z(n318) );
  MUX2_X1 U334 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(N10), .Z(n319) );
  MUX2_X1 U335 ( .A(n319), .B(n318), .S(n399), .Z(n320) );
  MUX2_X1 U336 ( .A(n320), .B(n317), .S(N12), .Z(n321) );
  MUX2_X1 U337 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n402), .Z(n322) );
  MUX2_X1 U338 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n402), .Z(n323) );
  MUX2_X1 U339 ( .A(n323), .B(n322), .S(n399), .Z(n324) );
  MUX2_X1 U340 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n400), .Z(n325) );
  MUX2_X1 U341 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(N10), .Z(n326) );
  MUX2_X1 U342 ( .A(n326), .B(n325), .S(n399), .Z(n327) );
  MUX2_X1 U343 ( .A(n327), .B(n324), .S(N12), .Z(n328) );
  MUX2_X1 U344 ( .A(n328), .B(n321), .S(N13), .Z(N19) );
  MUX2_X1 U345 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(N10), .Z(n329) );
  MUX2_X1 U346 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n400), .Z(n330) );
  MUX2_X1 U347 ( .A(n330), .B(n329), .S(n399), .Z(n331) );
  MUX2_X1 U348 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n401), .Z(n332) );
  MUX2_X1 U349 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n333) );
  MUX2_X1 U350 ( .A(n333), .B(n332), .S(n399), .Z(n334) );
  MUX2_X1 U351 ( .A(n334), .B(n331), .S(N12), .Z(n335) );
  MUX2_X1 U352 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n400), .Z(n336) );
  MUX2_X1 U353 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n400), .Z(n337) );
  MUX2_X1 U354 ( .A(n337), .B(n336), .S(n399), .Z(n338) );
  MUX2_X1 U355 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n400), .Z(n339) );
  MUX2_X1 U356 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n400), .Z(n340) );
  MUX2_X1 U357 ( .A(n340), .B(n339), .S(n399), .Z(n341) );
  MUX2_X1 U358 ( .A(n341), .B(n338), .S(N12), .Z(n342) );
  MUX2_X1 U359 ( .A(n342), .B(n335), .S(N13), .Z(N18) );
  MUX2_X1 U360 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n400), .Z(n343) );
  MUX2_X1 U361 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n400), .Z(n344) );
  MUX2_X1 U362 ( .A(n344), .B(n343), .S(n399), .Z(n345) );
  MUX2_X1 U363 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n400), .Z(n346) );
  MUX2_X1 U364 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n400), .Z(n347) );
  MUX2_X1 U365 ( .A(n347), .B(n346), .S(n399), .Z(n348) );
  MUX2_X1 U366 ( .A(n348), .B(n345), .S(N12), .Z(n349) );
  MUX2_X1 U367 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n400), .Z(n350) );
  MUX2_X1 U368 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n400), .Z(n351) );
  MUX2_X1 U369 ( .A(n351), .B(n350), .S(n399), .Z(n352) );
  MUX2_X1 U370 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n400), .Z(n353) );
  MUX2_X1 U371 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n400), .Z(n354) );
  MUX2_X1 U372 ( .A(n354), .B(n353), .S(n399), .Z(n355) );
  MUX2_X1 U373 ( .A(n355), .B(n352), .S(N12), .Z(n356) );
  MUX2_X1 U374 ( .A(n356), .B(n349), .S(N13), .Z(N17) );
  MUX2_X1 U375 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n401), .Z(n357) );
  MUX2_X1 U376 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n401), .Z(n358) );
  MUX2_X1 U377 ( .A(n358), .B(n357), .S(N11), .Z(n359) );
  MUX2_X1 U378 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n401), .Z(n360) );
  MUX2_X1 U379 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n401), .Z(n361) );
  MUX2_X1 U380 ( .A(n361), .B(n360), .S(N11), .Z(n362) );
  MUX2_X1 U381 ( .A(n362), .B(n359), .S(N12), .Z(n363) );
  MUX2_X1 U382 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n401), .Z(n364) );
  MUX2_X1 U383 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n401), .Z(n365) );
  MUX2_X1 U384 ( .A(n365), .B(n364), .S(N11), .Z(n366) );
  MUX2_X1 U385 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n401), .Z(n367) );
  MUX2_X1 U386 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n401), .Z(n368) );
  MUX2_X1 U387 ( .A(n368), .B(n367), .S(N11), .Z(n369) );
  MUX2_X1 U388 ( .A(n369), .B(n366), .S(N12), .Z(n370) );
  MUX2_X1 U389 ( .A(n370), .B(n363), .S(N13), .Z(N16) );
  MUX2_X1 U390 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n401), .Z(n371) );
  MUX2_X1 U391 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n401), .Z(n372) );
  MUX2_X1 U392 ( .A(n372), .B(n371), .S(N11), .Z(n373) );
  MUX2_X1 U393 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n401), .Z(n374) );
  MUX2_X1 U394 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n401), .Z(n375) );
  MUX2_X1 U395 ( .A(n375), .B(n374), .S(N11), .Z(n376) );
  MUX2_X1 U396 ( .A(n376), .B(n373), .S(N12), .Z(n377) );
  MUX2_X1 U397 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n402), .Z(n378) );
  MUX2_X1 U398 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n402), .Z(n379) );
  MUX2_X1 U399 ( .A(n379), .B(n378), .S(N11), .Z(n380) );
  MUX2_X1 U400 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n402), .Z(n381) );
  MUX2_X1 U401 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n402), .Z(n382) );
  MUX2_X1 U402 ( .A(n382), .B(n381), .S(N11), .Z(n383) );
  MUX2_X1 U403 ( .A(n383), .B(n380), .S(N12), .Z(n384) );
  MUX2_X1 U404 ( .A(n384), .B(n377), .S(N13), .Z(N15) );
  MUX2_X1 U405 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n402), .Z(n385) );
  MUX2_X1 U406 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n402), .Z(n386) );
  MUX2_X1 U407 ( .A(n386), .B(n385), .S(N11), .Z(n387) );
  MUX2_X1 U408 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n402), .Z(n388) );
  MUX2_X1 U409 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n402), .Z(n389) );
  MUX2_X1 U410 ( .A(n389), .B(n388), .S(N11), .Z(n390) );
  MUX2_X1 U411 ( .A(n390), .B(n387), .S(N12), .Z(n391) );
  MUX2_X1 U412 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n402), .Z(n392) );
  MUX2_X1 U413 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n402), .Z(n393) );
  MUX2_X1 U414 ( .A(n393), .B(n392), .S(N11), .Z(n394) );
  MUX2_X1 U415 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n402), .Z(n395) );
  MUX2_X1 U416 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n402), .Z(n396) );
  MUX2_X1 U417 ( .A(n396), .B(n395), .S(n399), .Z(n397) );
  MUX2_X1 U418 ( .A(n397), .B(n394), .S(N12), .Z(n398) );
  MUX2_X1 U419 ( .A(n398), .B(n391), .S(N13), .Z(N14) );
  INV_X1 U420 ( .A(N10), .ZN(n403) );
  INV_X1 U421 ( .A(N11), .ZN(n404) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_5 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, N19, N20, N21, n1, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n413), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n414), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n415), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n416), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n417), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n418), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n419), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n420), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n421), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n422), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n423), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n424), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n425), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n426), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n427), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n428), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n429), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n430), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n431), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n432), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n433), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n434), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n435), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n436), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n437), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n438), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n439), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n440), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n441), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n442), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n443), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n444), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n445), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n446), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n447), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n448), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n449), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n450), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n451), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n452), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n453), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n454), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n455), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n456), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n457), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n458), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n459), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n460), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n461), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n462), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n463), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n464), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n465), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n466), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n467), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n468), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n469), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n470), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n471), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n472), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n473), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n474), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n475), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n476), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n477), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n478), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n479), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n480), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n481), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n482), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n483), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n484), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n485), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n486), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n487), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n488), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n489), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n490), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n491), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n492), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n493), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n494), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n495), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n496), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n497), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n498), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n499), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n500), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n501), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n502), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n503), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n504), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n505), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n506), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n507), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n508), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n509), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n510), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n511), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n512), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n513), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n514), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n515), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n516), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n517), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n518), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n519), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n520), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n521), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n522), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n523), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n524), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n525), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n526), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n527), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n528), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n529), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n530), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n531), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n532), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n533), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n534), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n535), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n536), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n537), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n538), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n539), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n540), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N20), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .QN(n1) );
  DFF_X1 \data_out_reg[5]  ( .D(N16), .CK(clk), .Q(data_out[5]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(N10), .Z(n398) );
  BUF_X1 U5 ( .A(N10), .Z(n399) );
  BUF_X1 U6 ( .A(N10), .Z(n400) );
  BUF_X1 U7 ( .A(N11), .Z(n397) );
  NAND2_X1 U8 ( .A1(n664), .A2(n684), .ZN(n673) );
  NAND2_X1 U9 ( .A1(n664), .A2(n674), .ZN(n663) );
  NAND2_X1 U10 ( .A1(n685), .A2(n684), .ZN(n694) );
  NAND2_X1 U11 ( .A1(n674), .A2(n685), .ZN(n683) );
  NAND2_X1 U12 ( .A1(n606), .A2(n685), .ZN(n615) );
  NAND2_X1 U13 ( .A1(n596), .A2(n685), .ZN(n605) );
  NAND2_X1 U14 ( .A1(n606), .A2(n664), .ZN(n595) );
  NAND2_X1 U15 ( .A1(n596), .A2(n664), .ZN(n586) );
  NAND2_X1 U16 ( .A1(n645), .A2(n684), .ZN(n654) );
  NAND2_X1 U17 ( .A1(n645), .A2(n674), .ZN(n644) );
  NAND2_X1 U18 ( .A1(n626), .A2(n684), .ZN(n635) );
  NAND2_X1 U19 ( .A1(n626), .A2(n674), .ZN(n624) );
  NAND2_X1 U20 ( .A1(n606), .A2(n645), .ZN(n577) );
  NAND2_X1 U21 ( .A1(n596), .A2(n645), .ZN(n568) );
  NAND2_X1 U22 ( .A1(n606), .A2(n626), .ZN(n559) );
  NAND2_X1 U23 ( .A1(n596), .A2(n626), .ZN(n549) );
  AND2_X1 U24 ( .A1(n550), .A2(N10), .ZN(n596) );
  AND2_X1 U25 ( .A1(n550), .A2(n402), .ZN(n606) );
  AND2_X1 U26 ( .A1(N10), .A2(n625), .ZN(n674) );
  AND2_X1 U27 ( .A1(n625), .A2(n402), .ZN(n684) );
  OAI21_X1 U28 ( .B1(n694), .B2(n412), .A(n693), .ZN(n540) );
  NAND2_X1 U29 ( .A1(\mem[0][0] ), .A2(n694), .ZN(n693) );
  OAI21_X1 U30 ( .B1(n694), .B2(n411), .A(n692), .ZN(n539) );
  NAND2_X1 U31 ( .A1(\mem[0][1] ), .A2(n694), .ZN(n692) );
  OAI21_X1 U32 ( .B1(n694), .B2(n410), .A(n691), .ZN(n538) );
  NAND2_X1 U33 ( .A1(\mem[0][2] ), .A2(n694), .ZN(n691) );
  OAI21_X1 U34 ( .B1(n694), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U35 ( .A1(\mem[0][3] ), .A2(n694), .ZN(n690) );
  OAI21_X1 U36 ( .B1(n694), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U37 ( .A1(\mem[0][4] ), .A2(n694), .ZN(n689) );
  OAI21_X1 U38 ( .B1(n694), .B2(n407), .A(n688), .ZN(n535) );
  NAND2_X1 U39 ( .A1(\mem[0][5] ), .A2(n694), .ZN(n688) );
  OAI21_X1 U40 ( .B1(n694), .B2(n406), .A(n687), .ZN(n534) );
  NAND2_X1 U41 ( .A1(\mem[0][6] ), .A2(n694), .ZN(n687) );
  OAI21_X1 U42 ( .B1(n694), .B2(n405), .A(n686), .ZN(n533) );
  NAND2_X1 U43 ( .A1(\mem[0][7] ), .A2(n694), .ZN(n686) );
  OAI21_X1 U44 ( .B1(n412), .B2(n673), .A(n672), .ZN(n524) );
  NAND2_X1 U45 ( .A1(\mem[2][0] ), .A2(n673), .ZN(n672) );
  OAI21_X1 U46 ( .B1(n411), .B2(n673), .A(n671), .ZN(n523) );
  NAND2_X1 U47 ( .A1(\mem[2][1] ), .A2(n673), .ZN(n671) );
  OAI21_X1 U48 ( .B1(n410), .B2(n673), .A(n670), .ZN(n522) );
  NAND2_X1 U49 ( .A1(\mem[2][2] ), .A2(n673), .ZN(n670) );
  OAI21_X1 U50 ( .B1(n409), .B2(n673), .A(n669), .ZN(n521) );
  NAND2_X1 U51 ( .A1(\mem[2][3] ), .A2(n673), .ZN(n669) );
  OAI21_X1 U52 ( .B1(n408), .B2(n673), .A(n668), .ZN(n520) );
  NAND2_X1 U53 ( .A1(\mem[2][4] ), .A2(n673), .ZN(n668) );
  OAI21_X1 U54 ( .B1(n407), .B2(n673), .A(n667), .ZN(n519) );
  NAND2_X1 U55 ( .A1(\mem[2][5] ), .A2(n673), .ZN(n667) );
  OAI21_X1 U56 ( .B1(n406), .B2(n673), .A(n666), .ZN(n518) );
  NAND2_X1 U57 ( .A1(\mem[2][6] ), .A2(n673), .ZN(n666) );
  OAI21_X1 U58 ( .B1(n405), .B2(n673), .A(n665), .ZN(n517) );
  NAND2_X1 U59 ( .A1(\mem[2][7] ), .A2(n673), .ZN(n665) );
  OAI21_X1 U60 ( .B1(n412), .B2(n663), .A(n662), .ZN(n516) );
  NAND2_X1 U61 ( .A1(\mem[3][0] ), .A2(n663), .ZN(n662) );
  OAI21_X1 U62 ( .B1(n411), .B2(n663), .A(n661), .ZN(n515) );
  NAND2_X1 U63 ( .A1(\mem[3][1] ), .A2(n663), .ZN(n661) );
  OAI21_X1 U64 ( .B1(n410), .B2(n663), .A(n660), .ZN(n514) );
  NAND2_X1 U65 ( .A1(\mem[3][2] ), .A2(n663), .ZN(n660) );
  OAI21_X1 U66 ( .B1(n409), .B2(n663), .A(n659), .ZN(n513) );
  NAND2_X1 U67 ( .A1(\mem[3][3] ), .A2(n663), .ZN(n659) );
  OAI21_X1 U68 ( .B1(n408), .B2(n663), .A(n658), .ZN(n512) );
  NAND2_X1 U69 ( .A1(\mem[3][4] ), .A2(n663), .ZN(n658) );
  OAI21_X1 U70 ( .B1(n407), .B2(n663), .A(n657), .ZN(n511) );
  NAND2_X1 U71 ( .A1(\mem[3][5] ), .A2(n663), .ZN(n657) );
  OAI21_X1 U72 ( .B1(n406), .B2(n663), .A(n656), .ZN(n510) );
  NAND2_X1 U73 ( .A1(\mem[3][6] ), .A2(n663), .ZN(n656) );
  OAI21_X1 U74 ( .B1(n405), .B2(n663), .A(n655), .ZN(n509) );
  NAND2_X1 U75 ( .A1(\mem[3][7] ), .A2(n663), .ZN(n655) );
  NOR2_X1 U76 ( .A1(n404), .A2(N13), .ZN(n625) );
  INV_X1 U77 ( .A(wr_en), .ZN(n404) );
  OAI21_X1 U78 ( .B1(n412), .B2(n683), .A(n682), .ZN(n532) );
  NAND2_X1 U79 ( .A1(\mem[1][0] ), .A2(n683), .ZN(n682) );
  OAI21_X1 U80 ( .B1(n411), .B2(n683), .A(n681), .ZN(n531) );
  NAND2_X1 U81 ( .A1(\mem[1][1] ), .A2(n683), .ZN(n681) );
  OAI21_X1 U82 ( .B1(n410), .B2(n683), .A(n680), .ZN(n530) );
  NAND2_X1 U83 ( .A1(\mem[1][2] ), .A2(n683), .ZN(n680) );
  OAI21_X1 U84 ( .B1(n409), .B2(n683), .A(n679), .ZN(n529) );
  NAND2_X1 U85 ( .A1(\mem[1][3] ), .A2(n683), .ZN(n679) );
  OAI21_X1 U86 ( .B1(n408), .B2(n683), .A(n678), .ZN(n528) );
  NAND2_X1 U87 ( .A1(\mem[1][4] ), .A2(n683), .ZN(n678) );
  OAI21_X1 U88 ( .B1(n407), .B2(n683), .A(n677), .ZN(n527) );
  NAND2_X1 U89 ( .A1(\mem[1][5] ), .A2(n683), .ZN(n677) );
  OAI21_X1 U90 ( .B1(n406), .B2(n683), .A(n676), .ZN(n526) );
  NAND2_X1 U91 ( .A1(\mem[1][6] ), .A2(n683), .ZN(n676) );
  OAI21_X1 U92 ( .B1(n405), .B2(n683), .A(n675), .ZN(n525) );
  NAND2_X1 U93 ( .A1(\mem[1][7] ), .A2(n683), .ZN(n675) );
  OAI21_X1 U94 ( .B1(n412), .B2(n654), .A(n653), .ZN(n508) );
  NAND2_X1 U95 ( .A1(\mem[4][0] ), .A2(n654), .ZN(n653) );
  OAI21_X1 U96 ( .B1(n411), .B2(n654), .A(n652), .ZN(n507) );
  NAND2_X1 U97 ( .A1(\mem[4][1] ), .A2(n654), .ZN(n652) );
  OAI21_X1 U98 ( .B1(n410), .B2(n654), .A(n651), .ZN(n506) );
  NAND2_X1 U99 ( .A1(\mem[4][2] ), .A2(n654), .ZN(n651) );
  OAI21_X1 U100 ( .B1(n409), .B2(n654), .A(n650), .ZN(n505) );
  NAND2_X1 U101 ( .A1(\mem[4][3] ), .A2(n654), .ZN(n650) );
  OAI21_X1 U102 ( .B1(n408), .B2(n654), .A(n649), .ZN(n504) );
  NAND2_X1 U103 ( .A1(\mem[4][4] ), .A2(n654), .ZN(n649) );
  OAI21_X1 U104 ( .B1(n407), .B2(n654), .A(n648), .ZN(n503) );
  NAND2_X1 U105 ( .A1(\mem[4][5] ), .A2(n654), .ZN(n648) );
  OAI21_X1 U106 ( .B1(n406), .B2(n654), .A(n647), .ZN(n502) );
  NAND2_X1 U107 ( .A1(\mem[4][6] ), .A2(n654), .ZN(n647) );
  OAI21_X1 U108 ( .B1(n405), .B2(n654), .A(n646), .ZN(n501) );
  NAND2_X1 U109 ( .A1(\mem[4][7] ), .A2(n654), .ZN(n646) );
  OAI21_X1 U110 ( .B1(n412), .B2(n644), .A(n643), .ZN(n500) );
  NAND2_X1 U111 ( .A1(\mem[5][0] ), .A2(n644), .ZN(n643) );
  OAI21_X1 U112 ( .B1(n411), .B2(n644), .A(n642), .ZN(n499) );
  NAND2_X1 U113 ( .A1(\mem[5][1] ), .A2(n644), .ZN(n642) );
  OAI21_X1 U114 ( .B1(n410), .B2(n644), .A(n641), .ZN(n498) );
  NAND2_X1 U115 ( .A1(\mem[5][2] ), .A2(n644), .ZN(n641) );
  OAI21_X1 U116 ( .B1(n409), .B2(n644), .A(n640), .ZN(n497) );
  NAND2_X1 U117 ( .A1(\mem[5][3] ), .A2(n644), .ZN(n640) );
  OAI21_X1 U118 ( .B1(n408), .B2(n644), .A(n639), .ZN(n496) );
  NAND2_X1 U119 ( .A1(\mem[5][4] ), .A2(n644), .ZN(n639) );
  OAI21_X1 U120 ( .B1(n407), .B2(n644), .A(n638), .ZN(n495) );
  NAND2_X1 U121 ( .A1(\mem[5][5] ), .A2(n644), .ZN(n638) );
  OAI21_X1 U122 ( .B1(n406), .B2(n644), .A(n637), .ZN(n494) );
  NAND2_X1 U123 ( .A1(\mem[5][6] ), .A2(n644), .ZN(n637) );
  OAI21_X1 U124 ( .B1(n405), .B2(n644), .A(n636), .ZN(n493) );
  NAND2_X1 U125 ( .A1(\mem[5][7] ), .A2(n644), .ZN(n636) );
  OAI21_X1 U126 ( .B1(n412), .B2(n635), .A(n634), .ZN(n492) );
  NAND2_X1 U127 ( .A1(\mem[6][0] ), .A2(n635), .ZN(n634) );
  OAI21_X1 U128 ( .B1(n411), .B2(n635), .A(n633), .ZN(n491) );
  NAND2_X1 U129 ( .A1(\mem[6][1] ), .A2(n635), .ZN(n633) );
  OAI21_X1 U130 ( .B1(n410), .B2(n635), .A(n632), .ZN(n490) );
  NAND2_X1 U131 ( .A1(\mem[6][2] ), .A2(n635), .ZN(n632) );
  OAI21_X1 U132 ( .B1(n409), .B2(n635), .A(n631), .ZN(n489) );
  NAND2_X1 U133 ( .A1(\mem[6][3] ), .A2(n635), .ZN(n631) );
  OAI21_X1 U134 ( .B1(n408), .B2(n635), .A(n630), .ZN(n488) );
  NAND2_X1 U135 ( .A1(\mem[6][4] ), .A2(n635), .ZN(n630) );
  OAI21_X1 U136 ( .B1(n407), .B2(n635), .A(n629), .ZN(n487) );
  NAND2_X1 U137 ( .A1(\mem[6][5] ), .A2(n635), .ZN(n629) );
  OAI21_X1 U138 ( .B1(n406), .B2(n635), .A(n628), .ZN(n486) );
  NAND2_X1 U139 ( .A1(\mem[6][6] ), .A2(n635), .ZN(n628) );
  OAI21_X1 U140 ( .B1(n405), .B2(n635), .A(n627), .ZN(n485) );
  NAND2_X1 U141 ( .A1(\mem[6][7] ), .A2(n635), .ZN(n627) );
  OAI21_X1 U142 ( .B1(n412), .B2(n624), .A(n623), .ZN(n484) );
  NAND2_X1 U143 ( .A1(\mem[7][0] ), .A2(n624), .ZN(n623) );
  OAI21_X1 U144 ( .B1(n411), .B2(n624), .A(n622), .ZN(n483) );
  NAND2_X1 U145 ( .A1(\mem[7][1] ), .A2(n624), .ZN(n622) );
  OAI21_X1 U146 ( .B1(n410), .B2(n624), .A(n621), .ZN(n482) );
  NAND2_X1 U147 ( .A1(\mem[7][2] ), .A2(n624), .ZN(n621) );
  OAI21_X1 U148 ( .B1(n409), .B2(n624), .A(n620), .ZN(n481) );
  NAND2_X1 U149 ( .A1(\mem[7][3] ), .A2(n624), .ZN(n620) );
  OAI21_X1 U150 ( .B1(n408), .B2(n624), .A(n619), .ZN(n480) );
  NAND2_X1 U151 ( .A1(\mem[7][4] ), .A2(n624), .ZN(n619) );
  OAI21_X1 U152 ( .B1(n407), .B2(n624), .A(n618), .ZN(n479) );
  NAND2_X1 U153 ( .A1(\mem[7][5] ), .A2(n624), .ZN(n618) );
  OAI21_X1 U154 ( .B1(n406), .B2(n624), .A(n617), .ZN(n478) );
  NAND2_X1 U155 ( .A1(\mem[7][6] ), .A2(n624), .ZN(n617) );
  OAI21_X1 U156 ( .B1(n405), .B2(n624), .A(n616), .ZN(n477) );
  NAND2_X1 U157 ( .A1(\mem[7][7] ), .A2(n624), .ZN(n616) );
  OAI21_X1 U158 ( .B1(n412), .B2(n615), .A(n614), .ZN(n476) );
  NAND2_X1 U159 ( .A1(\mem[8][0] ), .A2(n615), .ZN(n614) );
  OAI21_X1 U160 ( .B1(n411), .B2(n615), .A(n613), .ZN(n475) );
  NAND2_X1 U161 ( .A1(\mem[8][1] ), .A2(n615), .ZN(n613) );
  OAI21_X1 U162 ( .B1(n410), .B2(n615), .A(n612), .ZN(n474) );
  NAND2_X1 U163 ( .A1(\mem[8][2] ), .A2(n615), .ZN(n612) );
  OAI21_X1 U164 ( .B1(n409), .B2(n615), .A(n611), .ZN(n473) );
  NAND2_X1 U165 ( .A1(\mem[8][3] ), .A2(n615), .ZN(n611) );
  OAI21_X1 U166 ( .B1(n408), .B2(n615), .A(n610), .ZN(n472) );
  NAND2_X1 U167 ( .A1(\mem[8][4] ), .A2(n615), .ZN(n610) );
  OAI21_X1 U168 ( .B1(n407), .B2(n615), .A(n609), .ZN(n471) );
  NAND2_X1 U169 ( .A1(\mem[8][5] ), .A2(n615), .ZN(n609) );
  OAI21_X1 U170 ( .B1(n406), .B2(n615), .A(n608), .ZN(n470) );
  NAND2_X1 U171 ( .A1(\mem[8][6] ), .A2(n615), .ZN(n608) );
  OAI21_X1 U172 ( .B1(n405), .B2(n615), .A(n607), .ZN(n469) );
  NAND2_X1 U173 ( .A1(\mem[8][7] ), .A2(n615), .ZN(n607) );
  OAI21_X1 U174 ( .B1(n412), .B2(n605), .A(n604), .ZN(n468) );
  NAND2_X1 U175 ( .A1(\mem[9][0] ), .A2(n605), .ZN(n604) );
  OAI21_X1 U176 ( .B1(n411), .B2(n605), .A(n603), .ZN(n467) );
  NAND2_X1 U177 ( .A1(\mem[9][1] ), .A2(n605), .ZN(n603) );
  OAI21_X1 U178 ( .B1(n410), .B2(n605), .A(n602), .ZN(n466) );
  NAND2_X1 U179 ( .A1(\mem[9][2] ), .A2(n605), .ZN(n602) );
  OAI21_X1 U180 ( .B1(n409), .B2(n605), .A(n601), .ZN(n465) );
  NAND2_X1 U181 ( .A1(\mem[9][3] ), .A2(n605), .ZN(n601) );
  OAI21_X1 U182 ( .B1(n408), .B2(n605), .A(n600), .ZN(n464) );
  NAND2_X1 U183 ( .A1(\mem[9][4] ), .A2(n605), .ZN(n600) );
  OAI21_X1 U184 ( .B1(n407), .B2(n605), .A(n599), .ZN(n463) );
  NAND2_X1 U185 ( .A1(\mem[9][5] ), .A2(n605), .ZN(n599) );
  OAI21_X1 U186 ( .B1(n406), .B2(n605), .A(n598), .ZN(n462) );
  NAND2_X1 U187 ( .A1(\mem[9][6] ), .A2(n605), .ZN(n598) );
  OAI21_X1 U188 ( .B1(n405), .B2(n605), .A(n597), .ZN(n461) );
  NAND2_X1 U189 ( .A1(\mem[9][7] ), .A2(n605), .ZN(n597) );
  OAI21_X1 U190 ( .B1(n412), .B2(n595), .A(n594), .ZN(n460) );
  NAND2_X1 U191 ( .A1(\mem[10][0] ), .A2(n595), .ZN(n594) );
  OAI21_X1 U192 ( .B1(n411), .B2(n595), .A(n593), .ZN(n459) );
  NAND2_X1 U193 ( .A1(\mem[10][1] ), .A2(n595), .ZN(n593) );
  OAI21_X1 U194 ( .B1(n410), .B2(n595), .A(n592), .ZN(n458) );
  NAND2_X1 U195 ( .A1(\mem[10][2] ), .A2(n595), .ZN(n592) );
  OAI21_X1 U196 ( .B1(n409), .B2(n595), .A(n591), .ZN(n457) );
  NAND2_X1 U197 ( .A1(\mem[10][3] ), .A2(n595), .ZN(n591) );
  OAI21_X1 U198 ( .B1(n408), .B2(n595), .A(n590), .ZN(n456) );
  NAND2_X1 U199 ( .A1(\mem[10][4] ), .A2(n595), .ZN(n590) );
  OAI21_X1 U200 ( .B1(n407), .B2(n595), .A(n589), .ZN(n455) );
  NAND2_X1 U201 ( .A1(\mem[10][5] ), .A2(n595), .ZN(n589) );
  OAI21_X1 U202 ( .B1(n406), .B2(n595), .A(n588), .ZN(n454) );
  NAND2_X1 U203 ( .A1(\mem[10][6] ), .A2(n595), .ZN(n588) );
  OAI21_X1 U204 ( .B1(n405), .B2(n595), .A(n587), .ZN(n453) );
  NAND2_X1 U205 ( .A1(\mem[10][7] ), .A2(n595), .ZN(n587) );
  OAI21_X1 U206 ( .B1(n412), .B2(n586), .A(n585), .ZN(n452) );
  NAND2_X1 U207 ( .A1(\mem[11][0] ), .A2(n586), .ZN(n585) );
  OAI21_X1 U208 ( .B1(n411), .B2(n586), .A(n584), .ZN(n451) );
  NAND2_X1 U209 ( .A1(\mem[11][1] ), .A2(n586), .ZN(n584) );
  OAI21_X1 U210 ( .B1(n410), .B2(n586), .A(n583), .ZN(n450) );
  NAND2_X1 U211 ( .A1(\mem[11][2] ), .A2(n586), .ZN(n583) );
  OAI21_X1 U212 ( .B1(n409), .B2(n586), .A(n582), .ZN(n449) );
  NAND2_X1 U213 ( .A1(\mem[11][3] ), .A2(n586), .ZN(n582) );
  OAI21_X1 U214 ( .B1(n408), .B2(n586), .A(n581), .ZN(n448) );
  NAND2_X1 U215 ( .A1(\mem[11][4] ), .A2(n586), .ZN(n581) );
  OAI21_X1 U216 ( .B1(n407), .B2(n586), .A(n580), .ZN(n447) );
  NAND2_X1 U217 ( .A1(\mem[11][5] ), .A2(n586), .ZN(n580) );
  OAI21_X1 U218 ( .B1(n406), .B2(n586), .A(n579), .ZN(n446) );
  NAND2_X1 U219 ( .A1(\mem[11][6] ), .A2(n586), .ZN(n579) );
  OAI21_X1 U220 ( .B1(n405), .B2(n586), .A(n578), .ZN(n445) );
  NAND2_X1 U221 ( .A1(\mem[11][7] ), .A2(n586), .ZN(n578) );
  OAI21_X1 U222 ( .B1(n412), .B2(n577), .A(n576), .ZN(n444) );
  NAND2_X1 U223 ( .A1(\mem[12][0] ), .A2(n577), .ZN(n576) );
  OAI21_X1 U224 ( .B1(n411), .B2(n577), .A(n575), .ZN(n443) );
  NAND2_X1 U225 ( .A1(\mem[12][1] ), .A2(n577), .ZN(n575) );
  OAI21_X1 U226 ( .B1(n410), .B2(n577), .A(n574), .ZN(n442) );
  NAND2_X1 U227 ( .A1(\mem[12][2] ), .A2(n577), .ZN(n574) );
  OAI21_X1 U228 ( .B1(n409), .B2(n577), .A(n573), .ZN(n441) );
  NAND2_X1 U229 ( .A1(\mem[12][3] ), .A2(n577), .ZN(n573) );
  OAI21_X1 U230 ( .B1(n408), .B2(n577), .A(n572), .ZN(n440) );
  NAND2_X1 U231 ( .A1(\mem[12][4] ), .A2(n577), .ZN(n572) );
  OAI21_X1 U232 ( .B1(n407), .B2(n577), .A(n571), .ZN(n439) );
  NAND2_X1 U233 ( .A1(\mem[12][5] ), .A2(n577), .ZN(n571) );
  OAI21_X1 U234 ( .B1(n406), .B2(n577), .A(n570), .ZN(n438) );
  NAND2_X1 U235 ( .A1(\mem[12][6] ), .A2(n577), .ZN(n570) );
  OAI21_X1 U236 ( .B1(n405), .B2(n577), .A(n569), .ZN(n437) );
  NAND2_X1 U237 ( .A1(\mem[12][7] ), .A2(n577), .ZN(n569) );
  OAI21_X1 U238 ( .B1(n412), .B2(n568), .A(n567), .ZN(n436) );
  NAND2_X1 U239 ( .A1(\mem[13][0] ), .A2(n568), .ZN(n567) );
  OAI21_X1 U240 ( .B1(n411), .B2(n568), .A(n566), .ZN(n435) );
  NAND2_X1 U241 ( .A1(\mem[13][1] ), .A2(n568), .ZN(n566) );
  OAI21_X1 U242 ( .B1(n410), .B2(n568), .A(n565), .ZN(n434) );
  NAND2_X1 U243 ( .A1(\mem[13][2] ), .A2(n568), .ZN(n565) );
  OAI21_X1 U244 ( .B1(n409), .B2(n568), .A(n564), .ZN(n433) );
  NAND2_X1 U245 ( .A1(\mem[13][3] ), .A2(n568), .ZN(n564) );
  OAI21_X1 U246 ( .B1(n408), .B2(n568), .A(n563), .ZN(n432) );
  NAND2_X1 U247 ( .A1(\mem[13][4] ), .A2(n568), .ZN(n563) );
  OAI21_X1 U248 ( .B1(n407), .B2(n568), .A(n562), .ZN(n431) );
  NAND2_X1 U249 ( .A1(\mem[13][5] ), .A2(n568), .ZN(n562) );
  OAI21_X1 U250 ( .B1(n406), .B2(n568), .A(n561), .ZN(n430) );
  NAND2_X1 U251 ( .A1(\mem[13][6] ), .A2(n568), .ZN(n561) );
  OAI21_X1 U252 ( .B1(n405), .B2(n568), .A(n560), .ZN(n429) );
  NAND2_X1 U253 ( .A1(\mem[13][7] ), .A2(n568), .ZN(n560) );
  OAI21_X1 U254 ( .B1(n412), .B2(n559), .A(n558), .ZN(n428) );
  NAND2_X1 U255 ( .A1(\mem[14][0] ), .A2(n559), .ZN(n558) );
  OAI21_X1 U256 ( .B1(n411), .B2(n559), .A(n557), .ZN(n427) );
  NAND2_X1 U257 ( .A1(\mem[14][1] ), .A2(n559), .ZN(n557) );
  OAI21_X1 U258 ( .B1(n410), .B2(n559), .A(n556), .ZN(n426) );
  NAND2_X1 U259 ( .A1(\mem[14][2] ), .A2(n559), .ZN(n556) );
  OAI21_X1 U260 ( .B1(n409), .B2(n559), .A(n555), .ZN(n425) );
  NAND2_X1 U261 ( .A1(\mem[14][3] ), .A2(n559), .ZN(n555) );
  OAI21_X1 U262 ( .B1(n408), .B2(n559), .A(n554), .ZN(n424) );
  NAND2_X1 U263 ( .A1(\mem[14][4] ), .A2(n559), .ZN(n554) );
  OAI21_X1 U264 ( .B1(n407), .B2(n559), .A(n553), .ZN(n423) );
  NAND2_X1 U265 ( .A1(\mem[14][5] ), .A2(n559), .ZN(n553) );
  OAI21_X1 U266 ( .B1(n406), .B2(n559), .A(n552), .ZN(n422) );
  NAND2_X1 U267 ( .A1(\mem[14][6] ), .A2(n559), .ZN(n552) );
  OAI21_X1 U268 ( .B1(n405), .B2(n559), .A(n551), .ZN(n421) );
  NAND2_X1 U269 ( .A1(\mem[14][7] ), .A2(n559), .ZN(n551) );
  OAI21_X1 U270 ( .B1(n412), .B2(n549), .A(n548), .ZN(n420) );
  NAND2_X1 U271 ( .A1(\mem[15][0] ), .A2(n549), .ZN(n548) );
  OAI21_X1 U272 ( .B1(n411), .B2(n549), .A(n547), .ZN(n419) );
  NAND2_X1 U273 ( .A1(\mem[15][1] ), .A2(n549), .ZN(n547) );
  OAI21_X1 U274 ( .B1(n410), .B2(n549), .A(n546), .ZN(n418) );
  NAND2_X1 U275 ( .A1(\mem[15][2] ), .A2(n549), .ZN(n546) );
  OAI21_X1 U276 ( .B1(n409), .B2(n549), .A(n545), .ZN(n417) );
  NAND2_X1 U277 ( .A1(\mem[15][3] ), .A2(n549), .ZN(n545) );
  OAI21_X1 U278 ( .B1(n408), .B2(n549), .A(n544), .ZN(n416) );
  NAND2_X1 U279 ( .A1(\mem[15][4] ), .A2(n549), .ZN(n544) );
  OAI21_X1 U280 ( .B1(n407), .B2(n549), .A(n543), .ZN(n415) );
  NAND2_X1 U281 ( .A1(\mem[15][5] ), .A2(n549), .ZN(n543) );
  OAI21_X1 U282 ( .B1(n406), .B2(n549), .A(n542), .ZN(n414) );
  NAND2_X1 U283 ( .A1(\mem[15][6] ), .A2(n549), .ZN(n542) );
  OAI21_X1 U284 ( .B1(n405), .B2(n549), .A(n541), .ZN(n413) );
  NAND2_X1 U285 ( .A1(\mem[15][7] ), .A2(n549), .ZN(n541) );
  AND2_X1 U286 ( .A1(N13), .A2(wr_en), .ZN(n550) );
  NOR2_X1 U287 ( .A1(N11), .A2(N12), .ZN(n685) );
  NOR2_X1 U288 ( .A1(n403), .A2(N12), .ZN(n664) );
  AND2_X1 U289 ( .A1(N12), .A2(n403), .ZN(n645) );
  AND2_X1 U290 ( .A1(N12), .A2(N11), .ZN(n626) );
  INV_X1 U291 ( .A(data_in[0]), .ZN(n412) );
  INV_X1 U292 ( .A(data_in[1]), .ZN(n411) );
  INV_X1 U293 ( .A(data_in[2]), .ZN(n410) );
  INV_X1 U294 ( .A(data_in[3]), .ZN(n409) );
  INV_X1 U295 ( .A(data_in[4]), .ZN(n408) );
  INV_X1 U296 ( .A(data_in[5]), .ZN(n407) );
  INV_X1 U297 ( .A(data_in[6]), .ZN(n406) );
  INV_X1 U298 ( .A(data_in[7]), .ZN(n405) );
  MUX2_X1 U299 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(N10), .Z(n3) );
  MUX2_X1 U300 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(N10), .Z(n4) );
  MUX2_X1 U301 ( .A(n4), .B(n3), .S(N11), .Z(n5) );
  MUX2_X1 U302 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(N10), .Z(n6) );
  MUX2_X1 U303 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n7) );
  MUX2_X1 U304 ( .A(n7), .B(n6), .S(N11), .Z(n8) );
  MUX2_X1 U305 ( .A(n8), .B(n5), .S(N12), .Z(n9) );
  MUX2_X1 U306 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n398), .Z(n10) );
  MUX2_X1 U307 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n398), .Z(n11) );
  MUX2_X1 U308 ( .A(n11), .B(n10), .S(N11), .Z(n294) );
  MUX2_X1 U309 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n398), .Z(n295) );
  MUX2_X1 U310 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n398), .Z(n296) );
  MUX2_X1 U311 ( .A(n296), .B(n295), .S(N11), .Z(n297) );
  MUX2_X1 U312 ( .A(n297), .B(n294), .S(N12), .Z(n298) );
  MUX2_X1 U313 ( .A(n298), .B(n9), .S(N13), .Z(N21) );
  MUX2_X1 U314 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n398), .Z(n299) );
  MUX2_X1 U315 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n398), .Z(n300) );
  MUX2_X1 U316 ( .A(n300), .B(n299), .S(N11), .Z(n301) );
  MUX2_X1 U317 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n398), .Z(n302) );
  MUX2_X1 U318 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n398), .Z(n303) );
  MUX2_X1 U319 ( .A(n303), .B(n302), .S(N11), .Z(n304) );
  MUX2_X1 U320 ( .A(n304), .B(n301), .S(N12), .Z(n305) );
  MUX2_X1 U321 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n398), .Z(n306) );
  MUX2_X1 U322 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n398), .Z(n307) );
  MUX2_X1 U323 ( .A(n307), .B(n306), .S(N11), .Z(n308) );
  MUX2_X1 U324 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n398), .Z(n309) );
  MUX2_X1 U325 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n398), .Z(n310) );
  MUX2_X1 U326 ( .A(n310), .B(n309), .S(N11), .Z(n311) );
  MUX2_X1 U327 ( .A(n311), .B(n308), .S(N12), .Z(n312) );
  MUX2_X1 U328 ( .A(n312), .B(n305), .S(N13), .Z(N20) );
  MUX2_X1 U329 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n399), .Z(n313) );
  MUX2_X1 U330 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n399), .Z(n314) );
  MUX2_X1 U331 ( .A(n314), .B(n313), .S(n397), .Z(n315) );
  MUX2_X1 U332 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n399), .Z(n316) );
  MUX2_X1 U333 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n399), .Z(n317) );
  MUX2_X1 U334 ( .A(n317), .B(n316), .S(n397), .Z(n318) );
  MUX2_X1 U335 ( .A(n318), .B(n315), .S(N12), .Z(n319) );
  MUX2_X1 U336 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n399), .Z(n320) );
  MUX2_X1 U337 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n399), .Z(n321) );
  MUX2_X1 U338 ( .A(n321), .B(n320), .S(n397), .Z(n322) );
  MUX2_X1 U339 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n399), .Z(n323) );
  MUX2_X1 U340 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n399), .Z(n324) );
  MUX2_X1 U341 ( .A(n324), .B(n323), .S(n397), .Z(n325) );
  MUX2_X1 U342 ( .A(n325), .B(n322), .S(N12), .Z(n326) );
  MUX2_X1 U343 ( .A(n326), .B(n319), .S(N13), .Z(N19) );
  MUX2_X1 U344 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n399), .Z(n327) );
  MUX2_X1 U345 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n399), .Z(n328) );
  MUX2_X1 U346 ( .A(n328), .B(n327), .S(n397), .Z(n329) );
  MUX2_X1 U347 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n399), .Z(n330) );
  MUX2_X1 U348 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n399), .Z(n331) );
  MUX2_X1 U349 ( .A(n331), .B(n330), .S(n397), .Z(n332) );
  MUX2_X1 U350 ( .A(n332), .B(n329), .S(N12), .Z(n333) );
  MUX2_X1 U351 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n400), .Z(n334) );
  MUX2_X1 U352 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n400), .Z(n335) );
  MUX2_X1 U353 ( .A(n335), .B(n334), .S(n397), .Z(n336) );
  MUX2_X1 U354 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n400), .Z(n337) );
  MUX2_X1 U355 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n400), .Z(n338) );
  MUX2_X1 U356 ( .A(n338), .B(n337), .S(n397), .Z(n339) );
  MUX2_X1 U357 ( .A(n339), .B(n336), .S(N12), .Z(n340) );
  MUX2_X1 U358 ( .A(n340), .B(n333), .S(N13), .Z(N18) );
  MUX2_X1 U359 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n400), .Z(n341) );
  MUX2_X1 U360 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n400), .Z(n342) );
  MUX2_X1 U361 ( .A(n342), .B(n341), .S(n397), .Z(n343) );
  MUX2_X1 U362 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n400), .Z(n344) );
  MUX2_X1 U363 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n400), .Z(n345) );
  MUX2_X1 U364 ( .A(n345), .B(n344), .S(n397), .Z(n346) );
  MUX2_X1 U365 ( .A(n346), .B(n343), .S(N12), .Z(n347) );
  MUX2_X1 U366 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n400), .Z(n348) );
  MUX2_X1 U367 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n400), .Z(n349) );
  MUX2_X1 U368 ( .A(n349), .B(n348), .S(n397), .Z(n350) );
  MUX2_X1 U369 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n400), .Z(n351) );
  MUX2_X1 U370 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n400), .Z(n352) );
  MUX2_X1 U371 ( .A(n352), .B(n351), .S(n397), .Z(n353) );
  MUX2_X1 U372 ( .A(n353), .B(n350), .S(N12), .Z(n354) );
  MUX2_X1 U373 ( .A(n354), .B(n347), .S(N13), .Z(N17) );
  MUX2_X1 U374 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n398), .Z(n355) );
  MUX2_X1 U375 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n399), .Z(n356) );
  MUX2_X1 U376 ( .A(n356), .B(n355), .S(N11), .Z(n357) );
  MUX2_X1 U377 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n399), .Z(n358) );
  MUX2_X1 U378 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n398), .Z(n359) );
  MUX2_X1 U379 ( .A(n359), .B(n358), .S(N11), .Z(n360) );
  MUX2_X1 U380 ( .A(n360), .B(n357), .S(N12), .Z(n361) );
  MUX2_X1 U381 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n398), .Z(n362) );
  MUX2_X1 U382 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n400), .Z(n363) );
  MUX2_X1 U383 ( .A(n363), .B(n362), .S(N11), .Z(n364) );
  MUX2_X1 U384 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n398), .Z(n365) );
  MUX2_X1 U385 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n399), .Z(n366) );
  MUX2_X1 U386 ( .A(n366), .B(n365), .S(n397), .Z(n367) );
  MUX2_X1 U387 ( .A(n367), .B(n364), .S(N12), .Z(n368) );
  MUX2_X1 U388 ( .A(n368), .B(n361), .S(N13), .Z(N16) );
  MUX2_X1 U389 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(N10), .Z(n369) );
  MUX2_X1 U390 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n400), .Z(n370) );
  MUX2_X1 U391 ( .A(n370), .B(n369), .S(N11), .Z(n371) );
  MUX2_X1 U392 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n400), .Z(n372) );
  MUX2_X1 U393 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n399), .Z(n373) );
  MUX2_X1 U394 ( .A(n373), .B(n372), .S(N11), .Z(n374) );
  MUX2_X1 U395 ( .A(n374), .B(n371), .S(N12), .Z(n375) );
  MUX2_X1 U396 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n376) );
  MUX2_X1 U397 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n377) );
  MUX2_X1 U398 ( .A(n377), .B(n376), .S(N11), .Z(n378) );
  MUX2_X1 U399 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n379) );
  MUX2_X1 U400 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n399), .Z(n380) );
  MUX2_X1 U401 ( .A(n380), .B(n379), .S(n397), .Z(n381) );
  MUX2_X1 U402 ( .A(n381), .B(n378), .S(N12), .Z(n382) );
  MUX2_X1 U403 ( .A(n382), .B(n375), .S(N13), .Z(N15) );
  MUX2_X1 U404 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(N10), .Z(n383) );
  MUX2_X1 U405 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n384) );
  MUX2_X1 U406 ( .A(n384), .B(n383), .S(N11), .Z(n385) );
  MUX2_X1 U407 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(N10), .Z(n386) );
  MUX2_X1 U408 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n387) );
  MUX2_X1 U409 ( .A(n387), .B(n386), .S(N11), .Z(n388) );
  MUX2_X1 U410 ( .A(n388), .B(n385), .S(N12), .Z(n389) );
  MUX2_X1 U411 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n390) );
  MUX2_X1 U412 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n391) );
  MUX2_X1 U413 ( .A(n391), .B(n390), .S(N11), .Z(n392) );
  MUX2_X1 U414 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n393) );
  MUX2_X1 U415 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n400), .Z(n394) );
  MUX2_X1 U416 ( .A(n394), .B(n393), .S(n397), .Z(n395) );
  MUX2_X1 U417 ( .A(n395), .B(n392), .S(N12), .Z(n396) );
  MUX2_X1 U418 ( .A(n396), .B(n389), .S(N13), .Z(N14) );
  INV_X1 U419 ( .A(N10), .ZN(n402) );
  INV_X1 U420 ( .A(N11), .ZN(n403) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_4 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, N19, N20, N21, n1, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N16), .CK(clk), .QN(n1) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n412), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n413), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n414), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n415), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n416), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n417), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n418), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n419), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n420), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n421), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n422), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n423), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n424), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n425), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n426), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n427), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n428), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n429), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n430), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n431), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n432), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n433), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n434), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n435), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n436), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n437), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n438), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n439), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n440), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n441), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n442), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n443), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n444), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n445), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n446), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n447), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n448), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n449), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n450), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n451), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n452), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n453), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n454), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n455), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n456), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n457), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n458), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n459), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n460), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n461), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n462), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n463), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n464), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n465), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n466), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n467), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n468), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n469), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n470), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n471), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n472), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n473), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n474), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n475), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n476), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n477), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n478), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n479), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n480), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n481), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n482), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n483), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n484), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n485), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n486), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n487), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n488), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n489), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n490), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n491), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n492), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n493), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n494), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n495), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n496), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n497), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n498), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n499), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n500), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n501), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n502), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n503), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n504), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n505), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n506), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n507), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n508), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n509), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n510), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n511), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n512), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n513), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n514), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n515), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n516), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n517), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n518), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n519), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n520), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n521), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n522), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n523), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n524), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n525), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n526), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n527), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n528), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n529), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n530), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n531), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n532), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n533), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n534), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n535), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n536), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n537), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n538), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n539), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N18), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[1]  ( .D(N20), .CK(clk), .Q(data_out[1]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[5]) );
  BUF_X1 U4 ( .A(N10), .Z(n398) );
  BUF_X1 U5 ( .A(N10), .Z(n399) );
  BUF_X1 U6 ( .A(N10), .Z(n400) );
  BUF_X1 U7 ( .A(N11), .Z(n397) );
  NAND2_X1 U8 ( .A1(n663), .A2(n683), .ZN(n672) );
  NAND2_X1 U9 ( .A1(n663), .A2(n673), .ZN(n662) );
  NAND2_X1 U10 ( .A1(n684), .A2(n683), .ZN(n693) );
  NAND2_X1 U11 ( .A1(n673), .A2(n684), .ZN(n682) );
  NAND2_X1 U12 ( .A1(n605), .A2(n684), .ZN(n614) );
  NAND2_X1 U13 ( .A1(n595), .A2(n684), .ZN(n604) );
  NAND2_X1 U14 ( .A1(n605), .A2(n663), .ZN(n594) );
  NAND2_X1 U15 ( .A1(n595), .A2(n663), .ZN(n585) );
  NAND2_X1 U16 ( .A1(n644), .A2(n683), .ZN(n653) );
  NAND2_X1 U17 ( .A1(n644), .A2(n673), .ZN(n643) );
  NAND2_X1 U18 ( .A1(n625), .A2(n683), .ZN(n634) );
  NAND2_X1 U19 ( .A1(n625), .A2(n673), .ZN(n623) );
  NAND2_X1 U20 ( .A1(n605), .A2(n644), .ZN(n576) );
  NAND2_X1 U21 ( .A1(n595), .A2(n644), .ZN(n567) );
  NAND2_X1 U22 ( .A1(n605), .A2(n625), .ZN(n558) );
  NAND2_X1 U23 ( .A1(n595), .A2(n625), .ZN(n548) );
  AND2_X1 U24 ( .A1(n549), .A2(N10), .ZN(n595) );
  AND2_X1 U25 ( .A1(n549), .A2(n401), .ZN(n605) );
  AND2_X1 U26 ( .A1(N10), .A2(n624), .ZN(n673) );
  AND2_X1 U27 ( .A1(n624), .A2(n401), .ZN(n683) );
  OAI21_X1 U28 ( .B1(n693), .B2(n411), .A(n692), .ZN(n539) );
  NAND2_X1 U29 ( .A1(\mem[0][0] ), .A2(n693), .ZN(n692) );
  OAI21_X1 U30 ( .B1(n693), .B2(n410), .A(n691), .ZN(n538) );
  NAND2_X1 U31 ( .A1(\mem[0][1] ), .A2(n693), .ZN(n691) );
  OAI21_X1 U32 ( .B1(n693), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U33 ( .A1(\mem[0][2] ), .A2(n693), .ZN(n690) );
  OAI21_X1 U34 ( .B1(n693), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U35 ( .A1(\mem[0][3] ), .A2(n693), .ZN(n689) );
  OAI21_X1 U36 ( .B1(n693), .B2(n407), .A(n688), .ZN(n535) );
  NAND2_X1 U37 ( .A1(\mem[0][4] ), .A2(n693), .ZN(n688) );
  OAI21_X1 U38 ( .B1(n693), .B2(n406), .A(n687), .ZN(n534) );
  NAND2_X1 U39 ( .A1(\mem[0][5] ), .A2(n693), .ZN(n687) );
  OAI21_X1 U40 ( .B1(n693), .B2(n405), .A(n686), .ZN(n533) );
  NAND2_X1 U41 ( .A1(\mem[0][6] ), .A2(n693), .ZN(n686) );
  OAI21_X1 U42 ( .B1(n693), .B2(n404), .A(n685), .ZN(n532) );
  NAND2_X1 U43 ( .A1(\mem[0][7] ), .A2(n693), .ZN(n685) );
  OAI21_X1 U44 ( .B1(n411), .B2(n672), .A(n671), .ZN(n523) );
  NAND2_X1 U45 ( .A1(\mem[2][0] ), .A2(n672), .ZN(n671) );
  OAI21_X1 U46 ( .B1(n410), .B2(n672), .A(n670), .ZN(n522) );
  NAND2_X1 U47 ( .A1(\mem[2][1] ), .A2(n672), .ZN(n670) );
  OAI21_X1 U48 ( .B1(n409), .B2(n672), .A(n669), .ZN(n521) );
  NAND2_X1 U49 ( .A1(\mem[2][2] ), .A2(n672), .ZN(n669) );
  OAI21_X1 U50 ( .B1(n408), .B2(n672), .A(n668), .ZN(n520) );
  NAND2_X1 U51 ( .A1(\mem[2][3] ), .A2(n672), .ZN(n668) );
  OAI21_X1 U52 ( .B1(n407), .B2(n672), .A(n667), .ZN(n519) );
  NAND2_X1 U53 ( .A1(\mem[2][4] ), .A2(n672), .ZN(n667) );
  OAI21_X1 U54 ( .B1(n406), .B2(n672), .A(n666), .ZN(n518) );
  NAND2_X1 U55 ( .A1(\mem[2][5] ), .A2(n672), .ZN(n666) );
  OAI21_X1 U56 ( .B1(n405), .B2(n672), .A(n665), .ZN(n517) );
  NAND2_X1 U57 ( .A1(\mem[2][6] ), .A2(n672), .ZN(n665) );
  OAI21_X1 U58 ( .B1(n404), .B2(n672), .A(n664), .ZN(n516) );
  NAND2_X1 U59 ( .A1(\mem[2][7] ), .A2(n672), .ZN(n664) );
  OAI21_X1 U60 ( .B1(n411), .B2(n662), .A(n661), .ZN(n515) );
  NAND2_X1 U61 ( .A1(\mem[3][0] ), .A2(n662), .ZN(n661) );
  OAI21_X1 U62 ( .B1(n410), .B2(n662), .A(n660), .ZN(n514) );
  NAND2_X1 U63 ( .A1(\mem[3][1] ), .A2(n662), .ZN(n660) );
  OAI21_X1 U64 ( .B1(n409), .B2(n662), .A(n659), .ZN(n513) );
  NAND2_X1 U65 ( .A1(\mem[3][2] ), .A2(n662), .ZN(n659) );
  OAI21_X1 U66 ( .B1(n408), .B2(n662), .A(n658), .ZN(n512) );
  NAND2_X1 U67 ( .A1(\mem[3][3] ), .A2(n662), .ZN(n658) );
  OAI21_X1 U68 ( .B1(n407), .B2(n662), .A(n657), .ZN(n511) );
  NAND2_X1 U69 ( .A1(\mem[3][4] ), .A2(n662), .ZN(n657) );
  OAI21_X1 U70 ( .B1(n406), .B2(n662), .A(n656), .ZN(n510) );
  NAND2_X1 U71 ( .A1(\mem[3][5] ), .A2(n662), .ZN(n656) );
  OAI21_X1 U72 ( .B1(n405), .B2(n662), .A(n655), .ZN(n509) );
  NAND2_X1 U73 ( .A1(\mem[3][6] ), .A2(n662), .ZN(n655) );
  OAI21_X1 U74 ( .B1(n404), .B2(n662), .A(n654), .ZN(n508) );
  NAND2_X1 U75 ( .A1(\mem[3][7] ), .A2(n662), .ZN(n654) );
  NOR2_X1 U76 ( .A1(n403), .A2(N13), .ZN(n624) );
  INV_X1 U77 ( .A(wr_en), .ZN(n403) );
  OAI21_X1 U78 ( .B1(n411), .B2(n682), .A(n681), .ZN(n531) );
  NAND2_X1 U79 ( .A1(\mem[1][0] ), .A2(n682), .ZN(n681) );
  OAI21_X1 U80 ( .B1(n410), .B2(n682), .A(n680), .ZN(n530) );
  NAND2_X1 U81 ( .A1(\mem[1][1] ), .A2(n682), .ZN(n680) );
  OAI21_X1 U82 ( .B1(n409), .B2(n682), .A(n679), .ZN(n529) );
  NAND2_X1 U83 ( .A1(\mem[1][2] ), .A2(n682), .ZN(n679) );
  OAI21_X1 U84 ( .B1(n408), .B2(n682), .A(n678), .ZN(n528) );
  NAND2_X1 U85 ( .A1(\mem[1][3] ), .A2(n682), .ZN(n678) );
  OAI21_X1 U86 ( .B1(n407), .B2(n682), .A(n677), .ZN(n527) );
  NAND2_X1 U87 ( .A1(\mem[1][4] ), .A2(n682), .ZN(n677) );
  OAI21_X1 U88 ( .B1(n406), .B2(n682), .A(n676), .ZN(n526) );
  NAND2_X1 U89 ( .A1(\mem[1][5] ), .A2(n682), .ZN(n676) );
  OAI21_X1 U90 ( .B1(n405), .B2(n682), .A(n675), .ZN(n525) );
  NAND2_X1 U91 ( .A1(\mem[1][6] ), .A2(n682), .ZN(n675) );
  OAI21_X1 U92 ( .B1(n404), .B2(n682), .A(n674), .ZN(n524) );
  NAND2_X1 U93 ( .A1(\mem[1][7] ), .A2(n682), .ZN(n674) );
  OAI21_X1 U94 ( .B1(n411), .B2(n653), .A(n652), .ZN(n507) );
  NAND2_X1 U95 ( .A1(\mem[4][0] ), .A2(n653), .ZN(n652) );
  OAI21_X1 U96 ( .B1(n410), .B2(n653), .A(n651), .ZN(n506) );
  NAND2_X1 U97 ( .A1(\mem[4][1] ), .A2(n653), .ZN(n651) );
  OAI21_X1 U98 ( .B1(n409), .B2(n653), .A(n650), .ZN(n505) );
  NAND2_X1 U99 ( .A1(\mem[4][2] ), .A2(n653), .ZN(n650) );
  OAI21_X1 U100 ( .B1(n408), .B2(n653), .A(n649), .ZN(n504) );
  NAND2_X1 U101 ( .A1(\mem[4][3] ), .A2(n653), .ZN(n649) );
  OAI21_X1 U102 ( .B1(n407), .B2(n653), .A(n648), .ZN(n503) );
  NAND2_X1 U103 ( .A1(\mem[4][4] ), .A2(n653), .ZN(n648) );
  OAI21_X1 U104 ( .B1(n406), .B2(n653), .A(n647), .ZN(n502) );
  NAND2_X1 U105 ( .A1(\mem[4][5] ), .A2(n653), .ZN(n647) );
  OAI21_X1 U106 ( .B1(n405), .B2(n653), .A(n646), .ZN(n501) );
  NAND2_X1 U107 ( .A1(\mem[4][6] ), .A2(n653), .ZN(n646) );
  OAI21_X1 U108 ( .B1(n404), .B2(n653), .A(n645), .ZN(n500) );
  NAND2_X1 U109 ( .A1(\mem[4][7] ), .A2(n653), .ZN(n645) );
  OAI21_X1 U110 ( .B1(n411), .B2(n643), .A(n642), .ZN(n499) );
  NAND2_X1 U111 ( .A1(\mem[5][0] ), .A2(n643), .ZN(n642) );
  OAI21_X1 U112 ( .B1(n410), .B2(n643), .A(n641), .ZN(n498) );
  NAND2_X1 U113 ( .A1(\mem[5][1] ), .A2(n643), .ZN(n641) );
  OAI21_X1 U114 ( .B1(n409), .B2(n643), .A(n640), .ZN(n497) );
  NAND2_X1 U115 ( .A1(\mem[5][2] ), .A2(n643), .ZN(n640) );
  OAI21_X1 U116 ( .B1(n408), .B2(n643), .A(n639), .ZN(n496) );
  NAND2_X1 U117 ( .A1(\mem[5][3] ), .A2(n643), .ZN(n639) );
  OAI21_X1 U118 ( .B1(n407), .B2(n643), .A(n638), .ZN(n495) );
  NAND2_X1 U119 ( .A1(\mem[5][4] ), .A2(n643), .ZN(n638) );
  OAI21_X1 U120 ( .B1(n406), .B2(n643), .A(n637), .ZN(n494) );
  NAND2_X1 U121 ( .A1(\mem[5][5] ), .A2(n643), .ZN(n637) );
  OAI21_X1 U122 ( .B1(n405), .B2(n643), .A(n636), .ZN(n493) );
  NAND2_X1 U123 ( .A1(\mem[5][6] ), .A2(n643), .ZN(n636) );
  OAI21_X1 U124 ( .B1(n404), .B2(n643), .A(n635), .ZN(n492) );
  NAND2_X1 U125 ( .A1(\mem[5][7] ), .A2(n643), .ZN(n635) );
  OAI21_X1 U126 ( .B1(n411), .B2(n634), .A(n633), .ZN(n491) );
  NAND2_X1 U127 ( .A1(\mem[6][0] ), .A2(n634), .ZN(n633) );
  OAI21_X1 U128 ( .B1(n410), .B2(n634), .A(n632), .ZN(n490) );
  NAND2_X1 U129 ( .A1(\mem[6][1] ), .A2(n634), .ZN(n632) );
  OAI21_X1 U130 ( .B1(n409), .B2(n634), .A(n631), .ZN(n489) );
  NAND2_X1 U131 ( .A1(\mem[6][2] ), .A2(n634), .ZN(n631) );
  OAI21_X1 U132 ( .B1(n408), .B2(n634), .A(n630), .ZN(n488) );
  NAND2_X1 U133 ( .A1(\mem[6][3] ), .A2(n634), .ZN(n630) );
  OAI21_X1 U134 ( .B1(n407), .B2(n634), .A(n629), .ZN(n487) );
  NAND2_X1 U135 ( .A1(\mem[6][4] ), .A2(n634), .ZN(n629) );
  OAI21_X1 U136 ( .B1(n406), .B2(n634), .A(n628), .ZN(n486) );
  NAND2_X1 U137 ( .A1(\mem[6][5] ), .A2(n634), .ZN(n628) );
  OAI21_X1 U138 ( .B1(n405), .B2(n634), .A(n627), .ZN(n485) );
  NAND2_X1 U139 ( .A1(\mem[6][6] ), .A2(n634), .ZN(n627) );
  OAI21_X1 U140 ( .B1(n404), .B2(n634), .A(n626), .ZN(n484) );
  NAND2_X1 U141 ( .A1(\mem[6][7] ), .A2(n634), .ZN(n626) );
  OAI21_X1 U142 ( .B1(n411), .B2(n623), .A(n622), .ZN(n483) );
  NAND2_X1 U143 ( .A1(\mem[7][0] ), .A2(n623), .ZN(n622) );
  OAI21_X1 U144 ( .B1(n410), .B2(n623), .A(n621), .ZN(n482) );
  NAND2_X1 U145 ( .A1(\mem[7][1] ), .A2(n623), .ZN(n621) );
  OAI21_X1 U146 ( .B1(n409), .B2(n623), .A(n620), .ZN(n481) );
  NAND2_X1 U147 ( .A1(\mem[7][2] ), .A2(n623), .ZN(n620) );
  OAI21_X1 U148 ( .B1(n408), .B2(n623), .A(n619), .ZN(n480) );
  NAND2_X1 U149 ( .A1(\mem[7][3] ), .A2(n623), .ZN(n619) );
  OAI21_X1 U150 ( .B1(n407), .B2(n623), .A(n618), .ZN(n479) );
  NAND2_X1 U151 ( .A1(\mem[7][4] ), .A2(n623), .ZN(n618) );
  OAI21_X1 U152 ( .B1(n406), .B2(n623), .A(n617), .ZN(n478) );
  NAND2_X1 U153 ( .A1(\mem[7][5] ), .A2(n623), .ZN(n617) );
  OAI21_X1 U154 ( .B1(n405), .B2(n623), .A(n616), .ZN(n477) );
  NAND2_X1 U155 ( .A1(\mem[7][6] ), .A2(n623), .ZN(n616) );
  OAI21_X1 U156 ( .B1(n404), .B2(n623), .A(n615), .ZN(n476) );
  NAND2_X1 U157 ( .A1(\mem[7][7] ), .A2(n623), .ZN(n615) );
  OAI21_X1 U158 ( .B1(n411), .B2(n614), .A(n613), .ZN(n475) );
  NAND2_X1 U159 ( .A1(\mem[8][0] ), .A2(n614), .ZN(n613) );
  OAI21_X1 U160 ( .B1(n410), .B2(n614), .A(n612), .ZN(n474) );
  NAND2_X1 U161 ( .A1(\mem[8][1] ), .A2(n614), .ZN(n612) );
  OAI21_X1 U162 ( .B1(n409), .B2(n614), .A(n611), .ZN(n473) );
  NAND2_X1 U163 ( .A1(\mem[8][2] ), .A2(n614), .ZN(n611) );
  OAI21_X1 U164 ( .B1(n408), .B2(n614), .A(n610), .ZN(n472) );
  NAND2_X1 U165 ( .A1(\mem[8][3] ), .A2(n614), .ZN(n610) );
  OAI21_X1 U166 ( .B1(n407), .B2(n614), .A(n609), .ZN(n471) );
  NAND2_X1 U167 ( .A1(\mem[8][4] ), .A2(n614), .ZN(n609) );
  OAI21_X1 U168 ( .B1(n406), .B2(n614), .A(n608), .ZN(n470) );
  NAND2_X1 U169 ( .A1(\mem[8][5] ), .A2(n614), .ZN(n608) );
  OAI21_X1 U170 ( .B1(n405), .B2(n614), .A(n607), .ZN(n469) );
  NAND2_X1 U171 ( .A1(\mem[8][6] ), .A2(n614), .ZN(n607) );
  OAI21_X1 U172 ( .B1(n404), .B2(n614), .A(n606), .ZN(n468) );
  NAND2_X1 U173 ( .A1(\mem[8][7] ), .A2(n614), .ZN(n606) );
  OAI21_X1 U174 ( .B1(n411), .B2(n604), .A(n603), .ZN(n467) );
  NAND2_X1 U175 ( .A1(\mem[9][0] ), .A2(n604), .ZN(n603) );
  OAI21_X1 U176 ( .B1(n410), .B2(n604), .A(n602), .ZN(n466) );
  NAND2_X1 U177 ( .A1(\mem[9][1] ), .A2(n604), .ZN(n602) );
  OAI21_X1 U178 ( .B1(n409), .B2(n604), .A(n601), .ZN(n465) );
  NAND2_X1 U179 ( .A1(\mem[9][2] ), .A2(n604), .ZN(n601) );
  OAI21_X1 U180 ( .B1(n408), .B2(n604), .A(n600), .ZN(n464) );
  NAND2_X1 U181 ( .A1(\mem[9][3] ), .A2(n604), .ZN(n600) );
  OAI21_X1 U182 ( .B1(n407), .B2(n604), .A(n599), .ZN(n463) );
  NAND2_X1 U183 ( .A1(\mem[9][4] ), .A2(n604), .ZN(n599) );
  OAI21_X1 U184 ( .B1(n406), .B2(n604), .A(n598), .ZN(n462) );
  NAND2_X1 U185 ( .A1(\mem[9][5] ), .A2(n604), .ZN(n598) );
  OAI21_X1 U186 ( .B1(n405), .B2(n604), .A(n597), .ZN(n461) );
  NAND2_X1 U187 ( .A1(\mem[9][6] ), .A2(n604), .ZN(n597) );
  OAI21_X1 U188 ( .B1(n404), .B2(n604), .A(n596), .ZN(n460) );
  NAND2_X1 U189 ( .A1(\mem[9][7] ), .A2(n604), .ZN(n596) );
  OAI21_X1 U190 ( .B1(n411), .B2(n594), .A(n593), .ZN(n459) );
  NAND2_X1 U191 ( .A1(\mem[10][0] ), .A2(n594), .ZN(n593) );
  OAI21_X1 U192 ( .B1(n410), .B2(n594), .A(n592), .ZN(n458) );
  NAND2_X1 U193 ( .A1(\mem[10][1] ), .A2(n594), .ZN(n592) );
  OAI21_X1 U194 ( .B1(n409), .B2(n594), .A(n591), .ZN(n457) );
  NAND2_X1 U195 ( .A1(\mem[10][2] ), .A2(n594), .ZN(n591) );
  OAI21_X1 U196 ( .B1(n408), .B2(n594), .A(n590), .ZN(n456) );
  NAND2_X1 U197 ( .A1(\mem[10][3] ), .A2(n594), .ZN(n590) );
  OAI21_X1 U198 ( .B1(n407), .B2(n594), .A(n589), .ZN(n455) );
  NAND2_X1 U199 ( .A1(\mem[10][4] ), .A2(n594), .ZN(n589) );
  OAI21_X1 U200 ( .B1(n406), .B2(n594), .A(n588), .ZN(n454) );
  NAND2_X1 U201 ( .A1(\mem[10][5] ), .A2(n594), .ZN(n588) );
  OAI21_X1 U202 ( .B1(n405), .B2(n594), .A(n587), .ZN(n453) );
  NAND2_X1 U203 ( .A1(\mem[10][6] ), .A2(n594), .ZN(n587) );
  OAI21_X1 U204 ( .B1(n404), .B2(n594), .A(n586), .ZN(n452) );
  NAND2_X1 U205 ( .A1(\mem[10][7] ), .A2(n594), .ZN(n586) );
  OAI21_X1 U206 ( .B1(n411), .B2(n585), .A(n584), .ZN(n451) );
  NAND2_X1 U207 ( .A1(\mem[11][0] ), .A2(n585), .ZN(n584) );
  OAI21_X1 U208 ( .B1(n410), .B2(n585), .A(n583), .ZN(n450) );
  NAND2_X1 U209 ( .A1(\mem[11][1] ), .A2(n585), .ZN(n583) );
  OAI21_X1 U210 ( .B1(n409), .B2(n585), .A(n582), .ZN(n449) );
  NAND2_X1 U211 ( .A1(\mem[11][2] ), .A2(n585), .ZN(n582) );
  OAI21_X1 U212 ( .B1(n408), .B2(n585), .A(n581), .ZN(n448) );
  NAND2_X1 U213 ( .A1(\mem[11][3] ), .A2(n585), .ZN(n581) );
  OAI21_X1 U214 ( .B1(n407), .B2(n585), .A(n580), .ZN(n447) );
  NAND2_X1 U215 ( .A1(\mem[11][4] ), .A2(n585), .ZN(n580) );
  OAI21_X1 U216 ( .B1(n406), .B2(n585), .A(n579), .ZN(n446) );
  NAND2_X1 U217 ( .A1(\mem[11][5] ), .A2(n585), .ZN(n579) );
  OAI21_X1 U218 ( .B1(n405), .B2(n585), .A(n578), .ZN(n445) );
  NAND2_X1 U219 ( .A1(\mem[11][6] ), .A2(n585), .ZN(n578) );
  OAI21_X1 U220 ( .B1(n404), .B2(n585), .A(n577), .ZN(n444) );
  NAND2_X1 U221 ( .A1(\mem[11][7] ), .A2(n585), .ZN(n577) );
  OAI21_X1 U222 ( .B1(n411), .B2(n576), .A(n575), .ZN(n443) );
  NAND2_X1 U223 ( .A1(\mem[12][0] ), .A2(n576), .ZN(n575) );
  OAI21_X1 U224 ( .B1(n410), .B2(n576), .A(n574), .ZN(n442) );
  NAND2_X1 U225 ( .A1(\mem[12][1] ), .A2(n576), .ZN(n574) );
  OAI21_X1 U226 ( .B1(n409), .B2(n576), .A(n573), .ZN(n441) );
  NAND2_X1 U227 ( .A1(\mem[12][2] ), .A2(n576), .ZN(n573) );
  OAI21_X1 U228 ( .B1(n408), .B2(n576), .A(n572), .ZN(n440) );
  NAND2_X1 U229 ( .A1(\mem[12][3] ), .A2(n576), .ZN(n572) );
  OAI21_X1 U230 ( .B1(n407), .B2(n576), .A(n571), .ZN(n439) );
  NAND2_X1 U231 ( .A1(\mem[12][4] ), .A2(n576), .ZN(n571) );
  OAI21_X1 U232 ( .B1(n406), .B2(n576), .A(n570), .ZN(n438) );
  NAND2_X1 U233 ( .A1(\mem[12][5] ), .A2(n576), .ZN(n570) );
  OAI21_X1 U234 ( .B1(n405), .B2(n576), .A(n569), .ZN(n437) );
  NAND2_X1 U235 ( .A1(\mem[12][6] ), .A2(n576), .ZN(n569) );
  OAI21_X1 U236 ( .B1(n404), .B2(n576), .A(n568), .ZN(n436) );
  NAND2_X1 U237 ( .A1(\mem[12][7] ), .A2(n576), .ZN(n568) );
  OAI21_X1 U238 ( .B1(n411), .B2(n567), .A(n566), .ZN(n435) );
  NAND2_X1 U239 ( .A1(\mem[13][0] ), .A2(n567), .ZN(n566) );
  OAI21_X1 U240 ( .B1(n410), .B2(n567), .A(n565), .ZN(n434) );
  NAND2_X1 U241 ( .A1(\mem[13][1] ), .A2(n567), .ZN(n565) );
  OAI21_X1 U242 ( .B1(n409), .B2(n567), .A(n564), .ZN(n433) );
  NAND2_X1 U243 ( .A1(\mem[13][2] ), .A2(n567), .ZN(n564) );
  OAI21_X1 U244 ( .B1(n408), .B2(n567), .A(n563), .ZN(n432) );
  NAND2_X1 U245 ( .A1(\mem[13][3] ), .A2(n567), .ZN(n563) );
  OAI21_X1 U246 ( .B1(n407), .B2(n567), .A(n562), .ZN(n431) );
  NAND2_X1 U247 ( .A1(\mem[13][4] ), .A2(n567), .ZN(n562) );
  OAI21_X1 U248 ( .B1(n406), .B2(n567), .A(n561), .ZN(n430) );
  NAND2_X1 U249 ( .A1(\mem[13][5] ), .A2(n567), .ZN(n561) );
  OAI21_X1 U250 ( .B1(n405), .B2(n567), .A(n560), .ZN(n429) );
  NAND2_X1 U251 ( .A1(\mem[13][6] ), .A2(n567), .ZN(n560) );
  OAI21_X1 U252 ( .B1(n404), .B2(n567), .A(n559), .ZN(n428) );
  NAND2_X1 U253 ( .A1(\mem[13][7] ), .A2(n567), .ZN(n559) );
  OAI21_X1 U254 ( .B1(n411), .B2(n558), .A(n557), .ZN(n427) );
  NAND2_X1 U255 ( .A1(\mem[14][0] ), .A2(n558), .ZN(n557) );
  OAI21_X1 U256 ( .B1(n410), .B2(n558), .A(n556), .ZN(n426) );
  NAND2_X1 U257 ( .A1(\mem[14][1] ), .A2(n558), .ZN(n556) );
  OAI21_X1 U258 ( .B1(n409), .B2(n558), .A(n555), .ZN(n425) );
  NAND2_X1 U259 ( .A1(\mem[14][2] ), .A2(n558), .ZN(n555) );
  OAI21_X1 U260 ( .B1(n408), .B2(n558), .A(n554), .ZN(n424) );
  NAND2_X1 U261 ( .A1(\mem[14][3] ), .A2(n558), .ZN(n554) );
  OAI21_X1 U262 ( .B1(n407), .B2(n558), .A(n553), .ZN(n423) );
  NAND2_X1 U263 ( .A1(\mem[14][4] ), .A2(n558), .ZN(n553) );
  OAI21_X1 U264 ( .B1(n406), .B2(n558), .A(n552), .ZN(n422) );
  NAND2_X1 U265 ( .A1(\mem[14][5] ), .A2(n558), .ZN(n552) );
  OAI21_X1 U266 ( .B1(n405), .B2(n558), .A(n551), .ZN(n421) );
  NAND2_X1 U267 ( .A1(\mem[14][6] ), .A2(n558), .ZN(n551) );
  OAI21_X1 U268 ( .B1(n404), .B2(n558), .A(n550), .ZN(n420) );
  NAND2_X1 U269 ( .A1(\mem[14][7] ), .A2(n558), .ZN(n550) );
  OAI21_X1 U270 ( .B1(n411), .B2(n548), .A(n547), .ZN(n419) );
  NAND2_X1 U271 ( .A1(\mem[15][0] ), .A2(n548), .ZN(n547) );
  OAI21_X1 U272 ( .B1(n410), .B2(n548), .A(n546), .ZN(n418) );
  NAND2_X1 U273 ( .A1(\mem[15][1] ), .A2(n548), .ZN(n546) );
  OAI21_X1 U274 ( .B1(n409), .B2(n548), .A(n545), .ZN(n417) );
  NAND2_X1 U275 ( .A1(\mem[15][2] ), .A2(n548), .ZN(n545) );
  OAI21_X1 U276 ( .B1(n408), .B2(n548), .A(n544), .ZN(n416) );
  NAND2_X1 U277 ( .A1(\mem[15][3] ), .A2(n548), .ZN(n544) );
  OAI21_X1 U278 ( .B1(n407), .B2(n548), .A(n543), .ZN(n415) );
  NAND2_X1 U279 ( .A1(\mem[15][4] ), .A2(n548), .ZN(n543) );
  OAI21_X1 U280 ( .B1(n406), .B2(n548), .A(n542), .ZN(n414) );
  NAND2_X1 U281 ( .A1(\mem[15][5] ), .A2(n548), .ZN(n542) );
  OAI21_X1 U282 ( .B1(n405), .B2(n548), .A(n541), .ZN(n413) );
  NAND2_X1 U283 ( .A1(\mem[15][6] ), .A2(n548), .ZN(n541) );
  OAI21_X1 U284 ( .B1(n404), .B2(n548), .A(n540), .ZN(n412) );
  NAND2_X1 U285 ( .A1(\mem[15][7] ), .A2(n548), .ZN(n540) );
  AND2_X1 U286 ( .A1(N13), .A2(wr_en), .ZN(n549) );
  NOR2_X1 U287 ( .A1(N11), .A2(N12), .ZN(n684) );
  NOR2_X1 U288 ( .A1(n402), .A2(N12), .ZN(n663) );
  AND2_X1 U289 ( .A1(N12), .A2(n402), .ZN(n644) );
  AND2_X1 U290 ( .A1(N12), .A2(N11), .ZN(n625) );
  INV_X1 U291 ( .A(data_in[0]), .ZN(n411) );
  INV_X1 U292 ( .A(data_in[1]), .ZN(n410) );
  INV_X1 U293 ( .A(data_in[2]), .ZN(n409) );
  INV_X1 U294 ( .A(data_in[3]), .ZN(n408) );
  INV_X1 U295 ( .A(data_in[4]), .ZN(n407) );
  INV_X1 U296 ( .A(data_in[5]), .ZN(n406) );
  INV_X1 U297 ( .A(data_in[6]), .ZN(n405) );
  INV_X1 U298 ( .A(data_in[7]), .ZN(n404) );
  MUX2_X1 U299 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n398), .Z(n3) );
  MUX2_X1 U300 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(N10), .Z(n4) );
  MUX2_X1 U301 ( .A(n4), .B(n3), .S(N11), .Z(n5) );
  MUX2_X1 U302 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(N10), .Z(n6) );
  MUX2_X1 U303 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n7) );
  MUX2_X1 U304 ( .A(n7), .B(n6), .S(N11), .Z(n8) );
  MUX2_X1 U305 ( .A(n8), .B(n5), .S(N12), .Z(n9) );
  MUX2_X1 U306 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n398), .Z(n10) );
  MUX2_X1 U307 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n398), .Z(n11) );
  MUX2_X1 U308 ( .A(n11), .B(n10), .S(N11), .Z(n294) );
  MUX2_X1 U309 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n398), .Z(n295) );
  MUX2_X1 U310 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n398), .Z(n296) );
  MUX2_X1 U311 ( .A(n296), .B(n295), .S(N11), .Z(n297) );
  MUX2_X1 U312 ( .A(n297), .B(n294), .S(N12), .Z(n298) );
  MUX2_X1 U313 ( .A(n298), .B(n9), .S(N13), .Z(N21) );
  MUX2_X1 U314 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n398), .Z(n299) );
  MUX2_X1 U315 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n398), .Z(n300) );
  MUX2_X1 U316 ( .A(n300), .B(n299), .S(N11), .Z(n301) );
  MUX2_X1 U317 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n398), .Z(n302) );
  MUX2_X1 U318 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n398), .Z(n303) );
  MUX2_X1 U319 ( .A(n303), .B(n302), .S(N11), .Z(n304) );
  MUX2_X1 U320 ( .A(n304), .B(n301), .S(N12), .Z(n305) );
  MUX2_X1 U321 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n398), .Z(n306) );
  MUX2_X1 U322 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n398), .Z(n307) );
  MUX2_X1 U323 ( .A(n307), .B(n306), .S(N11), .Z(n308) );
  MUX2_X1 U324 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n398), .Z(n309) );
  MUX2_X1 U325 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n398), .Z(n310) );
  MUX2_X1 U326 ( .A(n310), .B(n309), .S(N11), .Z(n311) );
  MUX2_X1 U327 ( .A(n311), .B(n308), .S(N12), .Z(n312) );
  MUX2_X1 U328 ( .A(n312), .B(n305), .S(N13), .Z(N20) );
  MUX2_X1 U329 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n399), .Z(n313) );
  MUX2_X1 U330 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n399), .Z(n314) );
  MUX2_X1 U331 ( .A(n314), .B(n313), .S(n397), .Z(n315) );
  MUX2_X1 U332 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n399), .Z(n316) );
  MUX2_X1 U333 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n399), .Z(n317) );
  MUX2_X1 U334 ( .A(n317), .B(n316), .S(n397), .Z(n318) );
  MUX2_X1 U335 ( .A(n318), .B(n315), .S(N12), .Z(n319) );
  MUX2_X1 U336 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n399), .Z(n320) );
  MUX2_X1 U337 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n399), .Z(n321) );
  MUX2_X1 U338 ( .A(n321), .B(n320), .S(n397), .Z(n322) );
  MUX2_X1 U339 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n399), .Z(n323) );
  MUX2_X1 U340 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n399), .Z(n324) );
  MUX2_X1 U341 ( .A(n324), .B(n323), .S(n397), .Z(n325) );
  MUX2_X1 U342 ( .A(n325), .B(n322), .S(N12), .Z(n326) );
  MUX2_X1 U343 ( .A(n326), .B(n319), .S(N13), .Z(N19) );
  MUX2_X1 U344 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n399), .Z(n327) );
  MUX2_X1 U345 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n399), .Z(n328) );
  MUX2_X1 U346 ( .A(n328), .B(n327), .S(n397), .Z(n329) );
  MUX2_X1 U347 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n399), .Z(n330) );
  MUX2_X1 U348 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n399), .Z(n331) );
  MUX2_X1 U349 ( .A(n331), .B(n330), .S(n397), .Z(n332) );
  MUX2_X1 U350 ( .A(n332), .B(n329), .S(N12), .Z(n333) );
  MUX2_X1 U351 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n400), .Z(n334) );
  MUX2_X1 U352 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n400), .Z(n335) );
  MUX2_X1 U353 ( .A(n335), .B(n334), .S(n397), .Z(n336) );
  MUX2_X1 U354 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n400), .Z(n337) );
  MUX2_X1 U355 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n400), .Z(n338) );
  MUX2_X1 U356 ( .A(n338), .B(n337), .S(n397), .Z(n339) );
  MUX2_X1 U357 ( .A(n339), .B(n336), .S(N12), .Z(n340) );
  MUX2_X1 U358 ( .A(n340), .B(n333), .S(N13), .Z(N18) );
  MUX2_X1 U359 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n400), .Z(n341) );
  MUX2_X1 U360 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n400), .Z(n342) );
  MUX2_X1 U361 ( .A(n342), .B(n341), .S(n397), .Z(n343) );
  MUX2_X1 U362 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n400), .Z(n344) );
  MUX2_X1 U363 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n400), .Z(n345) );
  MUX2_X1 U364 ( .A(n345), .B(n344), .S(n397), .Z(n346) );
  MUX2_X1 U365 ( .A(n346), .B(n343), .S(N12), .Z(n347) );
  MUX2_X1 U366 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n400), .Z(n348) );
  MUX2_X1 U367 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n400), .Z(n349) );
  MUX2_X1 U368 ( .A(n349), .B(n348), .S(n397), .Z(n350) );
  MUX2_X1 U369 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n400), .Z(n351) );
  MUX2_X1 U370 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n400), .Z(n352) );
  MUX2_X1 U371 ( .A(n352), .B(n351), .S(n397), .Z(n353) );
  MUX2_X1 U372 ( .A(n353), .B(n350), .S(N12), .Z(n354) );
  MUX2_X1 U373 ( .A(n354), .B(n347), .S(N13), .Z(N17) );
  MUX2_X1 U374 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n398), .Z(n355) );
  MUX2_X1 U375 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n399), .Z(n356) );
  MUX2_X1 U376 ( .A(n356), .B(n355), .S(N11), .Z(n357) );
  MUX2_X1 U377 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(N10), .Z(n358) );
  MUX2_X1 U378 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n399), .Z(n359) );
  MUX2_X1 U379 ( .A(n359), .B(n358), .S(N11), .Z(n360) );
  MUX2_X1 U380 ( .A(n360), .B(n357), .S(N12), .Z(n361) );
  MUX2_X1 U381 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n400), .Z(n362) );
  MUX2_X1 U382 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n400), .Z(n363) );
  MUX2_X1 U383 ( .A(n363), .B(n362), .S(N11), .Z(n364) );
  MUX2_X1 U384 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n400), .Z(n365) );
  MUX2_X1 U385 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n399), .Z(n366) );
  MUX2_X1 U386 ( .A(n366), .B(n365), .S(N11), .Z(n367) );
  MUX2_X1 U387 ( .A(n367), .B(n364), .S(N12), .Z(n368) );
  MUX2_X1 U388 ( .A(n368), .B(n361), .S(N13), .Z(N16) );
  MUX2_X1 U389 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(N10), .Z(n369) );
  MUX2_X1 U390 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n398), .Z(n370) );
  MUX2_X1 U391 ( .A(n370), .B(n369), .S(N11), .Z(n371) );
  MUX2_X1 U392 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(N10), .Z(n372) );
  MUX2_X1 U393 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n398), .Z(n373) );
  MUX2_X1 U394 ( .A(n373), .B(n372), .S(N11), .Z(n374) );
  MUX2_X1 U395 ( .A(n374), .B(n371), .S(N12), .Z(n375) );
  MUX2_X1 U396 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n376) );
  MUX2_X1 U397 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n377) );
  MUX2_X1 U398 ( .A(n377), .B(n376), .S(N11), .Z(n378) );
  MUX2_X1 U399 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n379) );
  MUX2_X1 U400 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n380) );
  MUX2_X1 U401 ( .A(n380), .B(n379), .S(n397), .Z(n381) );
  MUX2_X1 U402 ( .A(n381), .B(n378), .S(N12), .Z(n382) );
  MUX2_X1 U403 ( .A(n382), .B(n375), .S(N13), .Z(N15) );
  MUX2_X1 U404 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n400), .Z(n383) );
  MUX2_X1 U405 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n384) );
  MUX2_X1 U406 ( .A(n384), .B(n383), .S(N11), .Z(n385) );
  MUX2_X1 U407 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n399), .Z(n386) );
  MUX2_X1 U408 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n387) );
  MUX2_X1 U409 ( .A(n387), .B(n386), .S(N11), .Z(n388) );
  MUX2_X1 U410 ( .A(n388), .B(n385), .S(N12), .Z(n389) );
  MUX2_X1 U411 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n390) );
  MUX2_X1 U412 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n391) );
  MUX2_X1 U413 ( .A(n391), .B(n390), .S(N11), .Z(n392) );
  MUX2_X1 U414 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n393) );
  MUX2_X1 U415 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n394) );
  MUX2_X1 U416 ( .A(n394), .B(n393), .S(n397), .Z(n395) );
  MUX2_X1 U417 ( .A(n395), .B(n392), .S(N12), .Z(n396) );
  MUX2_X1 U418 ( .A(n396), .B(n389), .S(N13), .Z(N14) );
  INV_X1 U419 ( .A(N10), .ZN(n401) );
  INV_X1 U420 ( .A(N11), .ZN(n402) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_3 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, N19, N20, N21, n1, n3, n5, n7, n8, n9, n10, n11,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n416), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n417), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n418), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n419), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n420), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n421), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n422), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n423), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n424), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n425), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n426), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n427), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n428), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n429), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n430), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n431), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n432), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n433), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n434), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n435), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n436), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n437), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n438), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n439), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n440), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n441), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n442), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n443), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n444), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n445), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n446), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n447), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n448), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n449), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n450), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n451), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n452), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n453), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n454), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n455), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n456), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n457), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n458), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n459), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n460), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n461), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n462), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n463), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n464), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n465), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n466), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n467), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n468), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n469), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n470), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n471), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n472), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n473), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n474), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n475), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n476), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n477), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n478), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n479), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n480), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n481), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n482), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n483), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n484), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n485), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n486), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n487), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n488), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n489), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n490), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n491), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n492), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n493), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n494), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n495), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n496), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n497), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n498), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n499), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n500), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n501), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n502), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n503), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n504), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n505), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n506), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n507), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n508), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n509), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n510), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n511), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n512), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n513), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n514), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n515), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n516), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n517), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n518), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n519), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n520), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n521), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n522), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n523), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n524), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n525), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n526), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n527), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n528), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n529), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n530), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n531), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n532), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n533), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n534), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n535), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n536), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n537), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n538), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n539), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n540), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n541), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n542), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n543), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N20), .CK(clk), .QN(n5) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .QN(n3) );
  DFF_X1 \data_out_reg[5]  ( .D(N16), .CK(clk), .QN(n1) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[5]) );
  INV_X2 U4 ( .A(n3), .ZN(data_out[3]) );
  INV_X2 U5 ( .A(n5), .ZN(data_out[1]) );
  BUF_X1 U6 ( .A(N10), .Z(n402) );
  BUF_X1 U7 ( .A(N10), .Z(n403) );
  BUF_X1 U8 ( .A(N10), .Z(n404) );
  BUF_X1 U9 ( .A(N11), .Z(n401) );
  NAND2_X1 U10 ( .A1(n667), .A2(n687), .ZN(n676) );
  NAND2_X1 U11 ( .A1(n667), .A2(n677), .ZN(n666) );
  NAND2_X1 U12 ( .A1(n688), .A2(n687), .ZN(n697) );
  NAND2_X1 U13 ( .A1(n677), .A2(n688), .ZN(n686) );
  NAND2_X1 U14 ( .A1(n609), .A2(n688), .ZN(n618) );
  NAND2_X1 U15 ( .A1(n599), .A2(n688), .ZN(n608) );
  NAND2_X1 U16 ( .A1(n609), .A2(n667), .ZN(n598) );
  NAND2_X1 U17 ( .A1(n599), .A2(n667), .ZN(n589) );
  NAND2_X1 U18 ( .A1(n648), .A2(n687), .ZN(n657) );
  NAND2_X1 U19 ( .A1(n648), .A2(n677), .ZN(n647) );
  NAND2_X1 U20 ( .A1(n629), .A2(n687), .ZN(n638) );
  NAND2_X1 U21 ( .A1(n629), .A2(n677), .ZN(n627) );
  NAND2_X1 U22 ( .A1(n609), .A2(n648), .ZN(n580) );
  NAND2_X1 U23 ( .A1(n599), .A2(n648), .ZN(n571) );
  NAND2_X1 U24 ( .A1(n609), .A2(n629), .ZN(n562) );
  NAND2_X1 U25 ( .A1(n599), .A2(n629), .ZN(n552) );
  AND2_X1 U26 ( .A1(n553), .A2(N10), .ZN(n599) );
  AND2_X1 U27 ( .A1(n553), .A2(n405), .ZN(n609) );
  AND2_X1 U28 ( .A1(N10), .A2(n628), .ZN(n677) );
  AND2_X1 U29 ( .A1(n628), .A2(n405), .ZN(n687) );
  OAI21_X1 U30 ( .B1(n697), .B2(n415), .A(n696), .ZN(n543) );
  NAND2_X1 U31 ( .A1(\mem[0][0] ), .A2(n697), .ZN(n696) );
  OAI21_X1 U32 ( .B1(n697), .B2(n414), .A(n695), .ZN(n542) );
  NAND2_X1 U33 ( .A1(\mem[0][1] ), .A2(n697), .ZN(n695) );
  OAI21_X1 U34 ( .B1(n697), .B2(n413), .A(n694), .ZN(n541) );
  NAND2_X1 U35 ( .A1(\mem[0][2] ), .A2(n697), .ZN(n694) );
  OAI21_X1 U36 ( .B1(n697), .B2(n412), .A(n693), .ZN(n540) );
  NAND2_X1 U37 ( .A1(\mem[0][3] ), .A2(n697), .ZN(n693) );
  OAI21_X1 U38 ( .B1(n697), .B2(n411), .A(n692), .ZN(n539) );
  NAND2_X1 U39 ( .A1(\mem[0][4] ), .A2(n697), .ZN(n692) );
  OAI21_X1 U40 ( .B1(n697), .B2(n410), .A(n691), .ZN(n538) );
  NAND2_X1 U41 ( .A1(\mem[0][5] ), .A2(n697), .ZN(n691) );
  OAI21_X1 U42 ( .B1(n697), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U43 ( .A1(\mem[0][6] ), .A2(n697), .ZN(n690) );
  OAI21_X1 U44 ( .B1(n697), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U45 ( .A1(\mem[0][7] ), .A2(n697), .ZN(n689) );
  OAI21_X1 U46 ( .B1(n415), .B2(n676), .A(n675), .ZN(n527) );
  NAND2_X1 U47 ( .A1(\mem[2][0] ), .A2(n676), .ZN(n675) );
  OAI21_X1 U48 ( .B1(n414), .B2(n676), .A(n674), .ZN(n526) );
  NAND2_X1 U49 ( .A1(\mem[2][1] ), .A2(n676), .ZN(n674) );
  OAI21_X1 U50 ( .B1(n413), .B2(n676), .A(n673), .ZN(n525) );
  NAND2_X1 U51 ( .A1(\mem[2][2] ), .A2(n676), .ZN(n673) );
  OAI21_X1 U52 ( .B1(n412), .B2(n676), .A(n672), .ZN(n524) );
  NAND2_X1 U53 ( .A1(\mem[2][3] ), .A2(n676), .ZN(n672) );
  OAI21_X1 U54 ( .B1(n411), .B2(n676), .A(n671), .ZN(n523) );
  NAND2_X1 U55 ( .A1(\mem[2][4] ), .A2(n676), .ZN(n671) );
  OAI21_X1 U56 ( .B1(n410), .B2(n676), .A(n670), .ZN(n522) );
  NAND2_X1 U57 ( .A1(\mem[2][5] ), .A2(n676), .ZN(n670) );
  OAI21_X1 U58 ( .B1(n409), .B2(n676), .A(n669), .ZN(n521) );
  NAND2_X1 U59 ( .A1(\mem[2][6] ), .A2(n676), .ZN(n669) );
  OAI21_X1 U60 ( .B1(n408), .B2(n676), .A(n668), .ZN(n520) );
  NAND2_X1 U61 ( .A1(\mem[2][7] ), .A2(n676), .ZN(n668) );
  OAI21_X1 U62 ( .B1(n415), .B2(n666), .A(n665), .ZN(n519) );
  NAND2_X1 U63 ( .A1(\mem[3][0] ), .A2(n666), .ZN(n665) );
  OAI21_X1 U64 ( .B1(n414), .B2(n666), .A(n664), .ZN(n518) );
  NAND2_X1 U65 ( .A1(\mem[3][1] ), .A2(n666), .ZN(n664) );
  OAI21_X1 U66 ( .B1(n413), .B2(n666), .A(n663), .ZN(n517) );
  NAND2_X1 U67 ( .A1(\mem[3][2] ), .A2(n666), .ZN(n663) );
  OAI21_X1 U68 ( .B1(n412), .B2(n666), .A(n662), .ZN(n516) );
  NAND2_X1 U69 ( .A1(\mem[3][3] ), .A2(n666), .ZN(n662) );
  OAI21_X1 U70 ( .B1(n411), .B2(n666), .A(n661), .ZN(n515) );
  NAND2_X1 U71 ( .A1(\mem[3][4] ), .A2(n666), .ZN(n661) );
  OAI21_X1 U72 ( .B1(n410), .B2(n666), .A(n660), .ZN(n514) );
  NAND2_X1 U73 ( .A1(\mem[3][5] ), .A2(n666), .ZN(n660) );
  OAI21_X1 U74 ( .B1(n409), .B2(n666), .A(n659), .ZN(n513) );
  NAND2_X1 U75 ( .A1(\mem[3][6] ), .A2(n666), .ZN(n659) );
  OAI21_X1 U76 ( .B1(n408), .B2(n666), .A(n658), .ZN(n512) );
  NAND2_X1 U77 ( .A1(\mem[3][7] ), .A2(n666), .ZN(n658) );
  NOR2_X1 U78 ( .A1(n407), .A2(N13), .ZN(n628) );
  INV_X1 U79 ( .A(wr_en), .ZN(n407) );
  OAI21_X1 U80 ( .B1(n415), .B2(n686), .A(n685), .ZN(n535) );
  NAND2_X1 U81 ( .A1(\mem[1][0] ), .A2(n686), .ZN(n685) );
  OAI21_X1 U82 ( .B1(n414), .B2(n686), .A(n684), .ZN(n534) );
  NAND2_X1 U83 ( .A1(\mem[1][1] ), .A2(n686), .ZN(n684) );
  OAI21_X1 U84 ( .B1(n413), .B2(n686), .A(n683), .ZN(n533) );
  NAND2_X1 U85 ( .A1(\mem[1][2] ), .A2(n686), .ZN(n683) );
  OAI21_X1 U86 ( .B1(n412), .B2(n686), .A(n682), .ZN(n532) );
  NAND2_X1 U87 ( .A1(\mem[1][3] ), .A2(n686), .ZN(n682) );
  OAI21_X1 U88 ( .B1(n411), .B2(n686), .A(n681), .ZN(n531) );
  NAND2_X1 U89 ( .A1(\mem[1][4] ), .A2(n686), .ZN(n681) );
  OAI21_X1 U90 ( .B1(n410), .B2(n686), .A(n680), .ZN(n530) );
  NAND2_X1 U91 ( .A1(\mem[1][5] ), .A2(n686), .ZN(n680) );
  OAI21_X1 U92 ( .B1(n409), .B2(n686), .A(n679), .ZN(n529) );
  NAND2_X1 U93 ( .A1(\mem[1][6] ), .A2(n686), .ZN(n679) );
  OAI21_X1 U94 ( .B1(n408), .B2(n686), .A(n678), .ZN(n528) );
  NAND2_X1 U95 ( .A1(\mem[1][7] ), .A2(n686), .ZN(n678) );
  OAI21_X1 U96 ( .B1(n415), .B2(n657), .A(n656), .ZN(n511) );
  NAND2_X1 U97 ( .A1(\mem[4][0] ), .A2(n657), .ZN(n656) );
  OAI21_X1 U98 ( .B1(n414), .B2(n657), .A(n655), .ZN(n510) );
  NAND2_X1 U99 ( .A1(\mem[4][1] ), .A2(n657), .ZN(n655) );
  OAI21_X1 U100 ( .B1(n413), .B2(n657), .A(n654), .ZN(n509) );
  NAND2_X1 U101 ( .A1(\mem[4][2] ), .A2(n657), .ZN(n654) );
  OAI21_X1 U102 ( .B1(n412), .B2(n657), .A(n653), .ZN(n508) );
  NAND2_X1 U103 ( .A1(\mem[4][3] ), .A2(n657), .ZN(n653) );
  OAI21_X1 U104 ( .B1(n411), .B2(n657), .A(n652), .ZN(n507) );
  NAND2_X1 U105 ( .A1(\mem[4][4] ), .A2(n657), .ZN(n652) );
  OAI21_X1 U106 ( .B1(n410), .B2(n657), .A(n651), .ZN(n506) );
  NAND2_X1 U107 ( .A1(\mem[4][5] ), .A2(n657), .ZN(n651) );
  OAI21_X1 U108 ( .B1(n409), .B2(n657), .A(n650), .ZN(n505) );
  NAND2_X1 U109 ( .A1(\mem[4][6] ), .A2(n657), .ZN(n650) );
  OAI21_X1 U110 ( .B1(n408), .B2(n657), .A(n649), .ZN(n504) );
  NAND2_X1 U111 ( .A1(\mem[4][7] ), .A2(n657), .ZN(n649) );
  OAI21_X1 U112 ( .B1(n415), .B2(n647), .A(n646), .ZN(n503) );
  NAND2_X1 U113 ( .A1(\mem[5][0] ), .A2(n647), .ZN(n646) );
  OAI21_X1 U114 ( .B1(n414), .B2(n647), .A(n645), .ZN(n502) );
  NAND2_X1 U115 ( .A1(\mem[5][1] ), .A2(n647), .ZN(n645) );
  OAI21_X1 U116 ( .B1(n413), .B2(n647), .A(n644), .ZN(n501) );
  NAND2_X1 U117 ( .A1(\mem[5][2] ), .A2(n647), .ZN(n644) );
  OAI21_X1 U118 ( .B1(n412), .B2(n647), .A(n643), .ZN(n500) );
  NAND2_X1 U119 ( .A1(\mem[5][3] ), .A2(n647), .ZN(n643) );
  OAI21_X1 U120 ( .B1(n411), .B2(n647), .A(n642), .ZN(n499) );
  NAND2_X1 U121 ( .A1(\mem[5][4] ), .A2(n647), .ZN(n642) );
  OAI21_X1 U122 ( .B1(n410), .B2(n647), .A(n641), .ZN(n498) );
  NAND2_X1 U123 ( .A1(\mem[5][5] ), .A2(n647), .ZN(n641) );
  OAI21_X1 U124 ( .B1(n409), .B2(n647), .A(n640), .ZN(n497) );
  NAND2_X1 U125 ( .A1(\mem[5][6] ), .A2(n647), .ZN(n640) );
  OAI21_X1 U126 ( .B1(n408), .B2(n647), .A(n639), .ZN(n496) );
  NAND2_X1 U127 ( .A1(\mem[5][7] ), .A2(n647), .ZN(n639) );
  OAI21_X1 U128 ( .B1(n415), .B2(n638), .A(n637), .ZN(n495) );
  NAND2_X1 U129 ( .A1(\mem[6][0] ), .A2(n638), .ZN(n637) );
  OAI21_X1 U130 ( .B1(n414), .B2(n638), .A(n636), .ZN(n494) );
  NAND2_X1 U131 ( .A1(\mem[6][1] ), .A2(n638), .ZN(n636) );
  OAI21_X1 U132 ( .B1(n413), .B2(n638), .A(n635), .ZN(n493) );
  NAND2_X1 U133 ( .A1(\mem[6][2] ), .A2(n638), .ZN(n635) );
  OAI21_X1 U134 ( .B1(n412), .B2(n638), .A(n634), .ZN(n492) );
  NAND2_X1 U135 ( .A1(\mem[6][3] ), .A2(n638), .ZN(n634) );
  OAI21_X1 U136 ( .B1(n411), .B2(n638), .A(n633), .ZN(n491) );
  NAND2_X1 U137 ( .A1(\mem[6][4] ), .A2(n638), .ZN(n633) );
  OAI21_X1 U138 ( .B1(n410), .B2(n638), .A(n632), .ZN(n490) );
  NAND2_X1 U139 ( .A1(\mem[6][5] ), .A2(n638), .ZN(n632) );
  OAI21_X1 U140 ( .B1(n409), .B2(n638), .A(n631), .ZN(n489) );
  NAND2_X1 U141 ( .A1(\mem[6][6] ), .A2(n638), .ZN(n631) );
  OAI21_X1 U142 ( .B1(n408), .B2(n638), .A(n630), .ZN(n488) );
  NAND2_X1 U143 ( .A1(\mem[6][7] ), .A2(n638), .ZN(n630) );
  OAI21_X1 U144 ( .B1(n415), .B2(n627), .A(n626), .ZN(n487) );
  NAND2_X1 U145 ( .A1(\mem[7][0] ), .A2(n627), .ZN(n626) );
  OAI21_X1 U146 ( .B1(n414), .B2(n627), .A(n625), .ZN(n486) );
  NAND2_X1 U147 ( .A1(\mem[7][1] ), .A2(n627), .ZN(n625) );
  OAI21_X1 U148 ( .B1(n413), .B2(n627), .A(n624), .ZN(n485) );
  NAND2_X1 U149 ( .A1(\mem[7][2] ), .A2(n627), .ZN(n624) );
  OAI21_X1 U150 ( .B1(n412), .B2(n627), .A(n623), .ZN(n484) );
  NAND2_X1 U151 ( .A1(\mem[7][3] ), .A2(n627), .ZN(n623) );
  OAI21_X1 U152 ( .B1(n411), .B2(n627), .A(n622), .ZN(n483) );
  NAND2_X1 U153 ( .A1(\mem[7][4] ), .A2(n627), .ZN(n622) );
  OAI21_X1 U154 ( .B1(n410), .B2(n627), .A(n621), .ZN(n482) );
  NAND2_X1 U155 ( .A1(\mem[7][5] ), .A2(n627), .ZN(n621) );
  OAI21_X1 U156 ( .B1(n409), .B2(n627), .A(n620), .ZN(n481) );
  NAND2_X1 U157 ( .A1(\mem[7][6] ), .A2(n627), .ZN(n620) );
  OAI21_X1 U158 ( .B1(n408), .B2(n627), .A(n619), .ZN(n480) );
  NAND2_X1 U159 ( .A1(\mem[7][7] ), .A2(n627), .ZN(n619) );
  OAI21_X1 U160 ( .B1(n415), .B2(n618), .A(n617), .ZN(n479) );
  NAND2_X1 U161 ( .A1(\mem[8][0] ), .A2(n618), .ZN(n617) );
  OAI21_X1 U162 ( .B1(n414), .B2(n618), .A(n616), .ZN(n478) );
  NAND2_X1 U163 ( .A1(\mem[8][1] ), .A2(n618), .ZN(n616) );
  OAI21_X1 U164 ( .B1(n413), .B2(n618), .A(n615), .ZN(n477) );
  NAND2_X1 U165 ( .A1(\mem[8][2] ), .A2(n618), .ZN(n615) );
  OAI21_X1 U166 ( .B1(n412), .B2(n618), .A(n614), .ZN(n476) );
  NAND2_X1 U167 ( .A1(\mem[8][3] ), .A2(n618), .ZN(n614) );
  OAI21_X1 U168 ( .B1(n411), .B2(n618), .A(n613), .ZN(n475) );
  NAND2_X1 U169 ( .A1(\mem[8][4] ), .A2(n618), .ZN(n613) );
  OAI21_X1 U170 ( .B1(n410), .B2(n618), .A(n612), .ZN(n474) );
  NAND2_X1 U171 ( .A1(\mem[8][5] ), .A2(n618), .ZN(n612) );
  OAI21_X1 U172 ( .B1(n409), .B2(n618), .A(n611), .ZN(n473) );
  NAND2_X1 U173 ( .A1(\mem[8][6] ), .A2(n618), .ZN(n611) );
  OAI21_X1 U174 ( .B1(n408), .B2(n618), .A(n610), .ZN(n472) );
  NAND2_X1 U175 ( .A1(\mem[8][7] ), .A2(n618), .ZN(n610) );
  OAI21_X1 U176 ( .B1(n415), .B2(n608), .A(n607), .ZN(n471) );
  NAND2_X1 U177 ( .A1(\mem[9][0] ), .A2(n608), .ZN(n607) );
  OAI21_X1 U178 ( .B1(n414), .B2(n608), .A(n606), .ZN(n470) );
  NAND2_X1 U179 ( .A1(\mem[9][1] ), .A2(n608), .ZN(n606) );
  OAI21_X1 U180 ( .B1(n413), .B2(n608), .A(n605), .ZN(n469) );
  NAND2_X1 U181 ( .A1(\mem[9][2] ), .A2(n608), .ZN(n605) );
  OAI21_X1 U182 ( .B1(n412), .B2(n608), .A(n604), .ZN(n468) );
  NAND2_X1 U183 ( .A1(\mem[9][3] ), .A2(n608), .ZN(n604) );
  OAI21_X1 U184 ( .B1(n411), .B2(n608), .A(n603), .ZN(n467) );
  NAND2_X1 U185 ( .A1(\mem[9][4] ), .A2(n608), .ZN(n603) );
  OAI21_X1 U186 ( .B1(n410), .B2(n608), .A(n602), .ZN(n466) );
  NAND2_X1 U187 ( .A1(\mem[9][5] ), .A2(n608), .ZN(n602) );
  OAI21_X1 U188 ( .B1(n409), .B2(n608), .A(n601), .ZN(n465) );
  NAND2_X1 U189 ( .A1(\mem[9][6] ), .A2(n608), .ZN(n601) );
  OAI21_X1 U190 ( .B1(n408), .B2(n608), .A(n600), .ZN(n464) );
  NAND2_X1 U191 ( .A1(\mem[9][7] ), .A2(n608), .ZN(n600) );
  OAI21_X1 U192 ( .B1(n415), .B2(n598), .A(n597), .ZN(n463) );
  NAND2_X1 U193 ( .A1(\mem[10][0] ), .A2(n598), .ZN(n597) );
  OAI21_X1 U194 ( .B1(n414), .B2(n598), .A(n596), .ZN(n462) );
  NAND2_X1 U195 ( .A1(\mem[10][1] ), .A2(n598), .ZN(n596) );
  OAI21_X1 U196 ( .B1(n413), .B2(n598), .A(n595), .ZN(n461) );
  NAND2_X1 U197 ( .A1(\mem[10][2] ), .A2(n598), .ZN(n595) );
  OAI21_X1 U198 ( .B1(n412), .B2(n598), .A(n594), .ZN(n460) );
  NAND2_X1 U199 ( .A1(\mem[10][3] ), .A2(n598), .ZN(n594) );
  OAI21_X1 U200 ( .B1(n411), .B2(n598), .A(n593), .ZN(n459) );
  NAND2_X1 U201 ( .A1(\mem[10][4] ), .A2(n598), .ZN(n593) );
  OAI21_X1 U202 ( .B1(n410), .B2(n598), .A(n592), .ZN(n458) );
  NAND2_X1 U203 ( .A1(\mem[10][5] ), .A2(n598), .ZN(n592) );
  OAI21_X1 U204 ( .B1(n409), .B2(n598), .A(n591), .ZN(n457) );
  NAND2_X1 U205 ( .A1(\mem[10][6] ), .A2(n598), .ZN(n591) );
  OAI21_X1 U206 ( .B1(n408), .B2(n598), .A(n590), .ZN(n456) );
  NAND2_X1 U207 ( .A1(\mem[10][7] ), .A2(n598), .ZN(n590) );
  OAI21_X1 U208 ( .B1(n415), .B2(n589), .A(n588), .ZN(n455) );
  NAND2_X1 U209 ( .A1(\mem[11][0] ), .A2(n589), .ZN(n588) );
  OAI21_X1 U210 ( .B1(n414), .B2(n589), .A(n587), .ZN(n454) );
  NAND2_X1 U211 ( .A1(\mem[11][1] ), .A2(n589), .ZN(n587) );
  OAI21_X1 U212 ( .B1(n413), .B2(n589), .A(n586), .ZN(n453) );
  NAND2_X1 U213 ( .A1(\mem[11][2] ), .A2(n589), .ZN(n586) );
  OAI21_X1 U214 ( .B1(n412), .B2(n589), .A(n585), .ZN(n452) );
  NAND2_X1 U215 ( .A1(\mem[11][3] ), .A2(n589), .ZN(n585) );
  OAI21_X1 U216 ( .B1(n411), .B2(n589), .A(n584), .ZN(n451) );
  NAND2_X1 U217 ( .A1(\mem[11][4] ), .A2(n589), .ZN(n584) );
  OAI21_X1 U218 ( .B1(n410), .B2(n589), .A(n583), .ZN(n450) );
  NAND2_X1 U219 ( .A1(\mem[11][5] ), .A2(n589), .ZN(n583) );
  OAI21_X1 U220 ( .B1(n409), .B2(n589), .A(n582), .ZN(n449) );
  NAND2_X1 U221 ( .A1(\mem[11][6] ), .A2(n589), .ZN(n582) );
  OAI21_X1 U222 ( .B1(n408), .B2(n589), .A(n581), .ZN(n448) );
  NAND2_X1 U223 ( .A1(\mem[11][7] ), .A2(n589), .ZN(n581) );
  OAI21_X1 U224 ( .B1(n415), .B2(n580), .A(n579), .ZN(n447) );
  NAND2_X1 U225 ( .A1(\mem[12][0] ), .A2(n580), .ZN(n579) );
  OAI21_X1 U226 ( .B1(n414), .B2(n580), .A(n578), .ZN(n446) );
  NAND2_X1 U227 ( .A1(\mem[12][1] ), .A2(n580), .ZN(n578) );
  OAI21_X1 U228 ( .B1(n413), .B2(n580), .A(n577), .ZN(n445) );
  NAND2_X1 U229 ( .A1(\mem[12][2] ), .A2(n580), .ZN(n577) );
  OAI21_X1 U230 ( .B1(n412), .B2(n580), .A(n576), .ZN(n444) );
  NAND2_X1 U231 ( .A1(\mem[12][3] ), .A2(n580), .ZN(n576) );
  OAI21_X1 U232 ( .B1(n411), .B2(n580), .A(n575), .ZN(n443) );
  NAND2_X1 U233 ( .A1(\mem[12][4] ), .A2(n580), .ZN(n575) );
  OAI21_X1 U234 ( .B1(n410), .B2(n580), .A(n574), .ZN(n442) );
  NAND2_X1 U235 ( .A1(\mem[12][5] ), .A2(n580), .ZN(n574) );
  OAI21_X1 U236 ( .B1(n409), .B2(n580), .A(n573), .ZN(n441) );
  NAND2_X1 U237 ( .A1(\mem[12][6] ), .A2(n580), .ZN(n573) );
  OAI21_X1 U238 ( .B1(n408), .B2(n580), .A(n572), .ZN(n440) );
  NAND2_X1 U239 ( .A1(\mem[12][7] ), .A2(n580), .ZN(n572) );
  OAI21_X1 U240 ( .B1(n415), .B2(n571), .A(n570), .ZN(n439) );
  NAND2_X1 U241 ( .A1(\mem[13][0] ), .A2(n571), .ZN(n570) );
  OAI21_X1 U242 ( .B1(n414), .B2(n571), .A(n569), .ZN(n438) );
  NAND2_X1 U243 ( .A1(\mem[13][1] ), .A2(n571), .ZN(n569) );
  OAI21_X1 U244 ( .B1(n413), .B2(n571), .A(n568), .ZN(n437) );
  NAND2_X1 U245 ( .A1(\mem[13][2] ), .A2(n571), .ZN(n568) );
  OAI21_X1 U246 ( .B1(n412), .B2(n571), .A(n567), .ZN(n436) );
  NAND2_X1 U247 ( .A1(\mem[13][3] ), .A2(n571), .ZN(n567) );
  OAI21_X1 U248 ( .B1(n411), .B2(n571), .A(n566), .ZN(n435) );
  NAND2_X1 U249 ( .A1(\mem[13][4] ), .A2(n571), .ZN(n566) );
  OAI21_X1 U250 ( .B1(n410), .B2(n571), .A(n565), .ZN(n434) );
  NAND2_X1 U251 ( .A1(\mem[13][5] ), .A2(n571), .ZN(n565) );
  OAI21_X1 U252 ( .B1(n409), .B2(n571), .A(n564), .ZN(n433) );
  NAND2_X1 U253 ( .A1(\mem[13][6] ), .A2(n571), .ZN(n564) );
  OAI21_X1 U254 ( .B1(n408), .B2(n571), .A(n563), .ZN(n432) );
  NAND2_X1 U255 ( .A1(\mem[13][7] ), .A2(n571), .ZN(n563) );
  OAI21_X1 U256 ( .B1(n415), .B2(n562), .A(n561), .ZN(n431) );
  NAND2_X1 U257 ( .A1(\mem[14][0] ), .A2(n562), .ZN(n561) );
  OAI21_X1 U258 ( .B1(n414), .B2(n562), .A(n560), .ZN(n430) );
  NAND2_X1 U259 ( .A1(\mem[14][1] ), .A2(n562), .ZN(n560) );
  OAI21_X1 U260 ( .B1(n413), .B2(n562), .A(n559), .ZN(n429) );
  NAND2_X1 U261 ( .A1(\mem[14][2] ), .A2(n562), .ZN(n559) );
  OAI21_X1 U262 ( .B1(n412), .B2(n562), .A(n558), .ZN(n428) );
  NAND2_X1 U263 ( .A1(\mem[14][3] ), .A2(n562), .ZN(n558) );
  OAI21_X1 U264 ( .B1(n411), .B2(n562), .A(n557), .ZN(n427) );
  NAND2_X1 U265 ( .A1(\mem[14][4] ), .A2(n562), .ZN(n557) );
  OAI21_X1 U266 ( .B1(n410), .B2(n562), .A(n556), .ZN(n426) );
  NAND2_X1 U267 ( .A1(\mem[14][5] ), .A2(n562), .ZN(n556) );
  OAI21_X1 U268 ( .B1(n409), .B2(n562), .A(n555), .ZN(n425) );
  NAND2_X1 U269 ( .A1(\mem[14][6] ), .A2(n562), .ZN(n555) );
  OAI21_X1 U270 ( .B1(n408), .B2(n562), .A(n554), .ZN(n424) );
  NAND2_X1 U271 ( .A1(\mem[14][7] ), .A2(n562), .ZN(n554) );
  OAI21_X1 U272 ( .B1(n415), .B2(n552), .A(n551), .ZN(n423) );
  NAND2_X1 U273 ( .A1(\mem[15][0] ), .A2(n552), .ZN(n551) );
  OAI21_X1 U274 ( .B1(n414), .B2(n552), .A(n550), .ZN(n422) );
  NAND2_X1 U275 ( .A1(\mem[15][1] ), .A2(n552), .ZN(n550) );
  OAI21_X1 U276 ( .B1(n413), .B2(n552), .A(n549), .ZN(n421) );
  NAND2_X1 U277 ( .A1(\mem[15][2] ), .A2(n552), .ZN(n549) );
  OAI21_X1 U278 ( .B1(n412), .B2(n552), .A(n548), .ZN(n420) );
  NAND2_X1 U279 ( .A1(\mem[15][3] ), .A2(n552), .ZN(n548) );
  OAI21_X1 U280 ( .B1(n411), .B2(n552), .A(n547), .ZN(n419) );
  NAND2_X1 U281 ( .A1(\mem[15][4] ), .A2(n552), .ZN(n547) );
  OAI21_X1 U282 ( .B1(n410), .B2(n552), .A(n546), .ZN(n418) );
  NAND2_X1 U283 ( .A1(\mem[15][5] ), .A2(n552), .ZN(n546) );
  OAI21_X1 U284 ( .B1(n409), .B2(n552), .A(n545), .ZN(n417) );
  NAND2_X1 U285 ( .A1(\mem[15][6] ), .A2(n552), .ZN(n545) );
  OAI21_X1 U286 ( .B1(n408), .B2(n552), .A(n544), .ZN(n416) );
  NAND2_X1 U287 ( .A1(\mem[15][7] ), .A2(n552), .ZN(n544) );
  AND2_X1 U288 ( .A1(N13), .A2(wr_en), .ZN(n553) );
  NOR2_X1 U289 ( .A1(N11), .A2(N12), .ZN(n688) );
  NOR2_X1 U290 ( .A1(n406), .A2(N12), .ZN(n667) );
  AND2_X1 U291 ( .A1(N12), .A2(n406), .ZN(n648) );
  AND2_X1 U292 ( .A1(N12), .A2(N11), .ZN(n629) );
  INV_X1 U293 ( .A(data_in[0]), .ZN(n415) );
  INV_X1 U294 ( .A(data_in[1]), .ZN(n414) );
  INV_X1 U295 ( .A(data_in[2]), .ZN(n413) );
  INV_X1 U296 ( .A(data_in[3]), .ZN(n412) );
  INV_X1 U297 ( .A(data_in[4]), .ZN(n411) );
  INV_X1 U298 ( .A(data_in[5]), .ZN(n410) );
  INV_X1 U299 ( .A(data_in[6]), .ZN(n409) );
  INV_X1 U300 ( .A(data_in[7]), .ZN(n408) );
  MUX2_X1 U301 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(N10), .Z(n7) );
  MUX2_X1 U302 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(N10), .Z(n8) );
  MUX2_X1 U303 ( .A(n8), .B(n7), .S(n401), .Z(n9) );
  MUX2_X1 U304 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(N10), .Z(n10) );
  MUX2_X1 U305 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n11) );
  MUX2_X1 U306 ( .A(n11), .B(n10), .S(n401), .Z(n294) );
  MUX2_X1 U307 ( .A(n294), .B(n9), .S(N12), .Z(n295) );
  MUX2_X1 U308 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n402), .Z(n296) );
  MUX2_X1 U309 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n402), .Z(n297) );
  MUX2_X1 U310 ( .A(n297), .B(n296), .S(n401), .Z(n298) );
  MUX2_X1 U311 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n402), .Z(n299) );
  MUX2_X1 U312 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n402), .Z(n300) );
  MUX2_X1 U313 ( .A(n300), .B(n299), .S(n401), .Z(n301) );
  MUX2_X1 U314 ( .A(n301), .B(n298), .S(N12), .Z(n302) );
  MUX2_X1 U315 ( .A(n302), .B(n295), .S(N13), .Z(N21) );
  MUX2_X1 U316 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n402), .Z(n303) );
  MUX2_X1 U317 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n402), .Z(n304) );
  MUX2_X1 U318 ( .A(n304), .B(n303), .S(n401), .Z(n305) );
  MUX2_X1 U319 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n402), .Z(n306) );
  MUX2_X1 U320 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n402), .Z(n307) );
  MUX2_X1 U321 ( .A(n307), .B(n306), .S(n401), .Z(n308) );
  MUX2_X1 U322 ( .A(n308), .B(n305), .S(N12), .Z(n309) );
  MUX2_X1 U323 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n402), .Z(n310) );
  MUX2_X1 U324 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n402), .Z(n311) );
  MUX2_X1 U325 ( .A(n311), .B(n310), .S(n401), .Z(n312) );
  MUX2_X1 U326 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n402), .Z(n313) );
  MUX2_X1 U327 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n402), .Z(n314) );
  MUX2_X1 U328 ( .A(n314), .B(n313), .S(n401), .Z(n315) );
  MUX2_X1 U329 ( .A(n315), .B(n312), .S(N12), .Z(n316) );
  MUX2_X1 U330 ( .A(n316), .B(n309), .S(N13), .Z(N20) );
  MUX2_X1 U331 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n403), .Z(n317) );
  MUX2_X1 U332 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n403), .Z(n318) );
  MUX2_X1 U333 ( .A(n318), .B(n317), .S(N11), .Z(n319) );
  MUX2_X1 U334 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n403), .Z(n320) );
  MUX2_X1 U335 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n403), .Z(n321) );
  MUX2_X1 U336 ( .A(n321), .B(n320), .S(N11), .Z(n322) );
  MUX2_X1 U337 ( .A(n322), .B(n319), .S(N12), .Z(n323) );
  MUX2_X1 U338 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n403), .Z(n324) );
  MUX2_X1 U339 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n403), .Z(n325) );
  MUX2_X1 U340 ( .A(n325), .B(n324), .S(N11), .Z(n326) );
  MUX2_X1 U341 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n403), .Z(n327) );
  MUX2_X1 U342 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n403), .Z(n328) );
  MUX2_X1 U343 ( .A(n328), .B(n327), .S(n401), .Z(n329) );
  MUX2_X1 U344 ( .A(n329), .B(n326), .S(N12), .Z(n330) );
  MUX2_X1 U345 ( .A(n330), .B(n323), .S(N13), .Z(N19) );
  MUX2_X1 U346 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n403), .Z(n331) );
  MUX2_X1 U347 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n403), .Z(n332) );
  MUX2_X1 U348 ( .A(n332), .B(n331), .S(N11), .Z(n333) );
  MUX2_X1 U349 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n403), .Z(n334) );
  MUX2_X1 U350 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n403), .Z(n335) );
  MUX2_X1 U351 ( .A(n335), .B(n334), .S(N11), .Z(n336) );
  MUX2_X1 U352 ( .A(n336), .B(n333), .S(N12), .Z(n337) );
  MUX2_X1 U353 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n404), .Z(n338) );
  MUX2_X1 U354 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n404), .Z(n339) );
  MUX2_X1 U355 ( .A(n339), .B(n338), .S(N11), .Z(n340) );
  MUX2_X1 U356 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n404), .Z(n341) );
  MUX2_X1 U357 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n404), .Z(n342) );
  MUX2_X1 U358 ( .A(n342), .B(n341), .S(n401), .Z(n343) );
  MUX2_X1 U359 ( .A(n343), .B(n340), .S(N12), .Z(n344) );
  MUX2_X1 U360 ( .A(n344), .B(n337), .S(N13), .Z(N18) );
  MUX2_X1 U361 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n404), .Z(n345) );
  MUX2_X1 U362 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n404), .Z(n346) );
  MUX2_X1 U363 ( .A(n346), .B(n345), .S(N11), .Z(n347) );
  MUX2_X1 U364 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n404), .Z(n348) );
  MUX2_X1 U365 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n404), .Z(n349) );
  MUX2_X1 U366 ( .A(n349), .B(n348), .S(N11), .Z(n350) );
  MUX2_X1 U367 ( .A(n350), .B(n347), .S(N12), .Z(n351) );
  MUX2_X1 U368 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n404), .Z(n352) );
  MUX2_X1 U369 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n404), .Z(n353) );
  MUX2_X1 U370 ( .A(n353), .B(n352), .S(N11), .Z(n354) );
  MUX2_X1 U371 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n404), .Z(n355) );
  MUX2_X1 U372 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n404), .Z(n356) );
  MUX2_X1 U373 ( .A(n356), .B(n355), .S(n401), .Z(n357) );
  MUX2_X1 U374 ( .A(n357), .B(n354), .S(N12), .Z(n358) );
  MUX2_X1 U375 ( .A(n358), .B(n351), .S(N13), .Z(N17) );
  MUX2_X1 U376 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(N10), .Z(n359) );
  MUX2_X1 U377 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n404), .Z(n360) );
  MUX2_X1 U378 ( .A(n360), .B(n359), .S(n401), .Z(n361) );
  MUX2_X1 U379 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n403), .Z(n362) );
  MUX2_X1 U380 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n404), .Z(n363) );
  MUX2_X1 U381 ( .A(n363), .B(n362), .S(N11), .Z(n364) );
  MUX2_X1 U382 ( .A(n364), .B(n361), .S(N12), .Z(n365) );
  MUX2_X1 U383 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n403), .Z(n366) );
  MUX2_X1 U384 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n402), .Z(n367) );
  MUX2_X1 U385 ( .A(n367), .B(n366), .S(n401), .Z(n368) );
  MUX2_X1 U386 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n403), .Z(n369) );
  MUX2_X1 U387 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n403), .Z(n370) );
  MUX2_X1 U388 ( .A(n370), .B(n369), .S(N11), .Z(n371) );
  MUX2_X1 U389 ( .A(n371), .B(n368), .S(N12), .Z(n372) );
  MUX2_X1 U390 ( .A(n372), .B(n365), .S(N13), .Z(N16) );
  MUX2_X1 U391 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n402), .Z(n373) );
  MUX2_X1 U392 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n402), .Z(n374) );
  MUX2_X1 U393 ( .A(n374), .B(n373), .S(n401), .Z(n375) );
  MUX2_X1 U394 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n404), .Z(n376) );
  MUX2_X1 U395 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n402), .Z(n377) );
  MUX2_X1 U396 ( .A(n377), .B(n376), .S(N11), .Z(n378) );
  MUX2_X1 U397 ( .A(n378), .B(n375), .S(N12), .Z(n379) );
  MUX2_X1 U398 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n380) );
  MUX2_X1 U399 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n381) );
  MUX2_X1 U400 ( .A(n381), .B(n380), .S(N11), .Z(n382) );
  MUX2_X1 U401 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n383) );
  MUX2_X1 U402 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n402), .Z(n384) );
  MUX2_X1 U403 ( .A(n384), .B(n383), .S(N11), .Z(n385) );
  MUX2_X1 U404 ( .A(n385), .B(n382), .S(N12), .Z(n386) );
  MUX2_X1 U405 ( .A(n386), .B(n379), .S(N13), .Z(N15) );
  MUX2_X1 U406 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(N10), .Z(n387) );
  MUX2_X1 U407 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n388) );
  MUX2_X1 U408 ( .A(n388), .B(n387), .S(n401), .Z(n389) );
  MUX2_X1 U409 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(N10), .Z(n390) );
  MUX2_X1 U410 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n391) );
  MUX2_X1 U411 ( .A(n391), .B(n390), .S(N11), .Z(n392) );
  MUX2_X1 U412 ( .A(n392), .B(n389), .S(N12), .Z(n393) );
  MUX2_X1 U413 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n394) );
  MUX2_X1 U414 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n395) );
  MUX2_X1 U415 ( .A(n395), .B(n394), .S(N11), .Z(n396) );
  MUX2_X1 U416 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n397) );
  MUX2_X1 U417 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n404), .Z(n398) );
  MUX2_X1 U418 ( .A(n398), .B(n397), .S(N11), .Z(n399) );
  MUX2_X1 U419 ( .A(n399), .B(n396), .S(N12), .Z(n400) );
  MUX2_X1 U420 ( .A(n400), .B(n393), .S(N13), .Z(N14) );
  INV_X1 U421 ( .A(N10), .ZN(n405) );
  INV_X1 U422 ( .A(N11), .ZN(n406) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_2 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N16, N17, N18, N19, N20, N21, n1, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N21), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n412), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n413), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n414), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n415), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n416), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n417), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n418), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n419), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n420), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n421), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n422), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n423), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n424), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n425), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n426), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n427), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n428), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n429), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n430), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n431), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n432), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n433), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n434), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n435), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n436), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n437), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n438), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n439), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n440), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n441), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n442), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n443), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n444), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n445), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n446), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n447), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n448), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n449), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n450), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n451), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n452), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n453), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n454), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n455), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n456), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n457), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n458), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n459), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n460), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n461), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n462), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n463), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n464), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n465), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n466), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n467), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n468), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n469), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n470), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n471), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n472), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n473), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n474), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n475), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n476), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n477), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n478), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n479), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n480), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n481), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n482), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n483), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n484), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n485), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n486), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n487), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n488), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n489), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n490), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n491), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n492), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n493), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n494), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n495), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n496), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n497), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n498), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n499), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n500), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n501), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n502), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n503), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n504), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n505), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n506), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n507), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n508), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n509), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n510), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n511), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n512), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n513), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n514), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n515), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n516), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n517), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n518), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n519), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n520), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n521), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n522), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n523), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n524), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n525), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n526), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n527), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n528), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n529), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n530), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n531), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n532), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n533), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n534), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n535), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n536), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n537), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n538), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n539), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N20), .CK(clk), .Q(data_out[1]) );
  DFF_X2 \data_out_reg[5]  ( .D(N16), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .QN(n1) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(N10), .Z(n398) );
  BUF_X1 U5 ( .A(N10), .Z(n399) );
  BUF_X1 U6 ( .A(N10), .Z(n400) );
  BUF_X1 U7 ( .A(N11), .Z(n397) );
  NAND2_X1 U8 ( .A1(n663), .A2(n683), .ZN(n672) );
  NAND2_X1 U9 ( .A1(n663), .A2(n673), .ZN(n662) );
  NAND2_X1 U10 ( .A1(n684), .A2(n683), .ZN(n693) );
  NAND2_X1 U11 ( .A1(n673), .A2(n684), .ZN(n682) );
  NAND2_X1 U12 ( .A1(n605), .A2(n684), .ZN(n614) );
  NAND2_X1 U13 ( .A1(n595), .A2(n684), .ZN(n604) );
  NAND2_X1 U14 ( .A1(n605), .A2(n663), .ZN(n594) );
  NAND2_X1 U15 ( .A1(n595), .A2(n663), .ZN(n585) );
  NAND2_X1 U16 ( .A1(n644), .A2(n683), .ZN(n653) );
  NAND2_X1 U17 ( .A1(n644), .A2(n673), .ZN(n643) );
  NAND2_X1 U18 ( .A1(n625), .A2(n683), .ZN(n634) );
  NAND2_X1 U19 ( .A1(n625), .A2(n673), .ZN(n623) );
  NAND2_X1 U20 ( .A1(n605), .A2(n644), .ZN(n576) );
  NAND2_X1 U21 ( .A1(n595), .A2(n644), .ZN(n567) );
  NAND2_X1 U22 ( .A1(n605), .A2(n625), .ZN(n558) );
  NAND2_X1 U23 ( .A1(n595), .A2(n625), .ZN(n548) );
  AND2_X1 U24 ( .A1(n549), .A2(N10), .ZN(n595) );
  AND2_X1 U25 ( .A1(n549), .A2(n401), .ZN(n605) );
  AND2_X1 U26 ( .A1(N10), .A2(n624), .ZN(n673) );
  AND2_X1 U27 ( .A1(n624), .A2(n401), .ZN(n683) );
  OAI21_X1 U28 ( .B1(n693), .B2(n411), .A(n692), .ZN(n539) );
  NAND2_X1 U29 ( .A1(\mem[0][0] ), .A2(n693), .ZN(n692) );
  OAI21_X1 U30 ( .B1(n693), .B2(n410), .A(n691), .ZN(n538) );
  NAND2_X1 U31 ( .A1(\mem[0][1] ), .A2(n693), .ZN(n691) );
  OAI21_X1 U32 ( .B1(n693), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U33 ( .A1(\mem[0][2] ), .A2(n693), .ZN(n690) );
  OAI21_X1 U34 ( .B1(n693), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U35 ( .A1(\mem[0][3] ), .A2(n693), .ZN(n689) );
  OAI21_X1 U36 ( .B1(n693), .B2(n407), .A(n688), .ZN(n535) );
  NAND2_X1 U37 ( .A1(\mem[0][4] ), .A2(n693), .ZN(n688) );
  OAI21_X1 U38 ( .B1(n693), .B2(n406), .A(n687), .ZN(n534) );
  NAND2_X1 U39 ( .A1(\mem[0][5] ), .A2(n693), .ZN(n687) );
  OAI21_X1 U40 ( .B1(n693), .B2(n405), .A(n686), .ZN(n533) );
  NAND2_X1 U41 ( .A1(\mem[0][6] ), .A2(n693), .ZN(n686) );
  OAI21_X1 U42 ( .B1(n693), .B2(n404), .A(n685), .ZN(n532) );
  NAND2_X1 U43 ( .A1(\mem[0][7] ), .A2(n693), .ZN(n685) );
  OAI21_X1 U44 ( .B1(n411), .B2(n672), .A(n671), .ZN(n523) );
  NAND2_X1 U45 ( .A1(\mem[2][0] ), .A2(n672), .ZN(n671) );
  OAI21_X1 U46 ( .B1(n410), .B2(n672), .A(n670), .ZN(n522) );
  NAND2_X1 U47 ( .A1(\mem[2][1] ), .A2(n672), .ZN(n670) );
  OAI21_X1 U48 ( .B1(n409), .B2(n672), .A(n669), .ZN(n521) );
  NAND2_X1 U49 ( .A1(\mem[2][2] ), .A2(n672), .ZN(n669) );
  OAI21_X1 U50 ( .B1(n408), .B2(n672), .A(n668), .ZN(n520) );
  NAND2_X1 U51 ( .A1(\mem[2][3] ), .A2(n672), .ZN(n668) );
  OAI21_X1 U52 ( .B1(n407), .B2(n672), .A(n667), .ZN(n519) );
  NAND2_X1 U53 ( .A1(\mem[2][4] ), .A2(n672), .ZN(n667) );
  OAI21_X1 U54 ( .B1(n406), .B2(n672), .A(n666), .ZN(n518) );
  NAND2_X1 U55 ( .A1(\mem[2][5] ), .A2(n672), .ZN(n666) );
  OAI21_X1 U56 ( .B1(n405), .B2(n672), .A(n665), .ZN(n517) );
  NAND2_X1 U57 ( .A1(\mem[2][6] ), .A2(n672), .ZN(n665) );
  OAI21_X1 U58 ( .B1(n404), .B2(n672), .A(n664), .ZN(n516) );
  NAND2_X1 U59 ( .A1(\mem[2][7] ), .A2(n672), .ZN(n664) );
  OAI21_X1 U60 ( .B1(n411), .B2(n662), .A(n661), .ZN(n515) );
  NAND2_X1 U61 ( .A1(\mem[3][0] ), .A2(n662), .ZN(n661) );
  OAI21_X1 U62 ( .B1(n410), .B2(n662), .A(n660), .ZN(n514) );
  NAND2_X1 U63 ( .A1(\mem[3][1] ), .A2(n662), .ZN(n660) );
  OAI21_X1 U64 ( .B1(n409), .B2(n662), .A(n659), .ZN(n513) );
  NAND2_X1 U65 ( .A1(\mem[3][2] ), .A2(n662), .ZN(n659) );
  OAI21_X1 U66 ( .B1(n408), .B2(n662), .A(n658), .ZN(n512) );
  NAND2_X1 U67 ( .A1(\mem[3][3] ), .A2(n662), .ZN(n658) );
  OAI21_X1 U68 ( .B1(n407), .B2(n662), .A(n657), .ZN(n511) );
  NAND2_X1 U69 ( .A1(\mem[3][4] ), .A2(n662), .ZN(n657) );
  OAI21_X1 U70 ( .B1(n406), .B2(n662), .A(n656), .ZN(n510) );
  NAND2_X1 U71 ( .A1(\mem[3][5] ), .A2(n662), .ZN(n656) );
  OAI21_X1 U72 ( .B1(n405), .B2(n662), .A(n655), .ZN(n509) );
  NAND2_X1 U73 ( .A1(\mem[3][6] ), .A2(n662), .ZN(n655) );
  OAI21_X1 U74 ( .B1(n404), .B2(n662), .A(n654), .ZN(n508) );
  NAND2_X1 U75 ( .A1(\mem[3][7] ), .A2(n662), .ZN(n654) );
  NOR2_X1 U76 ( .A1(n403), .A2(N13), .ZN(n624) );
  INV_X1 U77 ( .A(wr_en), .ZN(n403) );
  OAI21_X1 U78 ( .B1(n411), .B2(n682), .A(n681), .ZN(n531) );
  NAND2_X1 U79 ( .A1(\mem[1][0] ), .A2(n682), .ZN(n681) );
  OAI21_X1 U80 ( .B1(n410), .B2(n682), .A(n680), .ZN(n530) );
  NAND2_X1 U81 ( .A1(\mem[1][1] ), .A2(n682), .ZN(n680) );
  OAI21_X1 U82 ( .B1(n409), .B2(n682), .A(n679), .ZN(n529) );
  NAND2_X1 U83 ( .A1(\mem[1][2] ), .A2(n682), .ZN(n679) );
  OAI21_X1 U84 ( .B1(n408), .B2(n682), .A(n678), .ZN(n528) );
  NAND2_X1 U85 ( .A1(\mem[1][3] ), .A2(n682), .ZN(n678) );
  OAI21_X1 U86 ( .B1(n407), .B2(n682), .A(n677), .ZN(n527) );
  NAND2_X1 U87 ( .A1(\mem[1][4] ), .A2(n682), .ZN(n677) );
  OAI21_X1 U88 ( .B1(n406), .B2(n682), .A(n676), .ZN(n526) );
  NAND2_X1 U89 ( .A1(\mem[1][5] ), .A2(n682), .ZN(n676) );
  OAI21_X1 U90 ( .B1(n405), .B2(n682), .A(n675), .ZN(n525) );
  NAND2_X1 U91 ( .A1(\mem[1][6] ), .A2(n682), .ZN(n675) );
  OAI21_X1 U92 ( .B1(n404), .B2(n682), .A(n674), .ZN(n524) );
  NAND2_X1 U93 ( .A1(\mem[1][7] ), .A2(n682), .ZN(n674) );
  OAI21_X1 U94 ( .B1(n411), .B2(n653), .A(n652), .ZN(n507) );
  NAND2_X1 U95 ( .A1(\mem[4][0] ), .A2(n653), .ZN(n652) );
  OAI21_X1 U96 ( .B1(n410), .B2(n653), .A(n651), .ZN(n506) );
  NAND2_X1 U97 ( .A1(\mem[4][1] ), .A2(n653), .ZN(n651) );
  OAI21_X1 U98 ( .B1(n409), .B2(n653), .A(n650), .ZN(n505) );
  NAND2_X1 U99 ( .A1(\mem[4][2] ), .A2(n653), .ZN(n650) );
  OAI21_X1 U100 ( .B1(n408), .B2(n653), .A(n649), .ZN(n504) );
  NAND2_X1 U101 ( .A1(\mem[4][3] ), .A2(n653), .ZN(n649) );
  OAI21_X1 U102 ( .B1(n407), .B2(n653), .A(n648), .ZN(n503) );
  NAND2_X1 U103 ( .A1(\mem[4][4] ), .A2(n653), .ZN(n648) );
  OAI21_X1 U104 ( .B1(n406), .B2(n653), .A(n647), .ZN(n502) );
  NAND2_X1 U105 ( .A1(\mem[4][5] ), .A2(n653), .ZN(n647) );
  OAI21_X1 U106 ( .B1(n405), .B2(n653), .A(n646), .ZN(n501) );
  NAND2_X1 U107 ( .A1(\mem[4][6] ), .A2(n653), .ZN(n646) );
  OAI21_X1 U108 ( .B1(n404), .B2(n653), .A(n645), .ZN(n500) );
  NAND2_X1 U109 ( .A1(\mem[4][7] ), .A2(n653), .ZN(n645) );
  OAI21_X1 U110 ( .B1(n411), .B2(n643), .A(n642), .ZN(n499) );
  NAND2_X1 U111 ( .A1(\mem[5][0] ), .A2(n643), .ZN(n642) );
  OAI21_X1 U112 ( .B1(n410), .B2(n643), .A(n641), .ZN(n498) );
  NAND2_X1 U113 ( .A1(\mem[5][1] ), .A2(n643), .ZN(n641) );
  OAI21_X1 U114 ( .B1(n409), .B2(n643), .A(n640), .ZN(n497) );
  NAND2_X1 U115 ( .A1(\mem[5][2] ), .A2(n643), .ZN(n640) );
  OAI21_X1 U116 ( .B1(n408), .B2(n643), .A(n639), .ZN(n496) );
  NAND2_X1 U117 ( .A1(\mem[5][3] ), .A2(n643), .ZN(n639) );
  OAI21_X1 U118 ( .B1(n407), .B2(n643), .A(n638), .ZN(n495) );
  NAND2_X1 U119 ( .A1(\mem[5][4] ), .A2(n643), .ZN(n638) );
  OAI21_X1 U120 ( .B1(n406), .B2(n643), .A(n637), .ZN(n494) );
  NAND2_X1 U121 ( .A1(\mem[5][5] ), .A2(n643), .ZN(n637) );
  OAI21_X1 U122 ( .B1(n405), .B2(n643), .A(n636), .ZN(n493) );
  NAND2_X1 U123 ( .A1(\mem[5][6] ), .A2(n643), .ZN(n636) );
  OAI21_X1 U124 ( .B1(n404), .B2(n643), .A(n635), .ZN(n492) );
  NAND2_X1 U125 ( .A1(\mem[5][7] ), .A2(n643), .ZN(n635) );
  OAI21_X1 U126 ( .B1(n411), .B2(n634), .A(n633), .ZN(n491) );
  NAND2_X1 U127 ( .A1(\mem[6][0] ), .A2(n634), .ZN(n633) );
  OAI21_X1 U128 ( .B1(n410), .B2(n634), .A(n632), .ZN(n490) );
  NAND2_X1 U129 ( .A1(\mem[6][1] ), .A2(n634), .ZN(n632) );
  OAI21_X1 U130 ( .B1(n409), .B2(n634), .A(n631), .ZN(n489) );
  NAND2_X1 U131 ( .A1(\mem[6][2] ), .A2(n634), .ZN(n631) );
  OAI21_X1 U132 ( .B1(n408), .B2(n634), .A(n630), .ZN(n488) );
  NAND2_X1 U133 ( .A1(\mem[6][3] ), .A2(n634), .ZN(n630) );
  OAI21_X1 U134 ( .B1(n407), .B2(n634), .A(n629), .ZN(n487) );
  NAND2_X1 U135 ( .A1(\mem[6][4] ), .A2(n634), .ZN(n629) );
  OAI21_X1 U136 ( .B1(n406), .B2(n634), .A(n628), .ZN(n486) );
  NAND2_X1 U137 ( .A1(\mem[6][5] ), .A2(n634), .ZN(n628) );
  OAI21_X1 U138 ( .B1(n405), .B2(n634), .A(n627), .ZN(n485) );
  NAND2_X1 U139 ( .A1(\mem[6][6] ), .A2(n634), .ZN(n627) );
  OAI21_X1 U140 ( .B1(n404), .B2(n634), .A(n626), .ZN(n484) );
  NAND2_X1 U141 ( .A1(\mem[6][7] ), .A2(n634), .ZN(n626) );
  OAI21_X1 U142 ( .B1(n411), .B2(n623), .A(n622), .ZN(n483) );
  NAND2_X1 U143 ( .A1(\mem[7][0] ), .A2(n623), .ZN(n622) );
  OAI21_X1 U144 ( .B1(n410), .B2(n623), .A(n621), .ZN(n482) );
  NAND2_X1 U145 ( .A1(\mem[7][1] ), .A2(n623), .ZN(n621) );
  OAI21_X1 U146 ( .B1(n409), .B2(n623), .A(n620), .ZN(n481) );
  NAND2_X1 U147 ( .A1(\mem[7][2] ), .A2(n623), .ZN(n620) );
  OAI21_X1 U148 ( .B1(n408), .B2(n623), .A(n619), .ZN(n480) );
  NAND2_X1 U149 ( .A1(\mem[7][3] ), .A2(n623), .ZN(n619) );
  OAI21_X1 U150 ( .B1(n407), .B2(n623), .A(n618), .ZN(n479) );
  NAND2_X1 U151 ( .A1(\mem[7][4] ), .A2(n623), .ZN(n618) );
  OAI21_X1 U152 ( .B1(n406), .B2(n623), .A(n617), .ZN(n478) );
  NAND2_X1 U153 ( .A1(\mem[7][5] ), .A2(n623), .ZN(n617) );
  OAI21_X1 U154 ( .B1(n405), .B2(n623), .A(n616), .ZN(n477) );
  NAND2_X1 U155 ( .A1(\mem[7][6] ), .A2(n623), .ZN(n616) );
  OAI21_X1 U156 ( .B1(n404), .B2(n623), .A(n615), .ZN(n476) );
  NAND2_X1 U157 ( .A1(\mem[7][7] ), .A2(n623), .ZN(n615) );
  OAI21_X1 U158 ( .B1(n411), .B2(n614), .A(n613), .ZN(n475) );
  NAND2_X1 U159 ( .A1(\mem[8][0] ), .A2(n614), .ZN(n613) );
  OAI21_X1 U160 ( .B1(n410), .B2(n614), .A(n612), .ZN(n474) );
  NAND2_X1 U161 ( .A1(\mem[8][1] ), .A2(n614), .ZN(n612) );
  OAI21_X1 U162 ( .B1(n409), .B2(n614), .A(n611), .ZN(n473) );
  NAND2_X1 U163 ( .A1(\mem[8][2] ), .A2(n614), .ZN(n611) );
  OAI21_X1 U164 ( .B1(n408), .B2(n614), .A(n610), .ZN(n472) );
  NAND2_X1 U165 ( .A1(\mem[8][3] ), .A2(n614), .ZN(n610) );
  OAI21_X1 U166 ( .B1(n407), .B2(n614), .A(n609), .ZN(n471) );
  NAND2_X1 U167 ( .A1(\mem[8][4] ), .A2(n614), .ZN(n609) );
  OAI21_X1 U168 ( .B1(n406), .B2(n614), .A(n608), .ZN(n470) );
  NAND2_X1 U169 ( .A1(\mem[8][5] ), .A2(n614), .ZN(n608) );
  OAI21_X1 U170 ( .B1(n405), .B2(n614), .A(n607), .ZN(n469) );
  NAND2_X1 U171 ( .A1(\mem[8][6] ), .A2(n614), .ZN(n607) );
  OAI21_X1 U172 ( .B1(n404), .B2(n614), .A(n606), .ZN(n468) );
  NAND2_X1 U173 ( .A1(\mem[8][7] ), .A2(n614), .ZN(n606) );
  OAI21_X1 U174 ( .B1(n411), .B2(n604), .A(n603), .ZN(n467) );
  NAND2_X1 U175 ( .A1(\mem[9][0] ), .A2(n604), .ZN(n603) );
  OAI21_X1 U176 ( .B1(n410), .B2(n604), .A(n602), .ZN(n466) );
  NAND2_X1 U177 ( .A1(\mem[9][1] ), .A2(n604), .ZN(n602) );
  OAI21_X1 U178 ( .B1(n409), .B2(n604), .A(n601), .ZN(n465) );
  NAND2_X1 U179 ( .A1(\mem[9][2] ), .A2(n604), .ZN(n601) );
  OAI21_X1 U180 ( .B1(n408), .B2(n604), .A(n600), .ZN(n464) );
  NAND2_X1 U181 ( .A1(\mem[9][3] ), .A2(n604), .ZN(n600) );
  OAI21_X1 U182 ( .B1(n407), .B2(n604), .A(n599), .ZN(n463) );
  NAND2_X1 U183 ( .A1(\mem[9][4] ), .A2(n604), .ZN(n599) );
  OAI21_X1 U184 ( .B1(n406), .B2(n604), .A(n598), .ZN(n462) );
  NAND2_X1 U185 ( .A1(\mem[9][5] ), .A2(n604), .ZN(n598) );
  OAI21_X1 U186 ( .B1(n405), .B2(n604), .A(n597), .ZN(n461) );
  NAND2_X1 U187 ( .A1(\mem[9][6] ), .A2(n604), .ZN(n597) );
  OAI21_X1 U188 ( .B1(n404), .B2(n604), .A(n596), .ZN(n460) );
  NAND2_X1 U189 ( .A1(\mem[9][7] ), .A2(n604), .ZN(n596) );
  OAI21_X1 U190 ( .B1(n411), .B2(n594), .A(n593), .ZN(n459) );
  NAND2_X1 U191 ( .A1(\mem[10][0] ), .A2(n594), .ZN(n593) );
  OAI21_X1 U192 ( .B1(n410), .B2(n594), .A(n592), .ZN(n458) );
  NAND2_X1 U193 ( .A1(\mem[10][1] ), .A2(n594), .ZN(n592) );
  OAI21_X1 U194 ( .B1(n409), .B2(n594), .A(n591), .ZN(n457) );
  NAND2_X1 U195 ( .A1(\mem[10][2] ), .A2(n594), .ZN(n591) );
  OAI21_X1 U196 ( .B1(n408), .B2(n594), .A(n590), .ZN(n456) );
  NAND2_X1 U197 ( .A1(\mem[10][3] ), .A2(n594), .ZN(n590) );
  OAI21_X1 U198 ( .B1(n407), .B2(n594), .A(n589), .ZN(n455) );
  NAND2_X1 U199 ( .A1(\mem[10][4] ), .A2(n594), .ZN(n589) );
  OAI21_X1 U200 ( .B1(n406), .B2(n594), .A(n588), .ZN(n454) );
  NAND2_X1 U201 ( .A1(\mem[10][5] ), .A2(n594), .ZN(n588) );
  OAI21_X1 U202 ( .B1(n405), .B2(n594), .A(n587), .ZN(n453) );
  NAND2_X1 U203 ( .A1(\mem[10][6] ), .A2(n594), .ZN(n587) );
  OAI21_X1 U204 ( .B1(n404), .B2(n594), .A(n586), .ZN(n452) );
  NAND2_X1 U205 ( .A1(\mem[10][7] ), .A2(n594), .ZN(n586) );
  OAI21_X1 U206 ( .B1(n411), .B2(n585), .A(n584), .ZN(n451) );
  NAND2_X1 U207 ( .A1(\mem[11][0] ), .A2(n585), .ZN(n584) );
  OAI21_X1 U208 ( .B1(n410), .B2(n585), .A(n583), .ZN(n450) );
  NAND2_X1 U209 ( .A1(\mem[11][1] ), .A2(n585), .ZN(n583) );
  OAI21_X1 U210 ( .B1(n409), .B2(n585), .A(n582), .ZN(n449) );
  NAND2_X1 U211 ( .A1(\mem[11][2] ), .A2(n585), .ZN(n582) );
  OAI21_X1 U212 ( .B1(n408), .B2(n585), .A(n581), .ZN(n448) );
  NAND2_X1 U213 ( .A1(\mem[11][3] ), .A2(n585), .ZN(n581) );
  OAI21_X1 U214 ( .B1(n407), .B2(n585), .A(n580), .ZN(n447) );
  NAND2_X1 U215 ( .A1(\mem[11][4] ), .A2(n585), .ZN(n580) );
  OAI21_X1 U216 ( .B1(n406), .B2(n585), .A(n579), .ZN(n446) );
  NAND2_X1 U217 ( .A1(\mem[11][5] ), .A2(n585), .ZN(n579) );
  OAI21_X1 U218 ( .B1(n405), .B2(n585), .A(n578), .ZN(n445) );
  NAND2_X1 U219 ( .A1(\mem[11][6] ), .A2(n585), .ZN(n578) );
  OAI21_X1 U220 ( .B1(n404), .B2(n585), .A(n577), .ZN(n444) );
  NAND2_X1 U221 ( .A1(\mem[11][7] ), .A2(n585), .ZN(n577) );
  OAI21_X1 U222 ( .B1(n411), .B2(n576), .A(n575), .ZN(n443) );
  NAND2_X1 U223 ( .A1(\mem[12][0] ), .A2(n576), .ZN(n575) );
  OAI21_X1 U224 ( .B1(n410), .B2(n576), .A(n574), .ZN(n442) );
  NAND2_X1 U225 ( .A1(\mem[12][1] ), .A2(n576), .ZN(n574) );
  OAI21_X1 U226 ( .B1(n409), .B2(n576), .A(n573), .ZN(n441) );
  NAND2_X1 U227 ( .A1(\mem[12][2] ), .A2(n576), .ZN(n573) );
  OAI21_X1 U228 ( .B1(n408), .B2(n576), .A(n572), .ZN(n440) );
  NAND2_X1 U229 ( .A1(\mem[12][3] ), .A2(n576), .ZN(n572) );
  OAI21_X1 U230 ( .B1(n407), .B2(n576), .A(n571), .ZN(n439) );
  NAND2_X1 U231 ( .A1(\mem[12][4] ), .A2(n576), .ZN(n571) );
  OAI21_X1 U232 ( .B1(n406), .B2(n576), .A(n570), .ZN(n438) );
  NAND2_X1 U233 ( .A1(\mem[12][5] ), .A2(n576), .ZN(n570) );
  OAI21_X1 U234 ( .B1(n405), .B2(n576), .A(n569), .ZN(n437) );
  NAND2_X1 U235 ( .A1(\mem[12][6] ), .A2(n576), .ZN(n569) );
  OAI21_X1 U236 ( .B1(n404), .B2(n576), .A(n568), .ZN(n436) );
  NAND2_X1 U237 ( .A1(\mem[12][7] ), .A2(n576), .ZN(n568) );
  OAI21_X1 U238 ( .B1(n411), .B2(n567), .A(n566), .ZN(n435) );
  NAND2_X1 U239 ( .A1(\mem[13][0] ), .A2(n567), .ZN(n566) );
  OAI21_X1 U240 ( .B1(n410), .B2(n567), .A(n565), .ZN(n434) );
  NAND2_X1 U241 ( .A1(\mem[13][1] ), .A2(n567), .ZN(n565) );
  OAI21_X1 U242 ( .B1(n409), .B2(n567), .A(n564), .ZN(n433) );
  NAND2_X1 U243 ( .A1(\mem[13][2] ), .A2(n567), .ZN(n564) );
  OAI21_X1 U244 ( .B1(n408), .B2(n567), .A(n563), .ZN(n432) );
  NAND2_X1 U245 ( .A1(\mem[13][3] ), .A2(n567), .ZN(n563) );
  OAI21_X1 U246 ( .B1(n407), .B2(n567), .A(n562), .ZN(n431) );
  NAND2_X1 U247 ( .A1(\mem[13][4] ), .A2(n567), .ZN(n562) );
  OAI21_X1 U248 ( .B1(n406), .B2(n567), .A(n561), .ZN(n430) );
  NAND2_X1 U249 ( .A1(\mem[13][5] ), .A2(n567), .ZN(n561) );
  OAI21_X1 U250 ( .B1(n405), .B2(n567), .A(n560), .ZN(n429) );
  NAND2_X1 U251 ( .A1(\mem[13][6] ), .A2(n567), .ZN(n560) );
  OAI21_X1 U252 ( .B1(n404), .B2(n567), .A(n559), .ZN(n428) );
  NAND2_X1 U253 ( .A1(\mem[13][7] ), .A2(n567), .ZN(n559) );
  OAI21_X1 U254 ( .B1(n411), .B2(n558), .A(n557), .ZN(n427) );
  NAND2_X1 U255 ( .A1(\mem[14][0] ), .A2(n558), .ZN(n557) );
  OAI21_X1 U256 ( .B1(n410), .B2(n558), .A(n556), .ZN(n426) );
  NAND2_X1 U257 ( .A1(\mem[14][1] ), .A2(n558), .ZN(n556) );
  OAI21_X1 U258 ( .B1(n409), .B2(n558), .A(n555), .ZN(n425) );
  NAND2_X1 U259 ( .A1(\mem[14][2] ), .A2(n558), .ZN(n555) );
  OAI21_X1 U260 ( .B1(n408), .B2(n558), .A(n554), .ZN(n424) );
  NAND2_X1 U261 ( .A1(\mem[14][3] ), .A2(n558), .ZN(n554) );
  OAI21_X1 U262 ( .B1(n407), .B2(n558), .A(n553), .ZN(n423) );
  NAND2_X1 U263 ( .A1(\mem[14][4] ), .A2(n558), .ZN(n553) );
  OAI21_X1 U264 ( .B1(n406), .B2(n558), .A(n552), .ZN(n422) );
  NAND2_X1 U265 ( .A1(\mem[14][5] ), .A2(n558), .ZN(n552) );
  OAI21_X1 U266 ( .B1(n405), .B2(n558), .A(n551), .ZN(n421) );
  NAND2_X1 U267 ( .A1(\mem[14][6] ), .A2(n558), .ZN(n551) );
  OAI21_X1 U268 ( .B1(n404), .B2(n558), .A(n550), .ZN(n420) );
  NAND2_X1 U269 ( .A1(\mem[14][7] ), .A2(n558), .ZN(n550) );
  OAI21_X1 U270 ( .B1(n411), .B2(n548), .A(n547), .ZN(n419) );
  NAND2_X1 U271 ( .A1(\mem[15][0] ), .A2(n548), .ZN(n547) );
  OAI21_X1 U272 ( .B1(n410), .B2(n548), .A(n546), .ZN(n418) );
  NAND2_X1 U273 ( .A1(\mem[15][1] ), .A2(n548), .ZN(n546) );
  OAI21_X1 U274 ( .B1(n409), .B2(n548), .A(n545), .ZN(n417) );
  NAND2_X1 U275 ( .A1(\mem[15][2] ), .A2(n548), .ZN(n545) );
  OAI21_X1 U276 ( .B1(n408), .B2(n548), .A(n544), .ZN(n416) );
  NAND2_X1 U277 ( .A1(\mem[15][3] ), .A2(n548), .ZN(n544) );
  OAI21_X1 U278 ( .B1(n407), .B2(n548), .A(n543), .ZN(n415) );
  NAND2_X1 U279 ( .A1(\mem[15][4] ), .A2(n548), .ZN(n543) );
  OAI21_X1 U280 ( .B1(n406), .B2(n548), .A(n542), .ZN(n414) );
  NAND2_X1 U281 ( .A1(\mem[15][5] ), .A2(n548), .ZN(n542) );
  OAI21_X1 U282 ( .B1(n405), .B2(n548), .A(n541), .ZN(n413) );
  NAND2_X1 U283 ( .A1(\mem[15][6] ), .A2(n548), .ZN(n541) );
  OAI21_X1 U284 ( .B1(n404), .B2(n548), .A(n540), .ZN(n412) );
  NAND2_X1 U285 ( .A1(\mem[15][7] ), .A2(n548), .ZN(n540) );
  AND2_X1 U286 ( .A1(N13), .A2(wr_en), .ZN(n549) );
  NOR2_X1 U287 ( .A1(N11), .A2(N12), .ZN(n684) );
  NOR2_X1 U288 ( .A1(n402), .A2(N12), .ZN(n663) );
  AND2_X1 U289 ( .A1(N12), .A2(n402), .ZN(n644) );
  AND2_X1 U290 ( .A1(N12), .A2(N11), .ZN(n625) );
  INV_X1 U291 ( .A(data_in[0]), .ZN(n411) );
  INV_X1 U292 ( .A(data_in[1]), .ZN(n410) );
  INV_X1 U293 ( .A(data_in[2]), .ZN(n409) );
  INV_X1 U294 ( .A(data_in[3]), .ZN(n408) );
  INV_X1 U295 ( .A(data_in[4]), .ZN(n407) );
  INV_X1 U296 ( .A(data_in[5]), .ZN(n406) );
  INV_X1 U297 ( .A(data_in[6]), .ZN(n405) );
  INV_X1 U298 ( .A(data_in[7]), .ZN(n404) );
  MUX2_X1 U299 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(N10), .Z(n3) );
  MUX2_X1 U300 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(N10), .Z(n4) );
  MUX2_X1 U301 ( .A(n4), .B(n3), .S(n397), .Z(n5) );
  MUX2_X1 U302 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(N10), .Z(n6) );
  MUX2_X1 U303 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n7) );
  MUX2_X1 U304 ( .A(n7), .B(n6), .S(N11), .Z(n8) );
  MUX2_X1 U305 ( .A(n8), .B(n5), .S(N12), .Z(n9) );
  MUX2_X1 U306 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(N10), .Z(n10) );
  MUX2_X1 U307 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n399), .Z(n11) );
  MUX2_X1 U308 ( .A(n11), .B(n10), .S(N11), .Z(n294) );
  MUX2_X1 U309 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(N10), .Z(n295) );
  MUX2_X1 U310 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n296) );
  MUX2_X1 U311 ( .A(n296), .B(n295), .S(N11), .Z(n297) );
  MUX2_X1 U312 ( .A(n297), .B(n294), .S(N12), .Z(n298) );
  MUX2_X1 U313 ( .A(n298), .B(n9), .S(N13), .Z(N21) );
  MUX2_X1 U314 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n400), .Z(n299) );
  MUX2_X1 U315 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(N10), .Z(n300) );
  MUX2_X1 U316 ( .A(n300), .B(n299), .S(N11), .Z(n301) );
  MUX2_X1 U317 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(N10), .Z(n302) );
  MUX2_X1 U318 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n398), .Z(n303) );
  MUX2_X1 U319 ( .A(n303), .B(n302), .S(N11), .Z(n304) );
  MUX2_X1 U320 ( .A(n304), .B(n301), .S(N12), .Z(n305) );
  MUX2_X1 U321 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(N10), .Z(n306) );
  MUX2_X1 U322 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n399), .Z(n307) );
  MUX2_X1 U323 ( .A(n307), .B(n306), .S(N11), .Z(n308) );
  MUX2_X1 U324 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(N10), .Z(n309) );
  MUX2_X1 U325 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(N10), .Z(n310) );
  MUX2_X1 U326 ( .A(n310), .B(n309), .S(N11), .Z(n311) );
  MUX2_X1 U327 ( .A(n311), .B(n308), .S(N12), .Z(n312) );
  MUX2_X1 U328 ( .A(n312), .B(n305), .S(N13), .Z(N20) );
  MUX2_X1 U329 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n398), .Z(n313) );
  MUX2_X1 U330 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n398), .Z(n314) );
  MUX2_X1 U331 ( .A(n314), .B(n313), .S(n397), .Z(n315) );
  MUX2_X1 U332 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n398), .Z(n316) );
  MUX2_X1 U333 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n398), .Z(n317) );
  MUX2_X1 U334 ( .A(n317), .B(n316), .S(n397), .Z(n318) );
  MUX2_X1 U335 ( .A(n318), .B(n315), .S(N12), .Z(n319) );
  MUX2_X1 U336 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n398), .Z(n320) );
  MUX2_X1 U337 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n398), .Z(n321) );
  MUX2_X1 U338 ( .A(n321), .B(n320), .S(n397), .Z(n322) );
  MUX2_X1 U339 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n398), .Z(n323) );
  MUX2_X1 U340 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n398), .Z(n324) );
  MUX2_X1 U341 ( .A(n324), .B(n323), .S(n397), .Z(n325) );
  MUX2_X1 U342 ( .A(n325), .B(n322), .S(N12), .Z(n326) );
  MUX2_X1 U343 ( .A(n326), .B(n319), .S(N13), .Z(N19) );
  MUX2_X1 U344 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n398), .Z(n327) );
  MUX2_X1 U345 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n398), .Z(n328) );
  MUX2_X1 U346 ( .A(n328), .B(n327), .S(n397), .Z(n329) );
  MUX2_X1 U347 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n398), .Z(n330) );
  MUX2_X1 U348 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n398), .Z(n331) );
  MUX2_X1 U349 ( .A(n331), .B(n330), .S(n397), .Z(n332) );
  MUX2_X1 U350 ( .A(n332), .B(n329), .S(N12), .Z(n333) );
  MUX2_X1 U351 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n399), .Z(n334) );
  MUX2_X1 U352 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n399), .Z(n335) );
  MUX2_X1 U353 ( .A(n335), .B(n334), .S(n397), .Z(n336) );
  MUX2_X1 U354 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n399), .Z(n337) );
  MUX2_X1 U355 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n399), .Z(n338) );
  MUX2_X1 U356 ( .A(n338), .B(n337), .S(n397), .Z(n339) );
  MUX2_X1 U357 ( .A(n339), .B(n336), .S(N12), .Z(n340) );
  MUX2_X1 U358 ( .A(n340), .B(n333), .S(N13), .Z(N18) );
  MUX2_X1 U359 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n399), .Z(n341) );
  MUX2_X1 U360 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n399), .Z(n342) );
  MUX2_X1 U361 ( .A(n342), .B(n341), .S(n397), .Z(n343) );
  MUX2_X1 U362 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n399), .Z(n344) );
  MUX2_X1 U363 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n399), .Z(n345) );
  MUX2_X1 U364 ( .A(n345), .B(n344), .S(n397), .Z(n346) );
  MUX2_X1 U365 ( .A(n346), .B(n343), .S(N12), .Z(n347) );
  MUX2_X1 U366 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n399), .Z(n348) );
  MUX2_X1 U367 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n399), .Z(n349) );
  MUX2_X1 U368 ( .A(n349), .B(n348), .S(n397), .Z(n350) );
  MUX2_X1 U369 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n399), .Z(n351) );
  MUX2_X1 U370 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n399), .Z(n352) );
  MUX2_X1 U371 ( .A(n352), .B(n351), .S(n397), .Z(n353) );
  MUX2_X1 U372 ( .A(n353), .B(n350), .S(N12), .Z(n354) );
  MUX2_X1 U373 ( .A(n354), .B(n347), .S(N13), .Z(N17) );
  MUX2_X1 U374 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n400), .Z(n355) );
  MUX2_X1 U375 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n400), .Z(n356) );
  MUX2_X1 U376 ( .A(n356), .B(n355), .S(N11), .Z(n357) );
  MUX2_X1 U377 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n400), .Z(n358) );
  MUX2_X1 U378 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n400), .Z(n359) );
  MUX2_X1 U379 ( .A(n359), .B(n358), .S(N11), .Z(n360) );
  MUX2_X1 U380 ( .A(n360), .B(n357), .S(N12), .Z(n361) );
  MUX2_X1 U381 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n400), .Z(n362) );
  MUX2_X1 U382 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n400), .Z(n363) );
  MUX2_X1 U383 ( .A(n363), .B(n362), .S(N11), .Z(n364) );
  MUX2_X1 U384 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n400), .Z(n365) );
  MUX2_X1 U385 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n400), .Z(n366) );
  MUX2_X1 U386 ( .A(n366), .B(n365), .S(N11), .Z(n367) );
  MUX2_X1 U387 ( .A(n367), .B(n364), .S(N12), .Z(n368) );
  MUX2_X1 U388 ( .A(n368), .B(n361), .S(N13), .Z(N16) );
  MUX2_X1 U389 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n400), .Z(n369) );
  MUX2_X1 U390 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n400), .Z(n370) );
  MUX2_X1 U391 ( .A(n370), .B(n369), .S(N11), .Z(n371) );
  MUX2_X1 U392 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n400), .Z(n372) );
  MUX2_X1 U393 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n400), .Z(n373) );
  MUX2_X1 U394 ( .A(n373), .B(n372), .S(N11), .Z(n374) );
  MUX2_X1 U395 ( .A(n374), .B(n371), .S(N12), .Z(n375) );
  MUX2_X1 U396 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n376) );
  MUX2_X1 U397 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n398), .Z(n377) );
  MUX2_X1 U398 ( .A(n377), .B(n376), .S(N11), .Z(n378) );
  MUX2_X1 U399 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n379) );
  MUX2_X1 U400 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n399), .Z(n380) );
  MUX2_X1 U401 ( .A(n380), .B(n379), .S(N11), .Z(n381) );
  MUX2_X1 U402 ( .A(n381), .B(n378), .S(N12), .Z(n382) );
  MUX2_X1 U403 ( .A(n382), .B(n375), .S(N13), .Z(N15) );
  MUX2_X1 U404 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n398), .Z(n383) );
  MUX2_X1 U405 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n384) );
  MUX2_X1 U406 ( .A(n384), .B(n383), .S(N11), .Z(n385) );
  MUX2_X1 U407 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n399), .Z(n386) );
  MUX2_X1 U408 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n400), .Z(n387) );
  MUX2_X1 U409 ( .A(n387), .B(n386), .S(N11), .Z(n388) );
  MUX2_X1 U410 ( .A(n388), .B(n385), .S(N12), .Z(n389) );
  MUX2_X1 U411 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n390) );
  MUX2_X1 U412 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n400), .Z(n391) );
  MUX2_X1 U413 ( .A(n391), .B(n390), .S(N11), .Z(n392) );
  MUX2_X1 U414 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n398), .Z(n393) );
  MUX2_X1 U415 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n400), .Z(n394) );
  MUX2_X1 U416 ( .A(n394), .B(n393), .S(n397), .Z(n395) );
  MUX2_X1 U417 ( .A(n395), .B(n392), .S(N12), .Z(n396) );
  MUX2_X1 U418 ( .A(n396), .B(n389), .S(N13), .Z(N14) );
  INV_X1 U419 ( .A(N10), .ZN(n401) );
  INV_X1 U420 ( .A(N11), .ZN(n402) );
endmodule


module memory_WIDTH8_SIZE16_LOGSIZE4_1 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][7] , \mem[15][6] , \mem[15][5] ,
         \mem[15][4] , \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] ,
         \mem[14][7] , \mem[14][6] , \mem[14][5] , \mem[14][4] , \mem[14][3] ,
         \mem[14][2] , \mem[14][1] , \mem[14][0] , \mem[13][7] , \mem[13][6] ,
         \mem[13][5] , \mem[13][4] , \mem[13][3] , \mem[13][2] , \mem[13][1] ,
         \mem[13][0] , \mem[12][7] , \mem[12][6] , \mem[12][5] , \mem[12][4] ,
         \mem[12][3] , \mem[12][2] , \mem[12][1] , \mem[12][0] , \mem[11][7] ,
         \mem[11][6] , \mem[11][5] , \mem[11][4] , \mem[11][3] , \mem[11][2] ,
         \mem[11][1] , \mem[11][0] , \mem[10][7] , \mem[10][6] , \mem[10][5] ,
         \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] , \mem[10][0] ,
         \mem[9][7] , \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] ,
         \mem[9][2] , \mem[9][1] , \mem[9][0] , \mem[8][7] , \mem[8][6] ,
         \mem[8][5] , \mem[8][4] , \mem[8][3] , \mem[8][2] , \mem[8][1] ,
         \mem[8][0] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][7] ,
         \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] , \mem[6][2] ,
         \mem[6][1] , \mem[6][0] , \mem[5][7] , \mem[5][6] , \mem[5][5] ,
         \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] ,
         \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] ,
         \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][7] ,
         \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] , \mem[1][2] ,
         \mem[1][1] , \mem[1][0] , \mem[0][7] , \mem[0][6] , \mem[0][5] ,
         \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14,
         N15, N17, N18, N19, N20, n3, n4, n5, n6, n7, n8, n9, n10, n11, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[7]  ( .D(N14), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N15), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N17), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N19), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[15][7]  ( .D(n414), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n415), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n416), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n417), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n418), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n419), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n420), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n421), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n422), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n423), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n424), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n425), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n426), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n427), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n428), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n429), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n430), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n431), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n432), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n433), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n434), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n435), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n436), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n437), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n438), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n439), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n440), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n441), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n442), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n443), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n444), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n445), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n446), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n447), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n448), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n449), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n450), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n451), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n452), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n453), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n454), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n455), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n456), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n457), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n458), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n459), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n460), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n461), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n462), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n463), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n464), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n465), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n466), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n467), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n468), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n469), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n470), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n471), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n472), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n473), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n474), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n475), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n476), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n477), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n478), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n479), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n480), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n481), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n482), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n483), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n484), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n485), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n486), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n487), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n488), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n489), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n490), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n491), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n492), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n493), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n494), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n495), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n496), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n497), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n498), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n499), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n500), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n501), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n502), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n503), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n504), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n505), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n506), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n507), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n508), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n509), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n510), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n511), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n512), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n513), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n514), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n515), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n516), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n517), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n518), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n519), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n520), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n521), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n522), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n523), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n524), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n525), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n526), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n527), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n528), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n529), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n530), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n531), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n532), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n533), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n534), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n535), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n536), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n537), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n538), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n539), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n540), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n541), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N20), .CK(clk), .QN(n401) );
  DFF_X1 \data_out_reg[3]  ( .D(N18), .CK(clk), .Q(data_out[3]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n368), .SI(n361), .SE(N13), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n298), .SI(n9), .SE(N13), .CK(clk), .Q(
        data_out[0]) );
  BUF_X1 U3 ( .A(N10), .Z(n399) );
  BUF_X1 U4 ( .A(N10), .Z(n400) );
  BUF_X1 U5 ( .A(N11), .Z(n397) );
  NAND2_X1 U6 ( .A1(n665), .A2(n685), .ZN(n674) );
  NAND2_X1 U7 ( .A1(n665), .A2(n675), .ZN(n664) );
  NAND2_X1 U8 ( .A1(n686), .A2(n685), .ZN(n695) );
  NAND2_X1 U9 ( .A1(n675), .A2(n686), .ZN(n684) );
  NAND2_X1 U10 ( .A1(n607), .A2(n686), .ZN(n616) );
  NAND2_X1 U11 ( .A1(n597), .A2(n686), .ZN(n606) );
  NAND2_X1 U12 ( .A1(n607), .A2(n665), .ZN(n596) );
  NAND2_X1 U13 ( .A1(n597), .A2(n665), .ZN(n587) );
  NAND2_X1 U14 ( .A1(n646), .A2(n685), .ZN(n655) );
  NAND2_X1 U15 ( .A1(n646), .A2(n675), .ZN(n645) );
  NAND2_X1 U16 ( .A1(n627), .A2(n685), .ZN(n636) );
  NAND2_X1 U17 ( .A1(n627), .A2(n675), .ZN(n625) );
  NAND2_X1 U18 ( .A1(n607), .A2(n646), .ZN(n578) );
  NAND2_X1 U19 ( .A1(n597), .A2(n646), .ZN(n569) );
  NAND2_X1 U20 ( .A1(n607), .A2(n627), .ZN(n560) );
  NAND2_X1 U21 ( .A1(n597), .A2(n627), .ZN(n550) );
  AND2_X1 U22 ( .A1(n551), .A2(N10), .ZN(n597) );
  AND2_X1 U23 ( .A1(n551), .A2(n403), .ZN(n607) );
  AND2_X1 U24 ( .A1(N10), .A2(n626), .ZN(n675) );
  AND2_X1 U25 ( .A1(n626), .A2(n403), .ZN(n685) );
  OAI21_X1 U26 ( .B1(n695), .B2(n413), .A(n694), .ZN(n541) );
  NAND2_X1 U27 ( .A1(\mem[0][0] ), .A2(n695), .ZN(n694) );
  OAI21_X1 U28 ( .B1(n695), .B2(n412), .A(n693), .ZN(n540) );
  NAND2_X1 U29 ( .A1(\mem[0][1] ), .A2(n695), .ZN(n693) );
  OAI21_X1 U30 ( .B1(n695), .B2(n411), .A(n692), .ZN(n539) );
  NAND2_X1 U31 ( .A1(\mem[0][2] ), .A2(n695), .ZN(n692) );
  OAI21_X1 U32 ( .B1(n695), .B2(n410), .A(n691), .ZN(n538) );
  NAND2_X1 U33 ( .A1(\mem[0][3] ), .A2(n695), .ZN(n691) );
  OAI21_X1 U34 ( .B1(n695), .B2(n409), .A(n690), .ZN(n537) );
  NAND2_X1 U35 ( .A1(\mem[0][4] ), .A2(n695), .ZN(n690) );
  OAI21_X1 U36 ( .B1(n695), .B2(n408), .A(n689), .ZN(n536) );
  NAND2_X1 U37 ( .A1(\mem[0][5] ), .A2(n695), .ZN(n689) );
  OAI21_X1 U38 ( .B1(n695), .B2(n407), .A(n688), .ZN(n535) );
  NAND2_X1 U39 ( .A1(\mem[0][6] ), .A2(n695), .ZN(n688) );
  OAI21_X1 U40 ( .B1(n695), .B2(n406), .A(n687), .ZN(n534) );
  NAND2_X1 U41 ( .A1(\mem[0][7] ), .A2(n695), .ZN(n687) );
  OAI21_X1 U42 ( .B1(n413), .B2(n674), .A(n673), .ZN(n525) );
  NAND2_X1 U43 ( .A1(\mem[2][0] ), .A2(n674), .ZN(n673) );
  OAI21_X1 U44 ( .B1(n412), .B2(n674), .A(n672), .ZN(n524) );
  NAND2_X1 U45 ( .A1(\mem[2][1] ), .A2(n674), .ZN(n672) );
  OAI21_X1 U46 ( .B1(n411), .B2(n674), .A(n671), .ZN(n523) );
  NAND2_X1 U47 ( .A1(\mem[2][2] ), .A2(n674), .ZN(n671) );
  OAI21_X1 U48 ( .B1(n410), .B2(n674), .A(n670), .ZN(n522) );
  NAND2_X1 U49 ( .A1(\mem[2][3] ), .A2(n674), .ZN(n670) );
  OAI21_X1 U50 ( .B1(n409), .B2(n674), .A(n669), .ZN(n521) );
  NAND2_X1 U51 ( .A1(\mem[2][4] ), .A2(n674), .ZN(n669) );
  OAI21_X1 U52 ( .B1(n408), .B2(n674), .A(n668), .ZN(n520) );
  NAND2_X1 U53 ( .A1(\mem[2][5] ), .A2(n674), .ZN(n668) );
  OAI21_X1 U54 ( .B1(n407), .B2(n674), .A(n667), .ZN(n519) );
  NAND2_X1 U55 ( .A1(\mem[2][6] ), .A2(n674), .ZN(n667) );
  OAI21_X1 U56 ( .B1(n406), .B2(n674), .A(n666), .ZN(n518) );
  NAND2_X1 U57 ( .A1(\mem[2][7] ), .A2(n674), .ZN(n666) );
  OAI21_X1 U58 ( .B1(n413), .B2(n664), .A(n663), .ZN(n517) );
  NAND2_X1 U59 ( .A1(\mem[3][0] ), .A2(n664), .ZN(n663) );
  OAI21_X1 U60 ( .B1(n412), .B2(n664), .A(n662), .ZN(n516) );
  NAND2_X1 U61 ( .A1(\mem[3][1] ), .A2(n664), .ZN(n662) );
  OAI21_X1 U62 ( .B1(n411), .B2(n664), .A(n661), .ZN(n515) );
  NAND2_X1 U63 ( .A1(\mem[3][2] ), .A2(n664), .ZN(n661) );
  OAI21_X1 U64 ( .B1(n410), .B2(n664), .A(n660), .ZN(n514) );
  NAND2_X1 U65 ( .A1(\mem[3][3] ), .A2(n664), .ZN(n660) );
  OAI21_X1 U66 ( .B1(n409), .B2(n664), .A(n659), .ZN(n513) );
  NAND2_X1 U67 ( .A1(\mem[3][4] ), .A2(n664), .ZN(n659) );
  OAI21_X1 U68 ( .B1(n408), .B2(n664), .A(n658), .ZN(n512) );
  NAND2_X1 U69 ( .A1(\mem[3][5] ), .A2(n664), .ZN(n658) );
  OAI21_X1 U70 ( .B1(n407), .B2(n664), .A(n657), .ZN(n511) );
  NAND2_X1 U71 ( .A1(\mem[3][6] ), .A2(n664), .ZN(n657) );
  OAI21_X1 U72 ( .B1(n406), .B2(n664), .A(n656), .ZN(n510) );
  NAND2_X1 U73 ( .A1(\mem[3][7] ), .A2(n664), .ZN(n656) );
  NOR2_X1 U74 ( .A1(n405), .A2(N13), .ZN(n626) );
  INV_X1 U75 ( .A(wr_en), .ZN(n405) );
  OAI21_X1 U76 ( .B1(n413), .B2(n684), .A(n683), .ZN(n533) );
  NAND2_X1 U77 ( .A1(\mem[1][0] ), .A2(n684), .ZN(n683) );
  OAI21_X1 U78 ( .B1(n412), .B2(n684), .A(n682), .ZN(n532) );
  NAND2_X1 U79 ( .A1(\mem[1][1] ), .A2(n684), .ZN(n682) );
  OAI21_X1 U80 ( .B1(n411), .B2(n684), .A(n681), .ZN(n531) );
  NAND2_X1 U81 ( .A1(\mem[1][2] ), .A2(n684), .ZN(n681) );
  OAI21_X1 U82 ( .B1(n410), .B2(n684), .A(n680), .ZN(n530) );
  NAND2_X1 U83 ( .A1(\mem[1][3] ), .A2(n684), .ZN(n680) );
  OAI21_X1 U84 ( .B1(n409), .B2(n684), .A(n679), .ZN(n529) );
  NAND2_X1 U85 ( .A1(\mem[1][4] ), .A2(n684), .ZN(n679) );
  OAI21_X1 U86 ( .B1(n408), .B2(n684), .A(n678), .ZN(n528) );
  NAND2_X1 U87 ( .A1(\mem[1][5] ), .A2(n684), .ZN(n678) );
  OAI21_X1 U88 ( .B1(n407), .B2(n684), .A(n677), .ZN(n527) );
  NAND2_X1 U89 ( .A1(\mem[1][6] ), .A2(n684), .ZN(n677) );
  OAI21_X1 U90 ( .B1(n406), .B2(n684), .A(n676), .ZN(n526) );
  NAND2_X1 U91 ( .A1(\mem[1][7] ), .A2(n684), .ZN(n676) );
  OAI21_X1 U92 ( .B1(n413), .B2(n655), .A(n654), .ZN(n509) );
  NAND2_X1 U93 ( .A1(\mem[4][0] ), .A2(n655), .ZN(n654) );
  OAI21_X1 U94 ( .B1(n412), .B2(n655), .A(n653), .ZN(n508) );
  NAND2_X1 U95 ( .A1(\mem[4][1] ), .A2(n655), .ZN(n653) );
  OAI21_X1 U96 ( .B1(n411), .B2(n655), .A(n652), .ZN(n507) );
  NAND2_X1 U97 ( .A1(\mem[4][2] ), .A2(n655), .ZN(n652) );
  OAI21_X1 U98 ( .B1(n410), .B2(n655), .A(n651), .ZN(n506) );
  NAND2_X1 U99 ( .A1(\mem[4][3] ), .A2(n655), .ZN(n651) );
  OAI21_X1 U100 ( .B1(n409), .B2(n655), .A(n650), .ZN(n505) );
  NAND2_X1 U101 ( .A1(\mem[4][4] ), .A2(n655), .ZN(n650) );
  OAI21_X1 U102 ( .B1(n408), .B2(n655), .A(n649), .ZN(n504) );
  NAND2_X1 U103 ( .A1(\mem[4][5] ), .A2(n655), .ZN(n649) );
  OAI21_X1 U104 ( .B1(n407), .B2(n655), .A(n648), .ZN(n503) );
  NAND2_X1 U105 ( .A1(\mem[4][6] ), .A2(n655), .ZN(n648) );
  OAI21_X1 U106 ( .B1(n406), .B2(n655), .A(n647), .ZN(n502) );
  NAND2_X1 U107 ( .A1(\mem[4][7] ), .A2(n655), .ZN(n647) );
  OAI21_X1 U108 ( .B1(n413), .B2(n645), .A(n644), .ZN(n501) );
  NAND2_X1 U109 ( .A1(\mem[5][0] ), .A2(n645), .ZN(n644) );
  OAI21_X1 U110 ( .B1(n412), .B2(n645), .A(n643), .ZN(n500) );
  NAND2_X1 U111 ( .A1(\mem[5][1] ), .A2(n645), .ZN(n643) );
  OAI21_X1 U112 ( .B1(n411), .B2(n645), .A(n642), .ZN(n499) );
  NAND2_X1 U113 ( .A1(\mem[5][2] ), .A2(n645), .ZN(n642) );
  OAI21_X1 U114 ( .B1(n410), .B2(n645), .A(n641), .ZN(n498) );
  NAND2_X1 U115 ( .A1(\mem[5][3] ), .A2(n645), .ZN(n641) );
  OAI21_X1 U116 ( .B1(n409), .B2(n645), .A(n640), .ZN(n497) );
  NAND2_X1 U117 ( .A1(\mem[5][4] ), .A2(n645), .ZN(n640) );
  OAI21_X1 U118 ( .B1(n408), .B2(n645), .A(n639), .ZN(n496) );
  NAND2_X1 U119 ( .A1(\mem[5][5] ), .A2(n645), .ZN(n639) );
  OAI21_X1 U120 ( .B1(n407), .B2(n645), .A(n638), .ZN(n495) );
  NAND2_X1 U121 ( .A1(\mem[5][6] ), .A2(n645), .ZN(n638) );
  OAI21_X1 U122 ( .B1(n406), .B2(n645), .A(n637), .ZN(n494) );
  NAND2_X1 U123 ( .A1(\mem[5][7] ), .A2(n645), .ZN(n637) );
  OAI21_X1 U124 ( .B1(n413), .B2(n636), .A(n635), .ZN(n493) );
  NAND2_X1 U125 ( .A1(\mem[6][0] ), .A2(n636), .ZN(n635) );
  OAI21_X1 U126 ( .B1(n412), .B2(n636), .A(n634), .ZN(n492) );
  NAND2_X1 U127 ( .A1(\mem[6][1] ), .A2(n636), .ZN(n634) );
  OAI21_X1 U128 ( .B1(n411), .B2(n636), .A(n633), .ZN(n491) );
  NAND2_X1 U129 ( .A1(\mem[6][2] ), .A2(n636), .ZN(n633) );
  OAI21_X1 U130 ( .B1(n410), .B2(n636), .A(n632), .ZN(n490) );
  NAND2_X1 U131 ( .A1(\mem[6][3] ), .A2(n636), .ZN(n632) );
  OAI21_X1 U132 ( .B1(n409), .B2(n636), .A(n631), .ZN(n489) );
  NAND2_X1 U133 ( .A1(\mem[6][4] ), .A2(n636), .ZN(n631) );
  OAI21_X1 U134 ( .B1(n408), .B2(n636), .A(n630), .ZN(n488) );
  NAND2_X1 U135 ( .A1(\mem[6][5] ), .A2(n636), .ZN(n630) );
  OAI21_X1 U136 ( .B1(n407), .B2(n636), .A(n629), .ZN(n487) );
  NAND2_X1 U137 ( .A1(\mem[6][6] ), .A2(n636), .ZN(n629) );
  OAI21_X1 U138 ( .B1(n406), .B2(n636), .A(n628), .ZN(n486) );
  NAND2_X1 U139 ( .A1(\mem[6][7] ), .A2(n636), .ZN(n628) );
  OAI21_X1 U140 ( .B1(n413), .B2(n625), .A(n624), .ZN(n485) );
  NAND2_X1 U141 ( .A1(\mem[7][0] ), .A2(n625), .ZN(n624) );
  OAI21_X1 U142 ( .B1(n412), .B2(n625), .A(n623), .ZN(n484) );
  NAND2_X1 U143 ( .A1(\mem[7][1] ), .A2(n625), .ZN(n623) );
  OAI21_X1 U144 ( .B1(n411), .B2(n625), .A(n622), .ZN(n483) );
  NAND2_X1 U145 ( .A1(\mem[7][2] ), .A2(n625), .ZN(n622) );
  OAI21_X1 U146 ( .B1(n410), .B2(n625), .A(n621), .ZN(n482) );
  NAND2_X1 U147 ( .A1(\mem[7][3] ), .A2(n625), .ZN(n621) );
  OAI21_X1 U148 ( .B1(n409), .B2(n625), .A(n620), .ZN(n481) );
  NAND2_X1 U149 ( .A1(\mem[7][4] ), .A2(n625), .ZN(n620) );
  OAI21_X1 U150 ( .B1(n408), .B2(n625), .A(n619), .ZN(n480) );
  NAND2_X1 U151 ( .A1(\mem[7][5] ), .A2(n625), .ZN(n619) );
  OAI21_X1 U152 ( .B1(n407), .B2(n625), .A(n618), .ZN(n479) );
  NAND2_X1 U153 ( .A1(\mem[7][6] ), .A2(n625), .ZN(n618) );
  OAI21_X1 U154 ( .B1(n406), .B2(n625), .A(n617), .ZN(n478) );
  NAND2_X1 U155 ( .A1(\mem[7][7] ), .A2(n625), .ZN(n617) );
  OAI21_X1 U156 ( .B1(n413), .B2(n616), .A(n615), .ZN(n477) );
  NAND2_X1 U157 ( .A1(\mem[8][0] ), .A2(n616), .ZN(n615) );
  OAI21_X1 U158 ( .B1(n412), .B2(n616), .A(n614), .ZN(n476) );
  NAND2_X1 U159 ( .A1(\mem[8][1] ), .A2(n616), .ZN(n614) );
  OAI21_X1 U160 ( .B1(n411), .B2(n616), .A(n613), .ZN(n475) );
  NAND2_X1 U161 ( .A1(\mem[8][2] ), .A2(n616), .ZN(n613) );
  OAI21_X1 U162 ( .B1(n410), .B2(n616), .A(n612), .ZN(n474) );
  NAND2_X1 U163 ( .A1(\mem[8][3] ), .A2(n616), .ZN(n612) );
  OAI21_X1 U164 ( .B1(n409), .B2(n616), .A(n611), .ZN(n473) );
  NAND2_X1 U165 ( .A1(\mem[8][4] ), .A2(n616), .ZN(n611) );
  OAI21_X1 U166 ( .B1(n408), .B2(n616), .A(n610), .ZN(n472) );
  NAND2_X1 U167 ( .A1(\mem[8][5] ), .A2(n616), .ZN(n610) );
  OAI21_X1 U168 ( .B1(n407), .B2(n616), .A(n609), .ZN(n471) );
  NAND2_X1 U169 ( .A1(\mem[8][6] ), .A2(n616), .ZN(n609) );
  OAI21_X1 U170 ( .B1(n406), .B2(n616), .A(n608), .ZN(n470) );
  NAND2_X1 U171 ( .A1(\mem[8][7] ), .A2(n616), .ZN(n608) );
  OAI21_X1 U172 ( .B1(n413), .B2(n606), .A(n605), .ZN(n469) );
  NAND2_X1 U173 ( .A1(\mem[9][0] ), .A2(n606), .ZN(n605) );
  OAI21_X1 U174 ( .B1(n412), .B2(n606), .A(n604), .ZN(n468) );
  NAND2_X1 U175 ( .A1(\mem[9][1] ), .A2(n606), .ZN(n604) );
  OAI21_X1 U176 ( .B1(n411), .B2(n606), .A(n603), .ZN(n467) );
  NAND2_X1 U177 ( .A1(\mem[9][2] ), .A2(n606), .ZN(n603) );
  OAI21_X1 U178 ( .B1(n410), .B2(n606), .A(n602), .ZN(n466) );
  NAND2_X1 U179 ( .A1(\mem[9][3] ), .A2(n606), .ZN(n602) );
  OAI21_X1 U180 ( .B1(n409), .B2(n606), .A(n601), .ZN(n465) );
  NAND2_X1 U181 ( .A1(\mem[9][4] ), .A2(n606), .ZN(n601) );
  OAI21_X1 U182 ( .B1(n408), .B2(n606), .A(n600), .ZN(n464) );
  NAND2_X1 U183 ( .A1(\mem[9][5] ), .A2(n606), .ZN(n600) );
  OAI21_X1 U184 ( .B1(n407), .B2(n606), .A(n599), .ZN(n463) );
  NAND2_X1 U185 ( .A1(\mem[9][6] ), .A2(n606), .ZN(n599) );
  OAI21_X1 U186 ( .B1(n406), .B2(n606), .A(n598), .ZN(n462) );
  NAND2_X1 U187 ( .A1(\mem[9][7] ), .A2(n606), .ZN(n598) );
  OAI21_X1 U188 ( .B1(n413), .B2(n596), .A(n595), .ZN(n461) );
  NAND2_X1 U189 ( .A1(\mem[10][0] ), .A2(n596), .ZN(n595) );
  OAI21_X1 U190 ( .B1(n412), .B2(n596), .A(n594), .ZN(n460) );
  NAND2_X1 U191 ( .A1(\mem[10][1] ), .A2(n596), .ZN(n594) );
  OAI21_X1 U192 ( .B1(n411), .B2(n596), .A(n593), .ZN(n459) );
  NAND2_X1 U193 ( .A1(\mem[10][2] ), .A2(n596), .ZN(n593) );
  OAI21_X1 U194 ( .B1(n410), .B2(n596), .A(n592), .ZN(n458) );
  NAND2_X1 U195 ( .A1(\mem[10][3] ), .A2(n596), .ZN(n592) );
  OAI21_X1 U196 ( .B1(n409), .B2(n596), .A(n591), .ZN(n457) );
  NAND2_X1 U197 ( .A1(\mem[10][4] ), .A2(n596), .ZN(n591) );
  OAI21_X1 U198 ( .B1(n408), .B2(n596), .A(n590), .ZN(n456) );
  NAND2_X1 U199 ( .A1(\mem[10][5] ), .A2(n596), .ZN(n590) );
  OAI21_X1 U200 ( .B1(n407), .B2(n596), .A(n589), .ZN(n455) );
  NAND2_X1 U201 ( .A1(\mem[10][6] ), .A2(n596), .ZN(n589) );
  OAI21_X1 U202 ( .B1(n406), .B2(n596), .A(n588), .ZN(n454) );
  NAND2_X1 U203 ( .A1(\mem[10][7] ), .A2(n596), .ZN(n588) );
  OAI21_X1 U204 ( .B1(n413), .B2(n587), .A(n586), .ZN(n453) );
  NAND2_X1 U205 ( .A1(\mem[11][0] ), .A2(n587), .ZN(n586) );
  OAI21_X1 U206 ( .B1(n412), .B2(n587), .A(n585), .ZN(n452) );
  NAND2_X1 U207 ( .A1(\mem[11][1] ), .A2(n587), .ZN(n585) );
  OAI21_X1 U208 ( .B1(n411), .B2(n587), .A(n584), .ZN(n451) );
  NAND2_X1 U209 ( .A1(\mem[11][2] ), .A2(n587), .ZN(n584) );
  OAI21_X1 U210 ( .B1(n410), .B2(n587), .A(n583), .ZN(n450) );
  NAND2_X1 U211 ( .A1(\mem[11][3] ), .A2(n587), .ZN(n583) );
  OAI21_X1 U212 ( .B1(n409), .B2(n587), .A(n582), .ZN(n449) );
  NAND2_X1 U213 ( .A1(\mem[11][4] ), .A2(n587), .ZN(n582) );
  OAI21_X1 U214 ( .B1(n408), .B2(n587), .A(n581), .ZN(n448) );
  NAND2_X1 U215 ( .A1(\mem[11][5] ), .A2(n587), .ZN(n581) );
  OAI21_X1 U216 ( .B1(n407), .B2(n587), .A(n580), .ZN(n447) );
  NAND2_X1 U217 ( .A1(\mem[11][6] ), .A2(n587), .ZN(n580) );
  OAI21_X1 U218 ( .B1(n406), .B2(n587), .A(n579), .ZN(n446) );
  NAND2_X1 U219 ( .A1(\mem[11][7] ), .A2(n587), .ZN(n579) );
  OAI21_X1 U220 ( .B1(n413), .B2(n578), .A(n577), .ZN(n445) );
  NAND2_X1 U221 ( .A1(\mem[12][0] ), .A2(n578), .ZN(n577) );
  OAI21_X1 U222 ( .B1(n412), .B2(n578), .A(n576), .ZN(n444) );
  NAND2_X1 U223 ( .A1(\mem[12][1] ), .A2(n578), .ZN(n576) );
  OAI21_X1 U224 ( .B1(n411), .B2(n578), .A(n575), .ZN(n443) );
  NAND2_X1 U225 ( .A1(\mem[12][2] ), .A2(n578), .ZN(n575) );
  OAI21_X1 U226 ( .B1(n410), .B2(n578), .A(n574), .ZN(n442) );
  NAND2_X1 U227 ( .A1(\mem[12][3] ), .A2(n578), .ZN(n574) );
  OAI21_X1 U228 ( .B1(n409), .B2(n578), .A(n573), .ZN(n441) );
  NAND2_X1 U229 ( .A1(\mem[12][4] ), .A2(n578), .ZN(n573) );
  OAI21_X1 U230 ( .B1(n408), .B2(n578), .A(n572), .ZN(n440) );
  NAND2_X1 U231 ( .A1(\mem[12][5] ), .A2(n578), .ZN(n572) );
  OAI21_X1 U232 ( .B1(n407), .B2(n578), .A(n571), .ZN(n439) );
  NAND2_X1 U233 ( .A1(\mem[12][6] ), .A2(n578), .ZN(n571) );
  OAI21_X1 U234 ( .B1(n406), .B2(n578), .A(n570), .ZN(n438) );
  NAND2_X1 U235 ( .A1(\mem[12][7] ), .A2(n578), .ZN(n570) );
  OAI21_X1 U236 ( .B1(n413), .B2(n569), .A(n568), .ZN(n437) );
  NAND2_X1 U237 ( .A1(\mem[13][0] ), .A2(n569), .ZN(n568) );
  OAI21_X1 U238 ( .B1(n412), .B2(n569), .A(n567), .ZN(n436) );
  NAND2_X1 U239 ( .A1(\mem[13][1] ), .A2(n569), .ZN(n567) );
  OAI21_X1 U240 ( .B1(n411), .B2(n569), .A(n566), .ZN(n435) );
  NAND2_X1 U241 ( .A1(\mem[13][2] ), .A2(n569), .ZN(n566) );
  OAI21_X1 U242 ( .B1(n410), .B2(n569), .A(n565), .ZN(n434) );
  NAND2_X1 U243 ( .A1(\mem[13][3] ), .A2(n569), .ZN(n565) );
  OAI21_X1 U244 ( .B1(n409), .B2(n569), .A(n564), .ZN(n433) );
  NAND2_X1 U245 ( .A1(\mem[13][4] ), .A2(n569), .ZN(n564) );
  OAI21_X1 U246 ( .B1(n408), .B2(n569), .A(n563), .ZN(n432) );
  NAND2_X1 U247 ( .A1(\mem[13][5] ), .A2(n569), .ZN(n563) );
  OAI21_X1 U248 ( .B1(n407), .B2(n569), .A(n562), .ZN(n431) );
  NAND2_X1 U249 ( .A1(\mem[13][6] ), .A2(n569), .ZN(n562) );
  OAI21_X1 U250 ( .B1(n406), .B2(n569), .A(n561), .ZN(n430) );
  NAND2_X1 U251 ( .A1(\mem[13][7] ), .A2(n569), .ZN(n561) );
  OAI21_X1 U252 ( .B1(n413), .B2(n560), .A(n559), .ZN(n429) );
  NAND2_X1 U253 ( .A1(\mem[14][0] ), .A2(n560), .ZN(n559) );
  OAI21_X1 U254 ( .B1(n412), .B2(n560), .A(n558), .ZN(n428) );
  NAND2_X1 U255 ( .A1(\mem[14][1] ), .A2(n560), .ZN(n558) );
  OAI21_X1 U256 ( .B1(n411), .B2(n560), .A(n557), .ZN(n427) );
  NAND2_X1 U257 ( .A1(\mem[14][2] ), .A2(n560), .ZN(n557) );
  OAI21_X1 U258 ( .B1(n410), .B2(n560), .A(n556), .ZN(n426) );
  NAND2_X1 U259 ( .A1(\mem[14][3] ), .A2(n560), .ZN(n556) );
  OAI21_X1 U260 ( .B1(n409), .B2(n560), .A(n555), .ZN(n425) );
  NAND2_X1 U261 ( .A1(\mem[14][4] ), .A2(n560), .ZN(n555) );
  OAI21_X1 U262 ( .B1(n408), .B2(n560), .A(n554), .ZN(n424) );
  NAND2_X1 U263 ( .A1(\mem[14][5] ), .A2(n560), .ZN(n554) );
  OAI21_X1 U264 ( .B1(n407), .B2(n560), .A(n553), .ZN(n423) );
  NAND2_X1 U265 ( .A1(\mem[14][6] ), .A2(n560), .ZN(n553) );
  OAI21_X1 U266 ( .B1(n406), .B2(n560), .A(n552), .ZN(n422) );
  NAND2_X1 U267 ( .A1(\mem[14][7] ), .A2(n560), .ZN(n552) );
  OAI21_X1 U268 ( .B1(n413), .B2(n550), .A(n549), .ZN(n421) );
  NAND2_X1 U269 ( .A1(\mem[15][0] ), .A2(n550), .ZN(n549) );
  OAI21_X1 U270 ( .B1(n412), .B2(n550), .A(n548), .ZN(n420) );
  NAND2_X1 U271 ( .A1(\mem[15][1] ), .A2(n550), .ZN(n548) );
  OAI21_X1 U272 ( .B1(n411), .B2(n550), .A(n547), .ZN(n419) );
  NAND2_X1 U273 ( .A1(\mem[15][2] ), .A2(n550), .ZN(n547) );
  OAI21_X1 U274 ( .B1(n410), .B2(n550), .A(n546), .ZN(n418) );
  NAND2_X1 U275 ( .A1(\mem[15][3] ), .A2(n550), .ZN(n546) );
  OAI21_X1 U276 ( .B1(n409), .B2(n550), .A(n545), .ZN(n417) );
  NAND2_X1 U277 ( .A1(\mem[15][4] ), .A2(n550), .ZN(n545) );
  OAI21_X1 U278 ( .B1(n408), .B2(n550), .A(n544), .ZN(n416) );
  NAND2_X1 U279 ( .A1(\mem[15][5] ), .A2(n550), .ZN(n544) );
  OAI21_X1 U280 ( .B1(n407), .B2(n550), .A(n543), .ZN(n415) );
  NAND2_X1 U281 ( .A1(\mem[15][6] ), .A2(n550), .ZN(n543) );
  OAI21_X1 U282 ( .B1(n406), .B2(n550), .A(n542), .ZN(n414) );
  NAND2_X1 U283 ( .A1(\mem[15][7] ), .A2(n550), .ZN(n542) );
  AND2_X1 U284 ( .A1(N13), .A2(wr_en), .ZN(n551) );
  NOR2_X1 U285 ( .A1(N11), .A2(N12), .ZN(n686) );
  NOR2_X1 U286 ( .A1(n404), .A2(N12), .ZN(n665) );
  AND2_X1 U287 ( .A1(N12), .A2(n404), .ZN(n646) );
  AND2_X1 U288 ( .A1(N12), .A2(N11), .ZN(n627) );
  INV_X1 U289 ( .A(data_in[0]), .ZN(n413) );
  INV_X1 U290 ( .A(data_in[1]), .ZN(n412) );
  INV_X1 U291 ( .A(data_in[2]), .ZN(n411) );
  INV_X1 U292 ( .A(data_in[3]), .ZN(n410) );
  INV_X1 U293 ( .A(data_in[4]), .ZN(n409) );
  INV_X1 U294 ( .A(data_in[5]), .ZN(n408) );
  INV_X1 U295 ( .A(data_in[6]), .ZN(n407) );
  INV_X1 U296 ( .A(data_in[7]), .ZN(n406) );
  MUX2_X1 U297 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n398), .Z(n3) );
  MUX2_X1 U298 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n398), .Z(n4) );
  MUX2_X1 U299 ( .A(n4), .B(n3), .S(n397), .Z(n5) );
  MUX2_X1 U300 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n398), .Z(n6) );
  MUX2_X1 U301 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n398), .Z(n7) );
  MUX2_X1 U302 ( .A(n7), .B(n6), .S(n397), .Z(n8) );
  MUX2_X1 U303 ( .A(n8), .B(n5), .S(N12), .Z(n9) );
  MUX2_X1 U304 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n400), .Z(n10) );
  MUX2_X1 U305 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n399), .Z(n11) );
  MUX2_X1 U306 ( .A(n11), .B(n10), .S(n397), .Z(n294) );
  MUX2_X1 U307 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n398), .Z(n295) );
  MUX2_X1 U308 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n400), .Z(n296) );
  MUX2_X1 U309 ( .A(n296), .B(n295), .S(n397), .Z(n297) );
  MUX2_X1 U310 ( .A(n297), .B(n294), .S(N12), .Z(n298) );
  MUX2_X1 U311 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n399), .Z(n299) );
  MUX2_X1 U312 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n398), .Z(n300) );
  MUX2_X1 U313 ( .A(n300), .B(n299), .S(n397), .Z(n301) );
  MUX2_X1 U314 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(N10), .Z(n302) );
  MUX2_X1 U315 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n398), .Z(n303) );
  MUX2_X1 U316 ( .A(n303), .B(n302), .S(n397), .Z(n304) );
  MUX2_X1 U317 ( .A(n304), .B(n301), .S(N12), .Z(n305) );
  MUX2_X1 U318 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(N10), .Z(n306) );
  MUX2_X1 U319 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n400), .Z(n307) );
  MUX2_X1 U320 ( .A(n307), .B(n306), .S(n397), .Z(n308) );
  MUX2_X1 U321 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n399), .Z(n309) );
  MUX2_X1 U322 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n399), .Z(n310) );
  MUX2_X1 U323 ( .A(n310), .B(n309), .S(n397), .Z(n311) );
  MUX2_X1 U324 ( .A(n311), .B(n308), .S(N12), .Z(n312) );
  MUX2_X1 U325 ( .A(n312), .B(n305), .S(N13), .Z(N20) );
  MUX2_X1 U326 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n400), .Z(n313) );
  MUX2_X1 U327 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(N10), .Z(n314) );
  MUX2_X1 U328 ( .A(n314), .B(n313), .S(n397), .Z(n315) );
  MUX2_X1 U329 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(N10), .Z(n316) );
  MUX2_X1 U330 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(N10), .Z(n317) );
  MUX2_X1 U331 ( .A(n317), .B(n316), .S(N11), .Z(n318) );
  MUX2_X1 U332 ( .A(n318), .B(n315), .S(N12), .Z(n319) );
  MUX2_X1 U333 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n400), .Z(n320) );
  MUX2_X1 U334 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(N10), .Z(n321) );
  MUX2_X1 U335 ( .A(n321), .B(n320), .S(n397), .Z(n322) );
  MUX2_X1 U336 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(N10), .Z(n323) );
  MUX2_X1 U337 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(N10), .Z(n324) );
  MUX2_X1 U338 ( .A(n324), .B(n323), .S(N11), .Z(n325) );
  MUX2_X1 U339 ( .A(n325), .B(n322), .S(N12), .Z(n326) );
  MUX2_X1 U340 ( .A(n326), .B(n319), .S(N13), .Z(N19) );
  MUX2_X1 U341 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n399), .Z(n327) );
  MUX2_X1 U342 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(N10), .Z(n328) );
  MUX2_X1 U343 ( .A(n328), .B(n327), .S(n397), .Z(n329) );
  MUX2_X1 U344 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(N10), .Z(n330) );
  MUX2_X1 U345 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n331) );
  MUX2_X1 U346 ( .A(n331), .B(n330), .S(N11), .Z(n332) );
  MUX2_X1 U347 ( .A(n332), .B(n329), .S(N12), .Z(n333) );
  MUX2_X1 U348 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n398), .Z(n334) );
  MUX2_X1 U349 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n335) );
  MUX2_X1 U350 ( .A(n335), .B(n334), .S(N11), .Z(n336) );
  MUX2_X1 U351 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n398), .Z(n337) );
  MUX2_X1 U352 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n338) );
  MUX2_X1 U353 ( .A(n338), .B(n337), .S(N11), .Z(n339) );
  MUX2_X1 U354 ( .A(n339), .B(n336), .S(N12), .Z(n340) );
  MUX2_X1 U355 ( .A(n340), .B(n333), .S(N13), .Z(N18) );
  MUX2_X1 U356 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n398), .Z(n341) );
  MUX2_X1 U357 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n398), .Z(n342) );
  MUX2_X1 U358 ( .A(n342), .B(n341), .S(n397), .Z(n343) );
  MUX2_X1 U359 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n398), .Z(n344) );
  MUX2_X1 U360 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(N10), .Z(n345) );
  MUX2_X1 U361 ( .A(n345), .B(n344), .S(N11), .Z(n346) );
  MUX2_X1 U362 ( .A(n346), .B(n343), .S(N12), .Z(n347) );
  MUX2_X1 U363 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n398), .Z(n348) );
  MUX2_X1 U364 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(N10), .Z(n349) );
  MUX2_X1 U365 ( .A(n349), .B(n348), .S(N11), .Z(n350) );
  MUX2_X1 U366 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n398), .Z(n351) );
  MUX2_X1 U367 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n352) );
  MUX2_X1 U368 ( .A(n352), .B(n351), .S(N11), .Z(n353) );
  MUX2_X1 U369 ( .A(n353), .B(n350), .S(N12), .Z(n354) );
  MUX2_X1 U370 ( .A(n354), .B(n347), .S(N13), .Z(N17) );
  MUX2_X1 U371 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n399), .Z(n355) );
  MUX2_X1 U372 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n399), .Z(n356) );
  MUX2_X1 U373 ( .A(n356), .B(n355), .S(N11), .Z(n357) );
  MUX2_X1 U374 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n399), .Z(n358) );
  MUX2_X1 U375 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n399), .Z(n359) );
  MUX2_X1 U376 ( .A(n359), .B(n358), .S(N11), .Z(n360) );
  MUX2_X1 U377 ( .A(n360), .B(n357), .S(N12), .Z(n361) );
  MUX2_X1 U378 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n399), .Z(n362) );
  MUX2_X1 U379 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n399), .Z(n363) );
  MUX2_X1 U380 ( .A(n363), .B(n362), .S(n397), .Z(n364) );
  MUX2_X1 U381 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n399), .Z(n365) );
  MUX2_X1 U382 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n399), .Z(n366) );
  MUX2_X1 U383 ( .A(n366), .B(n365), .S(n397), .Z(n367) );
  MUX2_X1 U384 ( .A(n367), .B(n364), .S(N12), .Z(n368) );
  MUX2_X1 U385 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n399), .Z(n369) );
  MUX2_X1 U386 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n399), .Z(n370) );
  MUX2_X1 U387 ( .A(n370), .B(n369), .S(N11), .Z(n371) );
  MUX2_X1 U388 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n399), .Z(n372) );
  MUX2_X1 U389 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n399), .Z(n373) );
  MUX2_X1 U390 ( .A(n373), .B(n372), .S(N11), .Z(n374) );
  MUX2_X1 U391 ( .A(n374), .B(n371), .S(N12), .Z(n375) );
  MUX2_X1 U392 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n400), .Z(n376) );
  MUX2_X1 U393 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n400), .Z(n377) );
  MUX2_X1 U394 ( .A(n377), .B(n376), .S(N11), .Z(n378) );
  MUX2_X1 U395 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n400), .Z(n379) );
  MUX2_X1 U396 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n400), .Z(n380) );
  MUX2_X1 U397 ( .A(n380), .B(n379), .S(N11), .Z(n381) );
  MUX2_X1 U398 ( .A(n381), .B(n378), .S(N12), .Z(n382) );
  MUX2_X1 U399 ( .A(n382), .B(n375), .S(N13), .Z(N15) );
  MUX2_X1 U400 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n400), .Z(n383) );
  MUX2_X1 U401 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n400), .Z(n384) );
  MUX2_X1 U402 ( .A(n384), .B(n383), .S(N11), .Z(n385) );
  MUX2_X1 U403 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n400), .Z(n386) );
  MUX2_X1 U404 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n400), .Z(n387) );
  MUX2_X1 U405 ( .A(n387), .B(n386), .S(N11), .Z(n388) );
  MUX2_X1 U406 ( .A(n388), .B(n385), .S(N12), .Z(n389) );
  MUX2_X1 U407 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n400), .Z(n390) );
  MUX2_X1 U408 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n400), .Z(n391) );
  MUX2_X1 U409 ( .A(n391), .B(n390), .S(N11), .Z(n392) );
  MUX2_X1 U410 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n400), .Z(n393) );
  MUX2_X1 U411 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n400), .Z(n394) );
  MUX2_X1 U412 ( .A(n394), .B(n393), .S(N11), .Z(n395) );
  MUX2_X1 U413 ( .A(n395), .B(n392), .S(N12), .Z(n396) );
  MUX2_X1 U414 ( .A(n396), .B(n389), .S(N13), .Z(N14) );
  CLKBUF_X1 U415 ( .A(N10), .Z(n398) );
  INV_X2 U416 ( .A(n401), .ZN(data_out[1]) );
  INV_X1 U417 ( .A(N10), .ZN(n403) );
  INV_X1 U418 ( .A(N11), .ZN(n404) );
endmodule


module memory_WIDTH16_SIZE16_LOGSIZE4 ( clk, data_in, data_out, addr, wr_en );
  input [15:0] data_in;
  output [15:0] data_out;
  input [3:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, \mem[15][15] , \mem[15][14] , \mem[15][13] ,
         \mem[15][12] , \mem[15][11] , \mem[15][10] , \mem[15][9] ,
         \mem[15][8] , \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] ,
         \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][15] ,
         \mem[14][14] , \mem[14][13] , \mem[14][12] , \mem[14][11] ,
         \mem[14][10] , \mem[14][9] , \mem[14][8] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][15] , \mem[13][14] , \mem[13][13] ,
         \mem[13][12] , \mem[13][11] , \mem[13][10] , \mem[13][9] ,
         \mem[13][8] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][15] ,
         \mem[12][14] , \mem[12][13] , \mem[12][12] , \mem[12][11] ,
         \mem[12][10] , \mem[12][9] , \mem[12][8] , \mem[12][7] , \mem[12][6] ,
         \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] , \mem[12][1] ,
         \mem[12][0] , \mem[11][15] , \mem[11][14] , \mem[11][13] ,
         \mem[11][12] , \mem[11][11] , \mem[11][10] , \mem[11][9] ,
         \mem[11][8] , \mem[11][7] , \mem[11][6] , \mem[11][5] , \mem[11][4] ,
         \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] , \mem[10][15] ,
         \mem[10][14] , \mem[10][13] , \mem[10][12] , \mem[10][11] ,
         \mem[10][10] , \mem[10][9] , \mem[10][8] , \mem[10][7] , \mem[10][6] ,
         \mem[10][5] , \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] ,
         \mem[10][0] , \mem[9][15] , \mem[9][14] , \mem[9][13] , \mem[9][12] ,
         \mem[9][11] , \mem[9][10] , \mem[9][9] , \mem[9][8] , \mem[9][7] ,
         \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] ,
         \mem[9][1] , \mem[9][0] , \mem[8][15] , \mem[8][14] , \mem[8][13] ,
         \mem[8][12] , \mem[8][11] , \mem[8][10] , \mem[8][9] , \mem[8][8] ,
         \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] , \mem[8][3] ,
         \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][15] , \mem[7][14] ,
         \mem[7][13] , \mem[7][12] , \mem[7][11] , \mem[7][10] , \mem[7][9] ,
         \mem[7][8] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][15] ,
         \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] ,
         \mem[4][11] , \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] ,
         \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] ,
         \mem[4][1] , \mem[4][0] , \mem[3][15] , \mem[3][14] , \mem[3][13] ,
         \mem[3][12] , \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] ,
         \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] ,
         \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][15] , \mem[2][14] ,
         \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] ,
         \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][15] ,
         \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24,
         N25, N26, N27, N28, N29, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];

  DFF_X1 \data_out_reg[15]  ( .D(N14), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N15), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(N16), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(N17), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(N18), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N19), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N20), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N21), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N22), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N23), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N24), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N25), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N26), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N27), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N28), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N29), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[15][15]  ( .D(n557), .CK(clk), .Q(\mem[15][15] ) );
  DFF_X1 \mem_reg[15][14]  ( .D(n556), .CK(clk), .Q(\mem[15][14] ) );
  DFF_X1 \mem_reg[15][13]  ( .D(n555), .CK(clk), .Q(\mem[15][13] ) );
  DFF_X1 \mem_reg[15][12]  ( .D(n554), .CK(clk), .Q(\mem[15][12] ) );
  DFF_X1 \mem_reg[15][11]  ( .D(n553), .CK(clk), .Q(\mem[15][11] ) );
  DFF_X1 \mem_reg[15][10]  ( .D(n552), .CK(clk), .Q(\mem[15][10] ) );
  DFF_X1 \mem_reg[15][9]  ( .D(n551), .CK(clk), .Q(\mem[15][9] ) );
  DFF_X1 \mem_reg[15][8]  ( .D(n550), .CK(clk), .Q(\mem[15][8] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n549), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n548), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n547), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n546), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n545), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n544), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n543), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n542), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][15]  ( .D(n541), .CK(clk), .Q(\mem[14][15] ) );
  DFF_X1 \mem_reg[14][14]  ( .D(n540), .CK(clk), .Q(\mem[14][14] ) );
  DFF_X1 \mem_reg[14][13]  ( .D(n539), .CK(clk), .Q(\mem[14][13] ) );
  DFF_X1 \mem_reg[14][12]  ( .D(n538), .CK(clk), .Q(\mem[14][12] ) );
  DFF_X1 \mem_reg[14][11]  ( .D(n537), .CK(clk), .Q(\mem[14][11] ) );
  DFF_X1 \mem_reg[14][10]  ( .D(n536), .CK(clk), .Q(\mem[14][10] ) );
  DFF_X1 \mem_reg[14][9]  ( .D(n535), .CK(clk), .Q(\mem[14][9] ) );
  DFF_X1 \mem_reg[14][8]  ( .D(n534), .CK(clk), .Q(\mem[14][8] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n533), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n532), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n531), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n530), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n529), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n528), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n527), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n526), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][15]  ( .D(n525), .CK(clk), .Q(\mem[13][15] ) );
  DFF_X1 \mem_reg[13][14]  ( .D(n524), .CK(clk), .Q(\mem[13][14] ) );
  DFF_X1 \mem_reg[13][13]  ( .D(n523), .CK(clk), .Q(\mem[13][13] ) );
  DFF_X1 \mem_reg[13][12]  ( .D(n522), .CK(clk), .Q(\mem[13][12] ) );
  DFF_X1 \mem_reg[13][11]  ( .D(n521), .CK(clk), .Q(\mem[13][11] ) );
  DFF_X1 \mem_reg[13][10]  ( .D(n520), .CK(clk), .Q(\mem[13][10] ) );
  DFF_X1 \mem_reg[13][9]  ( .D(n519), .CK(clk), .Q(\mem[13][9] ) );
  DFF_X1 \mem_reg[13][8]  ( .D(n518), .CK(clk), .Q(\mem[13][8] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n517), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n516), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n515), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n514), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n513), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n512), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n511), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n510), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][15]  ( .D(n509), .CK(clk), .Q(\mem[12][15] ) );
  DFF_X1 \mem_reg[12][14]  ( .D(n508), .CK(clk), .Q(\mem[12][14] ) );
  DFF_X1 \mem_reg[12][13]  ( .D(n507), .CK(clk), .Q(\mem[12][13] ) );
  DFF_X1 \mem_reg[12][12]  ( .D(n506), .CK(clk), .Q(\mem[12][12] ) );
  DFF_X1 \mem_reg[12][11]  ( .D(n505), .CK(clk), .Q(\mem[12][11] ) );
  DFF_X1 \mem_reg[12][10]  ( .D(n504), .CK(clk), .Q(\mem[12][10] ) );
  DFF_X1 \mem_reg[12][9]  ( .D(n503), .CK(clk), .Q(\mem[12][9] ) );
  DFF_X1 \mem_reg[12][8]  ( .D(n502), .CK(clk), .Q(\mem[12][8] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n501), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n500), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n499), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n498), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n497), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n496), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n495), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n494), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][15]  ( .D(n493), .CK(clk), .Q(\mem[11][15] ) );
  DFF_X1 \mem_reg[11][14]  ( .D(n492), .CK(clk), .Q(\mem[11][14] ) );
  DFF_X1 \mem_reg[11][13]  ( .D(n491), .CK(clk), .Q(\mem[11][13] ) );
  DFF_X1 \mem_reg[11][12]  ( .D(n490), .CK(clk), .Q(\mem[11][12] ) );
  DFF_X1 \mem_reg[11][11]  ( .D(n489), .CK(clk), .Q(\mem[11][11] ) );
  DFF_X1 \mem_reg[11][10]  ( .D(n488), .CK(clk), .Q(\mem[11][10] ) );
  DFF_X1 \mem_reg[11][9]  ( .D(n487), .CK(clk), .Q(\mem[11][9] ) );
  DFF_X1 \mem_reg[11][8]  ( .D(n486), .CK(clk), .Q(\mem[11][8] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n485), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n484), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n483), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n482), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n481), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n480), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n479), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n478), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][15]  ( .D(n477), .CK(clk), .Q(\mem[10][15] ) );
  DFF_X1 \mem_reg[10][14]  ( .D(n476), .CK(clk), .Q(\mem[10][14] ) );
  DFF_X1 \mem_reg[10][13]  ( .D(n475), .CK(clk), .Q(\mem[10][13] ) );
  DFF_X1 \mem_reg[10][12]  ( .D(n474), .CK(clk), .Q(\mem[10][12] ) );
  DFF_X1 \mem_reg[10][11]  ( .D(n473), .CK(clk), .Q(\mem[10][11] ) );
  DFF_X1 \mem_reg[10][10]  ( .D(n472), .CK(clk), .Q(\mem[10][10] ) );
  DFF_X1 \mem_reg[10][9]  ( .D(n471), .CK(clk), .Q(\mem[10][9] ) );
  DFF_X1 \mem_reg[10][8]  ( .D(n470), .CK(clk), .Q(\mem[10][8] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n469), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n468), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n467), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n466), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n465), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n464), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n463), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n462), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][15]  ( .D(n461), .CK(clk), .Q(\mem[9][15] ) );
  DFF_X1 \mem_reg[9][14]  ( .D(n460), .CK(clk), .Q(\mem[9][14] ) );
  DFF_X1 \mem_reg[9][13]  ( .D(n459), .CK(clk), .Q(\mem[9][13] ) );
  DFF_X1 \mem_reg[9][12]  ( .D(n458), .CK(clk), .Q(\mem[9][12] ) );
  DFF_X1 \mem_reg[9][11]  ( .D(n457), .CK(clk), .Q(\mem[9][11] ) );
  DFF_X1 \mem_reg[9][10]  ( .D(n456), .CK(clk), .Q(\mem[9][10] ) );
  DFF_X1 \mem_reg[9][9]  ( .D(n455), .CK(clk), .Q(\mem[9][9] ) );
  DFF_X1 \mem_reg[9][8]  ( .D(n454), .CK(clk), .Q(\mem[9][8] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n453), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n452), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n451), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n450), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n449), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n448), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n447), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n446), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][15]  ( .D(n445), .CK(clk), .Q(\mem[8][15] ) );
  DFF_X1 \mem_reg[8][14]  ( .D(n444), .CK(clk), .Q(\mem[8][14] ) );
  DFF_X1 \mem_reg[8][13]  ( .D(n443), .CK(clk), .Q(\mem[8][13] ) );
  DFF_X1 \mem_reg[8][12]  ( .D(n442), .CK(clk), .Q(\mem[8][12] ) );
  DFF_X1 \mem_reg[8][11]  ( .D(n441), .CK(clk), .Q(\mem[8][11] ) );
  DFF_X1 \mem_reg[8][10]  ( .D(n440), .CK(clk), .Q(\mem[8][10] ) );
  DFF_X1 \mem_reg[8][9]  ( .D(n439), .CK(clk), .Q(\mem[8][9] ) );
  DFF_X1 \mem_reg[8][8]  ( .D(n438), .CK(clk), .Q(\mem[8][8] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n437), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n436), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n435), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n434), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n433), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n432), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n431), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n430), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n429), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n428), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n427), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n426), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n425), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n424), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n423), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n422), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n421), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n420), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n419), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n418), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n417), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n416), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n415), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n414), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n413), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n412), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n411), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n410), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n409), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n408), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n407), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n406), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n405), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n404), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n403), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n402), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n401), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n400), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n399), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n398), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n397), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n396), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n395), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n394), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n393), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n392), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n391), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n390), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n389), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n388), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n387), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n386), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n385), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n384), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n383), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n382), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n381), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n380), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n379), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n378), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n377), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n376), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n375), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n374), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n373), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n372), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n371), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n370), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n369), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n368), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n367), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n366), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n365), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n364), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n363), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n362), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n361), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n360), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n359), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n358), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n357), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n356), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n355), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n354), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n353), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n352), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n351), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n350), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n349), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n348), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n347), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n346), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n345), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n344), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n343), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n342), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n341), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n340), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n339), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n338), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n337), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n336), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n335), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n334), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n333), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n332), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n331), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n330), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n329), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n328), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n327), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n326), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n325), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n324), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n323), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n322), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n321), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n320), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n319), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n318), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n317), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n316), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n315), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n314), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n313), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n312), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n311), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n310), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n309), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n308), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n307), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n306), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n305), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n304), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n303), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n302), .CK(clk), .Q(\mem[0][0] ) );
  BUF_X1 U3 ( .A(N11), .Z(n764) );
  BUF_X1 U4 ( .A(N11), .Z(n765) );
  BUF_X1 U5 ( .A(N11), .Z(n766) );
  BUF_X1 U6 ( .A(n772), .Z(n770) );
  BUF_X1 U7 ( .A(n772), .Z(n771) );
  BUF_X1 U8 ( .A(n772), .Z(n768) );
  BUF_X1 U9 ( .A(n772), .Z(n769) );
  BUF_X1 U10 ( .A(n20), .Z(n788) );
  BUF_X1 U11 ( .A(n39), .Z(n787) );
  BUF_X1 U12 ( .A(n181), .Z(n779) );
  BUF_X1 U13 ( .A(n199), .Z(n778) );
  BUF_X1 U14 ( .A(n57), .Z(n786) );
  BUF_X1 U15 ( .A(n75), .Z(n785) );
  BUF_X1 U16 ( .A(n127), .Z(n782) );
  BUF_X1 U17 ( .A(n146), .Z(n781) );
  BUF_X1 U18 ( .A(n233), .Z(n776) );
  BUF_X1 U19 ( .A(n250), .Z(n775) );
  BUF_X1 U20 ( .A(n267), .Z(n774) );
  BUF_X1 U21 ( .A(n285), .Z(n773) );
  BUF_X1 U22 ( .A(n92), .Z(n784) );
  BUF_X1 U23 ( .A(n110), .Z(n783) );
  BUF_X1 U24 ( .A(n163), .Z(n780) );
  BUF_X1 U25 ( .A(n216), .Z(n777) );
  BUF_X1 U26 ( .A(N10), .Z(n772) );
  AND2_X1 U27 ( .A1(n145), .A2(n789), .ZN(n38) );
  AND2_X1 U28 ( .A1(N10), .A2(n145), .ZN(n56) );
  AND2_X1 U29 ( .A1(n284), .A2(N10), .ZN(n198) );
  AND2_X1 U30 ( .A1(n284), .A2(n789), .ZN(n180) );
  NAND2_X1 U31 ( .A1(n56), .A2(n37), .ZN(n39) );
  NAND2_X1 U32 ( .A1(n180), .A2(n37), .ZN(n163) );
  NAND2_X1 U33 ( .A1(n198), .A2(n37), .ZN(n181) );
  NAND2_X1 U34 ( .A1(n180), .A2(n74), .ZN(n199) );
  NAND2_X1 U35 ( .A1(n198), .A2(n74), .ZN(n216) );
  NAND2_X1 U36 ( .A1(n37), .A2(n38), .ZN(n20) );
  NAND2_X1 U37 ( .A1(n74), .A2(n38), .ZN(n57) );
  NAND2_X1 U38 ( .A1(n74), .A2(n56), .ZN(n75) );
  NAND2_X1 U39 ( .A1(n180), .A2(n109), .ZN(n233) );
  NAND2_X1 U40 ( .A1(n198), .A2(n109), .ZN(n250) );
  NAND2_X1 U41 ( .A1(n180), .A2(n144), .ZN(n267) );
  NAND2_X1 U42 ( .A1(n198), .A2(n144), .ZN(n285) );
  NAND2_X1 U43 ( .A1(n109), .A2(n38), .ZN(n92) );
  NAND2_X1 U44 ( .A1(n109), .A2(n56), .ZN(n110) );
  NAND2_X1 U45 ( .A1(n144), .A2(n38), .ZN(n127) );
  NAND2_X1 U46 ( .A1(n144), .A2(n56), .ZN(n146) );
  NOR2_X1 U47 ( .A1(N11), .A2(N12), .ZN(n37) );
  NOR2_X1 U48 ( .A1(n791), .A2(N13), .ZN(n145) );
  INV_X1 U49 ( .A(wr_en), .ZN(n791) );
  AND2_X1 U50 ( .A1(N12), .A2(N11), .ZN(n144) );
  OAI21_X1 U51 ( .B1(n800), .B2(n57), .A(n65), .ZN(n341) );
  NAND2_X1 U52 ( .A1(\mem[2][7] ), .A2(n786), .ZN(n65) );
  OAI21_X1 U53 ( .B1(n799), .B2(n786), .A(n66), .ZN(n342) );
  NAND2_X1 U54 ( .A1(\mem[2][8] ), .A2(n786), .ZN(n66) );
  OAI21_X1 U55 ( .B1(n798), .B2(n57), .A(n67), .ZN(n343) );
  NAND2_X1 U56 ( .A1(\mem[2][9] ), .A2(n786), .ZN(n67) );
  OAI21_X1 U57 ( .B1(n797), .B2(n57), .A(n68), .ZN(n344) );
  NAND2_X1 U58 ( .A1(\mem[2][10] ), .A2(n786), .ZN(n68) );
  OAI21_X1 U59 ( .B1(n796), .B2(n57), .A(n69), .ZN(n345) );
  NAND2_X1 U60 ( .A1(\mem[2][11] ), .A2(n786), .ZN(n69) );
  OAI21_X1 U61 ( .B1(n795), .B2(n57), .A(n70), .ZN(n346) );
  NAND2_X1 U62 ( .A1(\mem[2][12] ), .A2(n786), .ZN(n70) );
  OAI21_X1 U63 ( .B1(n794), .B2(n57), .A(n71), .ZN(n347) );
  NAND2_X1 U64 ( .A1(\mem[2][13] ), .A2(n786), .ZN(n71) );
  OAI21_X1 U65 ( .B1(n793), .B2(n57), .A(n72), .ZN(n348) );
  NAND2_X1 U66 ( .A1(\mem[2][14] ), .A2(n786), .ZN(n72) );
  OAI21_X1 U67 ( .B1(n800), .B2(n75), .A(n83), .ZN(n357) );
  NAND2_X1 U68 ( .A1(\mem[3][7] ), .A2(n785), .ZN(n83) );
  OAI21_X1 U69 ( .B1(n799), .B2(n785), .A(n84), .ZN(n358) );
  NAND2_X1 U70 ( .A1(\mem[3][8] ), .A2(n785), .ZN(n84) );
  OAI21_X1 U71 ( .B1(n798), .B2(n75), .A(n85), .ZN(n359) );
  NAND2_X1 U72 ( .A1(\mem[3][9] ), .A2(n785), .ZN(n85) );
  OAI21_X1 U73 ( .B1(n797), .B2(n75), .A(n86), .ZN(n360) );
  NAND2_X1 U74 ( .A1(\mem[3][10] ), .A2(n785), .ZN(n86) );
  OAI21_X1 U75 ( .B1(n796), .B2(n75), .A(n87), .ZN(n361) );
  NAND2_X1 U76 ( .A1(\mem[3][11] ), .A2(n785), .ZN(n87) );
  OAI21_X1 U77 ( .B1(n795), .B2(n75), .A(n88), .ZN(n362) );
  NAND2_X1 U78 ( .A1(\mem[3][12] ), .A2(n785), .ZN(n88) );
  OAI21_X1 U79 ( .B1(n794), .B2(n75), .A(n89), .ZN(n363) );
  NAND2_X1 U80 ( .A1(\mem[3][13] ), .A2(n785), .ZN(n89) );
  OAI21_X1 U81 ( .B1(n793), .B2(n75), .A(n90), .ZN(n364) );
  NAND2_X1 U82 ( .A1(\mem[3][14] ), .A2(n785), .ZN(n90) );
  OAI21_X1 U83 ( .B1(n800), .B2(n39), .A(n47), .ZN(n325) );
  NAND2_X1 U84 ( .A1(\mem[1][7] ), .A2(n787), .ZN(n47) );
  OAI21_X1 U85 ( .B1(n799), .B2(n787), .A(n48), .ZN(n326) );
  NAND2_X1 U86 ( .A1(\mem[1][8] ), .A2(n787), .ZN(n48) );
  OAI21_X1 U87 ( .B1(n798), .B2(n39), .A(n49), .ZN(n327) );
  NAND2_X1 U88 ( .A1(\mem[1][9] ), .A2(n787), .ZN(n49) );
  OAI21_X1 U89 ( .B1(n797), .B2(n39), .A(n50), .ZN(n328) );
  NAND2_X1 U90 ( .A1(\mem[1][10] ), .A2(n787), .ZN(n50) );
  OAI21_X1 U91 ( .B1(n796), .B2(n39), .A(n51), .ZN(n329) );
  NAND2_X1 U92 ( .A1(\mem[1][11] ), .A2(n787), .ZN(n51) );
  OAI21_X1 U93 ( .B1(n795), .B2(n39), .A(n52), .ZN(n330) );
  NAND2_X1 U94 ( .A1(\mem[1][12] ), .A2(n787), .ZN(n52) );
  OAI21_X1 U95 ( .B1(n794), .B2(n39), .A(n53), .ZN(n331) );
  NAND2_X1 U96 ( .A1(\mem[1][13] ), .A2(n787), .ZN(n53) );
  OAI21_X1 U97 ( .B1(n793), .B2(n39), .A(n54), .ZN(n332) );
  NAND2_X1 U98 ( .A1(\mem[1][14] ), .A2(n787), .ZN(n54) );
  OAI21_X1 U99 ( .B1(n800), .B2(n92), .A(n100), .ZN(n373) );
  NAND2_X1 U100 ( .A1(\mem[4][7] ), .A2(n784), .ZN(n100) );
  OAI21_X1 U101 ( .B1(n799), .B2(n92), .A(n101), .ZN(n374) );
  NAND2_X1 U102 ( .A1(\mem[4][8] ), .A2(n784), .ZN(n101) );
  OAI21_X1 U103 ( .B1(n798), .B2(n92), .A(n102), .ZN(n375) );
  NAND2_X1 U104 ( .A1(\mem[4][9] ), .A2(n92), .ZN(n102) );
  OAI21_X1 U105 ( .B1(n797), .B2(n92), .A(n103), .ZN(n376) );
  NAND2_X1 U106 ( .A1(\mem[4][10] ), .A2(n92), .ZN(n103) );
  OAI21_X1 U107 ( .B1(n796), .B2(n92), .A(n104), .ZN(n377) );
  NAND2_X1 U108 ( .A1(\mem[4][11] ), .A2(n92), .ZN(n104) );
  OAI21_X1 U109 ( .B1(n795), .B2(n92), .A(n105), .ZN(n378) );
  NAND2_X1 U110 ( .A1(\mem[4][12] ), .A2(n784), .ZN(n105) );
  OAI21_X1 U111 ( .B1(n794), .B2(n92), .A(n106), .ZN(n379) );
  NAND2_X1 U112 ( .A1(\mem[4][13] ), .A2(n92), .ZN(n106) );
  OAI21_X1 U113 ( .B1(n793), .B2(n92), .A(n107), .ZN(n380) );
  NAND2_X1 U114 ( .A1(\mem[4][14] ), .A2(n92), .ZN(n107) );
  OAI21_X1 U115 ( .B1(n800), .B2(n110), .A(n118), .ZN(n389) );
  NAND2_X1 U116 ( .A1(\mem[5][7] ), .A2(n783), .ZN(n118) );
  OAI21_X1 U117 ( .B1(n799), .B2(n110), .A(n119), .ZN(n390) );
  NAND2_X1 U118 ( .A1(\mem[5][8] ), .A2(n783), .ZN(n119) );
  OAI21_X1 U119 ( .B1(n798), .B2(n110), .A(n120), .ZN(n391) );
  NAND2_X1 U120 ( .A1(\mem[5][9] ), .A2(n110), .ZN(n120) );
  OAI21_X1 U121 ( .B1(n797), .B2(n110), .A(n121), .ZN(n392) );
  NAND2_X1 U122 ( .A1(\mem[5][10] ), .A2(n110), .ZN(n121) );
  OAI21_X1 U123 ( .B1(n796), .B2(n110), .A(n122), .ZN(n393) );
  NAND2_X1 U124 ( .A1(\mem[5][11] ), .A2(n110), .ZN(n122) );
  OAI21_X1 U125 ( .B1(n795), .B2(n110), .A(n123), .ZN(n394) );
  NAND2_X1 U126 ( .A1(\mem[5][12] ), .A2(n783), .ZN(n123) );
  OAI21_X1 U127 ( .B1(n794), .B2(n110), .A(n124), .ZN(n395) );
  NAND2_X1 U128 ( .A1(\mem[5][13] ), .A2(n110), .ZN(n124) );
  OAI21_X1 U129 ( .B1(n793), .B2(n110), .A(n125), .ZN(n396) );
  NAND2_X1 U130 ( .A1(\mem[5][14] ), .A2(n110), .ZN(n125) );
  OAI21_X1 U131 ( .B1(n800), .B2(n127), .A(n135), .ZN(n405) );
  NAND2_X1 U132 ( .A1(\mem[6][7] ), .A2(n782), .ZN(n135) );
  OAI21_X1 U133 ( .B1(n799), .B2(n782), .A(n136), .ZN(n406) );
  NAND2_X1 U134 ( .A1(\mem[6][8] ), .A2(n782), .ZN(n136) );
  OAI21_X1 U135 ( .B1(n798), .B2(n127), .A(n137), .ZN(n407) );
  NAND2_X1 U136 ( .A1(\mem[6][9] ), .A2(n782), .ZN(n137) );
  OAI21_X1 U137 ( .B1(n797), .B2(n127), .A(n138), .ZN(n408) );
  NAND2_X1 U138 ( .A1(\mem[6][10] ), .A2(n782), .ZN(n138) );
  OAI21_X1 U139 ( .B1(n796), .B2(n127), .A(n139), .ZN(n409) );
  NAND2_X1 U140 ( .A1(\mem[6][11] ), .A2(n782), .ZN(n139) );
  OAI21_X1 U141 ( .B1(n795), .B2(n127), .A(n140), .ZN(n410) );
  NAND2_X1 U142 ( .A1(\mem[6][12] ), .A2(n782), .ZN(n140) );
  OAI21_X1 U143 ( .B1(n794), .B2(n127), .A(n141), .ZN(n411) );
  NAND2_X1 U144 ( .A1(\mem[6][13] ), .A2(n782), .ZN(n141) );
  OAI21_X1 U145 ( .B1(n793), .B2(n127), .A(n142), .ZN(n412) );
  NAND2_X1 U146 ( .A1(\mem[6][14] ), .A2(n782), .ZN(n142) );
  OAI21_X1 U147 ( .B1(n800), .B2(n146), .A(n154), .ZN(n421) );
  NAND2_X1 U148 ( .A1(\mem[7][7] ), .A2(n781), .ZN(n154) );
  OAI21_X1 U149 ( .B1(n799), .B2(n781), .A(n155), .ZN(n422) );
  NAND2_X1 U150 ( .A1(\mem[7][8] ), .A2(n781), .ZN(n155) );
  OAI21_X1 U151 ( .B1(n798), .B2(n146), .A(n156), .ZN(n423) );
  NAND2_X1 U152 ( .A1(\mem[7][9] ), .A2(n781), .ZN(n156) );
  OAI21_X1 U153 ( .B1(n797), .B2(n146), .A(n157), .ZN(n424) );
  NAND2_X1 U154 ( .A1(\mem[7][10] ), .A2(n781), .ZN(n157) );
  OAI21_X1 U155 ( .B1(n796), .B2(n146), .A(n158), .ZN(n425) );
  NAND2_X1 U156 ( .A1(\mem[7][11] ), .A2(n781), .ZN(n158) );
  OAI21_X1 U157 ( .B1(n795), .B2(n146), .A(n159), .ZN(n426) );
  NAND2_X1 U158 ( .A1(\mem[7][12] ), .A2(n781), .ZN(n159) );
  OAI21_X1 U159 ( .B1(n794), .B2(n146), .A(n160), .ZN(n427) );
  NAND2_X1 U160 ( .A1(\mem[7][13] ), .A2(n781), .ZN(n160) );
  OAI21_X1 U161 ( .B1(n793), .B2(n146), .A(n161), .ZN(n428) );
  NAND2_X1 U162 ( .A1(\mem[7][14] ), .A2(n781), .ZN(n161) );
  OAI21_X1 U163 ( .B1(n800), .B2(n780), .A(n171), .ZN(n437) );
  NAND2_X1 U164 ( .A1(\mem[8][7] ), .A2(n780), .ZN(n171) );
  OAI21_X1 U165 ( .B1(n799), .B2(n780), .A(n172), .ZN(n438) );
  NAND2_X1 U166 ( .A1(\mem[8][8] ), .A2(n163), .ZN(n172) );
  OAI21_X1 U167 ( .B1(n798), .B2(n780), .A(n173), .ZN(n439) );
  NAND2_X1 U168 ( .A1(\mem[8][9] ), .A2(n163), .ZN(n173) );
  OAI21_X1 U169 ( .B1(n797), .B2(n780), .A(n174), .ZN(n440) );
  NAND2_X1 U170 ( .A1(\mem[8][10] ), .A2(n163), .ZN(n174) );
  OAI21_X1 U171 ( .B1(n796), .B2(n780), .A(n175), .ZN(n441) );
  NAND2_X1 U172 ( .A1(\mem[8][11] ), .A2(n163), .ZN(n175) );
  OAI21_X1 U173 ( .B1(n795), .B2(n780), .A(n176), .ZN(n442) );
  NAND2_X1 U174 ( .A1(\mem[8][12] ), .A2(n163), .ZN(n176) );
  OAI21_X1 U175 ( .B1(n794), .B2(n780), .A(n177), .ZN(n443) );
  NAND2_X1 U176 ( .A1(\mem[8][13] ), .A2(n163), .ZN(n177) );
  OAI21_X1 U177 ( .B1(n793), .B2(n780), .A(n178), .ZN(n444) );
  NAND2_X1 U178 ( .A1(\mem[8][14] ), .A2(n163), .ZN(n178) );
  OAI21_X1 U179 ( .B1(n800), .B2(n181), .A(n189), .ZN(n453) );
  NAND2_X1 U180 ( .A1(\mem[9][7] ), .A2(n779), .ZN(n189) );
  OAI21_X1 U181 ( .B1(n799), .B2(n779), .A(n190), .ZN(n454) );
  NAND2_X1 U182 ( .A1(\mem[9][8] ), .A2(n779), .ZN(n190) );
  OAI21_X1 U183 ( .B1(n798), .B2(n181), .A(n191), .ZN(n455) );
  NAND2_X1 U184 ( .A1(\mem[9][9] ), .A2(n779), .ZN(n191) );
  OAI21_X1 U185 ( .B1(n797), .B2(n181), .A(n192), .ZN(n456) );
  NAND2_X1 U186 ( .A1(\mem[9][10] ), .A2(n779), .ZN(n192) );
  OAI21_X1 U187 ( .B1(n796), .B2(n181), .A(n193), .ZN(n457) );
  NAND2_X1 U188 ( .A1(\mem[9][11] ), .A2(n779), .ZN(n193) );
  OAI21_X1 U189 ( .B1(n795), .B2(n181), .A(n194), .ZN(n458) );
  NAND2_X1 U190 ( .A1(\mem[9][12] ), .A2(n779), .ZN(n194) );
  OAI21_X1 U191 ( .B1(n794), .B2(n181), .A(n195), .ZN(n459) );
  NAND2_X1 U192 ( .A1(\mem[9][13] ), .A2(n779), .ZN(n195) );
  OAI21_X1 U193 ( .B1(n793), .B2(n181), .A(n196), .ZN(n460) );
  NAND2_X1 U194 ( .A1(\mem[9][14] ), .A2(n779), .ZN(n196) );
  OAI21_X1 U195 ( .B1(n800), .B2(n199), .A(n207), .ZN(n469) );
  NAND2_X1 U196 ( .A1(\mem[10][7] ), .A2(n778), .ZN(n207) );
  OAI21_X1 U197 ( .B1(n799), .B2(n778), .A(n208), .ZN(n470) );
  NAND2_X1 U198 ( .A1(\mem[10][8] ), .A2(n778), .ZN(n208) );
  OAI21_X1 U199 ( .B1(n798), .B2(n199), .A(n209), .ZN(n471) );
  NAND2_X1 U200 ( .A1(\mem[10][9] ), .A2(n778), .ZN(n209) );
  OAI21_X1 U201 ( .B1(n797), .B2(n199), .A(n210), .ZN(n472) );
  NAND2_X1 U202 ( .A1(\mem[10][10] ), .A2(n778), .ZN(n210) );
  OAI21_X1 U203 ( .B1(n796), .B2(n199), .A(n211), .ZN(n473) );
  NAND2_X1 U204 ( .A1(\mem[10][11] ), .A2(n778), .ZN(n211) );
  OAI21_X1 U205 ( .B1(n795), .B2(n199), .A(n212), .ZN(n474) );
  NAND2_X1 U206 ( .A1(\mem[10][12] ), .A2(n778), .ZN(n212) );
  OAI21_X1 U207 ( .B1(n794), .B2(n199), .A(n213), .ZN(n475) );
  NAND2_X1 U208 ( .A1(\mem[10][13] ), .A2(n778), .ZN(n213) );
  OAI21_X1 U209 ( .B1(n793), .B2(n199), .A(n214), .ZN(n476) );
  NAND2_X1 U210 ( .A1(\mem[10][14] ), .A2(n778), .ZN(n214) );
  OAI21_X1 U211 ( .B1(n800), .B2(n777), .A(n224), .ZN(n485) );
  NAND2_X1 U212 ( .A1(\mem[11][7] ), .A2(n777), .ZN(n224) );
  OAI21_X1 U213 ( .B1(n799), .B2(n777), .A(n225), .ZN(n486) );
  NAND2_X1 U214 ( .A1(\mem[11][8] ), .A2(n216), .ZN(n225) );
  OAI21_X1 U215 ( .B1(n798), .B2(n777), .A(n226), .ZN(n487) );
  NAND2_X1 U216 ( .A1(\mem[11][9] ), .A2(n216), .ZN(n226) );
  OAI21_X1 U217 ( .B1(n797), .B2(n777), .A(n227), .ZN(n488) );
  NAND2_X1 U218 ( .A1(\mem[11][10] ), .A2(n216), .ZN(n227) );
  OAI21_X1 U219 ( .B1(n796), .B2(n777), .A(n228), .ZN(n489) );
  NAND2_X1 U220 ( .A1(\mem[11][11] ), .A2(n216), .ZN(n228) );
  OAI21_X1 U221 ( .B1(n795), .B2(n777), .A(n229), .ZN(n490) );
  NAND2_X1 U222 ( .A1(\mem[11][12] ), .A2(n216), .ZN(n229) );
  OAI21_X1 U223 ( .B1(n794), .B2(n777), .A(n230), .ZN(n491) );
  NAND2_X1 U224 ( .A1(\mem[11][13] ), .A2(n216), .ZN(n230) );
  OAI21_X1 U225 ( .B1(n793), .B2(n777), .A(n231), .ZN(n492) );
  NAND2_X1 U226 ( .A1(\mem[11][14] ), .A2(n216), .ZN(n231) );
  OAI21_X1 U227 ( .B1(n800), .B2(n233), .A(n241), .ZN(n501) );
  NAND2_X1 U228 ( .A1(\mem[12][7] ), .A2(n776), .ZN(n241) );
  OAI21_X1 U229 ( .B1(n799), .B2(n776), .A(n242), .ZN(n502) );
  NAND2_X1 U230 ( .A1(\mem[12][8] ), .A2(n776), .ZN(n242) );
  OAI21_X1 U231 ( .B1(n798), .B2(n233), .A(n243), .ZN(n503) );
  NAND2_X1 U232 ( .A1(\mem[12][9] ), .A2(n776), .ZN(n243) );
  OAI21_X1 U233 ( .B1(n797), .B2(n233), .A(n244), .ZN(n504) );
  NAND2_X1 U234 ( .A1(\mem[12][10] ), .A2(n776), .ZN(n244) );
  OAI21_X1 U235 ( .B1(n796), .B2(n233), .A(n245), .ZN(n505) );
  NAND2_X1 U236 ( .A1(\mem[12][11] ), .A2(n776), .ZN(n245) );
  OAI21_X1 U237 ( .B1(n795), .B2(n233), .A(n246), .ZN(n506) );
  NAND2_X1 U238 ( .A1(\mem[12][12] ), .A2(n776), .ZN(n246) );
  OAI21_X1 U239 ( .B1(n794), .B2(n233), .A(n247), .ZN(n507) );
  NAND2_X1 U240 ( .A1(\mem[12][13] ), .A2(n776), .ZN(n247) );
  OAI21_X1 U241 ( .B1(n793), .B2(n233), .A(n248), .ZN(n508) );
  NAND2_X1 U242 ( .A1(\mem[12][14] ), .A2(n776), .ZN(n248) );
  OAI21_X1 U243 ( .B1(n800), .B2(n250), .A(n258), .ZN(n517) );
  NAND2_X1 U244 ( .A1(\mem[13][7] ), .A2(n775), .ZN(n258) );
  OAI21_X1 U245 ( .B1(n799), .B2(n775), .A(n259), .ZN(n518) );
  NAND2_X1 U246 ( .A1(\mem[13][8] ), .A2(n775), .ZN(n259) );
  OAI21_X1 U247 ( .B1(n798), .B2(n250), .A(n260), .ZN(n519) );
  NAND2_X1 U248 ( .A1(\mem[13][9] ), .A2(n775), .ZN(n260) );
  OAI21_X1 U249 ( .B1(n797), .B2(n250), .A(n261), .ZN(n520) );
  NAND2_X1 U250 ( .A1(\mem[13][10] ), .A2(n775), .ZN(n261) );
  OAI21_X1 U251 ( .B1(n796), .B2(n250), .A(n262), .ZN(n521) );
  NAND2_X1 U252 ( .A1(\mem[13][11] ), .A2(n775), .ZN(n262) );
  OAI21_X1 U253 ( .B1(n795), .B2(n250), .A(n263), .ZN(n522) );
  NAND2_X1 U254 ( .A1(\mem[13][12] ), .A2(n775), .ZN(n263) );
  OAI21_X1 U255 ( .B1(n794), .B2(n250), .A(n264), .ZN(n523) );
  NAND2_X1 U256 ( .A1(\mem[13][13] ), .A2(n775), .ZN(n264) );
  OAI21_X1 U257 ( .B1(n793), .B2(n250), .A(n265), .ZN(n524) );
  NAND2_X1 U258 ( .A1(\mem[13][14] ), .A2(n775), .ZN(n265) );
  OAI21_X1 U259 ( .B1(n800), .B2(n267), .A(n275), .ZN(n533) );
  NAND2_X1 U260 ( .A1(\mem[14][7] ), .A2(n774), .ZN(n275) );
  OAI21_X1 U261 ( .B1(n799), .B2(n774), .A(n276), .ZN(n534) );
  NAND2_X1 U262 ( .A1(\mem[14][8] ), .A2(n774), .ZN(n276) );
  OAI21_X1 U263 ( .B1(n798), .B2(n267), .A(n277), .ZN(n535) );
  NAND2_X1 U264 ( .A1(\mem[14][9] ), .A2(n774), .ZN(n277) );
  OAI21_X1 U265 ( .B1(n797), .B2(n267), .A(n278), .ZN(n536) );
  NAND2_X1 U266 ( .A1(\mem[14][10] ), .A2(n774), .ZN(n278) );
  OAI21_X1 U267 ( .B1(n796), .B2(n267), .A(n279), .ZN(n537) );
  NAND2_X1 U268 ( .A1(\mem[14][11] ), .A2(n774), .ZN(n279) );
  OAI21_X1 U269 ( .B1(n795), .B2(n267), .A(n280), .ZN(n538) );
  NAND2_X1 U270 ( .A1(\mem[14][12] ), .A2(n774), .ZN(n280) );
  OAI21_X1 U271 ( .B1(n794), .B2(n267), .A(n281), .ZN(n539) );
  NAND2_X1 U272 ( .A1(\mem[14][13] ), .A2(n774), .ZN(n281) );
  OAI21_X1 U273 ( .B1(n793), .B2(n267), .A(n282), .ZN(n540) );
  NAND2_X1 U274 ( .A1(\mem[14][14] ), .A2(n774), .ZN(n282) );
  OAI21_X1 U275 ( .B1(n800), .B2(n285), .A(n293), .ZN(n549) );
  NAND2_X1 U276 ( .A1(\mem[15][7] ), .A2(n773), .ZN(n293) );
  OAI21_X1 U277 ( .B1(n799), .B2(n773), .A(n294), .ZN(n550) );
  NAND2_X1 U278 ( .A1(\mem[15][8] ), .A2(n773), .ZN(n294) );
  OAI21_X1 U279 ( .B1(n798), .B2(n285), .A(n295), .ZN(n551) );
  NAND2_X1 U280 ( .A1(\mem[15][9] ), .A2(n773), .ZN(n295) );
  OAI21_X1 U281 ( .B1(n797), .B2(n285), .A(n296), .ZN(n552) );
  NAND2_X1 U282 ( .A1(\mem[15][10] ), .A2(n773), .ZN(n296) );
  OAI21_X1 U283 ( .B1(n796), .B2(n285), .A(n297), .ZN(n553) );
  NAND2_X1 U284 ( .A1(\mem[15][11] ), .A2(n773), .ZN(n297) );
  OAI21_X1 U285 ( .B1(n795), .B2(n285), .A(n298), .ZN(n554) );
  NAND2_X1 U286 ( .A1(\mem[15][12] ), .A2(n773), .ZN(n298) );
  OAI21_X1 U287 ( .B1(n794), .B2(n285), .A(n299), .ZN(n555) );
  NAND2_X1 U288 ( .A1(\mem[15][13] ), .A2(n773), .ZN(n299) );
  OAI21_X1 U289 ( .B1(n793), .B2(n285), .A(n300), .ZN(n556) );
  NAND2_X1 U290 ( .A1(\mem[15][14] ), .A2(n773), .ZN(n300) );
  OAI21_X1 U291 ( .B1(n20), .B2(n799), .A(n29), .ZN(n310) );
  NAND2_X1 U292 ( .A1(\mem[0][8] ), .A2(n788), .ZN(n29) );
  OAI21_X1 U293 ( .B1(n20), .B2(n798), .A(n30), .ZN(n311) );
  NAND2_X1 U294 ( .A1(\mem[0][9] ), .A2(n20), .ZN(n30) );
  OAI21_X1 U295 ( .B1(n788), .B2(n797), .A(n31), .ZN(n312) );
  NAND2_X1 U296 ( .A1(\mem[0][10] ), .A2(n20), .ZN(n31) );
  OAI21_X1 U297 ( .B1(n20), .B2(n796), .A(n32), .ZN(n313) );
  NAND2_X1 U298 ( .A1(\mem[0][11] ), .A2(n20), .ZN(n32) );
  OAI21_X1 U299 ( .B1(n20), .B2(n795), .A(n33), .ZN(n314) );
  NAND2_X1 U300 ( .A1(\mem[0][12] ), .A2(n20), .ZN(n33) );
  OAI21_X1 U301 ( .B1(n20), .B2(n794), .A(n34), .ZN(n315) );
  NAND2_X1 U302 ( .A1(\mem[0][13] ), .A2(n20), .ZN(n34) );
  OAI21_X1 U303 ( .B1(n20), .B2(n793), .A(n35), .ZN(n316) );
  NAND2_X1 U304 ( .A1(\mem[0][14] ), .A2(n20), .ZN(n35) );
  OAI21_X1 U305 ( .B1(n807), .B2(n39), .A(n40), .ZN(n318) );
  NAND2_X1 U306 ( .A1(\mem[1][0] ), .A2(n787), .ZN(n40) );
  OAI21_X1 U307 ( .B1(n806), .B2(n39), .A(n41), .ZN(n319) );
  NAND2_X1 U308 ( .A1(\mem[1][1] ), .A2(n787), .ZN(n41) );
  OAI21_X1 U309 ( .B1(n805), .B2(n39), .A(n42), .ZN(n320) );
  NAND2_X1 U310 ( .A1(\mem[1][2] ), .A2(n787), .ZN(n42) );
  OAI21_X1 U311 ( .B1(n804), .B2(n39), .A(n43), .ZN(n321) );
  NAND2_X1 U312 ( .A1(\mem[1][3] ), .A2(n787), .ZN(n43) );
  OAI21_X1 U313 ( .B1(n803), .B2(n39), .A(n44), .ZN(n322) );
  NAND2_X1 U314 ( .A1(\mem[1][4] ), .A2(n39), .ZN(n44) );
  OAI21_X1 U315 ( .B1(n802), .B2(n39), .A(n45), .ZN(n323) );
  NAND2_X1 U316 ( .A1(\mem[1][5] ), .A2(n39), .ZN(n45) );
  OAI21_X1 U317 ( .B1(n801), .B2(n39), .A(n46), .ZN(n324) );
  NAND2_X1 U318 ( .A1(\mem[1][6] ), .A2(n39), .ZN(n46) );
  OAI21_X1 U319 ( .B1(n792), .B2(n39), .A(n55), .ZN(n333) );
  NAND2_X1 U320 ( .A1(\mem[1][15] ), .A2(n787), .ZN(n55) );
  OAI21_X1 U321 ( .B1(n807), .B2(n57), .A(n58), .ZN(n334) );
  NAND2_X1 U322 ( .A1(\mem[2][0] ), .A2(n786), .ZN(n58) );
  OAI21_X1 U323 ( .B1(n806), .B2(n57), .A(n59), .ZN(n335) );
  NAND2_X1 U324 ( .A1(\mem[2][1] ), .A2(n786), .ZN(n59) );
  OAI21_X1 U325 ( .B1(n805), .B2(n57), .A(n60), .ZN(n336) );
  NAND2_X1 U326 ( .A1(\mem[2][2] ), .A2(n786), .ZN(n60) );
  OAI21_X1 U327 ( .B1(n804), .B2(n57), .A(n61), .ZN(n337) );
  NAND2_X1 U328 ( .A1(\mem[2][3] ), .A2(n786), .ZN(n61) );
  OAI21_X1 U329 ( .B1(n803), .B2(n57), .A(n62), .ZN(n338) );
  NAND2_X1 U330 ( .A1(\mem[2][4] ), .A2(n57), .ZN(n62) );
  OAI21_X1 U331 ( .B1(n802), .B2(n57), .A(n63), .ZN(n339) );
  NAND2_X1 U332 ( .A1(\mem[2][5] ), .A2(n57), .ZN(n63) );
  OAI21_X1 U333 ( .B1(n801), .B2(n57), .A(n64), .ZN(n340) );
  NAND2_X1 U334 ( .A1(\mem[2][6] ), .A2(n57), .ZN(n64) );
  OAI21_X1 U335 ( .B1(n792), .B2(n57), .A(n73), .ZN(n349) );
  NAND2_X1 U336 ( .A1(\mem[2][15] ), .A2(n786), .ZN(n73) );
  OAI21_X1 U337 ( .B1(n807), .B2(n75), .A(n76), .ZN(n350) );
  NAND2_X1 U338 ( .A1(\mem[3][0] ), .A2(n785), .ZN(n76) );
  OAI21_X1 U339 ( .B1(n806), .B2(n75), .A(n77), .ZN(n351) );
  NAND2_X1 U340 ( .A1(\mem[3][1] ), .A2(n785), .ZN(n77) );
  OAI21_X1 U341 ( .B1(n805), .B2(n75), .A(n78), .ZN(n352) );
  NAND2_X1 U342 ( .A1(\mem[3][2] ), .A2(n785), .ZN(n78) );
  OAI21_X1 U343 ( .B1(n804), .B2(n75), .A(n79), .ZN(n353) );
  NAND2_X1 U344 ( .A1(\mem[3][3] ), .A2(n785), .ZN(n79) );
  OAI21_X1 U345 ( .B1(n803), .B2(n75), .A(n80), .ZN(n354) );
  NAND2_X1 U346 ( .A1(\mem[3][4] ), .A2(n75), .ZN(n80) );
  OAI21_X1 U347 ( .B1(n802), .B2(n75), .A(n81), .ZN(n355) );
  NAND2_X1 U348 ( .A1(\mem[3][5] ), .A2(n75), .ZN(n81) );
  OAI21_X1 U349 ( .B1(n801), .B2(n75), .A(n82), .ZN(n356) );
  NAND2_X1 U350 ( .A1(\mem[3][6] ), .A2(n75), .ZN(n82) );
  OAI21_X1 U351 ( .B1(n792), .B2(n75), .A(n91), .ZN(n365) );
  NAND2_X1 U352 ( .A1(\mem[3][15] ), .A2(n785), .ZN(n91) );
  OAI21_X1 U353 ( .B1(n807), .B2(n784), .A(n93), .ZN(n366) );
  NAND2_X1 U354 ( .A1(\mem[4][0] ), .A2(n92), .ZN(n93) );
  OAI21_X1 U355 ( .B1(n806), .B2(n784), .A(n94), .ZN(n367) );
  NAND2_X1 U356 ( .A1(\mem[4][1] ), .A2(n92), .ZN(n94) );
  OAI21_X1 U357 ( .B1(n805), .B2(n784), .A(n95), .ZN(n368) );
  NAND2_X1 U358 ( .A1(\mem[4][2] ), .A2(n92), .ZN(n95) );
  OAI21_X1 U359 ( .B1(n804), .B2(n784), .A(n96), .ZN(n369) );
  NAND2_X1 U360 ( .A1(\mem[4][3] ), .A2(n92), .ZN(n96) );
  OAI21_X1 U361 ( .B1(n803), .B2(n784), .A(n97), .ZN(n370) );
  NAND2_X1 U362 ( .A1(\mem[4][4] ), .A2(n784), .ZN(n97) );
  OAI21_X1 U363 ( .B1(n802), .B2(n784), .A(n98), .ZN(n371) );
  NAND2_X1 U364 ( .A1(\mem[4][5] ), .A2(n784), .ZN(n98) );
  OAI21_X1 U365 ( .B1(n801), .B2(n784), .A(n99), .ZN(n372) );
  NAND2_X1 U366 ( .A1(\mem[4][6] ), .A2(n784), .ZN(n99) );
  OAI21_X1 U367 ( .B1(n792), .B2(n784), .A(n108), .ZN(n381) );
  NAND2_X1 U368 ( .A1(\mem[4][15] ), .A2(n92), .ZN(n108) );
  OAI21_X1 U369 ( .B1(n807), .B2(n783), .A(n111), .ZN(n382) );
  NAND2_X1 U370 ( .A1(\mem[5][0] ), .A2(n110), .ZN(n111) );
  OAI21_X1 U371 ( .B1(n806), .B2(n783), .A(n112), .ZN(n383) );
  NAND2_X1 U372 ( .A1(\mem[5][1] ), .A2(n110), .ZN(n112) );
  OAI21_X1 U373 ( .B1(n805), .B2(n783), .A(n113), .ZN(n384) );
  NAND2_X1 U374 ( .A1(\mem[5][2] ), .A2(n110), .ZN(n113) );
  OAI21_X1 U375 ( .B1(n804), .B2(n783), .A(n114), .ZN(n385) );
  NAND2_X1 U376 ( .A1(\mem[5][3] ), .A2(n110), .ZN(n114) );
  OAI21_X1 U377 ( .B1(n803), .B2(n783), .A(n115), .ZN(n386) );
  NAND2_X1 U378 ( .A1(\mem[5][4] ), .A2(n783), .ZN(n115) );
  OAI21_X1 U379 ( .B1(n802), .B2(n783), .A(n116), .ZN(n387) );
  NAND2_X1 U380 ( .A1(\mem[5][5] ), .A2(n783), .ZN(n116) );
  OAI21_X1 U381 ( .B1(n801), .B2(n783), .A(n117), .ZN(n388) );
  NAND2_X1 U382 ( .A1(\mem[5][6] ), .A2(n783), .ZN(n117) );
  OAI21_X1 U383 ( .B1(n792), .B2(n783), .A(n126), .ZN(n397) );
  NAND2_X1 U384 ( .A1(\mem[5][15] ), .A2(n110), .ZN(n126) );
  OAI21_X1 U385 ( .B1(n807), .B2(n127), .A(n128), .ZN(n398) );
  NAND2_X1 U386 ( .A1(\mem[6][0] ), .A2(n782), .ZN(n128) );
  OAI21_X1 U387 ( .B1(n806), .B2(n127), .A(n129), .ZN(n399) );
  NAND2_X1 U388 ( .A1(\mem[6][1] ), .A2(n782), .ZN(n129) );
  OAI21_X1 U389 ( .B1(n805), .B2(n127), .A(n130), .ZN(n400) );
  NAND2_X1 U390 ( .A1(\mem[6][2] ), .A2(n782), .ZN(n130) );
  OAI21_X1 U391 ( .B1(n804), .B2(n127), .A(n131), .ZN(n401) );
  NAND2_X1 U392 ( .A1(\mem[6][3] ), .A2(n782), .ZN(n131) );
  OAI21_X1 U393 ( .B1(n803), .B2(n127), .A(n132), .ZN(n402) );
  NAND2_X1 U394 ( .A1(\mem[6][4] ), .A2(n127), .ZN(n132) );
  OAI21_X1 U395 ( .B1(n802), .B2(n127), .A(n133), .ZN(n403) );
  NAND2_X1 U396 ( .A1(\mem[6][5] ), .A2(n127), .ZN(n133) );
  OAI21_X1 U397 ( .B1(n801), .B2(n127), .A(n134), .ZN(n404) );
  NAND2_X1 U398 ( .A1(\mem[6][6] ), .A2(n127), .ZN(n134) );
  OAI21_X1 U399 ( .B1(n792), .B2(n127), .A(n143), .ZN(n413) );
  NAND2_X1 U400 ( .A1(\mem[6][15] ), .A2(n782), .ZN(n143) );
  OAI21_X1 U401 ( .B1(n807), .B2(n146), .A(n147), .ZN(n414) );
  NAND2_X1 U402 ( .A1(\mem[7][0] ), .A2(n781), .ZN(n147) );
  OAI21_X1 U403 ( .B1(n806), .B2(n146), .A(n148), .ZN(n415) );
  NAND2_X1 U404 ( .A1(\mem[7][1] ), .A2(n781), .ZN(n148) );
  OAI21_X1 U405 ( .B1(n805), .B2(n146), .A(n149), .ZN(n416) );
  NAND2_X1 U406 ( .A1(\mem[7][2] ), .A2(n781), .ZN(n149) );
  OAI21_X1 U407 ( .B1(n804), .B2(n146), .A(n150), .ZN(n417) );
  NAND2_X1 U408 ( .A1(\mem[7][3] ), .A2(n781), .ZN(n150) );
  OAI21_X1 U409 ( .B1(n803), .B2(n146), .A(n151), .ZN(n418) );
  NAND2_X1 U410 ( .A1(\mem[7][4] ), .A2(n146), .ZN(n151) );
  OAI21_X1 U411 ( .B1(n802), .B2(n146), .A(n152), .ZN(n419) );
  NAND2_X1 U412 ( .A1(\mem[7][5] ), .A2(n146), .ZN(n152) );
  OAI21_X1 U413 ( .B1(n801), .B2(n146), .A(n153), .ZN(n420) );
  NAND2_X1 U414 ( .A1(\mem[7][6] ), .A2(n146), .ZN(n153) );
  OAI21_X1 U415 ( .B1(n792), .B2(n146), .A(n162), .ZN(n429) );
  NAND2_X1 U416 ( .A1(\mem[7][15] ), .A2(n781), .ZN(n162) );
  OAI21_X1 U417 ( .B1(n807), .B2(n780), .A(n164), .ZN(n430) );
  NAND2_X1 U418 ( .A1(\mem[8][0] ), .A2(n780), .ZN(n164) );
  OAI21_X1 U419 ( .B1(n806), .B2(n163), .A(n165), .ZN(n431) );
  NAND2_X1 U420 ( .A1(\mem[8][1] ), .A2(n163), .ZN(n165) );
  OAI21_X1 U421 ( .B1(n805), .B2(n163), .A(n166), .ZN(n432) );
  NAND2_X1 U422 ( .A1(\mem[8][2] ), .A2(n163), .ZN(n166) );
  OAI21_X1 U423 ( .B1(n804), .B2(n163), .A(n167), .ZN(n433) );
  NAND2_X1 U424 ( .A1(\mem[8][3] ), .A2(n163), .ZN(n167) );
  OAI21_X1 U425 ( .B1(n803), .B2(n163), .A(n168), .ZN(n434) );
  NAND2_X1 U426 ( .A1(\mem[8][4] ), .A2(n780), .ZN(n168) );
  OAI21_X1 U427 ( .B1(n802), .B2(n163), .A(n169), .ZN(n435) );
  NAND2_X1 U428 ( .A1(\mem[8][5] ), .A2(n780), .ZN(n169) );
  OAI21_X1 U429 ( .B1(n801), .B2(n163), .A(n170), .ZN(n436) );
  NAND2_X1 U430 ( .A1(\mem[8][6] ), .A2(n780), .ZN(n170) );
  OAI21_X1 U431 ( .B1(n792), .B2(n163), .A(n179), .ZN(n445) );
  NAND2_X1 U432 ( .A1(\mem[8][15] ), .A2(n163), .ZN(n179) );
  OAI21_X1 U433 ( .B1(n807), .B2(n181), .A(n182), .ZN(n446) );
  NAND2_X1 U434 ( .A1(\mem[9][0] ), .A2(n779), .ZN(n182) );
  OAI21_X1 U435 ( .B1(n806), .B2(n181), .A(n183), .ZN(n447) );
  NAND2_X1 U436 ( .A1(\mem[9][1] ), .A2(n779), .ZN(n183) );
  OAI21_X1 U437 ( .B1(n805), .B2(n181), .A(n184), .ZN(n448) );
  NAND2_X1 U438 ( .A1(\mem[9][2] ), .A2(n779), .ZN(n184) );
  OAI21_X1 U439 ( .B1(n804), .B2(n181), .A(n185), .ZN(n449) );
  NAND2_X1 U440 ( .A1(\mem[9][3] ), .A2(n779), .ZN(n185) );
  OAI21_X1 U441 ( .B1(n803), .B2(n181), .A(n186), .ZN(n450) );
  NAND2_X1 U442 ( .A1(\mem[9][4] ), .A2(n181), .ZN(n186) );
  OAI21_X1 U443 ( .B1(n802), .B2(n181), .A(n187), .ZN(n451) );
  NAND2_X1 U444 ( .A1(\mem[9][5] ), .A2(n181), .ZN(n187) );
  OAI21_X1 U445 ( .B1(n801), .B2(n181), .A(n188), .ZN(n452) );
  NAND2_X1 U446 ( .A1(\mem[9][6] ), .A2(n181), .ZN(n188) );
  OAI21_X1 U447 ( .B1(n792), .B2(n181), .A(n197), .ZN(n461) );
  NAND2_X1 U448 ( .A1(\mem[9][15] ), .A2(n779), .ZN(n197) );
  OAI21_X1 U449 ( .B1(n807), .B2(n199), .A(n200), .ZN(n462) );
  NAND2_X1 U450 ( .A1(\mem[10][0] ), .A2(n778), .ZN(n200) );
  OAI21_X1 U451 ( .B1(n806), .B2(n199), .A(n201), .ZN(n463) );
  NAND2_X1 U452 ( .A1(\mem[10][1] ), .A2(n778), .ZN(n201) );
  OAI21_X1 U453 ( .B1(n805), .B2(n199), .A(n202), .ZN(n464) );
  NAND2_X1 U454 ( .A1(\mem[10][2] ), .A2(n778), .ZN(n202) );
  OAI21_X1 U455 ( .B1(n804), .B2(n199), .A(n203), .ZN(n465) );
  NAND2_X1 U456 ( .A1(\mem[10][3] ), .A2(n778), .ZN(n203) );
  OAI21_X1 U457 ( .B1(n803), .B2(n199), .A(n204), .ZN(n466) );
  NAND2_X1 U458 ( .A1(\mem[10][4] ), .A2(n199), .ZN(n204) );
  OAI21_X1 U459 ( .B1(n802), .B2(n199), .A(n205), .ZN(n467) );
  NAND2_X1 U460 ( .A1(\mem[10][5] ), .A2(n199), .ZN(n205) );
  OAI21_X1 U461 ( .B1(n801), .B2(n199), .A(n206), .ZN(n468) );
  NAND2_X1 U462 ( .A1(\mem[10][6] ), .A2(n199), .ZN(n206) );
  OAI21_X1 U463 ( .B1(n792), .B2(n199), .A(n215), .ZN(n477) );
  NAND2_X1 U464 ( .A1(\mem[10][15] ), .A2(n778), .ZN(n215) );
  OAI21_X1 U465 ( .B1(n807), .B2(n777), .A(n217), .ZN(n478) );
  NAND2_X1 U466 ( .A1(\mem[11][0] ), .A2(n777), .ZN(n217) );
  OAI21_X1 U467 ( .B1(n806), .B2(n216), .A(n218), .ZN(n479) );
  NAND2_X1 U468 ( .A1(\mem[11][1] ), .A2(n216), .ZN(n218) );
  OAI21_X1 U469 ( .B1(n805), .B2(n216), .A(n219), .ZN(n480) );
  NAND2_X1 U470 ( .A1(\mem[11][2] ), .A2(n216), .ZN(n219) );
  OAI21_X1 U471 ( .B1(n804), .B2(n216), .A(n220), .ZN(n481) );
  NAND2_X1 U472 ( .A1(\mem[11][3] ), .A2(n216), .ZN(n220) );
  OAI21_X1 U473 ( .B1(n803), .B2(n216), .A(n221), .ZN(n482) );
  NAND2_X1 U474 ( .A1(\mem[11][4] ), .A2(n777), .ZN(n221) );
  OAI21_X1 U475 ( .B1(n802), .B2(n216), .A(n222), .ZN(n483) );
  NAND2_X1 U476 ( .A1(\mem[11][5] ), .A2(n777), .ZN(n222) );
  OAI21_X1 U477 ( .B1(n801), .B2(n216), .A(n223), .ZN(n484) );
  NAND2_X1 U478 ( .A1(\mem[11][6] ), .A2(n777), .ZN(n223) );
  OAI21_X1 U479 ( .B1(n792), .B2(n216), .A(n232), .ZN(n493) );
  NAND2_X1 U480 ( .A1(\mem[11][15] ), .A2(n216), .ZN(n232) );
  OAI21_X1 U481 ( .B1(n807), .B2(n233), .A(n234), .ZN(n494) );
  NAND2_X1 U482 ( .A1(\mem[12][0] ), .A2(n776), .ZN(n234) );
  OAI21_X1 U483 ( .B1(n806), .B2(n233), .A(n235), .ZN(n495) );
  NAND2_X1 U484 ( .A1(\mem[12][1] ), .A2(n776), .ZN(n235) );
  OAI21_X1 U485 ( .B1(n805), .B2(n233), .A(n236), .ZN(n496) );
  NAND2_X1 U486 ( .A1(\mem[12][2] ), .A2(n776), .ZN(n236) );
  OAI21_X1 U487 ( .B1(n804), .B2(n233), .A(n237), .ZN(n497) );
  NAND2_X1 U488 ( .A1(\mem[12][3] ), .A2(n776), .ZN(n237) );
  OAI21_X1 U489 ( .B1(n803), .B2(n233), .A(n238), .ZN(n498) );
  NAND2_X1 U490 ( .A1(\mem[12][4] ), .A2(n233), .ZN(n238) );
  OAI21_X1 U491 ( .B1(n802), .B2(n233), .A(n239), .ZN(n499) );
  NAND2_X1 U492 ( .A1(\mem[12][5] ), .A2(n233), .ZN(n239) );
  OAI21_X1 U493 ( .B1(n801), .B2(n233), .A(n240), .ZN(n500) );
  NAND2_X1 U494 ( .A1(\mem[12][6] ), .A2(n233), .ZN(n240) );
  OAI21_X1 U495 ( .B1(n792), .B2(n233), .A(n249), .ZN(n509) );
  NAND2_X1 U496 ( .A1(\mem[12][15] ), .A2(n776), .ZN(n249) );
  OAI21_X1 U497 ( .B1(n807), .B2(n250), .A(n251), .ZN(n510) );
  NAND2_X1 U498 ( .A1(\mem[13][0] ), .A2(n775), .ZN(n251) );
  OAI21_X1 U499 ( .B1(n806), .B2(n250), .A(n252), .ZN(n511) );
  NAND2_X1 U500 ( .A1(\mem[13][1] ), .A2(n775), .ZN(n252) );
  OAI21_X1 U501 ( .B1(n805), .B2(n250), .A(n253), .ZN(n512) );
  NAND2_X1 U502 ( .A1(\mem[13][2] ), .A2(n775), .ZN(n253) );
  OAI21_X1 U503 ( .B1(n804), .B2(n250), .A(n254), .ZN(n513) );
  NAND2_X1 U504 ( .A1(\mem[13][3] ), .A2(n775), .ZN(n254) );
  OAI21_X1 U505 ( .B1(n803), .B2(n250), .A(n255), .ZN(n514) );
  NAND2_X1 U506 ( .A1(\mem[13][4] ), .A2(n250), .ZN(n255) );
  OAI21_X1 U507 ( .B1(n802), .B2(n250), .A(n256), .ZN(n515) );
  NAND2_X1 U508 ( .A1(\mem[13][5] ), .A2(n250), .ZN(n256) );
  OAI21_X1 U509 ( .B1(n801), .B2(n250), .A(n257), .ZN(n516) );
  NAND2_X1 U510 ( .A1(\mem[13][6] ), .A2(n250), .ZN(n257) );
  OAI21_X1 U511 ( .B1(n792), .B2(n250), .A(n266), .ZN(n525) );
  NAND2_X1 U512 ( .A1(\mem[13][15] ), .A2(n775), .ZN(n266) );
  OAI21_X1 U513 ( .B1(n807), .B2(n267), .A(n268), .ZN(n526) );
  NAND2_X1 U514 ( .A1(\mem[14][0] ), .A2(n774), .ZN(n268) );
  OAI21_X1 U515 ( .B1(n806), .B2(n267), .A(n269), .ZN(n527) );
  NAND2_X1 U516 ( .A1(\mem[14][1] ), .A2(n774), .ZN(n269) );
  OAI21_X1 U517 ( .B1(n805), .B2(n267), .A(n270), .ZN(n528) );
  NAND2_X1 U518 ( .A1(\mem[14][2] ), .A2(n774), .ZN(n270) );
  OAI21_X1 U519 ( .B1(n804), .B2(n267), .A(n271), .ZN(n529) );
  NAND2_X1 U520 ( .A1(\mem[14][3] ), .A2(n774), .ZN(n271) );
  OAI21_X1 U521 ( .B1(n803), .B2(n267), .A(n272), .ZN(n530) );
  NAND2_X1 U522 ( .A1(\mem[14][4] ), .A2(n267), .ZN(n272) );
  OAI21_X1 U523 ( .B1(n802), .B2(n267), .A(n273), .ZN(n531) );
  NAND2_X1 U524 ( .A1(\mem[14][5] ), .A2(n267), .ZN(n273) );
  OAI21_X1 U525 ( .B1(n801), .B2(n267), .A(n274), .ZN(n532) );
  NAND2_X1 U526 ( .A1(\mem[14][6] ), .A2(n267), .ZN(n274) );
  OAI21_X1 U527 ( .B1(n792), .B2(n267), .A(n283), .ZN(n541) );
  NAND2_X1 U528 ( .A1(\mem[14][15] ), .A2(n774), .ZN(n283) );
  OAI21_X1 U529 ( .B1(n807), .B2(n285), .A(n286), .ZN(n542) );
  NAND2_X1 U530 ( .A1(\mem[15][0] ), .A2(n773), .ZN(n286) );
  OAI21_X1 U531 ( .B1(n806), .B2(n285), .A(n287), .ZN(n543) );
  NAND2_X1 U532 ( .A1(\mem[15][1] ), .A2(n773), .ZN(n287) );
  OAI21_X1 U533 ( .B1(n805), .B2(n285), .A(n288), .ZN(n544) );
  NAND2_X1 U534 ( .A1(\mem[15][2] ), .A2(n773), .ZN(n288) );
  OAI21_X1 U535 ( .B1(n804), .B2(n285), .A(n289), .ZN(n545) );
  NAND2_X1 U536 ( .A1(\mem[15][3] ), .A2(n773), .ZN(n289) );
  OAI21_X1 U537 ( .B1(n803), .B2(n285), .A(n290), .ZN(n546) );
  NAND2_X1 U538 ( .A1(\mem[15][4] ), .A2(n285), .ZN(n290) );
  OAI21_X1 U539 ( .B1(n802), .B2(n285), .A(n291), .ZN(n547) );
  NAND2_X1 U540 ( .A1(\mem[15][5] ), .A2(n285), .ZN(n291) );
  OAI21_X1 U541 ( .B1(n801), .B2(n285), .A(n292), .ZN(n548) );
  NAND2_X1 U542 ( .A1(\mem[15][6] ), .A2(n285), .ZN(n292) );
  OAI21_X1 U543 ( .B1(n792), .B2(n285), .A(n301), .ZN(n557) );
  NAND2_X1 U544 ( .A1(\mem[15][15] ), .A2(n773), .ZN(n301) );
  OAI21_X1 U545 ( .B1(n788), .B2(n807), .A(n21), .ZN(n302) );
  NAND2_X1 U546 ( .A1(\mem[0][0] ), .A2(n20), .ZN(n21) );
  OAI21_X1 U547 ( .B1(n788), .B2(n806), .A(n22), .ZN(n303) );
  NAND2_X1 U548 ( .A1(\mem[0][1] ), .A2(n20), .ZN(n22) );
  OAI21_X1 U549 ( .B1(n788), .B2(n805), .A(n23), .ZN(n304) );
  NAND2_X1 U550 ( .A1(\mem[0][2] ), .A2(n20), .ZN(n23) );
  OAI21_X1 U551 ( .B1(n788), .B2(n804), .A(n24), .ZN(n305) );
  NAND2_X1 U552 ( .A1(\mem[0][3] ), .A2(n20), .ZN(n24) );
  OAI21_X1 U553 ( .B1(n788), .B2(n803), .A(n25), .ZN(n306) );
  NAND2_X1 U554 ( .A1(\mem[0][4] ), .A2(n788), .ZN(n25) );
  OAI21_X1 U555 ( .B1(n788), .B2(n802), .A(n26), .ZN(n307) );
  NAND2_X1 U556 ( .A1(\mem[0][5] ), .A2(n788), .ZN(n26) );
  OAI21_X1 U557 ( .B1(n788), .B2(n801), .A(n27), .ZN(n308) );
  NAND2_X1 U558 ( .A1(\mem[0][6] ), .A2(n788), .ZN(n27) );
  OAI21_X1 U559 ( .B1(n788), .B2(n800), .A(n28), .ZN(n309) );
  NAND2_X1 U560 ( .A1(\mem[0][7] ), .A2(n788), .ZN(n28) );
  OAI21_X1 U561 ( .B1(n788), .B2(n792), .A(n36), .ZN(n317) );
  NAND2_X1 U562 ( .A1(\mem[0][15] ), .A2(n20), .ZN(n36) );
  AND2_X1 U563 ( .A1(N13), .A2(wr_en), .ZN(n284) );
  NOR2_X1 U564 ( .A1(n790), .A2(N12), .ZN(n74) );
  INV_X1 U565 ( .A(data_in[0]), .ZN(n807) );
  INV_X1 U566 ( .A(data_in[1]), .ZN(n806) );
  INV_X1 U567 ( .A(data_in[2]), .ZN(n805) );
  INV_X1 U568 ( .A(data_in[3]), .ZN(n804) );
  INV_X1 U569 ( .A(data_in[4]), .ZN(n803) );
  INV_X1 U570 ( .A(data_in[5]), .ZN(n802) );
  INV_X1 U571 ( .A(data_in[6]), .ZN(n801) );
  INV_X1 U572 ( .A(data_in[7]), .ZN(n800) );
  INV_X1 U573 ( .A(data_in[8]), .ZN(n799) );
  INV_X1 U574 ( .A(data_in[9]), .ZN(n798) );
  INV_X1 U575 ( .A(data_in[10]), .ZN(n797) );
  INV_X1 U576 ( .A(data_in[11]), .ZN(n796) );
  INV_X1 U577 ( .A(data_in[12]), .ZN(n795) );
  INV_X1 U578 ( .A(data_in[13]), .ZN(n794) );
  INV_X1 U579 ( .A(data_in[14]), .ZN(n793) );
  INV_X1 U580 ( .A(data_in[15]), .ZN(n792) );
  AND2_X1 U581 ( .A1(N12), .A2(n790), .ZN(n109) );
  BUF_X1 U582 ( .A(N12), .Z(n763) );
  MUX2_X1 U583 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n767), .Z(n1) );
  MUX2_X1 U584 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n767), .Z(n2) );
  MUX2_X1 U585 ( .A(n2), .B(n1), .S(n764), .Z(n3) );
  MUX2_X1 U586 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n767), .Z(n4) );
  MUX2_X1 U587 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n767), .Z(n5) );
  MUX2_X1 U588 ( .A(n5), .B(n4), .S(n766), .Z(n6) );
  MUX2_X1 U589 ( .A(n6), .B(n3), .S(n763), .Z(n7) );
  MUX2_X1 U590 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n767), .Z(n8) );
  MUX2_X1 U591 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n767), .Z(n9) );
  MUX2_X1 U592 ( .A(n9), .B(n8), .S(n765), .Z(n10) );
  MUX2_X1 U593 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n767), .Z(n11) );
  MUX2_X1 U594 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n767), .Z(n12) );
  MUX2_X1 U595 ( .A(n12), .B(n11), .S(n765), .Z(n13) );
  MUX2_X1 U596 ( .A(n13), .B(n10), .S(n763), .Z(n14) );
  MUX2_X1 U597 ( .A(n14), .B(n7), .S(N13), .Z(N29) );
  MUX2_X1 U598 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n772), .Z(n15) );
  MUX2_X1 U599 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(N10), .Z(n16) );
  MUX2_X1 U600 ( .A(n16), .B(n15), .S(n764), .Z(n17) );
  MUX2_X1 U601 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(N10), .Z(n18) );
  MUX2_X1 U602 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(N10), .Z(n19) );
  MUX2_X1 U603 ( .A(n19), .B(n18), .S(n764), .Z(n558) );
  MUX2_X1 U604 ( .A(n558), .B(n17), .S(n763), .Z(n559) );
  MUX2_X1 U605 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(N10), .Z(n560) );
  MUX2_X1 U606 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(N10), .Z(n561) );
  MUX2_X1 U607 ( .A(n561), .B(n560), .S(n764), .Z(n562) );
  MUX2_X1 U608 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(N10), .Z(n563) );
  MUX2_X1 U609 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n772), .Z(n564) );
  MUX2_X1 U610 ( .A(n564), .B(n563), .S(n764), .Z(n565) );
  MUX2_X1 U611 ( .A(n565), .B(n562), .S(n763), .Z(n566) );
  MUX2_X1 U612 ( .A(n566), .B(n559), .S(N13), .Z(N28) );
  MUX2_X1 U613 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n772), .Z(n567) );
  MUX2_X1 U614 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(N10), .Z(n568) );
  MUX2_X1 U615 ( .A(n568), .B(n567), .S(n764), .Z(n569) );
  MUX2_X1 U616 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(N10), .Z(n570) );
  MUX2_X1 U617 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n772), .Z(n571) );
  MUX2_X1 U618 ( .A(n571), .B(n570), .S(n764), .Z(n572) );
  MUX2_X1 U619 ( .A(n572), .B(n569), .S(n763), .Z(n573) );
  MUX2_X1 U620 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n767), .Z(n574) );
  MUX2_X1 U621 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(N10), .Z(n575) );
  MUX2_X1 U622 ( .A(n575), .B(n574), .S(n764), .Z(n576) );
  MUX2_X1 U623 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n772), .Z(n577) );
  MUX2_X1 U624 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(N10), .Z(n578) );
  MUX2_X1 U625 ( .A(n578), .B(n577), .S(n764), .Z(n579) );
  MUX2_X1 U626 ( .A(n579), .B(n576), .S(n763), .Z(n580) );
  MUX2_X1 U627 ( .A(n580), .B(n573), .S(N13), .Z(N27) );
  MUX2_X1 U628 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n767), .Z(n581) );
  MUX2_X1 U629 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n772), .Z(n582) );
  MUX2_X1 U630 ( .A(n582), .B(n581), .S(n764), .Z(n583) );
  MUX2_X1 U631 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n772), .Z(n584) );
  MUX2_X1 U632 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n585) );
  MUX2_X1 U633 ( .A(n585), .B(n584), .S(n764), .Z(n586) );
  MUX2_X1 U634 ( .A(n586), .B(n583), .S(n763), .Z(n587) );
  MUX2_X1 U635 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n767), .Z(n588) );
  MUX2_X1 U636 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n589) );
  MUX2_X1 U637 ( .A(n589), .B(n588), .S(n764), .Z(n590) );
  MUX2_X1 U638 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n591) );
  MUX2_X1 U639 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n592) );
  MUX2_X1 U640 ( .A(n592), .B(n591), .S(n764), .Z(n593) );
  MUX2_X1 U641 ( .A(n593), .B(n590), .S(n763), .Z(n594) );
  MUX2_X1 U642 ( .A(n594), .B(n587), .S(N13), .Z(N26) );
  MUX2_X1 U643 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n768), .Z(n595) );
  MUX2_X1 U644 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n768), .Z(n596) );
  MUX2_X1 U645 ( .A(n596), .B(n595), .S(n765), .Z(n597) );
  MUX2_X1 U646 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n768), .Z(n598) );
  MUX2_X1 U647 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n768), .Z(n599) );
  MUX2_X1 U648 ( .A(n599), .B(n598), .S(n765), .Z(n600) );
  MUX2_X1 U649 ( .A(n600), .B(n597), .S(n763), .Z(n601) );
  MUX2_X1 U650 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n768), .Z(n602) );
  MUX2_X1 U651 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n768), .Z(n603) );
  MUX2_X1 U652 ( .A(n603), .B(n602), .S(n765), .Z(n604) );
  MUX2_X1 U653 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n768), .Z(n605) );
  MUX2_X1 U654 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n768), .Z(n606) );
  MUX2_X1 U655 ( .A(n606), .B(n605), .S(n765), .Z(n607) );
  MUX2_X1 U656 ( .A(n607), .B(n604), .S(N12), .Z(n608) );
  MUX2_X1 U657 ( .A(n608), .B(n601), .S(N13), .Z(N25) );
  MUX2_X1 U658 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n768), .Z(n609) );
  MUX2_X1 U659 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n768), .Z(n610) );
  MUX2_X1 U660 ( .A(n610), .B(n609), .S(n765), .Z(n611) );
  MUX2_X1 U661 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n768), .Z(n612) );
  MUX2_X1 U662 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n768), .Z(n613) );
  MUX2_X1 U663 ( .A(n613), .B(n612), .S(n765), .Z(n614) );
  MUX2_X1 U664 ( .A(n614), .B(n611), .S(n763), .Z(n615) );
  MUX2_X1 U665 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n769), .Z(n616) );
  MUX2_X1 U666 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n769), .Z(n617) );
  MUX2_X1 U667 ( .A(n617), .B(n616), .S(n765), .Z(n618) );
  MUX2_X1 U668 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n769), .Z(n619) );
  MUX2_X1 U669 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n769), .Z(n620) );
  MUX2_X1 U670 ( .A(n620), .B(n619), .S(n765), .Z(n621) );
  MUX2_X1 U671 ( .A(n621), .B(n618), .S(N12), .Z(n622) );
  MUX2_X1 U672 ( .A(n622), .B(n615), .S(N13), .Z(N24) );
  MUX2_X1 U673 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n769), .Z(n623) );
  MUX2_X1 U674 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n769), .Z(n624) );
  MUX2_X1 U675 ( .A(n624), .B(n623), .S(n765), .Z(n625) );
  MUX2_X1 U676 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n769), .Z(n626) );
  MUX2_X1 U677 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n769), .Z(n627) );
  MUX2_X1 U678 ( .A(n627), .B(n626), .S(n765), .Z(n628) );
  MUX2_X1 U679 ( .A(n628), .B(n625), .S(n763), .Z(n629) );
  MUX2_X1 U680 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n769), .Z(n630) );
  MUX2_X1 U681 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n769), .Z(n631) );
  MUX2_X1 U682 ( .A(n631), .B(n630), .S(n765), .Z(n632) );
  MUX2_X1 U683 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n769), .Z(n633) );
  MUX2_X1 U684 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n769), .Z(n634) );
  MUX2_X1 U685 ( .A(n634), .B(n633), .S(n765), .Z(n635) );
  MUX2_X1 U686 ( .A(n635), .B(n632), .S(N12), .Z(n636) );
  MUX2_X1 U687 ( .A(n636), .B(n629), .S(N13), .Z(N23) );
  MUX2_X1 U688 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n772), .Z(n637) );
  MUX2_X1 U689 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n770), .Z(n638) );
  MUX2_X1 U690 ( .A(n638), .B(n637), .S(n766), .Z(n639) );
  MUX2_X1 U691 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n769), .Z(n640) );
  MUX2_X1 U692 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n771), .Z(n641) );
  MUX2_X1 U693 ( .A(n641), .B(n640), .S(n766), .Z(n642) );
  MUX2_X1 U694 ( .A(n642), .B(n639), .S(n763), .Z(n643) );
  MUX2_X1 U695 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n768), .Z(n644) );
  MUX2_X1 U696 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n770), .Z(n645) );
  MUX2_X1 U697 ( .A(n645), .B(n644), .S(n766), .Z(n646) );
  MUX2_X1 U698 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n769), .Z(n647) );
  MUX2_X1 U699 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n768), .Z(n648) );
  MUX2_X1 U700 ( .A(n648), .B(n647), .S(n766), .Z(n649) );
  MUX2_X1 U701 ( .A(n649), .B(n646), .S(N12), .Z(n650) );
  MUX2_X1 U702 ( .A(n650), .B(n643), .S(N13), .Z(N22) );
  MUX2_X1 U703 ( .A(\mem[14][8] ), .B(\mem[15][8] ), .S(n770), .Z(n651) );
  MUX2_X1 U704 ( .A(\mem[12][8] ), .B(\mem[13][8] ), .S(n768), .Z(n652) );
  MUX2_X1 U705 ( .A(n652), .B(n651), .S(n766), .Z(n653) );
  MUX2_X1 U706 ( .A(\mem[10][8] ), .B(\mem[11][8] ), .S(n771), .Z(n654) );
  MUX2_X1 U707 ( .A(\mem[8][8] ), .B(\mem[9][8] ), .S(n769), .Z(n655) );
  MUX2_X1 U708 ( .A(n655), .B(n654), .S(n766), .Z(n656) );
  MUX2_X1 U709 ( .A(n656), .B(n653), .S(n763), .Z(n657) );
  MUX2_X1 U710 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n772), .Z(n658) );
  MUX2_X1 U711 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n772), .Z(n659) );
  MUX2_X1 U712 ( .A(n659), .B(n658), .S(n766), .Z(n660) );
  MUX2_X1 U713 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n772), .Z(n661) );
  MUX2_X1 U714 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n772), .Z(n662) );
  MUX2_X1 U715 ( .A(n662), .B(n661), .S(n766), .Z(n663) );
  MUX2_X1 U716 ( .A(n663), .B(n660), .S(N12), .Z(n664) );
  MUX2_X1 U717 ( .A(n664), .B(n657), .S(N13), .Z(N21) );
  MUX2_X1 U718 ( .A(\mem[14][9] ), .B(\mem[15][9] ), .S(n772), .Z(n665) );
  MUX2_X1 U719 ( .A(\mem[12][9] ), .B(\mem[13][9] ), .S(n772), .Z(n666) );
  MUX2_X1 U720 ( .A(n666), .B(n665), .S(n766), .Z(n667) );
  MUX2_X1 U721 ( .A(\mem[10][9] ), .B(\mem[11][9] ), .S(n772), .Z(n668) );
  MUX2_X1 U722 ( .A(\mem[8][9] ), .B(\mem[9][9] ), .S(n772), .Z(n669) );
  MUX2_X1 U723 ( .A(n669), .B(n668), .S(n766), .Z(n670) );
  MUX2_X1 U724 ( .A(n670), .B(n667), .S(n763), .Z(n671) );
  MUX2_X1 U725 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n772), .Z(n672) );
  MUX2_X1 U726 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n772), .Z(n673) );
  MUX2_X1 U727 ( .A(n673), .B(n672), .S(n766), .Z(n674) );
  MUX2_X1 U728 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n772), .Z(n675) );
  MUX2_X1 U729 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n772), .Z(n676) );
  MUX2_X1 U730 ( .A(n676), .B(n675), .S(n766), .Z(n677) );
  MUX2_X1 U731 ( .A(n677), .B(n674), .S(N12), .Z(n678) );
  MUX2_X1 U732 ( .A(n678), .B(n671), .S(N13), .Z(N20) );
  MUX2_X1 U733 ( .A(\mem[14][10] ), .B(\mem[15][10] ), .S(n767), .Z(n679) );
  MUX2_X1 U734 ( .A(\mem[12][10] ), .B(\mem[13][10] ), .S(n767), .Z(n680) );
  MUX2_X1 U735 ( .A(n680), .B(n679), .S(n764), .Z(n681) );
  MUX2_X1 U736 ( .A(\mem[10][10] ), .B(\mem[11][10] ), .S(n767), .Z(n682) );
  MUX2_X1 U737 ( .A(\mem[8][10] ), .B(\mem[9][10] ), .S(n767), .Z(n683) );
  MUX2_X1 U738 ( .A(n683), .B(n682), .S(n766), .Z(n684) );
  MUX2_X1 U739 ( .A(n684), .B(n681), .S(n763), .Z(n685) );
  MUX2_X1 U740 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n767), .Z(n686) );
  MUX2_X1 U741 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n767), .Z(n687) );
  MUX2_X1 U742 ( .A(n687), .B(n686), .S(n766), .Z(n688) );
  MUX2_X1 U743 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n767), .Z(n689) );
  MUX2_X1 U744 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n767), .Z(n690) );
  MUX2_X1 U745 ( .A(n690), .B(n689), .S(n765), .Z(n691) );
  MUX2_X1 U746 ( .A(n691), .B(n688), .S(N12), .Z(n692) );
  MUX2_X1 U747 ( .A(n692), .B(n685), .S(N13), .Z(N19) );
  MUX2_X1 U748 ( .A(\mem[14][11] ), .B(\mem[15][11] ), .S(n767), .Z(n693) );
  MUX2_X1 U749 ( .A(\mem[12][11] ), .B(\mem[13][11] ), .S(n767), .Z(n694) );
  MUX2_X1 U750 ( .A(n694), .B(n693), .S(n765), .Z(n695) );
  MUX2_X1 U751 ( .A(\mem[10][11] ), .B(\mem[11][11] ), .S(n767), .Z(n696) );
  MUX2_X1 U752 ( .A(\mem[8][11] ), .B(\mem[9][11] ), .S(n767), .Z(n697) );
  MUX2_X1 U753 ( .A(n697), .B(n696), .S(n764), .Z(n698) );
  MUX2_X1 U754 ( .A(n698), .B(n695), .S(n763), .Z(n699) );
  MUX2_X1 U755 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n770), .Z(n700) );
  MUX2_X1 U756 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n770), .Z(n701) );
  MUX2_X1 U757 ( .A(n701), .B(n700), .S(n764), .Z(n702) );
  MUX2_X1 U758 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n770), .Z(n703) );
  MUX2_X1 U759 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n770), .Z(n704) );
  MUX2_X1 U760 ( .A(n704), .B(n703), .S(n764), .Z(n705) );
  MUX2_X1 U761 ( .A(n705), .B(n702), .S(n763), .Z(n706) );
  MUX2_X1 U762 ( .A(n706), .B(n699), .S(N13), .Z(N18) );
  MUX2_X1 U763 ( .A(\mem[14][12] ), .B(\mem[15][12] ), .S(n770), .Z(n707) );
  MUX2_X1 U764 ( .A(\mem[12][12] ), .B(\mem[13][12] ), .S(n770), .Z(n708) );
  MUX2_X1 U765 ( .A(n708), .B(n707), .S(n766), .Z(n709) );
  MUX2_X1 U766 ( .A(\mem[10][12] ), .B(\mem[11][12] ), .S(n770), .Z(n710) );
  MUX2_X1 U767 ( .A(\mem[8][12] ), .B(\mem[9][12] ), .S(n770), .Z(n711) );
  MUX2_X1 U768 ( .A(n711), .B(n710), .S(n765), .Z(n712) );
  MUX2_X1 U769 ( .A(n712), .B(n709), .S(n763), .Z(n713) );
  MUX2_X1 U770 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n770), .Z(n714) );
  MUX2_X1 U771 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n770), .Z(n715) );
  MUX2_X1 U772 ( .A(n715), .B(n714), .S(n764), .Z(n716) );
  MUX2_X1 U773 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n770), .Z(n717) );
  MUX2_X1 U774 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n770), .Z(n718) );
  MUX2_X1 U775 ( .A(n718), .B(n717), .S(n766), .Z(n719) );
  MUX2_X1 U776 ( .A(n719), .B(n716), .S(N12), .Z(n720) );
  MUX2_X1 U777 ( .A(n720), .B(n713), .S(N13), .Z(N17) );
  MUX2_X1 U778 ( .A(\mem[14][13] ), .B(\mem[15][13] ), .S(n771), .Z(n721) );
  MUX2_X1 U779 ( .A(\mem[12][13] ), .B(\mem[13][13] ), .S(n771), .Z(n722) );
  MUX2_X1 U780 ( .A(n722), .B(n721), .S(n764), .Z(n723) );
  MUX2_X1 U781 ( .A(\mem[10][13] ), .B(\mem[11][13] ), .S(n771), .Z(n724) );
  MUX2_X1 U782 ( .A(\mem[8][13] ), .B(\mem[9][13] ), .S(n771), .Z(n725) );
  MUX2_X1 U783 ( .A(n725), .B(n724), .S(n765), .Z(n726) );
  MUX2_X1 U784 ( .A(n726), .B(n723), .S(n763), .Z(n727) );
  MUX2_X1 U785 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n771), .Z(n728) );
  MUX2_X1 U786 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n771), .Z(n729) );
  MUX2_X1 U787 ( .A(n729), .B(n728), .S(n765), .Z(n730) );
  MUX2_X1 U788 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n771), .Z(n731) );
  MUX2_X1 U789 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n771), .Z(n732) );
  MUX2_X1 U790 ( .A(n732), .B(n731), .S(n764), .Z(n733) );
  MUX2_X1 U791 ( .A(n733), .B(n730), .S(n763), .Z(n734) );
  MUX2_X1 U792 ( .A(n734), .B(n727), .S(N13), .Z(N16) );
  MUX2_X1 U793 ( .A(\mem[14][14] ), .B(\mem[15][14] ), .S(n771), .Z(n735) );
  MUX2_X1 U794 ( .A(\mem[12][14] ), .B(\mem[13][14] ), .S(n771), .Z(n736) );
  MUX2_X1 U795 ( .A(n736), .B(n735), .S(n765), .Z(n737) );
  MUX2_X1 U796 ( .A(\mem[10][14] ), .B(\mem[11][14] ), .S(n771), .Z(n738) );
  MUX2_X1 U797 ( .A(\mem[8][14] ), .B(\mem[9][14] ), .S(n771), .Z(n739) );
  MUX2_X1 U798 ( .A(n739), .B(n738), .S(n766), .Z(n740) );
  MUX2_X1 U799 ( .A(n740), .B(n737), .S(n763), .Z(n741) );
  MUX2_X1 U800 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n769), .Z(n742) );
  MUX2_X1 U801 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n768), .Z(n743) );
  MUX2_X1 U802 ( .A(n743), .B(n742), .S(n766), .Z(n744) );
  MUX2_X1 U803 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n771), .Z(n745) );
  MUX2_X1 U804 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n768), .Z(n746) );
  MUX2_X1 U805 ( .A(n746), .B(n745), .S(n764), .Z(n747) );
  MUX2_X1 U806 ( .A(n747), .B(n744), .S(N12), .Z(n748) );
  MUX2_X1 U807 ( .A(n748), .B(n741), .S(N13), .Z(N15) );
  MUX2_X1 U808 ( .A(\mem[14][15] ), .B(\mem[15][15] ), .S(n770), .Z(n749) );
  MUX2_X1 U809 ( .A(\mem[12][15] ), .B(\mem[13][15] ), .S(n768), .Z(n750) );
  MUX2_X1 U810 ( .A(n750), .B(n749), .S(n766), .Z(n751) );
  MUX2_X1 U811 ( .A(\mem[10][15] ), .B(\mem[11][15] ), .S(n769), .Z(n752) );
  MUX2_X1 U812 ( .A(\mem[8][15] ), .B(\mem[9][15] ), .S(n771), .Z(n753) );
  MUX2_X1 U813 ( .A(n753), .B(n752), .S(n766), .Z(n754) );
  MUX2_X1 U814 ( .A(n754), .B(n751), .S(n763), .Z(n755) );
  MUX2_X1 U815 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n771), .Z(n756) );
  MUX2_X1 U816 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n770), .Z(n757) );
  MUX2_X1 U817 ( .A(n757), .B(n756), .S(n764), .Z(n758) );
  MUX2_X1 U818 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n769), .Z(n759) );
  MUX2_X1 U819 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n770), .Z(n760) );
  MUX2_X1 U820 ( .A(n760), .B(n759), .S(n765), .Z(n761) );
  MUX2_X1 U821 ( .A(n761), .B(n758), .S(n763), .Z(n762) );
  MUX2_X1 U822 ( .A(n762), .B(n755), .S(N13), .Z(N14) );
  CLKBUF_X1 U823 ( .A(N10), .Z(n767) );
  INV_X1 U824 ( .A(N10), .ZN(n789) );
  INV_X1 U825 ( .A(N11), .ZN(n790) );
endmodule


module datapath_DW_mult_tc_15 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346;

  FA_X1 U11 ( .A(n50), .B(n53), .CI(n11), .CO(n10), .S(product[5]) );
  FA_X1 U12 ( .A(n54), .B(n55), .CI(n12), .CO(n11), .S(product[4]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n289), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n288), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n292), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n291), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n294), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  INV_X2 U157 ( .A(n295), .ZN(n216) );
  BUF_X2 U158 ( .A(a[3]), .Z(n213) );
  INV_X1 U159 ( .A(n15), .ZN(n285) );
  XNOR2_X1 U160 ( .A(n260), .B(n220), .ZN(product[11]) );
  CLKBUF_X1 U161 ( .A(b[1]), .Z(n206) );
  XNOR2_X1 U162 ( .A(n286), .B(n15), .ZN(n207) );
  AND3_X1 U163 ( .A1(n221), .A2(n222), .A3(n223), .ZN(product[15]) );
  XNOR2_X1 U164 ( .A(n17), .B(n285), .ZN(n209) );
  NAND3_X1 U165 ( .A1(n263), .A2(n262), .A3(n261), .ZN(n210) );
  AND2_X1 U166 ( .A1(n104), .A2(n72), .ZN(n211) );
  INV_X1 U167 ( .A(a[0]), .ZN(n212) );
  INV_X1 U168 ( .A(a[0]), .ZN(n296) );
  XOR2_X1 U169 ( .A(a[5]), .B(a[4]), .Z(n341) );
  XNOR2_X1 U170 ( .A(b[1]), .B(a[1]), .ZN(n214) );
  NAND2_X1 U171 ( .A1(n282), .A2(n340), .ZN(n215) );
  NAND2_X1 U172 ( .A1(n282), .A2(n340), .ZN(n304) );
  NAND3_X1 U173 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n217) );
  XNOR2_X1 U174 ( .A(n256), .B(n218), .ZN(product[10]) );
  AND3_X1 U175 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n218) );
  XNOR2_X1 U176 ( .A(n3), .B(n209), .ZN(product[13]) );
  XNOR2_X1 U177 ( .A(n2), .B(n207), .ZN(product[14]) );
  NAND3_X1 U178 ( .A1(n274), .A2(n275), .A3(n276), .ZN(n219) );
  NAND2_X1 U179 ( .A1(a[1]), .A2(n296), .ZN(n298) );
  AND3_X1 U180 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n220) );
  NAND2_X1 U181 ( .A1(n217), .A2(n286), .ZN(n221) );
  NAND2_X1 U182 ( .A1(n217), .A2(n15), .ZN(n222) );
  NAND2_X1 U183 ( .A1(n286), .A2(n15), .ZN(n223) );
  XNOR2_X1 U184 ( .A(a[2]), .B(a[1]), .ZN(n224) );
  NAND3_X1 U185 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n225) );
  NAND3_X1 U186 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n226) );
  CLKBUF_X1 U187 ( .A(b[0]), .Z(n227) );
  CLKBUF_X1 U188 ( .A(n302), .Z(n283) );
  XNOR2_X1 U189 ( .A(n211), .B(n228), .ZN(product[2]) );
  XNOR2_X1 U190 ( .A(n96), .B(n103), .ZN(n228) );
  NAND3_X1 U191 ( .A1(n274), .A2(n275), .A3(n276), .ZN(n229) );
  XNOR2_X1 U192 ( .A(n247), .B(n230), .ZN(product[3]) );
  XNOR2_X1 U193 ( .A(n56), .B(n71), .ZN(n230) );
  XOR2_X1 U194 ( .A(n46), .B(n49), .Z(n231) );
  XOR2_X1 U195 ( .A(n10), .B(n231), .Z(product[6]) );
  NAND2_X1 U196 ( .A1(n10), .A2(n46), .ZN(n232) );
  NAND2_X1 U197 ( .A1(n10), .A2(n49), .ZN(n233) );
  NAND2_X1 U198 ( .A1(n46), .A2(n49), .ZN(n234) );
  NAND3_X1 U199 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n9) );
  NAND3_X1 U200 ( .A1(n263), .A2(n262), .A3(n261), .ZN(n235) );
  NAND3_X1 U201 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n236) );
  NAND3_X1 U202 ( .A1(n245), .A2(n244), .A3(n246), .ZN(n237) );
  CLKBUF_X1 U203 ( .A(n227), .Z(n238) );
  XOR2_X1 U204 ( .A(n18), .B(n19), .Z(n239) );
  XOR2_X1 U205 ( .A(n236), .B(n239), .Z(product[12]) );
  NAND2_X1 U206 ( .A1(n210), .A2(n18), .ZN(n240) );
  NAND2_X1 U207 ( .A1(n235), .A2(n19), .ZN(n241) );
  NAND2_X1 U208 ( .A1(n18), .A2(n19), .ZN(n242) );
  NAND3_X1 U209 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n3) );
  XOR2_X1 U210 ( .A(n33), .B(n28), .Z(n243) );
  XOR2_X1 U211 ( .A(n219), .B(n243), .Z(product[9]) );
  NAND2_X1 U212 ( .A1(n229), .A2(n33), .ZN(n244) );
  NAND2_X1 U213 ( .A1(n7), .A2(n28), .ZN(n245) );
  NAND2_X1 U214 ( .A1(n33), .A2(n28), .ZN(n246) );
  NAND3_X1 U215 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n6) );
  NAND3_X1 U216 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n247) );
  NAND2_X1 U217 ( .A1(n3), .A2(n17), .ZN(n248) );
  NAND2_X1 U218 ( .A1(n225), .A2(n285), .ZN(n249) );
  NAND2_X1 U219 ( .A1(n17), .A2(n285), .ZN(n250) );
  NAND3_X1 U220 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n2) );
  NAND3_X1 U221 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n251) );
  NAND2_X1 U222 ( .A1(a[4]), .A2(a[3]), .ZN(n254) );
  NAND2_X1 U223 ( .A1(n252), .A2(n253), .ZN(n255) );
  NAND2_X2 U224 ( .A1(n254), .A2(n255), .ZN(n312) );
  INV_X1 U225 ( .A(a[4]), .ZN(n252) );
  INV_X1 U226 ( .A(a[3]), .ZN(n253) );
  XOR2_X1 U227 ( .A(n24), .B(n27), .Z(n256) );
  NAND2_X1 U228 ( .A1(n24), .A2(n27), .ZN(n257) );
  NAND2_X1 U229 ( .A1(n24), .A2(n6), .ZN(n258) );
  NAND2_X1 U230 ( .A1(n27), .A2(n237), .ZN(n259) );
  NAND3_X1 U231 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n5) );
  XOR2_X1 U232 ( .A(n20), .B(n23), .Z(n260) );
  NAND2_X1 U233 ( .A1(n20), .A2(n23), .ZN(n261) );
  NAND2_X1 U234 ( .A1(n20), .A2(n251), .ZN(n262) );
  NAND2_X1 U235 ( .A1(n23), .A2(n5), .ZN(n263) );
  NAND2_X1 U236 ( .A1(n211), .A2(n96), .ZN(n264) );
  NAND2_X1 U237 ( .A1(n14), .A2(n103), .ZN(n265) );
  NAND2_X1 U238 ( .A1(n96), .A2(n103), .ZN(n266) );
  NAND3_X1 U239 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n13) );
  NAND3_X1 U240 ( .A1(n271), .A2(n270), .A3(n272), .ZN(n267) );
  NAND3_X1 U241 ( .A1(n270), .A2(n271), .A3(n272), .ZN(n268) );
  XOR2_X1 U242 ( .A(n40), .B(n45), .Z(n269) );
  XOR2_X1 U243 ( .A(n269), .B(n9), .Z(product[7]) );
  NAND2_X1 U244 ( .A1(n40), .A2(n45), .ZN(n270) );
  NAND2_X1 U245 ( .A1(n40), .A2(n226), .ZN(n271) );
  NAND2_X1 U246 ( .A1(n45), .A2(n226), .ZN(n272) );
  NAND3_X1 U247 ( .A1(n272), .A2(n271), .A3(n270), .ZN(n8) );
  XOR2_X1 U248 ( .A(n34), .B(n39), .Z(n273) );
  XOR2_X1 U249 ( .A(n273), .B(n268), .Z(product[8]) );
  NAND2_X1 U250 ( .A1(n34), .A2(n39), .ZN(n274) );
  NAND2_X1 U251 ( .A1(n34), .A2(n267), .ZN(n275) );
  NAND2_X1 U252 ( .A1(n39), .A2(n8), .ZN(n276) );
  NAND3_X1 U253 ( .A1(n276), .A2(n275), .A3(n274), .ZN(n7) );
  XOR2_X1 U254 ( .A(n213), .B(n284), .Z(n303) );
  XOR2_X1 U255 ( .A(n278), .B(n102), .Z(n277) );
  OAI22_X1 U256 ( .A1(n303), .A2(n304), .B1(n224), .B2(n305), .ZN(n278) );
  NAND2_X1 U257 ( .A1(n247), .A2(n277), .ZN(n279) );
  NAND2_X1 U258 ( .A1(n13), .A2(n71), .ZN(n280) );
  NAND2_X1 U259 ( .A1(n277), .A2(n71), .ZN(n281) );
  NAND3_X1 U260 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n12) );
  INV_X1 U261 ( .A(n31), .ZN(n291) );
  INV_X1 U262 ( .A(n21), .ZN(n288) );
  INV_X1 U263 ( .A(n321), .ZN(n289) );
  INV_X1 U264 ( .A(n332), .ZN(n286) );
  INV_X1 U265 ( .A(n301), .ZN(n294) );
  INV_X1 U266 ( .A(n310), .ZN(n292) );
  INV_X1 U267 ( .A(b[0]), .ZN(n284) );
  INV_X1 U268 ( .A(a[5]), .ZN(n290) );
  INV_X1 U269 ( .A(a[7]), .ZN(n287) );
  BUF_X1 U270 ( .A(n302), .Z(n282) );
  XNOR2_X1 U271 ( .A(a[2]), .B(a[1]), .ZN(n302) );
  INV_X1 U272 ( .A(a[3]), .ZN(n293) );
  NAND2_X2 U273 ( .A1(n312), .A2(n341), .ZN(n314) );
  INV_X1 U274 ( .A(a[1]), .ZN(n295) );
  XOR2_X2 U275 ( .A(a[6]), .B(n290), .Z(n323) );
  NOR2_X1 U276 ( .A1(n212), .A2(n284), .ZN(product[0]) );
  OAI22_X1 U277 ( .A1(n297), .A2(n298), .B1(n299), .B2(n212), .ZN(n99) );
  OAI22_X1 U278 ( .A1(n299), .A2(n298), .B1(n300), .B2(n212), .ZN(n98) );
  XNOR2_X1 U279 ( .A(b[6]), .B(n216), .ZN(n299) );
  OAI22_X1 U280 ( .A1(n212), .A2(n300), .B1(n298), .B2(n300), .ZN(n301) );
  XNOR2_X1 U281 ( .A(b[7]), .B(n216), .ZN(n300) );
  NOR2_X1 U282 ( .A1(n283), .A2(n284), .ZN(n96) );
  OAI22_X1 U283 ( .A1(n303), .A2(n304), .B1(n224), .B2(n305), .ZN(n95) );
  OAI22_X1 U284 ( .A1(n305), .A2(n304), .B1(n283), .B2(n306), .ZN(n94) );
  XNOR2_X1 U285 ( .A(b[1]), .B(n213), .ZN(n305) );
  OAI22_X1 U286 ( .A1(n306), .A2(n215), .B1(n283), .B2(n307), .ZN(n93) );
  XNOR2_X1 U287 ( .A(b[2]), .B(n213), .ZN(n306) );
  OAI22_X1 U288 ( .A1(n307), .A2(n215), .B1(n224), .B2(n308), .ZN(n92) );
  XNOR2_X1 U289 ( .A(b[3]), .B(n213), .ZN(n307) );
  OAI22_X1 U290 ( .A1(n308), .A2(n215), .B1(n224), .B2(n309), .ZN(n91) );
  XNOR2_X1 U291 ( .A(b[4]), .B(n213), .ZN(n308) );
  OAI22_X1 U292 ( .A1(n311), .A2(n283), .B1(n215), .B2(n311), .ZN(n310) );
  NOR2_X1 U293 ( .A1(n312), .A2(n284), .ZN(n88) );
  OAI22_X1 U294 ( .A1(n313), .A2(n314), .B1(n312), .B2(n315), .ZN(n87) );
  XNOR2_X1 U295 ( .A(a[5]), .B(n227), .ZN(n313) );
  OAI22_X1 U296 ( .A1(n315), .A2(n314), .B1(n312), .B2(n316), .ZN(n86) );
  XNOR2_X1 U297 ( .A(n206), .B(a[5]), .ZN(n315) );
  OAI22_X1 U298 ( .A1(n316), .A2(n314), .B1(n312), .B2(n317), .ZN(n85) );
  XNOR2_X1 U299 ( .A(b[2]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U300 ( .A1(n317), .A2(n314), .B1(n312), .B2(n318), .ZN(n84) );
  XNOR2_X1 U301 ( .A(b[3]), .B(a[5]), .ZN(n317) );
  OAI22_X1 U302 ( .A1(n318), .A2(n314), .B1(n312), .B2(n319), .ZN(n83) );
  XNOR2_X1 U303 ( .A(b[4]), .B(a[5]), .ZN(n318) );
  OAI22_X1 U304 ( .A1(n319), .A2(n314), .B1(n312), .B2(n320), .ZN(n82) );
  XNOR2_X1 U305 ( .A(b[5]), .B(a[5]), .ZN(n319) );
  OAI22_X1 U306 ( .A1(n322), .A2(n312), .B1(n314), .B2(n322), .ZN(n321) );
  NOR2_X1 U307 ( .A1(n323), .A2(n284), .ZN(n80) );
  OAI22_X1 U308 ( .A1(n324), .A2(n325), .B1(n323), .B2(n326), .ZN(n79) );
  XNOR2_X1 U309 ( .A(a[7]), .B(n238), .ZN(n324) );
  OAI22_X1 U310 ( .A1(n327), .A2(n325), .B1(n323), .B2(n328), .ZN(n77) );
  OAI22_X1 U311 ( .A1(n328), .A2(n325), .B1(n323), .B2(n329), .ZN(n76) );
  XNOR2_X1 U312 ( .A(b[3]), .B(a[7]), .ZN(n328) );
  OAI22_X1 U313 ( .A1(n329), .A2(n325), .B1(n323), .B2(n330), .ZN(n75) );
  XNOR2_X1 U314 ( .A(b[4]), .B(a[7]), .ZN(n329) );
  OAI22_X1 U315 ( .A1(n330), .A2(n325), .B1(n323), .B2(n331), .ZN(n74) );
  XNOR2_X1 U316 ( .A(b[5]), .B(a[7]), .ZN(n330) );
  OAI22_X1 U317 ( .A1(n333), .A2(n323), .B1(n325), .B2(n333), .ZN(n332) );
  OAI21_X1 U318 ( .B1(n227), .B2(n295), .A(n298), .ZN(n72) );
  OAI21_X1 U319 ( .B1(n293), .B2(n215), .A(n334), .ZN(n71) );
  OR3_X1 U320 ( .A1(n224), .A2(n227), .A3(n293), .ZN(n334) );
  OAI21_X1 U321 ( .B1(n290), .B2(n314), .A(n335), .ZN(n70) );
  OR3_X1 U322 ( .A1(n312), .A2(n227), .A3(n290), .ZN(n335) );
  OAI21_X1 U323 ( .B1(n287), .B2(n325), .A(n336), .ZN(n69) );
  OR3_X1 U324 ( .A1(n323), .A2(n238), .A3(n287), .ZN(n336) );
  XNOR2_X1 U325 ( .A(n337), .B(n338), .ZN(n38) );
  OR2_X1 U326 ( .A1(n337), .A2(n338), .ZN(n37) );
  OAI22_X1 U327 ( .A1(n309), .A2(n215), .B1(n224), .B2(n339), .ZN(n338) );
  XNOR2_X1 U328 ( .A(b[5]), .B(n213), .ZN(n309) );
  OAI22_X1 U329 ( .A1(n326), .A2(n325), .B1(n323), .B2(n327), .ZN(n337) );
  XNOR2_X1 U330 ( .A(b[2]), .B(a[7]), .ZN(n327) );
  XNOR2_X1 U331 ( .A(n206), .B(a[7]), .ZN(n326) );
  OAI22_X1 U332 ( .A1(n339), .A2(n215), .B1(n283), .B2(n311), .ZN(n31) );
  XNOR2_X1 U333 ( .A(b[7]), .B(n213), .ZN(n311) );
  XNOR2_X1 U334 ( .A(n293), .B(a[2]), .ZN(n340) );
  XNOR2_X1 U335 ( .A(b[6]), .B(n213), .ZN(n339) );
  OAI22_X1 U336 ( .A1(n320), .A2(n314), .B1(n312), .B2(n322), .ZN(n21) );
  XNOR2_X1 U337 ( .A(b[7]), .B(a[5]), .ZN(n322) );
  XNOR2_X1 U338 ( .A(b[6]), .B(a[5]), .ZN(n320) );
  OAI22_X1 U339 ( .A1(n331), .A2(n325), .B1(n323), .B2(n333), .ZN(n15) );
  XNOR2_X1 U340 ( .A(b[7]), .B(a[7]), .ZN(n333) );
  NAND2_X1 U341 ( .A1(n323), .A2(n342), .ZN(n325) );
  XNOR2_X1 U342 ( .A(n287), .B(a[6]), .ZN(n342) );
  XNOR2_X1 U343 ( .A(b[6]), .B(a[7]), .ZN(n331) );
  OAI22_X1 U344 ( .A1(n227), .A2(n298), .B1(n343), .B2(n296), .ZN(n104) );
  OAI22_X1 U345 ( .A1(n214), .A2(n298), .B1(n344), .B2(n296), .ZN(n103) );
  XNOR2_X1 U346 ( .A(b[1]), .B(a[1]), .ZN(n343) );
  OAI22_X1 U347 ( .A1(n344), .A2(n298), .B1(n345), .B2(n296), .ZN(n102) );
  XNOR2_X1 U348 ( .A(b[2]), .B(a[1]), .ZN(n344) );
  OAI22_X1 U349 ( .A1(n345), .A2(n298), .B1(n346), .B2(n296), .ZN(n101) );
  XNOR2_X1 U350 ( .A(b[3]), .B(a[1]), .ZN(n345) );
  OAI22_X1 U351 ( .A1(n346), .A2(n298), .B1(n297), .B2(n212), .ZN(n100) );
  XNOR2_X1 U352 ( .A(b[5]), .B(n216), .ZN(n297) );
  XNOR2_X1 U353 ( .A(b[4]), .B(n216), .ZN(n346) );
endmodule


module datapath_DW01_add_15 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n69;
  wire   [15:1] carry;

  FA_X1 U1_4 ( .A(B[4]), .B(A[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n69), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  XNOR2_X1 U1 ( .A(n2), .B(n1), .ZN(SUM[14]) );
  XNOR2_X1 U2 ( .A(B[14]), .B(A[14]), .ZN(n1) );
  XNOR2_X1 U3 ( .A(B[15]), .B(A[15]), .ZN(n59) );
  CLKBUF_X1 U4 ( .A(n15), .Z(n2) );
  XOR2_X1 U5 ( .A(carry[2]), .B(A[2]), .Z(n3) );
  XOR2_X1 U6 ( .A(B[2]), .B(n3), .Z(SUM[2]) );
  NAND2_X1 U7 ( .A1(carry[2]), .A2(B[2]), .ZN(n4) );
  NAND2_X1 U8 ( .A1(B[2]), .A2(A[2]), .ZN(n5) );
  NAND2_X1 U9 ( .A1(carry[2]), .A2(A[2]), .ZN(n6) );
  NAND3_X1 U10 ( .A1(n4), .A2(n5), .A3(n6), .ZN(carry[3]) );
  CLKBUF_X1 U11 ( .A(carry[5]), .Z(n7) );
  NAND3_X1 U12 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n8) );
  NAND3_X1 U13 ( .A1(n40), .A2(n41), .A3(n42), .ZN(n9) );
  CLKBUF_X1 U14 ( .A(n51), .Z(n10) );
  NAND3_X1 U15 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n11) );
  NAND3_X1 U16 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n12) );
  NAND3_X1 U17 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n13) );
  NAND3_X1 U18 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n14) );
  NAND3_X1 U19 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n15) );
  CLKBUF_X1 U20 ( .A(n11), .Z(n16) );
  NAND2_X1 U21 ( .A1(n15), .A2(B[14]), .ZN(n17) );
  NAND2_X1 U22 ( .A1(carry[14]), .A2(A[14]), .ZN(n18) );
  NAND2_X1 U23 ( .A1(B[14]), .A2(A[14]), .ZN(n19) );
  NAND3_X1 U24 ( .A1(n17), .A2(n18), .A3(n19), .ZN(carry[15]) );
  XOR2_X1 U25 ( .A(carry[3]), .B(A[3]), .Z(n20) );
  XOR2_X1 U26 ( .A(B[3]), .B(n20), .Z(SUM[3]) );
  NAND2_X1 U27 ( .A1(B[3]), .A2(carry[3]), .ZN(n21) );
  NAND2_X1 U28 ( .A1(B[3]), .A2(A[3]), .ZN(n22) );
  NAND2_X1 U29 ( .A1(carry[3]), .A2(A[3]), .ZN(n23) );
  NAND3_X1 U30 ( .A1(n21), .A2(n22), .A3(n23), .ZN(carry[4]) );
  CLKBUF_X1 U31 ( .A(n43), .Z(n24) );
  XOR2_X1 U32 ( .A(B[5]), .B(A[5]), .Z(n25) );
  XOR2_X1 U33 ( .A(n7), .B(n25), .Z(SUM[5]) );
  NAND2_X1 U34 ( .A1(carry[5]), .A2(B[5]), .ZN(n26) );
  NAND2_X1 U35 ( .A1(carry[5]), .A2(A[5]), .ZN(n27) );
  NAND2_X1 U36 ( .A1(B[5]), .A2(A[5]), .ZN(n28) );
  NAND3_X1 U37 ( .A1(n26), .A2(n27), .A3(n28), .ZN(carry[6]) );
  XOR2_X1 U38 ( .A(B[13]), .B(A[13]), .Z(n29) );
  XOR2_X1 U39 ( .A(n16), .B(n29), .Z(SUM[13]) );
  NAND2_X1 U40 ( .A1(B[13]), .A2(n11), .ZN(n30) );
  NAND2_X1 U41 ( .A1(carry[13]), .A2(A[13]), .ZN(n31) );
  NAND2_X1 U42 ( .A1(B[13]), .A2(A[13]), .ZN(n32) );
  NAND3_X1 U43 ( .A1(n31), .A2(n32), .A3(n30), .ZN(carry[14]) );
  XOR2_X1 U44 ( .A(B[6]), .B(A[6]), .Z(n33) );
  XOR2_X1 U45 ( .A(n8), .B(n33), .Z(SUM[6]) );
  NAND2_X1 U46 ( .A1(n8), .A2(B[6]), .ZN(n34) );
  NAND2_X1 U47 ( .A1(carry[6]), .A2(A[6]), .ZN(n35) );
  NAND2_X1 U48 ( .A1(B[6]), .A2(A[6]), .ZN(n36) );
  NAND3_X1 U49 ( .A1(n34), .A2(n35), .A3(n36), .ZN(carry[7]) );
  NAND3_X1 U50 ( .A1(n40), .A2(n41), .A3(n42), .ZN(n37) );
  CLKBUF_X1 U51 ( .A(carry[12]), .Z(n38) );
  XOR2_X1 U52 ( .A(B[7]), .B(A[7]), .Z(n39) );
  XOR2_X1 U53 ( .A(carry[7]), .B(n39), .Z(SUM[7]) );
  NAND2_X1 U54 ( .A1(carry[7]), .A2(B[7]), .ZN(n40) );
  NAND2_X1 U55 ( .A1(n14), .A2(A[7]), .ZN(n41) );
  NAND2_X1 U56 ( .A1(B[7]), .A2(A[7]), .ZN(n42) );
  NAND3_X1 U57 ( .A1(n40), .A2(n41), .A3(n42), .ZN(carry[8]) );
  NAND3_X1 U58 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n43) );
  XOR2_X1 U59 ( .A(B[8]), .B(A[8]), .Z(n44) );
  XOR2_X1 U60 ( .A(carry[8]), .B(n44), .Z(SUM[8]) );
  NAND2_X1 U61 ( .A1(n9), .A2(B[8]), .ZN(n45) );
  NAND2_X1 U62 ( .A1(n37), .A2(A[8]), .ZN(n46) );
  NAND2_X1 U63 ( .A1(B[8]), .A2(A[8]), .ZN(n47) );
  NAND3_X1 U64 ( .A1(n46), .A2(n45), .A3(n47), .ZN(carry[9]) );
  NAND3_X1 U65 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n48) );
  CLKBUF_X1 U66 ( .A(n13), .Z(n49) );
  XOR2_X1 U67 ( .A(B[10]), .B(A[10]), .Z(n50) );
  XOR2_X1 U68 ( .A(n49), .B(n50), .Z(SUM[10]) );
  NAND2_X1 U69 ( .A1(B[10]), .A2(n13), .ZN(n51) );
  NAND2_X1 U70 ( .A1(carry[10]), .A2(A[10]), .ZN(n52) );
  NAND2_X1 U71 ( .A1(B[10]), .A2(A[10]), .ZN(n53) );
  NAND3_X1 U72 ( .A1(n10), .A2(n52), .A3(n53), .ZN(carry[11]) );
  NAND3_X1 U73 ( .A1(n57), .A2(n56), .A3(n58), .ZN(n54) );
  XOR2_X1 U74 ( .A(B[11]), .B(A[11]), .Z(n55) );
  XOR2_X1 U75 ( .A(carry[11]), .B(n55), .Z(SUM[11]) );
  NAND2_X1 U76 ( .A1(n12), .A2(B[11]), .ZN(n56) );
  NAND2_X1 U77 ( .A1(n48), .A2(A[11]), .ZN(n57) );
  NAND2_X1 U78 ( .A1(B[11]), .A2(A[11]), .ZN(n58) );
  NAND3_X1 U79 ( .A1(n56), .A2(n57), .A3(n58), .ZN(carry[12]) );
  XNOR2_X1 U80 ( .A(carry[15]), .B(n59), .ZN(SUM[15]) );
  XOR2_X1 U81 ( .A(B[9]), .B(A[9]), .Z(n60) );
  XOR2_X1 U82 ( .A(n24), .B(n60), .Z(SUM[9]) );
  NAND2_X1 U83 ( .A1(n43), .A2(B[9]), .ZN(n61) );
  NAND2_X1 U84 ( .A1(carry[9]), .A2(A[9]), .ZN(n62) );
  NAND2_X1 U85 ( .A1(B[9]), .A2(A[9]), .ZN(n63) );
  NAND3_X1 U86 ( .A1(n61), .A2(n62), .A3(n63), .ZN(carry[10]) );
  XOR2_X1 U87 ( .A(B[12]), .B(A[12]), .Z(n64) );
  XOR2_X1 U88 ( .A(n38), .B(n64), .Z(SUM[12]) );
  NAND2_X1 U89 ( .A1(carry[12]), .A2(B[12]), .ZN(n65) );
  NAND2_X1 U90 ( .A1(n54), .A2(A[12]), .ZN(n66) );
  NAND2_X1 U91 ( .A1(B[12]), .A2(A[12]), .ZN(n67) );
  NAND3_X1 U92 ( .A1(n65), .A2(n66), .A3(n67), .ZN(carry[13]) );
  XOR2_X1 U93 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U94 ( .A1(B[0]), .A2(A[0]), .ZN(n69) );
endmodule


module datapath_DW_mult_tc_14 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n296), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n295), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n299), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n298), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n301), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n207), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  BUF_X2 U157 ( .A(a[5]), .Z(n233) );
  AND3_X1 U158 ( .A1(n282), .A2(n283), .A3(n284), .ZN(product[15]) );
  AND2_X1 U159 ( .A1(n87), .A2(n70), .ZN(n207) );
  NAND3_X1 U160 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n208) );
  NAND3_X1 U161 ( .A1(n276), .A2(n275), .A3(n277), .ZN(n209) );
  XNOR2_X1 U162 ( .A(n250), .B(n210), .ZN(product[10]) );
  XNOR2_X1 U163 ( .A(n27), .B(n24), .ZN(n210) );
  NAND2_X2 U164 ( .A1(a[1]), .A2(n303), .ZN(n305) );
  XNOR2_X1 U165 ( .A(a[4]), .B(a[3]), .ZN(n319) );
  NAND2_X2 U166 ( .A1(n309), .A2(n347), .ZN(n311) );
  XNOR2_X2 U167 ( .A(a[2]), .B(a[1]), .ZN(n287) );
  OAI22_X1 U168 ( .A1(n274), .A2(n305), .B1(n351), .B2(n303), .ZN(n211) );
  XNOR2_X1 U169 ( .A(n288), .B(n262), .ZN(n212) );
  XNOR2_X1 U170 ( .A(n213), .B(n2), .ZN(product[14]) );
  XNOR2_X1 U171 ( .A(n293), .B(n15), .ZN(n213) );
  OAI22_X1 U172 ( .A1(n212), .A2(n311), .B1(n287), .B2(n312), .ZN(n214) );
  XNOR2_X1 U173 ( .A(n219), .B(n215), .ZN(product[5]) );
  XNOR2_X1 U174 ( .A(n50), .B(n53), .ZN(n215) );
  NAND3_X1 U175 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n216) );
  NAND3_X1 U176 ( .A1(n222), .A2(n223), .A3(n224), .ZN(n217) );
  NAND3_X1 U177 ( .A1(n268), .A2(n269), .A3(n267), .ZN(n218) );
  NAND3_X1 U178 ( .A1(n268), .A2(n269), .A3(n267), .ZN(n219) );
  NAND3_X1 U179 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n220) );
  XOR2_X1 U180 ( .A(n23), .B(n20), .Z(n221) );
  XOR2_X1 U181 ( .A(n209), .B(n221), .Z(product[11]) );
  NAND2_X1 U182 ( .A1(n209), .A2(n23), .ZN(n222) );
  NAND2_X1 U183 ( .A1(n5), .A2(n20), .ZN(n223) );
  NAND2_X1 U184 ( .A1(n23), .A2(n20), .ZN(n224) );
  NAND3_X1 U185 ( .A1(n222), .A2(n223), .A3(n224), .ZN(n4) );
  NAND2_X1 U186 ( .A1(n218), .A2(n50), .ZN(n225) );
  NAND2_X1 U187 ( .A1(n11), .A2(n53), .ZN(n226) );
  NAND2_X1 U188 ( .A1(n50), .A2(n53), .ZN(n227) );
  NAND3_X1 U189 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n10) );
  NAND3_X1 U190 ( .A1(n237), .A2(n236), .A3(n238), .ZN(n228) );
  XOR2_X1 U191 ( .A(n70), .B(n87), .Z(n52) );
  CLKBUF_X1 U192 ( .A(n208), .Z(n229) );
  NAND3_X1 U193 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n230) );
  NAND3_X1 U194 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n231) );
  XNOR2_X1 U195 ( .A(n232), .B(n229), .ZN(product[3]) );
  XNOR2_X1 U196 ( .A(n56), .B(n71), .ZN(n232) );
  NAND2_X1 U197 ( .A1(n319), .A2(n348), .ZN(n321) );
  XNOR2_X1 U198 ( .A(n262), .B(n288), .ZN(n310) );
  XNOR2_X1 U199 ( .A(n14), .B(n234), .ZN(product[2]) );
  XNOR2_X1 U200 ( .A(n103), .B(n96), .ZN(n234) );
  XOR2_X1 U201 ( .A(n18), .B(n19), .Z(n235) );
  XOR2_X1 U202 ( .A(n217), .B(n235), .Z(product[12]) );
  NAND2_X1 U203 ( .A1(n217), .A2(n18), .ZN(n236) );
  NAND2_X1 U204 ( .A1(n4), .A2(n19), .ZN(n237) );
  NAND2_X1 U205 ( .A1(n18), .A2(n19), .ZN(n238) );
  NAND3_X1 U206 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n3) );
  NAND2_X1 U207 ( .A1(n14), .A2(n103), .ZN(n239) );
  NAND2_X1 U208 ( .A1(n14), .A2(n96), .ZN(n240) );
  NAND2_X1 U209 ( .A1(n211), .A2(n96), .ZN(n241) );
  NAND3_X1 U210 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n13) );
  NAND3_X1 U211 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n242) );
  XOR2_X1 U212 ( .A(n34), .B(n39), .Z(n243) );
  XOR2_X1 U213 ( .A(n231), .B(n243), .Z(product[8]) );
  NAND2_X1 U214 ( .A1(n230), .A2(n34), .ZN(n244) );
  NAND2_X1 U215 ( .A1(n8), .A2(n39), .ZN(n245) );
  NAND2_X1 U216 ( .A1(n34), .A2(n39), .ZN(n246) );
  NAND3_X1 U217 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n7) );
  NAND3_X1 U218 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n247) );
  NAND3_X1 U219 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n248) );
  NAND3_X1 U220 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n249) );
  NAND3_X1 U221 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n250) );
  XOR2_X1 U222 ( .A(n214), .B(n102), .Z(n251) );
  XOR2_X1 U223 ( .A(n46), .B(n49), .Z(n252) );
  XOR2_X1 U224 ( .A(n10), .B(n252), .Z(product[6]) );
  NAND2_X1 U225 ( .A1(n220), .A2(n46), .ZN(n253) );
  NAND2_X1 U226 ( .A1(n10), .A2(n49), .ZN(n254) );
  NAND2_X1 U227 ( .A1(n46), .A2(n49), .ZN(n255) );
  NAND3_X1 U228 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n9) );
  XOR2_X1 U229 ( .A(n33), .B(n28), .Z(n256) );
  XOR2_X1 U230 ( .A(n242), .B(n256), .Z(product[9]) );
  NAND2_X1 U231 ( .A1(n242), .A2(n33), .ZN(n257) );
  NAND2_X1 U232 ( .A1(n7), .A2(n28), .ZN(n258) );
  NAND2_X1 U233 ( .A1(n33), .A2(n28), .ZN(n259) );
  NAND3_X1 U234 ( .A1(n265), .A2(n264), .A3(n263), .ZN(n260) );
  NAND3_X1 U235 ( .A1(n263), .A2(n264), .A3(n265), .ZN(n261) );
  BUF_X2 U236 ( .A(n291), .Z(n262) );
  NAND2_X1 U237 ( .A1(n251), .A2(n71), .ZN(n263) );
  NAND2_X1 U238 ( .A1(n251), .A2(n13), .ZN(n264) );
  NAND2_X1 U239 ( .A1(n71), .A2(n208), .ZN(n265) );
  NAND3_X1 U240 ( .A1(n263), .A2(n264), .A3(n265), .ZN(n12) );
  XOR2_X1 U241 ( .A(n54), .B(n55), .Z(n266) );
  XOR2_X1 U242 ( .A(n266), .B(n261), .Z(product[4]) );
  NAND2_X1 U243 ( .A1(n54), .A2(n55), .ZN(n267) );
  NAND2_X1 U244 ( .A1(n260), .A2(n54), .ZN(n268) );
  NAND2_X1 U245 ( .A1(n12), .A2(n55), .ZN(n269) );
  NAND3_X1 U246 ( .A1(n268), .A2(n269), .A3(n267), .ZN(n11) );
  XOR2_X1 U247 ( .A(n40), .B(n45), .Z(n270) );
  XOR2_X1 U248 ( .A(n248), .B(n270), .Z(product[7]) );
  NAND2_X1 U249 ( .A1(n247), .A2(n40), .ZN(n271) );
  NAND2_X1 U250 ( .A1(n9), .A2(n45), .ZN(n272) );
  NAND2_X1 U251 ( .A1(n40), .A2(n45), .ZN(n273) );
  NAND3_X1 U252 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n8) );
  BUF_X1 U253 ( .A(n350), .Z(n274) );
  NAND2_X1 U254 ( .A1(n249), .A2(n27), .ZN(n275) );
  NAND2_X1 U255 ( .A1(n249), .A2(n24), .ZN(n276) );
  NAND2_X1 U256 ( .A1(n27), .A2(n24), .ZN(n277) );
  NAND3_X1 U257 ( .A1(n276), .A2(n275), .A3(n277), .ZN(n5) );
  INV_X1 U258 ( .A(b[0]), .ZN(n291) );
  INV_X2 U259 ( .A(n291), .ZN(n290) );
  XOR2_X1 U260 ( .A(n17), .B(n292), .Z(n278) );
  XOR2_X1 U261 ( .A(n278), .B(n228), .Z(product[13]) );
  NAND2_X1 U262 ( .A1(n17), .A2(n292), .ZN(n279) );
  NAND2_X1 U263 ( .A1(n17), .A2(n216), .ZN(n280) );
  NAND2_X1 U264 ( .A1(n292), .A2(n3), .ZN(n281) );
  NAND3_X1 U265 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n2) );
  NAND2_X1 U266 ( .A1(n293), .A2(n15), .ZN(n282) );
  NAND2_X1 U267 ( .A1(n293), .A2(n2), .ZN(n283) );
  NAND2_X1 U268 ( .A1(n15), .A2(n2), .ZN(n284) );
  INV_X1 U269 ( .A(n319), .ZN(n285) );
  INV_X2 U270 ( .A(n285), .ZN(n286) );
  INV_X1 U271 ( .A(n15), .ZN(n292) );
  INV_X1 U272 ( .A(n317), .ZN(n299) );
  INV_X1 U273 ( .A(n31), .ZN(n298) );
  INV_X1 U274 ( .A(n21), .ZN(n295) );
  INV_X1 U275 ( .A(n328), .ZN(n296) );
  INV_X1 U276 ( .A(n339), .ZN(n293) );
  INV_X1 U277 ( .A(n308), .ZN(n301) );
  INV_X1 U278 ( .A(a[5]), .ZN(n297) );
  INV_X1 U279 ( .A(a[7]), .ZN(n294) );
  XNOR2_X1 U280 ( .A(a[2]), .B(a[1]), .ZN(n309) );
  INV_X1 U281 ( .A(a[3]), .ZN(n288) );
  INV_X2 U282 ( .A(n288), .ZN(n289) );
  INV_X1 U283 ( .A(a[3]), .ZN(n300) );
  INV_X1 U284 ( .A(a[1]), .ZN(n302) );
  XOR2_X2 U285 ( .A(a[6]), .B(n297), .Z(n330) );
  INV_X2 U286 ( .A(a[0]), .ZN(n303) );
  NOR2_X1 U287 ( .A1(n303), .A2(n262), .ZN(product[0]) );
  OAI22_X1 U288 ( .A1(n304), .A2(n305), .B1(n306), .B2(n303), .ZN(n99) );
  OAI22_X1 U289 ( .A1(n306), .A2(n305), .B1(n307), .B2(n303), .ZN(n98) );
  XNOR2_X1 U290 ( .A(b[6]), .B(a[1]), .ZN(n306) );
  OAI22_X1 U291 ( .A1(n303), .A2(n307), .B1(n305), .B2(n307), .ZN(n308) );
  XNOR2_X1 U292 ( .A(b[7]), .B(a[1]), .ZN(n307) );
  NOR2_X1 U293 ( .A1(n287), .A2(n262), .ZN(n96) );
  OAI22_X1 U294 ( .A1(n310), .A2(n311), .B1(n287), .B2(n312), .ZN(n95) );
  OAI22_X1 U295 ( .A1(n312), .A2(n311), .B1(n287), .B2(n313), .ZN(n94) );
  XNOR2_X1 U296 ( .A(b[1]), .B(n289), .ZN(n312) );
  OAI22_X1 U297 ( .A1(n313), .A2(n311), .B1(n287), .B2(n314), .ZN(n93) );
  XNOR2_X1 U298 ( .A(b[2]), .B(n289), .ZN(n313) );
  OAI22_X1 U299 ( .A1(n314), .A2(n311), .B1(n287), .B2(n315), .ZN(n92) );
  XNOR2_X1 U300 ( .A(b[3]), .B(n289), .ZN(n314) );
  OAI22_X1 U301 ( .A1(n315), .A2(n311), .B1(n287), .B2(n316), .ZN(n91) );
  XNOR2_X1 U302 ( .A(b[4]), .B(n289), .ZN(n315) );
  OAI22_X1 U303 ( .A1(n318), .A2(n287), .B1(n311), .B2(n318), .ZN(n317) );
  NOR2_X1 U304 ( .A1(n319), .A2(n262), .ZN(n88) );
  OAI22_X1 U305 ( .A1(n320), .A2(n321), .B1(n286), .B2(n322), .ZN(n87) );
  XNOR2_X1 U306 ( .A(n233), .B(n290), .ZN(n320) );
  OAI22_X1 U307 ( .A1(n322), .A2(n321), .B1(n286), .B2(n323), .ZN(n86) );
  XNOR2_X1 U308 ( .A(b[1]), .B(n233), .ZN(n322) );
  OAI22_X1 U309 ( .A1(n323), .A2(n321), .B1(n286), .B2(n324), .ZN(n85) );
  XNOR2_X1 U310 ( .A(b[2]), .B(n233), .ZN(n323) );
  OAI22_X1 U311 ( .A1(n324), .A2(n321), .B1(n286), .B2(n325), .ZN(n84) );
  XNOR2_X1 U312 ( .A(b[3]), .B(n233), .ZN(n324) );
  OAI22_X1 U313 ( .A1(n325), .A2(n321), .B1(n286), .B2(n326), .ZN(n83) );
  XNOR2_X1 U314 ( .A(b[4]), .B(n233), .ZN(n325) );
  OAI22_X1 U315 ( .A1(n326), .A2(n321), .B1(n286), .B2(n327), .ZN(n82) );
  XNOR2_X1 U316 ( .A(b[5]), .B(n233), .ZN(n326) );
  OAI22_X1 U317 ( .A1(n329), .A2(n286), .B1(n321), .B2(n329), .ZN(n328) );
  NOR2_X1 U318 ( .A1(n330), .A2(n262), .ZN(n80) );
  OAI22_X1 U319 ( .A1(n331), .A2(n332), .B1(n330), .B2(n333), .ZN(n79) );
  XNOR2_X1 U320 ( .A(a[7]), .B(n290), .ZN(n331) );
  OAI22_X1 U321 ( .A1(n334), .A2(n332), .B1(n330), .B2(n335), .ZN(n77) );
  OAI22_X1 U322 ( .A1(n335), .A2(n332), .B1(n330), .B2(n336), .ZN(n76) );
  XNOR2_X1 U323 ( .A(b[3]), .B(a[7]), .ZN(n335) );
  OAI22_X1 U324 ( .A1(n336), .A2(n332), .B1(n330), .B2(n337), .ZN(n75) );
  XNOR2_X1 U325 ( .A(b[4]), .B(a[7]), .ZN(n336) );
  OAI22_X1 U326 ( .A1(n337), .A2(n332), .B1(n330), .B2(n338), .ZN(n74) );
  XNOR2_X1 U327 ( .A(b[5]), .B(a[7]), .ZN(n337) );
  OAI22_X1 U328 ( .A1(n340), .A2(n330), .B1(n332), .B2(n340), .ZN(n339) );
  OAI21_X1 U329 ( .B1(n290), .B2(n302), .A(n305), .ZN(n72) );
  OAI21_X1 U330 ( .B1(n300), .B2(n311), .A(n341), .ZN(n71) );
  OR3_X1 U331 ( .A1(n287), .A2(n290), .A3(n300), .ZN(n341) );
  OAI21_X1 U332 ( .B1(n297), .B2(n321), .A(n342), .ZN(n70) );
  OR3_X1 U333 ( .A1(n319), .A2(n290), .A3(n297), .ZN(n342) );
  OAI21_X1 U334 ( .B1(n294), .B2(n332), .A(n343), .ZN(n69) );
  OR3_X1 U335 ( .A1(n330), .A2(n290), .A3(n294), .ZN(n343) );
  XNOR2_X1 U336 ( .A(n344), .B(n345), .ZN(n38) );
  OR2_X1 U337 ( .A1(n344), .A2(n345), .ZN(n37) );
  OAI22_X1 U338 ( .A1(n316), .A2(n311), .B1(n287), .B2(n346), .ZN(n345) );
  XNOR2_X1 U339 ( .A(b[5]), .B(n289), .ZN(n316) );
  OAI22_X1 U340 ( .A1(n333), .A2(n332), .B1(n330), .B2(n334), .ZN(n344) );
  XNOR2_X1 U341 ( .A(b[2]), .B(a[7]), .ZN(n334) );
  XNOR2_X1 U342 ( .A(b[1]), .B(a[7]), .ZN(n333) );
  OAI22_X1 U343 ( .A1(n346), .A2(n311), .B1(n287), .B2(n318), .ZN(n31) );
  XNOR2_X1 U344 ( .A(b[7]), .B(n289), .ZN(n318) );
  XNOR2_X1 U345 ( .A(n300), .B(a[2]), .ZN(n347) );
  XNOR2_X1 U346 ( .A(b[6]), .B(n289), .ZN(n346) );
  OAI22_X1 U347 ( .A1(n327), .A2(n321), .B1(n286), .B2(n329), .ZN(n21) );
  XNOR2_X1 U348 ( .A(b[7]), .B(n233), .ZN(n329) );
  XNOR2_X1 U349 ( .A(n297), .B(a[4]), .ZN(n348) );
  XNOR2_X1 U350 ( .A(b[6]), .B(n233), .ZN(n327) );
  OAI22_X1 U351 ( .A1(n338), .A2(n332), .B1(n330), .B2(n340), .ZN(n15) );
  XNOR2_X1 U352 ( .A(b[7]), .B(a[7]), .ZN(n340) );
  NAND2_X1 U353 ( .A1(n330), .A2(n349), .ZN(n332) );
  XNOR2_X1 U354 ( .A(n294), .B(a[6]), .ZN(n349) );
  XNOR2_X1 U355 ( .A(b[6]), .B(a[7]), .ZN(n338) );
  OAI22_X1 U356 ( .A1(n290), .A2(n305), .B1(n350), .B2(n303), .ZN(n104) );
  OAI22_X1 U357 ( .A1(n274), .A2(n305), .B1(n351), .B2(n303), .ZN(n103) );
  XNOR2_X1 U358 ( .A(b[1]), .B(a[1]), .ZN(n350) );
  OAI22_X1 U359 ( .A1(n351), .A2(n305), .B1(n352), .B2(n303), .ZN(n102) );
  XNOR2_X1 U360 ( .A(b[2]), .B(a[1]), .ZN(n351) );
  OAI22_X1 U361 ( .A1(n352), .A2(n305), .B1(n353), .B2(n303), .ZN(n101) );
  XNOR2_X1 U362 ( .A(b[3]), .B(a[1]), .ZN(n352) );
  OAI22_X1 U363 ( .A1(n353), .A2(n305), .B1(n304), .B2(n303), .ZN(n100) );
  XNOR2_X1 U364 ( .A(b[5]), .B(a[1]), .ZN(n304) );
  XNOR2_X1 U365 ( .A(b[4]), .B(a[1]), .ZN(n353) );
endmodule


module datapath_DW01_add_14 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n75;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n75), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(carry[2]), .Z(n1) );
  XNOR2_X1 U2 ( .A(B[15]), .B(A[15]), .ZN(n38) );
  CLKBUF_X1 U3 ( .A(n55), .Z(n2) );
  CLKBUF_X1 U4 ( .A(carry[7]), .Z(n3) );
  CLKBUF_X1 U5 ( .A(B[4]), .Z(n4) );
  CLKBUF_X1 U6 ( .A(n40), .Z(n5) );
  NAND3_X1 U7 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n6) );
  NAND3_X1 U8 ( .A1(n53), .A2(n54), .A3(n2), .ZN(n7) );
  NAND3_X1 U9 ( .A1(n13), .A2(n14), .A3(n15), .ZN(n8) );
  NAND3_X1 U10 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n9) );
  NAND3_X1 U11 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n10) );
  NAND3_X1 U12 ( .A1(n5), .A2(n41), .A3(n42), .ZN(n11) );
  XOR2_X1 U13 ( .A(n11), .B(A[11]), .Z(n12) );
  XOR2_X1 U14 ( .A(B[11]), .B(n12), .Z(SUM[11]) );
  NAND2_X1 U15 ( .A1(B[11]), .A2(carry[11]), .ZN(n13) );
  NAND2_X1 U16 ( .A1(B[11]), .A2(A[11]), .ZN(n14) );
  NAND2_X1 U17 ( .A1(carry[11]), .A2(A[11]), .ZN(n15) );
  NAND3_X1 U18 ( .A1(n13), .A2(n15), .A3(n14), .ZN(carry[12]) );
  NAND3_X1 U19 ( .A1(n44), .A2(n45), .A3(n46), .ZN(n16) );
  XOR2_X1 U20 ( .A(n7), .B(A[5]), .Z(n17) );
  XOR2_X1 U21 ( .A(B[5]), .B(n17), .Z(SUM[5]) );
  NAND2_X1 U22 ( .A1(B[5]), .A2(n6), .ZN(n18) );
  NAND2_X1 U23 ( .A1(B[5]), .A2(A[5]), .ZN(n19) );
  NAND2_X1 U24 ( .A1(carry[5]), .A2(A[5]), .ZN(n20) );
  NAND3_X1 U25 ( .A1(n18), .A2(n19), .A3(n20), .ZN(carry[6]) );
  NAND3_X1 U26 ( .A1(n26), .A2(n25), .A3(n27), .ZN(n21) );
  CLKBUF_X1 U27 ( .A(n45), .Z(n22) );
  NAND3_X1 U28 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n23) );
  XOR2_X1 U29 ( .A(B[7]), .B(A[7]), .Z(n24) );
  XOR2_X1 U30 ( .A(n3), .B(n24), .Z(SUM[7]) );
  NAND2_X1 U31 ( .A1(n23), .A2(B[7]), .ZN(n25) );
  NAND2_X1 U32 ( .A1(carry[7]), .A2(A[7]), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[7]), .A2(A[7]), .ZN(n27) );
  NAND3_X1 U34 ( .A1(n26), .A2(n25), .A3(n27), .ZN(carry[8]) );
  NAND3_X1 U35 ( .A1(n63), .A2(n65), .A3(n64), .ZN(n28) );
  XOR2_X1 U36 ( .A(B[6]), .B(A[6]), .Z(n29) );
  XOR2_X1 U37 ( .A(n10), .B(n29), .Z(SUM[6]) );
  NAND2_X1 U38 ( .A1(n9), .A2(B[6]), .ZN(n30) );
  NAND2_X1 U39 ( .A1(carry[6]), .A2(A[6]), .ZN(n31) );
  NAND2_X1 U40 ( .A1(B[6]), .A2(A[6]), .ZN(n32) );
  NAND3_X1 U41 ( .A1(n30), .A2(n31), .A3(n32), .ZN(carry[7]) );
  CLKBUF_X1 U42 ( .A(n35), .Z(n33) );
  CLKBUF_X1 U43 ( .A(n47), .Z(n34) );
  NAND3_X1 U44 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n35) );
  NAND3_X1 U45 ( .A1(n44), .A2(n45), .A3(n46), .ZN(n36) );
  CLKBUF_X1 U46 ( .A(carry[12]), .Z(n37) );
  XNOR2_X1 U47 ( .A(carry[15]), .B(n38), .ZN(SUM[15]) );
  XOR2_X1 U48 ( .A(B[10]), .B(A[10]), .Z(n39) );
  XOR2_X1 U49 ( .A(n33), .B(n39), .Z(SUM[10]) );
  NAND2_X1 U50 ( .A1(n35), .A2(B[10]), .ZN(n40) );
  NAND2_X1 U51 ( .A1(carry[10]), .A2(A[10]), .ZN(n41) );
  NAND2_X1 U52 ( .A1(B[10]), .A2(A[10]), .ZN(n42) );
  NAND3_X1 U53 ( .A1(n40), .A2(n41), .A3(n42), .ZN(carry[11]) );
  XOR2_X1 U54 ( .A(B[8]), .B(A[8]), .Z(n43) );
  XOR2_X1 U55 ( .A(carry[8]), .B(n43), .Z(SUM[8]) );
  NAND2_X1 U56 ( .A1(n21), .A2(B[8]), .ZN(n44) );
  NAND2_X1 U57 ( .A1(n21), .A2(A[8]), .ZN(n45) );
  NAND2_X1 U58 ( .A1(B[8]), .A2(A[8]), .ZN(n46) );
  NAND3_X1 U59 ( .A1(n44), .A2(n22), .A3(n46), .ZN(carry[9]) );
  NAND3_X1 U60 ( .A1(n69), .A2(n68), .A3(n67), .ZN(n47) );
  XOR2_X1 U61 ( .A(B[9]), .B(A[9]), .Z(n48) );
  XOR2_X1 U62 ( .A(carry[9]), .B(n48), .Z(SUM[9]) );
  NAND2_X1 U63 ( .A1(n16), .A2(B[9]), .ZN(n49) );
  NAND2_X1 U64 ( .A1(n36), .A2(A[9]), .ZN(n50) );
  NAND2_X1 U65 ( .A1(B[9]), .A2(A[9]), .ZN(n51) );
  NAND3_X1 U66 ( .A1(n50), .A2(n49), .A3(n51), .ZN(carry[10]) );
  XOR2_X1 U67 ( .A(n4), .B(A[4]), .Z(n52) );
  XOR2_X1 U68 ( .A(carry[4]), .B(n52), .Z(SUM[4]) );
  NAND2_X1 U69 ( .A1(B[4]), .A2(n28), .ZN(n53) );
  NAND2_X1 U70 ( .A1(carry[4]), .A2(A[4]), .ZN(n54) );
  NAND2_X1 U71 ( .A1(B[4]), .A2(A[4]), .ZN(n55) );
  NAND3_X1 U72 ( .A1(n53), .A2(n54), .A3(n55), .ZN(carry[5]) );
  NAND3_X1 U73 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n56) );
  NAND3_X1 U74 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n57) );
  XOR2_X1 U75 ( .A(A[2]), .B(B[2]), .Z(n58) );
  XOR2_X1 U76 ( .A(n58), .B(n1), .Z(SUM[2]) );
  NAND2_X1 U77 ( .A1(A[2]), .A2(B[2]), .ZN(n59) );
  NAND2_X1 U78 ( .A1(A[2]), .A2(carry[2]), .ZN(n60) );
  NAND2_X1 U79 ( .A1(B[2]), .A2(carry[2]), .ZN(n61) );
  NAND3_X1 U80 ( .A1(n59), .A2(n60), .A3(n61), .ZN(carry[3]) );
  XOR2_X1 U81 ( .A(A[3]), .B(B[3]), .Z(n62) );
  XOR2_X1 U82 ( .A(n62), .B(n57), .Z(SUM[3]) );
  NAND2_X1 U83 ( .A1(A[3]), .A2(B[3]), .ZN(n63) );
  NAND2_X1 U84 ( .A1(A[3]), .A2(n56), .ZN(n64) );
  NAND2_X1 U85 ( .A1(B[3]), .A2(carry[3]), .ZN(n65) );
  NAND3_X1 U86 ( .A1(n63), .A2(n65), .A3(n64), .ZN(carry[4]) );
  XOR2_X1 U87 ( .A(A[12]), .B(B[12]), .Z(n66) );
  XOR2_X1 U88 ( .A(n66), .B(n37), .Z(SUM[12]) );
  NAND2_X1 U89 ( .A1(A[12]), .A2(B[12]), .ZN(n67) );
  NAND2_X1 U90 ( .A1(A[12]), .A2(n8), .ZN(n68) );
  NAND2_X1 U91 ( .A1(carry[12]), .A2(B[12]), .ZN(n69) );
  NAND3_X1 U92 ( .A1(n67), .A2(n68), .A3(n69), .ZN(carry[13]) );
  XOR2_X1 U93 ( .A(A[13]), .B(B[13]), .Z(n70) );
  XOR2_X1 U94 ( .A(n70), .B(n34), .Z(SUM[13]) );
  NAND2_X1 U95 ( .A1(A[13]), .A2(B[13]), .ZN(n71) );
  NAND2_X1 U96 ( .A1(A[13]), .A2(carry[13]), .ZN(n72) );
  NAND2_X1 U97 ( .A1(n47), .A2(B[13]), .ZN(n73) );
  NAND3_X1 U98 ( .A1(n73), .A2(n72), .A3(n71), .ZN(carry[14]) );
  XOR2_X1 U99 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U100 ( .A1(B[0]), .A2(A[0]), .ZN(n75) );
endmodule


module datapath_DW_mult_tc_13 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345;

  FA_X1 U12 ( .A(n54), .B(n206), .CI(n12), .CO(n11), .S(product[4]) );
  FA_X1 U13 ( .A(n13), .B(n71), .CI(n56), .CO(n12), .S(product[3]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n288), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n287), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n291), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n290), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n293), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  NAND2_X2 U157 ( .A1(n311), .A2(n340), .ZN(n313) );
  AND2_X1 U158 ( .A1(n95), .A2(n102), .ZN(n206) );
  XNOR2_X1 U159 ( .A(n17), .B(n284), .ZN(n207) );
  AND3_X1 U160 ( .A1(n260), .A2(n261), .A3(n262), .ZN(product[15]) );
  NAND3_X1 U161 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n209) );
  NAND2_X1 U162 ( .A1(n4), .A2(n19), .ZN(n210) );
  NAND2_X2 U163 ( .A1(n322), .A2(n341), .ZN(n324) );
  CLKBUF_X1 U164 ( .A(b[1]), .Z(n211) );
  NAND2_X2 U165 ( .A1(a[1]), .A2(n295), .ZN(n297) );
  NAND3_X1 U166 ( .A1(n249), .A2(n250), .A3(n248), .ZN(n212) );
  CLKBUF_X3 U167 ( .A(a[1]), .Z(n281) );
  NAND2_X1 U168 ( .A1(n301), .A2(n339), .ZN(n213) );
  XOR2_X1 U169 ( .A(n95), .B(n102), .Z(n56) );
  NAND2_X1 U170 ( .A1(n301), .A2(n339), .ZN(n303) );
  NAND2_X2 U171 ( .A1(n278), .A2(n279), .ZN(n214) );
  NAND2_X1 U172 ( .A1(n278), .A2(n279), .ZN(n311) );
  XOR2_X1 U173 ( .A(a[3]), .B(a[2]), .Z(n339) );
  AND2_X1 U174 ( .A1(n104), .A2(n72), .ZN(n215) );
  XNOR2_X1 U175 ( .A(n207), .B(n220), .ZN(product[13]) );
  OAI22_X1 U176 ( .A1(n275), .A2(n297), .B1(n343), .B2(n295), .ZN(n216) );
  CLKBUF_X1 U177 ( .A(n11), .Z(n217) );
  BUF_X2 U178 ( .A(n280), .Z(n218) );
  XNOR2_X1 U179 ( .A(a[2]), .B(n281), .ZN(n280) );
  XNOR2_X1 U180 ( .A(n247), .B(n219), .ZN(product[11]) );
  AND3_X1 U181 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n219) );
  NAND3_X1 U182 ( .A1(n210), .A2(n230), .A3(n232), .ZN(n220) );
  XNOR2_X1 U183 ( .A(n217), .B(n221), .ZN(product[5]) );
  XNOR2_X1 U184 ( .A(n50), .B(n53), .ZN(n221) );
  NAND3_X1 U185 ( .A1(n249), .A2(n250), .A3(n248), .ZN(n222) );
  NAND3_X1 U186 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n223) );
  NAND3_X1 U187 ( .A1(n274), .A2(n272), .A3(n273), .ZN(n224) );
  NAND3_X1 U188 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n225) );
  NAND3_X1 U189 ( .A1(n230), .A2(n231), .A3(n232), .ZN(n226) );
  NAND3_X1 U190 ( .A1(n270), .A2(n269), .A3(n268), .ZN(n227) );
  NAND3_X1 U191 ( .A1(n269), .A2(n270), .A3(n268), .ZN(n228) );
  XOR2_X1 U192 ( .A(n18), .B(n19), .Z(n229) );
  XOR2_X1 U193 ( .A(n212), .B(n229), .Z(product[12]) );
  NAND2_X1 U194 ( .A1(n222), .A2(n18), .ZN(n230) );
  NAND2_X1 U195 ( .A1(n4), .A2(n19), .ZN(n231) );
  NAND2_X1 U196 ( .A1(n18), .A2(n19), .ZN(n232) );
  NAND3_X1 U197 ( .A1(n210), .A2(n230), .A3(n232), .ZN(n3) );
  NAND2_X1 U198 ( .A1(n11), .A2(n50), .ZN(n233) );
  NAND2_X1 U199 ( .A1(n11), .A2(n53), .ZN(n234) );
  NAND2_X1 U200 ( .A1(n50), .A2(n53), .ZN(n235) );
  NAND3_X1 U201 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n10) );
  NAND3_X1 U202 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n236) );
  NAND3_X1 U203 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n237) );
  NAND3_X1 U204 ( .A1(n246), .A2(n245), .A3(n244), .ZN(n238) );
  XOR2_X1 U205 ( .A(n216), .B(n96), .Z(n239) );
  XOR2_X1 U206 ( .A(n215), .B(n239), .Z(product[2]) );
  NAND2_X1 U207 ( .A1(n215), .A2(n96), .ZN(n240) );
  NAND2_X1 U208 ( .A1(n14), .A2(n103), .ZN(n241) );
  NAND2_X1 U209 ( .A1(n96), .A2(n103), .ZN(n242) );
  NAND3_X1 U210 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n13) );
  XOR2_X1 U211 ( .A(n24), .B(n27), .Z(n243) );
  XOR2_X1 U212 ( .A(n243), .B(n225), .Z(product[10]) );
  NAND2_X1 U213 ( .A1(n24), .A2(n27), .ZN(n244) );
  NAND2_X1 U214 ( .A1(n24), .A2(n6), .ZN(n245) );
  NAND2_X1 U215 ( .A1(n27), .A2(n224), .ZN(n246) );
  NAND3_X1 U216 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n5) );
  XOR2_X1 U217 ( .A(n20), .B(n23), .Z(n247) );
  NAND2_X1 U218 ( .A1(n20), .A2(n23), .ZN(n248) );
  NAND2_X1 U219 ( .A1(n20), .A2(n5), .ZN(n249) );
  NAND2_X1 U220 ( .A1(n238), .A2(n23), .ZN(n250) );
  NAND3_X1 U221 ( .A1(n249), .A2(n250), .A3(n248), .ZN(n4) );
  XOR2_X1 U222 ( .A(n46), .B(n49), .Z(n251) );
  XOR2_X1 U223 ( .A(n223), .B(n251), .Z(product[6]) );
  NAND2_X1 U224 ( .A1(n223), .A2(n46), .ZN(n252) );
  NAND2_X1 U225 ( .A1(n10), .A2(n49), .ZN(n253) );
  NAND2_X1 U226 ( .A1(n46), .A2(n49), .ZN(n254) );
  NAND3_X1 U227 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n9) );
  NAND3_X1 U228 ( .A1(n258), .A2(n257), .A3(n256), .ZN(n255) );
  BUF_X2 U229 ( .A(b[0]), .Z(n276) );
  NAND2_X1 U230 ( .A1(n17), .A2(n284), .ZN(n256) );
  NAND2_X1 U231 ( .A1(n17), .A2(n226), .ZN(n257) );
  NAND2_X1 U232 ( .A1(n284), .A2(n3), .ZN(n258) );
  NAND3_X1 U233 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n2) );
  XOR2_X1 U234 ( .A(n285), .B(n15), .Z(n259) );
  XOR2_X1 U235 ( .A(n259), .B(n2), .Z(product[14]) );
  NAND2_X1 U236 ( .A1(n285), .A2(n15), .ZN(n260) );
  NAND2_X1 U237 ( .A1(n255), .A2(n285), .ZN(n261) );
  NAND2_X1 U238 ( .A1(n255), .A2(n15), .ZN(n262) );
  XOR2_X1 U239 ( .A(n40), .B(n45), .Z(n263) );
  XOR2_X1 U240 ( .A(n209), .B(n263), .Z(product[7]) );
  NAND2_X1 U241 ( .A1(n236), .A2(n40), .ZN(n264) );
  NAND2_X1 U242 ( .A1(n9), .A2(n45), .ZN(n265) );
  NAND2_X1 U243 ( .A1(n40), .A2(n45), .ZN(n266) );
  NAND3_X1 U244 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n8) );
  XOR2_X1 U245 ( .A(n34), .B(n39), .Z(n267) );
  XOR2_X1 U246 ( .A(n267), .B(n237), .Z(product[8]) );
  NAND2_X1 U247 ( .A1(n34), .A2(n39), .ZN(n268) );
  NAND2_X1 U248 ( .A1(n34), .A2(n8), .ZN(n269) );
  NAND2_X1 U249 ( .A1(n39), .A2(n8), .ZN(n270) );
  NAND3_X1 U250 ( .A1(n269), .A2(n268), .A3(n270), .ZN(n7) );
  XOR2_X1 U251 ( .A(n28), .B(n33), .Z(n271) );
  XOR2_X1 U252 ( .A(n271), .B(n228), .Z(product[9]) );
  NAND2_X1 U253 ( .A1(n28), .A2(n33), .ZN(n272) );
  NAND2_X1 U254 ( .A1(n28), .A2(n227), .ZN(n273) );
  NAND2_X1 U255 ( .A1(n33), .A2(n7), .ZN(n274) );
  NAND3_X1 U256 ( .A1(n274), .A2(n273), .A3(n272), .ZN(n6) );
  XNOR2_X1 U257 ( .A(b[1]), .B(n281), .ZN(n275) );
  NAND2_X1 U258 ( .A1(a[4]), .A2(a[3]), .ZN(n278) );
  NAND2_X1 U259 ( .A1(n277), .A2(n292), .ZN(n279) );
  INV_X1 U260 ( .A(a[4]), .ZN(n277) );
  INV_X1 U261 ( .A(n15), .ZN(n284) );
  INV_X1 U262 ( .A(n31), .ZN(n290) );
  INV_X1 U263 ( .A(n21), .ZN(n287) );
  INV_X1 U264 ( .A(n320), .ZN(n288) );
  INV_X1 U265 ( .A(n331), .ZN(n285) );
  INV_X1 U266 ( .A(n300), .ZN(n293) );
  INV_X1 U267 ( .A(n309), .ZN(n291) );
  INV_X1 U268 ( .A(b[0]), .ZN(n283) );
  INV_X1 U269 ( .A(a[5]), .ZN(n289) );
  INV_X1 U270 ( .A(a[7]), .ZN(n286) );
  CLKBUF_X1 U271 ( .A(a[1]), .Z(n282) );
  XNOR2_X1 U272 ( .A(a[2]), .B(n282), .ZN(n301) );
  INV_X1 U273 ( .A(a[3]), .ZN(n292) );
  INV_X1 U274 ( .A(n281), .ZN(n294) );
  XOR2_X2 U275 ( .A(a[6]), .B(n289), .Z(n322) );
  INV_X2 U276 ( .A(a[0]), .ZN(n295) );
  NOR2_X1 U277 ( .A1(n295), .A2(n283), .ZN(product[0]) );
  OAI22_X1 U278 ( .A1(n296), .A2(n297), .B1(n298), .B2(n295), .ZN(n99) );
  OAI22_X1 U279 ( .A1(n298), .A2(n297), .B1(n299), .B2(n295), .ZN(n98) );
  XNOR2_X1 U280 ( .A(b[6]), .B(n281), .ZN(n298) );
  OAI22_X1 U281 ( .A1(n295), .A2(n299), .B1(n297), .B2(n299), .ZN(n300) );
  XNOR2_X1 U282 ( .A(b[7]), .B(n281), .ZN(n299) );
  NOR2_X1 U283 ( .A1(n280), .A2(n283), .ZN(n96) );
  OAI22_X1 U284 ( .A1(n302), .A2(n303), .B1(n280), .B2(n304), .ZN(n95) );
  XNOR2_X1 U285 ( .A(a[3]), .B(n276), .ZN(n302) );
  OAI22_X1 U286 ( .A1(n304), .A2(n303), .B1(n218), .B2(n305), .ZN(n94) );
  XNOR2_X1 U287 ( .A(b[1]), .B(a[3]), .ZN(n304) );
  OAI22_X1 U288 ( .A1(n305), .A2(n213), .B1(n218), .B2(n306), .ZN(n93) );
  XNOR2_X1 U289 ( .A(b[2]), .B(a[3]), .ZN(n305) );
  OAI22_X1 U290 ( .A1(n306), .A2(n213), .B1(n218), .B2(n307), .ZN(n92) );
  XNOR2_X1 U291 ( .A(b[3]), .B(a[3]), .ZN(n306) );
  OAI22_X1 U292 ( .A1(n307), .A2(n213), .B1(n218), .B2(n308), .ZN(n91) );
  XNOR2_X1 U293 ( .A(b[4]), .B(a[3]), .ZN(n307) );
  OAI22_X1 U294 ( .A1(n310), .A2(n218), .B1(n213), .B2(n310), .ZN(n309) );
  NOR2_X1 U295 ( .A1(n214), .A2(n283), .ZN(n88) );
  OAI22_X1 U296 ( .A1(n312), .A2(n313), .B1(n214), .B2(n314), .ZN(n87) );
  XNOR2_X1 U297 ( .A(a[5]), .B(n276), .ZN(n312) );
  OAI22_X1 U298 ( .A1(n314), .A2(n313), .B1(n214), .B2(n315), .ZN(n86) );
  XNOR2_X1 U299 ( .A(n211), .B(a[5]), .ZN(n314) );
  OAI22_X1 U300 ( .A1(n315), .A2(n313), .B1(n214), .B2(n316), .ZN(n85) );
  XNOR2_X1 U301 ( .A(b[2]), .B(a[5]), .ZN(n315) );
  OAI22_X1 U302 ( .A1(n316), .A2(n313), .B1(n214), .B2(n317), .ZN(n84) );
  XNOR2_X1 U303 ( .A(b[3]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U304 ( .A1(n317), .A2(n313), .B1(n214), .B2(n318), .ZN(n83) );
  XNOR2_X1 U305 ( .A(b[4]), .B(a[5]), .ZN(n317) );
  OAI22_X1 U306 ( .A1(n318), .A2(n313), .B1(n214), .B2(n319), .ZN(n82) );
  XNOR2_X1 U307 ( .A(b[5]), .B(a[5]), .ZN(n318) );
  OAI22_X1 U308 ( .A1(n321), .A2(n214), .B1(n313), .B2(n321), .ZN(n320) );
  NOR2_X1 U309 ( .A1(n322), .A2(n283), .ZN(n80) );
  OAI22_X1 U310 ( .A1(n323), .A2(n324), .B1(n322), .B2(n325), .ZN(n79) );
  XNOR2_X1 U311 ( .A(a[7]), .B(n276), .ZN(n323) );
  OAI22_X1 U312 ( .A1(n326), .A2(n324), .B1(n322), .B2(n327), .ZN(n77) );
  OAI22_X1 U313 ( .A1(n327), .A2(n324), .B1(n322), .B2(n328), .ZN(n76) );
  XNOR2_X1 U314 ( .A(b[3]), .B(a[7]), .ZN(n327) );
  OAI22_X1 U315 ( .A1(n328), .A2(n324), .B1(n322), .B2(n329), .ZN(n75) );
  XNOR2_X1 U316 ( .A(b[4]), .B(a[7]), .ZN(n328) );
  OAI22_X1 U317 ( .A1(n329), .A2(n324), .B1(n322), .B2(n330), .ZN(n74) );
  XNOR2_X1 U318 ( .A(b[5]), .B(a[7]), .ZN(n329) );
  OAI22_X1 U319 ( .A1(n332), .A2(n322), .B1(n324), .B2(n332), .ZN(n331) );
  OAI21_X1 U320 ( .B1(n276), .B2(n294), .A(n297), .ZN(n72) );
  OAI21_X1 U321 ( .B1(n292), .B2(n213), .A(n333), .ZN(n71) );
  OR3_X1 U322 ( .A1(n218), .A2(n276), .A3(n292), .ZN(n333) );
  OAI21_X1 U323 ( .B1(n289), .B2(n313), .A(n334), .ZN(n70) );
  OR3_X1 U324 ( .A1(n311), .A2(n276), .A3(n289), .ZN(n334) );
  OAI21_X1 U325 ( .B1(n286), .B2(n324), .A(n335), .ZN(n69) );
  OR3_X1 U326 ( .A1(n322), .A2(n276), .A3(n286), .ZN(n335) );
  XNOR2_X1 U327 ( .A(n336), .B(n337), .ZN(n38) );
  OR2_X1 U328 ( .A1(n336), .A2(n337), .ZN(n37) );
  OAI22_X1 U329 ( .A1(n308), .A2(n213), .B1(n218), .B2(n338), .ZN(n337) );
  XNOR2_X1 U330 ( .A(b[5]), .B(a[3]), .ZN(n308) );
  OAI22_X1 U331 ( .A1(n325), .A2(n324), .B1(n322), .B2(n326), .ZN(n336) );
  XNOR2_X1 U332 ( .A(b[2]), .B(a[7]), .ZN(n326) );
  XNOR2_X1 U333 ( .A(n211), .B(a[7]), .ZN(n325) );
  OAI22_X1 U334 ( .A1(n338), .A2(n213), .B1(n218), .B2(n310), .ZN(n31) );
  XNOR2_X1 U335 ( .A(b[7]), .B(a[3]), .ZN(n310) );
  XNOR2_X1 U336 ( .A(b[6]), .B(a[3]), .ZN(n338) );
  OAI22_X1 U337 ( .A1(n319), .A2(n313), .B1(n214), .B2(n321), .ZN(n21) );
  XNOR2_X1 U338 ( .A(b[7]), .B(a[5]), .ZN(n321) );
  XNOR2_X1 U339 ( .A(n289), .B(a[4]), .ZN(n340) );
  XNOR2_X1 U340 ( .A(b[6]), .B(a[5]), .ZN(n319) );
  OAI22_X1 U341 ( .A1(n330), .A2(n324), .B1(n322), .B2(n332), .ZN(n15) );
  XNOR2_X1 U342 ( .A(b[7]), .B(a[7]), .ZN(n332) );
  XNOR2_X1 U343 ( .A(n286), .B(a[6]), .ZN(n341) );
  XNOR2_X1 U344 ( .A(b[6]), .B(a[7]), .ZN(n330) );
  OAI22_X1 U345 ( .A1(n276), .A2(n297), .B1(n342), .B2(n295), .ZN(n104) );
  OAI22_X1 U346 ( .A1(n275), .A2(n297), .B1(n343), .B2(n295), .ZN(n103) );
  XNOR2_X1 U347 ( .A(b[1]), .B(n281), .ZN(n342) );
  OAI22_X1 U348 ( .A1(n343), .A2(n297), .B1(n344), .B2(n295), .ZN(n102) );
  XNOR2_X1 U349 ( .A(b[2]), .B(n282), .ZN(n343) );
  OAI22_X1 U350 ( .A1(n344), .A2(n297), .B1(n345), .B2(n295), .ZN(n101) );
  XNOR2_X1 U351 ( .A(b[3]), .B(n281), .ZN(n344) );
  OAI22_X1 U352 ( .A1(n345), .A2(n297), .B1(n296), .B2(n295), .ZN(n100) );
  XNOR2_X1 U353 ( .A(b[5]), .B(n282), .ZN(n296) );
  XNOR2_X1 U354 ( .A(b[4]), .B(n282), .ZN(n345) );
endmodule


module datapath_DW01_add_13 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n82;
  wire   [15:1] carry;

  FA_X1 U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n82), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(carry[3]), .Z(n1) );
  NAND3_X1 U2 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n2) );
  CLKBUF_X1 U3 ( .A(n66), .Z(n3) );
  NAND2_X1 U4 ( .A1(n47), .A2(B[11]), .ZN(n4) );
  CLKBUF_X1 U5 ( .A(B[11]), .Z(n5) );
  NAND2_X1 U6 ( .A1(n22), .A2(B[9]), .ZN(n6) );
  CLKBUF_X1 U7 ( .A(n22), .Z(n7) );
  CLKBUF_X1 U8 ( .A(n79), .Z(n8) );
  CLKBUF_X1 U9 ( .A(n44), .Z(n9) );
  CLKBUF_X1 U10 ( .A(n6), .Z(n10) );
  NAND2_X1 U11 ( .A1(B[11]), .A2(A[11]), .ZN(n11) );
  NAND2_X1 U12 ( .A1(n5), .A2(A[11]), .ZN(n12) );
  NAND3_X1 U13 ( .A1(n10), .A2(n31), .A3(n32), .ZN(n13) );
  NAND3_X1 U14 ( .A1(n19), .A2(n20), .A3(n21), .ZN(n14) );
  NAND2_X1 U15 ( .A1(n47), .A2(B[11]), .ZN(n15) );
  CLKBUF_X1 U16 ( .A(n33), .Z(n16) );
  CLKBUF_X1 U17 ( .A(B[5]), .Z(n17) );
  XOR2_X1 U18 ( .A(n1), .B(A[3]), .Z(n18) );
  XOR2_X1 U19 ( .A(B[3]), .B(n18), .Z(SUM[3]) );
  NAND2_X1 U20 ( .A1(B[3]), .A2(carry[3]), .ZN(n19) );
  NAND2_X1 U21 ( .A1(B[3]), .A2(A[3]), .ZN(n20) );
  NAND2_X1 U22 ( .A1(carry[3]), .A2(A[3]), .ZN(n21) );
  NAND3_X1 U23 ( .A1(n19), .A2(n20), .A3(n21), .ZN(carry[4]) );
  NAND3_X1 U24 ( .A1(n69), .A2(n70), .A3(n71), .ZN(n22) );
  NAND3_X1 U25 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n23) );
  XOR2_X1 U26 ( .A(B[4]), .B(A[4]), .Z(n24) );
  XOR2_X1 U27 ( .A(n14), .B(n24), .Z(SUM[4]) );
  NAND2_X1 U28 ( .A1(n14), .A2(B[4]), .ZN(n25) );
  NAND2_X1 U29 ( .A1(carry[4]), .A2(A[4]), .ZN(n26) );
  NAND2_X1 U30 ( .A1(B[4]), .A2(A[4]), .ZN(n27) );
  NAND3_X1 U31 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[5]) );
  NAND3_X1 U32 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n28) );
  XOR2_X1 U33 ( .A(B[9]), .B(A[9]), .Z(n29) );
  XOR2_X1 U34 ( .A(n7), .B(n29), .Z(SUM[9]) );
  NAND2_X1 U35 ( .A1(n22), .A2(B[9]), .ZN(n30) );
  NAND2_X1 U36 ( .A1(carry[9]), .A2(A[9]), .ZN(n31) );
  NAND2_X1 U37 ( .A1(B[9]), .A2(A[9]), .ZN(n32) );
  NAND3_X1 U38 ( .A1(n6), .A2(n31), .A3(n32), .ZN(carry[10]) );
  NAND3_X1 U39 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n33) );
  NAND3_X1 U40 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n34) );
  CLKBUF_X1 U41 ( .A(n4), .Z(n35) );
  XOR2_X1 U42 ( .A(B[6]), .B(A[6]), .Z(n36) );
  XOR2_X1 U43 ( .A(carry[6]), .B(n36), .Z(SUM[6]) );
  NAND2_X1 U44 ( .A1(n2), .A2(B[6]), .ZN(n37) );
  NAND2_X1 U45 ( .A1(n34), .A2(A[6]), .ZN(n38) );
  NAND2_X1 U46 ( .A1(B[6]), .A2(A[6]), .ZN(n39) );
  NAND3_X1 U47 ( .A1(n38), .A2(n37), .A3(n39), .ZN(carry[7]) );
  NAND3_X1 U48 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n40) );
  XOR2_X1 U49 ( .A(n17), .B(A[5]), .Z(n41) );
  XOR2_X1 U50 ( .A(n23), .B(n41), .Z(SUM[5]) );
  NAND2_X1 U51 ( .A1(B[5]), .A2(carry[5]), .ZN(n42) );
  NAND2_X1 U52 ( .A1(n23), .A2(A[5]), .ZN(n43) );
  NAND2_X1 U53 ( .A1(B[5]), .A2(A[5]), .ZN(n44) );
  NAND3_X1 U54 ( .A1(n42), .A2(n43), .A3(n9), .ZN(carry[6]) );
  CLKBUF_X1 U55 ( .A(n47), .Z(n45) );
  XNOR2_X1 U56 ( .A(n49), .B(n46), .ZN(SUM[14]) );
  XNOR2_X1 U57 ( .A(B[14]), .B(A[14]), .ZN(n46) );
  NAND3_X1 U58 ( .A1(n55), .A2(n54), .A3(n56), .ZN(n47) );
  NAND3_X1 U59 ( .A1(n78), .A2(n79), .A3(n80), .ZN(n48) );
  NAND3_X1 U60 ( .A1(n8), .A2(n78), .A3(n80), .ZN(n49) );
  NAND3_X1 U61 ( .A1(n15), .A2(n66), .A3(n67), .ZN(n50) );
  NAND3_X1 U62 ( .A1(n35), .A2(n3), .A3(n12), .ZN(n51) );
  NAND3_X1 U63 ( .A1(n76), .A2(n74), .A3(n75), .ZN(n52) );
  XOR2_X1 U64 ( .A(B[10]), .B(A[10]), .Z(n53) );
  XOR2_X1 U65 ( .A(n13), .B(n53), .Z(SUM[10]) );
  NAND2_X1 U66 ( .A1(n28), .A2(B[10]), .ZN(n54) );
  NAND2_X1 U67 ( .A1(carry[10]), .A2(A[10]), .ZN(n55) );
  NAND2_X1 U68 ( .A1(B[10]), .A2(A[10]), .ZN(n56) );
  NAND3_X1 U69 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[11]) );
  XNOR2_X1 U70 ( .A(carry[15]), .B(n57), .ZN(SUM[15]) );
  XNOR2_X1 U71 ( .A(B[15]), .B(A[15]), .ZN(n57) );
  NAND2_X1 U72 ( .A1(B[14]), .A2(carry[14]), .ZN(n58) );
  NAND2_X1 U73 ( .A1(n48), .A2(A[14]), .ZN(n59) );
  NAND2_X1 U74 ( .A1(B[14]), .A2(A[14]), .ZN(n60) );
  NAND3_X1 U75 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[15]) );
  XOR2_X1 U76 ( .A(B[7]), .B(A[7]), .Z(n61) );
  XOR2_X1 U77 ( .A(n16), .B(n61), .Z(SUM[7]) );
  NAND2_X1 U78 ( .A1(n33), .A2(B[7]), .ZN(n62) );
  NAND2_X1 U79 ( .A1(carry[7]), .A2(A[7]), .ZN(n63) );
  NAND2_X1 U80 ( .A1(B[7]), .A2(A[7]), .ZN(n64) );
  NAND3_X1 U81 ( .A1(n62), .A2(n63), .A3(n64), .ZN(carry[8]) );
  XOR2_X1 U82 ( .A(n5), .B(A[11]), .Z(n65) );
  XOR2_X1 U83 ( .A(n45), .B(n65), .Z(SUM[11]) );
  NAND2_X1 U84 ( .A1(carry[11]), .A2(A[11]), .ZN(n66) );
  NAND2_X1 U85 ( .A1(B[11]), .A2(A[11]), .ZN(n67) );
  NAND3_X1 U86 ( .A1(n4), .A2(n66), .A3(n11), .ZN(carry[12]) );
  XOR2_X1 U87 ( .A(B[8]), .B(A[8]), .Z(n68) );
  XOR2_X1 U88 ( .A(carry[8]), .B(n68), .Z(SUM[8]) );
  NAND2_X1 U89 ( .A1(n40), .A2(B[8]), .ZN(n69) );
  NAND2_X1 U90 ( .A1(n40), .A2(A[8]), .ZN(n70) );
  NAND2_X1 U91 ( .A1(B[8]), .A2(A[8]), .ZN(n71) );
  NAND3_X1 U92 ( .A1(n69), .A2(n70), .A3(n71), .ZN(carry[9]) );
  CLKBUF_X1 U93 ( .A(n52), .Z(n72) );
  XOR2_X1 U94 ( .A(A[12]), .B(B[12]), .Z(n73) );
  XOR2_X1 U95 ( .A(n73), .B(n51), .Z(SUM[12]) );
  NAND2_X1 U96 ( .A1(A[12]), .A2(B[12]), .ZN(n74) );
  NAND2_X1 U97 ( .A1(A[12]), .A2(n50), .ZN(n75) );
  NAND2_X1 U98 ( .A1(B[12]), .A2(carry[12]), .ZN(n76) );
  NAND3_X1 U99 ( .A1(n74), .A2(n75), .A3(n76), .ZN(carry[13]) );
  XOR2_X1 U100 ( .A(B[13]), .B(A[13]), .Z(n77) );
  XOR2_X1 U101 ( .A(n77), .B(n72), .Z(SUM[13]) );
  NAND2_X1 U102 ( .A1(A[13]), .A2(B[13]), .ZN(n78) );
  NAND2_X1 U103 ( .A1(n52), .A2(A[13]), .ZN(n79) );
  NAND2_X1 U104 ( .A1(B[13]), .A2(carry[13]), .ZN(n80) );
  NAND3_X1 U105 ( .A1(n79), .A2(n78), .A3(n80), .ZN(carry[14]) );
  XOR2_X1 U106 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U107 ( .A1(B[0]), .A2(A[0]), .ZN(n82) );
endmodule


module datapath_DW_mult_tc_12 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n210, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351;

  FA_X1 U12 ( .A(n54), .B(n209), .CI(n12), .CO(n11), .S(product[4]) );
  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n294), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n293), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n297), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n296), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n299), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  BUF_X2 U157 ( .A(a[1]), .Z(n208) );
  INV_X1 U158 ( .A(n281), .ZN(n288) );
  NAND2_X1 U159 ( .A1(n206), .A2(n301), .ZN(n303) );
  NAND3_X1 U160 ( .A1(n283), .A2(n284), .A3(n285), .ZN(n49) );
  NAND2_X1 U161 ( .A1(n317), .A2(n346), .ZN(n319) );
  INV_X1 U162 ( .A(n15), .ZN(n290) );
  CLKBUF_X1 U163 ( .A(a[1]), .Z(n206) );
  BUF_X1 U164 ( .A(a[1]), .Z(n207) );
  AND2_X1 U165 ( .A1(n95), .A2(n102), .ZN(n209) );
  XNOR2_X1 U166 ( .A(n291), .B(n15), .ZN(n210) );
  AND3_X1 U167 ( .A1(n258), .A2(n259), .A3(n260), .ZN(product[15]) );
  XOR2_X1 U168 ( .A(n19), .B(n18), .Z(n212) );
  XOR2_X1 U169 ( .A(n4), .B(n212), .Z(product[12]) );
  NAND2_X1 U170 ( .A1(n4), .A2(n19), .ZN(n213) );
  NAND2_X1 U171 ( .A1(n4), .A2(n18), .ZN(n214) );
  NAND2_X1 U172 ( .A1(n19), .A2(n18), .ZN(n215) );
  NAND3_X1 U173 ( .A1(n213), .A2(n214), .A3(n215), .ZN(n3) );
  XOR2_X1 U174 ( .A(n216), .B(n217), .Z(product[6]) );
  AND3_X1 U175 ( .A1(n265), .A2(n266), .A3(n267), .ZN(n216) );
  XNOR2_X1 U176 ( .A(n46), .B(n49), .ZN(n217) );
  CLKBUF_X1 U177 ( .A(b[1]), .Z(n218) );
  XOR2_X1 U178 ( .A(a[3]), .B(a[2]), .Z(n219) );
  XOR2_X1 U179 ( .A(a[3]), .B(a[2]), .Z(n345) );
  NAND2_X1 U180 ( .A1(n6), .A2(n24), .ZN(n220) );
  BUF_X2 U181 ( .A(n317), .Z(n221) );
  XNOR2_X1 U182 ( .A(a[4]), .B(a[3]), .ZN(n317) );
  NAND2_X1 U183 ( .A1(n10), .A2(n49), .ZN(n222) );
  BUF_X1 U184 ( .A(n289), .Z(n223) );
  BUF_X2 U185 ( .A(n328), .Z(n224) );
  XOR2_X1 U186 ( .A(a[6]), .B(n295), .Z(n328) );
  AND2_X1 U187 ( .A1(n104), .A2(n72), .ZN(n225) );
  NAND3_X1 U188 ( .A1(n256), .A2(n255), .A3(n257), .ZN(n226) );
  NAND3_X1 U189 ( .A1(n278), .A2(n279), .A3(n280), .ZN(n227) );
  XNOR2_X1 U190 ( .A(n249), .B(n228), .ZN(product[5]) );
  XNOR2_X1 U191 ( .A(n50), .B(n53), .ZN(n228) );
  NAND3_X1 U192 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n229) );
  NAND3_X1 U193 ( .A1(n246), .A2(n220), .A3(n248), .ZN(n230) );
  XNOR2_X1 U194 ( .A(n2), .B(n210), .ZN(product[14]) );
  NAND3_X1 U195 ( .A1(n279), .A2(n278), .A3(n280), .ZN(n231) );
  NAND3_X1 U196 ( .A1(n280), .A2(n279), .A3(n278), .ZN(n232) );
  OR2_X1 U197 ( .A1(n349), .A2(n303), .ZN(n233) );
  OR2_X1 U198 ( .A1(n350), .A2(n301), .ZN(n234) );
  NAND2_X1 U199 ( .A1(n233), .A2(n234), .ZN(n102) );
  XNOR2_X1 U200 ( .A(n225), .B(n235), .ZN(product[2]) );
  XNOR2_X1 U201 ( .A(n103), .B(n96), .ZN(n235) );
  XOR2_X1 U202 ( .A(n23), .B(n20), .Z(n236) );
  XOR2_X1 U203 ( .A(n230), .B(n236), .Z(product[11]) );
  NAND2_X1 U204 ( .A1(n229), .A2(n23), .ZN(n237) );
  NAND2_X1 U205 ( .A1(n5), .A2(n20), .ZN(n238) );
  NAND2_X1 U206 ( .A1(n23), .A2(n20), .ZN(n239) );
  NAND3_X1 U207 ( .A1(n238), .A2(n237), .A3(n239), .ZN(n4) );
  XOR2_X1 U208 ( .A(n17), .B(n290), .Z(n240) );
  XOR2_X1 U209 ( .A(n3), .B(n240), .Z(product[13]) );
  NAND2_X1 U210 ( .A1(n3), .A2(n17), .ZN(n241) );
  NAND2_X1 U211 ( .A1(n3), .A2(n290), .ZN(n242) );
  NAND2_X1 U212 ( .A1(n17), .A2(n290), .ZN(n243) );
  NAND3_X1 U213 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n2) );
  NAND3_X1 U214 ( .A1(n255), .A2(n257), .A3(n256), .ZN(n244) );
  XOR2_X1 U215 ( .A(n27), .B(n24), .Z(n245) );
  XOR2_X1 U216 ( .A(n226), .B(n245), .Z(product[10]) );
  NAND2_X1 U217 ( .A1(n244), .A2(n27), .ZN(n246) );
  NAND2_X1 U218 ( .A1(n6), .A2(n24), .ZN(n247) );
  NAND2_X1 U219 ( .A1(n27), .A2(n24), .ZN(n248) );
  NAND3_X1 U220 ( .A1(n220), .A2(n246), .A3(n248), .ZN(n5) );
  CLKBUF_X1 U221 ( .A(n11), .Z(n249) );
  NAND3_X1 U222 ( .A1(n269), .A2(n222), .A3(n271), .ZN(n250) );
  NAND3_X1 U223 ( .A1(n266), .A2(n267), .A3(n265), .ZN(n251) );
  XOR2_X1 U224 ( .A(a[3]), .B(n289), .Z(n308) );
  XNOR2_X1 U225 ( .A(a[2]), .B(n208), .ZN(n252) );
  XNOR2_X1 U226 ( .A(a[2]), .B(n206), .ZN(n253) );
  XNOR2_X1 U227 ( .A(a[2]), .B(n207), .ZN(n307) );
  XOR2_X1 U228 ( .A(n33), .B(n28), .Z(n254) );
  XOR2_X1 U229 ( .A(n227), .B(n254), .Z(product[9]) );
  NAND2_X1 U230 ( .A1(n232), .A2(n33), .ZN(n255) );
  NAND2_X1 U231 ( .A1(n231), .A2(n28), .ZN(n256) );
  NAND2_X1 U232 ( .A1(n33), .A2(n28), .ZN(n257) );
  NAND3_X1 U233 ( .A1(n256), .A2(n255), .A3(n257), .ZN(n6) );
  NAND2_X1 U234 ( .A1(n2), .A2(n291), .ZN(n258) );
  NAND2_X1 U235 ( .A1(n2), .A2(n15), .ZN(n259) );
  NAND2_X1 U236 ( .A1(n291), .A2(n15), .ZN(n260) );
  XOR2_X1 U237 ( .A(n95), .B(n102), .Z(n56) );
  NAND2_X1 U238 ( .A1(n225), .A2(n103), .ZN(n261) );
  NAND2_X1 U239 ( .A1(n14), .A2(n96), .ZN(n262) );
  NAND2_X1 U240 ( .A1(n103), .A2(n96), .ZN(n263) );
  NAND3_X1 U241 ( .A1(n262), .A2(n261), .A3(n263), .ZN(n13) );
  BUF_X1 U242 ( .A(n275), .Z(n264) );
  NAND2_X1 U243 ( .A1(n11), .A2(n50), .ZN(n265) );
  NAND2_X1 U244 ( .A1(n11), .A2(n53), .ZN(n266) );
  NAND2_X1 U245 ( .A1(n50), .A2(n53), .ZN(n267) );
  NAND3_X1 U246 ( .A1(n265), .A2(n266), .A3(n267), .ZN(n10) );
  NAND3_X1 U247 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n268) );
  NAND2_X1 U248 ( .A1(n251), .A2(n46), .ZN(n269) );
  NAND2_X1 U249 ( .A1(n10), .A2(n49), .ZN(n270) );
  NAND2_X1 U250 ( .A1(n46), .A2(n49), .ZN(n271) );
  NAND3_X1 U251 ( .A1(n222), .A2(n269), .A3(n271), .ZN(n9) );
  NAND3_X1 U252 ( .A1(n274), .A2(n264), .A3(n276), .ZN(n272) );
  XOR2_X1 U253 ( .A(n40), .B(n45), .Z(n273) );
  XOR2_X1 U254 ( .A(n273), .B(n250), .Z(product[7]) );
  NAND2_X1 U255 ( .A1(n40), .A2(n45), .ZN(n274) );
  NAND2_X1 U256 ( .A1(n9), .A2(n40), .ZN(n275) );
  NAND2_X1 U257 ( .A1(n45), .A2(n268), .ZN(n276) );
  NAND3_X1 U258 ( .A1(n276), .A2(n275), .A3(n274), .ZN(n8) );
  XOR2_X1 U259 ( .A(n34), .B(n39), .Z(n277) );
  XOR2_X1 U260 ( .A(n277), .B(n272), .Z(product[8]) );
  NAND2_X1 U261 ( .A1(n34), .A2(n39), .ZN(n278) );
  NAND2_X1 U262 ( .A1(n8), .A2(n34), .ZN(n279) );
  NAND2_X1 U263 ( .A1(n8), .A2(n39), .ZN(n280) );
  INV_X1 U264 ( .A(b[0]), .ZN(n281) );
  XNOR2_X1 U265 ( .A(n52), .B(n282), .ZN(n50) );
  XNOR2_X1 U266 ( .A(n93), .B(n100), .ZN(n282) );
  INV_X1 U267 ( .A(n31), .ZN(n296) );
  INV_X1 U268 ( .A(n21), .ZN(n293) );
  INV_X1 U269 ( .A(n326), .ZN(n294) );
  INV_X1 U270 ( .A(n337), .ZN(n291) );
  INV_X1 U271 ( .A(n306), .ZN(n299) );
  INV_X1 U272 ( .A(n315), .ZN(n297) );
  INV_X1 U273 ( .A(b[0]), .ZN(n289) );
  INV_X1 U274 ( .A(a[5]), .ZN(n295) );
  INV_X1 U275 ( .A(a[7]), .ZN(n292) );
  NAND2_X1 U276 ( .A1(n52), .A2(n93), .ZN(n283) );
  NAND2_X1 U277 ( .A1(n52), .A2(n100), .ZN(n284) );
  NAND2_X1 U278 ( .A1(n93), .A2(n100), .ZN(n285) );
  INV_X1 U279 ( .A(a[3]), .ZN(n298) );
  NAND2_X1 U280 ( .A1(n307), .A2(n219), .ZN(n286) );
  NAND2_X1 U281 ( .A1(n252), .A2(n345), .ZN(n287) );
  NAND2_X1 U282 ( .A1(n307), .A2(n345), .ZN(n309) );
  INV_X1 U283 ( .A(n207), .ZN(n300) );
  INV_X2 U284 ( .A(a[0]), .ZN(n301) );
  NOR2_X1 U285 ( .A1(n301), .A2(n223), .ZN(product[0]) );
  OAI22_X1 U286 ( .A1(n302), .A2(n303), .B1(n304), .B2(n301), .ZN(n99) );
  OAI22_X1 U287 ( .A1(n304), .A2(n303), .B1(n305), .B2(n301), .ZN(n98) );
  XNOR2_X1 U288 ( .A(b[6]), .B(n207), .ZN(n304) );
  OAI22_X1 U289 ( .A1(n301), .A2(n305), .B1(n303), .B2(n305), .ZN(n306) );
  XNOR2_X1 U290 ( .A(b[7]), .B(n207), .ZN(n305) );
  NOR2_X1 U291 ( .A1(n252), .A2(n223), .ZN(n96) );
  OAI22_X1 U292 ( .A1(n309), .A2(n308), .B1(n253), .B2(n310), .ZN(n95) );
  OAI22_X1 U293 ( .A1(n310), .A2(n286), .B1(n253), .B2(n311), .ZN(n94) );
  XNOR2_X1 U294 ( .A(b[1]), .B(a[3]), .ZN(n310) );
  OAI22_X1 U295 ( .A1(n311), .A2(n287), .B1(n252), .B2(n312), .ZN(n93) );
  XNOR2_X1 U296 ( .A(b[2]), .B(a[3]), .ZN(n311) );
  OAI22_X1 U297 ( .A1(n312), .A2(n286), .B1(n253), .B2(n313), .ZN(n92) );
  XNOR2_X1 U298 ( .A(b[3]), .B(a[3]), .ZN(n312) );
  OAI22_X1 U299 ( .A1(n313), .A2(n286), .B1(n253), .B2(n314), .ZN(n91) );
  XNOR2_X1 U300 ( .A(b[4]), .B(a[3]), .ZN(n313) );
  OAI22_X1 U301 ( .A1(n316), .A2(n252), .B1(n286), .B2(n316), .ZN(n315) );
  NOR2_X1 U302 ( .A1(n221), .A2(n223), .ZN(n88) );
  OAI22_X1 U303 ( .A1(n318), .A2(n319), .B1(n221), .B2(n320), .ZN(n87) );
  XNOR2_X1 U304 ( .A(a[5]), .B(n288), .ZN(n318) );
  OAI22_X1 U305 ( .A1(n320), .A2(n319), .B1(n221), .B2(n321), .ZN(n86) );
  XNOR2_X1 U306 ( .A(n218), .B(a[5]), .ZN(n320) );
  OAI22_X1 U307 ( .A1(n321), .A2(n319), .B1(n221), .B2(n322), .ZN(n85) );
  XNOR2_X1 U308 ( .A(b[2]), .B(a[5]), .ZN(n321) );
  OAI22_X1 U309 ( .A1(n322), .A2(n319), .B1(n221), .B2(n323), .ZN(n84) );
  XNOR2_X1 U310 ( .A(b[3]), .B(a[5]), .ZN(n322) );
  OAI22_X1 U311 ( .A1(n323), .A2(n319), .B1(n221), .B2(n324), .ZN(n83) );
  XNOR2_X1 U312 ( .A(b[4]), .B(a[5]), .ZN(n323) );
  OAI22_X1 U313 ( .A1(n324), .A2(n319), .B1(n221), .B2(n325), .ZN(n82) );
  XNOR2_X1 U314 ( .A(b[5]), .B(a[5]), .ZN(n324) );
  OAI22_X1 U315 ( .A1(n327), .A2(n221), .B1(n319), .B2(n327), .ZN(n326) );
  NOR2_X1 U316 ( .A1(n328), .A2(n223), .ZN(n80) );
  OAI22_X1 U317 ( .A1(n329), .A2(n330), .B1(n224), .B2(n331), .ZN(n79) );
  XNOR2_X1 U318 ( .A(a[7]), .B(n288), .ZN(n329) );
  OAI22_X1 U319 ( .A1(n332), .A2(n330), .B1(n224), .B2(n333), .ZN(n77) );
  OAI22_X1 U320 ( .A1(n333), .A2(n330), .B1(n224), .B2(n334), .ZN(n76) );
  XNOR2_X1 U321 ( .A(b[3]), .B(a[7]), .ZN(n333) );
  OAI22_X1 U322 ( .A1(n334), .A2(n330), .B1(n224), .B2(n335), .ZN(n75) );
  XNOR2_X1 U323 ( .A(b[4]), .B(a[7]), .ZN(n334) );
  OAI22_X1 U324 ( .A1(n335), .A2(n330), .B1(n224), .B2(n336), .ZN(n74) );
  XNOR2_X1 U325 ( .A(b[5]), .B(a[7]), .ZN(n335) );
  OAI22_X1 U326 ( .A1(n338), .A2(n224), .B1(n330), .B2(n338), .ZN(n337) );
  OAI21_X1 U327 ( .B1(n288), .B2(n300), .A(n303), .ZN(n72) );
  OAI21_X1 U328 ( .B1(n298), .B2(n287), .A(n339), .ZN(n71) );
  OR3_X1 U329 ( .A1(n253), .A2(n288), .A3(n298), .ZN(n339) );
  OAI21_X1 U330 ( .B1(n295), .B2(n319), .A(n340), .ZN(n70) );
  OR3_X1 U331 ( .A1(n221), .A2(n288), .A3(n295), .ZN(n340) );
  OAI21_X1 U332 ( .B1(n292), .B2(n330), .A(n341), .ZN(n69) );
  OR3_X1 U333 ( .A1(n328), .A2(n288), .A3(n292), .ZN(n341) );
  XNOR2_X1 U334 ( .A(n342), .B(n343), .ZN(n38) );
  OR2_X1 U335 ( .A1(n342), .A2(n343), .ZN(n37) );
  OAI22_X1 U336 ( .A1(n314), .A2(n287), .B1(n252), .B2(n344), .ZN(n343) );
  XNOR2_X1 U337 ( .A(b[5]), .B(a[3]), .ZN(n314) );
  OAI22_X1 U338 ( .A1(n331), .A2(n330), .B1(n224), .B2(n332), .ZN(n342) );
  XNOR2_X1 U339 ( .A(b[2]), .B(a[7]), .ZN(n332) );
  XNOR2_X1 U340 ( .A(n218), .B(a[7]), .ZN(n331) );
  OAI22_X1 U341 ( .A1(n344), .A2(n287), .B1(n253), .B2(n316), .ZN(n31) );
  XNOR2_X1 U342 ( .A(b[7]), .B(a[3]), .ZN(n316) );
  XNOR2_X1 U343 ( .A(b[6]), .B(a[3]), .ZN(n344) );
  OAI22_X1 U344 ( .A1(n325), .A2(n319), .B1(n221), .B2(n327), .ZN(n21) );
  XNOR2_X1 U345 ( .A(b[7]), .B(a[5]), .ZN(n327) );
  XNOR2_X1 U346 ( .A(n295), .B(a[4]), .ZN(n346) );
  XNOR2_X1 U347 ( .A(b[6]), .B(a[5]), .ZN(n325) );
  OAI22_X1 U348 ( .A1(n336), .A2(n330), .B1(n224), .B2(n338), .ZN(n15) );
  XNOR2_X1 U349 ( .A(b[7]), .B(a[7]), .ZN(n338) );
  NAND2_X1 U350 ( .A1(n328), .A2(n347), .ZN(n330) );
  XNOR2_X1 U351 ( .A(n292), .B(a[6]), .ZN(n347) );
  XNOR2_X1 U352 ( .A(b[6]), .B(a[7]), .ZN(n336) );
  OAI22_X1 U353 ( .A1(n288), .A2(n303), .B1(n348), .B2(n301), .ZN(n104) );
  OAI22_X1 U354 ( .A1(n348), .A2(n303), .B1(n301), .B2(n349), .ZN(n103) );
  XNOR2_X1 U355 ( .A(b[1]), .B(n208), .ZN(n348) );
  XNOR2_X1 U356 ( .A(b[2]), .B(n208), .ZN(n349) );
  OAI22_X1 U357 ( .A1(n350), .A2(n303), .B1(n351), .B2(n301), .ZN(n101) );
  XNOR2_X1 U358 ( .A(b[3]), .B(n207), .ZN(n350) );
  OAI22_X1 U359 ( .A1(n351), .A2(n303), .B1(n302), .B2(n301), .ZN(n100) );
  XNOR2_X1 U360 ( .A(b[5]), .B(n208), .ZN(n302) );
  XNOR2_X1 U361 ( .A(b[4]), .B(n208), .ZN(n351) );
endmodule


module datapath_DW01_add_12 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n82;
  wire   [15:1] carry;

  CLKBUF_X1 U1 ( .A(B[5]), .Z(n1) );
  CLKBUF_X1 U2 ( .A(B[8]), .Z(n2) );
  XNOR2_X1 U3 ( .A(B[14]), .B(A[14]), .ZN(n3) );
  XNOR2_X1 U4 ( .A(n3), .B(n8), .ZN(SUM[14]) );
  CLKBUF_X1 U5 ( .A(n35), .Z(n4) );
  CLKBUF_X1 U6 ( .A(n36), .Z(n5) );
  CLKBUF_X1 U7 ( .A(n33), .Z(n6) );
  CLKBUF_X1 U8 ( .A(n16), .Z(n7) );
  NAND3_X1 U9 ( .A1(n80), .A2(n79), .A3(n78), .ZN(n8) );
  NAND2_X1 U10 ( .A1(n8), .A2(B[14]), .ZN(n9) );
  NAND2_X1 U11 ( .A1(carry[14]), .A2(A[14]), .ZN(n10) );
  NAND2_X1 U12 ( .A1(B[14]), .A2(A[14]), .ZN(n11) );
  NAND3_X1 U13 ( .A1(n9), .A2(n10), .A3(n11), .ZN(carry[15]) );
  XOR2_X1 U14 ( .A(n82), .B(A[1]), .Z(n12) );
  XOR2_X1 U15 ( .A(B[1]), .B(n12), .Z(SUM[1]) );
  NAND2_X1 U16 ( .A1(B[1]), .A2(n82), .ZN(n13) );
  NAND2_X1 U17 ( .A1(B[1]), .A2(A[1]), .ZN(n14) );
  NAND2_X1 U18 ( .A1(n82), .A2(A[1]), .ZN(n15) );
  NAND3_X1 U19 ( .A1(n13), .A2(n14), .A3(n15), .ZN(carry[2]) );
  NAND2_X1 U20 ( .A1(n35), .A2(B[10]), .ZN(n16) );
  NAND3_X1 U21 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n17) );
  NAND3_X1 U22 ( .A1(n74), .A2(n75), .A3(n76), .ZN(n18) );
  NAND3_X1 U23 ( .A1(n66), .A2(n67), .A3(n68), .ZN(n19) );
  NAND3_X1 U24 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n20) );
  NAND3_X1 U25 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n21) );
  NAND3_X1 U26 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n22) );
  XOR2_X1 U27 ( .A(n22), .B(A[4]), .Z(n23) );
  XOR2_X1 U28 ( .A(B[4]), .B(n23), .Z(SUM[4]) );
  NAND2_X1 U29 ( .A1(B[4]), .A2(n21), .ZN(n24) );
  NAND2_X1 U30 ( .A1(B[4]), .A2(A[4]), .ZN(n25) );
  NAND2_X1 U31 ( .A1(carry[4]), .A2(A[4]), .ZN(n26) );
  NAND3_X1 U32 ( .A1(n24), .A2(n25), .A3(n26), .ZN(carry[5]) );
  NAND3_X1 U33 ( .A1(n16), .A2(n47), .A3(n48), .ZN(n27) );
  NAND3_X1 U34 ( .A1(n7), .A2(n47), .A3(n48), .ZN(n28) );
  XOR2_X1 U35 ( .A(B[11]), .B(A[11]), .Z(n29) );
  XOR2_X1 U36 ( .A(n28), .B(n29), .Z(SUM[11]) );
  NAND2_X1 U37 ( .A1(n27), .A2(B[11]), .ZN(n30) );
  NAND2_X1 U38 ( .A1(carry[11]), .A2(A[11]), .ZN(n31) );
  NAND2_X1 U39 ( .A1(B[11]), .A2(A[11]), .ZN(n32) );
  NAND3_X1 U40 ( .A1(n30), .A2(n31), .A3(n32), .ZN(carry[12]) );
  NAND3_X1 U41 ( .A1(n39), .A2(n41), .A3(n40), .ZN(n33) );
  NAND3_X1 U42 ( .A1(n50), .A2(n51), .A3(n52), .ZN(n34) );
  NAND3_X1 U43 ( .A1(n70), .A2(n71), .A3(n72), .ZN(n35) );
  NAND3_X1 U44 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n36) );
  NAND3_X1 U45 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n37) );
  XOR2_X1 U46 ( .A(n2), .B(A[8]), .Z(n38) );
  XOR2_X1 U47 ( .A(carry[8]), .B(n38), .Z(SUM[8]) );
  NAND2_X1 U48 ( .A1(B[8]), .A2(n19), .ZN(n39) );
  NAND2_X1 U49 ( .A1(n19), .A2(A[8]), .ZN(n40) );
  NAND2_X1 U50 ( .A1(B[8]), .A2(A[8]), .ZN(n41) );
  NAND3_X1 U51 ( .A1(n41), .A2(n40), .A3(n39), .ZN(carry[9]) );
  XNOR2_X1 U52 ( .A(carry[15]), .B(n42), .ZN(SUM[15]) );
  XNOR2_X1 U53 ( .A(B[15]), .B(A[15]), .ZN(n42) );
  NAND3_X1 U54 ( .A1(n74), .A2(n75), .A3(n76), .ZN(n43) );
  NAND3_X1 U55 ( .A1(n75), .A2(n74), .A3(n76), .ZN(n44) );
  XOR2_X1 U56 ( .A(B[10]), .B(A[10]), .Z(n45) );
  XOR2_X1 U57 ( .A(n4), .B(n45), .Z(SUM[10]) );
  NAND2_X1 U58 ( .A1(n35), .A2(B[10]), .ZN(n46) );
  NAND2_X1 U59 ( .A1(carry[10]), .A2(A[10]), .ZN(n47) );
  NAND2_X1 U60 ( .A1(B[10]), .A2(A[10]), .ZN(n48) );
  NAND3_X1 U61 ( .A1(n46), .A2(n47), .A3(n48), .ZN(carry[11]) );
  XOR2_X1 U62 ( .A(n1), .B(A[5]), .Z(n49) );
  XOR2_X1 U63 ( .A(carry[5]), .B(n49), .Z(SUM[5]) );
  NAND2_X1 U64 ( .A1(n20), .A2(B[5]), .ZN(n50) );
  NAND2_X1 U65 ( .A1(n20), .A2(A[5]), .ZN(n51) );
  NAND2_X1 U66 ( .A1(B[5]), .A2(A[5]), .ZN(n52) );
  NAND3_X1 U67 ( .A1(n51), .A2(n50), .A3(n52), .ZN(carry[6]) );
  XOR2_X1 U68 ( .A(B[2]), .B(A[2]), .Z(n53) );
  XOR2_X1 U69 ( .A(carry[2]), .B(n53), .Z(SUM[2]) );
  NAND2_X1 U70 ( .A1(carry[2]), .A2(B[2]), .ZN(n54) );
  NAND2_X1 U71 ( .A1(carry[2]), .A2(A[2]), .ZN(n55) );
  NAND2_X1 U72 ( .A1(B[2]), .A2(A[2]), .ZN(n56) );
  NAND3_X1 U73 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[3]) );
  NAND2_X1 U74 ( .A1(B[12]), .A2(A[12]), .ZN(n74) );
  XOR2_X1 U75 ( .A(B[3]), .B(A[3]), .Z(n57) );
  XOR2_X1 U76 ( .A(n37), .B(n57), .Z(SUM[3]) );
  NAND2_X1 U77 ( .A1(n37), .A2(B[3]), .ZN(n58) );
  NAND2_X1 U78 ( .A1(carry[3]), .A2(A[3]), .ZN(n59) );
  NAND2_X1 U79 ( .A1(B[3]), .A2(A[3]), .ZN(n60) );
  NAND3_X1 U80 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[4]) );
  XOR2_X1 U81 ( .A(B[6]), .B(A[6]), .Z(n61) );
  XOR2_X1 U82 ( .A(n34), .B(n61), .Z(SUM[6]) );
  NAND2_X1 U83 ( .A1(n34), .A2(B[6]), .ZN(n62) );
  NAND2_X1 U84 ( .A1(carry[6]), .A2(A[6]), .ZN(n63) );
  NAND2_X1 U85 ( .A1(B[6]), .A2(A[6]), .ZN(n64) );
  NAND3_X1 U86 ( .A1(n62), .A2(n63), .A3(n64), .ZN(carry[7]) );
  XOR2_X1 U87 ( .A(B[7]), .B(A[7]), .Z(n65) );
  XOR2_X1 U88 ( .A(n5), .B(n65), .Z(SUM[7]) );
  NAND2_X1 U89 ( .A1(n36), .A2(B[7]), .ZN(n66) );
  NAND2_X1 U90 ( .A1(carry[7]), .A2(A[7]), .ZN(n67) );
  NAND2_X1 U91 ( .A1(B[7]), .A2(A[7]), .ZN(n68) );
  NAND3_X1 U92 ( .A1(n66), .A2(n67), .A3(n68), .ZN(carry[8]) );
  XOR2_X1 U93 ( .A(B[9]), .B(A[9]), .Z(n69) );
  XOR2_X1 U94 ( .A(n6), .B(n69), .Z(SUM[9]) );
  NAND2_X1 U95 ( .A1(n33), .A2(B[9]), .ZN(n70) );
  NAND2_X1 U96 ( .A1(carry[9]), .A2(A[9]), .ZN(n71) );
  NAND2_X1 U97 ( .A1(B[9]), .A2(A[9]), .ZN(n72) );
  NAND3_X1 U98 ( .A1(n70), .A2(n71), .A3(n72), .ZN(carry[10]) );
  XOR2_X1 U99 ( .A(A[12]), .B(B[12]), .Z(n73) );
  XOR2_X1 U100 ( .A(n73), .B(n17), .Z(SUM[12]) );
  NAND2_X1 U101 ( .A1(A[12]), .A2(n17), .ZN(n75) );
  NAND2_X1 U102 ( .A1(B[12]), .A2(carry[12]), .ZN(n76) );
  XOR2_X1 U103 ( .A(A[13]), .B(B[13]), .Z(n77) );
  XOR2_X1 U104 ( .A(n77), .B(n18), .Z(SUM[13]) );
  NAND2_X1 U105 ( .A1(A[13]), .A2(B[13]), .ZN(n78) );
  NAND2_X1 U106 ( .A1(n44), .A2(A[13]), .ZN(n79) );
  NAND2_X1 U107 ( .A1(n43), .A2(B[13]), .ZN(n80) );
  NAND3_X1 U108 ( .A1(n80), .A2(n79), .A3(n78), .ZN(carry[14]) );
  XOR2_X1 U109 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U110 ( .A1(B[0]), .A2(A[0]), .ZN(n82) );
endmodule


module datapath_DW_mult_tc_11 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347;

  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n290), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n289), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n293), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n292), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n295), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n94), .B(n88), .CI(n101), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  INV_X1 U157 ( .A(n15), .ZN(n286) );
  AND3_X1 U158 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n216) );
  BUF_X2 U159 ( .A(b[0]), .Z(n279) );
  AND3_X1 U160 ( .A1(n246), .A2(n247), .A3(n248), .ZN(product[15]) );
  CLKBUF_X1 U161 ( .A(n12), .Z(n207) );
  NAND3_X1 U162 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n208) );
  NAND3_X1 U163 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n209) );
  XOR2_X1 U164 ( .A(a[5]), .B(a[4]), .Z(n342) );
  XNOR2_X1 U165 ( .A(n210), .B(n217), .ZN(product[6]) );
  AND3_X1 U166 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n210) );
  NAND2_X2 U167 ( .A1(n324), .A2(n343), .ZN(n326) );
  XNOR2_X1 U168 ( .A(n211), .B(n207), .ZN(product[4]) );
  XNOR2_X1 U169 ( .A(n54), .B(n55), .ZN(n211) );
  NAND3_X1 U170 ( .A1(n218), .A2(n219), .A3(n220), .ZN(n212) );
  NAND3_X1 U171 ( .A1(n218), .A2(n219), .A3(n220), .ZN(n213) );
  BUF_X2 U172 ( .A(a[3]), .Z(n214) );
  NAND3_X1 U173 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n215) );
  XNOR2_X1 U174 ( .A(n216), .B(n245), .ZN(product[14]) );
  XOR2_X1 U175 ( .A(n46), .B(n49), .Z(n217) );
  NAND2_X1 U176 ( .A1(n215), .A2(n46), .ZN(n218) );
  NAND2_X1 U177 ( .A1(n10), .A2(n49), .ZN(n219) );
  NAND2_X1 U178 ( .A1(n46), .A2(n49), .ZN(n220) );
  NAND3_X1 U179 ( .A1(n218), .A2(n219), .A3(n220), .ZN(n9) );
  NAND3_X1 U180 ( .A1(n271), .A2(n270), .A3(n269), .ZN(n221) );
  XNOR2_X1 U181 ( .A(n222), .B(n225), .ZN(product[5]) );
  XNOR2_X1 U182 ( .A(n50), .B(n53), .ZN(n222) );
  CLKBUF_X1 U183 ( .A(n344), .Z(n226) );
  NAND3_X1 U184 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n223) );
  NAND3_X1 U185 ( .A1(n235), .A2(n234), .A3(n233), .ZN(n224) );
  NAND3_X1 U186 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n225) );
  XOR2_X1 U187 ( .A(n27), .B(n24), .Z(n227) );
  XOR2_X1 U188 ( .A(n221), .B(n227), .Z(product[10]) );
  NAND2_X1 U189 ( .A1(n223), .A2(n27), .ZN(n228) );
  NAND2_X1 U190 ( .A1(n6), .A2(n24), .ZN(n229) );
  NAND2_X1 U191 ( .A1(n27), .A2(n24), .ZN(n230) );
  NAND3_X1 U192 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n5) );
  NAND3_X1 U193 ( .A1(n241), .A2(n242), .A3(n240), .ZN(n231) );
  NAND3_X1 U194 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n232) );
  NAND2_X1 U195 ( .A1(n54), .A2(n55), .ZN(n233) );
  NAND2_X1 U196 ( .A1(n54), .A2(n12), .ZN(n234) );
  NAND2_X1 U197 ( .A1(n55), .A2(n12), .ZN(n235) );
  NAND3_X1 U198 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n11) );
  NAND2_X1 U199 ( .A1(n50), .A2(n53), .ZN(n236) );
  NAND2_X1 U200 ( .A1(n224), .A2(n50), .ZN(n237) );
  NAND2_X1 U201 ( .A1(n11), .A2(n53), .ZN(n238) );
  NAND3_X1 U202 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n10) );
  XOR2_X1 U203 ( .A(n40), .B(n45), .Z(n239) );
  XOR2_X1 U204 ( .A(n213), .B(n239), .Z(product[7]) );
  NAND2_X1 U205 ( .A1(n9), .A2(n40), .ZN(n240) );
  NAND2_X1 U206 ( .A1(n212), .A2(n45), .ZN(n241) );
  NAND2_X1 U207 ( .A1(n40), .A2(n45), .ZN(n242) );
  NAND3_X1 U208 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n8) );
  XOR2_X1 U209 ( .A(n243), .B(n244), .Z(product[9]) );
  XNOR2_X1 U210 ( .A(n28), .B(n33), .ZN(n243) );
  AND3_X1 U211 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n244) );
  XOR2_X1 U212 ( .A(n287), .B(n15), .Z(n245) );
  NAND2_X1 U213 ( .A1(n2), .A2(n287), .ZN(n246) );
  NAND2_X1 U214 ( .A1(n2), .A2(n15), .ZN(n247) );
  NAND2_X1 U215 ( .A1(n287), .A2(n15), .ZN(n248) );
  NAND2_X1 U216 ( .A1(a[4]), .A2(a[3]), .ZN(n251) );
  NAND2_X1 U217 ( .A1(n249), .A2(n250), .ZN(n252) );
  NAND2_X2 U218 ( .A1(n251), .A2(n252), .ZN(n313) );
  INV_X1 U219 ( .A(a[4]), .ZN(n249) );
  INV_X1 U220 ( .A(a[3]), .ZN(n250) );
  XNOR2_X1 U221 ( .A(n253), .B(n232), .ZN(product[8]) );
  XNOR2_X1 U222 ( .A(n34), .B(n39), .ZN(n253) );
  NAND3_X1 U223 ( .A1(n259), .A2(n258), .A3(n260), .ZN(n254) );
  NAND3_X1 U224 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n255) );
  NAND3_X1 U225 ( .A1(n263), .A2(n262), .A3(n264), .ZN(n256) );
  XOR2_X1 U226 ( .A(n23), .B(n20), .Z(n257) );
  XOR2_X1 U227 ( .A(n209), .B(n257), .Z(product[11]) );
  NAND2_X1 U228 ( .A1(n5), .A2(n23), .ZN(n258) );
  NAND2_X1 U229 ( .A1(n208), .A2(n20), .ZN(n259) );
  NAND2_X1 U230 ( .A1(n23), .A2(n20), .ZN(n260) );
  XOR2_X1 U231 ( .A(n18), .B(n19), .Z(n261) );
  XOR2_X1 U232 ( .A(n255), .B(n261), .Z(product[12]) );
  NAND2_X1 U233 ( .A1(n254), .A2(n18), .ZN(n262) );
  NAND2_X1 U234 ( .A1(n254), .A2(n19), .ZN(n263) );
  NAND2_X1 U235 ( .A1(n18), .A2(n19), .ZN(n264) );
  NAND3_X1 U236 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n3) );
  NAND3_X1 U237 ( .A1(n267), .A2(n266), .A3(n268), .ZN(n265) );
  NAND2_X1 U238 ( .A1(n34), .A2(n39), .ZN(n266) );
  NAND2_X1 U239 ( .A1(n34), .A2(n231), .ZN(n267) );
  NAND2_X1 U240 ( .A1(n8), .A2(n39), .ZN(n268) );
  NAND3_X1 U241 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n7) );
  NAND2_X1 U242 ( .A1(n28), .A2(n33), .ZN(n269) );
  NAND2_X1 U243 ( .A1(n265), .A2(n28), .ZN(n270) );
  NAND2_X1 U244 ( .A1(n33), .A2(n7), .ZN(n271) );
  NAND3_X1 U245 ( .A1(n271), .A2(n270), .A3(n269), .ZN(n6) );
  XOR2_X1 U246 ( .A(n17), .B(n286), .Z(n272) );
  XOR2_X1 U247 ( .A(n3), .B(n272), .Z(product[13]) );
  NAND2_X1 U248 ( .A1(n256), .A2(n17), .ZN(n273) );
  NAND2_X1 U249 ( .A1(n256), .A2(n286), .ZN(n274) );
  NAND2_X1 U250 ( .A1(n17), .A2(n286), .ZN(n275) );
  NAND3_X1 U251 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n2) );
  CLKBUF_X1 U252 ( .A(b[3]), .Z(n276) );
  NAND2_X1 U253 ( .A1(n283), .A2(n284), .ZN(n277) );
  NAND2_X1 U254 ( .A1(n283), .A2(n284), .ZN(n278) );
  NAND2_X1 U255 ( .A1(n283), .A2(n284), .ZN(n303) );
  INV_X1 U256 ( .A(n31), .ZN(n292) );
  INV_X1 U257 ( .A(n21), .ZN(n289) );
  INV_X1 U258 ( .A(n322), .ZN(n290) );
  INV_X1 U259 ( .A(n333), .ZN(n287) );
  INV_X1 U260 ( .A(n302), .ZN(n295) );
  INV_X1 U261 ( .A(n311), .ZN(n293) );
  INV_X1 U262 ( .A(a[5]), .ZN(n291) );
  INV_X1 U263 ( .A(a[7]), .ZN(n288) );
  INV_X1 U264 ( .A(b[0]), .ZN(n285) );
  NAND2_X1 U265 ( .A1(n277), .A2(n341), .ZN(n280) );
  NAND2_X1 U266 ( .A1(a[2]), .A2(a[1]), .ZN(n283) );
  NAND2_X1 U267 ( .A1(n281), .A2(n282), .ZN(n284) );
  INV_X1 U268 ( .A(a[2]), .ZN(n281) );
  INV_X1 U269 ( .A(a[1]), .ZN(n282) );
  NAND2_X1 U270 ( .A1(n303), .A2(n341), .ZN(n305) );
  INV_X1 U271 ( .A(a[3]), .ZN(n294) );
  NAND2_X2 U272 ( .A1(n313), .A2(n342), .ZN(n315) );
  INV_X1 U273 ( .A(a[1]), .ZN(n296) );
  XOR2_X2 U274 ( .A(a[6]), .B(n291), .Z(n324) );
  INV_X2 U275 ( .A(a[0]), .ZN(n297) );
  NOR2_X1 U276 ( .A1(n297), .A2(n285), .ZN(product[0]) );
  OAI22_X1 U277 ( .A1(n298), .A2(n299), .B1(n300), .B2(n297), .ZN(n99) );
  OAI22_X1 U278 ( .A1(n300), .A2(n299), .B1(n301), .B2(n297), .ZN(n98) );
  XNOR2_X1 U279 ( .A(b[6]), .B(a[1]), .ZN(n300) );
  OAI22_X1 U280 ( .A1(n297), .A2(n301), .B1(n299), .B2(n301), .ZN(n302) );
  XNOR2_X1 U281 ( .A(b[7]), .B(a[1]), .ZN(n301) );
  NOR2_X1 U282 ( .A1(n278), .A2(n285), .ZN(n96) );
  OAI22_X1 U283 ( .A1(n304), .A2(n305), .B1(n278), .B2(n306), .ZN(n95) );
  XNOR2_X1 U284 ( .A(n214), .B(n279), .ZN(n304) );
  OAI22_X1 U285 ( .A1(n306), .A2(n280), .B1(n277), .B2(n307), .ZN(n94) );
  XNOR2_X1 U286 ( .A(b[1]), .B(n214), .ZN(n306) );
  OAI22_X1 U287 ( .A1(n307), .A2(n305), .B1(n277), .B2(n308), .ZN(n93) );
  XNOR2_X1 U288 ( .A(b[2]), .B(n214), .ZN(n307) );
  OAI22_X1 U289 ( .A1(n308), .A2(n280), .B1(n278), .B2(n309), .ZN(n92) );
  XNOR2_X1 U290 ( .A(b[3]), .B(n214), .ZN(n308) );
  OAI22_X1 U291 ( .A1(n309), .A2(n280), .B1(n278), .B2(n310), .ZN(n91) );
  XNOR2_X1 U292 ( .A(b[4]), .B(n214), .ZN(n309) );
  OAI22_X1 U293 ( .A1(n312), .A2(n277), .B1(n305), .B2(n312), .ZN(n311) );
  NOR2_X1 U294 ( .A1(n313), .A2(n285), .ZN(n88) );
  OAI22_X1 U295 ( .A1(n314), .A2(n315), .B1(n313), .B2(n316), .ZN(n87) );
  XNOR2_X1 U296 ( .A(a[5]), .B(n279), .ZN(n314) );
  OAI22_X1 U297 ( .A1(n316), .A2(n315), .B1(n313), .B2(n317), .ZN(n86) );
  XNOR2_X1 U298 ( .A(b[1]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U299 ( .A1(n317), .A2(n315), .B1(n313), .B2(n318), .ZN(n85) );
  XNOR2_X1 U300 ( .A(b[2]), .B(a[5]), .ZN(n317) );
  OAI22_X1 U301 ( .A1(n318), .A2(n315), .B1(n313), .B2(n319), .ZN(n84) );
  XNOR2_X1 U302 ( .A(b[3]), .B(a[5]), .ZN(n318) );
  OAI22_X1 U303 ( .A1(n319), .A2(n315), .B1(n313), .B2(n320), .ZN(n83) );
  XNOR2_X1 U304 ( .A(b[4]), .B(a[5]), .ZN(n319) );
  OAI22_X1 U305 ( .A1(n320), .A2(n315), .B1(n313), .B2(n321), .ZN(n82) );
  XNOR2_X1 U306 ( .A(b[5]), .B(a[5]), .ZN(n320) );
  OAI22_X1 U307 ( .A1(n323), .A2(n313), .B1(n315), .B2(n323), .ZN(n322) );
  NOR2_X1 U308 ( .A1(n324), .A2(n285), .ZN(n80) );
  OAI22_X1 U309 ( .A1(n325), .A2(n326), .B1(n324), .B2(n327), .ZN(n79) );
  XNOR2_X1 U310 ( .A(a[7]), .B(n279), .ZN(n325) );
  OAI22_X1 U311 ( .A1(n328), .A2(n326), .B1(n324), .B2(n329), .ZN(n77) );
  OAI22_X1 U312 ( .A1(n329), .A2(n326), .B1(n324), .B2(n330), .ZN(n76) );
  XNOR2_X1 U313 ( .A(n276), .B(a[7]), .ZN(n329) );
  OAI22_X1 U314 ( .A1(n330), .A2(n326), .B1(n324), .B2(n331), .ZN(n75) );
  XNOR2_X1 U315 ( .A(b[4]), .B(a[7]), .ZN(n330) );
  OAI22_X1 U316 ( .A1(n331), .A2(n326), .B1(n324), .B2(n332), .ZN(n74) );
  XNOR2_X1 U317 ( .A(b[5]), .B(a[7]), .ZN(n331) );
  OAI22_X1 U318 ( .A1(n334), .A2(n324), .B1(n326), .B2(n334), .ZN(n333) );
  OAI21_X1 U319 ( .B1(n279), .B2(n296), .A(n299), .ZN(n72) );
  OAI21_X1 U320 ( .B1(n294), .B2(n305), .A(n335), .ZN(n71) );
  OR3_X1 U321 ( .A1(n278), .A2(n279), .A3(n294), .ZN(n335) );
  OAI21_X1 U322 ( .B1(n291), .B2(n315), .A(n336), .ZN(n70) );
  OR3_X1 U323 ( .A1(n313), .A2(n279), .A3(n291), .ZN(n336) );
  OAI21_X1 U324 ( .B1(n288), .B2(n326), .A(n337), .ZN(n69) );
  OR3_X1 U325 ( .A1(n324), .A2(n279), .A3(n288), .ZN(n337) );
  XNOR2_X1 U326 ( .A(n338), .B(n339), .ZN(n38) );
  OR2_X1 U327 ( .A1(n338), .A2(n339), .ZN(n37) );
  OAI22_X1 U328 ( .A1(n310), .A2(n280), .B1(n277), .B2(n340), .ZN(n339) );
  XNOR2_X1 U329 ( .A(b[5]), .B(n214), .ZN(n310) );
  OAI22_X1 U330 ( .A1(n327), .A2(n326), .B1(n324), .B2(n328), .ZN(n338) );
  XNOR2_X1 U331 ( .A(b[2]), .B(a[7]), .ZN(n328) );
  XNOR2_X1 U332 ( .A(b[1]), .B(a[7]), .ZN(n327) );
  OAI22_X1 U333 ( .A1(n340), .A2(n305), .B1(n278), .B2(n312), .ZN(n31) );
  XNOR2_X1 U334 ( .A(b[7]), .B(n214), .ZN(n312) );
  XNOR2_X1 U335 ( .A(n294), .B(a[2]), .ZN(n341) );
  XNOR2_X1 U336 ( .A(b[6]), .B(n214), .ZN(n340) );
  OAI22_X1 U337 ( .A1(n321), .A2(n315), .B1(n313), .B2(n323), .ZN(n21) );
  XNOR2_X1 U338 ( .A(b[7]), .B(a[5]), .ZN(n323) );
  XNOR2_X1 U339 ( .A(b[6]), .B(a[5]), .ZN(n321) );
  OAI22_X1 U340 ( .A1(n332), .A2(n326), .B1(n324), .B2(n334), .ZN(n15) );
  XNOR2_X1 U341 ( .A(b[7]), .B(a[7]), .ZN(n334) );
  XNOR2_X1 U342 ( .A(n288), .B(a[6]), .ZN(n343) );
  XNOR2_X1 U343 ( .A(b[6]), .B(a[7]), .ZN(n332) );
  OAI22_X1 U344 ( .A1(n279), .A2(n299), .B1(n344), .B2(n297), .ZN(n104) );
  OAI22_X1 U345 ( .A1(n226), .A2(n299), .B1(n345), .B2(n297), .ZN(n103) );
  XNOR2_X1 U346 ( .A(b[1]), .B(a[1]), .ZN(n344) );
  OAI22_X1 U347 ( .A1(n345), .A2(n299), .B1(n346), .B2(n297), .ZN(n102) );
  XNOR2_X1 U348 ( .A(b[2]), .B(a[1]), .ZN(n345) );
  OAI22_X1 U349 ( .A1(n346), .A2(n299), .B1(n347), .B2(n297), .ZN(n101) );
  XNOR2_X1 U350 ( .A(b[3]), .B(a[1]), .ZN(n346) );
  OAI22_X1 U351 ( .A1(n347), .A2(n299), .B1(n298), .B2(n297), .ZN(n100) );
  XNOR2_X1 U352 ( .A(b[5]), .B(a[1]), .ZN(n298) );
  NAND2_X1 U353 ( .A1(a[1]), .A2(n297), .ZN(n299) );
  XNOR2_X1 U354 ( .A(b[4]), .B(a[1]), .ZN(n347) );
endmodule


module datapath_DW01_add_11 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n80;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n80), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(n37), .Z(n1) );
  NAND3_X1 U2 ( .A1(n77), .A2(n76), .A3(n75), .ZN(n2) );
  NAND3_X1 U3 ( .A1(n10), .A2(n11), .A3(n12), .ZN(n3) );
  NAND3_X1 U4 ( .A1(n10), .A2(n11), .A3(n12), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n18), .A2(B[10]), .ZN(n5) );
  CLKBUF_X1 U6 ( .A(n18), .Z(n6) );
  CLKBUF_X1 U7 ( .A(n67), .Z(n7) );
  CLKBUF_X1 U8 ( .A(B[4]), .Z(n8) );
  XOR2_X1 U9 ( .A(carry[2]), .B(A[2]), .Z(n9) );
  XOR2_X1 U10 ( .A(B[2]), .B(n9), .Z(SUM[2]) );
  NAND2_X1 U11 ( .A1(B[2]), .A2(carry[2]), .ZN(n10) );
  NAND2_X1 U12 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  NAND2_X1 U13 ( .A1(carry[2]), .A2(A[2]), .ZN(n12) );
  NAND3_X1 U14 ( .A1(n10), .A2(n11), .A3(n12), .ZN(carry[3]) );
  CLKBUF_X1 U15 ( .A(n5), .Z(n13) );
  CLKBUF_X1 U16 ( .A(n43), .Z(n14) );
  XNOR2_X1 U17 ( .A(B[15]), .B(A[15]), .ZN(n78) );
  NAND3_X1 U18 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n15) );
  NAND3_X1 U19 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n16) );
  NAND3_X1 U20 ( .A1(n42), .A2(n14), .A3(n44), .ZN(n17) );
  NAND3_X1 U21 ( .A1(n23), .A2(n24), .A3(n25), .ZN(n18) );
  NAND3_X1 U22 ( .A1(n36), .A2(n37), .A3(n38), .ZN(n19) );
  CLKBUF_X1 U23 ( .A(n72), .Z(n20) );
  CLKBUF_X1 U24 ( .A(n15), .Z(n21) );
  XOR2_X1 U25 ( .A(B[9]), .B(A[9]), .Z(n22) );
  XOR2_X1 U26 ( .A(n17), .B(n22), .Z(SUM[9]) );
  NAND2_X1 U27 ( .A1(n16), .A2(B[9]), .ZN(n23) );
  NAND2_X1 U28 ( .A1(carry[9]), .A2(A[9]), .ZN(n24) );
  NAND2_X1 U29 ( .A1(B[9]), .A2(A[9]), .ZN(n25) );
  NAND3_X1 U30 ( .A1(n24), .A2(n23), .A3(n25), .ZN(carry[10]) );
  CLKBUF_X1 U31 ( .A(n76), .Z(n26) );
  XOR2_X1 U32 ( .A(n8), .B(A[4]), .Z(n27) );
  XOR2_X1 U33 ( .A(carry[4]), .B(n27), .Z(SUM[4]) );
  NAND2_X1 U34 ( .A1(n19), .A2(B[4]), .ZN(n28) );
  NAND2_X1 U35 ( .A1(n19), .A2(A[4]), .ZN(n29) );
  NAND2_X1 U36 ( .A1(B[4]), .A2(A[4]), .ZN(n30) );
  NAND3_X1 U37 ( .A1(n29), .A2(n28), .A3(n30), .ZN(carry[5]) );
  CLKBUF_X1 U38 ( .A(n40), .Z(n31) );
  NAND3_X1 U39 ( .A1(n77), .A2(n76), .A3(n75), .ZN(n32) );
  NAND3_X1 U40 ( .A1(n5), .A2(n51), .A3(n52), .ZN(n33) );
  NAND3_X1 U41 ( .A1(n13), .A2(n51), .A3(n52), .ZN(n34) );
  XOR2_X1 U42 ( .A(B[3]), .B(A[3]), .Z(n35) );
  XOR2_X1 U43 ( .A(n4), .B(n35), .Z(SUM[3]) );
  NAND2_X1 U44 ( .A1(n3), .A2(B[3]), .ZN(n36) );
  NAND2_X1 U45 ( .A1(carry[3]), .A2(A[3]), .ZN(n37) );
  NAND2_X1 U46 ( .A1(B[3]), .A2(A[3]), .ZN(n38) );
  NAND3_X1 U47 ( .A1(n36), .A2(n1), .A3(n38), .ZN(carry[4]) );
  NAND3_X1 U48 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n39) );
  NAND3_X1 U49 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n40) );
  XOR2_X1 U50 ( .A(B[8]), .B(A[8]), .Z(n41) );
  XOR2_X1 U51 ( .A(carry[8]), .B(n41), .Z(SUM[8]) );
  NAND2_X1 U52 ( .A1(n2), .A2(B[8]), .ZN(n42) );
  NAND2_X1 U53 ( .A1(n32), .A2(A[8]), .ZN(n43) );
  NAND2_X1 U54 ( .A1(B[8]), .A2(A[8]), .ZN(n44) );
  NAND3_X1 U55 ( .A1(n42), .A2(n43), .A3(n44), .ZN(carry[9]) );
  XOR2_X1 U56 ( .A(B[12]), .B(A[12]), .Z(n45) );
  XOR2_X1 U57 ( .A(n31), .B(n45), .Z(SUM[12]) );
  NAND2_X1 U58 ( .A1(n40), .A2(B[12]), .ZN(n46) );
  NAND2_X1 U59 ( .A1(carry[12]), .A2(A[12]), .ZN(n47) );
  NAND2_X1 U60 ( .A1(B[12]), .A2(A[12]), .ZN(n48) );
  NAND3_X1 U61 ( .A1(n46), .A2(n47), .A3(n48), .ZN(carry[13]) );
  XOR2_X1 U62 ( .A(B[10]), .B(A[10]), .Z(n49) );
  XOR2_X1 U63 ( .A(n6), .B(n49), .Z(SUM[10]) );
  NAND2_X1 U64 ( .A1(n18), .A2(B[10]), .ZN(n50) );
  NAND2_X1 U65 ( .A1(carry[10]), .A2(A[10]), .ZN(n51) );
  NAND2_X1 U66 ( .A1(B[10]), .A2(A[10]), .ZN(n52) );
  NAND3_X1 U67 ( .A1(n50), .A2(n51), .A3(n52), .ZN(carry[11]) );
  XOR2_X1 U68 ( .A(B[11]), .B(A[11]), .Z(n53) );
  XOR2_X1 U69 ( .A(n34), .B(n53), .Z(SUM[11]) );
  NAND2_X1 U70 ( .A1(n33), .A2(B[11]), .ZN(n54) );
  NAND2_X1 U71 ( .A1(carry[11]), .A2(A[11]), .ZN(n55) );
  NAND2_X1 U72 ( .A1(B[11]), .A2(A[11]), .ZN(n56) );
  NAND3_X1 U73 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[12]) );
  CLKBUF_X1 U74 ( .A(n39), .Z(n57) );
  XOR2_X1 U75 ( .A(B[13]), .B(A[13]), .Z(n58) );
  XOR2_X1 U76 ( .A(n57), .B(n58), .Z(SUM[13]) );
  NAND2_X1 U77 ( .A1(n39), .A2(B[13]), .ZN(n59) );
  NAND2_X1 U78 ( .A1(carry[13]), .A2(A[13]), .ZN(n60) );
  NAND2_X1 U79 ( .A1(B[13]), .A2(A[13]), .ZN(n61) );
  NAND3_X1 U80 ( .A1(n59), .A2(n60), .A3(n61), .ZN(carry[14]) );
  NAND3_X1 U81 ( .A1(n73), .A2(n72), .A3(n71), .ZN(n62) );
  NAND3_X1 U82 ( .A1(n73), .A2(n20), .A3(n71), .ZN(n63) );
  NAND3_X1 U83 ( .A1(n67), .A2(n69), .A3(n68), .ZN(n64) );
  NAND3_X1 U84 ( .A1(n7), .A2(n68), .A3(n69), .ZN(n65) );
  XOR2_X1 U85 ( .A(B[5]), .B(A[5]), .Z(n66) );
  XOR2_X1 U86 ( .A(n21), .B(n66), .Z(SUM[5]) );
  NAND2_X1 U87 ( .A1(n15), .A2(B[5]), .ZN(n67) );
  NAND2_X1 U88 ( .A1(carry[5]), .A2(A[5]), .ZN(n68) );
  NAND2_X1 U89 ( .A1(B[5]), .A2(A[5]), .ZN(n69) );
  NAND3_X1 U90 ( .A1(n67), .A2(n68), .A3(n69), .ZN(carry[6]) );
  XOR2_X1 U91 ( .A(A[6]), .B(B[6]), .Z(n70) );
  XOR2_X1 U92 ( .A(n70), .B(n65), .Z(SUM[6]) );
  NAND2_X1 U93 ( .A1(A[6]), .A2(B[6]), .ZN(n71) );
  NAND2_X1 U94 ( .A1(A[6]), .A2(carry[6]), .ZN(n72) );
  NAND2_X1 U95 ( .A1(B[6]), .A2(n64), .ZN(n73) );
  NAND3_X1 U96 ( .A1(n73), .A2(n72), .A3(n71), .ZN(carry[7]) );
  XOR2_X1 U97 ( .A(A[7]), .B(B[7]), .Z(n74) );
  XOR2_X1 U98 ( .A(n74), .B(n63), .Z(SUM[7]) );
  NAND2_X1 U99 ( .A1(A[7]), .A2(B[7]), .ZN(n75) );
  NAND2_X1 U100 ( .A1(A[7]), .A2(n62), .ZN(n76) );
  NAND2_X1 U101 ( .A1(B[7]), .A2(carry[7]), .ZN(n77) );
  NAND3_X1 U102 ( .A1(n77), .A2(n26), .A3(n75), .ZN(carry[8]) );
  XNOR2_X1 U103 ( .A(carry[15]), .B(n78), .ZN(SUM[15]) );
  XOR2_X1 U104 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U105 ( .A1(B[0]), .A2(A[0]), .ZN(n80) );
endmodule


module datapath_DW_mult_tc_10 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n6, n7, n9, n10, n11, n12, n13, n14, n15, n17, n18, n19,
         n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76, n77,
         n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94, n95,
         n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208, n209,
         n210, n211, n212, n213, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355;

  FA_X1 U13 ( .A(n13), .B(n71), .CI(n56), .CO(n12), .S(product[3]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n298), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n297), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n301), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n300), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n303), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n92), .B(n80), .CI(n99), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n94), .B(n88), .CI(n101), .CO(n53), .S(n54) );
  CLKBUF_X1 U157 ( .A(b[2]), .Z(n206) );
  XNOR2_X1 U158 ( .A(n207), .B(n221), .ZN(product[8]) );
  XNOR2_X1 U159 ( .A(n34), .B(n39), .ZN(n207) );
  BUF_X2 U160 ( .A(a[3]), .Z(n227) );
  NAND3_X1 U161 ( .A1(n289), .A2(n290), .A3(n291), .ZN(n49) );
  NAND2_X1 U162 ( .A1(n311), .A2(n349), .ZN(n313) );
  AND2_X1 U163 ( .A1(n104), .A2(n72), .ZN(n208) );
  CLKBUF_X1 U164 ( .A(n52), .Z(n209) );
  OAI22_X1 U165 ( .A1(n231), .A2(n307), .B1(n353), .B2(n305), .ZN(n210) );
  CLKBUF_X1 U166 ( .A(n293), .Z(n271) );
  NAND2_X2 U167 ( .A1(a[1]), .A2(n211), .ZN(n307) );
  NAND2_X2 U168 ( .A1(n321), .A2(n350), .ZN(n323) );
  BUF_X2 U169 ( .A(n311), .Z(n292) );
  INV_X1 U170 ( .A(a[0]), .ZN(n211) );
  INV_X1 U171 ( .A(a[0]), .ZN(n305) );
  AND2_X1 U172 ( .A1(n250), .A2(n102), .ZN(n212) );
  XNOR2_X1 U173 ( .A(n295), .B(n15), .ZN(n213) );
  AND3_X1 U174 ( .A1(n267), .A2(n268), .A3(n269), .ZN(product[15]) );
  XNOR2_X1 U175 ( .A(n14), .B(n215), .ZN(product[2]) );
  XNOR2_X1 U176 ( .A(n210), .B(n96), .ZN(n215) );
  NAND2_X1 U177 ( .A1(n208), .A2(n103), .ZN(n216) );
  NAND2_X1 U178 ( .A1(n208), .A2(n96), .ZN(n217) );
  NAND2_X1 U179 ( .A1(n103), .A2(n96), .ZN(n218) );
  NAND3_X1 U180 ( .A1(n216), .A2(n217), .A3(n218), .ZN(n13) );
  XNOR2_X1 U181 ( .A(a[6]), .B(a[5]), .ZN(n332) );
  XNOR2_X1 U182 ( .A(a[6]), .B(a[5]), .ZN(n219) );
  XNOR2_X1 U183 ( .A(n220), .B(n12), .ZN(product[4]) );
  XNOR2_X1 U184 ( .A(n54), .B(n212), .ZN(n220) );
  NAND3_X1 U185 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n221) );
  NAND2_X1 U186 ( .A1(n266), .A2(n39), .ZN(n222) );
  CLKBUF_X1 U187 ( .A(b[1]), .Z(n223) );
  INV_X1 U188 ( .A(n304), .ZN(n224) );
  INV_X1 U189 ( .A(n293), .ZN(n225) );
  NAND3_X1 U190 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n226) );
  NAND3_X1 U191 ( .A1(n283), .A2(n284), .A3(n285), .ZN(n228) );
  NAND3_X1 U192 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n229) );
  NAND3_X1 U193 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n230) );
  XNOR2_X1 U194 ( .A(b[1]), .B(a[1]), .ZN(n231) );
  NAND3_X1 U195 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n232) );
  NAND3_X1 U196 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n233) );
  NAND3_X1 U197 ( .A1(n246), .A2(n245), .A3(n247), .ZN(n234) );
  NAND3_X1 U198 ( .A1(n246), .A2(n245), .A3(n247), .ZN(n235) );
  CLKBUF_X1 U199 ( .A(n95), .Z(n250) );
  XOR2_X1 U200 ( .A(n19), .B(n18), .Z(n236) );
  XOR2_X1 U201 ( .A(n236), .B(n232), .Z(product[12]) );
  NAND2_X1 U202 ( .A1(n19), .A2(n18), .ZN(n237) );
  NAND2_X1 U203 ( .A1(n19), .A2(n4), .ZN(n238) );
  NAND2_X1 U204 ( .A1(n18), .A2(n4), .ZN(n239) );
  NAND3_X1 U205 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n3) );
  XOR2_X1 U206 ( .A(n17), .B(n294), .Z(n240) );
  XOR2_X1 U207 ( .A(n240), .B(n233), .Z(product[13]) );
  NAND2_X1 U208 ( .A1(n17), .A2(n294), .ZN(n241) );
  NAND2_X1 U209 ( .A1(n17), .A2(n3), .ZN(n242) );
  NAND2_X1 U210 ( .A1(n294), .A2(n3), .ZN(n243) );
  NAND3_X1 U211 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n2) );
  XNOR2_X1 U212 ( .A(n2), .B(n213), .ZN(product[14]) );
  XOR2_X1 U213 ( .A(n46), .B(n49), .Z(n244) );
  XOR2_X1 U214 ( .A(n10), .B(n244), .Z(product[6]) );
  NAND2_X1 U215 ( .A1(n228), .A2(n46), .ZN(n245) );
  NAND2_X1 U216 ( .A1(n10), .A2(n49), .ZN(n246) );
  NAND2_X1 U217 ( .A1(n46), .A2(n49), .ZN(n247) );
  NAND3_X1 U218 ( .A1(n246), .A2(n245), .A3(n247), .ZN(n9) );
  NAND3_X1 U219 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n248) );
  NAND3_X1 U220 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n249) );
  XOR2_X1 U221 ( .A(n95), .B(n102), .Z(n56) );
  XOR2_X1 U222 ( .A(n27), .B(n24), .Z(n251) );
  XOR2_X1 U223 ( .A(n229), .B(n251), .Z(product[10]) );
  NAND2_X1 U224 ( .A1(n229), .A2(n27), .ZN(n252) );
  NAND2_X1 U225 ( .A1(n6), .A2(n24), .ZN(n253) );
  NAND2_X1 U226 ( .A1(n27), .A2(n24), .ZN(n254) );
  NAND3_X1 U227 ( .A1(n277), .A2(n222), .A3(n276), .ZN(n255) );
  NAND3_X1 U228 ( .A1(n277), .A2(n276), .A3(n222), .ZN(n256) );
  XOR2_X1 U229 ( .A(n33), .B(n28), .Z(n257) );
  XOR2_X1 U230 ( .A(n256), .B(n257), .Z(product[9]) );
  NAND2_X1 U231 ( .A1(n255), .A2(n33), .ZN(n258) );
  NAND2_X1 U232 ( .A1(n7), .A2(n28), .ZN(n259) );
  NAND2_X1 U233 ( .A1(n33), .A2(n28), .ZN(n260) );
  NAND3_X1 U234 ( .A1(n259), .A2(n258), .A3(n260), .ZN(n6) );
  XOR2_X1 U235 ( .A(n23), .B(n20), .Z(n261) );
  XOR2_X1 U236 ( .A(n248), .B(n261), .Z(product[11]) );
  NAND2_X1 U237 ( .A1(n248), .A2(n23), .ZN(n262) );
  NAND2_X1 U238 ( .A1(n249), .A2(n20), .ZN(n263) );
  NAND2_X1 U239 ( .A1(n23), .A2(n20), .ZN(n264) );
  NAND3_X1 U240 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n4) );
  NAND3_X1 U241 ( .A1(n275), .A2(n274), .A3(n273), .ZN(n265) );
  NAND3_X1 U242 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n266) );
  NAND2_X1 U243 ( .A1(n230), .A2(n295), .ZN(n267) );
  NAND2_X1 U244 ( .A1(n230), .A2(n15), .ZN(n268) );
  NAND2_X1 U245 ( .A1(n295), .A2(n15), .ZN(n269) );
  NAND3_X1 U246 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n270) );
  XOR2_X1 U247 ( .A(n40), .B(n45), .Z(n272) );
  XOR2_X1 U248 ( .A(n272), .B(n235), .Z(product[7]) );
  NAND2_X1 U249 ( .A1(n40), .A2(n45), .ZN(n273) );
  NAND2_X1 U250 ( .A1(n40), .A2(n234), .ZN(n274) );
  NAND2_X1 U251 ( .A1(n45), .A2(n9), .ZN(n275) );
  NAND2_X1 U252 ( .A1(n34), .A2(n39), .ZN(n276) );
  NAND2_X1 U253 ( .A1(n34), .A2(n265), .ZN(n277) );
  NAND2_X1 U254 ( .A1(n221), .A2(n39), .ZN(n278) );
  NAND3_X1 U255 ( .A1(n277), .A2(n278), .A3(n276), .ZN(n7) );
  NAND2_X1 U256 ( .A1(n54), .A2(n212), .ZN(n279) );
  NAND2_X1 U257 ( .A1(n54), .A2(n12), .ZN(n280) );
  NAND2_X1 U258 ( .A1(n12), .A2(n212), .ZN(n281) );
  NAND3_X1 U259 ( .A1(n280), .A2(n279), .A3(n281), .ZN(n11) );
  XOR2_X1 U260 ( .A(n50), .B(n53), .Z(n282) );
  XOR2_X1 U261 ( .A(n282), .B(n226), .Z(product[5]) );
  NAND2_X1 U262 ( .A1(n50), .A2(n53), .ZN(n283) );
  NAND2_X1 U263 ( .A1(n270), .A2(n50), .ZN(n284) );
  NAND2_X1 U264 ( .A1(n53), .A2(n11), .ZN(n285) );
  NAND3_X1 U265 ( .A1(n284), .A2(n283), .A3(n285), .ZN(n10) );
  CLKBUF_X1 U266 ( .A(n313), .Z(n286) );
  INV_X1 U267 ( .A(n293), .ZN(n287) );
  XNOR2_X2 U268 ( .A(a[4]), .B(a[3]), .ZN(n321) );
  XNOR2_X1 U269 ( .A(n52), .B(n288), .ZN(n50) );
  XNOR2_X1 U270 ( .A(n93), .B(n100), .ZN(n288) );
  INV_X1 U271 ( .A(n15), .ZN(n294) );
  INV_X1 U272 ( .A(n319), .ZN(n301) );
  INV_X1 U273 ( .A(n31), .ZN(n300) );
  INV_X1 U274 ( .A(n21), .ZN(n297) );
  INV_X1 U275 ( .A(n330), .ZN(n298) );
  INV_X1 U276 ( .A(n341), .ZN(n295) );
  INV_X1 U277 ( .A(n310), .ZN(n303) );
  INV_X1 U278 ( .A(a[5]), .ZN(n299) );
  INV_X1 U279 ( .A(a[7]), .ZN(n296) );
  INV_X1 U280 ( .A(b[0]), .ZN(n293) );
  NAND2_X1 U281 ( .A1(n209), .A2(n93), .ZN(n289) );
  NAND2_X1 U282 ( .A1(n209), .A2(n100), .ZN(n290) );
  NAND2_X1 U283 ( .A1(n93), .A2(n100), .ZN(n291) );
  XNOR2_X1 U284 ( .A(a[2]), .B(a[1]), .ZN(n311) );
  INV_X1 U285 ( .A(a[3]), .ZN(n302) );
  INV_X1 U286 ( .A(a[1]), .ZN(n304) );
  NOR2_X1 U287 ( .A1(n305), .A2(n271), .ZN(product[0]) );
  OAI22_X1 U288 ( .A1(n306), .A2(n307), .B1(n308), .B2(n305), .ZN(n99) );
  OAI22_X1 U289 ( .A1(n308), .A2(n307), .B1(n309), .B2(n305), .ZN(n98) );
  XNOR2_X1 U290 ( .A(b[6]), .B(n224), .ZN(n308) );
  OAI22_X1 U291 ( .A1(n305), .A2(n309), .B1(n307), .B2(n309), .ZN(n310) );
  XNOR2_X1 U292 ( .A(b[7]), .B(n224), .ZN(n309) );
  NOR2_X1 U293 ( .A1(n292), .A2(n271), .ZN(n96) );
  OAI22_X1 U294 ( .A1(n312), .A2(n313), .B1(n292), .B2(n314), .ZN(n95) );
  XNOR2_X1 U295 ( .A(n227), .B(n225), .ZN(n312) );
  OAI22_X1 U296 ( .A1(n314), .A2(n313), .B1(n292), .B2(n315), .ZN(n94) );
  XNOR2_X1 U297 ( .A(b[1]), .B(n227), .ZN(n314) );
  OAI22_X1 U298 ( .A1(n315), .A2(n313), .B1(n292), .B2(n316), .ZN(n93) );
  XNOR2_X1 U299 ( .A(b[2]), .B(n227), .ZN(n315) );
  OAI22_X1 U300 ( .A1(n316), .A2(n313), .B1(n292), .B2(n317), .ZN(n92) );
  XNOR2_X1 U301 ( .A(b[3]), .B(n227), .ZN(n316) );
  OAI22_X1 U302 ( .A1(n317), .A2(n313), .B1(n292), .B2(n318), .ZN(n91) );
  XNOR2_X1 U303 ( .A(b[4]), .B(n227), .ZN(n317) );
  OAI22_X1 U304 ( .A1(n320), .A2(n292), .B1(n286), .B2(n320), .ZN(n319) );
  NOR2_X1 U305 ( .A1(n321), .A2(n271), .ZN(n88) );
  OAI22_X1 U306 ( .A1(n322), .A2(n323), .B1(n321), .B2(n324), .ZN(n87) );
  XNOR2_X1 U307 ( .A(a[5]), .B(n287), .ZN(n322) );
  OAI22_X1 U308 ( .A1(n324), .A2(n323), .B1(n321), .B2(n325), .ZN(n86) );
  XNOR2_X1 U309 ( .A(b[1]), .B(a[5]), .ZN(n324) );
  OAI22_X1 U310 ( .A1(n325), .A2(n323), .B1(n321), .B2(n326), .ZN(n85) );
  XNOR2_X1 U311 ( .A(n206), .B(a[5]), .ZN(n325) );
  OAI22_X1 U312 ( .A1(n326), .A2(n323), .B1(n321), .B2(n327), .ZN(n84) );
  XNOR2_X1 U313 ( .A(b[3]), .B(a[5]), .ZN(n326) );
  OAI22_X1 U314 ( .A1(n327), .A2(n323), .B1(n321), .B2(n328), .ZN(n83) );
  XNOR2_X1 U315 ( .A(b[4]), .B(a[5]), .ZN(n327) );
  OAI22_X1 U316 ( .A1(n328), .A2(n323), .B1(n321), .B2(n329), .ZN(n82) );
  XNOR2_X1 U317 ( .A(b[5]), .B(a[5]), .ZN(n328) );
  OAI22_X1 U318 ( .A1(n331), .A2(n321), .B1(n323), .B2(n331), .ZN(n330) );
  NOR2_X1 U319 ( .A1(n332), .A2(n271), .ZN(n80) );
  OAI22_X1 U320 ( .A1(n333), .A2(n334), .B1(n219), .B2(n335), .ZN(n79) );
  XNOR2_X1 U321 ( .A(a[7]), .B(n287), .ZN(n333) );
  OAI22_X1 U322 ( .A1(n336), .A2(n334), .B1(n219), .B2(n337), .ZN(n77) );
  OAI22_X1 U323 ( .A1(n337), .A2(n334), .B1(n219), .B2(n338), .ZN(n76) );
  XNOR2_X1 U324 ( .A(b[3]), .B(a[7]), .ZN(n337) );
  OAI22_X1 U325 ( .A1(n338), .A2(n334), .B1(n219), .B2(n339), .ZN(n75) );
  XNOR2_X1 U326 ( .A(b[4]), .B(a[7]), .ZN(n338) );
  OAI22_X1 U327 ( .A1(n339), .A2(n334), .B1(n219), .B2(n340), .ZN(n74) );
  XNOR2_X1 U328 ( .A(b[5]), .B(a[7]), .ZN(n339) );
  OAI22_X1 U329 ( .A1(n342), .A2(n219), .B1(n334), .B2(n342), .ZN(n341) );
  OAI21_X1 U330 ( .B1(n287), .B2(n304), .A(n307), .ZN(n72) );
  OAI21_X1 U331 ( .B1(n302), .B2(n313), .A(n343), .ZN(n71) );
  OR3_X1 U332 ( .A1(n292), .A2(n225), .A3(n302), .ZN(n343) );
  OAI21_X1 U333 ( .B1(n299), .B2(n323), .A(n344), .ZN(n70) );
  OR3_X1 U334 ( .A1(n321), .A2(n287), .A3(n299), .ZN(n344) );
  OAI21_X1 U335 ( .B1(n296), .B2(n334), .A(n345), .ZN(n69) );
  OR3_X1 U336 ( .A1(n219), .A2(n287), .A3(n296), .ZN(n345) );
  XNOR2_X1 U337 ( .A(n346), .B(n347), .ZN(n38) );
  OR2_X1 U338 ( .A1(n346), .A2(n347), .ZN(n37) );
  OAI22_X1 U339 ( .A1(n318), .A2(n286), .B1(n292), .B2(n348), .ZN(n347) );
  XNOR2_X1 U340 ( .A(b[5]), .B(n227), .ZN(n318) );
  OAI22_X1 U341 ( .A1(n335), .A2(n334), .B1(n219), .B2(n336), .ZN(n346) );
  XNOR2_X1 U342 ( .A(n206), .B(a[7]), .ZN(n336) );
  XNOR2_X1 U343 ( .A(n223), .B(a[7]), .ZN(n335) );
  OAI22_X1 U344 ( .A1(n348), .A2(n286), .B1(n292), .B2(n320), .ZN(n31) );
  XNOR2_X1 U345 ( .A(b[7]), .B(n227), .ZN(n320) );
  XNOR2_X1 U346 ( .A(n302), .B(a[2]), .ZN(n349) );
  XNOR2_X1 U347 ( .A(b[6]), .B(n227), .ZN(n348) );
  OAI22_X1 U348 ( .A1(n329), .A2(n323), .B1(n321), .B2(n331), .ZN(n21) );
  XNOR2_X1 U349 ( .A(b[7]), .B(a[5]), .ZN(n331) );
  XNOR2_X1 U350 ( .A(n299), .B(a[4]), .ZN(n350) );
  XNOR2_X1 U351 ( .A(b[6]), .B(a[5]), .ZN(n329) );
  OAI22_X1 U352 ( .A1(n340), .A2(n334), .B1(n219), .B2(n342), .ZN(n15) );
  XNOR2_X1 U353 ( .A(b[7]), .B(a[7]), .ZN(n342) );
  NAND2_X1 U354 ( .A1(n332), .A2(n351), .ZN(n334) );
  XNOR2_X1 U355 ( .A(n296), .B(a[6]), .ZN(n351) );
  XNOR2_X1 U356 ( .A(b[6]), .B(a[7]), .ZN(n340) );
  OAI22_X1 U357 ( .A1(n225), .A2(n307), .B1(n352), .B2(n305), .ZN(n104) );
  OAI22_X1 U358 ( .A1(n231), .A2(n307), .B1(n353), .B2(n305), .ZN(n103) );
  XNOR2_X1 U359 ( .A(b[1]), .B(a[1]), .ZN(n352) );
  OAI22_X1 U360 ( .A1(n353), .A2(n307), .B1(n354), .B2(n305), .ZN(n102) );
  XNOR2_X1 U361 ( .A(b[2]), .B(a[1]), .ZN(n353) );
  OAI22_X1 U362 ( .A1(n354), .A2(n307), .B1(n355), .B2(n305), .ZN(n101) );
  XNOR2_X1 U363 ( .A(b[3]), .B(a[1]), .ZN(n354) );
  OAI22_X1 U364 ( .A1(n355), .A2(n307), .B1(n306), .B2(n305), .ZN(n100) );
  XNOR2_X1 U365 ( .A(b[5]), .B(n224), .ZN(n306) );
  XNOR2_X1 U366 ( .A(b[4]), .B(n224), .ZN(n355) );
endmodule


module datapath_DW01_add_10 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n77;
  wire   [15:1] carry;

  FA_X1 U1_1 ( .A(A[1]), .B(n77), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(n64), .Z(n1) );
  CLKBUF_X1 U2 ( .A(carry[2]), .Z(n2) );
  CLKBUF_X1 U3 ( .A(n31), .Z(n3) );
  CLKBUF_X1 U4 ( .A(B[5]), .Z(n4) );
  XNOR2_X1 U5 ( .A(carry[14]), .B(n5), .ZN(SUM[14]) );
  XNOR2_X1 U6 ( .A(B[14]), .B(A[14]), .ZN(n5) );
  CLKBUF_X1 U7 ( .A(B[6]), .Z(n6) );
  NAND3_X1 U8 ( .A1(n20), .A2(n21), .A3(n22), .ZN(n7) );
  NAND3_X1 U9 ( .A1(n20), .A2(n21), .A3(n22), .ZN(n8) );
  CLKBUF_X1 U10 ( .A(B[3]), .Z(n9) );
  NAND3_X1 U11 ( .A1(n75), .A2(n74), .A3(n73), .ZN(n10) );
  NAND2_X1 U12 ( .A1(n10), .A2(B[14]), .ZN(n11) );
  NAND2_X1 U13 ( .A1(carry[14]), .A2(A[14]), .ZN(n12) );
  NAND2_X1 U14 ( .A1(B[14]), .A2(A[14]), .ZN(n13) );
  NAND3_X1 U15 ( .A1(n11), .A2(n12), .A3(n13), .ZN(carry[15]) );
  NAND3_X1 U16 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n14) );
  NAND3_X1 U17 ( .A1(n30), .A2(n3), .A3(n32), .ZN(n15) );
  NAND3_X1 U18 ( .A1(n36), .A2(n37), .A3(n38), .ZN(n16) );
  NAND3_X1 U19 ( .A1(n36), .A2(n37), .A3(n38), .ZN(n17) );
  NAND3_X1 U20 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n18) );
  XOR2_X1 U21 ( .A(n2), .B(A[2]), .Z(n19) );
  XOR2_X1 U22 ( .A(B[2]), .B(n19), .Z(SUM[2]) );
  NAND2_X1 U23 ( .A1(B[2]), .A2(carry[2]), .ZN(n20) );
  NAND2_X1 U24 ( .A1(B[2]), .A2(A[2]), .ZN(n21) );
  NAND2_X1 U25 ( .A1(carry[2]), .A2(A[2]), .ZN(n22) );
  NAND3_X1 U26 ( .A1(n20), .A2(n21), .A3(n22), .ZN(carry[3]) );
  NAND3_X1 U27 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n23) );
  XOR2_X1 U28 ( .A(B[7]), .B(A[7]), .Z(n24) );
  XOR2_X1 U29 ( .A(n17), .B(n24), .Z(SUM[7]) );
  NAND2_X1 U30 ( .A1(n16), .A2(B[7]), .ZN(n25) );
  NAND2_X1 U31 ( .A1(carry[7]), .A2(A[7]), .ZN(n26) );
  NAND2_X1 U32 ( .A1(B[7]), .A2(A[7]), .ZN(n27) );
  NAND3_X1 U33 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[8]) );
  NAND3_X1 U34 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n28) );
  XOR2_X1 U35 ( .A(n8), .B(A[3]), .Z(n29) );
  XOR2_X1 U36 ( .A(n9), .B(n29), .Z(SUM[3]) );
  NAND2_X1 U37 ( .A1(B[3]), .A2(n7), .ZN(n30) );
  NAND2_X1 U38 ( .A1(B[3]), .A2(A[3]), .ZN(n31) );
  NAND2_X1 U39 ( .A1(carry[3]), .A2(A[3]), .ZN(n32) );
  NAND3_X1 U40 ( .A1(n30), .A2(n31), .A3(n32), .ZN(carry[4]) );
  NAND3_X1 U41 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n33) );
  NAND3_X1 U42 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n34) );
  XOR2_X1 U43 ( .A(n6), .B(A[6]), .Z(n35) );
  XOR2_X1 U44 ( .A(n33), .B(n35), .Z(SUM[6]) );
  NAND2_X1 U45 ( .A1(n33), .A2(B[6]), .ZN(n36) );
  NAND2_X1 U46 ( .A1(carry[6]), .A2(A[6]), .ZN(n37) );
  NAND2_X1 U47 ( .A1(B[6]), .A2(A[6]), .ZN(n38) );
  NAND3_X1 U48 ( .A1(n36), .A2(n37), .A3(n38), .ZN(carry[7]) );
  NAND3_X1 U49 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n39) );
  NAND3_X1 U50 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n40) );
  XOR2_X1 U51 ( .A(B[11]), .B(A[11]), .Z(n41) );
  XOR2_X1 U52 ( .A(carry[11]), .B(n41), .Z(SUM[11]) );
  NAND2_X1 U53 ( .A1(n14), .A2(B[11]), .ZN(n42) );
  NAND2_X1 U54 ( .A1(n40), .A2(A[11]), .ZN(n43) );
  NAND2_X1 U55 ( .A1(B[11]), .A2(A[11]), .ZN(n44) );
  NAND3_X1 U56 ( .A1(n43), .A2(n42), .A3(n44), .ZN(carry[12]) );
  NAND3_X1 U57 ( .A1(n60), .A2(n61), .A3(n62), .ZN(n45) );
  XOR2_X1 U58 ( .A(B[8]), .B(A[8]), .Z(n46) );
  XOR2_X1 U59 ( .A(carry[8]), .B(n46), .Z(SUM[8]) );
  NAND2_X1 U60 ( .A1(n18), .A2(B[8]), .ZN(n47) );
  NAND2_X1 U61 ( .A1(n18), .A2(A[8]), .ZN(n48) );
  NAND2_X1 U62 ( .A1(B[8]), .A2(A[8]), .ZN(n49) );
  NAND3_X1 U63 ( .A1(n48), .A2(n47), .A3(n49), .ZN(carry[9]) );
  XOR2_X1 U64 ( .A(B[4]), .B(A[4]), .Z(n50) );
  XOR2_X1 U65 ( .A(n15), .B(n50), .Z(SUM[4]) );
  NAND2_X1 U66 ( .A1(carry[4]), .A2(B[4]), .ZN(n51) );
  NAND2_X1 U67 ( .A1(n28), .A2(A[4]), .ZN(n52) );
  NAND2_X1 U68 ( .A1(B[4]), .A2(A[4]), .ZN(n53) );
  NAND3_X1 U69 ( .A1(n52), .A2(n51), .A3(n53), .ZN(carry[5]) );
  XOR2_X1 U70 ( .A(n4), .B(A[5]), .Z(n54) );
  XOR2_X1 U71 ( .A(n23), .B(n54), .Z(SUM[5]) );
  NAND2_X1 U72 ( .A1(n23), .A2(B[5]), .ZN(n55) );
  NAND2_X1 U73 ( .A1(carry[5]), .A2(A[5]), .ZN(n56) );
  NAND2_X1 U74 ( .A1(B[5]), .A2(A[5]), .ZN(n57) );
  NAND3_X1 U75 ( .A1(n55), .A2(n56), .A3(n57), .ZN(carry[6]) );
  NAND3_X1 U76 ( .A1(n71), .A2(n69), .A3(n70), .ZN(n58) );
  XOR2_X1 U77 ( .A(B[9]), .B(A[9]), .Z(n59) );
  XOR2_X1 U78 ( .A(n34), .B(n59), .Z(SUM[9]) );
  NAND2_X1 U79 ( .A1(n34), .A2(B[9]), .ZN(n60) );
  NAND2_X1 U80 ( .A1(carry[9]), .A2(A[9]), .ZN(n61) );
  NAND2_X1 U81 ( .A1(B[9]), .A2(A[9]), .ZN(n62) );
  NAND3_X1 U82 ( .A1(n60), .A2(n61), .A3(n62), .ZN(carry[10]) );
  XOR2_X1 U83 ( .A(B[10]), .B(A[10]), .Z(n63) );
  XOR2_X1 U84 ( .A(n45), .B(n63), .Z(SUM[10]) );
  NAND2_X1 U85 ( .A1(n45), .A2(B[10]), .ZN(n64) );
  NAND2_X1 U86 ( .A1(carry[10]), .A2(A[10]), .ZN(n65) );
  NAND2_X1 U87 ( .A1(B[10]), .A2(A[10]), .ZN(n66) );
  NAND3_X1 U88 ( .A1(n1), .A2(n65), .A3(n66), .ZN(carry[11]) );
  NAND2_X1 U89 ( .A1(A[12]), .A2(B[12]), .ZN(n69) );
  XNOR2_X1 U90 ( .A(carry[15]), .B(n67), .ZN(SUM[15]) );
  XNOR2_X1 U91 ( .A(B[15]), .B(A[15]), .ZN(n67) );
  XOR2_X1 U92 ( .A(A[12]), .B(B[12]), .Z(n68) );
  XOR2_X1 U93 ( .A(n39), .B(n68), .Z(SUM[12]) );
  NAND2_X1 U94 ( .A1(A[12]), .A2(carry[12]), .ZN(n70) );
  NAND2_X1 U95 ( .A1(n39), .A2(B[12]), .ZN(n71) );
  NAND3_X1 U96 ( .A1(n71), .A2(n70), .A3(n69), .ZN(carry[13]) );
  XOR2_X1 U97 ( .A(A[13]), .B(B[13]), .Z(n72) );
  XOR2_X1 U98 ( .A(n72), .B(carry[13]), .Z(SUM[13]) );
  NAND2_X1 U99 ( .A1(A[13]), .A2(B[13]), .ZN(n73) );
  NAND2_X1 U100 ( .A1(A[13]), .A2(n58), .ZN(n74) );
  NAND2_X1 U101 ( .A1(carry[13]), .A2(B[13]), .ZN(n75) );
  NAND3_X1 U102 ( .A1(n75), .A2(n74), .A3(n73), .ZN(carry[14]) );
  XOR2_X1 U103 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U104 ( .A1(B[0]), .A2(A[0]), .ZN(n77) );
endmodule


module datapath_DW_mult_tc_9 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n210, n211, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362;

  FA_X1 U11 ( .A(n50), .B(n53), .CI(n11), .CO(n10), .S(product[5]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n306), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n305), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n309), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n308), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n311), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n92), .B(n80), .CI(n99), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  NAND3_X1 U157 ( .A1(n294), .A2(n295), .A3(n296), .ZN(n49) );
  INV_X1 U158 ( .A(n15), .ZN(n302) );
  CLKBUF_X1 U159 ( .A(b[1]), .Z(n206) );
  NAND3_X1 U160 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n207) );
  NAND3_X1 U161 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n208) );
  NAND3_X1 U162 ( .A1(n288), .A2(n289), .A3(n290), .ZN(n209) );
  CLKBUF_X1 U163 ( .A(n359), .Z(n234) );
  AND2_X1 U164 ( .A1(n95), .A2(n224), .ZN(n210) );
  AND2_X1 U165 ( .A1(n329), .A2(n357), .ZN(n211) );
  AND3_X1 U166 ( .A1(n227), .A2(n228), .A3(n229), .ZN(product[15]) );
  BUF_X1 U167 ( .A(a[1]), .Z(n220) );
  NAND3_X1 U168 ( .A1(n231), .A2(n232), .A3(n233), .ZN(n213) );
  NAND3_X1 U169 ( .A1(n231), .A2(n232), .A3(n233), .ZN(n214) );
  NAND3_X1 U170 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n215) );
  NAND3_X1 U171 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n216) );
  CLKBUF_X1 U172 ( .A(b[2]), .Z(n217) );
  INV_X1 U173 ( .A(n310), .ZN(n218) );
  INV_X1 U174 ( .A(n312), .ZN(n219) );
  NAND2_X2 U175 ( .A1(a[1]), .A2(n313), .ZN(n315) );
  BUF_X2 U176 ( .A(n339), .Z(n221) );
  XOR2_X1 U177 ( .A(a[6]), .B(n307), .Z(n339) );
  BUF_X1 U178 ( .A(n301), .Z(n222) );
  XNOR2_X1 U179 ( .A(n223), .B(n262), .ZN(product[4]) );
  XNOR2_X1 U180 ( .A(n54), .B(n210), .ZN(n223) );
  OAI22_X1 U181 ( .A1(n360), .A2(n315), .B1(n361), .B2(n313), .ZN(n224) );
  CLKBUF_X1 U182 ( .A(n329), .Z(n225) );
  XNOR2_X1 U183 ( .A(a[4]), .B(a[3]), .ZN(n329) );
  XOR2_X1 U184 ( .A(n303), .B(n15), .Z(n226) );
  XOR2_X1 U185 ( .A(n2), .B(n226), .Z(product[14]) );
  NAND2_X1 U186 ( .A1(n209), .A2(n303), .ZN(n227) );
  NAND2_X1 U187 ( .A1(n209), .A2(n15), .ZN(n228) );
  NAND2_X1 U188 ( .A1(n303), .A2(n15), .ZN(n229) );
  XOR2_X1 U189 ( .A(n23), .B(n20), .Z(n230) );
  XOR2_X1 U190 ( .A(n5), .B(n230), .Z(product[11]) );
  NAND2_X1 U191 ( .A1(n208), .A2(n23), .ZN(n231) );
  NAND2_X1 U192 ( .A1(n207), .A2(n20), .ZN(n232) );
  NAND2_X1 U193 ( .A1(n23), .A2(n20), .ZN(n233) );
  NAND3_X1 U194 ( .A1(n231), .A2(n232), .A3(n233), .ZN(n4) );
  INV_X1 U195 ( .A(n211), .ZN(n235) );
  INV_X1 U196 ( .A(n211), .ZN(n236) );
  NAND2_X1 U197 ( .A1(n14), .A2(n96), .ZN(n237) );
  AND2_X1 U198 ( .A1(n104), .A2(n72), .ZN(n238) );
  OAI22_X1 U199 ( .A1(n320), .A2(n321), .B1(n298), .B2(n322), .ZN(n239) );
  XOR2_X1 U200 ( .A(n46), .B(n49), .Z(n240) );
  XOR2_X1 U201 ( .A(n10), .B(n240), .Z(product[6]) );
  NAND2_X1 U202 ( .A1(n10), .A2(n46), .ZN(n241) );
  NAND2_X1 U203 ( .A1(n10), .A2(n49), .ZN(n242) );
  NAND2_X1 U204 ( .A1(n46), .A2(n49), .ZN(n243) );
  NAND3_X1 U205 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n9) );
  XOR2_X1 U206 ( .A(a[3]), .B(n301), .Z(n320) );
  XOR2_X1 U207 ( .A(n95), .B(n224), .Z(n244) );
  XNOR2_X1 U208 ( .A(n238), .B(n245), .ZN(product[2]) );
  XNOR2_X1 U209 ( .A(n103), .B(n96), .ZN(n245) );
  NAND3_X1 U210 ( .A1(n275), .A2(n276), .A3(n277), .ZN(n246) );
  NAND3_X1 U211 ( .A1(n275), .A2(n276), .A3(n277), .ZN(n247) );
  NAND3_X1 U212 ( .A1(n254), .A2(n253), .A3(n255), .ZN(n248) );
  NAND3_X1 U213 ( .A1(n237), .A2(n256), .A3(n258), .ZN(n249) );
  NAND3_X1 U214 ( .A1(n256), .A2(n237), .A3(n258), .ZN(n250) );
  OAI22_X1 U215 ( .A1(n234), .A2(n315), .B1(n360), .B2(n313), .ZN(n251) );
  XOR2_X1 U216 ( .A(n33), .B(n28), .Z(n252) );
  XOR2_X1 U217 ( .A(n247), .B(n252), .Z(product[9]) );
  NAND2_X1 U218 ( .A1(n246), .A2(n33), .ZN(n253) );
  NAND2_X1 U219 ( .A1(n246), .A2(n28), .ZN(n254) );
  NAND2_X1 U220 ( .A1(n33), .A2(n28), .ZN(n255) );
  NAND3_X1 U221 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n6) );
  NAND2_X1 U222 ( .A1(n238), .A2(n251), .ZN(n256) );
  NAND2_X1 U223 ( .A1(n14), .A2(n96), .ZN(n257) );
  NAND2_X1 U224 ( .A1(n251), .A2(n96), .ZN(n258) );
  NAND3_X1 U225 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n13) );
  CLKBUF_X1 U226 ( .A(b[1]), .Z(n259) );
  NAND3_X1 U227 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n260) );
  NAND3_X1 U228 ( .A1(n266), .A2(n265), .A3(n264), .ZN(n261) );
  NAND3_X1 U229 ( .A1(n265), .A2(n264), .A3(n266), .ZN(n262) );
  XNOR2_X1 U230 ( .A(n263), .B(n250), .ZN(product[3]) );
  XNOR2_X1 U231 ( .A(n244), .B(n71), .ZN(n263) );
  NAND2_X1 U232 ( .A1(n56), .A2(n71), .ZN(n264) );
  NAND2_X1 U233 ( .A1(n249), .A2(n56), .ZN(n265) );
  NAND2_X1 U234 ( .A1(n13), .A2(n71), .ZN(n266) );
  NAND3_X1 U235 ( .A1(n266), .A2(n265), .A3(n264), .ZN(n12) );
  NAND2_X1 U236 ( .A1(n54), .A2(n210), .ZN(n267) );
  NAND2_X1 U237 ( .A1(n261), .A2(n54), .ZN(n268) );
  NAND2_X1 U238 ( .A1(n12), .A2(n210), .ZN(n269) );
  NAND3_X1 U239 ( .A1(n268), .A2(n269), .A3(n267), .ZN(n11) );
  XOR2_X1 U240 ( .A(n40), .B(n45), .Z(n270) );
  XOR2_X1 U241 ( .A(n216), .B(n270), .Z(product[7]) );
  NAND2_X1 U242 ( .A1(n215), .A2(n40), .ZN(n271) );
  NAND2_X1 U243 ( .A1(n9), .A2(n45), .ZN(n272) );
  NAND2_X1 U244 ( .A1(n40), .A2(n45), .ZN(n273) );
  NAND3_X1 U245 ( .A1(n272), .A2(n271), .A3(n273), .ZN(n8) );
  XOR2_X1 U246 ( .A(n34), .B(n39), .Z(n274) );
  XOR2_X1 U247 ( .A(n260), .B(n274), .Z(product[8]) );
  NAND2_X1 U248 ( .A1(n260), .A2(n34), .ZN(n275) );
  NAND2_X1 U249 ( .A1(n8), .A2(n39), .ZN(n276) );
  NAND2_X1 U250 ( .A1(n34), .A2(n39), .ZN(n277) );
  XOR2_X1 U251 ( .A(n27), .B(n24), .Z(n278) );
  XOR2_X1 U252 ( .A(n248), .B(n278), .Z(product[10]) );
  NAND2_X1 U253 ( .A1(n248), .A2(n27), .ZN(n279) );
  NAND2_X1 U254 ( .A1(n6), .A2(n24), .ZN(n280) );
  NAND2_X1 U255 ( .A1(n27), .A2(n24), .ZN(n281) );
  NAND3_X1 U256 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n5) );
  NAND3_X1 U257 ( .A1(n284), .A2(n285), .A3(n286), .ZN(n282) );
  XOR2_X1 U258 ( .A(n239), .B(n102), .Z(n56) );
  XOR2_X1 U259 ( .A(n18), .B(n19), .Z(n283) );
  XOR2_X1 U260 ( .A(n214), .B(n283), .Z(product[12]) );
  NAND2_X1 U261 ( .A1(n213), .A2(n18), .ZN(n284) );
  NAND2_X1 U262 ( .A1(n4), .A2(n19), .ZN(n285) );
  NAND2_X1 U263 ( .A1(n18), .A2(n19), .ZN(n286) );
  NAND3_X1 U264 ( .A1(n285), .A2(n284), .A3(n286), .ZN(n3) );
  XOR2_X1 U265 ( .A(n17), .B(n302), .Z(n287) );
  XOR2_X1 U266 ( .A(n3), .B(n287), .Z(product[13]) );
  NAND2_X1 U267 ( .A1(n282), .A2(n17), .ZN(n288) );
  NAND2_X1 U268 ( .A1(n282), .A2(n302), .ZN(n289) );
  NAND2_X1 U269 ( .A1(n17), .A2(n302), .ZN(n290) );
  NAND3_X1 U270 ( .A1(n288), .A2(n289), .A3(n290), .ZN(n2) );
  NAND2_X1 U271 ( .A1(n297), .A2(n356), .ZN(n291) );
  INV_X1 U272 ( .A(n301), .ZN(n292) );
  XNOR2_X1 U273 ( .A(n52), .B(n293), .ZN(n50) );
  XNOR2_X1 U274 ( .A(n93), .B(n100), .ZN(n293) );
  INV_X1 U275 ( .A(n327), .ZN(n309) );
  INV_X1 U276 ( .A(n31), .ZN(n308) );
  INV_X1 U277 ( .A(n21), .ZN(n305) );
  INV_X1 U278 ( .A(n337), .ZN(n306) );
  INV_X1 U279 ( .A(n348), .ZN(n303) );
  INV_X1 U280 ( .A(n318), .ZN(n311) );
  CLKBUF_X1 U281 ( .A(n319), .Z(n299) );
  NAND2_X1 U282 ( .A1(n297), .A2(n356), .ZN(n321) );
  INV_X1 U283 ( .A(a[5]), .ZN(n307) );
  INV_X1 U284 ( .A(a[7]), .ZN(n304) );
  INV_X1 U285 ( .A(b[0]), .ZN(n301) );
  NAND2_X1 U286 ( .A1(n52), .A2(n93), .ZN(n294) );
  NAND2_X1 U287 ( .A1(n52), .A2(n100), .ZN(n295) );
  NAND2_X1 U288 ( .A1(n93), .A2(n100), .ZN(n296) );
  BUF_X1 U289 ( .A(n319), .Z(n297) );
  BUF_X1 U290 ( .A(n319), .Z(n298) );
  XNOR2_X1 U291 ( .A(a[2]), .B(a[1]), .ZN(n319) );
  INV_X1 U292 ( .A(a[3]), .ZN(n310) );
  INV_X1 U293 ( .A(a[1]), .ZN(n312) );
  INV_X1 U294 ( .A(n301), .ZN(n300) );
  INV_X2 U295 ( .A(a[0]), .ZN(n313) );
  NOR2_X1 U296 ( .A1(n313), .A2(n222), .ZN(product[0]) );
  OAI22_X1 U297 ( .A1(n314), .A2(n315), .B1(n316), .B2(n313), .ZN(n99) );
  OAI22_X1 U298 ( .A1(n316), .A2(n315), .B1(n317), .B2(n313), .ZN(n98) );
  XNOR2_X1 U299 ( .A(b[6]), .B(n220), .ZN(n316) );
  OAI22_X1 U300 ( .A1(n313), .A2(n317), .B1(n315), .B2(n317), .ZN(n318) );
  XNOR2_X1 U301 ( .A(b[7]), .B(n219), .ZN(n317) );
  NOR2_X1 U302 ( .A1(n299), .A2(n222), .ZN(n96) );
  OAI22_X1 U303 ( .A1(n320), .A2(n321), .B1(n298), .B2(n322), .ZN(n95) );
  OAI22_X1 U304 ( .A1(n322), .A2(n291), .B1(n298), .B2(n323), .ZN(n94) );
  XNOR2_X1 U305 ( .A(n206), .B(a[3]), .ZN(n322) );
  OAI22_X1 U306 ( .A1(n323), .A2(n321), .B1(n298), .B2(n324), .ZN(n93) );
  XNOR2_X1 U307 ( .A(b[2]), .B(a[3]), .ZN(n323) );
  OAI22_X1 U308 ( .A1(n324), .A2(n291), .B1(n299), .B2(n325), .ZN(n92) );
  XNOR2_X1 U309 ( .A(b[3]), .B(n218), .ZN(n324) );
  OAI22_X1 U310 ( .A1(n325), .A2(n291), .B1(n299), .B2(n326), .ZN(n91) );
  XNOR2_X1 U311 ( .A(b[4]), .B(n218), .ZN(n325) );
  OAI22_X1 U312 ( .A1(n328), .A2(n298), .B1(n321), .B2(n328), .ZN(n327) );
  NOR2_X1 U313 ( .A1(n329), .A2(n222), .ZN(n88) );
  OAI22_X1 U314 ( .A1(n330), .A2(n235), .B1(n329), .B2(n331), .ZN(n87) );
  XNOR2_X1 U315 ( .A(a[5]), .B(n292), .ZN(n330) );
  OAI22_X1 U316 ( .A1(n331), .A2(n236), .B1(n329), .B2(n332), .ZN(n86) );
  XNOR2_X1 U317 ( .A(n259), .B(a[5]), .ZN(n331) );
  OAI22_X1 U318 ( .A1(n332), .A2(n236), .B1(n329), .B2(n333), .ZN(n85) );
  XNOR2_X1 U319 ( .A(n217), .B(a[5]), .ZN(n332) );
  OAI22_X1 U320 ( .A1(n333), .A2(n236), .B1(n225), .B2(n334), .ZN(n84) );
  XNOR2_X1 U321 ( .A(b[3]), .B(a[5]), .ZN(n333) );
  OAI22_X1 U322 ( .A1(n334), .A2(n236), .B1(n225), .B2(n335), .ZN(n83) );
  XNOR2_X1 U323 ( .A(b[4]), .B(a[5]), .ZN(n334) );
  OAI22_X1 U324 ( .A1(n335), .A2(n236), .B1(n225), .B2(n336), .ZN(n82) );
  XNOR2_X1 U325 ( .A(b[5]), .B(a[5]), .ZN(n335) );
  OAI22_X1 U326 ( .A1(n338), .A2(n225), .B1(n236), .B2(n338), .ZN(n337) );
  NOR2_X1 U327 ( .A1(n339), .A2(n222), .ZN(n80) );
  OAI22_X1 U328 ( .A1(n340), .A2(n341), .B1(n221), .B2(n342), .ZN(n79) );
  XNOR2_X1 U329 ( .A(a[7]), .B(n292), .ZN(n340) );
  OAI22_X1 U330 ( .A1(n343), .A2(n341), .B1(n221), .B2(n344), .ZN(n77) );
  OAI22_X1 U331 ( .A1(n344), .A2(n341), .B1(n221), .B2(n345), .ZN(n76) );
  XNOR2_X1 U332 ( .A(b[3]), .B(a[7]), .ZN(n344) );
  OAI22_X1 U333 ( .A1(n345), .A2(n341), .B1(n221), .B2(n346), .ZN(n75) );
  XNOR2_X1 U334 ( .A(b[4]), .B(a[7]), .ZN(n345) );
  OAI22_X1 U335 ( .A1(n346), .A2(n341), .B1(n221), .B2(n347), .ZN(n74) );
  XNOR2_X1 U336 ( .A(b[5]), .B(a[7]), .ZN(n346) );
  OAI22_X1 U337 ( .A1(n349), .A2(n221), .B1(n341), .B2(n349), .ZN(n348) );
  OAI21_X1 U338 ( .B1(n300), .B2(n312), .A(n315), .ZN(n72) );
  OAI21_X1 U339 ( .B1(n310), .B2(n321), .A(n350), .ZN(n71) );
  OR3_X1 U340 ( .A1(n299), .A2(n292), .A3(n310), .ZN(n350) );
  OAI21_X1 U341 ( .B1(n307), .B2(n235), .A(n351), .ZN(n70) );
  OR3_X1 U342 ( .A1(n329), .A2(n292), .A3(n307), .ZN(n351) );
  OAI21_X1 U343 ( .B1(n304), .B2(n341), .A(n352), .ZN(n69) );
  OR3_X1 U344 ( .A1(n339), .A2(n292), .A3(n304), .ZN(n352) );
  XNOR2_X1 U345 ( .A(n353), .B(n354), .ZN(n38) );
  OR2_X1 U346 ( .A1(n353), .A2(n354), .ZN(n37) );
  OAI22_X1 U347 ( .A1(n326), .A2(n321), .B1(n299), .B2(n355), .ZN(n354) );
  XNOR2_X1 U348 ( .A(b[5]), .B(n218), .ZN(n326) );
  OAI22_X1 U349 ( .A1(n342), .A2(n341), .B1(n221), .B2(n343), .ZN(n353) );
  XNOR2_X1 U350 ( .A(n217), .B(a[7]), .ZN(n343) );
  XNOR2_X1 U351 ( .A(n259), .B(a[7]), .ZN(n342) );
  OAI22_X1 U352 ( .A1(n355), .A2(n291), .B1(n298), .B2(n328), .ZN(n31) );
  XNOR2_X1 U353 ( .A(b[7]), .B(n218), .ZN(n328) );
  XNOR2_X1 U354 ( .A(n310), .B(a[2]), .ZN(n356) );
  XNOR2_X1 U355 ( .A(b[6]), .B(n218), .ZN(n355) );
  OAI22_X1 U356 ( .A1(n336), .A2(n236), .B1(n225), .B2(n338), .ZN(n21) );
  XNOR2_X1 U357 ( .A(b[7]), .B(a[5]), .ZN(n338) );
  XNOR2_X1 U358 ( .A(n307), .B(a[4]), .ZN(n357) );
  XNOR2_X1 U359 ( .A(b[6]), .B(a[5]), .ZN(n336) );
  OAI22_X1 U360 ( .A1(n347), .A2(n341), .B1(n221), .B2(n349), .ZN(n15) );
  XNOR2_X1 U361 ( .A(b[7]), .B(a[7]), .ZN(n349) );
  NAND2_X1 U362 ( .A1(n339), .A2(n358), .ZN(n341) );
  XNOR2_X1 U363 ( .A(n304), .B(a[6]), .ZN(n358) );
  XNOR2_X1 U364 ( .A(b[6]), .B(a[7]), .ZN(n347) );
  OAI22_X1 U365 ( .A1(n300), .A2(n315), .B1(n359), .B2(n313), .ZN(n104) );
  OAI22_X1 U366 ( .A1(n234), .A2(n315), .B1(n360), .B2(n313), .ZN(n103) );
  XNOR2_X1 U367 ( .A(b[1]), .B(a[1]), .ZN(n359) );
  OAI22_X1 U368 ( .A1(n360), .A2(n315), .B1(n361), .B2(n313), .ZN(n102) );
  XNOR2_X1 U369 ( .A(b[2]), .B(n220), .ZN(n360) );
  OAI22_X1 U370 ( .A1(n361), .A2(n315), .B1(n362), .B2(n313), .ZN(n101) );
  XNOR2_X1 U371 ( .A(b[3]), .B(n220), .ZN(n361) );
  OAI22_X1 U372 ( .A1(n362), .A2(n315), .B1(n314), .B2(n313), .ZN(n100) );
  XNOR2_X1 U373 ( .A(b[5]), .B(n219), .ZN(n314) );
  XNOR2_X1 U374 ( .A(b[4]), .B(n220), .ZN(n362) );
endmodule


module datapath_DW01_add_9 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n82;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n82), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(n65), .Z(n1) );
  CLKBUF_X1 U2 ( .A(n64), .Z(n2) );
  CLKBUF_X1 U3 ( .A(n13), .Z(n3) );
  NAND3_X1 U4 ( .A1(n2), .A2(n1), .A3(n66), .ZN(n4) );
  CLKBUF_X1 U5 ( .A(n22), .Z(n5) );
  CLKBUF_X1 U6 ( .A(n59), .Z(n6) );
  CLKBUF_X1 U7 ( .A(carry[2]), .Z(n7) );
  NAND3_X1 U8 ( .A1(n11), .A2(n12), .A3(n13), .ZN(n8) );
  NAND3_X1 U9 ( .A1(n11), .A2(n12), .A3(n3), .ZN(n9) );
  XOR2_X1 U10 ( .A(n7), .B(A[2]), .Z(n10) );
  XOR2_X1 U11 ( .A(B[2]), .B(n10), .Z(SUM[2]) );
  NAND2_X1 U12 ( .A1(carry[2]), .A2(B[2]), .ZN(n11) );
  NAND2_X1 U13 ( .A1(B[2]), .A2(A[2]), .ZN(n12) );
  NAND2_X1 U14 ( .A1(carry[2]), .A2(A[2]), .ZN(n13) );
  NAND3_X1 U15 ( .A1(n11), .A2(n12), .A3(n13), .ZN(carry[3]) );
  NAND3_X1 U16 ( .A1(n76), .A2(n75), .A3(n74), .ZN(n14) );
  NAND3_X1 U17 ( .A1(n18), .A2(n17), .A3(n19), .ZN(n15) );
  XOR2_X1 U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  XOR2_X1 U19 ( .A(n9), .B(n16), .Z(SUM[3]) );
  NAND2_X1 U20 ( .A1(n8), .A2(B[3]), .ZN(n17) );
  NAND2_X1 U21 ( .A1(carry[3]), .A2(A[3]), .ZN(n18) );
  NAND2_X1 U22 ( .A1(B[3]), .A2(A[3]), .ZN(n19) );
  NAND3_X1 U23 ( .A1(n17), .A2(n18), .A3(n19), .ZN(carry[4]) );
  NAND3_X1 U24 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n20) );
  NAND2_X1 U25 ( .A1(carry[9]), .A2(A[9]), .ZN(n21) );
  NAND3_X1 U26 ( .A1(n40), .A2(n41), .A3(n42), .ZN(n22) );
  NAND3_X1 U27 ( .A1(n70), .A2(n69), .A3(n71), .ZN(n23) );
  CLKBUF_X1 U28 ( .A(n51), .Z(n24) );
  XOR2_X1 U29 ( .A(B[6]), .B(A[6]), .Z(n25) );
  XOR2_X1 U30 ( .A(n5), .B(n25), .Z(SUM[6]) );
  NAND2_X1 U31 ( .A1(n22), .A2(B[6]), .ZN(n26) );
  NAND2_X1 U32 ( .A1(carry[6]), .A2(A[6]), .ZN(n27) );
  NAND2_X1 U33 ( .A1(B[6]), .A2(A[6]), .ZN(n28) );
  NAND3_X1 U34 ( .A1(n26), .A2(n27), .A3(n28), .ZN(carry[7]) );
  NAND3_X1 U35 ( .A1(n76), .A2(n75), .A3(n74), .ZN(n29) );
  NAND3_X1 U36 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n30) );
  NAND3_X1 U37 ( .A1(n35), .A2(n36), .A3(n37), .ZN(n31) );
  NAND3_X1 U38 ( .A1(n50), .A2(n51), .A3(n52), .ZN(n32) );
  NAND3_X1 U39 ( .A1(n50), .A2(n24), .A3(n52), .ZN(n33) );
  XOR2_X1 U40 ( .A(B[4]), .B(A[4]), .Z(n34) );
  XOR2_X1 U41 ( .A(n15), .B(n34), .Z(SUM[4]) );
  NAND2_X1 U42 ( .A1(n15), .A2(B[4]), .ZN(n35) );
  NAND2_X1 U43 ( .A1(carry[4]), .A2(A[4]), .ZN(n36) );
  NAND2_X1 U44 ( .A1(B[4]), .A2(A[4]), .ZN(n37) );
  NAND3_X1 U45 ( .A1(n35), .A2(n36), .A3(n37), .ZN(carry[5]) );
  CLKBUF_X1 U46 ( .A(n75), .Z(n38) );
  XOR2_X1 U47 ( .A(B[5]), .B(A[5]), .Z(n39) );
  XOR2_X1 U48 ( .A(carry[5]), .B(n39), .Z(SUM[5]) );
  NAND2_X1 U49 ( .A1(n31), .A2(B[5]), .ZN(n40) );
  NAND2_X1 U50 ( .A1(n31), .A2(A[5]), .ZN(n41) );
  NAND2_X1 U51 ( .A1(B[5]), .A2(A[5]), .ZN(n42) );
  NAND3_X1 U52 ( .A1(n41), .A2(n40), .A3(n42), .ZN(carry[6]) );
  CLKBUF_X1 U53 ( .A(n69), .Z(n43) );
  CLKBUF_X1 U54 ( .A(n21), .Z(n44) );
  XOR2_X1 U55 ( .A(B[7]), .B(A[7]), .Z(n45) );
  XOR2_X1 U56 ( .A(carry[7]), .B(n45), .Z(SUM[7]) );
  NAND2_X1 U57 ( .A1(n20), .A2(B[7]), .ZN(n46) );
  NAND2_X1 U58 ( .A1(n20), .A2(A[7]), .ZN(n47) );
  NAND2_X1 U59 ( .A1(B[7]), .A2(A[7]), .ZN(n48) );
  NAND3_X1 U60 ( .A1(n46), .A2(n47), .A3(n48), .ZN(carry[8]) );
  XOR2_X1 U61 ( .A(B[8]), .B(A[8]), .Z(n49) );
  XOR2_X1 U62 ( .A(carry[8]), .B(n49), .Z(SUM[8]) );
  NAND2_X1 U63 ( .A1(n30), .A2(B[8]), .ZN(n50) );
  NAND2_X1 U64 ( .A1(n30), .A2(A[8]), .ZN(n51) );
  NAND2_X1 U65 ( .A1(B[8]), .A2(A[8]), .ZN(n52) );
  NAND3_X1 U66 ( .A1(n50), .A2(n51), .A3(n52), .ZN(carry[9]) );
  CLKBUF_X1 U67 ( .A(n70), .Z(n53) );
  NAND3_X1 U68 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n54) );
  NAND3_X1 U69 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n55) );
  NAND3_X1 U70 ( .A1(n59), .A2(n21), .A3(n61), .ZN(n56) );
  NAND3_X1 U71 ( .A1(n6), .A2(n44), .A3(n61), .ZN(n57) );
  XOR2_X1 U72 ( .A(B[9]), .B(A[9]), .Z(n58) );
  XOR2_X1 U73 ( .A(n33), .B(n58), .Z(SUM[9]) );
  NAND2_X1 U74 ( .A1(n32), .A2(B[9]), .ZN(n59) );
  NAND2_X1 U75 ( .A1(carry[9]), .A2(A[9]), .ZN(n60) );
  NAND2_X1 U76 ( .A1(B[9]), .A2(A[9]), .ZN(n61) );
  NAND3_X1 U77 ( .A1(n59), .A2(n60), .A3(n61), .ZN(carry[10]) );
  NAND3_X1 U78 ( .A1(n76), .A2(n38), .A3(n74), .ZN(n62) );
  XOR2_X1 U79 ( .A(B[10]), .B(A[10]), .Z(n63) );
  XOR2_X1 U80 ( .A(n57), .B(n63), .Z(SUM[10]) );
  NAND2_X1 U81 ( .A1(n56), .A2(B[10]), .ZN(n64) );
  NAND2_X1 U82 ( .A1(carry[10]), .A2(A[10]), .ZN(n65) );
  NAND2_X1 U83 ( .A1(B[10]), .A2(A[10]), .ZN(n66) );
  NAND3_X1 U84 ( .A1(n43), .A2(n53), .A3(n71), .ZN(n67) );
  XOR2_X1 U85 ( .A(B[11]), .B(A[11]), .Z(n68) );
  XOR2_X1 U86 ( .A(n4), .B(n68), .Z(SUM[11]) );
  NAND2_X1 U87 ( .A1(n54), .A2(B[11]), .ZN(n69) );
  NAND2_X1 U88 ( .A1(n55), .A2(A[11]), .ZN(n70) );
  NAND2_X1 U89 ( .A1(B[11]), .A2(A[11]), .ZN(n71) );
  NAND3_X1 U90 ( .A1(n69), .A2(n70), .A3(n71), .ZN(carry[12]) );
  XNOR2_X1 U91 ( .A(carry[15]), .B(n72), .ZN(SUM[15]) );
  XNOR2_X1 U92 ( .A(B[15]), .B(A[15]), .ZN(n72) );
  XOR2_X1 U93 ( .A(A[12]), .B(B[12]), .Z(n73) );
  XOR2_X1 U94 ( .A(n73), .B(n67), .Z(SUM[12]) );
  NAND2_X1 U95 ( .A1(A[12]), .A2(B[12]), .ZN(n74) );
  NAND2_X1 U96 ( .A1(A[12]), .A2(carry[12]), .ZN(n75) );
  NAND2_X1 U97 ( .A1(B[12]), .A2(n23), .ZN(n76) );
  XOR2_X1 U98 ( .A(A[13]), .B(B[13]), .Z(n77) );
  XOR2_X1 U99 ( .A(n77), .B(n62), .Z(SUM[13]) );
  NAND2_X1 U100 ( .A1(A[13]), .A2(B[13]), .ZN(n78) );
  NAND2_X1 U101 ( .A1(n29), .A2(A[13]), .ZN(n79) );
  NAND2_X1 U102 ( .A1(B[13]), .A2(n14), .ZN(n80) );
  NAND3_X1 U103 ( .A1(n80), .A2(n79), .A3(n78), .ZN(carry[14]) );
  XOR2_X1 U104 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U105 ( .A1(B[0]), .A2(A[0]), .ZN(n82) );
endmodule


module datapath_DW_mult_tc_8 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343;

  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n286), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n285), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n289), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n288), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n291), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  BUF_X1 U157 ( .A(n301), .Z(n209) );
  INV_X1 U158 ( .A(n15), .ZN(n282) );
  NAND2_X2 U159 ( .A1(n227), .A2(n293), .ZN(n295) );
  AND2_X1 U160 ( .A1(n95), .A2(n102), .ZN(n206) );
  XNOR2_X1 U161 ( .A(n283), .B(n15), .ZN(n207) );
  AND3_X1 U162 ( .A1(n255), .A2(n256), .A3(n257), .ZN(product[15]) );
  CLKBUF_X1 U163 ( .A(n12), .Z(n242) );
  XOR2_X1 U164 ( .A(n210), .B(n211), .Z(product[11]) );
  XNOR2_X1 U165 ( .A(n20), .B(n23), .ZN(n210) );
  AND3_X1 U166 ( .A1(n263), .A2(n264), .A3(n265), .ZN(n211) );
  XNOR2_X1 U167 ( .A(n249), .B(n212), .ZN(product[10]) );
  XNOR2_X1 U168 ( .A(n27), .B(n24), .ZN(n212) );
  XNOR2_X1 U169 ( .A(n213), .B(n234), .ZN(product[13]) );
  AND3_X1 U170 ( .A1(n270), .A2(n271), .A3(n272), .ZN(n213) );
  XNOR2_X1 U171 ( .A(n269), .B(n214), .ZN(product[12]) );
  AND3_X1 U172 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n214) );
  CLKBUF_X1 U173 ( .A(n320), .Z(n215) );
  XOR2_X1 U174 ( .A(a[6]), .B(n287), .Z(n320) );
  XNOR2_X1 U175 ( .A(n216), .B(n233), .ZN(product[5]) );
  XNOR2_X1 U176 ( .A(n50), .B(n53), .ZN(n216) );
  NAND3_X1 U177 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n217) );
  NAND3_X1 U178 ( .A1(n248), .A2(n247), .A3(n246), .ZN(n218) );
  NAND3_X1 U179 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n219) );
  NAND3_X1 U180 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n220) );
  XNOR2_X1 U181 ( .A(n221), .B(n242), .ZN(product[4]) );
  XNOR2_X1 U182 ( .A(n54), .B(n206), .ZN(n221) );
  NAND3_X1 U183 ( .A1(n261), .A2(n262), .A3(n260), .ZN(n222) );
  XOR2_X1 U184 ( .A(n46), .B(n49), .Z(n223) );
  XOR2_X1 U185 ( .A(n218), .B(n223), .Z(product[6]) );
  NAND2_X1 U186 ( .A1(n218), .A2(n46), .ZN(n224) );
  NAND2_X1 U187 ( .A1(n10), .A2(n49), .ZN(n225) );
  NAND2_X1 U188 ( .A1(n46), .A2(n49), .ZN(n226) );
  NAND3_X1 U189 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n9) );
  CLKBUF_X1 U190 ( .A(a[1]), .Z(n227) );
  NAND3_X1 U191 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n228) );
  NAND3_X1 U192 ( .A1(n270), .A2(n271), .A3(n272), .ZN(n229) );
  NAND3_X1 U193 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n230) );
  NAND3_X1 U194 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n231) );
  NAND3_X1 U195 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n232) );
  NAND3_X1 U196 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n233) );
  XOR2_X1 U197 ( .A(n17), .B(n282), .Z(n234) );
  NAND2_X1 U198 ( .A1(n229), .A2(n17), .ZN(n235) );
  NAND2_X1 U199 ( .A1(n3), .A2(n282), .ZN(n236) );
  NAND2_X1 U200 ( .A1(n17), .A2(n282), .ZN(n237) );
  NAND3_X1 U201 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n2) );
  XOR2_X1 U202 ( .A(n40), .B(n45), .Z(n238) );
  XOR2_X1 U203 ( .A(n220), .B(n238), .Z(product[7]) );
  NAND2_X1 U204 ( .A1(n219), .A2(n40), .ZN(n239) );
  NAND2_X1 U205 ( .A1(n9), .A2(n45), .ZN(n240) );
  NAND2_X1 U206 ( .A1(n40), .A2(n45), .ZN(n241) );
  NAND2_X1 U207 ( .A1(n54), .A2(n206), .ZN(n243) );
  NAND2_X1 U208 ( .A1(n54), .A2(n12), .ZN(n244) );
  NAND2_X1 U209 ( .A1(n206), .A2(n12), .ZN(n245) );
  NAND3_X1 U210 ( .A1(n245), .A2(n244), .A3(n243), .ZN(n11) );
  NAND2_X1 U211 ( .A1(n50), .A2(n53), .ZN(n246) );
  NAND2_X1 U212 ( .A1(n232), .A2(n50), .ZN(n247) );
  NAND2_X1 U213 ( .A1(n53), .A2(n11), .ZN(n248) );
  NAND3_X1 U214 ( .A1(n248), .A2(n247), .A3(n246), .ZN(n10) );
  XOR2_X1 U215 ( .A(a[3]), .B(n281), .Z(n300) );
  NAND3_X1 U216 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n249) );
  XNOR2_X1 U217 ( .A(n2), .B(n207), .ZN(product[14]) );
  XOR2_X1 U218 ( .A(n33), .B(n28), .Z(n250) );
  XOR2_X1 U219 ( .A(n222), .B(n250), .Z(product[9]) );
  NAND2_X1 U220 ( .A1(n228), .A2(n33), .ZN(n251) );
  NAND2_X1 U221 ( .A1(n7), .A2(n28), .ZN(n252) );
  NAND2_X1 U222 ( .A1(n33), .A2(n28), .ZN(n253) );
  NAND3_X1 U223 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n6) );
  CLKBUF_X1 U224 ( .A(n340), .Z(n254) );
  NAND2_X1 U225 ( .A1(n217), .A2(n283), .ZN(n255) );
  NAND2_X1 U226 ( .A1(n217), .A2(n15), .ZN(n256) );
  NAND2_X1 U227 ( .A1(n283), .A2(n15), .ZN(n257) );
  NAND3_X1 U228 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n258) );
  XOR2_X1 U229 ( .A(n34), .B(n39), .Z(n259) );
  XOR2_X1 U230 ( .A(n230), .B(n259), .Z(product[8]) );
  NAND2_X1 U231 ( .A1(n231), .A2(n34), .ZN(n260) );
  NAND2_X1 U232 ( .A1(n231), .A2(n39), .ZN(n261) );
  NAND2_X1 U233 ( .A1(n34), .A2(n39), .ZN(n262) );
  NAND3_X1 U234 ( .A1(n261), .A2(n260), .A3(n262), .ZN(n7) );
  NAND2_X1 U235 ( .A1(n249), .A2(n27), .ZN(n263) );
  NAND2_X1 U236 ( .A1(n6), .A2(n24), .ZN(n264) );
  NAND2_X1 U237 ( .A1(n27), .A2(n24), .ZN(n265) );
  NAND3_X1 U238 ( .A1(n263), .A2(n264), .A3(n265), .ZN(n5) );
  BUF_X2 U239 ( .A(a[1]), .Z(n275) );
  NAND2_X1 U240 ( .A1(n20), .A2(n23), .ZN(n266) );
  NAND2_X1 U241 ( .A1(n5), .A2(n20), .ZN(n267) );
  NAND2_X1 U242 ( .A1(n5), .A2(n23), .ZN(n268) );
  NAND3_X1 U243 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n4) );
  XOR2_X1 U244 ( .A(n19), .B(n18), .Z(n269) );
  NAND2_X1 U245 ( .A1(n19), .A2(n18), .ZN(n270) );
  NAND2_X1 U246 ( .A1(n19), .A2(n258), .ZN(n271) );
  NAND2_X1 U247 ( .A1(n4), .A2(n18), .ZN(n272) );
  NAND3_X1 U248 ( .A1(n271), .A2(n270), .A3(n272), .ZN(n3) );
  XOR2_X1 U249 ( .A(n95), .B(n102), .Z(n56) );
  BUF_X1 U250 ( .A(n281), .Z(n273) );
  NAND2_X1 U251 ( .A1(n309), .A2(n338), .ZN(n274) );
  NAND2_X2 U252 ( .A1(n276), .A2(n277), .ZN(n309) );
  NAND2_X1 U253 ( .A1(n309), .A2(n338), .ZN(n311) );
  OR2_X1 U254 ( .A1(a[4]), .A2(a[3]), .ZN(n277) );
  NAND2_X1 U255 ( .A1(a[4]), .A2(a[3]), .ZN(n276) );
  INV_X1 U256 ( .A(n31), .ZN(n288) );
  INV_X1 U257 ( .A(n21), .ZN(n285) );
  INV_X1 U258 ( .A(n318), .ZN(n286) );
  INV_X1 U259 ( .A(n329), .ZN(n283) );
  INV_X1 U260 ( .A(n298), .ZN(n291) );
  INV_X1 U261 ( .A(n307), .ZN(n289) );
  NAND2_X1 U262 ( .A1(n299), .A2(n337), .ZN(n301) );
  INV_X1 U263 ( .A(a[5]), .ZN(n287) );
  INV_X1 U264 ( .A(a[7]), .ZN(n284) );
  XNOR2_X1 U265 ( .A(a[2]), .B(a[1]), .ZN(n299) );
  INV_X1 U266 ( .A(n299), .ZN(n278) );
  INV_X1 U267 ( .A(n278), .ZN(n279) );
  INV_X1 U268 ( .A(b[0]), .ZN(n281) );
  INV_X1 U269 ( .A(a[3]), .ZN(n290) );
  INV_X1 U270 ( .A(n227), .ZN(n292) );
  INV_X1 U271 ( .A(n281), .ZN(n280) );
  INV_X2 U272 ( .A(a[0]), .ZN(n293) );
  NOR2_X1 U273 ( .A1(n293), .A2(n273), .ZN(product[0]) );
  OAI22_X1 U274 ( .A1(n294), .A2(n295), .B1(n296), .B2(n293), .ZN(n99) );
  OAI22_X1 U275 ( .A1(n296), .A2(n295), .B1(n297), .B2(n293), .ZN(n98) );
  XNOR2_X1 U276 ( .A(b[6]), .B(n275), .ZN(n296) );
  OAI22_X1 U277 ( .A1(n293), .A2(n297), .B1(n295), .B2(n297), .ZN(n298) );
  XNOR2_X1 U278 ( .A(b[7]), .B(n275), .ZN(n297) );
  NOR2_X1 U279 ( .A1(n299), .A2(n273), .ZN(n96) );
  OAI22_X1 U280 ( .A1(n300), .A2(n301), .B1(n299), .B2(n302), .ZN(n95) );
  OAI22_X1 U281 ( .A1(n302), .A2(n301), .B1(n279), .B2(n303), .ZN(n94) );
  XNOR2_X1 U282 ( .A(b[1]), .B(a[3]), .ZN(n302) );
  OAI22_X1 U283 ( .A1(n303), .A2(n209), .B1(n279), .B2(n304), .ZN(n93) );
  XNOR2_X1 U284 ( .A(b[2]), .B(a[3]), .ZN(n303) );
  OAI22_X1 U285 ( .A1(n304), .A2(n301), .B1(n279), .B2(n305), .ZN(n92) );
  XNOR2_X1 U286 ( .A(b[3]), .B(a[3]), .ZN(n304) );
  OAI22_X1 U287 ( .A1(n305), .A2(n209), .B1(n279), .B2(n306), .ZN(n91) );
  XNOR2_X1 U288 ( .A(b[4]), .B(a[3]), .ZN(n305) );
  OAI22_X1 U289 ( .A1(n308), .A2(n279), .B1(n209), .B2(n308), .ZN(n307) );
  NOR2_X1 U290 ( .A1(n309), .A2(n273), .ZN(n88) );
  OAI22_X1 U291 ( .A1(n310), .A2(n311), .B1(n309), .B2(n312), .ZN(n87) );
  XNOR2_X1 U292 ( .A(a[5]), .B(n280), .ZN(n310) );
  OAI22_X1 U293 ( .A1(n312), .A2(n274), .B1(n309), .B2(n313), .ZN(n86) );
  XNOR2_X1 U294 ( .A(b[1]), .B(a[5]), .ZN(n312) );
  OAI22_X1 U295 ( .A1(n313), .A2(n274), .B1(n309), .B2(n314), .ZN(n85) );
  XNOR2_X1 U296 ( .A(b[2]), .B(a[5]), .ZN(n313) );
  OAI22_X1 U297 ( .A1(n314), .A2(n274), .B1(n309), .B2(n315), .ZN(n84) );
  XNOR2_X1 U298 ( .A(b[3]), .B(a[5]), .ZN(n314) );
  OAI22_X1 U299 ( .A1(n315), .A2(n274), .B1(n309), .B2(n316), .ZN(n83) );
  XNOR2_X1 U300 ( .A(b[4]), .B(a[5]), .ZN(n315) );
  OAI22_X1 U301 ( .A1(n316), .A2(n274), .B1(n309), .B2(n317), .ZN(n82) );
  XNOR2_X1 U302 ( .A(b[5]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U303 ( .A1(n319), .A2(n309), .B1(n274), .B2(n319), .ZN(n318) );
  NOR2_X1 U304 ( .A1(n320), .A2(n273), .ZN(n80) );
  OAI22_X1 U305 ( .A1(n321), .A2(n322), .B1(n320), .B2(n323), .ZN(n79) );
  XNOR2_X1 U306 ( .A(a[7]), .B(n280), .ZN(n321) );
  OAI22_X1 U307 ( .A1(n324), .A2(n322), .B1(n215), .B2(n325), .ZN(n77) );
  OAI22_X1 U308 ( .A1(n325), .A2(n322), .B1(n215), .B2(n326), .ZN(n76) );
  XNOR2_X1 U309 ( .A(b[3]), .B(a[7]), .ZN(n325) );
  OAI22_X1 U310 ( .A1(n326), .A2(n322), .B1(n215), .B2(n327), .ZN(n75) );
  XNOR2_X1 U311 ( .A(b[4]), .B(a[7]), .ZN(n326) );
  OAI22_X1 U312 ( .A1(n327), .A2(n322), .B1(n215), .B2(n328), .ZN(n74) );
  XNOR2_X1 U313 ( .A(b[5]), .B(a[7]), .ZN(n327) );
  OAI22_X1 U314 ( .A1(n330), .A2(n215), .B1(n322), .B2(n330), .ZN(n329) );
  OAI21_X1 U315 ( .B1(b[0]), .B2(n292), .A(n295), .ZN(n72) );
  OAI21_X1 U316 ( .B1(n290), .B2(n209), .A(n331), .ZN(n71) );
  OR3_X1 U317 ( .A1(n299), .A2(n280), .A3(n290), .ZN(n331) );
  OAI21_X1 U318 ( .B1(n287), .B2(n311), .A(n332), .ZN(n70) );
  OR3_X1 U319 ( .A1(n309), .A2(n280), .A3(n287), .ZN(n332) );
  OAI21_X1 U320 ( .B1(n284), .B2(n322), .A(n333), .ZN(n69) );
  OR3_X1 U321 ( .A1(n320), .A2(n280), .A3(n284), .ZN(n333) );
  XNOR2_X1 U322 ( .A(n334), .B(n335), .ZN(n38) );
  OR2_X1 U323 ( .A1(n334), .A2(n335), .ZN(n37) );
  OAI22_X1 U324 ( .A1(n306), .A2(n209), .B1(n279), .B2(n336), .ZN(n335) );
  XNOR2_X1 U325 ( .A(b[5]), .B(a[3]), .ZN(n306) );
  OAI22_X1 U326 ( .A1(n323), .A2(n322), .B1(n215), .B2(n324), .ZN(n334) );
  XNOR2_X1 U327 ( .A(b[2]), .B(a[7]), .ZN(n324) );
  XNOR2_X1 U328 ( .A(b[1]), .B(a[7]), .ZN(n323) );
  OAI22_X1 U329 ( .A1(n336), .A2(n209), .B1(n279), .B2(n308), .ZN(n31) );
  XNOR2_X1 U330 ( .A(b[7]), .B(a[3]), .ZN(n308) );
  XNOR2_X1 U331 ( .A(n290), .B(a[2]), .ZN(n337) );
  XNOR2_X1 U332 ( .A(b[6]), .B(a[3]), .ZN(n336) );
  OAI22_X1 U333 ( .A1(n317), .A2(n274), .B1(n309), .B2(n319), .ZN(n21) );
  XNOR2_X1 U334 ( .A(b[7]), .B(a[5]), .ZN(n319) );
  XNOR2_X1 U335 ( .A(n287), .B(a[4]), .ZN(n338) );
  XNOR2_X1 U336 ( .A(b[6]), .B(a[5]), .ZN(n317) );
  OAI22_X1 U337 ( .A1(n328), .A2(n322), .B1(n215), .B2(n330), .ZN(n15) );
  XNOR2_X1 U338 ( .A(b[7]), .B(a[7]), .ZN(n330) );
  NAND2_X1 U339 ( .A1(n320), .A2(n339), .ZN(n322) );
  XNOR2_X1 U340 ( .A(n284), .B(a[6]), .ZN(n339) );
  XNOR2_X1 U341 ( .A(b[6]), .B(a[7]), .ZN(n328) );
  OAI22_X1 U342 ( .A1(b[0]), .A2(n295), .B1(n340), .B2(n293), .ZN(n104) );
  OAI22_X1 U343 ( .A1(n254), .A2(n295), .B1(n341), .B2(n293), .ZN(n103) );
  XNOR2_X1 U344 ( .A(b[1]), .B(n275), .ZN(n340) );
  OAI22_X1 U345 ( .A1(n341), .A2(n295), .B1(n342), .B2(n293), .ZN(n102) );
  XNOR2_X1 U346 ( .A(b[2]), .B(n275), .ZN(n341) );
  OAI22_X1 U347 ( .A1(n342), .A2(n295), .B1(n343), .B2(n293), .ZN(n101) );
  XNOR2_X1 U348 ( .A(b[3]), .B(n275), .ZN(n342) );
  OAI22_X1 U349 ( .A1(n343), .A2(n295), .B1(n294), .B2(n293), .ZN(n100) );
  XNOR2_X1 U350 ( .A(b[5]), .B(n275), .ZN(n294) );
  XNOR2_X1 U351 ( .A(b[4]), .B(n275), .ZN(n343) );
endmodule


module datapath_DW01_add_8 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n84;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n84), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND3_X1 U1 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n1) );
  CLKBUF_X1 U2 ( .A(B[9]), .Z(n2) );
  CLKBUF_X1 U3 ( .A(n31), .Z(n3) );
  NAND3_X1 U4 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n4) );
  CLKBUF_X1 U5 ( .A(n38), .Z(n5) );
  CLKBUF_X1 U6 ( .A(n60), .Z(n6) );
  NAND3_X1 U7 ( .A1(n60), .A2(n61), .A3(n62), .ZN(n7) );
  CLKBUF_X1 U8 ( .A(n56), .Z(n8) );
  CLKBUF_X1 U9 ( .A(n66), .Z(n9) );
  CLKBUF_X1 U10 ( .A(B[11]), .Z(n10) );
  CLKBUF_X1 U11 ( .A(n53), .Z(n11) );
  NAND3_X1 U12 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n12) );
  CLKBUF_X1 U13 ( .A(B[5]), .Z(n13) );
  CLKBUF_X1 U14 ( .A(n40), .Z(n14) );
  NAND3_X1 U15 ( .A1(n20), .A2(n19), .A3(n21), .ZN(n15) );
  NAND3_X1 U16 ( .A1(n65), .A2(n9), .A3(n67), .ZN(n16) );
  CLKBUF_X1 U17 ( .A(B[4]), .Z(n17) );
  XOR2_X1 U18 ( .A(B[8]), .B(A[8]), .Z(n18) );
  XOR2_X1 U19 ( .A(n16), .B(n18), .Z(SUM[8]) );
  NAND2_X1 U20 ( .A1(n4), .A2(B[8]), .ZN(n19) );
  NAND2_X1 U21 ( .A1(carry[8]), .A2(A[8]), .ZN(n20) );
  NAND2_X1 U22 ( .A1(B[8]), .A2(A[8]), .ZN(n21) );
  NAND3_X1 U23 ( .A1(n19), .A2(n20), .A3(n21), .ZN(carry[9]) );
  CLKBUF_X1 U24 ( .A(n41), .Z(n22) );
  CLKBUF_X1 U25 ( .A(carry[13]), .Z(n23) );
  XOR2_X1 U26 ( .A(carry[2]), .B(A[2]), .Z(n24) );
  XOR2_X1 U27 ( .A(B[2]), .B(n24), .Z(SUM[2]) );
  NAND2_X1 U28 ( .A1(B[2]), .A2(carry[2]), .ZN(n25) );
  NAND2_X1 U29 ( .A1(B[2]), .A2(A[2]), .ZN(n26) );
  NAND2_X1 U30 ( .A1(carry[2]), .A2(A[2]), .ZN(n27) );
  NAND3_X1 U31 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[3]) );
  CLKBUF_X1 U32 ( .A(carry[9]), .Z(n28) );
  NAND3_X1 U33 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n29) );
  NAND3_X1 U34 ( .A1(n8), .A2(n57), .A3(n58), .ZN(n30) );
  NAND3_X1 U35 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n31) );
  XOR2_X1 U36 ( .A(B[3]), .B(A[3]), .Z(n32) );
  XOR2_X1 U37 ( .A(n12), .B(n32), .Z(SUM[3]) );
  NAND2_X1 U38 ( .A1(B[3]), .A2(n12), .ZN(n33) );
  NAND2_X1 U39 ( .A1(carry[3]), .A2(A[3]), .ZN(n34) );
  NAND2_X1 U40 ( .A1(B[3]), .A2(A[3]), .ZN(n35) );
  NAND3_X1 U41 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[4]) );
  NAND3_X1 U42 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n36) );
  XOR2_X1 U43 ( .A(n17), .B(A[4]), .Z(n37) );
  XOR2_X1 U44 ( .A(n3), .B(n37), .Z(SUM[4]) );
  NAND2_X1 U45 ( .A1(n31), .A2(B[4]), .ZN(n38) );
  NAND2_X1 U46 ( .A1(carry[4]), .A2(A[4]), .ZN(n39) );
  NAND2_X1 U47 ( .A1(B[4]), .A2(A[4]), .ZN(n40) );
  NAND3_X1 U48 ( .A1(n5), .A2(n39), .A3(n14), .ZN(carry[5]) );
  NAND3_X1 U49 ( .A1(n44), .A2(n45), .A3(n46), .ZN(n41) );
  CLKBUF_X1 U50 ( .A(n61), .Z(n42) );
  XOR2_X1 U51 ( .A(n13), .B(A[5]), .Z(n43) );
  XOR2_X1 U52 ( .A(carry[5]), .B(n43), .Z(SUM[5]) );
  NAND2_X1 U53 ( .A1(n1), .A2(B[5]), .ZN(n44) );
  NAND2_X1 U54 ( .A1(n36), .A2(A[5]), .ZN(n45) );
  NAND2_X1 U55 ( .A1(B[5]), .A2(A[5]), .ZN(n46) );
  NAND3_X1 U56 ( .A1(n44), .A2(n45), .A3(n46), .ZN(carry[6]) );
  NAND3_X1 U57 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n47) );
  NAND3_X1 U58 ( .A1(n51), .A2(n52), .A3(n11), .ZN(n48) );
  CLKBUF_X1 U59 ( .A(n72), .Z(n49) );
  XOR2_X1 U60 ( .A(n28), .B(A[9]), .Z(n50) );
  XOR2_X1 U61 ( .A(n2), .B(n50), .Z(SUM[9]) );
  NAND2_X1 U62 ( .A1(B[9]), .A2(n15), .ZN(n51) );
  NAND2_X1 U63 ( .A1(B[9]), .A2(A[9]), .ZN(n52) );
  NAND2_X1 U64 ( .A1(carry[9]), .A2(A[9]), .ZN(n53) );
  NAND3_X1 U65 ( .A1(n53), .A2(n52), .A3(n51), .ZN(carry[10]) );
  NAND3_X1 U66 ( .A1(n6), .A2(n42), .A3(n62), .ZN(n54) );
  XOR2_X1 U67 ( .A(B[6]), .B(A[6]), .Z(n55) );
  XOR2_X1 U68 ( .A(n22), .B(n55), .Z(SUM[6]) );
  NAND2_X1 U69 ( .A1(n41), .A2(B[6]), .ZN(n56) );
  NAND2_X1 U70 ( .A1(carry[6]), .A2(A[6]), .ZN(n57) );
  NAND2_X1 U71 ( .A1(B[6]), .A2(A[6]), .ZN(n58) );
  NAND3_X1 U72 ( .A1(n56), .A2(n57), .A3(n58), .ZN(carry[7]) );
  XOR2_X1 U73 ( .A(B[10]), .B(A[10]), .Z(n59) );
  XOR2_X1 U74 ( .A(n48), .B(n59), .Z(SUM[10]) );
  NAND2_X1 U75 ( .A1(n47), .A2(B[10]), .ZN(n60) );
  NAND2_X1 U76 ( .A1(carry[10]), .A2(A[10]), .ZN(n61) );
  NAND2_X1 U77 ( .A1(B[10]), .A2(A[10]), .ZN(n62) );
  NAND3_X1 U78 ( .A1(n60), .A2(n61), .A3(n62), .ZN(carry[11]) );
  NAND3_X1 U79 ( .A1(n77), .A2(n76), .A3(n78), .ZN(n63) );
  XOR2_X1 U80 ( .A(B[7]), .B(A[7]), .Z(n64) );
  XOR2_X1 U81 ( .A(n30), .B(n64), .Z(SUM[7]) );
  NAND2_X1 U82 ( .A1(n29), .A2(B[7]), .ZN(n65) );
  NAND2_X1 U83 ( .A1(carry[7]), .A2(A[7]), .ZN(n66) );
  NAND2_X1 U84 ( .A1(B[7]), .A2(A[7]), .ZN(n67) );
  NAND3_X1 U85 ( .A1(n65), .A2(n66), .A3(n67), .ZN(carry[8]) );
  NAND3_X1 U86 ( .A1(n71), .A2(n72), .A3(n73), .ZN(n68) );
  NAND3_X1 U87 ( .A1(n71), .A2(n49), .A3(n73), .ZN(n69) );
  XOR2_X1 U88 ( .A(n10), .B(A[11]), .Z(n70) );
  XOR2_X1 U89 ( .A(n54), .B(n70), .Z(SUM[11]) );
  NAND2_X1 U90 ( .A1(n7), .A2(B[11]), .ZN(n71) );
  NAND2_X1 U91 ( .A1(carry[11]), .A2(A[11]), .ZN(n72) );
  NAND2_X1 U92 ( .A1(B[11]), .A2(A[11]), .ZN(n73) );
  NAND3_X1 U93 ( .A1(n71), .A2(n72), .A3(n73), .ZN(carry[12]) );
  XNOR2_X1 U94 ( .A(carry[15]), .B(n74), .ZN(SUM[15]) );
  XNOR2_X1 U95 ( .A(B[15]), .B(A[15]), .ZN(n74) );
  XOR2_X1 U96 ( .A(A[12]), .B(B[12]), .Z(n75) );
  XOR2_X1 U97 ( .A(n75), .B(n69), .Z(SUM[12]) );
  NAND2_X1 U98 ( .A1(B[12]), .A2(A[12]), .ZN(n76) );
  NAND2_X1 U99 ( .A1(n68), .A2(A[12]), .ZN(n77) );
  NAND2_X1 U100 ( .A1(B[12]), .A2(carry[12]), .ZN(n78) );
  NAND3_X1 U101 ( .A1(n78), .A2(n77), .A3(n76), .ZN(carry[13]) );
  XOR2_X1 U102 ( .A(A[13]), .B(B[13]), .Z(n79) );
  XOR2_X1 U103 ( .A(n79), .B(n23), .Z(SUM[13]) );
  NAND2_X1 U104 ( .A1(A[13]), .A2(B[13]), .ZN(n80) );
  NAND2_X1 U105 ( .A1(A[13]), .A2(n63), .ZN(n81) );
  NAND2_X1 U106 ( .A1(carry[13]), .A2(B[13]), .ZN(n82) );
  NAND3_X1 U107 ( .A1(n80), .A2(n81), .A3(n82), .ZN(carry[14]) );
  XOR2_X1 U108 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U109 ( .A1(B[0]), .A2(A[0]), .ZN(n84) );
endmodule


module datapath_DW_mult_tc_7 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n6, n7, n8, n10, n11, n12, n13, n14, n15, n17, n18, n19, n20,
         n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76, n77, n79,
         n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94, n95, n96,
         n98, n99, n100, n101, n102, n103, n104, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342;

  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n287), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n286), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n290), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n289), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n292), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n94), .B(n88), .CI(n101), .CO(n53), .S(n54) );
  NAND2_X1 U157 ( .A1(n309), .A2(n337), .ZN(n311) );
  INV_X1 U158 ( .A(n15), .ZN(n283) );
  AND2_X1 U159 ( .A1(n95), .A2(n102), .ZN(n206) );
  XNOR2_X1 U160 ( .A(n284), .B(n15), .ZN(n207) );
  XNOR2_X1 U161 ( .A(n17), .B(n283), .ZN(n208) );
  NAND3_X1 U162 ( .A1(n270), .A2(n269), .A3(n271), .ZN(n209) );
  NAND3_X1 U163 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n210) );
  XNOR2_X1 U164 ( .A(n3), .B(n208), .ZN(product[13]) );
  AND3_X1 U165 ( .A1(n263), .A2(n264), .A3(n265), .ZN(product[15]) );
  NAND3_X1 U166 ( .A1(n223), .A2(n224), .A3(n225), .ZN(n211) );
  NAND3_X1 U167 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n212) );
  NAND3_X1 U168 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n213) );
  NAND3_X1 U169 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n214) );
  NAND3_X1 U170 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n215) );
  NAND3_X1 U171 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n216) );
  BUF_X1 U172 ( .A(b[1]), .Z(n266) );
  INV_X1 U173 ( .A(n288), .ZN(n218) );
  INV_X2 U174 ( .A(a[5]), .ZN(n288) );
  BUF_X1 U175 ( .A(n12), .Z(n219) );
  XOR2_X1 U176 ( .A(n95), .B(n102), .Z(n56) );
  CLKBUF_X1 U177 ( .A(n309), .Z(n220) );
  BUF_X2 U178 ( .A(n309), .Z(n221) );
  XOR2_X1 U179 ( .A(a[4]), .B(n291), .Z(n309) );
  XOR2_X1 U180 ( .A(n34), .B(n39), .Z(n222) );
  XOR2_X1 U181 ( .A(n216), .B(n222), .Z(product[8]) );
  NAND2_X1 U182 ( .A1(n216), .A2(n34), .ZN(n223) );
  NAND2_X1 U183 ( .A1(n8), .A2(n39), .ZN(n224) );
  NAND2_X1 U184 ( .A1(n34), .A2(n39), .ZN(n225) );
  NAND3_X1 U185 ( .A1(n223), .A2(n224), .A3(n225), .ZN(n7) );
  NAND3_X1 U186 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n226) );
  NAND3_X1 U187 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n227) );
  XOR2_X1 U188 ( .A(n33), .B(n28), .Z(n228) );
  XOR2_X1 U189 ( .A(n7), .B(n228), .Z(product[9]) );
  NAND2_X1 U190 ( .A1(n211), .A2(n33), .ZN(n229) );
  NAND2_X1 U191 ( .A1(n211), .A2(n28), .ZN(n230) );
  NAND2_X1 U192 ( .A1(n33), .A2(n28), .ZN(n231) );
  NAND3_X1 U193 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n6) );
  NAND3_X1 U194 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n232) );
  NAND3_X1 U195 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n233) );
  XNOR2_X1 U196 ( .A(n239), .B(n234), .ZN(product[5]) );
  XNOR2_X1 U197 ( .A(n50), .B(n53), .ZN(n234) );
  XOR2_X1 U198 ( .A(n46), .B(n49), .Z(n235) );
  XOR2_X1 U199 ( .A(n226), .B(n235), .Z(product[6]) );
  NAND2_X1 U200 ( .A1(n226), .A2(n46), .ZN(n236) );
  NAND2_X1 U201 ( .A1(n10), .A2(n49), .ZN(n237) );
  NAND2_X1 U202 ( .A1(n46), .A2(n49), .ZN(n238) );
  CLKBUF_X1 U203 ( .A(n11), .Z(n239) );
  NAND2_X1 U204 ( .A1(n11), .A2(n50), .ZN(n240) );
  NAND2_X1 U205 ( .A1(n210), .A2(n53), .ZN(n241) );
  NAND2_X1 U206 ( .A1(n50), .A2(n53), .ZN(n242) );
  NAND3_X1 U207 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n10) );
  XOR2_X1 U208 ( .A(n40), .B(n45), .Z(n243) );
  XOR2_X1 U209 ( .A(n233), .B(n243), .Z(product[7]) );
  NAND2_X1 U210 ( .A1(n232), .A2(n40), .ZN(n244) );
  NAND2_X1 U211 ( .A1(n232), .A2(n45), .ZN(n245) );
  NAND2_X1 U212 ( .A1(n40), .A2(n45), .ZN(n246) );
  NAND3_X1 U213 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n8) );
  XNOR2_X1 U214 ( .A(n2), .B(n207), .ZN(product[14]) );
  XOR2_X1 U215 ( .A(n18), .B(n19), .Z(n247) );
  XOR2_X1 U216 ( .A(n215), .B(n247), .Z(product[12]) );
  NAND2_X1 U217 ( .A1(n214), .A2(n18), .ZN(n248) );
  NAND2_X1 U218 ( .A1(n214), .A2(n19), .ZN(n249) );
  NAND2_X1 U219 ( .A1(n18), .A2(n19), .ZN(n250) );
  NAND3_X1 U220 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n3) );
  NAND2_X1 U221 ( .A1(n213), .A2(n17), .ZN(n251) );
  NAND2_X1 U222 ( .A1(n3), .A2(n283), .ZN(n252) );
  NAND2_X1 U223 ( .A1(n17), .A2(n283), .ZN(n253) );
  NAND3_X1 U224 ( .A1(n252), .A2(n251), .A3(n253), .ZN(n2) );
  INV_X1 U225 ( .A(n267), .ZN(n254) );
  INV_X1 U226 ( .A(n267), .ZN(n281) );
  OR2_X1 U227 ( .A1(n340), .A2(n296), .ZN(n255) );
  OR2_X1 U228 ( .A1(n341), .A2(n294), .ZN(n256) );
  NAND2_X1 U229 ( .A1(n255), .A2(n256), .ZN(n102) );
  NAND2_X2 U230 ( .A1(a[1]), .A2(n294), .ZN(n296) );
  INV_X1 U231 ( .A(a[3]), .ZN(n291) );
  NAND3_X1 U232 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n257) );
  NAND3_X1 U233 ( .A1(n270), .A2(n269), .A3(n271), .ZN(n258) );
  XOR2_X1 U234 ( .A(n54), .B(n206), .Z(n259) );
  XOR2_X1 U235 ( .A(n219), .B(n259), .Z(product[4]) );
  NAND2_X1 U236 ( .A1(n12), .A2(n54), .ZN(n260) );
  NAND2_X1 U237 ( .A1(n12), .A2(n206), .ZN(n261) );
  NAND2_X1 U238 ( .A1(n54), .A2(n206), .ZN(n262) );
  NAND3_X1 U239 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n11) );
  NAND2_X1 U240 ( .A1(n227), .A2(n284), .ZN(n263) );
  NAND2_X1 U241 ( .A1(n227), .A2(n15), .ZN(n264) );
  NAND2_X1 U242 ( .A1(n284), .A2(n15), .ZN(n265) );
  INV_X1 U243 ( .A(b[0]), .ZN(n267) );
  XOR2_X1 U244 ( .A(n27), .B(n24), .Z(n268) );
  XOR2_X1 U245 ( .A(n6), .B(n268), .Z(product[10]) );
  NAND2_X1 U246 ( .A1(n212), .A2(n27), .ZN(n269) );
  NAND2_X1 U247 ( .A1(n212), .A2(n24), .ZN(n270) );
  NAND2_X1 U248 ( .A1(n27), .A2(n24), .ZN(n271) );
  XOR2_X1 U249 ( .A(n23), .B(n20), .Z(n272) );
  XOR2_X1 U250 ( .A(n209), .B(n272), .Z(product[11]) );
  NAND2_X1 U251 ( .A1(n258), .A2(n23), .ZN(n273) );
  NAND2_X1 U252 ( .A1(n257), .A2(n20), .ZN(n274) );
  NAND2_X1 U253 ( .A1(n23), .A2(n20), .ZN(n275) );
  INV_X1 U254 ( .A(n31), .ZN(n289) );
  INV_X1 U255 ( .A(n21), .ZN(n286) );
  INV_X1 U256 ( .A(n318), .ZN(n287) );
  INV_X1 U257 ( .A(n329), .ZN(n284) );
  INV_X1 U258 ( .A(n299), .ZN(n292) );
  INV_X1 U259 ( .A(n307), .ZN(n290) );
  OR2_X2 U260 ( .A1(n276), .A2(n277), .ZN(n301) );
  XOR2_X1 U261 ( .A(a[2]), .B(a[1]), .Z(n276) );
  XOR2_X1 U262 ( .A(n279), .B(a[2]), .Z(n277) );
  INV_X1 U263 ( .A(a[7]), .ZN(n285) );
  XNOR2_X1 U264 ( .A(a[1]), .B(a[2]), .ZN(n278) );
  INV_X1 U265 ( .A(b[0]), .ZN(n282) );
  INV_X1 U266 ( .A(a[3]), .ZN(n279) );
  INV_X2 U267 ( .A(n279), .ZN(n280) );
  INV_X1 U268 ( .A(a[1]), .ZN(n293) );
  XOR2_X2 U269 ( .A(a[6]), .B(n288), .Z(n320) );
  INV_X2 U270 ( .A(a[0]), .ZN(n294) );
  NOR2_X1 U271 ( .A1(n294), .A2(n282), .ZN(product[0]) );
  OAI22_X1 U272 ( .A1(n295), .A2(n296), .B1(n297), .B2(n294), .ZN(n99) );
  OAI22_X1 U273 ( .A1(n297), .A2(n296), .B1(n298), .B2(n294), .ZN(n98) );
  XNOR2_X1 U274 ( .A(b[6]), .B(a[1]), .ZN(n297) );
  OAI22_X1 U275 ( .A1(n294), .A2(n298), .B1(n296), .B2(n298), .ZN(n299) );
  XNOR2_X1 U276 ( .A(b[7]), .B(a[1]), .ZN(n298) );
  NOR2_X1 U277 ( .A1(n278), .A2(n282), .ZN(n96) );
  OAI22_X1 U278 ( .A1(n300), .A2(n301), .B1(n302), .B2(n278), .ZN(n95) );
  XNOR2_X1 U279 ( .A(n280), .B(n281), .ZN(n300) );
  OAI22_X1 U280 ( .A1(n302), .A2(n301), .B1(n278), .B2(n303), .ZN(n94) );
  XNOR2_X1 U281 ( .A(n266), .B(n280), .ZN(n302) );
  OAI22_X1 U282 ( .A1(n303), .A2(n301), .B1(n278), .B2(n304), .ZN(n93) );
  XNOR2_X1 U283 ( .A(b[2]), .B(n280), .ZN(n303) );
  OAI22_X1 U284 ( .A1(n304), .A2(n301), .B1(n278), .B2(n305), .ZN(n92) );
  XNOR2_X1 U285 ( .A(b[3]), .B(n280), .ZN(n304) );
  OAI22_X1 U286 ( .A1(n305), .A2(n301), .B1(n278), .B2(n306), .ZN(n91) );
  XNOR2_X1 U287 ( .A(b[4]), .B(n280), .ZN(n305) );
  OAI22_X1 U288 ( .A1(n308), .A2(n278), .B1(n301), .B2(n308), .ZN(n307) );
  NOR2_X1 U289 ( .A1(n220), .A2(n282), .ZN(n88) );
  OAI22_X1 U290 ( .A1(n310), .A2(n311), .B1(n221), .B2(n312), .ZN(n87) );
  XNOR2_X1 U291 ( .A(n218), .B(n254), .ZN(n310) );
  OAI22_X1 U292 ( .A1(n312), .A2(n311), .B1(n221), .B2(n313), .ZN(n86) );
  XNOR2_X1 U293 ( .A(n266), .B(a[5]), .ZN(n312) );
  OAI22_X1 U294 ( .A1(n313), .A2(n311), .B1(n220), .B2(n314), .ZN(n85) );
  XNOR2_X1 U295 ( .A(b[2]), .B(n218), .ZN(n313) );
  OAI22_X1 U296 ( .A1(n314), .A2(n311), .B1(n220), .B2(n315), .ZN(n84) );
  XNOR2_X1 U297 ( .A(b[3]), .B(n218), .ZN(n314) );
  OAI22_X1 U298 ( .A1(n315), .A2(n311), .B1(n221), .B2(n316), .ZN(n83) );
  XNOR2_X1 U299 ( .A(b[4]), .B(n218), .ZN(n315) );
  OAI22_X1 U300 ( .A1(n316), .A2(n311), .B1(n220), .B2(n317), .ZN(n82) );
  XNOR2_X1 U301 ( .A(b[5]), .B(n218), .ZN(n316) );
  OAI22_X1 U302 ( .A1(n319), .A2(n220), .B1(n311), .B2(n319), .ZN(n318) );
  NOR2_X1 U303 ( .A1(n320), .A2(n282), .ZN(n80) );
  OAI22_X1 U304 ( .A1(n321), .A2(n322), .B1(n320), .B2(n323), .ZN(n79) );
  XNOR2_X1 U305 ( .A(a[7]), .B(n254), .ZN(n321) );
  OAI22_X1 U306 ( .A1(n324), .A2(n322), .B1(n320), .B2(n325), .ZN(n77) );
  OAI22_X1 U307 ( .A1(n325), .A2(n322), .B1(n320), .B2(n326), .ZN(n76) );
  XNOR2_X1 U308 ( .A(b[3]), .B(a[7]), .ZN(n325) );
  OAI22_X1 U309 ( .A1(n326), .A2(n322), .B1(n320), .B2(n327), .ZN(n75) );
  XNOR2_X1 U310 ( .A(b[4]), .B(a[7]), .ZN(n326) );
  OAI22_X1 U311 ( .A1(n327), .A2(n322), .B1(n320), .B2(n328), .ZN(n74) );
  XNOR2_X1 U312 ( .A(b[5]), .B(a[7]), .ZN(n327) );
  OAI22_X1 U313 ( .A1(n330), .A2(n320), .B1(n322), .B2(n330), .ZN(n329) );
  OAI21_X1 U314 ( .B1(n281), .B2(n293), .A(n296), .ZN(n72) );
  OAI21_X1 U315 ( .B1(n279), .B2(n301), .A(n331), .ZN(n71) );
  OR3_X1 U316 ( .A1(n278), .A2(n254), .A3(n279), .ZN(n331) );
  OAI21_X1 U317 ( .B1(n288), .B2(n311), .A(n332), .ZN(n70) );
  OR3_X1 U318 ( .A1(n221), .A2(n254), .A3(n288), .ZN(n332) );
  OAI21_X1 U319 ( .B1(n285), .B2(n322), .A(n333), .ZN(n69) );
  OR3_X1 U320 ( .A1(n320), .A2(n254), .A3(n285), .ZN(n333) );
  XNOR2_X1 U321 ( .A(n334), .B(n335), .ZN(n38) );
  OR2_X1 U322 ( .A1(n334), .A2(n335), .ZN(n37) );
  OAI22_X1 U323 ( .A1(n306), .A2(n301), .B1(n278), .B2(n336), .ZN(n335) );
  XNOR2_X1 U324 ( .A(b[5]), .B(n280), .ZN(n306) );
  OAI22_X1 U325 ( .A1(n323), .A2(n322), .B1(n320), .B2(n324), .ZN(n334) );
  XNOR2_X1 U326 ( .A(b[2]), .B(a[7]), .ZN(n324) );
  XNOR2_X1 U327 ( .A(n266), .B(a[7]), .ZN(n323) );
  OAI22_X1 U328 ( .A1(n336), .A2(n301), .B1(n278), .B2(n308), .ZN(n31) );
  XNOR2_X1 U329 ( .A(b[7]), .B(n280), .ZN(n308) );
  XNOR2_X1 U330 ( .A(b[6]), .B(n280), .ZN(n336) );
  OAI22_X1 U331 ( .A1(n317), .A2(n311), .B1(n221), .B2(n319), .ZN(n21) );
  XNOR2_X1 U332 ( .A(b[7]), .B(n218), .ZN(n319) );
  XNOR2_X1 U333 ( .A(n288), .B(a[4]), .ZN(n337) );
  XNOR2_X1 U334 ( .A(b[6]), .B(n218), .ZN(n317) );
  OAI22_X1 U335 ( .A1(n328), .A2(n322), .B1(n320), .B2(n330), .ZN(n15) );
  XNOR2_X1 U336 ( .A(b[7]), .B(a[7]), .ZN(n330) );
  NAND2_X1 U337 ( .A1(n320), .A2(n338), .ZN(n322) );
  XNOR2_X1 U338 ( .A(n285), .B(a[6]), .ZN(n338) );
  XNOR2_X1 U339 ( .A(b[6]), .B(a[7]), .ZN(n328) );
  OAI22_X1 U340 ( .A1(n281), .A2(n296), .B1(n339), .B2(n294), .ZN(n104) );
  OAI22_X1 U341 ( .A1(n339), .A2(n296), .B1(n340), .B2(n294), .ZN(n103) );
  XNOR2_X1 U342 ( .A(b[1]), .B(a[1]), .ZN(n339) );
  XNOR2_X1 U343 ( .A(b[2]), .B(a[1]), .ZN(n340) );
  OAI22_X1 U344 ( .A1(n341), .A2(n296), .B1(n342), .B2(n294), .ZN(n101) );
  XNOR2_X1 U345 ( .A(b[3]), .B(a[1]), .ZN(n341) );
  OAI22_X1 U346 ( .A1(n342), .A2(n296), .B1(n295), .B2(n294), .ZN(n100) );
  XNOR2_X1 U347 ( .A(b[5]), .B(a[1]), .ZN(n295) );
  XNOR2_X1 U348 ( .A(b[4]), .B(a[1]), .ZN(n342) );
endmodule


module datapath_DW01_add_7 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n80;
  wire   [15:1] carry;

  FA_X1 U1_1 ( .A(A[1]), .B(n80), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[14]), .ZN(n24) );
  NAND3_X1 U2 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n1) );
  CLKBUF_X1 U3 ( .A(n42), .Z(n2) );
  CLKBUF_X1 U4 ( .A(B[3]), .Z(n3) );
  XOR2_X1 U5 ( .A(n4), .B(n18), .Z(SUM[14]) );
  XNOR2_X1 U6 ( .A(B[14]), .B(n24), .ZN(n4) );
  XNOR2_X1 U7 ( .A(B[15]), .B(A[15]), .ZN(n70) );
  CLKBUF_X1 U8 ( .A(n47), .Z(n5) );
  CLKBUF_X1 U9 ( .A(n73), .Z(n6) );
  NAND3_X1 U10 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n7) );
  NAND3_X1 U11 ( .A1(n2), .A2(n43), .A3(n44), .ZN(n8) );
  NAND3_X1 U12 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n9) );
  CLKBUF_X1 U13 ( .A(n23), .Z(n10) );
  CLKBUF_X1 U14 ( .A(n74), .Z(n11) );
  CLKBUF_X1 U15 ( .A(n17), .Z(n12) );
  NAND3_X1 U16 ( .A1(n20), .A2(n21), .A3(n22), .ZN(n13) );
  NAND3_X1 U17 ( .A1(n52), .A2(n54), .A3(n53), .ZN(n14) );
  CLKBUF_X1 U18 ( .A(B[4]), .Z(n15) );
  CLKBUF_X1 U19 ( .A(n13), .Z(n16) );
  NAND3_X1 U20 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n17) );
  NAND3_X1 U21 ( .A1(n78), .A2(n77), .A3(n76), .ZN(n18) );
  XOR2_X1 U22 ( .A(B[7]), .B(A[7]), .Z(n19) );
  XOR2_X1 U23 ( .A(n8), .B(n19), .Z(SUM[7]) );
  NAND2_X1 U24 ( .A1(n7), .A2(B[7]), .ZN(n20) );
  NAND2_X1 U25 ( .A1(carry[7]), .A2(A[7]), .ZN(n21) );
  NAND2_X1 U26 ( .A1(B[7]), .A2(A[7]), .ZN(n22) );
  NAND3_X1 U27 ( .A1(n20), .A2(n21), .A3(n22), .ZN(carry[8]) );
  NAND3_X1 U28 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n23) );
  XOR2_X1 U29 ( .A(carry[2]), .B(A[2]), .Z(n25) );
  XOR2_X1 U30 ( .A(B[2]), .B(n25), .Z(SUM[2]) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(carry[2]), .ZN(n26) );
  NAND2_X1 U32 ( .A1(B[2]), .A2(A[2]), .ZN(n27) );
  NAND2_X1 U33 ( .A1(carry[2]), .A2(A[2]), .ZN(n28) );
  NAND3_X1 U34 ( .A1(n26), .A2(n27), .A3(n28), .ZN(carry[3]) );
  XOR2_X1 U35 ( .A(n15), .B(A[4]), .Z(n29) );
  XOR2_X1 U36 ( .A(n9), .B(n29), .Z(SUM[4]) );
  NAND2_X1 U37 ( .A1(n9), .A2(B[4]), .ZN(n30) );
  NAND2_X1 U38 ( .A1(carry[4]), .A2(A[4]), .ZN(n31) );
  NAND2_X1 U39 ( .A1(B[4]), .A2(A[4]), .ZN(n32) );
  NAND3_X1 U40 ( .A1(n31), .A2(n30), .A3(n32), .ZN(carry[5]) );
  NAND3_X1 U41 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n33) );
  NAND2_X1 U42 ( .A1(n18), .A2(B[14]), .ZN(n34) );
  NAND2_X1 U43 ( .A1(carry[14]), .A2(A[14]), .ZN(n35) );
  NAND2_X1 U44 ( .A1(B[14]), .A2(A[14]), .ZN(n36) );
  NAND3_X1 U45 ( .A1(n34), .A2(n35), .A3(n36), .ZN(carry[15]) );
  XOR2_X1 U46 ( .A(n3), .B(A[3]), .Z(n37) );
  XOR2_X1 U47 ( .A(carry[3]), .B(n37), .Z(SUM[3]) );
  NAND2_X1 U48 ( .A1(carry[3]), .A2(B[3]), .ZN(n38) );
  NAND2_X1 U49 ( .A1(carry[3]), .A2(A[3]), .ZN(n39) );
  NAND2_X1 U50 ( .A1(B[3]), .A2(A[3]), .ZN(n40) );
  NAND3_X1 U51 ( .A1(n38), .A2(n39), .A3(n40), .ZN(carry[4]) );
  XOR2_X1 U52 ( .A(B[6]), .B(A[6]), .Z(n41) );
  XOR2_X1 U53 ( .A(n14), .B(n41), .Z(SUM[6]) );
  NAND2_X1 U54 ( .A1(n14), .A2(B[6]), .ZN(n42) );
  NAND2_X1 U55 ( .A1(carry[6]), .A2(A[6]), .ZN(n43) );
  NAND2_X1 U56 ( .A1(B[6]), .A2(A[6]), .ZN(n44) );
  NAND3_X1 U57 ( .A1(n42), .A2(n43), .A3(n44), .ZN(carry[7]) );
  NAND3_X1 U58 ( .A1(n74), .A2(n73), .A3(n72), .ZN(n45) );
  XOR2_X1 U59 ( .A(B[8]), .B(A[8]), .Z(n46) );
  XOR2_X1 U60 ( .A(n16), .B(n46), .Z(SUM[8]) );
  NAND2_X1 U61 ( .A1(n13), .A2(B[8]), .ZN(n47) );
  NAND2_X1 U62 ( .A1(carry[8]), .A2(A[8]), .ZN(n48) );
  NAND2_X1 U63 ( .A1(B[8]), .A2(A[8]), .ZN(n49) );
  NAND3_X1 U64 ( .A1(n5), .A2(n48), .A3(n49), .ZN(carry[9]) );
  CLKBUF_X1 U65 ( .A(carry[12]), .Z(n50) );
  NAND2_X1 U66 ( .A1(A[12]), .A2(B[12]), .ZN(n72) );
  XOR2_X1 U67 ( .A(B[5]), .B(A[5]), .Z(n51) );
  XOR2_X1 U68 ( .A(n10), .B(n51), .Z(SUM[5]) );
  NAND2_X1 U69 ( .A1(n23), .A2(B[5]), .ZN(n52) );
  NAND2_X1 U70 ( .A1(carry[5]), .A2(A[5]), .ZN(n53) );
  NAND2_X1 U71 ( .A1(B[5]), .A2(A[5]), .ZN(n54) );
  NAND3_X1 U72 ( .A1(n52), .A2(n54), .A3(n53), .ZN(carry[6]) );
  XOR2_X1 U73 ( .A(B[9]), .B(A[9]), .Z(n55) );
  XOR2_X1 U74 ( .A(carry[9]), .B(n55), .Z(SUM[9]) );
  NAND2_X1 U75 ( .A1(n33), .A2(B[9]), .ZN(n56) );
  NAND2_X1 U76 ( .A1(n33), .A2(A[9]), .ZN(n57) );
  NAND2_X1 U77 ( .A1(B[9]), .A2(A[9]), .ZN(n58) );
  NAND3_X1 U78 ( .A1(n57), .A2(n56), .A3(n58), .ZN(carry[10]) );
  NAND3_X1 U79 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n59) );
  XOR2_X1 U80 ( .A(B[10]), .B(A[10]), .Z(n60) );
  XOR2_X1 U81 ( .A(n12), .B(n60), .Z(SUM[10]) );
  NAND2_X1 U82 ( .A1(n17), .A2(B[10]), .ZN(n61) );
  NAND2_X1 U83 ( .A1(carry[10]), .A2(A[10]), .ZN(n62) );
  NAND2_X1 U84 ( .A1(B[10]), .A2(A[10]), .ZN(n63) );
  NAND3_X1 U85 ( .A1(n61), .A2(n62), .A3(n63), .ZN(carry[11]) );
  NAND3_X1 U86 ( .A1(n66), .A2(n67), .A3(n68), .ZN(n64) );
  XOR2_X1 U87 ( .A(B[11]), .B(A[11]), .Z(n65) );
  XOR2_X1 U88 ( .A(n1), .B(n65), .Z(SUM[11]) );
  NAND2_X1 U89 ( .A1(carry[11]), .A2(B[11]), .ZN(n66) );
  NAND2_X1 U90 ( .A1(n59), .A2(A[11]), .ZN(n67) );
  NAND2_X1 U91 ( .A1(B[11]), .A2(A[11]), .ZN(n68) );
  NAND3_X1 U92 ( .A1(n67), .A2(n66), .A3(n68), .ZN(carry[12]) );
  NAND3_X1 U93 ( .A1(n72), .A2(n6), .A3(n11), .ZN(n69) );
  XNOR2_X1 U94 ( .A(carry[15]), .B(n70), .ZN(SUM[15]) );
  XOR2_X1 U95 ( .A(A[12]), .B(B[12]), .Z(n71) );
  XOR2_X1 U96 ( .A(n71), .B(n50), .Z(SUM[12]) );
  NAND2_X1 U97 ( .A1(A[12]), .A2(n64), .ZN(n73) );
  NAND2_X1 U98 ( .A1(carry[12]), .A2(B[12]), .ZN(n74) );
  NAND3_X1 U99 ( .A1(n74), .A2(n73), .A3(n72), .ZN(carry[13]) );
  XOR2_X1 U100 ( .A(A[13]), .B(B[13]), .Z(n75) );
  XOR2_X1 U101 ( .A(n75), .B(n69), .Z(SUM[13]) );
  NAND2_X1 U102 ( .A1(A[13]), .A2(B[13]), .ZN(n76) );
  NAND2_X1 U103 ( .A1(n45), .A2(A[13]), .ZN(n77) );
  NAND2_X1 U104 ( .A1(B[13]), .A2(carry[13]), .ZN(n78) );
  NAND3_X1 U105 ( .A1(n78), .A2(n77), .A3(n76), .ZN(carry[14]) );
  XOR2_X1 U106 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U107 ( .A1(B[0]), .A2(A[0]), .ZN(n80) );
endmodule


module datapath_DW_mult_tc_6 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n7, n9, n10, n11, n12, n13, n14, n15, n17, n18, n19, n20,
         n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76, n77, n79,
         n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94, n96, n98,
         n99, n100, n101, n102, n103, n104, n206, n207, n208, n209, n210, n211,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350;

  FA_X1 U10 ( .A(n46), .B(n49), .CI(n10), .CO(n9), .S(product[6]) );
  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n293), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n292), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n296), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n295), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n298), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  INV_X1 U157 ( .A(n15), .ZN(n289) );
  NAND3_X1 U158 ( .A1(n280), .A2(n281), .A3(n279), .ZN(n206) );
  NAND2_X1 U159 ( .A1(n243), .A2(n27), .ZN(n207) );
  CLKBUF_X1 U160 ( .A(b[1]), .Z(n208) );
  CLKBUF_X1 U161 ( .A(b[1]), .Z(n209) );
  AND2_X1 U162 ( .A1(n265), .A2(n102), .ZN(n210) );
  XNOR2_X1 U163 ( .A(n290), .B(n15), .ZN(n211) );
  AND3_X1 U164 ( .A1(n266), .A2(n267), .A3(n268), .ZN(product[15]) );
  BUF_X1 U165 ( .A(n9), .Z(n214) );
  CLKBUF_X1 U166 ( .A(n225), .Z(n213) );
  INV_X1 U167 ( .A(n297), .ZN(n215) );
  CLKBUF_X1 U168 ( .A(n234), .Z(n216) );
  OAI22_X1 U169 ( .A1(n307), .A2(n308), .B1(n286), .B2(n309), .ZN(n217) );
  NAND2_X2 U170 ( .A1(n327), .A2(n346), .ZN(n329) );
  NAND3_X1 U171 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n218) );
  NAND3_X1 U172 ( .A1(n213), .A2(n224), .A3(n226), .ZN(n219) );
  XOR2_X1 U173 ( .A(n217), .B(n102), .Z(n220) );
  XOR2_X1 U174 ( .A(n221), .B(n222), .Z(product[5]) );
  AND3_X1 U175 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n221) );
  XNOR2_X1 U176 ( .A(n50), .B(n53), .ZN(n222) );
  XOR2_X1 U177 ( .A(n40), .B(n45), .Z(n223) );
  XOR2_X1 U178 ( .A(n214), .B(n223), .Z(product[7]) );
  NAND2_X1 U179 ( .A1(n9), .A2(n40), .ZN(n224) );
  NAND2_X1 U180 ( .A1(n9), .A2(n45), .ZN(n225) );
  NAND2_X1 U181 ( .A1(n40), .A2(n45), .ZN(n226) );
  CLKBUF_X1 U182 ( .A(n13), .Z(n227) );
  NAND3_X1 U183 ( .A1(n280), .A2(n281), .A3(n279), .ZN(n228) );
  NAND3_X1 U184 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n229) );
  NAND3_X1 U185 ( .A1(n235), .A2(n234), .A3(n233), .ZN(n230) );
  NAND3_X1 U186 ( .A1(n235), .A2(n216), .A3(n233), .ZN(n231) );
  XNOR2_X1 U187 ( .A(n232), .B(n227), .ZN(product[3]) );
  XNOR2_X1 U188 ( .A(n56), .B(n71), .ZN(n232) );
  NAND2_X1 U189 ( .A1(n220), .A2(n71), .ZN(n233) );
  NAND2_X1 U190 ( .A1(n13), .A2(n220), .ZN(n234) );
  NAND2_X1 U191 ( .A1(n13), .A2(n71), .ZN(n235) );
  NAND3_X1 U192 ( .A1(n235), .A2(n234), .A3(n233), .ZN(n12) );
  XOR2_X1 U193 ( .A(n54), .B(n210), .Z(n236) );
  XOR2_X1 U194 ( .A(n236), .B(n231), .Z(product[4]) );
  NAND2_X1 U195 ( .A1(n54), .A2(n210), .ZN(n237) );
  NAND2_X1 U196 ( .A1(n54), .A2(n230), .ZN(n238) );
  NAND2_X1 U197 ( .A1(n12), .A2(n210), .ZN(n239) );
  NAND3_X1 U198 ( .A1(n238), .A2(n237), .A3(n239), .ZN(n11) );
  NAND2_X1 U199 ( .A1(n229), .A2(n50), .ZN(n240) );
  NAND2_X1 U200 ( .A1(n11), .A2(n53), .ZN(n241) );
  NAND2_X1 U201 ( .A1(n50), .A2(n53), .ZN(n242) );
  NAND3_X1 U202 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n10) );
  NAND3_X1 U203 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n243) );
  NAND3_X1 U204 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n244) );
  XOR2_X1 U205 ( .A(n34), .B(n39), .Z(n245) );
  XOR2_X1 U206 ( .A(n219), .B(n245), .Z(product[8]) );
  NAND2_X1 U207 ( .A1(n218), .A2(n34), .ZN(n246) );
  NAND2_X1 U208 ( .A1(n218), .A2(n39), .ZN(n247) );
  NAND2_X1 U209 ( .A1(n34), .A2(n39), .ZN(n248) );
  NAND3_X1 U210 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n7) );
  XNOR2_X1 U211 ( .A(n2), .B(n211), .ZN(product[14]) );
  NAND2_X1 U212 ( .A1(n316), .A2(n345), .ZN(n249) );
  NAND2_X1 U213 ( .A1(n316), .A2(n345), .ZN(n318) );
  NAND3_X1 U214 ( .A1(n270), .A2(n271), .A3(n272), .ZN(n250) );
  NAND3_X1 U215 ( .A1(n207), .A2(n271), .A3(n272), .ZN(n251) );
  NAND3_X1 U216 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n252) );
  XOR2_X1 U217 ( .A(n33), .B(n28), .Z(n253) );
  XOR2_X1 U218 ( .A(n244), .B(n253), .Z(product[9]) );
  NAND2_X1 U219 ( .A1(n244), .A2(n33), .ZN(n254) );
  NAND2_X1 U220 ( .A1(n7), .A2(n28), .ZN(n255) );
  NAND2_X1 U221 ( .A1(n33), .A2(n28), .ZN(n256) );
  NAND3_X1 U222 ( .A1(n262), .A2(n261), .A3(n263), .ZN(n257) );
  NAND3_X1 U223 ( .A1(n207), .A2(n271), .A3(n272), .ZN(n258) );
  NAND3_X1 U224 ( .A1(n275), .A2(n276), .A3(n277), .ZN(n259) );
  XOR2_X1 U225 ( .A(n17), .B(n289), .Z(n260) );
  XOR2_X1 U226 ( .A(n3), .B(n260), .Z(product[13]) );
  NAND2_X1 U227 ( .A1(n206), .A2(n17), .ZN(n261) );
  NAND2_X1 U228 ( .A1(n228), .A2(n289), .ZN(n262) );
  NAND2_X1 U229 ( .A1(n17), .A2(n289), .ZN(n263) );
  NAND3_X1 U230 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n2) );
  CLKBUF_X1 U231 ( .A(b[3]), .Z(n264) );
  OAI22_X1 U232 ( .A1(n307), .A2(n308), .B1(n286), .B2(n309), .ZN(n265) );
  NAND2_X1 U233 ( .A1(n257), .A2(n290), .ZN(n266) );
  NAND2_X1 U234 ( .A1(n257), .A2(n15), .ZN(n267) );
  NAND2_X1 U235 ( .A1(n290), .A2(n15), .ZN(n268) );
  XOR2_X1 U236 ( .A(n27), .B(n24), .Z(n269) );
  XOR2_X1 U237 ( .A(n243), .B(n269), .Z(product[10]) );
  NAND2_X1 U238 ( .A1(n243), .A2(n27), .ZN(n270) );
  NAND2_X1 U239 ( .A1(n252), .A2(n24), .ZN(n271) );
  NAND2_X1 U240 ( .A1(n27), .A2(n24), .ZN(n272) );
  NAND3_X1 U241 ( .A1(n275), .A2(n276), .A3(n277), .ZN(n273) );
  XOR2_X1 U242 ( .A(n20), .B(n23), .Z(n274) );
  XOR2_X1 U243 ( .A(n274), .B(n251), .Z(product[11]) );
  NAND2_X1 U244 ( .A1(n20), .A2(n23), .ZN(n275) );
  NAND2_X1 U245 ( .A1(n258), .A2(n20), .ZN(n276) );
  NAND2_X1 U246 ( .A1(n23), .A2(n250), .ZN(n277) );
  NAND3_X1 U247 ( .A1(n276), .A2(n275), .A3(n277), .ZN(n4) );
  XOR2_X1 U248 ( .A(n19), .B(n18), .Z(n278) );
  XOR2_X1 U249 ( .A(n278), .B(n259), .Z(product[12]) );
  NAND2_X1 U250 ( .A1(n19), .A2(n18), .ZN(n279) );
  NAND2_X1 U251 ( .A1(n19), .A2(n273), .ZN(n280) );
  NAND2_X1 U252 ( .A1(n4), .A2(n18), .ZN(n281) );
  NAND3_X1 U253 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n3) );
  XOR2_X1 U254 ( .A(n265), .B(n102), .Z(n56) );
  NAND2_X1 U255 ( .A1(n285), .A2(n344), .ZN(n282) );
  INV_X1 U256 ( .A(n288), .ZN(n283) );
  BUF_X2 U257 ( .A(a[1]), .Z(n284) );
  INV_X1 U258 ( .A(n31), .ZN(n295) );
  INV_X1 U259 ( .A(n21), .ZN(n292) );
  INV_X1 U260 ( .A(n325), .ZN(n293) );
  INV_X1 U261 ( .A(n336), .ZN(n290) );
  INV_X1 U262 ( .A(n305), .ZN(n298) );
  INV_X1 U263 ( .A(n314), .ZN(n296) );
  NAND2_X1 U264 ( .A1(n285), .A2(n344), .ZN(n308) );
  INV_X1 U265 ( .A(a[5]), .ZN(n294) );
  INV_X1 U266 ( .A(a[7]), .ZN(n291) );
  INV_X1 U267 ( .A(b[0]), .ZN(n288) );
  XNOR2_X2 U268 ( .A(a[4]), .B(a[3]), .ZN(n316) );
  BUF_X1 U269 ( .A(n306), .Z(n285) );
  BUF_X1 U270 ( .A(n306), .Z(n286) );
  XNOR2_X1 U271 ( .A(a[2]), .B(a[1]), .ZN(n306) );
  INV_X1 U272 ( .A(a[3]), .ZN(n297) );
  INV_X1 U273 ( .A(n284), .ZN(n299) );
  XOR2_X2 U274 ( .A(a[6]), .B(n294), .Z(n327) );
  INV_X1 U275 ( .A(n288), .ZN(n287) );
  INV_X2 U276 ( .A(a[0]), .ZN(n300) );
  NOR2_X1 U277 ( .A1(n300), .A2(n288), .ZN(product[0]) );
  OAI22_X1 U278 ( .A1(n301), .A2(n302), .B1(n303), .B2(n300), .ZN(n99) );
  OAI22_X1 U279 ( .A1(n303), .A2(n302), .B1(n304), .B2(n300), .ZN(n98) );
  XNOR2_X1 U280 ( .A(b[6]), .B(n284), .ZN(n303) );
  OAI22_X1 U281 ( .A1(n300), .A2(n304), .B1(n302), .B2(n304), .ZN(n305) );
  XNOR2_X1 U282 ( .A(b[7]), .B(n284), .ZN(n304) );
  NOR2_X1 U283 ( .A1(n286), .A2(n288), .ZN(n96) );
  XNOR2_X1 U284 ( .A(a[3]), .B(n287), .ZN(n307) );
  OAI22_X1 U285 ( .A1(n309), .A2(n282), .B1(n286), .B2(n310), .ZN(n94) );
  XNOR2_X1 U286 ( .A(n208), .B(a[3]), .ZN(n309) );
  OAI22_X1 U287 ( .A1(n310), .A2(n308), .B1(n306), .B2(n311), .ZN(n93) );
  XNOR2_X1 U288 ( .A(b[2]), .B(a[3]), .ZN(n310) );
  OAI22_X1 U289 ( .A1(n311), .A2(n282), .B1(n286), .B2(n312), .ZN(n92) );
  XNOR2_X1 U290 ( .A(n264), .B(n215), .ZN(n311) );
  OAI22_X1 U291 ( .A1(n312), .A2(n282), .B1(n286), .B2(n313), .ZN(n91) );
  XNOR2_X1 U292 ( .A(b[4]), .B(a[3]), .ZN(n312) );
  OAI22_X1 U293 ( .A1(n315), .A2(n306), .B1(n308), .B2(n315), .ZN(n314) );
  NOR2_X1 U294 ( .A1(n316), .A2(n288), .ZN(n88) );
  OAI22_X1 U295 ( .A1(n317), .A2(n318), .B1(n316), .B2(n319), .ZN(n87) );
  XNOR2_X1 U296 ( .A(a[5]), .B(n287), .ZN(n317) );
  OAI22_X1 U297 ( .A1(n319), .A2(n249), .B1(n316), .B2(n320), .ZN(n86) );
  XNOR2_X1 U298 ( .A(n209), .B(a[5]), .ZN(n319) );
  OAI22_X1 U299 ( .A1(n320), .A2(n249), .B1(n316), .B2(n321), .ZN(n85) );
  XNOR2_X1 U300 ( .A(b[2]), .B(a[5]), .ZN(n320) );
  OAI22_X1 U301 ( .A1(n321), .A2(n249), .B1(n316), .B2(n322), .ZN(n84) );
  XNOR2_X1 U302 ( .A(n264), .B(a[5]), .ZN(n321) );
  OAI22_X1 U303 ( .A1(n322), .A2(n249), .B1(n316), .B2(n323), .ZN(n83) );
  XNOR2_X1 U304 ( .A(b[4]), .B(a[5]), .ZN(n322) );
  OAI22_X1 U305 ( .A1(n323), .A2(n249), .B1(n316), .B2(n324), .ZN(n82) );
  XNOR2_X1 U306 ( .A(b[5]), .B(a[5]), .ZN(n323) );
  OAI22_X1 U307 ( .A1(n326), .A2(n316), .B1(n249), .B2(n326), .ZN(n325) );
  NOR2_X1 U308 ( .A1(n327), .A2(n288), .ZN(n80) );
  OAI22_X1 U309 ( .A1(n328), .A2(n329), .B1(n327), .B2(n330), .ZN(n79) );
  XNOR2_X1 U310 ( .A(a[7]), .B(n283), .ZN(n328) );
  OAI22_X1 U311 ( .A1(n331), .A2(n329), .B1(n327), .B2(n332), .ZN(n77) );
  OAI22_X1 U312 ( .A1(n332), .A2(n329), .B1(n327), .B2(n333), .ZN(n76) );
  XNOR2_X1 U313 ( .A(n264), .B(a[7]), .ZN(n332) );
  OAI22_X1 U314 ( .A1(n333), .A2(n329), .B1(n327), .B2(n334), .ZN(n75) );
  XNOR2_X1 U315 ( .A(b[4]), .B(a[7]), .ZN(n333) );
  OAI22_X1 U316 ( .A1(n334), .A2(n329), .B1(n327), .B2(n335), .ZN(n74) );
  XNOR2_X1 U317 ( .A(b[5]), .B(a[7]), .ZN(n334) );
  OAI22_X1 U318 ( .A1(n337), .A2(n327), .B1(n329), .B2(n337), .ZN(n336) );
  OAI21_X1 U319 ( .B1(n283), .B2(n299), .A(n302), .ZN(n72) );
  OAI21_X1 U320 ( .B1(n297), .B2(n308), .A(n338), .ZN(n71) );
  OR3_X1 U321 ( .A1(n286), .A2(n283), .A3(n297), .ZN(n338) );
  OAI21_X1 U322 ( .B1(n294), .B2(n318), .A(n339), .ZN(n70) );
  OR3_X1 U323 ( .A1(n316), .A2(n283), .A3(n294), .ZN(n339) );
  OAI21_X1 U324 ( .B1(n291), .B2(n329), .A(n340), .ZN(n69) );
  OR3_X1 U325 ( .A1(n327), .A2(n287), .A3(n291), .ZN(n340) );
  XNOR2_X1 U326 ( .A(n341), .B(n342), .ZN(n38) );
  OR2_X1 U327 ( .A1(n341), .A2(n342), .ZN(n37) );
  OAI22_X1 U328 ( .A1(n313), .A2(n308), .B1(n286), .B2(n343), .ZN(n342) );
  XNOR2_X1 U329 ( .A(b[5]), .B(n215), .ZN(n313) );
  OAI22_X1 U330 ( .A1(n330), .A2(n329), .B1(n327), .B2(n331), .ZN(n341) );
  XNOR2_X1 U331 ( .A(b[2]), .B(a[7]), .ZN(n331) );
  XNOR2_X1 U332 ( .A(n209), .B(a[7]), .ZN(n330) );
  OAI22_X1 U333 ( .A1(n343), .A2(n282), .B1(n306), .B2(n315), .ZN(n31) );
  XNOR2_X1 U334 ( .A(b[7]), .B(n215), .ZN(n315) );
  XNOR2_X1 U335 ( .A(n297), .B(a[2]), .ZN(n344) );
  XNOR2_X1 U336 ( .A(b[6]), .B(n215), .ZN(n343) );
  OAI22_X1 U337 ( .A1(n324), .A2(n249), .B1(n316), .B2(n326), .ZN(n21) );
  XNOR2_X1 U338 ( .A(b[7]), .B(a[5]), .ZN(n326) );
  XNOR2_X1 U339 ( .A(n294), .B(a[4]), .ZN(n345) );
  XNOR2_X1 U340 ( .A(b[6]), .B(a[5]), .ZN(n324) );
  OAI22_X1 U341 ( .A1(n335), .A2(n329), .B1(n327), .B2(n337), .ZN(n15) );
  XNOR2_X1 U342 ( .A(b[7]), .B(a[7]), .ZN(n337) );
  XNOR2_X1 U343 ( .A(n291), .B(a[6]), .ZN(n346) );
  XNOR2_X1 U344 ( .A(b[6]), .B(a[7]), .ZN(n335) );
  OAI22_X1 U345 ( .A1(n287), .A2(n302), .B1(n347), .B2(n300), .ZN(n104) );
  OAI22_X1 U346 ( .A1(n347), .A2(n302), .B1(n348), .B2(n300), .ZN(n103) );
  XNOR2_X1 U347 ( .A(b[1]), .B(a[1]), .ZN(n347) );
  OAI22_X1 U348 ( .A1(n348), .A2(n302), .B1(n349), .B2(n300), .ZN(n102) );
  XNOR2_X1 U349 ( .A(b[2]), .B(n284), .ZN(n348) );
  OAI22_X1 U350 ( .A1(n349), .A2(n302), .B1(n350), .B2(n300), .ZN(n101) );
  XNOR2_X1 U351 ( .A(b[3]), .B(n284), .ZN(n349) );
  OAI22_X1 U352 ( .A1(n350), .A2(n302), .B1(n301), .B2(n300), .ZN(n100) );
  XNOR2_X1 U353 ( .A(b[5]), .B(n284), .ZN(n301) );
  NAND2_X1 U354 ( .A1(a[1]), .A2(n300), .ZN(n302) );
  XNOR2_X1 U355 ( .A(b[4]), .B(n284), .ZN(n350) );
endmodule


module datapath_DW01_add_6 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n89;
  wire   [15:1] carry;

  FA_X1 U1_1 ( .A(A[1]), .B(n89), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(B[5]), .Z(n1) );
  CLKBUF_X1 U2 ( .A(n34), .Z(n2) );
  CLKBUF_X1 U3 ( .A(n26), .Z(n3) );
  CLKBUF_X1 U4 ( .A(n24), .Z(n4) );
  CLKBUF_X1 U5 ( .A(n33), .Z(n5) );
  CLKBUF_X1 U6 ( .A(n83), .Z(n6) );
  CLKBUF_X1 U7 ( .A(n58), .Z(n7) );
  NAND3_X1 U8 ( .A1(n87), .A2(n86), .A3(n85), .ZN(n8) );
  NAND3_X1 U9 ( .A1(n33), .A2(n32), .A3(n34), .ZN(n9) );
  NAND3_X1 U10 ( .A1(n32), .A2(n2), .A3(n5), .ZN(n10) );
  BUF_X1 U11 ( .A(B[14]), .Z(n11) );
  XOR2_X1 U12 ( .A(B[14]), .B(A[14]), .Z(n12) );
  XOR2_X1 U13 ( .A(n8), .B(n12), .Z(SUM[14]) );
  NAND2_X1 U14 ( .A1(n8), .A2(n11), .ZN(n13) );
  NAND2_X1 U15 ( .A1(carry[14]), .A2(A[14]), .ZN(n14) );
  NAND2_X1 U16 ( .A1(n11), .A2(A[14]), .ZN(n15) );
  NAND3_X1 U17 ( .A1(n13), .A2(n14), .A3(n15), .ZN(carry[15]) );
  NAND3_X1 U18 ( .A1(n44), .A2(n46), .A3(n45), .ZN(n16) );
  NAND3_X1 U19 ( .A1(n22), .A2(n23), .A3(n24), .ZN(n17) );
  NAND3_X1 U20 ( .A1(n22), .A2(n23), .A3(n4), .ZN(n18) );
  NAND3_X1 U21 ( .A1(n40), .A2(n41), .A3(n42), .ZN(n19) );
  NAND3_X1 U22 ( .A1(n40), .A2(n41), .A3(n42), .ZN(n20) );
  XOR2_X1 U23 ( .A(n10), .B(A[6]), .Z(n21) );
  XOR2_X1 U24 ( .A(B[6]), .B(n21), .Z(SUM[6]) );
  NAND2_X1 U25 ( .A1(B[6]), .A2(n9), .ZN(n22) );
  NAND2_X1 U26 ( .A1(B[6]), .A2(A[6]), .ZN(n23) );
  NAND2_X1 U27 ( .A1(carry[6]), .A2(A[6]), .ZN(n24) );
  NAND3_X1 U28 ( .A1(n22), .A2(n23), .A3(n24), .ZN(carry[7]) );
  NAND2_X1 U29 ( .A1(n53), .A2(A[8]), .ZN(n25) );
  NAND3_X1 U30 ( .A1(n29), .A2(n28), .A3(n30), .ZN(n26) );
  XOR2_X1 U31 ( .A(A[4]), .B(B[4]), .Z(n27) );
  XOR2_X1 U32 ( .A(n27), .B(n16), .Z(SUM[4]) );
  NAND2_X1 U33 ( .A1(A[4]), .A2(B[4]), .ZN(n28) );
  NAND2_X1 U34 ( .A1(A[4]), .A2(n16), .ZN(n29) );
  NAND2_X1 U35 ( .A1(B[4]), .A2(carry[4]), .ZN(n30) );
  NAND3_X1 U36 ( .A1(n28), .A2(n29), .A3(n30), .ZN(carry[5]) );
  XOR2_X1 U37 ( .A(A[5]), .B(n1), .Z(n31) );
  XOR2_X1 U38 ( .A(n31), .B(n3), .Z(SUM[5]) );
  NAND2_X1 U39 ( .A1(B[5]), .A2(A[5]), .ZN(n32) );
  NAND2_X1 U40 ( .A1(A[5]), .A2(n26), .ZN(n33) );
  NAND2_X1 U41 ( .A1(B[5]), .A2(carry[5]), .ZN(n34) );
  NAND3_X1 U42 ( .A1(n32), .A2(n33), .A3(n34), .ZN(carry[6]) );
  CLKBUF_X1 U43 ( .A(n76), .Z(n35) );
  CLKBUF_X1 U44 ( .A(n62), .Z(n36) );
  CLKBUF_X1 U45 ( .A(n25), .Z(n37) );
  NAND3_X1 U46 ( .A1(n35), .A2(n77), .A3(n78), .ZN(n38) );
  XOR2_X1 U47 ( .A(B[2]), .B(A[2]), .Z(n39) );
  XOR2_X1 U48 ( .A(n39), .B(carry[2]), .Z(SUM[2]) );
  NAND2_X1 U49 ( .A1(B[2]), .A2(A[2]), .ZN(n40) );
  NAND2_X1 U50 ( .A1(B[2]), .A2(carry[2]), .ZN(n41) );
  NAND2_X1 U51 ( .A1(A[2]), .A2(carry[2]), .ZN(n42) );
  NAND3_X1 U52 ( .A1(n40), .A2(n41), .A3(n42), .ZN(carry[3]) );
  XOR2_X1 U53 ( .A(A[3]), .B(B[3]), .Z(n43) );
  XOR2_X1 U54 ( .A(n43), .B(n20), .Z(SUM[3]) );
  NAND2_X1 U55 ( .A1(A[3]), .A2(B[3]), .ZN(n44) );
  NAND2_X1 U56 ( .A1(A[3]), .A2(n19), .ZN(n45) );
  NAND2_X1 U57 ( .A1(B[3]), .A2(carry[3]), .ZN(n46) );
  NAND3_X1 U58 ( .A1(n44), .A2(n45), .A3(n46), .ZN(carry[4]) );
  NAND2_X1 U59 ( .A1(A[12]), .A2(B[12]), .ZN(n81) );
  CLKBUF_X1 U60 ( .A(n52), .Z(n47) );
  CLKBUF_X1 U61 ( .A(n82), .Z(n48) );
  NAND3_X1 U62 ( .A1(n71), .A2(n72), .A3(n73), .ZN(n49) );
  NAND3_X1 U63 ( .A1(n25), .A2(n62), .A3(n60), .ZN(n50) );
  NAND3_X1 U64 ( .A1(n60), .A2(n37), .A3(n36), .ZN(n51) );
  NAND3_X1 U65 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n52) );
  NAND3_X1 U66 ( .A1(n57), .A2(n58), .A3(n56), .ZN(n53) );
  NAND3_X1 U67 ( .A1(n56), .A2(n57), .A3(n7), .ZN(n54) );
  XOR2_X1 U68 ( .A(A[7]), .B(B[7]), .Z(n55) );
  XOR2_X1 U69 ( .A(n55), .B(n18), .Z(SUM[7]) );
  NAND2_X1 U70 ( .A1(A[7]), .A2(B[7]), .ZN(n56) );
  NAND2_X1 U71 ( .A1(A[7]), .A2(n17), .ZN(n57) );
  NAND2_X1 U72 ( .A1(B[7]), .A2(carry[7]), .ZN(n58) );
  NAND3_X1 U73 ( .A1(n58), .A2(n57), .A3(n56), .ZN(carry[8]) );
  XOR2_X1 U74 ( .A(A[8]), .B(B[8]), .Z(n59) );
  XOR2_X1 U75 ( .A(n59), .B(n54), .Z(SUM[8]) );
  NAND2_X1 U76 ( .A1(A[8]), .A2(B[8]), .ZN(n60) );
  NAND2_X1 U77 ( .A1(n53), .A2(A[8]), .ZN(n61) );
  NAND2_X1 U78 ( .A1(carry[8]), .A2(B[8]), .ZN(n62) );
  NAND3_X1 U79 ( .A1(n62), .A2(n61), .A3(n60), .ZN(carry[9]) );
  XOR2_X1 U80 ( .A(B[9]), .B(A[9]), .Z(n63) );
  XOR2_X1 U81 ( .A(n51), .B(n63), .Z(SUM[9]) );
  NAND2_X1 U82 ( .A1(n50), .A2(B[9]), .ZN(n64) );
  NAND2_X1 U83 ( .A1(carry[9]), .A2(A[9]), .ZN(n65) );
  NAND2_X1 U84 ( .A1(B[9]), .A2(A[9]), .ZN(n66) );
  NAND3_X1 U85 ( .A1(n65), .A2(n64), .A3(n66), .ZN(carry[10]) );
  CLKBUF_X1 U86 ( .A(n49), .Z(n67) );
  NAND3_X1 U87 ( .A1(n81), .A2(n82), .A3(n83), .ZN(n68) );
  NAND3_X1 U88 ( .A1(n81), .A2(n48), .A3(n6), .ZN(n69) );
  XOR2_X1 U89 ( .A(B[10]), .B(A[10]), .Z(n70) );
  XOR2_X1 U90 ( .A(n47), .B(n70), .Z(SUM[10]) );
  NAND2_X1 U91 ( .A1(n52), .A2(B[10]), .ZN(n71) );
  NAND2_X1 U92 ( .A1(carry[10]), .A2(A[10]), .ZN(n72) );
  NAND2_X1 U93 ( .A1(B[10]), .A2(A[10]), .ZN(n73) );
  NAND3_X1 U94 ( .A1(n71), .A2(n72), .A3(n73), .ZN(carry[11]) );
  NAND3_X1 U95 ( .A1(n76), .A2(n77), .A3(n78), .ZN(n74) );
  XOR2_X1 U96 ( .A(B[11]), .B(A[11]), .Z(n75) );
  XOR2_X1 U97 ( .A(n67), .B(n75), .Z(SUM[11]) );
  NAND2_X1 U98 ( .A1(n49), .A2(B[11]), .ZN(n76) );
  NAND2_X1 U99 ( .A1(carry[11]), .A2(A[11]), .ZN(n77) );
  NAND2_X1 U100 ( .A1(B[11]), .A2(A[11]), .ZN(n78) );
  NAND3_X1 U101 ( .A1(n76), .A2(n77), .A3(n78), .ZN(carry[12]) );
  XNOR2_X1 U102 ( .A(carry[15]), .B(n79), .ZN(SUM[15]) );
  XNOR2_X1 U103 ( .A(B[15]), .B(A[15]), .ZN(n79) );
  XOR2_X1 U104 ( .A(A[12]), .B(B[12]), .Z(n80) );
  XOR2_X1 U105 ( .A(n80), .B(n38), .Z(SUM[12]) );
  NAND2_X1 U106 ( .A1(n74), .A2(A[12]), .ZN(n82) );
  NAND2_X1 U107 ( .A1(carry[12]), .A2(B[12]), .ZN(n83) );
  NAND3_X1 U108 ( .A1(n83), .A2(n82), .A3(n81), .ZN(carry[13]) );
  XOR2_X1 U109 ( .A(A[13]), .B(B[13]), .Z(n84) );
  XOR2_X1 U110 ( .A(n84), .B(n69), .Z(SUM[13]) );
  NAND2_X1 U111 ( .A1(A[13]), .A2(B[13]), .ZN(n85) );
  NAND2_X1 U112 ( .A1(n68), .A2(A[13]), .ZN(n86) );
  NAND2_X1 U113 ( .A1(B[13]), .A2(carry[13]), .ZN(n87) );
  NAND3_X1 U114 ( .A1(n86), .A2(n87), .A3(n85), .ZN(carry[14]) );
  XOR2_X1 U115 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U116 ( .A1(B[0]), .A2(A[0]), .ZN(n89) );
endmodule


module datapath_DW_mult_tc_5 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343;

  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n286), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n285), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n289), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n288), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n291), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  INV_X1 U157 ( .A(n292), .ZN(n213) );
  INV_X1 U158 ( .A(n15), .ZN(n282) );
  BUF_X2 U159 ( .A(n299), .Z(n279) );
  NAND2_X2 U160 ( .A1(n293), .A2(a[1]), .ZN(n295) );
  AND2_X1 U161 ( .A1(n95), .A2(n102), .ZN(n206) );
  XNOR2_X1 U162 ( .A(n283), .B(n15), .ZN(n207) );
  AND3_X1 U163 ( .A1(n275), .A2(n276), .A3(n277), .ZN(product[15]) );
  XNOR2_X1 U164 ( .A(n209), .B(n258), .ZN(product[13]) );
  AND3_X1 U165 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n209) );
  INV_X1 U166 ( .A(a[3]), .ZN(n210) );
  XNOR2_X1 U167 ( .A(a[6]), .B(a[5]), .ZN(n320) );
  BUF_X1 U168 ( .A(b[1]), .Z(n212) );
  XNOR2_X1 U169 ( .A(n212), .B(a[1]), .ZN(n211) );
  XNOR2_X1 U170 ( .A(a[4]), .B(a[3]), .ZN(n222) );
  XNOR2_X1 U171 ( .A(n210), .B(a[2]), .ZN(n337) );
  CLKBUF_X1 U172 ( .A(n12), .Z(n214) );
  XNOR2_X1 U173 ( .A(n214), .B(n215), .ZN(product[4]) );
  XNOR2_X1 U174 ( .A(n54), .B(n206), .ZN(n215) );
  XNOR2_X1 U175 ( .A(n228), .B(n216), .ZN(product[5]) );
  XNOR2_X1 U176 ( .A(n50), .B(n53), .ZN(n216) );
  NAND3_X1 U177 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n217) );
  NAND3_X1 U178 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n218) );
  NAND3_X1 U179 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n219) );
  XOR2_X1 U180 ( .A(n220), .B(n221), .Z(product[8]) );
  XNOR2_X1 U181 ( .A(n34), .B(n39), .ZN(n220) );
  AND3_X1 U182 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n221) );
  XNOR2_X1 U183 ( .A(a[4]), .B(a[3]), .ZN(n309) );
  CLKBUF_X1 U184 ( .A(b[1]), .Z(n223) );
  NAND3_X1 U185 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n224) );
  NAND3_X1 U186 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n225) );
  NAND3_X1 U187 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n226) );
  NAND3_X1 U188 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n227) );
  NAND3_X1 U189 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n228) );
  NAND2_X1 U190 ( .A1(n12), .A2(n54), .ZN(n229) );
  NAND2_X1 U191 ( .A1(n12), .A2(n206), .ZN(n230) );
  NAND2_X1 U192 ( .A1(n54), .A2(n206), .ZN(n231) );
  NAND3_X1 U193 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n11) );
  XOR2_X1 U194 ( .A(n23), .B(n20), .Z(n232) );
  XOR2_X1 U195 ( .A(n218), .B(n232), .Z(product[11]) );
  NAND2_X1 U196 ( .A1(n217), .A2(n23), .ZN(n233) );
  NAND2_X1 U197 ( .A1(n5), .A2(n20), .ZN(n234) );
  NAND2_X1 U198 ( .A1(n23), .A2(n20), .ZN(n235) );
  NAND3_X1 U199 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n4) );
  NAND3_X1 U200 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n236) );
  NAND3_X1 U201 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n237) );
  NAND3_X1 U202 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n238) );
  XOR2_X1 U203 ( .A(n27), .B(n24), .Z(n239) );
  XOR2_X1 U204 ( .A(n238), .B(n239), .Z(product[10]) );
  NAND2_X1 U205 ( .A1(n237), .A2(n27), .ZN(n240) );
  NAND2_X1 U206 ( .A1(n6), .A2(n24), .ZN(n241) );
  NAND2_X1 U207 ( .A1(n27), .A2(n24), .ZN(n242) );
  NAND3_X1 U208 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n5) );
  XOR2_X1 U209 ( .A(n18), .B(n19), .Z(n243) );
  XOR2_X1 U210 ( .A(n226), .B(n243), .Z(product[12]) );
  NAND2_X1 U211 ( .A1(n225), .A2(n18), .ZN(n244) );
  NAND2_X1 U212 ( .A1(n4), .A2(n19), .ZN(n245) );
  NAND2_X1 U213 ( .A1(n18), .A2(n19), .ZN(n246) );
  NAND3_X1 U214 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n3) );
  NAND2_X1 U215 ( .A1(n228), .A2(n50), .ZN(n247) );
  NAND2_X1 U216 ( .A1(n11), .A2(n53), .ZN(n248) );
  NAND2_X1 U217 ( .A1(n50), .A2(n53), .ZN(n249) );
  NAND3_X1 U218 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n10) );
  XOR2_X1 U219 ( .A(n46), .B(n49), .Z(n250) );
  XOR2_X1 U220 ( .A(n236), .B(n250), .Z(product[6]) );
  NAND2_X1 U221 ( .A1(n236), .A2(n46), .ZN(n251) );
  NAND2_X1 U222 ( .A1(n10), .A2(n49), .ZN(n252) );
  NAND2_X1 U223 ( .A1(n46), .A2(n49), .ZN(n253) );
  NAND3_X1 U224 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n9) );
  XOR2_X1 U225 ( .A(n40), .B(n45), .Z(n254) );
  XOR2_X1 U226 ( .A(n224), .B(n254), .Z(product[7]) );
  NAND2_X1 U227 ( .A1(n9), .A2(n40), .ZN(n255) );
  NAND2_X1 U228 ( .A1(n9), .A2(n45), .ZN(n256) );
  NAND2_X1 U229 ( .A1(n40), .A2(n45), .ZN(n257) );
  NAND3_X1 U230 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n8) );
  XOR2_X1 U231 ( .A(n17), .B(n282), .Z(n258) );
  NAND2_X1 U232 ( .A1(n227), .A2(n17), .ZN(n259) );
  NAND2_X1 U233 ( .A1(n3), .A2(n282), .ZN(n260) );
  NAND2_X1 U234 ( .A1(n17), .A2(n282), .ZN(n261) );
  NAND3_X1 U235 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n2) );
  NAND2_X1 U236 ( .A1(n222), .A2(n338), .ZN(n262) );
  NAND2_X1 U237 ( .A1(n222), .A2(n338), .ZN(n263) );
  NAND2_X1 U238 ( .A1(n309), .A2(n338), .ZN(n311) );
  XNOR2_X1 U239 ( .A(n219), .B(n207), .ZN(product[14]) );
  XOR2_X1 U240 ( .A(n102), .B(n95), .Z(n56) );
  NAND3_X1 U241 ( .A1(n270), .A2(n269), .A3(n268), .ZN(n264) );
  NAND3_X1 U242 ( .A1(n270), .A2(n269), .A3(n268), .ZN(n265) );
  NAND2_X1 U243 ( .A1(n278), .A2(n337), .ZN(n266) );
  NAND2_X1 U244 ( .A1(n278), .A2(n337), .ZN(n267) );
  NAND2_X1 U245 ( .A1(n278), .A2(n337), .ZN(n301) );
  NAND2_X1 U246 ( .A1(n34), .A2(n39), .ZN(n268) );
  NAND2_X1 U247 ( .A1(n34), .A2(n8), .ZN(n269) );
  NAND2_X1 U248 ( .A1(n39), .A2(n8), .ZN(n270) );
  NAND3_X1 U249 ( .A1(n269), .A2(n268), .A3(n270), .ZN(n7) );
  XOR2_X1 U250 ( .A(n28), .B(n33), .Z(n271) );
  XOR2_X1 U251 ( .A(n271), .B(n265), .Z(product[9]) );
  NAND2_X1 U252 ( .A1(n28), .A2(n33), .ZN(n272) );
  NAND2_X1 U253 ( .A1(n28), .A2(n264), .ZN(n273) );
  NAND2_X1 U254 ( .A1(n33), .A2(n7), .ZN(n274) );
  NAND3_X1 U255 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n6) );
  NAND2_X1 U256 ( .A1(n2), .A2(n283), .ZN(n275) );
  NAND2_X1 U257 ( .A1(n2), .A2(n15), .ZN(n276) );
  NAND2_X1 U258 ( .A1(n283), .A2(n15), .ZN(n277) );
  INV_X1 U259 ( .A(n31), .ZN(n288) );
  INV_X1 U260 ( .A(n21), .ZN(n285) );
  INV_X1 U261 ( .A(n318), .ZN(n286) );
  INV_X1 U262 ( .A(n329), .ZN(n283) );
  INV_X1 U263 ( .A(n298), .ZN(n291) );
  INV_X1 U264 ( .A(n307), .ZN(n289) );
  INV_X1 U265 ( .A(a[5]), .ZN(n287) );
  INV_X1 U266 ( .A(a[7]), .ZN(n284) );
  INV_X1 U267 ( .A(b[0]), .ZN(n281) );
  BUF_X1 U268 ( .A(n299), .Z(n278) );
  XNOR2_X1 U269 ( .A(a[2]), .B(a[1]), .ZN(n299) );
  INV_X1 U270 ( .A(a[3]), .ZN(n290) );
  INV_X1 U271 ( .A(a[1]), .ZN(n292) );
  INV_X1 U272 ( .A(n281), .ZN(n280) );
  INV_X2 U273 ( .A(a[0]), .ZN(n293) );
  NOR2_X1 U274 ( .A1(n293), .A2(n281), .ZN(product[0]) );
  OAI22_X1 U275 ( .A1(n294), .A2(n295), .B1(n296), .B2(n293), .ZN(n99) );
  OAI22_X1 U276 ( .A1(n296), .A2(n295), .B1(n297), .B2(n293), .ZN(n98) );
  XNOR2_X1 U277 ( .A(b[6]), .B(n213), .ZN(n296) );
  OAI22_X1 U278 ( .A1(n293), .A2(n297), .B1(n295), .B2(n297), .ZN(n298) );
  XNOR2_X1 U279 ( .A(b[7]), .B(n213), .ZN(n297) );
  NOR2_X1 U280 ( .A1(n279), .A2(n281), .ZN(n96) );
  OAI22_X1 U281 ( .A1(n300), .A2(n301), .B1(n302), .B2(n279), .ZN(n95) );
  XNOR2_X1 U282 ( .A(a[3]), .B(n280), .ZN(n300) );
  OAI22_X1 U283 ( .A1(n302), .A2(n266), .B1(n279), .B2(n303), .ZN(n94) );
  XNOR2_X1 U284 ( .A(n212), .B(a[3]), .ZN(n302) );
  OAI22_X1 U285 ( .A1(n303), .A2(n267), .B1(n279), .B2(n304), .ZN(n93) );
  XNOR2_X1 U286 ( .A(b[2]), .B(a[3]), .ZN(n303) );
  OAI22_X1 U287 ( .A1(n304), .A2(n266), .B1(n279), .B2(n305), .ZN(n92) );
  XNOR2_X1 U288 ( .A(b[3]), .B(a[3]), .ZN(n304) );
  OAI22_X1 U289 ( .A1(n305), .A2(n266), .B1(n279), .B2(n306), .ZN(n91) );
  XNOR2_X1 U290 ( .A(b[4]), .B(a[3]), .ZN(n305) );
  OAI22_X1 U291 ( .A1(n308), .A2(n279), .B1(n266), .B2(n308), .ZN(n307) );
  NOR2_X1 U292 ( .A1(n222), .A2(n281), .ZN(n88) );
  OAI22_X1 U293 ( .A1(n310), .A2(n311), .B1(n222), .B2(n312), .ZN(n87) );
  XNOR2_X1 U294 ( .A(a[5]), .B(n280), .ZN(n310) );
  OAI22_X1 U295 ( .A1(n312), .A2(n262), .B1(n222), .B2(n313), .ZN(n86) );
  XNOR2_X1 U296 ( .A(n223), .B(a[5]), .ZN(n312) );
  OAI22_X1 U297 ( .A1(n313), .A2(n263), .B1(n222), .B2(n314), .ZN(n85) );
  XNOR2_X1 U298 ( .A(b[2]), .B(a[5]), .ZN(n313) );
  OAI22_X1 U299 ( .A1(n314), .A2(n263), .B1(n222), .B2(n315), .ZN(n84) );
  XNOR2_X1 U300 ( .A(b[3]), .B(a[5]), .ZN(n314) );
  OAI22_X1 U301 ( .A1(n315), .A2(n262), .B1(n222), .B2(n316), .ZN(n83) );
  XNOR2_X1 U302 ( .A(b[4]), .B(a[5]), .ZN(n315) );
  OAI22_X1 U303 ( .A1(n316), .A2(n263), .B1(n222), .B2(n317), .ZN(n82) );
  XNOR2_X1 U304 ( .A(b[5]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U305 ( .A1(n319), .A2(n222), .B1(n262), .B2(n319), .ZN(n318) );
  NOR2_X1 U306 ( .A1(n320), .A2(n281), .ZN(n80) );
  OAI22_X1 U307 ( .A1(n321), .A2(n322), .B1(n320), .B2(n323), .ZN(n79) );
  XNOR2_X1 U308 ( .A(a[7]), .B(n280), .ZN(n321) );
  OAI22_X1 U309 ( .A1(n324), .A2(n322), .B1(n320), .B2(n325), .ZN(n77) );
  OAI22_X1 U310 ( .A1(n325), .A2(n322), .B1(n320), .B2(n326), .ZN(n76) );
  XNOR2_X1 U311 ( .A(b[3]), .B(a[7]), .ZN(n325) );
  OAI22_X1 U312 ( .A1(n326), .A2(n322), .B1(n320), .B2(n327), .ZN(n75) );
  XNOR2_X1 U313 ( .A(b[4]), .B(a[7]), .ZN(n326) );
  OAI22_X1 U314 ( .A1(n327), .A2(n322), .B1(n320), .B2(n328), .ZN(n74) );
  XNOR2_X1 U315 ( .A(b[5]), .B(a[7]), .ZN(n327) );
  OAI22_X1 U316 ( .A1(n330), .A2(n320), .B1(n322), .B2(n330), .ZN(n329) );
  OAI21_X1 U317 ( .B1(n280), .B2(n292), .A(n295), .ZN(n72) );
  OAI21_X1 U318 ( .B1(n290), .B2(n267), .A(n331), .ZN(n71) );
  OR3_X1 U319 ( .A1(n279), .A2(n280), .A3(n290), .ZN(n331) );
  OAI21_X1 U320 ( .B1(n287), .B2(n311), .A(n332), .ZN(n70) );
  OR3_X1 U321 ( .A1(n309), .A2(n280), .A3(n287), .ZN(n332) );
  OAI21_X1 U322 ( .B1(n284), .B2(n322), .A(n333), .ZN(n69) );
  OR3_X1 U323 ( .A1(n320), .A2(n280), .A3(n284), .ZN(n333) );
  XNOR2_X1 U324 ( .A(n334), .B(n335), .ZN(n38) );
  OR2_X1 U325 ( .A1(n334), .A2(n335), .ZN(n37) );
  OAI22_X1 U326 ( .A1(n306), .A2(n267), .B1(n279), .B2(n336), .ZN(n335) );
  XNOR2_X1 U327 ( .A(b[5]), .B(a[3]), .ZN(n306) );
  OAI22_X1 U328 ( .A1(n323), .A2(n322), .B1(n320), .B2(n324), .ZN(n334) );
  XNOR2_X1 U329 ( .A(b[2]), .B(a[7]), .ZN(n324) );
  XNOR2_X1 U330 ( .A(n223), .B(a[7]), .ZN(n323) );
  OAI22_X1 U331 ( .A1(n336), .A2(n267), .B1(n279), .B2(n308), .ZN(n31) );
  XNOR2_X1 U332 ( .A(b[7]), .B(a[3]), .ZN(n308) );
  XNOR2_X1 U333 ( .A(b[6]), .B(a[3]), .ZN(n336) );
  OAI22_X1 U334 ( .A1(n317), .A2(n263), .B1(n222), .B2(n319), .ZN(n21) );
  XNOR2_X1 U335 ( .A(b[7]), .B(a[5]), .ZN(n319) );
  XNOR2_X1 U336 ( .A(n287), .B(a[4]), .ZN(n338) );
  XNOR2_X1 U337 ( .A(b[6]), .B(a[5]), .ZN(n317) );
  OAI22_X1 U338 ( .A1(n328), .A2(n322), .B1(n320), .B2(n330), .ZN(n15) );
  XNOR2_X1 U339 ( .A(b[7]), .B(a[7]), .ZN(n330) );
  NAND2_X1 U340 ( .A1(n320), .A2(n339), .ZN(n322) );
  XNOR2_X1 U341 ( .A(n284), .B(a[6]), .ZN(n339) );
  XNOR2_X1 U342 ( .A(b[6]), .B(a[7]), .ZN(n328) );
  OAI22_X1 U343 ( .A1(n280), .A2(n295), .B1(n340), .B2(n293), .ZN(n104) );
  OAI22_X1 U344 ( .A1(n211), .A2(n295), .B1(n341), .B2(n293), .ZN(n103) );
  XNOR2_X1 U345 ( .A(b[1]), .B(a[1]), .ZN(n340) );
  OAI22_X1 U346 ( .A1(n341), .A2(n295), .B1(n342), .B2(n293), .ZN(n102) );
  XNOR2_X1 U347 ( .A(b[2]), .B(a[1]), .ZN(n341) );
  OAI22_X1 U348 ( .A1(n342), .A2(n295), .B1(n343), .B2(n293), .ZN(n101) );
  XNOR2_X1 U349 ( .A(b[3]), .B(a[1]), .ZN(n342) );
  OAI22_X1 U350 ( .A1(n343), .A2(n295), .B1(n293), .B2(n294), .ZN(n100) );
  XNOR2_X1 U351 ( .A(b[5]), .B(n213), .ZN(n294) );
  XNOR2_X1 U352 ( .A(b[4]), .B(n213), .ZN(n343) );
endmodule


module datapath_DW01_add_5 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n82;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n82), .CO(carry[2]), .S(SUM[1]) );
  NAND3_X1 U1 ( .A1(n5), .A2(n6), .A3(n7), .ZN(n1) );
  NAND3_X1 U2 ( .A1(n5), .A2(n6), .A3(n7), .ZN(n2) );
  NAND3_X1 U3 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n3) );
  XOR2_X1 U4 ( .A(carry[2]), .B(A[2]), .Z(n4) );
  XOR2_X1 U5 ( .A(B[2]), .B(n4), .Z(SUM[2]) );
  NAND2_X1 U6 ( .A1(B[2]), .A2(carry[2]), .ZN(n5) );
  NAND2_X1 U7 ( .A1(B[2]), .A2(A[2]), .ZN(n6) );
  NAND2_X1 U8 ( .A1(carry[2]), .A2(A[2]), .ZN(n7) );
  NAND3_X1 U9 ( .A1(n5), .A2(n6), .A3(n7), .ZN(carry[3]) );
  CLKBUF_X1 U10 ( .A(B[3]), .Z(n8) );
  XNOR2_X1 U11 ( .A(B[15]), .B(A[15]), .ZN(n80) );
  CLKBUF_X1 U12 ( .A(carry[6]), .Z(n9) );
  CLKBUF_X1 U13 ( .A(n51), .Z(n10) );
  NAND3_X1 U14 ( .A1(n49), .A2(n48), .A3(n50), .ZN(n11) );
  CLKBUF_X1 U15 ( .A(n65), .Z(n12) );
  NAND3_X1 U16 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n13) );
  NAND3_X1 U17 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n14) );
  CLKBUF_X1 U18 ( .A(n45), .Z(n15) );
  CLKBUF_X1 U19 ( .A(n79), .Z(n16) );
  NAND3_X1 U20 ( .A1(n36), .A2(n38), .A3(n37), .ZN(n17) );
  CLKBUF_X1 U21 ( .A(n13), .Z(n18) );
  CLKBUF_X1 U22 ( .A(n78), .Z(n19) );
  XOR2_X1 U23 ( .A(B[4]), .B(A[4]), .Z(n20) );
  XOR2_X1 U24 ( .A(n14), .B(n20), .Z(SUM[4]) );
  NAND2_X1 U25 ( .A1(n3), .A2(B[4]), .ZN(n21) );
  NAND2_X1 U26 ( .A1(carry[4]), .A2(A[4]), .ZN(n22) );
  NAND2_X1 U27 ( .A1(B[4]), .A2(A[4]), .ZN(n23) );
  NAND3_X1 U28 ( .A1(n22), .A2(n21), .A3(n23), .ZN(carry[5]) );
  XOR2_X1 U29 ( .A(n8), .B(A[3]), .Z(n24) );
  XOR2_X1 U30 ( .A(carry[3]), .B(n24), .Z(SUM[3]) );
  NAND2_X1 U31 ( .A1(n2), .A2(B[3]), .ZN(n25) );
  NAND2_X1 U32 ( .A1(n1), .A2(A[3]), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[3]), .A2(A[3]), .ZN(n27) );
  NAND3_X1 U34 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[4]) );
  NAND3_X1 U35 ( .A1(n49), .A2(n48), .A3(n50), .ZN(n28) );
  NAND3_X1 U36 ( .A1(n77), .A2(n19), .A3(n16), .ZN(n29) );
  CLKBUF_X1 U37 ( .A(n75), .Z(n30) );
  NAND3_X1 U38 ( .A1(n44), .A2(n45), .A3(n46), .ZN(n31) );
  NAND3_X1 U39 ( .A1(n44), .A2(n15), .A3(n46), .ZN(n32) );
  CLKBUF_X1 U40 ( .A(n74), .Z(n33) );
  CLKBUF_X1 U41 ( .A(n49), .Z(n34) );
  XOR2_X1 U42 ( .A(B[5]), .B(A[5]), .Z(n35) );
  XOR2_X1 U43 ( .A(n18), .B(n35), .Z(SUM[5]) );
  NAND2_X1 U44 ( .A1(n13), .A2(B[5]), .ZN(n36) );
  NAND2_X1 U45 ( .A1(carry[5]), .A2(A[5]), .ZN(n37) );
  NAND2_X1 U46 ( .A1(B[5]), .A2(A[5]), .ZN(n38) );
  NAND3_X1 U47 ( .A1(n36), .A2(n37), .A3(n38), .ZN(carry[6]) );
  NAND3_X1 U48 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n39) );
  NAND3_X1 U49 ( .A1(n64), .A2(n12), .A3(n66), .ZN(n40) );
  NAND3_X1 U50 ( .A1(n48), .A2(n34), .A3(n50), .ZN(n41) );
  NAND3_X1 U51 ( .A1(n57), .A2(n58), .A3(n59), .ZN(n42) );
  XOR2_X1 U52 ( .A(B[10]), .B(A[10]), .Z(n43) );
  XOR2_X1 U53 ( .A(n40), .B(n43), .Z(SUM[10]) );
  NAND2_X1 U54 ( .A1(n39), .A2(B[10]), .ZN(n44) );
  NAND2_X1 U55 ( .A1(carry[10]), .A2(A[10]), .ZN(n45) );
  NAND2_X1 U56 ( .A1(B[10]), .A2(A[10]), .ZN(n46) );
  NAND3_X1 U57 ( .A1(n44), .A2(n45), .A3(n46), .ZN(carry[11]) );
  XOR2_X1 U58 ( .A(B[6]), .B(A[6]), .Z(n47) );
  XOR2_X1 U59 ( .A(n9), .B(n47), .Z(SUM[6]) );
  NAND2_X1 U60 ( .A1(n17), .A2(B[6]), .ZN(n48) );
  NAND2_X1 U61 ( .A1(carry[6]), .A2(A[6]), .ZN(n49) );
  NAND2_X1 U62 ( .A1(B[6]), .A2(A[6]), .ZN(n50) );
  NAND3_X1 U63 ( .A1(n53), .A2(n55), .A3(n54), .ZN(n51) );
  XOR2_X1 U64 ( .A(n32), .B(A[11]), .Z(n52) );
  XOR2_X1 U65 ( .A(B[11]), .B(n52), .Z(SUM[11]) );
  NAND2_X1 U66 ( .A1(B[11]), .A2(n31), .ZN(n53) );
  NAND2_X1 U67 ( .A1(B[11]), .A2(A[11]), .ZN(n54) );
  NAND2_X1 U68 ( .A1(carry[11]), .A2(A[11]), .ZN(n55) );
  NAND3_X1 U69 ( .A1(n53), .A2(n55), .A3(n54), .ZN(carry[12]) );
  XOR2_X1 U70 ( .A(B[12]), .B(A[12]), .Z(n56) );
  XOR2_X1 U71 ( .A(n10), .B(n56), .Z(SUM[12]) );
  NAND2_X1 U72 ( .A1(n51), .A2(B[12]), .ZN(n57) );
  NAND2_X1 U73 ( .A1(carry[12]), .A2(A[12]), .ZN(n58) );
  NAND2_X1 U74 ( .A1(B[12]), .A2(A[12]), .ZN(n59) );
  NAND3_X1 U75 ( .A1(n57), .A2(n58), .A3(n59), .ZN(carry[13]) );
  NAND3_X1 U76 ( .A1(n79), .A2(n77), .A3(n78), .ZN(n60) );
  NAND3_X1 U77 ( .A1(n75), .A2(n74), .A3(n73), .ZN(n61) );
  NAND3_X1 U78 ( .A1(n73), .A2(n33), .A3(n30), .ZN(n62) );
  XOR2_X1 U79 ( .A(B[9]), .B(A[9]), .Z(n63) );
  XOR2_X1 U80 ( .A(n29), .B(n63), .Z(SUM[9]) );
  NAND2_X1 U81 ( .A1(carry[9]), .A2(B[9]), .ZN(n64) );
  NAND2_X1 U82 ( .A1(n60), .A2(A[9]), .ZN(n65) );
  NAND2_X1 U83 ( .A1(B[9]), .A2(A[9]), .ZN(n66) );
  NAND3_X1 U84 ( .A1(n64), .A2(n65), .A3(n66), .ZN(carry[10]) );
  CLKBUF_X1 U85 ( .A(n42), .Z(n67) );
  XOR2_X1 U86 ( .A(B[13]), .B(A[13]), .Z(n68) );
  XOR2_X1 U87 ( .A(n67), .B(n68), .Z(SUM[13]) );
  NAND2_X1 U88 ( .A1(B[13]), .A2(n42), .ZN(n69) );
  NAND2_X1 U89 ( .A1(carry[13]), .A2(A[13]), .ZN(n70) );
  NAND2_X1 U90 ( .A1(B[13]), .A2(A[13]), .ZN(n71) );
  NAND3_X1 U91 ( .A1(n69), .A2(n70), .A3(n71), .ZN(carry[14]) );
  XOR2_X1 U92 ( .A(A[7]), .B(B[7]), .Z(n72) );
  XOR2_X1 U93 ( .A(n72), .B(n41), .Z(SUM[7]) );
  NAND2_X1 U94 ( .A1(B[7]), .A2(A[7]), .ZN(n73) );
  NAND2_X1 U95 ( .A1(n28), .A2(A[7]), .ZN(n74) );
  NAND2_X1 U96 ( .A1(B[7]), .A2(n11), .ZN(n75) );
  NAND3_X1 U97 ( .A1(n75), .A2(n73), .A3(n74), .ZN(carry[8]) );
  XOR2_X1 U98 ( .A(A[8]), .B(B[8]), .Z(n76) );
  XOR2_X1 U99 ( .A(n76), .B(n62), .Z(SUM[8]) );
  NAND2_X1 U100 ( .A1(A[8]), .A2(B[8]), .ZN(n77) );
  NAND2_X1 U101 ( .A1(n61), .A2(A[8]), .ZN(n78) );
  NAND2_X1 U102 ( .A1(carry[8]), .A2(B[8]), .ZN(n79) );
  NAND3_X1 U103 ( .A1(n77), .A2(n78), .A3(n79), .ZN(carry[9]) );
  XNOR2_X1 U104 ( .A(carry[15]), .B(n80), .ZN(SUM[15]) );
  XOR2_X1 U105 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U106 ( .A1(B[0]), .A2(A[0]), .ZN(n82) );
endmodule


module datapath_DW_mult_tc_4 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350;

  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n293), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n292), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n296), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n295), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n298), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  BUF_X2 U157 ( .A(a[1]), .Z(n280) );
  AND2_X1 U158 ( .A1(n95), .A2(n102), .ZN(n206) );
  AND3_X1 U159 ( .A1(n276), .A2(n277), .A3(n278), .ZN(product[15]) );
  XNOR2_X1 U160 ( .A(a[6]), .B(a[5]), .ZN(n327) );
  NAND3_X1 U161 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n208) );
  CLKBUF_X1 U162 ( .A(b[3]), .Z(n260) );
  CLKBUF_X1 U163 ( .A(n52), .Z(n209) );
  NAND3_X1 U164 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n210) );
  NAND3_X1 U165 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n211) );
  XNOR2_X1 U166 ( .A(n212), .B(n2), .ZN(product[14]) );
  XNOR2_X1 U167 ( .A(n290), .B(n15), .ZN(n212) );
  NAND3_X1 U168 ( .A1(n226), .A2(n227), .A3(n228), .ZN(n213) );
  NAND3_X1 U169 ( .A1(n226), .A2(n227), .A3(n228), .ZN(n214) );
  CLKBUF_X1 U170 ( .A(b[1]), .Z(n215) );
  CLKBUF_X1 U171 ( .A(n12), .Z(n216) );
  NAND3_X1 U172 ( .A1(n270), .A2(n269), .A3(n271), .ZN(n217) );
  NAND3_X1 U173 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n218) );
  XNOR2_X1 U174 ( .A(n216), .B(n219), .ZN(product[4]) );
  XNOR2_X1 U175 ( .A(n54), .B(n206), .ZN(n219) );
  XNOR2_X1 U176 ( .A(n220), .B(n224), .ZN(product[5]) );
  XNOR2_X1 U177 ( .A(n50), .B(n53), .ZN(n220) );
  INV_X1 U178 ( .A(n299), .ZN(n221) );
  CLKBUF_X1 U179 ( .A(n347), .Z(n231) );
  NAND3_X1 U180 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n222) );
  NAND3_X1 U181 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n223) );
  NAND3_X1 U182 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n224) );
  NAND2_X2 U183 ( .A1(n327), .A2(n346), .ZN(n329) );
  XOR2_X1 U184 ( .A(a[3]), .B(a[2]), .Z(n344) );
  XOR2_X1 U185 ( .A(n27), .B(n24), .Z(n225) );
  XOR2_X1 U186 ( .A(n211), .B(n225), .Z(product[10]) );
  NAND2_X1 U187 ( .A1(n210), .A2(n27), .ZN(n226) );
  NAND2_X1 U188 ( .A1(n6), .A2(n24), .ZN(n227) );
  NAND2_X1 U189 ( .A1(n27), .A2(n24), .ZN(n228) );
  NAND3_X1 U190 ( .A1(n226), .A2(n227), .A3(n228), .ZN(n5) );
  NAND3_X1 U191 ( .A1(n262), .A2(n261), .A3(n263), .ZN(n229) );
  NAND3_X1 U192 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n230) );
  XNOR2_X1 U193 ( .A(n14), .B(n232), .ZN(product[2]) );
  XNOR2_X1 U194 ( .A(n103), .B(n96), .ZN(n232) );
  NAND2_X2 U195 ( .A1(n316), .A2(n345), .ZN(n318) );
  XOR2_X1 U196 ( .A(a[3]), .B(n288), .Z(n307) );
  NAND2_X1 U197 ( .A1(n12), .A2(n54), .ZN(n233) );
  NAND2_X1 U198 ( .A1(n12), .A2(n206), .ZN(n234) );
  NAND2_X1 U199 ( .A1(n54), .A2(n206), .ZN(n235) );
  NAND3_X1 U200 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n11) );
  BUF_X1 U201 ( .A(n288), .Z(n236) );
  XOR2_X1 U202 ( .A(n18), .B(n19), .Z(n237) );
  XOR2_X1 U203 ( .A(n218), .B(n237), .Z(product[12]) );
  NAND2_X1 U204 ( .A1(n217), .A2(n18), .ZN(n238) );
  NAND2_X1 U205 ( .A1(n217), .A2(n19), .ZN(n239) );
  NAND2_X1 U206 ( .A1(n18), .A2(n19), .ZN(n240) );
  NAND3_X1 U207 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n3) );
  NAND3_X1 U208 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n241) );
  NAND3_X1 U209 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n242) );
  NAND2_X1 U210 ( .A1(n14), .A2(n103), .ZN(n243) );
  NAND2_X1 U211 ( .A1(n14), .A2(n96), .ZN(n244) );
  NAND2_X1 U212 ( .A1(n103), .A2(n96), .ZN(n245) );
  NAND3_X1 U213 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n13) );
  XOR2_X1 U214 ( .A(n34), .B(n39), .Z(n246) );
  XOR2_X1 U215 ( .A(n241), .B(n246), .Z(product[8]) );
  NAND2_X1 U216 ( .A1(n241), .A2(n34), .ZN(n247) );
  NAND2_X1 U217 ( .A1(n8), .A2(n39), .ZN(n248) );
  NAND2_X1 U218 ( .A1(n34), .A2(n39), .ZN(n249) );
  NAND3_X1 U219 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n7) );
  NAND3_X1 U220 ( .A1(n265), .A2(n266), .A3(n267), .ZN(n250) );
  XOR2_X1 U221 ( .A(n40), .B(n45), .Z(n251) );
  XOR2_X1 U222 ( .A(n250), .B(n251), .Z(product[7]) );
  NAND2_X1 U223 ( .A1(n250), .A2(n40), .ZN(n252) );
  NAND2_X1 U224 ( .A1(n9), .A2(n45), .ZN(n253) );
  NAND2_X1 U225 ( .A1(n40), .A2(n45), .ZN(n254) );
  NAND3_X1 U226 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n8) );
  XOR2_X1 U227 ( .A(n33), .B(n28), .Z(n255) );
  XOR2_X1 U228 ( .A(n242), .B(n255), .Z(product[9]) );
  NAND2_X1 U229 ( .A1(n242), .A2(n33), .ZN(n256) );
  NAND2_X1 U230 ( .A1(n7), .A2(n28), .ZN(n257) );
  NAND2_X1 U231 ( .A1(n33), .A2(n28), .ZN(n258) );
  NAND3_X1 U232 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n6) );
  XNOR2_X1 U233 ( .A(b[3]), .B(n280), .ZN(n259) );
  XOR2_X1 U234 ( .A(n95), .B(n102), .Z(n56) );
  XNOR2_X2 U235 ( .A(a[2]), .B(a[1]), .ZN(n306) );
  NAND2_X1 U236 ( .A1(n50), .A2(n53), .ZN(n261) );
  NAND2_X1 U237 ( .A1(n50), .A2(n223), .ZN(n262) );
  NAND2_X1 U238 ( .A1(n53), .A2(n11), .ZN(n263) );
  NAND3_X1 U239 ( .A1(n263), .A2(n262), .A3(n261), .ZN(n10) );
  XOR2_X1 U240 ( .A(n46), .B(n49), .Z(n264) );
  XOR2_X1 U241 ( .A(n264), .B(n230), .Z(product[6]) );
  NAND2_X1 U242 ( .A1(n46), .A2(n49), .ZN(n265) );
  NAND2_X1 U243 ( .A1(n46), .A2(n229), .ZN(n266) );
  NAND2_X1 U244 ( .A1(n49), .A2(n10), .ZN(n267) );
  NAND3_X1 U245 ( .A1(n265), .A2(n266), .A3(n267), .ZN(n9) );
  XOR2_X1 U246 ( .A(n23), .B(n20), .Z(n268) );
  XOR2_X1 U247 ( .A(n214), .B(n268), .Z(product[11]) );
  NAND2_X1 U248 ( .A1(n5), .A2(n23), .ZN(n269) );
  NAND2_X1 U249 ( .A1(n213), .A2(n20), .ZN(n270) );
  NAND2_X1 U250 ( .A1(n23), .A2(n20), .ZN(n271) );
  XOR2_X1 U251 ( .A(n17), .B(n289), .Z(n272) );
  XOR2_X1 U252 ( .A(n272), .B(n222), .Z(product[13]) );
  NAND2_X1 U253 ( .A1(n17), .A2(n289), .ZN(n273) );
  NAND2_X1 U254 ( .A1(n17), .A2(n3), .ZN(n274) );
  NAND2_X1 U255 ( .A1(n289), .A2(n3), .ZN(n275) );
  NAND3_X1 U256 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n2) );
  NAND2_X1 U257 ( .A1(n290), .A2(n15), .ZN(n276) );
  NAND2_X1 U258 ( .A1(n290), .A2(n208), .ZN(n277) );
  NAND2_X1 U259 ( .A1(n15), .A2(n208), .ZN(n278) );
  INV_X1 U260 ( .A(n288), .ZN(n279) );
  XNOR2_X2 U261 ( .A(a[4]), .B(a[3]), .ZN(n316) );
  XNOR2_X1 U262 ( .A(n52), .B(n281), .ZN(n50) );
  XNOR2_X1 U263 ( .A(n93), .B(n100), .ZN(n281) );
  INV_X1 U264 ( .A(n15), .ZN(n289) );
  INV_X1 U265 ( .A(n31), .ZN(n295) );
  INV_X1 U266 ( .A(n21), .ZN(n292) );
  INV_X1 U267 ( .A(n325), .ZN(n293) );
  INV_X1 U268 ( .A(n336), .ZN(n290) );
  INV_X1 U269 ( .A(n305), .ZN(n298) );
  INV_X1 U270 ( .A(n314), .ZN(n296) );
  INV_X1 U271 ( .A(a[5]), .ZN(n294) );
  INV_X1 U272 ( .A(a[7]), .ZN(n291) );
  INV_X1 U273 ( .A(a[1]), .ZN(n299) );
  INV_X1 U274 ( .A(b[0]), .ZN(n288) );
  NAND2_X1 U275 ( .A1(n209), .A2(n93), .ZN(n282) );
  NAND2_X1 U276 ( .A1(n209), .A2(n100), .ZN(n283) );
  NAND2_X1 U277 ( .A1(n93), .A2(n100), .ZN(n284) );
  NAND3_X1 U278 ( .A1(n282), .A2(n283), .A3(n284), .ZN(n49) );
  INV_X1 U279 ( .A(a[3]), .ZN(n297) );
  NAND2_X1 U280 ( .A1(n306), .A2(n344), .ZN(n285) );
  NAND2_X1 U281 ( .A1(n306), .A2(n344), .ZN(n286) );
  NAND2_X1 U282 ( .A1(n344), .A2(n306), .ZN(n308) );
  INV_X1 U283 ( .A(n288), .ZN(n287) );
  INV_X2 U284 ( .A(a[0]), .ZN(n300) );
  NOR2_X1 U285 ( .A1(n300), .A2(n236), .ZN(product[0]) );
  OAI22_X1 U286 ( .A1(n301), .A2(n302), .B1(n303), .B2(n300), .ZN(n99) );
  OAI22_X1 U287 ( .A1(n303), .A2(n302), .B1(n304), .B2(n300), .ZN(n98) );
  XNOR2_X1 U288 ( .A(b[6]), .B(n280), .ZN(n303) );
  OAI22_X1 U289 ( .A1(n300), .A2(n304), .B1(n302), .B2(n304), .ZN(n305) );
  XNOR2_X1 U290 ( .A(b[7]), .B(n280), .ZN(n304) );
  NOR2_X1 U291 ( .A1(n306), .A2(n236), .ZN(n96) );
  OAI22_X1 U292 ( .A1(n307), .A2(n308), .B1(n306), .B2(n309), .ZN(n95) );
  OAI22_X1 U293 ( .A1(n309), .A2(n285), .B1(n306), .B2(n310), .ZN(n94) );
  XNOR2_X1 U294 ( .A(b[1]), .B(a[3]), .ZN(n309) );
  OAI22_X1 U295 ( .A1(n310), .A2(n286), .B1(n306), .B2(n311), .ZN(n93) );
  XNOR2_X1 U296 ( .A(b[2]), .B(a[3]), .ZN(n310) );
  OAI22_X1 U297 ( .A1(n311), .A2(n285), .B1(n306), .B2(n312), .ZN(n92) );
  XNOR2_X1 U298 ( .A(n260), .B(a[3]), .ZN(n311) );
  OAI22_X1 U299 ( .A1(n312), .A2(n285), .B1(n306), .B2(n313), .ZN(n91) );
  XNOR2_X1 U300 ( .A(b[4]), .B(a[3]), .ZN(n312) );
  OAI22_X1 U301 ( .A1(n315), .A2(n306), .B1(n285), .B2(n315), .ZN(n314) );
  NOR2_X1 U302 ( .A1(n316), .A2(n236), .ZN(n88) );
  OAI22_X1 U303 ( .A1(n317), .A2(n318), .B1(n316), .B2(n319), .ZN(n87) );
  XNOR2_X1 U304 ( .A(a[5]), .B(n279), .ZN(n317) );
  OAI22_X1 U305 ( .A1(n319), .A2(n318), .B1(n316), .B2(n320), .ZN(n86) );
  XNOR2_X1 U306 ( .A(n215), .B(a[5]), .ZN(n319) );
  OAI22_X1 U307 ( .A1(n320), .A2(n318), .B1(n316), .B2(n321), .ZN(n85) );
  XNOR2_X1 U308 ( .A(b[2]), .B(a[5]), .ZN(n320) );
  OAI22_X1 U309 ( .A1(n321), .A2(n318), .B1(n316), .B2(n322), .ZN(n84) );
  XNOR2_X1 U310 ( .A(n260), .B(a[5]), .ZN(n321) );
  OAI22_X1 U311 ( .A1(n322), .A2(n318), .B1(n316), .B2(n323), .ZN(n83) );
  XNOR2_X1 U312 ( .A(b[4]), .B(a[5]), .ZN(n322) );
  OAI22_X1 U313 ( .A1(n323), .A2(n318), .B1(n316), .B2(n324), .ZN(n82) );
  XNOR2_X1 U314 ( .A(b[5]), .B(a[5]), .ZN(n323) );
  OAI22_X1 U315 ( .A1(n326), .A2(n316), .B1(n318), .B2(n326), .ZN(n325) );
  NOR2_X1 U316 ( .A1(n327), .A2(n236), .ZN(n80) );
  OAI22_X1 U317 ( .A1(n328), .A2(n329), .B1(n327), .B2(n330), .ZN(n79) );
  XNOR2_X1 U318 ( .A(a[7]), .B(n279), .ZN(n328) );
  OAI22_X1 U319 ( .A1(n331), .A2(n329), .B1(n327), .B2(n332), .ZN(n77) );
  OAI22_X1 U320 ( .A1(n332), .A2(n329), .B1(n327), .B2(n333), .ZN(n76) );
  XNOR2_X1 U321 ( .A(b[3]), .B(a[7]), .ZN(n332) );
  OAI22_X1 U322 ( .A1(n333), .A2(n329), .B1(n327), .B2(n334), .ZN(n75) );
  XNOR2_X1 U323 ( .A(b[4]), .B(a[7]), .ZN(n333) );
  OAI22_X1 U324 ( .A1(n334), .A2(n329), .B1(n327), .B2(n335), .ZN(n74) );
  XNOR2_X1 U325 ( .A(b[5]), .B(a[7]), .ZN(n334) );
  OAI22_X1 U326 ( .A1(n337), .A2(n327), .B1(n329), .B2(n337), .ZN(n336) );
  OAI21_X1 U327 ( .B1(n287), .B2(n299), .A(n302), .ZN(n72) );
  OAI21_X1 U328 ( .B1(n297), .B2(n286), .A(n338), .ZN(n71) );
  OR3_X1 U329 ( .A1(n306), .A2(n279), .A3(n297), .ZN(n338) );
  OAI21_X1 U330 ( .B1(n294), .B2(n318), .A(n339), .ZN(n70) );
  OR3_X1 U331 ( .A1(n316), .A2(n279), .A3(n294), .ZN(n339) );
  OAI21_X1 U332 ( .B1(n291), .B2(n329), .A(n340), .ZN(n69) );
  OR3_X1 U333 ( .A1(n327), .A2(n279), .A3(n291), .ZN(n340) );
  XNOR2_X1 U334 ( .A(n341), .B(n342), .ZN(n38) );
  OR2_X1 U335 ( .A1(n341), .A2(n342), .ZN(n37) );
  OAI22_X1 U336 ( .A1(n313), .A2(n286), .B1(n306), .B2(n343), .ZN(n342) );
  XNOR2_X1 U337 ( .A(b[5]), .B(a[3]), .ZN(n313) );
  OAI22_X1 U338 ( .A1(n330), .A2(n329), .B1(n327), .B2(n331), .ZN(n341) );
  XNOR2_X1 U339 ( .A(b[2]), .B(a[7]), .ZN(n331) );
  XNOR2_X1 U340 ( .A(n215), .B(a[7]), .ZN(n330) );
  OAI22_X1 U341 ( .A1(n343), .A2(n286), .B1(n306), .B2(n315), .ZN(n31) );
  XNOR2_X1 U342 ( .A(b[7]), .B(a[3]), .ZN(n315) );
  XNOR2_X1 U343 ( .A(b[6]), .B(a[3]), .ZN(n343) );
  OAI22_X1 U344 ( .A1(n324), .A2(n318), .B1(n316), .B2(n326), .ZN(n21) );
  XNOR2_X1 U345 ( .A(b[7]), .B(a[5]), .ZN(n326) );
  XNOR2_X1 U346 ( .A(n294), .B(a[4]), .ZN(n345) );
  XNOR2_X1 U347 ( .A(b[6]), .B(a[5]), .ZN(n324) );
  OAI22_X1 U348 ( .A1(n335), .A2(n329), .B1(n327), .B2(n337), .ZN(n15) );
  XNOR2_X1 U349 ( .A(b[7]), .B(a[7]), .ZN(n337) );
  XNOR2_X1 U350 ( .A(n291), .B(a[6]), .ZN(n346) );
  XNOR2_X1 U351 ( .A(b[6]), .B(a[7]), .ZN(n335) );
  OAI22_X1 U352 ( .A1(n287), .A2(n302), .B1(n347), .B2(n300), .ZN(n104) );
  OAI22_X1 U353 ( .A1(n231), .A2(n302), .B1(n348), .B2(n300), .ZN(n103) );
  XNOR2_X1 U354 ( .A(b[1]), .B(n221), .ZN(n347) );
  OAI22_X1 U355 ( .A1(n348), .A2(n302), .B1(n349), .B2(n300), .ZN(n102) );
  XNOR2_X1 U356 ( .A(b[2]), .B(n280), .ZN(n348) );
  OAI22_X1 U357 ( .A1(n259), .A2(n302), .B1(n350), .B2(n300), .ZN(n101) );
  XNOR2_X1 U358 ( .A(b[3]), .B(n280), .ZN(n349) );
  OAI22_X1 U359 ( .A1(n350), .A2(n302), .B1(n301), .B2(n300), .ZN(n100) );
  XNOR2_X1 U360 ( .A(b[5]), .B(n280), .ZN(n301) );
  NAND2_X1 U361 ( .A1(a[1]), .A2(n300), .ZN(n302) );
  XNOR2_X1 U362 ( .A(b[4]), .B(n280), .ZN(n350) );
endmodule


module datapath_DW01_add_4 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n83;
  wire   [15:1] carry;

  INV_X1 U1 ( .A(A[14]), .ZN(n2) );
  CLKBUF_X1 U2 ( .A(n52), .Z(n1) );
  XNOR2_X1 U3 ( .A(B[14]), .B(n2), .ZN(n3) );
  XOR2_X1 U4 ( .A(n3), .B(carry[14]), .Z(SUM[14]) );
  NAND2_X1 U5 ( .A1(carry[14]), .A2(B[14]), .ZN(n4) );
  NAND2_X1 U6 ( .A1(carry[14]), .A2(A[14]), .ZN(n5) );
  NAND2_X1 U7 ( .A1(B[14]), .A2(A[14]), .ZN(n6) );
  NAND3_X1 U8 ( .A1(n4), .A2(n5), .A3(n6), .ZN(carry[15]) );
  NAND3_X1 U9 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n7) );
  CLKBUF_X1 U10 ( .A(n34), .Z(n8) );
  NAND3_X1 U11 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n9) );
  NAND3_X1 U12 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n10) );
  CLKBUF_X1 U13 ( .A(n70), .Z(n11) );
  NAND3_X1 U14 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n12) );
  XOR2_X1 U15 ( .A(B[7]), .B(A[7]), .Z(n13) );
  XOR2_X1 U16 ( .A(n10), .B(n13), .Z(SUM[7]) );
  NAND2_X1 U17 ( .A1(n9), .A2(B[7]), .ZN(n14) );
  NAND2_X1 U18 ( .A1(carry[7]), .A2(A[7]), .ZN(n15) );
  NAND2_X1 U19 ( .A1(B[7]), .A2(A[7]), .ZN(n16) );
  NAND3_X1 U20 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[8]) );
  NAND3_X1 U21 ( .A1(n11), .A2(n71), .A3(n72), .ZN(n17) );
  NAND3_X1 U22 ( .A1(n77), .A2(n76), .A3(n75), .ZN(n18) );
  NAND3_X1 U23 ( .A1(n1), .A2(n53), .A3(n54), .ZN(n19) );
  XOR2_X1 U24 ( .A(n83), .B(A[1]), .Z(n20) );
  XOR2_X1 U25 ( .A(B[1]), .B(n20), .Z(SUM[1]) );
  NAND2_X1 U26 ( .A1(B[1]), .A2(n83), .ZN(n21) );
  NAND2_X1 U27 ( .A1(B[1]), .A2(A[1]), .ZN(n22) );
  NAND2_X1 U28 ( .A1(n83), .A2(A[1]), .ZN(n23) );
  NAND3_X1 U29 ( .A1(n21), .A2(n22), .A3(n23), .ZN(carry[2]) );
  NAND3_X1 U30 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n24) );
  CLKBUF_X1 U31 ( .A(n33), .Z(n25) );
  XOR2_X1 U32 ( .A(B[11]), .B(A[11]), .Z(n26) );
  XOR2_X1 U33 ( .A(n17), .B(n26), .Z(SUM[11]) );
  NAND2_X1 U34 ( .A1(carry[11]), .A2(B[11]), .ZN(n27) );
  NAND2_X1 U35 ( .A1(carry[11]), .A2(A[11]), .ZN(n28) );
  NAND2_X1 U36 ( .A1(B[11]), .A2(A[11]), .ZN(n29) );
  NAND3_X1 U37 ( .A1(n28), .A2(n27), .A3(n29), .ZN(carry[12]) );
  NAND3_X1 U38 ( .A1(n58), .A2(n57), .A3(n59), .ZN(n30) );
  CLKBUF_X1 U39 ( .A(n12), .Z(n31) );
  NAND3_X1 U40 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n32) );
  NAND3_X1 U41 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n33) );
  NAND3_X1 U42 ( .A1(n77), .A2(n76), .A3(n75), .ZN(n34) );
  NAND3_X1 U43 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n35) );
  NAND3_X1 U44 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n36) );
  NAND3_X1 U45 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n37) );
  XOR2_X1 U46 ( .A(B[2]), .B(A[2]), .Z(n38) );
  XOR2_X1 U47 ( .A(n38), .B(carry[2]), .Z(SUM[2]) );
  NAND2_X1 U48 ( .A1(B[2]), .A2(A[2]), .ZN(n39) );
  NAND2_X1 U49 ( .A1(B[2]), .A2(carry[2]), .ZN(n40) );
  NAND2_X1 U50 ( .A1(A[2]), .A2(carry[2]), .ZN(n41) );
  NAND3_X1 U51 ( .A1(n39), .A2(n40), .A3(n41), .ZN(carry[3]) );
  XOR2_X1 U52 ( .A(A[3]), .B(B[3]), .Z(n42) );
  XOR2_X1 U53 ( .A(n42), .B(n37), .Z(SUM[3]) );
  NAND2_X1 U54 ( .A1(A[3]), .A2(B[3]), .ZN(n43) );
  NAND2_X1 U55 ( .A1(A[3]), .A2(n36), .ZN(n44) );
  NAND2_X1 U56 ( .A1(B[3]), .A2(carry[3]), .ZN(n45) );
  NAND3_X1 U57 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[4]) );
  XOR2_X1 U58 ( .A(B[9]), .B(A[9]), .Z(n46) );
  XOR2_X1 U59 ( .A(n25), .B(n46), .Z(SUM[9]) );
  NAND2_X1 U60 ( .A1(n33), .A2(B[9]), .ZN(n47) );
  NAND2_X1 U61 ( .A1(carry[9]), .A2(A[9]), .ZN(n48) );
  NAND2_X1 U62 ( .A1(B[9]), .A2(A[9]), .ZN(n49) );
  NAND3_X1 U63 ( .A1(n47), .A2(n48), .A3(n49), .ZN(carry[10]) );
  NAND3_X1 U64 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n50) );
  XOR2_X1 U65 ( .A(B[4]), .B(A[4]), .Z(n51) );
  XOR2_X1 U66 ( .A(n35), .B(n51), .Z(SUM[4]) );
  NAND2_X1 U67 ( .A1(n35), .A2(B[4]), .ZN(n52) );
  NAND2_X1 U68 ( .A1(carry[4]), .A2(A[4]), .ZN(n53) );
  NAND2_X1 U69 ( .A1(B[4]), .A2(A[4]), .ZN(n54) );
  CLKBUF_X1 U70 ( .A(n30), .Z(n55) );
  XOR2_X1 U71 ( .A(B[5]), .B(A[5]), .Z(n56) );
  XOR2_X1 U72 ( .A(n19), .B(n56), .Z(SUM[5]) );
  NAND2_X1 U73 ( .A1(n50), .A2(B[5]), .ZN(n57) );
  NAND2_X1 U74 ( .A1(n32), .A2(A[5]), .ZN(n58) );
  NAND2_X1 U75 ( .A1(B[5]), .A2(A[5]), .ZN(n59) );
  NAND3_X1 U76 ( .A1(n57), .A2(n58), .A3(n59), .ZN(carry[6]) );
  XOR2_X1 U77 ( .A(B[6]), .B(A[6]), .Z(n60) );
  XOR2_X1 U78 ( .A(n55), .B(n60), .Z(SUM[6]) );
  NAND2_X1 U79 ( .A1(n30), .A2(B[6]), .ZN(n61) );
  NAND2_X1 U80 ( .A1(carry[6]), .A2(A[6]), .ZN(n62) );
  NAND2_X1 U81 ( .A1(B[6]), .A2(A[6]), .ZN(n63) );
  NAND3_X1 U82 ( .A1(n61), .A2(n62), .A3(n63), .ZN(carry[7]) );
  XOR2_X1 U83 ( .A(B[8]), .B(A[8]), .Z(n64) );
  XOR2_X1 U84 ( .A(carry[8]), .B(n64), .Z(SUM[8]) );
  NAND2_X1 U85 ( .A1(n7), .A2(B[8]), .ZN(n65) );
  NAND2_X1 U86 ( .A1(n7), .A2(A[8]), .ZN(n66) );
  NAND2_X1 U87 ( .A1(B[8]), .A2(A[8]), .ZN(n67) );
  NAND3_X1 U88 ( .A1(n66), .A2(n65), .A3(n67), .ZN(carry[9]) );
  CLKBUF_X1 U89 ( .A(n24), .Z(n68) );
  XOR2_X1 U90 ( .A(B[10]), .B(A[10]), .Z(n69) );
  XOR2_X1 U91 ( .A(n68), .B(n69), .Z(SUM[10]) );
  NAND2_X1 U92 ( .A1(n24), .A2(B[10]), .ZN(n70) );
  NAND2_X1 U93 ( .A1(carry[10]), .A2(A[10]), .ZN(n71) );
  NAND2_X1 U94 ( .A1(B[10]), .A2(A[10]), .ZN(n72) );
  NAND3_X1 U95 ( .A1(n70), .A2(n71), .A3(n72), .ZN(carry[11]) );
  NAND2_X1 U96 ( .A1(A[12]), .A2(B[12]), .ZN(n75) );
  XNOR2_X1 U97 ( .A(carry[15]), .B(n73), .ZN(SUM[15]) );
  XNOR2_X1 U98 ( .A(B[15]), .B(A[15]), .ZN(n73) );
  XOR2_X1 U99 ( .A(A[12]), .B(B[12]), .Z(n74) );
  XOR2_X1 U100 ( .A(n74), .B(n31), .Z(SUM[12]) );
  NAND2_X1 U101 ( .A1(A[12]), .A2(carry[12]), .ZN(n76) );
  NAND2_X1 U102 ( .A1(B[12]), .A2(n12), .ZN(n77) );
  XOR2_X1 U103 ( .A(A[13]), .B(B[13]), .Z(n78) );
  XOR2_X1 U104 ( .A(n78), .B(n8), .Z(SUM[13]) );
  NAND2_X1 U105 ( .A1(B[13]), .A2(A[13]), .ZN(n79) );
  NAND2_X1 U106 ( .A1(A[13]), .A2(n34), .ZN(n80) );
  NAND2_X1 U107 ( .A1(B[13]), .A2(n18), .ZN(n81) );
  NAND3_X1 U108 ( .A1(n80), .A2(n81), .A3(n79), .ZN(carry[14]) );
  XOR2_X1 U109 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U110 ( .A1(B[0]), .A2(A[0]), .ZN(n83) );
endmodule


module datapath_DW_mult_tc_3 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n7, n9, n10, n11, n12, n13, n14, n15, n17, n18, n19,
         n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76, n77,
         n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94, n95,
         n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349;

  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n292), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n291), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n295), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n294), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n297), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  AND2_X1 U157 ( .A1(n268), .A2(n102), .ZN(n206) );
  XNOR2_X1 U158 ( .A(n289), .B(n15), .ZN(n207) );
  AND3_X1 U159 ( .A1(n265), .A2(n266), .A3(n267), .ZN(product[15]) );
  XNOR2_X1 U160 ( .A(n242), .B(n209), .ZN(product[13]) );
  AND3_X1 U161 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n209) );
  XNOR2_X1 U162 ( .A(n238), .B(n210), .ZN(product[12]) );
  AND3_X1 U163 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n210) );
  XNOR2_X1 U164 ( .A(b[2]), .B(a[1]), .ZN(n347) );
  NAND3_X1 U165 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n211) );
  NAND3_X1 U166 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n212) );
  NAND2_X2 U167 ( .A1(n326), .A2(n345), .ZN(n328) );
  XNOR2_X1 U168 ( .A(n218), .B(n213), .ZN(product[4]) );
  XNOR2_X1 U169 ( .A(n54), .B(n206), .ZN(n213) );
  XNOR2_X1 U170 ( .A(n13), .B(n214), .ZN(product[3]) );
  XNOR2_X1 U171 ( .A(n56), .B(n71), .ZN(n214) );
  NAND3_X1 U172 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n215) );
  NAND3_X1 U173 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n216) );
  OAI22_X1 U174 ( .A1(n306), .A2(n307), .B1(n305), .B2(n308), .ZN(n217) );
  NAND3_X1 U175 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n218) );
  XOR2_X1 U176 ( .A(n217), .B(n102), .Z(n219) );
  NAND3_X1 U177 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n220) );
  NAND3_X1 U178 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n221) );
  NAND3_X1 U179 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n222) );
  NAND3_X1 U180 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n223) );
  XOR2_X1 U181 ( .A(n23), .B(n20), .Z(n224) );
  XOR2_X1 U182 ( .A(n221), .B(n224), .Z(product[11]) );
  NAND2_X1 U183 ( .A1(n5), .A2(n23), .ZN(n225) );
  NAND2_X1 U184 ( .A1(n5), .A2(n20), .ZN(n226) );
  NAND2_X1 U185 ( .A1(n23), .A2(n20), .ZN(n227) );
  NAND3_X1 U186 ( .A1(n226), .A2(n225), .A3(n227), .ZN(n4) );
  CLKBUF_X1 U187 ( .A(b[1]), .Z(n228) );
  NAND2_X1 U188 ( .A1(n13), .A2(n219), .ZN(n229) );
  NAND2_X1 U189 ( .A1(n13), .A2(n71), .ZN(n230) );
  NAND2_X1 U190 ( .A1(n219), .A2(n71), .ZN(n231) );
  NAND3_X1 U191 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n12) );
  NAND3_X1 U192 ( .A1(n234), .A2(n235), .A3(n236), .ZN(n232) );
  XNOR2_X1 U193 ( .A(a[4]), .B(a[3]), .ZN(n233) );
  XNOR2_X1 U194 ( .A(a[4]), .B(a[3]), .ZN(n315) );
  NAND2_X1 U195 ( .A1(n218), .A2(n54), .ZN(n234) );
  NAND2_X1 U196 ( .A1(n12), .A2(n206), .ZN(n235) );
  NAND2_X1 U197 ( .A1(n54), .A2(n206), .ZN(n236) );
  NAND3_X1 U198 ( .A1(n234), .A2(n235), .A3(n236), .ZN(n11) );
  BUF_X1 U199 ( .A(n287), .Z(n237) );
  XOR2_X1 U200 ( .A(n19), .B(n18), .Z(n238) );
  NAND2_X1 U201 ( .A1(n19), .A2(n18), .ZN(n239) );
  NAND2_X1 U202 ( .A1(n19), .A2(n222), .ZN(n240) );
  NAND2_X1 U203 ( .A1(n18), .A2(n4), .ZN(n241) );
  NAND3_X1 U204 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n3) );
  XOR2_X1 U205 ( .A(n17), .B(n288), .Z(n242) );
  NAND2_X1 U206 ( .A1(n17), .A2(n288), .ZN(n243) );
  NAND2_X1 U207 ( .A1(n17), .A2(n223), .ZN(n244) );
  NAND2_X1 U208 ( .A1(n288), .A2(n3), .ZN(n245) );
  NAND3_X1 U209 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n2) );
  XOR2_X1 U210 ( .A(n33), .B(n28), .Z(n246) );
  XOR2_X1 U211 ( .A(n212), .B(n246), .Z(product[9]) );
  NAND2_X1 U212 ( .A1(n211), .A2(n33), .ZN(n247) );
  NAND2_X1 U213 ( .A1(n7), .A2(n28), .ZN(n248) );
  NAND2_X1 U214 ( .A1(n33), .A2(n28), .ZN(n249) );
  NAND3_X1 U215 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n250) );
  INV_X1 U216 ( .A(b[0]), .ZN(n287) );
  CLKBUF_X1 U217 ( .A(n217), .Z(n268) );
  XOR2_X1 U218 ( .A(n27), .B(n24), .Z(n251) );
  XOR2_X1 U219 ( .A(n216), .B(n251), .Z(product[10]) );
  NAND2_X1 U220 ( .A1(n215), .A2(n27), .ZN(n252) );
  NAND2_X1 U221 ( .A1(n215), .A2(n24), .ZN(n253) );
  NAND2_X1 U222 ( .A1(n27), .A2(n24), .ZN(n254) );
  NAND3_X1 U223 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n5) );
  NAND3_X1 U224 ( .A1(n276), .A2(n277), .A3(n275), .ZN(n255) );
  NAND3_X1 U225 ( .A1(n276), .A2(n277), .A3(n275), .ZN(n256) );
  XNOR2_X1 U226 ( .A(n11), .B(n257), .ZN(product[5]) );
  XNOR2_X1 U227 ( .A(n50), .B(n53), .ZN(n257) );
  XOR2_X1 U228 ( .A(n34), .B(n39), .Z(n258) );
  XOR2_X1 U229 ( .A(n256), .B(n258), .Z(product[8]) );
  NAND2_X1 U230 ( .A1(n255), .A2(n34), .ZN(n259) );
  NAND2_X1 U231 ( .A1(n255), .A2(n39), .ZN(n260) );
  NAND2_X1 U232 ( .A1(n34), .A2(n39), .ZN(n261) );
  NAND3_X1 U233 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n7) );
  XNOR2_X1 U234 ( .A(n220), .B(n207), .ZN(product[14]) );
  NAND2_X1 U235 ( .A1(n232), .A2(n50), .ZN(n262) );
  NAND2_X1 U236 ( .A1(n11), .A2(n53), .ZN(n263) );
  NAND2_X1 U237 ( .A1(n50), .A2(n53), .ZN(n264) );
  NAND3_X1 U238 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n10) );
  NAND2_X1 U239 ( .A1(n2), .A2(n289), .ZN(n265) );
  NAND2_X1 U240 ( .A1(n2), .A2(n15), .ZN(n266) );
  NAND2_X1 U241 ( .A1(n289), .A2(n15), .ZN(n267) );
  XOR2_X1 U242 ( .A(n95), .B(n102), .Z(n56) );
  NAND3_X1 U243 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n269) );
  XOR2_X1 U244 ( .A(n46), .B(n49), .Z(n270) );
  XOR2_X1 U245 ( .A(n270), .B(n250), .Z(product[6]) );
  NAND2_X1 U246 ( .A1(n46), .A2(n49), .ZN(n271) );
  NAND2_X1 U247 ( .A1(n46), .A2(n10), .ZN(n272) );
  NAND2_X1 U248 ( .A1(n250), .A2(n49), .ZN(n273) );
  NAND3_X1 U249 ( .A1(n273), .A2(n272), .A3(n271), .ZN(n9) );
  XOR2_X1 U250 ( .A(n40), .B(n45), .Z(n274) );
  XOR2_X1 U251 ( .A(n274), .B(n269), .Z(product[7]) );
  NAND2_X1 U252 ( .A1(n40), .A2(n45), .ZN(n275) );
  NAND2_X1 U253 ( .A1(n9), .A2(n40), .ZN(n276) );
  NAND2_X1 U254 ( .A1(n9), .A2(n45), .ZN(n277) );
  CLKBUF_X1 U255 ( .A(b[3]), .Z(n278) );
  CLKBUF_X1 U256 ( .A(n305), .Z(n279) );
  INV_X2 U257 ( .A(n298), .ZN(n280) );
  INV_X1 U258 ( .A(n287), .ZN(n281) );
  INV_X1 U259 ( .A(n15), .ZN(n288) );
  INV_X1 U260 ( .A(n31), .ZN(n294) );
  INV_X1 U261 ( .A(n21), .ZN(n291) );
  INV_X1 U262 ( .A(n324), .ZN(n292) );
  INV_X1 U263 ( .A(n335), .ZN(n289) );
  INV_X1 U264 ( .A(n304), .ZN(n297) );
  INV_X1 U265 ( .A(n313), .ZN(n295) );
  INV_X1 U266 ( .A(a[5]), .ZN(n293) );
  INV_X1 U267 ( .A(a[7]), .ZN(n290) );
  NAND2_X1 U268 ( .A1(n305), .A2(n343), .ZN(n282) );
  NAND2_X1 U269 ( .A1(a[2]), .A2(a[1]), .ZN(n284) );
  NAND2_X1 U270 ( .A1(n283), .A2(n298), .ZN(n285) );
  NAND2_X2 U271 ( .A1(n284), .A2(n285), .ZN(n305) );
  INV_X1 U272 ( .A(a[2]), .ZN(n283) );
  NAND2_X1 U273 ( .A1(n305), .A2(n343), .ZN(n307) );
  INV_X1 U274 ( .A(a[3]), .ZN(n296) );
  NAND2_X2 U275 ( .A1(n315), .A2(n344), .ZN(n317) );
  INV_X1 U276 ( .A(a[1]), .ZN(n298) );
  XOR2_X2 U277 ( .A(a[6]), .B(n293), .Z(n326) );
  INV_X1 U278 ( .A(n287), .ZN(n286) );
  INV_X2 U279 ( .A(a[0]), .ZN(n299) );
  NOR2_X1 U280 ( .A1(n299), .A2(n237), .ZN(product[0]) );
  OAI22_X1 U281 ( .A1(n300), .A2(n301), .B1(n302), .B2(n299), .ZN(n99) );
  OAI22_X1 U282 ( .A1(n302), .A2(n301), .B1(n303), .B2(n299), .ZN(n98) );
  XNOR2_X1 U283 ( .A(b[6]), .B(n280), .ZN(n302) );
  OAI22_X1 U284 ( .A1(n299), .A2(n303), .B1(n301), .B2(n303), .ZN(n304) );
  XNOR2_X1 U285 ( .A(b[7]), .B(n280), .ZN(n303) );
  NOR2_X1 U286 ( .A1(n305), .A2(n237), .ZN(n96) );
  OAI22_X1 U287 ( .A1(n306), .A2(n307), .B1(n305), .B2(n308), .ZN(n95) );
  XNOR2_X1 U288 ( .A(a[3]), .B(n286), .ZN(n306) );
  OAI22_X1 U289 ( .A1(n308), .A2(n282), .B1(n305), .B2(n309), .ZN(n94) );
  XNOR2_X1 U290 ( .A(b[1]), .B(a[3]), .ZN(n308) );
  OAI22_X1 U291 ( .A1(n309), .A2(n307), .B1(n305), .B2(n310), .ZN(n93) );
  XNOR2_X1 U292 ( .A(b[2]), .B(a[3]), .ZN(n309) );
  OAI22_X1 U293 ( .A1(n310), .A2(n282), .B1(n305), .B2(n311), .ZN(n92) );
  XNOR2_X1 U294 ( .A(b[3]), .B(a[3]), .ZN(n310) );
  OAI22_X1 U295 ( .A1(n311), .A2(n282), .B1(n305), .B2(n312), .ZN(n91) );
  XNOR2_X1 U296 ( .A(b[4]), .B(a[3]), .ZN(n311) );
  OAI22_X1 U297 ( .A1(n314), .A2(n279), .B1(n307), .B2(n314), .ZN(n313) );
  NOR2_X1 U298 ( .A1(n233), .A2(n237), .ZN(n88) );
  OAI22_X1 U299 ( .A1(n316), .A2(n317), .B1(n233), .B2(n318), .ZN(n87) );
  XNOR2_X1 U300 ( .A(a[5]), .B(n281), .ZN(n316) );
  OAI22_X1 U301 ( .A1(n318), .A2(n317), .B1(n233), .B2(n319), .ZN(n86) );
  XNOR2_X1 U302 ( .A(n228), .B(a[5]), .ZN(n318) );
  OAI22_X1 U303 ( .A1(n319), .A2(n317), .B1(n233), .B2(n320), .ZN(n85) );
  XNOR2_X1 U304 ( .A(b[2]), .B(a[5]), .ZN(n319) );
  OAI22_X1 U305 ( .A1(n320), .A2(n317), .B1(n233), .B2(n321), .ZN(n84) );
  XNOR2_X1 U306 ( .A(b[3]), .B(a[5]), .ZN(n320) );
  OAI22_X1 U307 ( .A1(n321), .A2(n317), .B1(n233), .B2(n322), .ZN(n83) );
  XNOR2_X1 U308 ( .A(b[4]), .B(a[5]), .ZN(n321) );
  OAI22_X1 U309 ( .A1(n322), .A2(n317), .B1(n233), .B2(n323), .ZN(n82) );
  XNOR2_X1 U310 ( .A(b[5]), .B(a[5]), .ZN(n322) );
  OAI22_X1 U311 ( .A1(n325), .A2(n233), .B1(n317), .B2(n325), .ZN(n324) );
  NOR2_X1 U312 ( .A1(n326), .A2(n237), .ZN(n80) );
  OAI22_X1 U313 ( .A1(n327), .A2(n328), .B1(n326), .B2(n329), .ZN(n79) );
  XNOR2_X1 U314 ( .A(a[7]), .B(n281), .ZN(n327) );
  OAI22_X1 U315 ( .A1(n330), .A2(n328), .B1(n326), .B2(n331), .ZN(n77) );
  OAI22_X1 U316 ( .A1(n331), .A2(n328), .B1(n326), .B2(n332), .ZN(n76) );
  XNOR2_X1 U317 ( .A(n278), .B(a[7]), .ZN(n331) );
  OAI22_X1 U318 ( .A1(n332), .A2(n328), .B1(n326), .B2(n333), .ZN(n75) );
  XNOR2_X1 U319 ( .A(b[4]), .B(a[7]), .ZN(n332) );
  OAI22_X1 U320 ( .A1(n333), .A2(n328), .B1(n326), .B2(n334), .ZN(n74) );
  XNOR2_X1 U321 ( .A(b[5]), .B(a[7]), .ZN(n333) );
  OAI22_X1 U322 ( .A1(n336), .A2(n326), .B1(n328), .B2(n336), .ZN(n335) );
  OAI21_X1 U323 ( .B1(n286), .B2(n298), .A(n301), .ZN(n72) );
  OAI21_X1 U324 ( .B1(n296), .B2(n307), .A(n337), .ZN(n71) );
  OR3_X1 U325 ( .A1(n305), .A2(n281), .A3(n296), .ZN(n337) );
  OAI21_X1 U326 ( .B1(n293), .B2(n317), .A(n338), .ZN(n70) );
  OR3_X1 U327 ( .A1(n233), .A2(n281), .A3(n293), .ZN(n338) );
  OAI21_X1 U328 ( .B1(n290), .B2(n328), .A(n339), .ZN(n69) );
  OR3_X1 U329 ( .A1(n326), .A2(n281), .A3(n290), .ZN(n339) );
  XNOR2_X1 U330 ( .A(n340), .B(n341), .ZN(n38) );
  OR2_X1 U331 ( .A1(n340), .A2(n341), .ZN(n37) );
  OAI22_X1 U332 ( .A1(n312), .A2(n282), .B1(n279), .B2(n342), .ZN(n341) );
  XNOR2_X1 U333 ( .A(b[5]), .B(a[3]), .ZN(n312) );
  OAI22_X1 U334 ( .A1(n329), .A2(n328), .B1(n326), .B2(n330), .ZN(n340) );
  XNOR2_X1 U335 ( .A(b[2]), .B(a[7]), .ZN(n330) );
  XNOR2_X1 U336 ( .A(n228), .B(a[7]), .ZN(n329) );
  OAI22_X1 U337 ( .A1(n342), .A2(n307), .B1(n279), .B2(n314), .ZN(n31) );
  XNOR2_X1 U338 ( .A(b[7]), .B(a[3]), .ZN(n314) );
  XNOR2_X1 U339 ( .A(n296), .B(a[2]), .ZN(n343) );
  XNOR2_X1 U340 ( .A(b[6]), .B(a[3]), .ZN(n342) );
  OAI22_X1 U341 ( .A1(n323), .A2(n317), .B1(n233), .B2(n325), .ZN(n21) );
  XNOR2_X1 U342 ( .A(b[7]), .B(a[5]), .ZN(n325) );
  XNOR2_X1 U343 ( .A(n293), .B(a[4]), .ZN(n344) );
  XNOR2_X1 U344 ( .A(b[6]), .B(a[5]), .ZN(n323) );
  OAI22_X1 U345 ( .A1(n334), .A2(n328), .B1(n326), .B2(n336), .ZN(n15) );
  XNOR2_X1 U346 ( .A(b[7]), .B(a[7]), .ZN(n336) );
  XNOR2_X1 U347 ( .A(n290), .B(a[6]), .ZN(n345) );
  XNOR2_X1 U348 ( .A(b[6]), .B(a[7]), .ZN(n334) );
  OAI22_X1 U349 ( .A1(n286), .A2(n301), .B1(n346), .B2(n299), .ZN(n104) );
  OAI22_X1 U350 ( .A1(n346), .A2(n301), .B1(n347), .B2(n299), .ZN(n103) );
  XNOR2_X1 U351 ( .A(b[1]), .B(a[1]), .ZN(n346) );
  OAI22_X1 U352 ( .A1(n347), .A2(n301), .B1(n348), .B2(n299), .ZN(n102) );
  OAI22_X1 U353 ( .A1(n348), .A2(n301), .B1(n349), .B2(n299), .ZN(n101) );
  XNOR2_X1 U354 ( .A(b[3]), .B(n280), .ZN(n348) );
  OAI22_X1 U355 ( .A1(n349), .A2(n301), .B1(n300), .B2(n299), .ZN(n100) );
  XNOR2_X1 U356 ( .A(b[5]), .B(n280), .ZN(n300) );
  NAND2_X1 U357 ( .A1(a[1]), .A2(n299), .ZN(n301) );
  XNOR2_X1 U358 ( .A(b[4]), .B(n280), .ZN(n349) );
endmodule


module datapath_DW01_add_3 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n84;
  wire   [15:1] carry;

  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n84), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[14]), .ZN(n53) );
  CLKBUF_X1 U2 ( .A(B[13]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(n34), .Z(n2) );
  NAND3_X1 U4 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n3) );
  NAND3_X1 U5 ( .A1(n71), .A2(n72), .A3(n73), .ZN(n4) );
  CLKBUF_X1 U6 ( .A(n78), .Z(n5) );
  NAND3_X1 U7 ( .A1(n9), .A2(n10), .A3(n11), .ZN(n6) );
  NAND3_X1 U8 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n7) );
  XOR2_X1 U9 ( .A(carry[2]), .B(A[2]), .Z(n8) );
  XOR2_X1 U10 ( .A(B[2]), .B(n8), .Z(SUM[2]) );
  NAND2_X1 U11 ( .A1(B[2]), .A2(carry[2]), .ZN(n9) );
  NAND2_X1 U12 ( .A1(B[2]), .A2(A[2]), .ZN(n10) );
  NAND2_X1 U13 ( .A1(carry[2]), .A2(A[2]), .ZN(n11) );
  NAND3_X1 U14 ( .A1(n9), .A2(n10), .A3(n11), .ZN(carry[3]) );
  CLKBUF_X1 U15 ( .A(carry[8]), .Z(n12) );
  NAND3_X1 U16 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n13) );
  NAND3_X1 U17 ( .A1(n33), .A2(n2), .A3(n35), .ZN(n14) );
  NAND3_X1 U18 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n15) );
  XOR2_X1 U19 ( .A(B[7]), .B(A[7]), .Z(n16) );
  XOR2_X1 U20 ( .A(n14), .B(n16), .Z(SUM[7]) );
  NAND2_X1 U21 ( .A1(n13), .A2(B[7]), .ZN(n17) );
  NAND2_X1 U22 ( .A1(carry[7]), .A2(A[7]), .ZN(n18) );
  NAND2_X1 U23 ( .A1(B[7]), .A2(A[7]), .ZN(n19) );
  NAND3_X1 U24 ( .A1(n17), .A2(n18), .A3(n19), .ZN(carry[8]) );
  NAND3_X1 U25 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n20) );
  NAND3_X1 U26 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n21) );
  CLKBUF_X1 U27 ( .A(n71), .Z(n22) );
  CLKBUF_X1 U28 ( .A(n42), .Z(n23) );
  NAND3_X1 U29 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n24) );
  NAND3_X1 U30 ( .A1(n41), .A2(n23), .A3(n43), .ZN(n25) );
  NAND3_X1 U31 ( .A1(n22), .A2(n72), .A3(n73), .ZN(n26) );
  XOR2_X1 U32 ( .A(n26), .B(A[11]), .Z(n27) );
  XOR2_X1 U33 ( .A(B[11]), .B(n27), .Z(SUM[11]) );
  NAND2_X1 U34 ( .A1(B[11]), .A2(n4), .ZN(n28) );
  NAND2_X1 U35 ( .A1(B[11]), .A2(A[11]), .ZN(n29) );
  NAND2_X1 U36 ( .A1(carry[11]), .A2(A[11]), .ZN(n30) );
  NAND3_X1 U37 ( .A1(n28), .A2(n29), .A3(n30), .ZN(carry[12]) );
  NAND3_X1 U38 ( .A1(n67), .A2(n68), .A3(n69), .ZN(n31) );
  XOR2_X1 U39 ( .A(B[6]), .B(A[6]), .Z(n32) );
  XOR2_X1 U40 ( .A(n21), .B(n32), .Z(SUM[6]) );
  NAND2_X1 U41 ( .A1(n20), .A2(B[6]), .ZN(n33) );
  NAND2_X1 U42 ( .A1(carry[6]), .A2(A[6]), .ZN(n34) );
  NAND2_X1 U43 ( .A1(B[6]), .A2(A[6]), .ZN(n35) );
  NAND3_X1 U44 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[7]) );
  XOR2_X1 U45 ( .A(B[3]), .B(A[3]), .Z(n36) );
  XOR2_X1 U46 ( .A(n6), .B(n36), .Z(SUM[3]) );
  NAND2_X1 U47 ( .A1(n6), .A2(B[3]), .ZN(n37) );
  NAND2_X1 U48 ( .A1(carry[3]), .A2(A[3]), .ZN(n38) );
  NAND2_X1 U49 ( .A1(B[3]), .A2(A[3]), .ZN(n39) );
  NAND3_X1 U50 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[4]) );
  XOR2_X1 U51 ( .A(B[8]), .B(A[8]), .Z(n40) );
  XOR2_X1 U52 ( .A(n12), .B(n40), .Z(SUM[8]) );
  NAND2_X1 U53 ( .A1(n7), .A2(B[8]), .ZN(n41) );
  NAND2_X1 U54 ( .A1(carry[8]), .A2(A[8]), .ZN(n42) );
  NAND2_X1 U55 ( .A1(B[8]), .A2(A[8]), .ZN(n43) );
  NAND3_X1 U56 ( .A1(n42), .A2(n41), .A3(n43), .ZN(carry[9]) );
  CLKBUF_X1 U57 ( .A(n15), .Z(n44) );
  NAND3_X1 U58 ( .A1(n81), .A2(n82), .A3(n80), .ZN(n45) );
  CLKBUF_X1 U59 ( .A(n31), .Z(n46) );
  NAND3_X1 U60 ( .A1(n78), .A2(n77), .A3(n76), .ZN(n47) );
  NAND3_X1 U61 ( .A1(n76), .A2(n77), .A3(n5), .ZN(n48) );
  CLKBUF_X1 U62 ( .A(n61), .Z(n49) );
  CLKBUF_X1 U63 ( .A(n24), .Z(n50) );
  CLKBUF_X1 U64 ( .A(B[5]), .Z(n51) );
  NAND3_X1 U65 ( .A1(n59), .A2(n60), .A3(n49), .ZN(n52) );
  XNOR2_X1 U66 ( .A(B[14]), .B(n53), .ZN(n54) );
  XOR2_X1 U67 ( .A(n54), .B(n45), .Z(SUM[14]) );
  NAND2_X1 U68 ( .A1(n45), .A2(B[14]), .ZN(n55) );
  NAND2_X1 U69 ( .A1(carry[14]), .A2(A[14]), .ZN(n56) );
  NAND2_X1 U70 ( .A1(B[14]), .A2(A[14]), .ZN(n57) );
  NAND3_X1 U71 ( .A1(n55), .A2(n56), .A3(n57), .ZN(carry[15]) );
  XOR2_X1 U72 ( .A(A[4]), .B(B[4]), .Z(n58) );
  XOR2_X1 U73 ( .A(n58), .B(n50), .Z(SUM[4]) );
  NAND2_X1 U74 ( .A1(A[4]), .A2(B[4]), .ZN(n59) );
  NAND2_X1 U75 ( .A1(A[4]), .A2(carry[4]), .ZN(n60) );
  NAND2_X1 U76 ( .A1(B[4]), .A2(n24), .ZN(n61) );
  NAND3_X1 U77 ( .A1(n61), .A2(n60), .A3(n59), .ZN(carry[5]) );
  XOR2_X1 U78 ( .A(A[5]), .B(n51), .Z(n62) );
  XOR2_X1 U79 ( .A(n62), .B(n52), .Z(SUM[5]) );
  NAND2_X1 U80 ( .A1(A[5]), .A2(B[5]), .ZN(n63) );
  NAND2_X1 U81 ( .A1(A[5]), .A2(carry[5]), .ZN(n64) );
  NAND2_X1 U82 ( .A1(B[5]), .A2(carry[5]), .ZN(n65) );
  NAND3_X1 U83 ( .A1(n63), .A2(n64), .A3(n65), .ZN(carry[6]) );
  XOR2_X1 U84 ( .A(B[9]), .B(A[9]), .Z(n66) );
  XOR2_X1 U85 ( .A(n25), .B(n66), .Z(SUM[9]) );
  NAND2_X1 U86 ( .A1(n3), .A2(B[9]), .ZN(n67) );
  NAND2_X1 U87 ( .A1(carry[9]), .A2(A[9]), .ZN(n68) );
  NAND2_X1 U88 ( .A1(B[9]), .A2(A[9]), .ZN(n69) );
  NAND3_X1 U89 ( .A1(n67), .A2(n68), .A3(n69), .ZN(carry[10]) );
  XOR2_X1 U90 ( .A(B[10]), .B(A[10]), .Z(n70) );
  XOR2_X1 U91 ( .A(n46), .B(n70), .Z(SUM[10]) );
  NAND2_X1 U92 ( .A1(n31), .A2(B[10]), .ZN(n71) );
  NAND2_X1 U93 ( .A1(carry[10]), .A2(A[10]), .ZN(n72) );
  NAND2_X1 U94 ( .A1(B[10]), .A2(A[10]), .ZN(n73) );
  NAND3_X1 U95 ( .A1(n71), .A2(n72), .A3(n73), .ZN(carry[11]) );
  NAND2_X1 U96 ( .A1(A[12]), .A2(B[12]), .ZN(n76) );
  XNOR2_X1 U97 ( .A(carry[15]), .B(n74), .ZN(SUM[15]) );
  XNOR2_X1 U98 ( .A(B[15]), .B(A[15]), .ZN(n74) );
  XOR2_X1 U99 ( .A(A[12]), .B(B[12]), .Z(n75) );
  XOR2_X1 U100 ( .A(n75), .B(n44), .Z(SUM[12]) );
  NAND2_X1 U101 ( .A1(A[12]), .A2(carry[12]), .ZN(n77) );
  NAND2_X1 U102 ( .A1(B[12]), .A2(n15), .ZN(n78) );
  NAND3_X1 U103 ( .A1(n78), .A2(n77), .A3(n76), .ZN(carry[13]) );
  XOR2_X1 U104 ( .A(A[13]), .B(n1), .Z(n79) );
  XOR2_X1 U105 ( .A(n79), .B(n48), .Z(SUM[13]) );
  NAND2_X1 U106 ( .A1(B[13]), .A2(A[13]), .ZN(n80) );
  NAND2_X1 U107 ( .A1(A[13]), .A2(carry[13]), .ZN(n81) );
  NAND2_X1 U108 ( .A1(B[13]), .A2(n47), .ZN(n82) );
  NAND3_X1 U109 ( .A1(n82), .A2(n81), .A3(n80), .ZN(carry[14]) );
  XOR2_X1 U110 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U111 ( .A1(B[0]), .A2(A[0]), .ZN(n84) );
endmodule


module datapath_DW_mult_tc_2 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343;

  FA_X1 U11 ( .A(n50), .B(n53), .CI(n11), .CO(n10), .S(product[5]) );
  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n286), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n285), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n289), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n288), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n291), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n208), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n215), .B(n102), .CO(n55), .S(n56) );
  NAND2_X1 U157 ( .A1(n309), .A2(n338), .ZN(n311) );
  AND3_X1 U158 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n224) );
  CLKBUF_X1 U159 ( .A(n243), .Z(n206) );
  NAND2_X1 U160 ( .A1(n231), .A2(n33), .ZN(n207) );
  AND2_X1 U161 ( .A1(n70), .A2(n87), .ZN(n208) );
  XOR2_X1 U162 ( .A(n283), .B(n15), .Z(n209) );
  AND3_X1 U163 ( .A1(n276), .A2(n277), .A3(n278), .ZN(product[15]) );
  XOR2_X1 U164 ( .A(n17), .B(n282), .Z(n211) );
  NAND3_X1 U165 ( .A1(n234), .A2(n235), .A3(n236), .ZN(n212) );
  NAND2_X2 U166 ( .A1(n320), .A2(n339), .ZN(n322) );
  NAND3_X1 U167 ( .A1(n262), .A2(n261), .A3(n260), .ZN(n213) );
  CLKBUF_X1 U168 ( .A(n252), .Z(n214) );
  BUF_X1 U169 ( .A(n309), .Z(n252) );
  OAI22_X1 U170 ( .A1(n300), .A2(n301), .B1(n280), .B2(n302), .ZN(n215) );
  XNOR2_X1 U171 ( .A(n211), .B(n216), .ZN(product[13]) );
  AND3_X1 U172 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n216) );
  NAND2_X1 U173 ( .A1(n218), .A2(n27), .ZN(n217) );
  NAND3_X1 U174 ( .A1(n207), .A2(n240), .A3(n241), .ZN(n218) );
  XOR2_X1 U175 ( .A(n70), .B(n87), .Z(n52) );
  CLKBUF_X1 U176 ( .A(n311), .Z(n219) );
  CLKBUF_X1 U177 ( .A(n13), .Z(n220) );
  AND3_X1 U178 ( .A1(n217), .A2(n250), .A3(n251), .ZN(n222) );
  NAND3_X1 U179 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n221) );
  XNOR2_X1 U180 ( .A(n222), .B(n223), .ZN(product[11]) );
  XOR2_X1 U181 ( .A(n23), .B(n20), .Z(n223) );
  XNOR2_X1 U182 ( .A(n209), .B(n224), .ZN(product[14]) );
  XOR2_X1 U183 ( .A(n95), .B(n102), .Z(n225) );
  XNOR2_X1 U184 ( .A(n226), .B(n220), .ZN(product[3]) );
  XNOR2_X1 U185 ( .A(n56), .B(n71), .ZN(n226) );
  NAND3_X1 U186 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n227) );
  NAND3_X1 U187 ( .A1(n242), .A2(n206), .A3(n244), .ZN(n228) );
  NAND3_X1 U188 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n229) );
  NAND3_X1 U189 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n230) );
  NAND3_X1 U190 ( .A1(n235), .A2(n234), .A3(n236), .ZN(n231) );
  NAND3_X1 U191 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n232) );
  XOR2_X1 U192 ( .A(n34), .B(n39), .Z(n233) );
  XOR2_X1 U193 ( .A(n230), .B(n233), .Z(product[8]) );
  NAND2_X1 U194 ( .A1(n229), .A2(n34), .ZN(n234) );
  NAND2_X1 U195 ( .A1(n8), .A2(n39), .ZN(n235) );
  NAND2_X1 U196 ( .A1(n34), .A2(n39), .ZN(n236) );
  NAND3_X1 U197 ( .A1(n234), .A2(n235), .A3(n236), .ZN(n7) );
  NAND3_X1 U198 ( .A1(n207), .A2(n240), .A3(n241), .ZN(n237) );
  XOR2_X1 U199 ( .A(n33), .B(n28), .Z(n238) );
  XOR2_X1 U200 ( .A(n212), .B(n238), .Z(product[9]) );
  NAND2_X1 U201 ( .A1(n231), .A2(n33), .ZN(n239) );
  NAND2_X1 U202 ( .A1(n7), .A2(n28), .ZN(n240) );
  NAND2_X1 U203 ( .A1(n33), .A2(n28), .ZN(n241) );
  NAND3_X1 U204 ( .A1(n240), .A2(n241), .A3(n239), .ZN(n6) );
  NAND2_X1 U205 ( .A1(n13), .A2(n225), .ZN(n242) );
  NAND2_X1 U206 ( .A1(n13), .A2(n71), .ZN(n243) );
  NAND2_X1 U207 ( .A1(n225), .A2(n71), .ZN(n244) );
  NAND3_X1 U208 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n12) );
  NAND3_X1 U209 ( .A1(n217), .A2(n250), .A3(n251), .ZN(n245) );
  CLKBUF_X1 U210 ( .A(b[0]), .Z(n246) );
  XNOR2_X1 U211 ( .A(n228), .B(n247), .ZN(product[4]) );
  XNOR2_X1 U212 ( .A(n54), .B(n55), .ZN(n247) );
  XOR2_X1 U213 ( .A(n27), .B(n24), .Z(n248) );
  XOR2_X1 U214 ( .A(n237), .B(n248), .Z(product[10]) );
  NAND2_X1 U215 ( .A1(n218), .A2(n27), .ZN(n249) );
  NAND2_X1 U216 ( .A1(n6), .A2(n24), .ZN(n250) );
  NAND2_X1 U217 ( .A1(n27), .A2(n24), .ZN(n251) );
  NAND3_X1 U218 ( .A1(n250), .A2(n249), .A3(n251), .ZN(n5) );
  XNOR2_X1 U219 ( .A(a[4]), .B(a[3]), .ZN(n309) );
  XOR2_X1 U220 ( .A(n18), .B(n19), .Z(n253) );
  XOR2_X1 U221 ( .A(n4), .B(n253), .Z(product[12]) );
  NAND2_X1 U222 ( .A1(n4), .A2(n18), .ZN(n254) );
  NAND2_X1 U223 ( .A1(n4), .A2(n19), .ZN(n255) );
  NAND2_X1 U224 ( .A1(n18), .A2(n19), .ZN(n256) );
  NAND3_X1 U225 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n3) );
  NAND3_X1 U226 ( .A1(n261), .A2(n260), .A3(n262), .ZN(n257) );
  CLKBUF_X1 U227 ( .A(n301), .Z(n258) );
  XOR2_X1 U228 ( .A(n46), .B(n49), .Z(n259) );
  XOR2_X1 U229 ( .A(n10), .B(n259), .Z(product[6]) );
  NAND2_X1 U230 ( .A1(n46), .A2(n49), .ZN(n260) );
  NAND2_X1 U231 ( .A1(n10), .A2(n46), .ZN(n261) );
  NAND2_X1 U232 ( .A1(n10), .A2(n49), .ZN(n262) );
  NAND3_X1 U233 ( .A1(n262), .A2(n261), .A3(n260), .ZN(n9) );
  XOR2_X1 U234 ( .A(n40), .B(n45), .Z(n263) );
  XOR2_X1 U235 ( .A(n263), .B(n257), .Z(product[7]) );
  NAND2_X1 U236 ( .A1(n40), .A2(n45), .ZN(n264) );
  NAND2_X1 U237 ( .A1(n213), .A2(n40), .ZN(n265) );
  NAND2_X1 U238 ( .A1(n9), .A2(n45), .ZN(n266) );
  NAND3_X1 U239 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n8) );
  NAND2_X1 U240 ( .A1(n227), .A2(n54), .ZN(n267) );
  NAND2_X1 U241 ( .A1(n12), .A2(n55), .ZN(n268) );
  NAND2_X1 U242 ( .A1(n54), .A2(n55), .ZN(n269) );
  NAND3_X1 U243 ( .A1(n267), .A2(n268), .A3(n269), .ZN(n11) );
  NAND2_X1 U244 ( .A1(n5), .A2(n23), .ZN(n270) );
  NAND2_X1 U245 ( .A1(n245), .A2(n20), .ZN(n271) );
  NAND2_X1 U246 ( .A1(n23), .A2(n20), .ZN(n272) );
  NAND3_X1 U247 ( .A1(n271), .A2(n270), .A3(n272), .ZN(n4) );
  NAND2_X1 U248 ( .A1(n17), .A2(n282), .ZN(n273) );
  NAND2_X1 U249 ( .A1(n17), .A2(n221), .ZN(n274) );
  NAND2_X1 U250 ( .A1(n3), .A2(n282), .ZN(n275) );
  NAND2_X1 U251 ( .A1(n283), .A2(n15), .ZN(n276) );
  NAND2_X1 U252 ( .A1(n283), .A2(n232), .ZN(n277) );
  NAND2_X1 U253 ( .A1(n15), .A2(n232), .ZN(n278) );
  INV_X1 U254 ( .A(n281), .ZN(n279) );
  INV_X1 U255 ( .A(n15), .ZN(n282) );
  INV_X1 U256 ( .A(n31), .ZN(n288) );
  INV_X1 U257 ( .A(n21), .ZN(n285) );
  INV_X1 U258 ( .A(n318), .ZN(n286) );
  INV_X1 U259 ( .A(n329), .ZN(n283) );
  INV_X1 U260 ( .A(n298), .ZN(n291) );
  INV_X1 U261 ( .A(n307), .ZN(n289) );
  INV_X1 U262 ( .A(a[5]), .ZN(n287) );
  INV_X1 U263 ( .A(a[7]), .ZN(n284) );
  INV_X1 U264 ( .A(b[0]), .ZN(n281) );
  BUF_X2 U265 ( .A(n299), .Z(n280) );
  XNOR2_X1 U266 ( .A(a[2]), .B(a[1]), .ZN(n299) );
  INV_X1 U267 ( .A(a[3]), .ZN(n290) );
  INV_X1 U268 ( .A(a[1]), .ZN(n292) );
  NAND2_X2 U269 ( .A1(n299), .A2(n337), .ZN(n301) );
  XOR2_X2 U270 ( .A(a[6]), .B(n287), .Z(n320) );
  INV_X2 U271 ( .A(a[0]), .ZN(n293) );
  NOR2_X1 U272 ( .A1(n293), .A2(n281), .ZN(product[0]) );
  OAI22_X1 U273 ( .A1(n294), .A2(n295), .B1(n296), .B2(n293), .ZN(n99) );
  OAI22_X1 U274 ( .A1(n296), .A2(n295), .B1(n297), .B2(n293), .ZN(n98) );
  XNOR2_X1 U275 ( .A(b[6]), .B(a[1]), .ZN(n296) );
  OAI22_X1 U276 ( .A1(n293), .A2(n297), .B1(n295), .B2(n297), .ZN(n298) );
  XNOR2_X1 U277 ( .A(b[7]), .B(a[1]), .ZN(n297) );
  NOR2_X1 U278 ( .A1(n280), .A2(n281), .ZN(n96) );
  OAI22_X1 U279 ( .A1(n300), .A2(n301), .B1(n280), .B2(n302), .ZN(n95) );
  XNOR2_X1 U280 ( .A(a[3]), .B(n246), .ZN(n300) );
  OAI22_X1 U281 ( .A1(n302), .A2(n301), .B1(n280), .B2(n303), .ZN(n94) );
  XNOR2_X1 U282 ( .A(b[1]), .B(a[3]), .ZN(n302) );
  OAI22_X1 U283 ( .A1(n303), .A2(n301), .B1(n280), .B2(n304), .ZN(n93) );
  XNOR2_X1 U284 ( .A(b[2]), .B(a[3]), .ZN(n303) );
  OAI22_X1 U285 ( .A1(n304), .A2(n301), .B1(n280), .B2(n305), .ZN(n92) );
  XNOR2_X1 U286 ( .A(b[3]), .B(a[3]), .ZN(n304) );
  OAI22_X1 U287 ( .A1(n305), .A2(n301), .B1(n280), .B2(n306), .ZN(n91) );
  XNOR2_X1 U288 ( .A(b[4]), .B(a[3]), .ZN(n305) );
  OAI22_X1 U289 ( .A1(n308), .A2(n280), .B1(n258), .B2(n308), .ZN(n307) );
  NOR2_X1 U290 ( .A1(n252), .A2(n281), .ZN(n88) );
  OAI22_X1 U291 ( .A1(n310), .A2(n311), .B1(n252), .B2(n312), .ZN(n87) );
  XNOR2_X1 U292 ( .A(a[5]), .B(n279), .ZN(n310) );
  OAI22_X1 U293 ( .A1(n312), .A2(n311), .B1(n214), .B2(n313), .ZN(n86) );
  XNOR2_X1 U294 ( .A(b[1]), .B(a[5]), .ZN(n312) );
  OAI22_X1 U295 ( .A1(n313), .A2(n311), .B1(n252), .B2(n314), .ZN(n85) );
  XNOR2_X1 U296 ( .A(b[2]), .B(a[5]), .ZN(n313) );
  OAI22_X1 U297 ( .A1(n314), .A2(n311), .B1(n214), .B2(n315), .ZN(n84) );
  XNOR2_X1 U298 ( .A(b[3]), .B(a[5]), .ZN(n314) );
  OAI22_X1 U299 ( .A1(n315), .A2(n219), .B1(n214), .B2(n316), .ZN(n83) );
  XNOR2_X1 U300 ( .A(b[4]), .B(a[5]), .ZN(n315) );
  OAI22_X1 U301 ( .A1(n316), .A2(n219), .B1(n214), .B2(n317), .ZN(n82) );
  XNOR2_X1 U302 ( .A(b[5]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U303 ( .A1(n319), .A2(n214), .B1(n219), .B2(n319), .ZN(n318) );
  NOR2_X1 U304 ( .A1(n320), .A2(n281), .ZN(n80) );
  OAI22_X1 U305 ( .A1(n321), .A2(n322), .B1(n320), .B2(n323), .ZN(n79) );
  XNOR2_X1 U306 ( .A(a[7]), .B(n279), .ZN(n321) );
  OAI22_X1 U307 ( .A1(n324), .A2(n322), .B1(n320), .B2(n325), .ZN(n77) );
  OAI22_X1 U308 ( .A1(n325), .A2(n322), .B1(n320), .B2(n326), .ZN(n76) );
  XNOR2_X1 U309 ( .A(b[3]), .B(a[7]), .ZN(n325) );
  OAI22_X1 U310 ( .A1(n326), .A2(n322), .B1(n320), .B2(n327), .ZN(n75) );
  XNOR2_X1 U311 ( .A(b[4]), .B(a[7]), .ZN(n326) );
  OAI22_X1 U312 ( .A1(n327), .A2(n322), .B1(n320), .B2(n328), .ZN(n74) );
  XNOR2_X1 U313 ( .A(b[5]), .B(a[7]), .ZN(n327) );
  OAI22_X1 U314 ( .A1(n330), .A2(n320), .B1(n322), .B2(n330), .ZN(n329) );
  OAI21_X1 U315 ( .B1(n246), .B2(n292), .A(n295), .ZN(n72) );
  OAI21_X1 U316 ( .B1(n290), .B2(n301), .A(n331), .ZN(n71) );
  OR3_X1 U317 ( .A1(n280), .A2(n279), .A3(n290), .ZN(n331) );
  OAI21_X1 U318 ( .B1(n287), .B2(n311), .A(n332), .ZN(n70) );
  OR3_X1 U319 ( .A1(n252), .A2(n279), .A3(n287), .ZN(n332) );
  OAI21_X1 U320 ( .B1(n284), .B2(n322), .A(n333), .ZN(n69) );
  OR3_X1 U321 ( .A1(n320), .A2(n279), .A3(n284), .ZN(n333) );
  XNOR2_X1 U322 ( .A(n334), .B(n335), .ZN(n38) );
  OR2_X1 U323 ( .A1(n334), .A2(n335), .ZN(n37) );
  OAI22_X1 U324 ( .A1(n306), .A2(n258), .B1(n280), .B2(n336), .ZN(n335) );
  XNOR2_X1 U325 ( .A(b[5]), .B(a[3]), .ZN(n306) );
  OAI22_X1 U326 ( .A1(n323), .A2(n322), .B1(n320), .B2(n324), .ZN(n334) );
  XNOR2_X1 U327 ( .A(b[2]), .B(a[7]), .ZN(n324) );
  XNOR2_X1 U328 ( .A(b[1]), .B(a[7]), .ZN(n323) );
  OAI22_X1 U329 ( .A1(n336), .A2(n258), .B1(n280), .B2(n308), .ZN(n31) );
  XNOR2_X1 U330 ( .A(b[7]), .B(a[3]), .ZN(n308) );
  XNOR2_X1 U331 ( .A(n290), .B(a[2]), .ZN(n337) );
  XNOR2_X1 U332 ( .A(b[6]), .B(a[3]), .ZN(n336) );
  OAI22_X1 U333 ( .A1(n317), .A2(n219), .B1(n214), .B2(n319), .ZN(n21) );
  XNOR2_X1 U334 ( .A(b[7]), .B(a[5]), .ZN(n319) );
  XNOR2_X1 U335 ( .A(n287), .B(a[4]), .ZN(n338) );
  XNOR2_X1 U336 ( .A(b[6]), .B(a[5]), .ZN(n317) );
  OAI22_X1 U337 ( .A1(n328), .A2(n322), .B1(n320), .B2(n330), .ZN(n15) );
  XNOR2_X1 U338 ( .A(b[7]), .B(a[7]), .ZN(n330) );
  XNOR2_X1 U339 ( .A(n284), .B(a[6]), .ZN(n339) );
  XNOR2_X1 U340 ( .A(b[6]), .B(a[7]), .ZN(n328) );
  OAI22_X1 U341 ( .A1(n246), .A2(n295), .B1(n340), .B2(n293), .ZN(n104) );
  OAI22_X1 U342 ( .A1(n340), .A2(n295), .B1(n341), .B2(n293), .ZN(n103) );
  XNOR2_X1 U343 ( .A(b[1]), .B(a[1]), .ZN(n340) );
  OAI22_X1 U344 ( .A1(n295), .A2(n341), .B1(n342), .B2(n293), .ZN(n102) );
  XNOR2_X1 U345 ( .A(b[2]), .B(a[1]), .ZN(n341) );
  OAI22_X1 U346 ( .A1(n342), .A2(n295), .B1(n343), .B2(n293), .ZN(n101) );
  XNOR2_X1 U347 ( .A(b[3]), .B(a[1]), .ZN(n342) );
  OAI22_X1 U348 ( .A1(n343), .A2(n295), .B1(n294), .B2(n293), .ZN(n100) );
  XNOR2_X1 U349 ( .A(b[5]), .B(a[1]), .ZN(n294) );
  NAND2_X1 U350 ( .A1(a[1]), .A2(n293), .ZN(n295) );
  XNOR2_X1 U351 ( .A(b[4]), .B(a[1]), .ZN(n343) );
endmodule


module datapath_DW01_add_2 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n72;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n72), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(B[2]), .Z(n1) );
  NAND3_X1 U2 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n2) );
  CLKBUF_X1 U3 ( .A(n7), .Z(n3) );
  NAND3_X1 U4 ( .A1(n23), .A2(n24), .A3(n25), .ZN(n4) );
  CLKBUF_X1 U5 ( .A(B[6]), .Z(n5) );
  NAND3_X1 U6 ( .A1(n60), .A2(n59), .A3(n61), .ZN(n6) );
  NAND3_X1 U7 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n7) );
  NAND3_X1 U8 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n8) );
  XOR2_X1 U9 ( .A(carry[2]), .B(A[2]), .Z(n9) );
  XOR2_X1 U10 ( .A(n1), .B(n9), .Z(SUM[2]) );
  NAND2_X1 U11 ( .A1(B[2]), .A2(carry[2]), .ZN(n10) );
  NAND2_X1 U12 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  NAND2_X1 U13 ( .A1(carry[2]), .A2(A[2]), .ZN(n12) );
  NAND3_X1 U14 ( .A1(n10), .A2(n11), .A3(n12), .ZN(carry[3]) );
  NAND3_X1 U15 ( .A1(n17), .A2(n19), .A3(n18), .ZN(n13) );
  CLKBUF_X1 U16 ( .A(n6), .Z(n14) );
  CLKBUF_X1 U17 ( .A(n4), .Z(n15) );
  XOR2_X1 U18 ( .A(B[11]), .B(A[11]), .Z(n16) );
  XOR2_X1 U19 ( .A(n14), .B(n16), .Z(SUM[11]) );
  NAND2_X1 U20 ( .A1(n6), .A2(B[11]), .ZN(n17) );
  NAND2_X1 U21 ( .A1(carry[11]), .A2(A[11]), .ZN(n18) );
  NAND2_X1 U22 ( .A1(B[11]), .A2(A[11]), .ZN(n19) );
  NAND3_X1 U23 ( .A1(n17), .A2(n19), .A3(n18), .ZN(carry[12]) );
  NAND3_X1 U24 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n20) );
  CLKBUF_X1 U25 ( .A(n53), .Z(n21) );
  XOR2_X1 U26 ( .A(B[4]), .B(A[4]), .Z(n22) );
  XOR2_X1 U27 ( .A(carry[4]), .B(n22), .Z(SUM[4]) );
  NAND2_X1 U28 ( .A1(n8), .A2(B[4]), .ZN(n23) );
  NAND2_X1 U29 ( .A1(carry[4]), .A2(A[4]), .ZN(n24) );
  NAND2_X1 U30 ( .A1(B[4]), .A2(A[4]), .ZN(n25) );
  NAND3_X1 U31 ( .A1(n23), .A2(n24), .A3(n25), .ZN(carry[5]) );
  NAND3_X1 U32 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n26) );
  NAND3_X1 U33 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n27) );
  XOR2_X1 U34 ( .A(B[5]), .B(A[5]), .Z(n28) );
  XOR2_X1 U35 ( .A(n15), .B(n28), .Z(SUM[5]) );
  NAND2_X1 U36 ( .A1(n4), .A2(B[5]), .ZN(n29) );
  NAND2_X1 U37 ( .A1(carry[5]), .A2(A[5]), .ZN(n30) );
  NAND2_X1 U38 ( .A1(B[5]), .A2(A[5]), .ZN(n31) );
  NAND3_X1 U39 ( .A1(n29), .A2(n30), .A3(n31), .ZN(carry[6]) );
  CLKBUF_X1 U40 ( .A(carry[3]), .Z(n32) );
  XOR2_X1 U41 ( .A(B[3]), .B(A[3]), .Z(n33) );
  XOR2_X1 U42 ( .A(n32), .B(n33), .Z(SUM[3]) );
  NAND2_X1 U43 ( .A1(B[3]), .A2(carry[3]), .ZN(n34) );
  NAND2_X1 U44 ( .A1(carry[3]), .A2(A[3]), .ZN(n35) );
  NAND2_X1 U45 ( .A1(B[3]), .A2(A[3]), .ZN(n36) );
  NAND3_X1 U46 ( .A1(n34), .A2(n35), .A3(n36), .ZN(carry[4]) );
  NAND3_X1 U47 ( .A1(n50), .A2(n51), .A3(n52), .ZN(n37) );
  XOR2_X1 U48 ( .A(B[7]), .B(A[7]), .Z(n38) );
  XOR2_X1 U49 ( .A(carry[7]), .B(n38), .Z(SUM[7]) );
  NAND2_X1 U50 ( .A1(n2), .A2(B[7]), .ZN(n39) );
  NAND2_X1 U51 ( .A1(n20), .A2(A[7]), .ZN(n40) );
  NAND2_X1 U52 ( .A1(B[7]), .A2(A[7]), .ZN(n41) );
  NAND3_X1 U53 ( .A1(n39), .A2(n40), .A3(n41), .ZN(carry[8]) );
  XOR2_X1 U54 ( .A(n5), .B(A[6]), .Z(n42) );
  XOR2_X1 U55 ( .A(n26), .B(n42), .Z(SUM[6]) );
  NAND2_X1 U56 ( .A1(n26), .A2(B[6]), .ZN(n43) );
  NAND2_X1 U57 ( .A1(carry[6]), .A2(A[6]), .ZN(n44) );
  NAND2_X1 U58 ( .A1(B[6]), .A2(A[6]), .ZN(n45) );
  NAND3_X1 U59 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[7]) );
  CLKBUF_X1 U60 ( .A(n13), .Z(n46) );
  CLKBUF_X1 U61 ( .A(carry[10]), .Z(n47) );
  CLKBUF_X1 U62 ( .A(n27), .Z(n48) );
  XOR2_X1 U63 ( .A(B[9]), .B(A[9]), .Z(n49) );
  XOR2_X1 U64 ( .A(n48), .B(n49), .Z(SUM[9]) );
  NAND2_X1 U65 ( .A1(n27), .A2(B[9]), .ZN(n50) );
  NAND2_X1 U66 ( .A1(carry[9]), .A2(A[9]), .ZN(n51) );
  NAND2_X1 U67 ( .A1(B[9]), .A2(A[9]), .ZN(n52) );
  NAND3_X1 U68 ( .A1(n50), .A2(n51), .A3(n52), .ZN(carry[10]) );
  NAND3_X1 U69 ( .A1(n66), .A2(n65), .A3(n64), .ZN(n53) );
  XOR2_X1 U70 ( .A(B[8]), .B(A[8]), .Z(n54) );
  XOR2_X1 U71 ( .A(n3), .B(n54), .Z(SUM[8]) );
  NAND2_X1 U72 ( .A1(n7), .A2(B[8]), .ZN(n55) );
  NAND2_X1 U73 ( .A1(carry[8]), .A2(A[8]), .ZN(n56) );
  NAND2_X1 U74 ( .A1(B[8]), .A2(A[8]), .ZN(n57) );
  NAND3_X1 U75 ( .A1(n55), .A2(n57), .A3(n56), .ZN(carry[9]) );
  XOR2_X1 U76 ( .A(B[10]), .B(A[10]), .Z(n58) );
  XOR2_X1 U77 ( .A(n47), .B(n58), .Z(SUM[10]) );
  NAND2_X1 U78 ( .A1(n37), .A2(B[10]), .ZN(n59) );
  NAND2_X1 U79 ( .A1(carry[10]), .A2(A[10]), .ZN(n60) );
  NAND2_X1 U80 ( .A1(B[10]), .A2(A[10]), .ZN(n61) );
  NAND3_X1 U81 ( .A1(n60), .A2(n59), .A3(n61), .ZN(carry[11]) );
  NAND2_X1 U82 ( .A1(B[12]), .A2(A[12]), .ZN(n64) );
  XNOR2_X1 U83 ( .A(carry[15]), .B(n62), .ZN(SUM[15]) );
  XNOR2_X1 U84 ( .A(B[15]), .B(A[15]), .ZN(n62) );
  XOR2_X1 U85 ( .A(A[12]), .B(B[12]), .Z(n63) );
  XOR2_X1 U86 ( .A(n63), .B(n46), .Z(SUM[12]) );
  NAND2_X1 U87 ( .A1(A[12]), .A2(carry[12]), .ZN(n65) );
  NAND2_X1 U88 ( .A1(B[12]), .A2(n13), .ZN(n66) );
  NAND3_X1 U89 ( .A1(n66), .A2(n65), .A3(n64), .ZN(carry[13]) );
  XOR2_X1 U90 ( .A(A[13]), .B(B[13]), .Z(n67) );
  XOR2_X1 U91 ( .A(n67), .B(n21), .Z(SUM[13]) );
  NAND2_X1 U92 ( .A1(B[13]), .A2(A[13]), .ZN(n68) );
  NAND2_X1 U93 ( .A1(n53), .A2(A[13]), .ZN(n69) );
  NAND2_X1 U94 ( .A1(carry[13]), .A2(B[13]), .ZN(n70) );
  NAND3_X1 U95 ( .A1(n69), .A2(n70), .A3(n68), .ZN(carry[14]) );
  XOR2_X1 U96 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U97 ( .A1(B[0]), .A2(A[0]), .ZN(n72) );
endmodule


module datapath_DW_mult_tc_1 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354;

  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n298), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n297), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n301), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n300), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n303), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  BUF_X2 U157 ( .A(a[1]), .Z(n283) );
  NAND3_X1 U158 ( .A1(n288), .A2(n289), .A3(n290), .ZN(n49) );
  INV_X1 U159 ( .A(n15), .ZN(n294) );
  NAND3_X1 U160 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n206) );
  CLKBUF_X1 U161 ( .A(b[1]), .Z(n207) );
  AND3_X1 U162 ( .A1(n267), .A2(n268), .A3(n269), .ZN(product[15]) );
  XNOR2_X1 U163 ( .A(n295), .B(n15), .ZN(n209) );
  NAND3_X1 U164 ( .A1(n230), .A2(n229), .A3(n231), .ZN(n210) );
  NAND3_X1 U165 ( .A1(n230), .A2(n229), .A3(n231), .ZN(n211) );
  NAND3_X1 U166 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n212) );
  NAND3_X1 U167 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n213) );
  NAND2_X1 U168 ( .A1(n310), .A2(n348), .ZN(n312) );
  NAND2_X2 U169 ( .A1(n331), .A2(n350), .ZN(n333) );
  NAND3_X1 U170 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n214) );
  XNOR2_X1 U171 ( .A(n236), .B(n215), .ZN(product[3]) );
  XNOR2_X1 U172 ( .A(n56), .B(n71), .ZN(n215) );
  NAND3_X1 U173 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n216) );
  NAND3_X1 U174 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n217) );
  OAI22_X1 U175 ( .A1(n311), .A2(n312), .B1(n285), .B2(n313), .ZN(n218) );
  XOR2_X1 U176 ( .A(n218), .B(n102), .Z(n219) );
  NAND3_X1 U177 ( .A1(n275), .A2(n276), .A3(n277), .ZN(n220) );
  NAND2_X2 U178 ( .A1(a[1]), .A2(n304), .ZN(n306) );
  BUF_X2 U179 ( .A(n285), .Z(n221) );
  NAND3_X1 U180 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n222) );
  XOR2_X1 U181 ( .A(n46), .B(n49), .Z(n223) );
  XOR2_X1 U182 ( .A(n217), .B(n223), .Z(product[6]) );
  NAND2_X1 U183 ( .A1(n216), .A2(n46), .ZN(n224) );
  NAND2_X1 U184 ( .A1(n10), .A2(n49), .ZN(n225) );
  NAND2_X1 U185 ( .A1(n46), .A2(n49), .ZN(n226) );
  NAND3_X1 U186 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n9) );
  NAND3_X1 U187 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n227) );
  XOR2_X1 U188 ( .A(n23), .B(n20), .Z(n228) );
  XOR2_X1 U189 ( .A(n5), .B(n228), .Z(product[11]) );
  NAND2_X1 U190 ( .A1(n5), .A2(n23), .ZN(n229) );
  NAND2_X1 U191 ( .A1(n5), .A2(n20), .ZN(n230) );
  NAND2_X1 U192 ( .A1(n23), .A2(n20), .ZN(n231) );
  NAND3_X1 U193 ( .A1(n229), .A2(n231), .A3(n230), .ZN(n4) );
  XOR2_X1 U194 ( .A(n40), .B(n45), .Z(n232) );
  XOR2_X1 U195 ( .A(n213), .B(n232), .Z(product[7]) );
  NAND2_X1 U196 ( .A1(n212), .A2(n40), .ZN(n233) );
  NAND2_X1 U197 ( .A1(n9), .A2(n45), .ZN(n234) );
  NAND2_X1 U198 ( .A1(n40), .A2(n45), .ZN(n235) );
  NAND3_X1 U199 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n8) );
  CLKBUF_X1 U200 ( .A(n13), .Z(n236) );
  NAND3_X1 U201 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n237) );
  XNOR2_X1 U202 ( .A(n220), .B(n209), .ZN(product[14]) );
  XOR2_X1 U203 ( .A(n34), .B(n39), .Z(n238) );
  XOR2_X1 U204 ( .A(n8), .B(n238), .Z(product[8]) );
  NAND2_X1 U205 ( .A1(n206), .A2(n34), .ZN(n239) );
  NAND2_X1 U206 ( .A1(n214), .A2(n39), .ZN(n240) );
  NAND2_X1 U207 ( .A1(n34), .A2(n39), .ZN(n241) );
  NAND3_X1 U208 ( .A1(n240), .A2(n239), .A3(n241), .ZN(n7) );
  NAND3_X1 U209 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n242) );
  NAND2_X1 U210 ( .A1(n13), .A2(n219), .ZN(n243) );
  NAND2_X1 U211 ( .A1(n13), .A2(n71), .ZN(n244) );
  NAND2_X1 U212 ( .A1(n219), .A2(n71), .ZN(n245) );
  NAND3_X1 U213 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n12) );
  NAND3_X1 U214 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n246) );
  NAND3_X1 U215 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n247) );
  NAND3_X1 U216 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n248) );
  XOR2_X1 U217 ( .A(n33), .B(n28), .Z(n249) );
  XOR2_X1 U218 ( .A(n237), .B(n249), .Z(product[9]) );
  NAND2_X1 U219 ( .A1(n237), .A2(n33), .ZN(n250) );
  NAND2_X1 U220 ( .A1(n7), .A2(n28), .ZN(n251) );
  NAND2_X1 U221 ( .A1(n33), .A2(n28), .ZN(n252) );
  XOR2_X1 U222 ( .A(n27), .B(n24), .Z(n253) );
  XOR2_X1 U223 ( .A(n222), .B(n253), .Z(product[10]) );
  NAND2_X1 U224 ( .A1(n247), .A2(n27), .ZN(n254) );
  NAND2_X1 U225 ( .A1(n222), .A2(n24), .ZN(n255) );
  NAND2_X1 U226 ( .A1(n27), .A2(n24), .ZN(n256) );
  NAND3_X1 U227 ( .A1(n255), .A2(n254), .A3(n256), .ZN(n5) );
  XNOR2_X1 U228 ( .A(b[3]), .B(n283), .ZN(n257) );
  CLKBUF_X1 U229 ( .A(n351), .Z(n258) );
  XOR2_X1 U230 ( .A(n54), .B(n55), .Z(n259) );
  XOR2_X1 U231 ( .A(n259), .B(n242), .Z(product[4]) );
  NAND2_X1 U232 ( .A1(n54), .A2(n55), .ZN(n260) );
  NAND2_X1 U233 ( .A1(n54), .A2(n242), .ZN(n261) );
  NAND2_X1 U234 ( .A1(n55), .A2(n12), .ZN(n262) );
  NAND3_X1 U235 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n11) );
  XOR2_X1 U236 ( .A(n50), .B(n53), .Z(n263) );
  XOR2_X1 U237 ( .A(n263), .B(n227), .Z(product[5]) );
  NAND2_X1 U238 ( .A1(n50), .A2(n53), .ZN(n264) );
  NAND2_X1 U239 ( .A1(n50), .A2(n248), .ZN(n265) );
  NAND2_X1 U240 ( .A1(n11), .A2(n53), .ZN(n266) );
  NAND3_X1 U241 ( .A1(n265), .A2(n264), .A3(n266), .ZN(n10) );
  NAND2_X1 U242 ( .A1(n2), .A2(n295), .ZN(n267) );
  NAND2_X1 U243 ( .A1(n2), .A2(n15), .ZN(n268) );
  NAND2_X1 U244 ( .A1(n295), .A2(n15), .ZN(n269) );
  XOR2_X1 U245 ( .A(n18), .B(n19), .Z(n270) );
  XOR2_X1 U246 ( .A(n211), .B(n270), .Z(product[12]) );
  NAND2_X1 U247 ( .A1(n210), .A2(n18), .ZN(n271) );
  NAND2_X1 U248 ( .A1(n4), .A2(n19), .ZN(n272) );
  NAND2_X1 U249 ( .A1(n18), .A2(n19), .ZN(n273) );
  NAND3_X1 U250 ( .A1(n272), .A2(n271), .A3(n273), .ZN(n3) );
  XOR2_X1 U251 ( .A(n17), .B(n294), .Z(n274) );
  XOR2_X1 U252 ( .A(n3), .B(n274), .Z(product[13]) );
  NAND2_X1 U253 ( .A1(n246), .A2(n17), .ZN(n275) );
  NAND2_X1 U254 ( .A1(n246), .A2(n294), .ZN(n276) );
  NAND2_X1 U255 ( .A1(n17), .A2(n294), .ZN(n277) );
  NAND3_X1 U256 ( .A1(n275), .A2(n276), .A3(n277), .ZN(n2) );
  CLKBUF_X1 U257 ( .A(b[3]), .Z(n278) );
  NAND2_X1 U258 ( .A1(a[4]), .A2(a[3]), .ZN(n281) );
  NAND2_X1 U259 ( .A1(n279), .A2(n280), .ZN(n282) );
  NAND2_X2 U260 ( .A1(n281), .A2(n282), .ZN(n320) );
  INV_X1 U261 ( .A(a[4]), .ZN(n279) );
  INV_X1 U262 ( .A(a[3]), .ZN(n280) );
  NAND2_X2 U263 ( .A1(n320), .A2(n349), .ZN(n322) );
  NAND2_X1 U264 ( .A1(n310), .A2(n348), .ZN(n284) );
  INV_X1 U265 ( .A(n31), .ZN(n300) );
  INV_X1 U266 ( .A(n21), .ZN(n297) );
  INV_X1 U267 ( .A(n329), .ZN(n298) );
  INV_X1 U268 ( .A(n340), .ZN(n295) );
  INV_X1 U269 ( .A(n309), .ZN(n303) );
  INV_X1 U270 ( .A(n318), .ZN(n301) );
  XOR2_X1 U271 ( .A(a[2]), .B(n291), .Z(n285) );
  XOR2_X1 U272 ( .A(a[2]), .B(n291), .Z(n310) );
  INV_X1 U273 ( .A(a[5]), .ZN(n299) );
  INV_X1 U274 ( .A(a[7]), .ZN(n296) );
  INV_X1 U275 ( .A(a[3]), .ZN(n302) );
  INV_X1 U276 ( .A(n293), .ZN(n286) );
  INV_X1 U277 ( .A(b[0]), .ZN(n293) );
  XNOR2_X1 U278 ( .A(n52), .B(n287), .ZN(n50) );
  XNOR2_X1 U279 ( .A(n93), .B(n100), .ZN(n287) );
  NAND2_X1 U280 ( .A1(n52), .A2(n93), .ZN(n288) );
  NAND2_X1 U281 ( .A1(n52), .A2(n100), .ZN(n289) );
  NAND2_X1 U282 ( .A1(n93), .A2(n100), .ZN(n290) );
  INV_X1 U283 ( .A(a[1]), .ZN(n291) );
  XOR2_X2 U284 ( .A(a[6]), .B(n299), .Z(n331) );
  INV_X1 U285 ( .A(n293), .ZN(n292) );
  INV_X2 U286 ( .A(a[0]), .ZN(n304) );
  NOR2_X1 U287 ( .A1(n304), .A2(n293), .ZN(product[0]) );
  OAI22_X1 U288 ( .A1(n305), .A2(n306), .B1(n307), .B2(n304), .ZN(n99) );
  OAI22_X1 U289 ( .A1(n307), .A2(n306), .B1(n308), .B2(n304), .ZN(n98) );
  XNOR2_X1 U290 ( .A(b[6]), .B(n283), .ZN(n307) );
  OAI22_X1 U291 ( .A1(n304), .A2(n308), .B1(n306), .B2(n308), .ZN(n309) );
  XNOR2_X1 U292 ( .A(b[7]), .B(n283), .ZN(n308) );
  NOR2_X1 U293 ( .A1(n285), .A2(n293), .ZN(n96) );
  OAI22_X1 U294 ( .A1(n311), .A2(n312), .B1(n285), .B2(n313), .ZN(n95) );
  XNOR2_X1 U295 ( .A(a[3]), .B(n292), .ZN(n311) );
  OAI22_X1 U296 ( .A1(n313), .A2(n284), .B1(n285), .B2(n314), .ZN(n94) );
  XNOR2_X1 U297 ( .A(n207), .B(a[3]), .ZN(n313) );
  OAI22_X1 U298 ( .A1(n314), .A2(n312), .B1(n221), .B2(n315), .ZN(n93) );
  XNOR2_X1 U299 ( .A(b[2]), .B(a[3]), .ZN(n314) );
  OAI22_X1 U300 ( .A1(n315), .A2(n284), .B1(n221), .B2(n316), .ZN(n92) );
  XNOR2_X1 U301 ( .A(b[3]), .B(a[3]), .ZN(n315) );
  OAI22_X1 U302 ( .A1(n316), .A2(n284), .B1(n221), .B2(n317), .ZN(n91) );
  XNOR2_X1 U303 ( .A(b[4]), .B(a[3]), .ZN(n316) );
  OAI22_X1 U304 ( .A1(n319), .A2(n221), .B1(n312), .B2(n319), .ZN(n318) );
  NOR2_X1 U305 ( .A1(n320), .A2(n293), .ZN(n88) );
  OAI22_X1 U306 ( .A1(n321), .A2(n322), .B1(n320), .B2(n323), .ZN(n87) );
  XNOR2_X1 U307 ( .A(a[5]), .B(n286), .ZN(n321) );
  OAI22_X1 U308 ( .A1(n323), .A2(n322), .B1(n320), .B2(n324), .ZN(n86) );
  XNOR2_X1 U309 ( .A(n207), .B(a[5]), .ZN(n323) );
  OAI22_X1 U310 ( .A1(n324), .A2(n322), .B1(n320), .B2(n325), .ZN(n85) );
  XNOR2_X1 U311 ( .A(b[2]), .B(a[5]), .ZN(n324) );
  OAI22_X1 U312 ( .A1(n325), .A2(n322), .B1(n320), .B2(n326), .ZN(n84) );
  XNOR2_X1 U313 ( .A(b[3]), .B(a[5]), .ZN(n325) );
  OAI22_X1 U314 ( .A1(n326), .A2(n322), .B1(n320), .B2(n327), .ZN(n83) );
  XNOR2_X1 U315 ( .A(b[4]), .B(a[5]), .ZN(n326) );
  OAI22_X1 U316 ( .A1(n327), .A2(n322), .B1(n320), .B2(n328), .ZN(n82) );
  XNOR2_X1 U317 ( .A(b[5]), .B(a[5]), .ZN(n327) );
  OAI22_X1 U318 ( .A1(n330), .A2(n320), .B1(n322), .B2(n330), .ZN(n329) );
  NOR2_X1 U319 ( .A1(n331), .A2(n293), .ZN(n80) );
  OAI22_X1 U320 ( .A1(n332), .A2(n333), .B1(n331), .B2(n334), .ZN(n79) );
  XNOR2_X1 U321 ( .A(a[7]), .B(n286), .ZN(n332) );
  OAI22_X1 U322 ( .A1(n335), .A2(n333), .B1(n331), .B2(n336), .ZN(n77) );
  OAI22_X1 U323 ( .A1(n336), .A2(n333), .B1(n331), .B2(n337), .ZN(n76) );
  XNOR2_X1 U324 ( .A(n278), .B(a[7]), .ZN(n336) );
  OAI22_X1 U325 ( .A1(n337), .A2(n333), .B1(n331), .B2(n338), .ZN(n75) );
  XNOR2_X1 U326 ( .A(b[4]), .B(a[7]), .ZN(n337) );
  OAI22_X1 U327 ( .A1(n338), .A2(n333), .B1(n331), .B2(n339), .ZN(n74) );
  XNOR2_X1 U328 ( .A(b[5]), .B(a[7]), .ZN(n338) );
  OAI22_X1 U329 ( .A1(n341), .A2(n331), .B1(n333), .B2(n341), .ZN(n340) );
  OAI21_X1 U330 ( .B1(n292), .B2(n291), .A(n306), .ZN(n72) );
  OAI21_X1 U331 ( .B1(n302), .B2(n312), .A(n342), .ZN(n71) );
  OR3_X1 U332 ( .A1(n221), .A2(n292), .A3(n302), .ZN(n342) );
  OAI21_X1 U333 ( .B1(n299), .B2(n322), .A(n343), .ZN(n70) );
  OR3_X1 U334 ( .A1(n320), .A2(n292), .A3(n299), .ZN(n343) );
  OAI21_X1 U335 ( .B1(n296), .B2(n333), .A(n344), .ZN(n69) );
  OR3_X1 U336 ( .A1(n331), .A2(n286), .A3(n296), .ZN(n344) );
  XNOR2_X1 U337 ( .A(n345), .B(n346), .ZN(n38) );
  OR2_X1 U338 ( .A1(n345), .A2(n346), .ZN(n37) );
  OAI22_X1 U339 ( .A1(n317), .A2(n312), .B1(n221), .B2(n347), .ZN(n346) );
  XNOR2_X1 U340 ( .A(b[5]), .B(a[3]), .ZN(n317) );
  OAI22_X1 U341 ( .A1(n334), .A2(n333), .B1(n331), .B2(n335), .ZN(n345) );
  XNOR2_X1 U342 ( .A(b[2]), .B(a[7]), .ZN(n335) );
  XNOR2_X1 U343 ( .A(n207), .B(a[7]), .ZN(n334) );
  OAI22_X1 U344 ( .A1(n347), .A2(n284), .B1(n221), .B2(n319), .ZN(n31) );
  XNOR2_X1 U345 ( .A(b[7]), .B(a[3]), .ZN(n319) );
  XNOR2_X1 U346 ( .A(n302), .B(a[2]), .ZN(n348) );
  XNOR2_X1 U347 ( .A(b[6]), .B(a[3]), .ZN(n347) );
  OAI22_X1 U348 ( .A1(n328), .A2(n322), .B1(n320), .B2(n330), .ZN(n21) );
  XNOR2_X1 U349 ( .A(b[7]), .B(a[5]), .ZN(n330) );
  XNOR2_X1 U350 ( .A(n299), .B(a[4]), .ZN(n349) );
  XNOR2_X1 U351 ( .A(b[6]), .B(a[5]), .ZN(n328) );
  OAI22_X1 U352 ( .A1(n339), .A2(n333), .B1(n331), .B2(n341), .ZN(n15) );
  XNOR2_X1 U353 ( .A(b[7]), .B(a[7]), .ZN(n341) );
  XNOR2_X1 U354 ( .A(n296), .B(a[6]), .ZN(n350) );
  XNOR2_X1 U355 ( .A(b[6]), .B(a[7]), .ZN(n339) );
  OAI22_X1 U356 ( .A1(n292), .A2(n306), .B1(n351), .B2(n304), .ZN(n104) );
  OAI22_X1 U357 ( .A1(n258), .A2(n306), .B1(n352), .B2(n304), .ZN(n103) );
  XNOR2_X1 U358 ( .A(b[1]), .B(a[1]), .ZN(n351) );
  OAI22_X1 U359 ( .A1(n352), .A2(n306), .B1(n353), .B2(n304), .ZN(n102) );
  XNOR2_X1 U360 ( .A(b[2]), .B(n283), .ZN(n352) );
  OAI22_X1 U361 ( .A1(n257), .A2(n306), .B1(n354), .B2(n304), .ZN(n101) );
  XNOR2_X1 U362 ( .A(b[3]), .B(n283), .ZN(n353) );
  OAI22_X1 U363 ( .A1(n354), .A2(n306), .B1(n305), .B2(n304), .ZN(n100) );
  XNOR2_X1 U364 ( .A(b[5]), .B(n283), .ZN(n305) );
  XNOR2_X1 U365 ( .A(b[4]), .B(n283), .ZN(n354) );
endmodule


module datapath_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n79;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n79), .CO(carry[2]), .S(SUM[1]) );
  XNOR2_X1 U1 ( .A(B[15]), .B(A[15]), .ZN(n69) );
  CLKBUF_X1 U2 ( .A(B[2]), .Z(n1) );
  NAND3_X1 U3 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n2) );
  NAND3_X1 U4 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n3) );
  NAND3_X1 U5 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n4) );
  CLKBUF_X1 U6 ( .A(n47), .Z(n5) );
  CLKBUF_X1 U7 ( .A(B[6]), .Z(n6) );
  CLKBUF_X1 U8 ( .A(carry[5]), .Z(n7) );
  NAND3_X1 U9 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n8) );
  NAND3_X1 U10 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n9) );
  NAND3_X1 U11 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n10) );
  CLKBUF_X1 U12 ( .A(n76), .Z(n11) );
  CLKBUF_X1 U13 ( .A(n42), .Z(n12) );
  XOR2_X1 U14 ( .A(carry[2]), .B(A[2]), .Z(n13) );
  XOR2_X1 U15 ( .A(n1), .B(n13), .Z(SUM[2]) );
  NAND2_X1 U16 ( .A1(B[2]), .A2(carry[2]), .ZN(n14) );
  NAND2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n15) );
  NAND2_X1 U18 ( .A1(carry[2]), .A2(A[2]), .ZN(n16) );
  NAND3_X1 U19 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[3]) );
  CLKBUF_X1 U20 ( .A(n45), .Z(n17) );
  NAND3_X1 U21 ( .A1(n35), .A2(n36), .A3(n37), .ZN(n18) );
  NAND3_X1 U22 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n19) );
  NAND3_X1 U23 ( .A1(n58), .A2(n59), .A3(n57), .ZN(n20) );
  CLKBUF_X1 U24 ( .A(carry[11]), .Z(n21) );
  NAND3_X1 U25 ( .A1(n75), .A2(n76), .A3(n77), .ZN(n22) );
  NAND3_X1 U26 ( .A1(n75), .A2(n11), .A3(n77), .ZN(n23) );
  CLKBUF_X1 U27 ( .A(carry[8]), .Z(n24) );
  CLKBUF_X1 U28 ( .A(B[3]), .Z(n25) );
  XOR2_X1 U29 ( .A(n25), .B(A[3]), .Z(n26) );
  XOR2_X1 U30 ( .A(n4), .B(n26), .Z(SUM[3]) );
  NAND2_X1 U31 ( .A1(B[3]), .A2(carry[3]), .ZN(n27) );
  NAND2_X1 U32 ( .A1(n3), .A2(A[3]), .ZN(n28) );
  NAND2_X1 U33 ( .A1(B[3]), .A2(A[3]), .ZN(n29) );
  NAND3_X1 U34 ( .A1(n27), .A2(n28), .A3(n29), .ZN(carry[4]) );
  NAND3_X1 U35 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n30) );
  NAND3_X1 U36 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n31) );
  CLKBUF_X1 U37 ( .A(n64), .Z(n32) );
  NAND3_X1 U38 ( .A1(n17), .A2(n46), .A3(n5), .ZN(n33) );
  XOR2_X1 U39 ( .A(B[10]), .B(A[10]), .Z(n34) );
  XOR2_X1 U40 ( .A(n23), .B(n34), .Z(SUM[10]) );
  NAND2_X1 U41 ( .A1(n22), .A2(B[10]), .ZN(n35) );
  NAND2_X1 U42 ( .A1(carry[10]), .A2(A[10]), .ZN(n36) );
  NAND2_X1 U43 ( .A1(B[10]), .A2(A[10]), .ZN(n37) );
  NAND3_X1 U44 ( .A1(n35), .A2(n36), .A3(n37), .ZN(carry[11]) );
  XOR2_X1 U45 ( .A(n33), .B(A[7]), .Z(n38) );
  XOR2_X1 U46 ( .A(B[7]), .B(n38), .Z(SUM[7]) );
  NAND2_X1 U47 ( .A1(B[7]), .A2(n10), .ZN(n39) );
  NAND2_X1 U48 ( .A1(B[7]), .A2(A[7]), .ZN(n40) );
  NAND2_X1 U49 ( .A1(carry[7]), .A2(A[7]), .ZN(n41) );
  NAND3_X1 U50 ( .A1(n39), .A2(n41), .A3(n40), .ZN(carry[8]) );
  NAND3_X1 U51 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n42) );
  CLKBUF_X1 U52 ( .A(n20), .Z(n43) );
  XOR2_X1 U53 ( .A(n6), .B(A[6]), .Z(n44) );
  XOR2_X1 U54 ( .A(n31), .B(n44), .Z(SUM[6]) );
  NAND2_X1 U55 ( .A1(n30), .A2(B[6]), .ZN(n45) );
  NAND2_X1 U56 ( .A1(n30), .A2(A[6]), .ZN(n46) );
  NAND2_X1 U57 ( .A1(B[6]), .A2(A[6]), .ZN(n47) );
  NAND3_X1 U58 ( .A1(n45), .A2(n46), .A3(n47), .ZN(carry[7]) );
  XOR2_X1 U59 ( .A(B[4]), .B(A[4]), .Z(n48) );
  XOR2_X1 U60 ( .A(n9), .B(n48), .Z(SUM[4]) );
  NAND2_X1 U61 ( .A1(n8), .A2(B[4]), .ZN(n49) );
  NAND2_X1 U62 ( .A1(carry[4]), .A2(A[4]), .ZN(n50) );
  NAND2_X1 U63 ( .A1(B[4]), .A2(A[4]), .ZN(n51) );
  NAND3_X1 U64 ( .A1(n49), .A2(n50), .A3(n51), .ZN(carry[5]) );
  XOR2_X1 U65 ( .A(B[5]), .B(A[5]), .Z(n52) );
  XOR2_X1 U66 ( .A(n7), .B(n52), .Z(SUM[5]) );
  NAND2_X1 U67 ( .A1(carry[5]), .A2(B[5]), .ZN(n53) );
  NAND2_X1 U68 ( .A1(n2), .A2(A[5]), .ZN(n54) );
  NAND2_X1 U69 ( .A1(B[5]), .A2(A[5]), .ZN(n55) );
  XOR2_X1 U70 ( .A(B[11]), .B(A[11]), .Z(n56) );
  XOR2_X1 U71 ( .A(n21), .B(n56), .Z(SUM[11]) );
  NAND2_X1 U72 ( .A1(B[11]), .A2(n18), .ZN(n57) );
  NAND2_X1 U73 ( .A1(carry[11]), .A2(A[11]), .ZN(n58) );
  NAND2_X1 U74 ( .A1(B[11]), .A2(A[11]), .ZN(n59) );
  NAND3_X1 U75 ( .A1(n57), .A2(n58), .A3(n59), .ZN(carry[12]) );
  XOR2_X1 U76 ( .A(B[12]), .B(A[12]), .Z(n60) );
  XOR2_X1 U77 ( .A(n43), .B(n60), .Z(SUM[12]) );
  NAND2_X1 U78 ( .A1(n20), .A2(B[12]), .ZN(n61) );
  NAND2_X1 U79 ( .A1(carry[12]), .A2(A[12]), .ZN(n62) );
  NAND2_X1 U80 ( .A1(B[12]), .A2(A[12]), .ZN(n63) );
  NAND3_X1 U81 ( .A1(n61), .A2(n62), .A3(n63), .ZN(carry[13]) );
  NAND3_X1 U82 ( .A1(n73), .A2(n72), .A3(n71), .ZN(n64) );
  XOR2_X1 U83 ( .A(B[13]), .B(A[13]), .Z(n65) );
  XOR2_X1 U84 ( .A(n12), .B(n65), .Z(SUM[13]) );
  NAND2_X1 U85 ( .A1(n42), .A2(B[13]), .ZN(n66) );
  NAND2_X1 U86 ( .A1(carry[13]), .A2(A[13]), .ZN(n67) );
  NAND2_X1 U87 ( .A1(B[13]), .A2(A[13]), .ZN(n68) );
  NAND3_X1 U88 ( .A1(n66), .A2(n67), .A3(n68), .ZN(carry[14]) );
  XNOR2_X1 U89 ( .A(carry[15]), .B(n69), .ZN(SUM[15]) );
  XOR2_X1 U90 ( .A(A[8]), .B(B[8]), .Z(n70) );
  XOR2_X1 U91 ( .A(n70), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U92 ( .A1(A[8]), .A2(B[8]), .ZN(n71) );
  NAND2_X1 U93 ( .A1(carry[8]), .A2(A[8]), .ZN(n72) );
  NAND2_X1 U94 ( .A1(B[8]), .A2(n19), .ZN(n73) );
  NAND3_X1 U95 ( .A1(n72), .A2(n71), .A3(n73), .ZN(carry[9]) );
  XOR2_X1 U96 ( .A(A[9]), .B(B[9]), .Z(n74) );
  XOR2_X1 U97 ( .A(n74), .B(n32), .Z(SUM[9]) );
  NAND2_X1 U98 ( .A1(A[9]), .A2(B[9]), .ZN(n75) );
  NAND2_X1 U99 ( .A1(n64), .A2(A[9]), .ZN(n76) );
  NAND2_X1 U100 ( .A1(B[9]), .A2(carry[9]), .ZN(n77) );
  NAND3_X1 U101 ( .A1(n76), .A2(n75), .A3(n77), .ZN(carry[10]) );
  XOR2_X1 U102 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U103 ( .A1(B[0]), .A2(A[0]), .ZN(n79) );
endmodule


module datapath_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n210, n211, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349;

  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n292), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n291), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n295), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n294), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n297), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  NAND2_X1 U157 ( .A1(n315), .A2(n344), .ZN(n317) );
  INV_X1 U158 ( .A(n15), .ZN(n288) );
  NAND3_X1 U159 ( .A1(n218), .A2(n219), .A3(n220), .ZN(n206) );
  OAI22_X1 U160 ( .A1(n306), .A2(n307), .B1(n255), .B2(n308), .ZN(n207) );
  BUF_X1 U161 ( .A(n12), .Z(n240) );
  CLKBUF_X1 U162 ( .A(b[1]), .Z(n208) );
  XOR2_X1 U163 ( .A(n209), .B(n210), .Z(product[8]) );
  AND3_X1 U164 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n209) );
  XNOR2_X1 U165 ( .A(n34), .B(n39), .ZN(n210) );
  AND2_X1 U166 ( .A1(n95), .A2(n102), .ZN(n211) );
  AND3_X1 U167 ( .A1(n267), .A2(n268), .A3(n269), .ZN(product[15]) );
  NAND2_X1 U168 ( .A1(n305), .A2(n343), .ZN(n307) );
  NAND3_X1 U169 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n213) );
  XNOR2_X1 U170 ( .A(n214), .B(n266), .ZN(product[14]) );
  AND3_X1 U171 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n214) );
  XOR2_X1 U172 ( .A(a[5]), .B(a[4]), .Z(n344) );
  XOR2_X1 U173 ( .A(n215), .B(n216), .Z(product[9]) );
  XNOR2_X1 U174 ( .A(n28), .B(n33), .ZN(n215) );
  AND3_X1 U175 ( .A1(n231), .A2(n230), .A3(n232), .ZN(n216) );
  XOR2_X1 U176 ( .A(n19), .B(n18), .Z(n217) );
  XOR2_X1 U177 ( .A(n4), .B(n217), .Z(product[12]) );
  NAND2_X1 U178 ( .A1(n4), .A2(n19), .ZN(n218) );
  NAND2_X1 U179 ( .A1(n4), .A2(n18), .ZN(n219) );
  NAND2_X1 U180 ( .A1(n19), .A2(n18), .ZN(n220) );
  NAND3_X1 U181 ( .A1(n218), .A2(n219), .A3(n220), .ZN(n3) );
  CLKBUF_X1 U182 ( .A(n346), .Z(n233) );
  NAND2_X2 U183 ( .A1(n326), .A2(n345), .ZN(n328) );
  OR2_X2 U184 ( .A1(a[2]), .A2(a[1]), .ZN(n284) );
  XOR2_X1 U185 ( .A(n221), .B(n222), .Z(product[7]) );
  AND3_X1 U186 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n221) );
  XNOR2_X1 U187 ( .A(n40), .B(n45), .ZN(n222) );
  NAND2_X1 U188 ( .A1(n28), .A2(n7), .ZN(n223) );
  XNOR2_X1 U189 ( .A(n240), .B(n224), .ZN(product[4]) );
  XNOR2_X1 U190 ( .A(n54), .B(n211), .ZN(n224) );
  INV_X1 U191 ( .A(a[3]), .ZN(n225) );
  INV_X2 U192 ( .A(n225), .ZN(n226) );
  XNOR2_X1 U193 ( .A(n227), .B(n250), .ZN(product[5]) );
  XNOR2_X1 U194 ( .A(n50), .B(n53), .ZN(n227) );
  XOR2_X1 U195 ( .A(a[3]), .B(a[2]), .Z(n343) );
  NAND3_X1 U196 ( .A1(n238), .A2(n237), .A3(n239), .ZN(n228) );
  NAND3_X1 U197 ( .A1(n230), .A2(n231), .A3(n232), .ZN(n229) );
  NAND2_X1 U198 ( .A1(n228), .A2(n34), .ZN(n230) );
  NAND2_X1 U199 ( .A1(n8), .A2(n39), .ZN(n231) );
  NAND2_X1 U200 ( .A1(n34), .A2(n39), .ZN(n232) );
  NAND3_X1 U201 ( .A1(n230), .A2(n231), .A3(n232), .ZN(n7) );
  NAND3_X1 U202 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n234) );
  NAND3_X1 U203 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n235) );
  NAND3_X1 U204 ( .A1(n279), .A2(n280), .A3(n281), .ZN(n236) );
  NAND2_X1 U205 ( .A1(n236), .A2(n40), .ZN(n237) );
  NAND2_X1 U206 ( .A1(n9), .A2(n45), .ZN(n238) );
  NAND2_X1 U207 ( .A1(n40), .A2(n45), .ZN(n239) );
  NAND3_X1 U208 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n8) );
  XOR2_X1 U209 ( .A(n23), .B(n20), .Z(n241) );
  XOR2_X1 U210 ( .A(n235), .B(n241), .Z(product[11]) );
  NAND2_X1 U211 ( .A1(n234), .A2(n23), .ZN(n242) );
  NAND2_X1 U212 ( .A1(n5), .A2(n20), .ZN(n243) );
  NAND2_X1 U213 ( .A1(n23), .A2(n20), .ZN(n244) );
  NAND3_X1 U214 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n4) );
  XOR2_X1 U215 ( .A(n17), .B(n288), .Z(n245) );
  XOR2_X1 U216 ( .A(n3), .B(n245), .Z(product[13]) );
  NAND2_X1 U217 ( .A1(n206), .A2(n17), .ZN(n246) );
  NAND2_X1 U218 ( .A1(n3), .A2(n288), .ZN(n247) );
  NAND2_X1 U219 ( .A1(n17), .A2(n288), .ZN(n248) );
  NAND3_X1 U220 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n249) );
  NAND3_X1 U221 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n250) );
  NAND3_X1 U222 ( .A1(n258), .A2(n256), .A3(n257), .ZN(n251) );
  NAND3_X1 U223 ( .A1(n223), .A2(n256), .A3(n258), .ZN(n252) );
  CLKBUF_X1 U224 ( .A(b[1]), .Z(n253) );
  NAND2_X1 U225 ( .A1(n283), .A2(n284), .ZN(n254) );
  NAND2_X1 U226 ( .A1(n283), .A2(n284), .ZN(n255) );
  NAND2_X1 U227 ( .A1(n283), .A2(n284), .ZN(n305) );
  NAND2_X2 U228 ( .A1(a[1]), .A2(n299), .ZN(n301) );
  NAND2_X1 U229 ( .A1(n28), .A2(n33), .ZN(n256) );
  NAND2_X1 U230 ( .A1(n28), .A2(n7), .ZN(n257) );
  NAND2_X1 U231 ( .A1(n33), .A2(n229), .ZN(n258) );
  NAND3_X1 U232 ( .A1(n223), .A2(n256), .A3(n258), .ZN(n6) );
  XOR2_X1 U233 ( .A(n24), .B(n27), .Z(n259) );
  XOR2_X1 U234 ( .A(n259), .B(n252), .Z(product[10]) );
  NAND2_X1 U235 ( .A1(n24), .A2(n27), .ZN(n260) );
  NAND2_X1 U236 ( .A1(n24), .A2(n251), .ZN(n261) );
  NAND2_X1 U237 ( .A1(n27), .A2(n6), .ZN(n262) );
  NAND3_X1 U238 ( .A1(n262), .A2(n261), .A3(n260), .ZN(n5) );
  NAND3_X1 U239 ( .A1(n277), .A2(n276), .A3(n275), .ZN(n263) );
  NAND3_X1 U240 ( .A1(n275), .A2(n276), .A3(n277), .ZN(n264) );
  BUF_X1 U241 ( .A(n287), .Z(n265) );
  XOR2_X1 U242 ( .A(n289), .B(n15), .Z(n266) );
  NAND2_X1 U243 ( .A1(n213), .A2(n289), .ZN(n267) );
  NAND2_X1 U244 ( .A1(n213), .A2(n15), .ZN(n268) );
  NAND2_X1 U245 ( .A1(n289), .A2(n15), .ZN(n269) );
  CLKBUF_X1 U246 ( .A(b[3]), .Z(n270) );
  XOR2_X1 U247 ( .A(n207), .B(n102), .Z(n56) );
  XNOR2_X1 U248 ( .A(a[4]), .B(a[3]), .ZN(n271) );
  XNOR2_X1 U249 ( .A(a[4]), .B(a[3]), .ZN(n315) );
  NAND2_X1 U250 ( .A1(n12), .A2(n54), .ZN(n272) );
  NAND2_X1 U251 ( .A1(n12), .A2(n211), .ZN(n273) );
  NAND2_X1 U252 ( .A1(n54), .A2(n211), .ZN(n274) );
  NAND3_X1 U253 ( .A1(n273), .A2(n272), .A3(n274), .ZN(n11) );
  NAND2_X1 U254 ( .A1(n50), .A2(n53), .ZN(n275) );
  NAND2_X1 U255 ( .A1(n249), .A2(n50), .ZN(n276) );
  NAND2_X1 U256 ( .A1(n53), .A2(n11), .ZN(n277) );
  NAND3_X1 U257 ( .A1(n277), .A2(n276), .A3(n275), .ZN(n10) );
  XOR2_X1 U258 ( .A(n46), .B(n49), .Z(n278) );
  XOR2_X1 U259 ( .A(n278), .B(n264), .Z(product[6]) );
  NAND2_X1 U260 ( .A1(n46), .A2(n49), .ZN(n279) );
  NAND2_X1 U261 ( .A1(n263), .A2(n46), .ZN(n280) );
  NAND2_X1 U262 ( .A1(n49), .A2(n10), .ZN(n281) );
  NAND3_X1 U263 ( .A1(n281), .A2(n280), .A3(n279), .ZN(n9) );
  INV_X1 U264 ( .A(n287), .ZN(n282) );
  NAND2_X1 U265 ( .A1(a[2]), .A2(a[1]), .ZN(n283) );
  INV_X1 U266 ( .A(n31), .ZN(n294) );
  NAND2_X1 U267 ( .A1(n254), .A2(n343), .ZN(n285) );
  INV_X1 U268 ( .A(n21), .ZN(n291) );
  INV_X1 U269 ( .A(n324), .ZN(n292) );
  INV_X1 U270 ( .A(n335), .ZN(n289) );
  INV_X1 U271 ( .A(n304), .ZN(n297) );
  INV_X1 U272 ( .A(n313), .ZN(n295) );
  INV_X1 U273 ( .A(a[5]), .ZN(n293) );
  INV_X1 U274 ( .A(a[7]), .ZN(n290) );
  INV_X1 U275 ( .A(b[0]), .ZN(n287) );
  INV_X1 U276 ( .A(n226), .ZN(n296) );
  INV_X1 U277 ( .A(a[1]), .ZN(n298) );
  XOR2_X2 U278 ( .A(a[6]), .B(n293), .Z(n326) );
  INV_X1 U279 ( .A(n287), .ZN(n286) );
  INV_X2 U280 ( .A(a[0]), .ZN(n299) );
  NOR2_X1 U281 ( .A1(n299), .A2(n265), .ZN(product[0]) );
  OAI22_X1 U282 ( .A1(n300), .A2(n301), .B1(n302), .B2(n299), .ZN(n99) );
  OAI22_X1 U283 ( .A1(n302), .A2(n301), .B1(n303), .B2(n299), .ZN(n98) );
  XNOR2_X1 U284 ( .A(b[6]), .B(a[1]), .ZN(n302) );
  OAI22_X1 U285 ( .A1(n299), .A2(n303), .B1(n301), .B2(n303), .ZN(n304) );
  XNOR2_X1 U286 ( .A(b[7]), .B(a[1]), .ZN(n303) );
  NOR2_X1 U287 ( .A1(n254), .A2(n265), .ZN(n96) );
  OAI22_X1 U288 ( .A1(n306), .A2(n307), .B1(n255), .B2(n308), .ZN(n95) );
  XNOR2_X1 U289 ( .A(n226), .B(n286), .ZN(n306) );
  OAI22_X1 U290 ( .A1(n308), .A2(n285), .B1(n255), .B2(n309), .ZN(n94) );
  XNOR2_X1 U291 ( .A(n208), .B(a[3]), .ZN(n308) );
  OAI22_X1 U292 ( .A1(n309), .A2(n307), .B1(n254), .B2(n310), .ZN(n93) );
  XNOR2_X1 U293 ( .A(b[2]), .B(n226), .ZN(n309) );
  OAI22_X1 U294 ( .A1(n310), .A2(n285), .B1(n255), .B2(n311), .ZN(n92) );
  XNOR2_X1 U295 ( .A(b[3]), .B(n226), .ZN(n310) );
  OAI22_X1 U296 ( .A1(n311), .A2(n285), .B1(n255), .B2(n312), .ZN(n91) );
  XNOR2_X1 U297 ( .A(b[4]), .B(n226), .ZN(n311) );
  OAI22_X1 U298 ( .A1(n314), .A2(n254), .B1(n307), .B2(n314), .ZN(n313) );
  NOR2_X1 U299 ( .A1(n271), .A2(n265), .ZN(n88) );
  OAI22_X1 U300 ( .A1(n316), .A2(n317), .B1(n271), .B2(n318), .ZN(n87) );
  XNOR2_X1 U301 ( .A(a[5]), .B(n282), .ZN(n316) );
  OAI22_X1 U302 ( .A1(n318), .A2(n317), .B1(n271), .B2(n319), .ZN(n86) );
  XNOR2_X1 U303 ( .A(n253), .B(a[5]), .ZN(n318) );
  OAI22_X1 U304 ( .A1(n319), .A2(n317), .B1(n271), .B2(n320), .ZN(n85) );
  XNOR2_X1 U305 ( .A(b[2]), .B(a[5]), .ZN(n319) );
  OAI22_X1 U306 ( .A1(n320), .A2(n317), .B1(n271), .B2(n321), .ZN(n84) );
  XNOR2_X1 U307 ( .A(n270), .B(a[5]), .ZN(n320) );
  OAI22_X1 U308 ( .A1(n321), .A2(n317), .B1(n271), .B2(n322), .ZN(n83) );
  XNOR2_X1 U309 ( .A(b[4]), .B(a[5]), .ZN(n321) );
  OAI22_X1 U310 ( .A1(n322), .A2(n317), .B1(n271), .B2(n323), .ZN(n82) );
  XNOR2_X1 U311 ( .A(b[5]), .B(a[5]), .ZN(n322) );
  OAI22_X1 U312 ( .A1(n325), .A2(n271), .B1(n317), .B2(n325), .ZN(n324) );
  NOR2_X1 U313 ( .A1(n326), .A2(n265), .ZN(n80) );
  OAI22_X1 U314 ( .A1(n327), .A2(n328), .B1(n326), .B2(n329), .ZN(n79) );
  XNOR2_X1 U315 ( .A(a[7]), .B(n282), .ZN(n327) );
  OAI22_X1 U316 ( .A1(n330), .A2(n328), .B1(n326), .B2(n331), .ZN(n77) );
  OAI22_X1 U317 ( .A1(n331), .A2(n328), .B1(n326), .B2(n332), .ZN(n76) );
  XNOR2_X1 U318 ( .A(n270), .B(a[7]), .ZN(n331) );
  OAI22_X1 U319 ( .A1(n332), .A2(n328), .B1(n326), .B2(n333), .ZN(n75) );
  XNOR2_X1 U320 ( .A(b[4]), .B(a[7]), .ZN(n332) );
  OAI22_X1 U321 ( .A1(n333), .A2(n328), .B1(n326), .B2(n334), .ZN(n74) );
  XNOR2_X1 U322 ( .A(b[5]), .B(a[7]), .ZN(n333) );
  OAI22_X1 U323 ( .A1(n336), .A2(n326), .B1(n328), .B2(n336), .ZN(n335) );
  OAI21_X1 U324 ( .B1(n286), .B2(n298), .A(n301), .ZN(n72) );
  OAI21_X1 U325 ( .B1(n296), .B2(n307), .A(n337), .ZN(n71) );
  OR3_X1 U326 ( .A1(n254), .A2(n282), .A3(n296), .ZN(n337) );
  OAI21_X1 U327 ( .B1(n293), .B2(n317), .A(n338), .ZN(n70) );
  OR3_X1 U328 ( .A1(n271), .A2(n282), .A3(n293), .ZN(n338) );
  OAI21_X1 U329 ( .B1(n290), .B2(n328), .A(n339), .ZN(n69) );
  OR3_X1 U330 ( .A1(n326), .A2(n282), .A3(n290), .ZN(n339) );
  XNOR2_X1 U331 ( .A(n340), .B(n341), .ZN(n38) );
  OR2_X1 U332 ( .A1(n340), .A2(n341), .ZN(n37) );
  OAI22_X1 U333 ( .A1(n312), .A2(n285), .B1(n254), .B2(n342), .ZN(n341) );
  XNOR2_X1 U334 ( .A(b[5]), .B(n226), .ZN(n312) );
  OAI22_X1 U335 ( .A1(n329), .A2(n328), .B1(n326), .B2(n330), .ZN(n340) );
  XNOR2_X1 U336 ( .A(b[2]), .B(a[7]), .ZN(n330) );
  XNOR2_X1 U337 ( .A(n253), .B(a[7]), .ZN(n329) );
  OAI22_X1 U338 ( .A1(n342), .A2(n307), .B1(n255), .B2(n314), .ZN(n31) );
  XNOR2_X1 U339 ( .A(b[7]), .B(n226), .ZN(n314) );
  XNOR2_X1 U340 ( .A(b[6]), .B(n226), .ZN(n342) );
  OAI22_X1 U341 ( .A1(n323), .A2(n317), .B1(n271), .B2(n325), .ZN(n21) );
  XNOR2_X1 U342 ( .A(b[7]), .B(a[5]), .ZN(n325) );
  XNOR2_X1 U343 ( .A(b[6]), .B(a[5]), .ZN(n323) );
  OAI22_X1 U344 ( .A1(n334), .A2(n328), .B1(n326), .B2(n336), .ZN(n15) );
  XNOR2_X1 U345 ( .A(b[7]), .B(a[7]), .ZN(n336) );
  XNOR2_X1 U346 ( .A(n290), .B(a[6]), .ZN(n345) );
  XNOR2_X1 U347 ( .A(b[6]), .B(a[7]), .ZN(n334) );
  OAI22_X1 U348 ( .A1(n286), .A2(n301), .B1(n346), .B2(n299), .ZN(n104) );
  OAI22_X1 U349 ( .A1(n233), .A2(n301), .B1(n347), .B2(n299), .ZN(n103) );
  XNOR2_X1 U350 ( .A(b[1]), .B(a[1]), .ZN(n346) );
  OAI22_X1 U351 ( .A1(n347), .A2(n301), .B1(n348), .B2(n299), .ZN(n102) );
  XNOR2_X1 U352 ( .A(b[2]), .B(a[1]), .ZN(n347) );
  OAI22_X1 U353 ( .A1(n348), .A2(n301), .B1(n349), .B2(n299), .ZN(n101) );
  XNOR2_X1 U354 ( .A(b[3]), .B(a[1]), .ZN(n348) );
  OAI22_X1 U355 ( .A1(n349), .A2(n301), .B1(n300), .B2(n299), .ZN(n100) );
  XNOR2_X1 U356 ( .A(b[5]), .B(a[1]), .ZN(n300) );
  XNOR2_X1 U357 ( .A(b[4]), .B(a[1]), .ZN(n349) );
endmodule


module datapath_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n76;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n76), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(B[13]), .Z(n1) );
  NAND3_X1 U2 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n2) );
  NAND3_X1 U3 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n3) );
  CLKBUF_X1 U4 ( .A(n28), .Z(n4) );
  CLKBUF_X1 U5 ( .A(n47), .Z(n5) );
  NAND3_X1 U6 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n6) );
  NAND3_X1 U7 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n7) );
  CLKBUF_X1 U8 ( .A(n63), .Z(n8) );
  CLKBUF_X1 U9 ( .A(n22), .Z(n9) );
  NAND3_X1 U10 ( .A1(n21), .A2(n9), .A3(n23), .ZN(n10) );
  NAND3_X1 U11 ( .A1(n17), .A2(n19), .A3(n18), .ZN(n11) );
  NAND3_X1 U12 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n12) );
  NAND3_X1 U13 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n13) );
  NAND3_X1 U14 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n14) );
  NAND3_X1 U15 ( .A1(n8), .A2(n64), .A3(n65), .ZN(n15) );
  XOR2_X1 U16 ( .A(n15), .B(A[11]), .Z(n16) );
  XOR2_X1 U17 ( .A(B[11]), .B(n16), .Z(SUM[11]) );
  NAND2_X1 U18 ( .A1(B[11]), .A2(n14), .ZN(n17) );
  NAND2_X1 U19 ( .A1(B[11]), .A2(A[11]), .ZN(n18) );
  NAND2_X1 U20 ( .A1(carry[11]), .A2(A[11]), .ZN(n19) );
  NAND3_X1 U21 ( .A1(n17), .A2(n19), .A3(n18), .ZN(carry[12]) );
  XOR2_X1 U22 ( .A(B[6]), .B(A[6]), .Z(n20) );
  XOR2_X1 U23 ( .A(carry[6]), .B(n20), .Z(SUM[6]) );
  NAND2_X1 U24 ( .A1(n2), .A2(B[6]), .ZN(n21) );
  NAND2_X1 U25 ( .A1(n12), .A2(A[6]), .ZN(n22) );
  NAND2_X1 U26 ( .A1(B[6]), .A2(A[6]), .ZN(n23) );
  NAND3_X1 U27 ( .A1(n21), .A2(n22), .A3(n23), .ZN(carry[7]) );
  XOR2_X1 U28 ( .A(carry[2]), .B(A[2]), .Z(n24) );
  XOR2_X1 U29 ( .A(B[2]), .B(n24), .Z(SUM[2]) );
  NAND2_X1 U30 ( .A1(B[2]), .A2(carry[2]), .ZN(n25) );
  NAND2_X1 U31 ( .A1(B[2]), .A2(A[2]), .ZN(n26) );
  NAND2_X1 U32 ( .A1(carry[2]), .A2(A[2]), .ZN(n27) );
  NAND3_X1 U33 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[3]) );
  NAND3_X1 U34 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n28) );
  CLKBUF_X1 U35 ( .A(n52), .Z(n29) );
  NAND3_X1 U36 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n30) );
  NAND3_X1 U37 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n31) );
  XOR2_X1 U38 ( .A(B[3]), .B(A[3]), .Z(n32) );
  XOR2_X1 U39 ( .A(n7), .B(n32), .Z(SUM[3]) );
  NAND2_X1 U40 ( .A1(n6), .A2(B[3]), .ZN(n33) );
  NAND2_X1 U41 ( .A1(carry[3]), .A2(A[3]), .ZN(n34) );
  NAND2_X1 U42 ( .A1(B[3]), .A2(A[3]), .ZN(n35) );
  NAND3_X1 U43 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[4]) );
  CLKBUF_X1 U44 ( .A(carry[13]), .Z(n36) );
  NAND3_X1 U45 ( .A1(n60), .A2(n59), .A3(n61), .ZN(n37) );
  XOR2_X1 U46 ( .A(B[7]), .B(A[7]), .Z(n38) );
  XOR2_X1 U47 ( .A(n10), .B(n38), .Z(SUM[7]) );
  NAND2_X1 U48 ( .A1(carry[7]), .A2(B[7]), .ZN(n39) );
  NAND2_X1 U49 ( .A1(n13), .A2(A[7]), .ZN(n40) );
  NAND2_X1 U50 ( .A1(B[7]), .A2(A[7]), .ZN(n41) );
  NAND3_X1 U51 ( .A1(n39), .A2(n40), .A3(n41), .ZN(carry[8]) );
  XOR2_X1 U52 ( .A(B[4]), .B(A[4]), .Z(n42) );
  XOR2_X1 U53 ( .A(carry[4]), .B(n42), .Z(SUM[4]) );
  NAND2_X1 U54 ( .A1(n31), .A2(B[4]), .ZN(n43) );
  NAND2_X1 U55 ( .A1(n31), .A2(A[4]), .ZN(n44) );
  NAND2_X1 U56 ( .A1(B[4]), .A2(A[4]), .ZN(n45) );
  NAND3_X1 U57 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[5]) );
  XOR2_X1 U58 ( .A(B[5]), .B(A[5]), .Z(n46) );
  XOR2_X1 U59 ( .A(n30), .B(n46), .Z(SUM[5]) );
  NAND2_X1 U60 ( .A1(B[5]), .A2(n30), .ZN(n47) );
  NAND2_X1 U61 ( .A1(carry[5]), .A2(A[5]), .ZN(n48) );
  NAND2_X1 U62 ( .A1(B[5]), .A2(A[5]), .ZN(n49) );
  NAND3_X1 U63 ( .A1(n5), .A2(n48), .A3(n49), .ZN(carry[6]) );
  NAND3_X1 U64 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n50) );
  XOR2_X1 U65 ( .A(B[8]), .B(A[8]), .Z(n51) );
  XOR2_X1 U66 ( .A(n4), .B(n51), .Z(SUM[8]) );
  NAND2_X1 U67 ( .A1(n28), .A2(B[8]), .ZN(n52) );
  NAND2_X1 U68 ( .A1(carry[8]), .A2(A[8]), .ZN(n53) );
  NAND2_X1 U69 ( .A1(B[8]), .A2(A[8]), .ZN(n54) );
  NAND3_X1 U70 ( .A1(n29), .A2(n53), .A3(n54), .ZN(carry[9]) );
  CLKBUF_X1 U71 ( .A(n11), .Z(n55) );
  CLKBUF_X1 U72 ( .A(n37), .Z(n56) );
  NAND3_X1 U73 ( .A1(n70), .A2(n69), .A3(n68), .ZN(n57) );
  XOR2_X1 U74 ( .A(B[9]), .B(A[9]), .Z(n58) );
  XOR2_X1 U75 ( .A(carry[9]), .B(n58), .Z(SUM[9]) );
  NAND2_X1 U76 ( .A1(n3), .A2(B[9]), .ZN(n59) );
  NAND2_X1 U77 ( .A1(n50), .A2(A[9]), .ZN(n60) );
  NAND2_X1 U78 ( .A1(B[9]), .A2(A[9]), .ZN(n61) );
  NAND3_X1 U79 ( .A1(n59), .A2(n60), .A3(n61), .ZN(carry[10]) );
  XOR2_X1 U80 ( .A(B[10]), .B(A[10]), .Z(n62) );
  XOR2_X1 U81 ( .A(n56), .B(n62), .Z(SUM[10]) );
  NAND2_X1 U82 ( .A1(n37), .A2(B[10]), .ZN(n63) );
  NAND2_X1 U83 ( .A1(carry[10]), .A2(A[10]), .ZN(n64) );
  NAND2_X1 U84 ( .A1(B[10]), .A2(A[10]), .ZN(n65) );
  NAND3_X1 U85 ( .A1(n63), .A2(n64), .A3(n65), .ZN(carry[11]) );
  NAND2_X1 U86 ( .A1(B[12]), .A2(A[12]), .ZN(n68) );
  XNOR2_X1 U87 ( .A(carry[15]), .B(n66), .ZN(SUM[15]) );
  XNOR2_X1 U88 ( .A(B[15]), .B(A[15]), .ZN(n66) );
  XOR2_X1 U89 ( .A(A[12]), .B(B[12]), .Z(n67) );
  XOR2_X1 U90 ( .A(n67), .B(n55), .Z(SUM[12]) );
  NAND2_X1 U91 ( .A1(A[12]), .A2(carry[12]), .ZN(n69) );
  NAND2_X1 U92 ( .A1(n11), .A2(B[12]), .ZN(n70) );
  NAND3_X1 U93 ( .A1(n70), .A2(n69), .A3(n68), .ZN(carry[13]) );
  XOR2_X1 U94 ( .A(A[13]), .B(n1), .Z(n71) );
  XOR2_X1 U95 ( .A(n71), .B(n36), .Z(SUM[13]) );
  NAND2_X1 U96 ( .A1(B[13]), .A2(A[13]), .ZN(n72) );
  NAND2_X1 U97 ( .A1(carry[13]), .A2(A[13]), .ZN(n73) );
  NAND2_X1 U98 ( .A1(B[13]), .A2(n57), .ZN(n74) );
  NAND3_X1 U99 ( .A1(n74), .A2(n72), .A3(n73), .ZN(carry[14]) );
  XOR2_X1 U100 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U101 ( .A1(B[0]), .A2(A[0]), .ZN(n76) );
endmodule


module datapath ( clk, data_in, addr_x, wr_en_x, addr_a1, addr_a2, addr_a3, 
        addr_a4, addr_a5, addr_a6, addr_a7, addr_a8, addr_a9, addr_a10, 
        addr_a11, addr_a12, addr_a13, addr_a14, addr_a15, addr_a16, wr_en_a1, 
        wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6, wr_en_a7, wr_en_a8, 
        wr_en_a9, wr_en_a10, wr_en_a11, wr_en_a12, wr_en_a13, wr_en_a14, 
        wr_en_a15, wr_en_a16, addr_y, wr_en_y, clear_acc, clc, clc1, data_out
 );
  input [7:0] data_in;
  input [3:0] addr_x;
  input [3:0] addr_a1;
  input [3:0] addr_a2;
  input [3:0] addr_a3;
  input [3:0] addr_a4;
  input [3:0] addr_a5;
  input [3:0] addr_a6;
  input [3:0] addr_a7;
  input [3:0] addr_a8;
  input [3:0] addr_a9;
  input [3:0] addr_a10;
  input [3:0] addr_a11;
  input [3:0] addr_a12;
  input [3:0] addr_a13;
  input [3:0] addr_a14;
  input [3:0] addr_a15;
  input [3:0] addr_a16;
  input [3:0] addr_y;
  output [15:0] data_out;
  input clk, wr_en_x, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5,
         wr_en_a6, wr_en_a7, wr_en_a8, wr_en_a9, wr_en_a10, wr_en_a11,
         wr_en_a12, wr_en_a13, wr_en_a14, wr_en_a15, wr_en_a16, wr_en_y,
         clear_acc, clc, clc1;
  wire   n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, \mul_out1[9] ,
         \mul_out1[8] , \mul_out1[7] , \mul_out1[6] , \mul_out1[5] ,
         \mul_out1[4] , \mul_out1[3] , \mul_out1[2] , \mul_out1[1] ,
         \mul_out1[15] , \mul_out1[14] , \mul_out1[13] , \mul_out1[12] ,
         \mul_out1[11] , \mul_out1[10] , \mul_out1[0] , \mul_out2[9] ,
         \mul_out2[8] , \mul_out2[7] , \mul_out2[6] , \mul_out2[5] ,
         \mul_out2[4] , \mul_out2[3] , \mul_out2[2] , \mul_out2[1] ,
         \mul_out2[15] , \mul_out2[14] , \mul_out2[13] , \mul_out2[12] ,
         \mul_out2[11] , \mul_out2[10] , \mul_out2[0] , \mul_out3[9] ,
         \mul_out3[8] , \mul_out3[7] , \mul_out3[6] , \mul_out3[5] ,
         \mul_out3[4] , \mul_out3[3] , \mul_out3[2] , \mul_out3[1] ,
         \mul_out3[15] , \mul_out3[14] , \mul_out3[13] , \mul_out3[12] ,
         \mul_out3[11] , \mul_out3[10] , \mul_out3[0] , \mul_out4[9] ,
         \mul_out4[8] , \mul_out4[7] , \mul_out4[6] , \mul_out4[5] ,
         \mul_out4[4] , \mul_out4[3] , \mul_out4[2] , \mul_out4[1] ,
         \mul_out4[15] , \mul_out4[14] , \mul_out4[13] , \mul_out4[12] ,
         \mul_out4[11] , \mul_out4[10] , \mul_out4[0] , \mul_out5[9] ,
         \mul_out5[8] , \mul_out5[7] , \mul_out5[6] , \mul_out5[5] ,
         \mul_out5[4] , \mul_out5[3] , \mul_out5[2] , \mul_out5[1] ,
         \mul_out5[15] , \mul_out5[14] , \mul_out5[13] , \mul_out5[12] ,
         \mul_out5[11] , \mul_out5[10] , \mul_out5[0] , \mul_out6[9] ,
         \mul_out6[8] , \mul_out6[7] , \mul_out6[6] , \mul_out6[5] ,
         \mul_out6[4] , \mul_out6[3] , \mul_out6[2] , \mul_out6[1] ,
         \mul_out6[15] , \mul_out6[14] , \mul_out6[13] , \mul_out6[12] ,
         \mul_out6[11] , \mul_out6[10] , \mul_out6[0] , \mul_out7[9] ,
         \mul_out7[8] , \mul_out7[7] , \mul_out7[6] , \mul_out7[5] ,
         \mul_out7[4] , \mul_out7[3] , \mul_out7[2] , \mul_out7[1] ,
         \mul_out7[15] , \mul_out7[14] , \mul_out7[13] , \mul_out7[12] ,
         \mul_out7[11] , \mul_out7[10] , \mul_out7[0] , \mul_out8[9] ,
         \mul_out8[8] , \mul_out8[7] , \mul_out8[6] , \mul_out8[5] ,
         \mul_out8[4] , \mul_out8[3] , \mul_out8[2] , \mul_out8[1] ,
         \mul_out8[15] , \mul_out8[14] , \mul_out8[13] , \mul_out8[12] ,
         \mul_out8[11] , \mul_out8[10] , \mul_out8[0] , \mul_out9[9] ,
         \mul_out9[8] , \mul_out9[7] , \mul_out9[6] , \mul_out9[5] ,
         \mul_out9[4] , \mul_out9[3] , \mul_out9[2] , \mul_out9[1] ,
         \mul_out9[15] , \mul_out9[14] , \mul_out9[13] , \mul_out9[12] ,
         \mul_out9[11] , \mul_out9[10] , \mul_out9[0] , \mul_out10[9] ,
         \mul_out10[8] , \mul_out10[7] , \mul_out10[6] , \mul_out10[5] ,
         \mul_out10[4] , \mul_out10[3] , \mul_out10[2] , \mul_out10[1] ,
         \mul_out10[15] , \mul_out10[14] , \mul_out10[13] , \mul_out10[12] ,
         \mul_out10[11] , \mul_out10[10] , \mul_out10[0] , \mul_out11[9] ,
         \mul_out11[8] , \mul_out11[7] , \mul_out11[6] , \mul_out11[5] ,
         \mul_out11[4] , \mul_out11[3] , \mul_out11[2] , \mul_out11[1] ,
         \mul_out11[15] , \mul_out11[14] , \mul_out11[13] , \mul_out11[12] ,
         \mul_out11[11] , \mul_out11[10] , \mul_out11[0] , \mul_out12[9] ,
         \mul_out12[8] , \mul_out12[7] , \mul_out12[6] , \mul_out12[5] ,
         \mul_out12[4] , \mul_out12[3] , \mul_out12[2] , \mul_out12[1] ,
         \mul_out12[15] , \mul_out12[14] , \mul_out12[13] , \mul_out12[12] ,
         \mul_out12[11] , \mul_out12[10] , \mul_out12[0] , \mul_out13[9] ,
         \mul_out13[8] , \mul_out13[7] , \mul_out13[6] , \mul_out13[5] ,
         \mul_out13[4] , \mul_out13[3] , \mul_out13[2] , \mul_out13[1] ,
         \mul_out13[15] , \mul_out13[14] , \mul_out13[13] , \mul_out13[12] ,
         \mul_out13[11] , \mul_out13[10] , \mul_out13[0] , \mul_out14[9] ,
         \mul_out14[8] , \mul_out14[7] , \mul_out14[6] , \mul_out14[5] ,
         \mul_out14[4] , \mul_out14[3] , \mul_out14[2] , \mul_out14[1] ,
         \mul_out14[15] , \mul_out14[14] , \mul_out14[13] , \mul_out14[12] ,
         \mul_out14[11] , \mul_out14[10] , \mul_out14[0] , \mul_out15[9] ,
         \mul_out15[8] , \mul_out15[7] , \mul_out15[6] , \mul_out15[5] ,
         \mul_out15[4] , \mul_out15[3] , \mul_out15[2] , \mul_out15[1] ,
         \mul_out15[15] , \mul_out15[14] , \mul_out15[13] , \mul_out15[12] ,
         \mul_out15[11] , \mul_out15[10] , \mul_out15[0] , \mul_out16[9] ,
         \mul_out16[8] , \mul_out16[7] , \mul_out16[6] , \mul_out16[5] ,
         \mul_out16[4] , \mul_out16[3] , \mul_out16[2] , \mul_out16[1] ,
         \mul_out16[15] , \mul_out16[14] , \mul_out16[13] , \mul_out16[12] ,
         \mul_out16[11] , \mul_out16[10] , \mul_out16[0] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101;
  wire   [7:0] data_out_x;
  wire   [7:0] data_out_a1;
  wire   [7:0] data_out_a2;
  wire   [7:0] data_out_a3;
  wire   [7:0] data_out_a4;
  wire   [7:0] data_out_a5;
  wire   [7:0] data_out_a6;
  wire   [7:0] data_out_a7;
  wire   [7:0] data_out_a8;
  wire   [7:0] data_out_a9;
  wire   [7:0] data_out_a10;
  wire   [7:0] data_out_a11;
  wire   [7:0] data_out_a12;
  wire   [7:0] data_out_a13;
  wire   [7:0] data_out_a14;
  wire   [7:0] data_out_a15;
  wire   [7:0] data_out_a16;
  wire   [15:0] f;
  wire   [15:0] f1;
  wire   [15:0] f2;
  wire   [15:0] f3;
  wire   [15:0] f4;
  wire   [15:0] f5;
  wire   [15:0] f6;
  wire   [15:0] f7;
  wire   [15:0] f8;
  wire   [15:0] f9;
  wire   [15:0] f10;
  wire   [15:0] f11;
  wire   [15:0] f12;
  wire   [15:0] f13;
  wire   [15:0] f14;
  wire   [15:0] f15;
  wire   [15:0] f16;
  wire   [15:0] add_r1;
  wire   [15:0] add_r2;
  wire   [15:0] add_r3;
  wire   [15:0] add_r4;
  wire   [15:0] add_r5;
  wire   [15:0] add_r6;
  wire   [15:0] add_r7;
  wire   [15:0] add_r8;
  wire   [15:0] add_r9;
  wire   [15:0] add_r10;
  wire   [15:0] add_r11;
  wire   [15:0] add_r12;
  wire   [15:0] add_r13;
  wire   [15:0] add_r14;
  wire   [15:0] add_r15;
  wire   [15:0] add_r16;

  DFF_X1 \f1_reg[15]  ( .D(n1020), .CK(clk), .Q(f1[15]), .QN(n17) );
  DFF_X1 \f1_reg[14]  ( .D(n1019), .CK(clk), .Q(f1[14]), .QN(n18) );
  DFF_X1 \f1_reg[11]  ( .D(n1016), .CK(clk), .Q(f1[11]), .QN(n21) );
  DFF_X1 \f1_reg[10]  ( .D(n1015), .CK(clk), .Q(f1[10]), .QN(n22) );
  DFF_X1 \f1_reg[9]  ( .D(n1014), .CK(clk), .Q(f1[9]), .QN(n23) );
  DFF_X1 \f1_reg[8]  ( .D(n1013), .CK(clk), .Q(f1[8]), .QN(n24) );
  DFF_X1 \f1_reg[7]  ( .D(n1012), .CK(clk), .Q(f1[7]), .QN(n25) );
  DFF_X1 \f1_reg[6]  ( .D(n1011), .CK(clk), .Q(f1[6]), .QN(n26) );
  DFF_X1 \f1_reg[5]  ( .D(n1010), .CK(clk), .Q(f1[5]), .QN(n27) );
  DFF_X1 \f1_reg[4]  ( .D(n1009), .CK(clk), .Q(f1[4]), .QN(n28) );
  DFF_X1 \f1_reg[3]  ( .D(n1008), .CK(clk), .Q(f1[3]), .QN(n29) );
  DFF_X1 \f1_reg[2]  ( .D(n1007), .CK(clk), .Q(f1[2]), .QN(n30) );
  DFF_X1 \f1_reg[1]  ( .D(n1006), .CK(clk), .Q(f1[1]), .QN(n31) );
  DFF_X1 \f1_reg[0]  ( .D(n1005), .CK(clk), .Q(f1[0]), .QN(n32) );
  DFF_X1 \f2_reg[14]  ( .D(n1003), .CK(clk), .Q(f2[14]), .QN(n34) );
  DFF_X1 \f2_reg[13]  ( .D(n1002), .CK(clk), .Q(f2[13]), .QN(n35) );
  DFF_X1 \f2_reg[12]  ( .D(n1001), .CK(clk), .Q(f2[12]), .QN(n36) );
  DFF_X1 \f2_reg[11]  ( .D(n1000), .CK(clk), .Q(f2[11]), .QN(n37) );
  DFF_X1 \f2_reg[10]  ( .D(n999), .CK(clk), .Q(f2[10]), .QN(n38) );
  DFF_X1 \f2_reg[9]  ( .D(n998), .CK(clk), .Q(f2[9]), .QN(n39) );
  DFF_X1 \f2_reg[8]  ( .D(n997), .CK(clk), .Q(f2[8]), .QN(n40) );
  DFF_X1 \f2_reg[7]  ( .D(n996), .CK(clk), .Q(f2[7]), .QN(n41) );
  DFF_X1 \f2_reg[6]  ( .D(n995), .CK(clk), .Q(f2[6]), .QN(n42) );
  DFF_X1 \f2_reg[5]  ( .D(n994), .CK(clk), .Q(f2[5]), .QN(n43) );
  DFF_X1 \f2_reg[4]  ( .D(n993), .CK(clk), .Q(f2[4]), .QN(n44) );
  DFF_X1 \f2_reg[3]  ( .D(n992), .CK(clk), .Q(f2[3]), .QN(n45) );
  DFF_X1 \f2_reg[2]  ( .D(n991), .CK(clk), .Q(f2[2]), .QN(n46) );
  DFF_X1 \f2_reg[1]  ( .D(n990), .CK(clk), .Q(f2[1]), .QN(n47) );
  DFF_X1 \f2_reg[0]  ( .D(n989), .CK(clk), .Q(f2[0]), .QN(n48) );
  DFF_X1 \f3_reg[14]  ( .D(n987), .CK(clk), .Q(f3[14]), .QN(n50) );
  DFF_X1 \f3_reg[13]  ( .D(n986), .CK(clk), .Q(f3[13]), .QN(n51) );
  DFF_X1 \f3_reg[12]  ( .D(n985), .CK(clk), .Q(f3[12]), .QN(n52) );
  DFF_X1 \f3_reg[11]  ( .D(n984), .CK(clk), .Q(f3[11]), .QN(n53) );
  DFF_X1 \f3_reg[10]  ( .D(n983), .CK(clk), .Q(f3[10]), .QN(n54) );
  DFF_X1 \f3_reg[9]  ( .D(n982), .CK(clk), .Q(f3[9]), .QN(n55) );
  DFF_X1 \f3_reg[8]  ( .D(n981), .CK(clk), .Q(f3[8]), .QN(n56) );
  DFF_X1 \f3_reg[7]  ( .D(n980), .CK(clk), .Q(f3[7]), .QN(n57) );
  DFF_X1 \f3_reg[6]  ( .D(n979), .CK(clk), .Q(f3[6]), .QN(n58) );
  DFF_X1 \f3_reg[5]  ( .D(n978), .CK(clk), .Q(f3[5]), .QN(n59) );
  DFF_X1 \f3_reg[4]  ( .D(n977), .CK(clk), .Q(f3[4]), .QN(n60) );
  DFF_X1 \f3_reg[3]  ( .D(n976), .CK(clk), .Q(f3[3]), .QN(n61) );
  DFF_X1 \f3_reg[2]  ( .D(n975), .CK(clk), .Q(f3[2]), .QN(n62) );
  DFF_X1 \f3_reg[1]  ( .D(n974), .CK(clk), .Q(f3[1]), .QN(n63) );
  DFF_X1 \f3_reg[0]  ( .D(n973), .CK(clk), .Q(f3[0]), .QN(n64) );
  DFF_X1 \f4_reg[13]  ( .D(n970), .CK(clk), .Q(f4[13]), .QN(n67) );
  DFF_X1 \f4_reg[12]  ( .D(n969), .CK(clk), .Q(f4[12]), .QN(n68) );
  DFF_X1 \f4_reg[11]  ( .D(n968), .CK(clk), .Q(f4[11]), .QN(n69) );
  DFF_X1 \f4_reg[10]  ( .D(n967), .CK(clk), .Q(f4[10]), .QN(n70) );
  DFF_X1 \f4_reg[9]  ( .D(n966), .CK(clk), .Q(f4[9]), .QN(n71) );
  DFF_X1 \f4_reg[8]  ( .D(n965), .CK(clk), .Q(f4[8]), .QN(n72) );
  DFF_X1 \f4_reg[7]  ( .D(n964), .CK(clk), .Q(f4[7]), .QN(n73) );
  DFF_X1 \f4_reg[6]  ( .D(n963), .CK(clk), .Q(f4[6]), .QN(n74) );
  DFF_X1 \f4_reg[5]  ( .D(n962), .CK(clk), .Q(f4[5]), .QN(n75) );
  DFF_X1 \f4_reg[4]  ( .D(n961), .CK(clk), .Q(f4[4]), .QN(n76) );
  DFF_X1 \f4_reg[3]  ( .D(n960), .CK(clk), .Q(f4[3]), .QN(n77) );
  DFF_X1 \f4_reg[2]  ( .D(n959), .CK(clk), .Q(f4[2]), .QN(n78) );
  DFF_X1 \f4_reg[1]  ( .D(n958), .CK(clk), .Q(f4[1]), .QN(n79) );
  DFF_X1 \f4_reg[0]  ( .D(n957), .CK(clk), .Q(f4[0]), .QN(n80) );
  DFF_X1 \f5_reg[14]  ( .D(n955), .CK(clk), .Q(f5[14]), .QN(n82) );
  DFF_X1 \f5_reg[13]  ( .D(n954), .CK(clk), .Q(f5[13]), .QN(n83) );
  DFF_X1 \f5_reg[12]  ( .D(n953), .CK(clk), .Q(f5[12]), .QN(n84) );
  DFF_X1 \f5_reg[11]  ( .D(n952), .CK(clk), .Q(f5[11]), .QN(n85) );
  DFF_X1 \f5_reg[10]  ( .D(n951), .CK(clk), .Q(f5[10]), .QN(n86) );
  DFF_X1 \f5_reg[9]  ( .D(n950), .CK(clk), .Q(f5[9]), .QN(n87) );
  DFF_X1 \f5_reg[8]  ( .D(n949), .CK(clk), .Q(f5[8]), .QN(n88) );
  DFF_X1 \f5_reg[7]  ( .D(n948), .CK(clk), .Q(f5[7]), .QN(n89) );
  DFF_X1 \f5_reg[6]  ( .D(n947), .CK(clk), .Q(f5[6]), .QN(n90) );
  DFF_X1 \f5_reg[5]  ( .D(n946), .CK(clk), .Q(f5[5]), .QN(n91) );
  DFF_X1 \f5_reg[4]  ( .D(n945), .CK(clk), .Q(f5[4]), .QN(n92) );
  DFF_X1 \f5_reg[3]  ( .D(n944), .CK(clk), .Q(f5[3]), .QN(n93) );
  DFF_X1 \f5_reg[2]  ( .D(n943), .CK(clk), .Q(f5[2]), .QN(n94) );
  DFF_X1 \f5_reg[1]  ( .D(n942), .CK(clk), .Q(f5[1]), .QN(n95) );
  DFF_X1 \f5_reg[0]  ( .D(n941), .CK(clk), .Q(f5[0]), .QN(n96) );
  DFF_X1 \f6_reg[13]  ( .D(n938), .CK(clk), .Q(f6[13]), .QN(n99) );
  DFF_X1 \f6_reg[12]  ( .D(n937), .CK(clk), .Q(f6[12]), .QN(n100) );
  DFF_X1 \f6_reg[11]  ( .D(n936), .CK(clk), .Q(f6[11]), .QN(n101) );
  DFF_X1 \f6_reg[10]  ( .D(n935), .CK(clk), .Q(f6[10]), .QN(n102) );
  DFF_X1 \f6_reg[9]  ( .D(n934), .CK(clk), .Q(f6[9]), .QN(n103) );
  DFF_X1 \f6_reg[8]  ( .D(n933), .CK(clk), .Q(f6[8]), .QN(n104) );
  DFF_X1 \f6_reg[7]  ( .D(n932), .CK(clk), .Q(f6[7]), .QN(n105) );
  DFF_X1 \f6_reg[6]  ( .D(n931), .CK(clk), .Q(f6[6]), .QN(n106) );
  DFF_X1 \f6_reg[5]  ( .D(n930), .CK(clk), .Q(f6[5]), .QN(n107) );
  DFF_X1 \f6_reg[4]  ( .D(n929), .CK(clk), .Q(f6[4]), .QN(n108) );
  DFF_X1 \f6_reg[3]  ( .D(n928), .CK(clk), .Q(f6[3]), .QN(n109) );
  DFF_X1 \f6_reg[2]  ( .D(n927), .CK(clk), .Q(f6[2]), .QN(n110) );
  DFF_X1 \f6_reg[1]  ( .D(n926), .CK(clk), .Q(f6[1]), .QN(n111) );
  DFF_X1 \f6_reg[0]  ( .D(n925), .CK(clk), .Q(f6[0]), .QN(n112) );
  DFF_X1 \f7_reg[14]  ( .D(n923), .CK(clk), .Q(f7[14]), .QN(n114) );
  DFF_X1 \f7_reg[13]  ( .D(n922), .CK(clk), .Q(f7[13]), .QN(n115) );
  DFF_X1 \f7_reg[12]  ( .D(n921), .CK(clk), .Q(f7[12]), .QN(n116) );
  DFF_X1 \f7_reg[11]  ( .D(n920), .CK(clk), .Q(f7[11]), .QN(n117) );
  DFF_X1 \f7_reg[10]  ( .D(n919), .CK(clk), .Q(f7[10]), .QN(n118) );
  DFF_X1 \f7_reg[9]  ( .D(n918), .CK(clk), .Q(f7[9]), .QN(n119) );
  DFF_X1 \f7_reg[8]  ( .D(n917), .CK(clk), .Q(f7[8]), .QN(n120) );
  DFF_X1 \f7_reg[7]  ( .D(n916), .CK(clk), .Q(f7[7]), .QN(n121) );
  DFF_X1 \f7_reg[6]  ( .D(n915), .CK(clk), .Q(f7[6]), .QN(n122) );
  DFF_X1 \f7_reg[5]  ( .D(n914), .CK(clk), .Q(f7[5]), .QN(n123) );
  DFF_X1 \f7_reg[4]  ( .D(n913), .CK(clk), .Q(f7[4]), .QN(n124) );
  DFF_X1 \f7_reg[3]  ( .D(n912), .CK(clk), .Q(f7[3]), .QN(n125) );
  DFF_X1 \f7_reg[2]  ( .D(n911), .CK(clk), .Q(f7[2]), .QN(n126) );
  DFF_X1 \f7_reg[1]  ( .D(n910), .CK(clk), .Q(f7[1]), .QN(n127) );
  DFF_X1 \f7_reg[0]  ( .D(n909), .CK(clk), .Q(f7[0]), .QN(n128) );
  DFF_X1 \f8_reg[14]  ( .D(n907), .CK(clk), .Q(f8[14]), .QN(n130) );
  DFF_X1 \f8_reg[13]  ( .D(n906), .CK(clk), .Q(f8[13]), .QN(n131) );
  DFF_X1 \f8_reg[12]  ( .D(n905), .CK(clk), .Q(f8[12]), .QN(n132) );
  DFF_X1 \f8_reg[11]  ( .D(n904), .CK(clk), .Q(f8[11]), .QN(n133) );
  DFF_X1 \f8_reg[10]  ( .D(n903), .CK(clk), .Q(f8[10]), .QN(n134) );
  DFF_X1 \f8_reg[9]  ( .D(n902), .CK(clk), .Q(f8[9]), .QN(n135) );
  DFF_X1 \f8_reg[8]  ( .D(n901), .CK(clk), .Q(f8[8]), .QN(n136) );
  DFF_X1 \f8_reg[7]  ( .D(n900), .CK(clk), .Q(f8[7]), .QN(n137) );
  DFF_X1 \f8_reg[6]  ( .D(n899), .CK(clk), .Q(f8[6]), .QN(n138) );
  DFF_X1 \f8_reg[5]  ( .D(n898), .CK(clk), .Q(f8[5]), .QN(n139) );
  DFF_X1 \f8_reg[4]  ( .D(n897), .CK(clk), .Q(f8[4]), .QN(n140) );
  DFF_X1 \f8_reg[3]  ( .D(n896), .CK(clk), .Q(f8[3]), .QN(n141) );
  DFF_X1 \f8_reg[2]  ( .D(n895), .CK(clk), .Q(f8[2]), .QN(n142) );
  DFF_X1 \f8_reg[1]  ( .D(n894), .CK(clk), .Q(f8[1]), .QN(n143) );
  DFF_X1 \f8_reg[0]  ( .D(n893), .CK(clk), .Q(f8[0]), .QN(n144) );
  DFF_X1 \f9_reg[15]  ( .D(n892), .CK(clk), .Q(f9[15]), .QN(n145) );
  DFF_X1 \f9_reg[14]  ( .D(n891), .CK(clk), .Q(f9[14]), .QN(n146) );
  DFF_X1 \f9_reg[13]  ( .D(n890), .CK(clk), .Q(f9[13]), .QN(n147) );
  DFF_X1 \f9_reg[12]  ( .D(n889), .CK(clk), .Q(f9[12]), .QN(n148) );
  DFF_X1 \f9_reg[11]  ( .D(n888), .CK(clk), .Q(f9[11]), .QN(n149) );
  DFF_X1 \f9_reg[10]  ( .D(n887), .CK(clk), .Q(f9[10]), .QN(n150) );
  DFF_X1 \f9_reg[9]  ( .D(n886), .CK(clk), .Q(f9[9]), .QN(n151) );
  DFF_X1 \f9_reg[8]  ( .D(n885), .CK(clk), .Q(f9[8]), .QN(n152) );
  DFF_X1 \f9_reg[7]  ( .D(n884), .CK(clk), .Q(f9[7]), .QN(n153) );
  DFF_X1 \f9_reg[6]  ( .D(n883), .CK(clk), .Q(f9[6]), .QN(n154) );
  DFF_X1 \f9_reg[5]  ( .D(n882), .CK(clk), .Q(f9[5]), .QN(n155) );
  DFF_X1 \f9_reg[4]  ( .D(n881), .CK(clk), .Q(f9[4]), .QN(n156) );
  DFF_X1 \f9_reg[3]  ( .D(n880), .CK(clk), .Q(f9[3]), .QN(n157) );
  DFF_X1 \f9_reg[2]  ( .D(n879), .CK(clk), .Q(f9[2]), .QN(n158) );
  DFF_X1 \f9_reg[1]  ( .D(n878), .CK(clk), .Q(f9[1]), .QN(n159) );
  DFF_X1 \f9_reg[0]  ( .D(n877), .CK(clk), .Q(f9[0]), .QN(n160) );
  DFF_X1 \f10_reg[14]  ( .D(n875), .CK(clk), .Q(f10[14]), .QN(n162) );
  DFF_X1 \f10_reg[13]  ( .D(n874), .CK(clk), .Q(f10[13]), .QN(n163) );
  DFF_X1 \f10_reg[12]  ( .D(n873), .CK(clk), .Q(f10[12]), .QN(n164) );
  DFF_X1 \f10_reg[11]  ( .D(n872), .CK(clk), .Q(f10[11]), .QN(n165) );
  DFF_X1 \f10_reg[10]  ( .D(n871), .CK(clk), .Q(f10[10]), .QN(n166) );
  DFF_X1 \f10_reg[9]  ( .D(n870), .CK(clk), .Q(f10[9]), .QN(n167) );
  DFF_X1 \f10_reg[8]  ( .D(n869), .CK(clk), .Q(f10[8]), .QN(n168) );
  DFF_X1 \f10_reg[7]  ( .D(n868), .CK(clk), .Q(f10[7]), .QN(n169) );
  DFF_X1 \f10_reg[6]  ( .D(n867), .CK(clk), .Q(f10[6]), .QN(n170) );
  DFF_X1 \f10_reg[5]  ( .D(n866), .CK(clk), .Q(f10[5]), .QN(n171) );
  DFF_X1 \f10_reg[4]  ( .D(n865), .CK(clk), .Q(f10[4]), .QN(n172) );
  DFF_X1 \f10_reg[3]  ( .D(n864), .CK(clk), .Q(f10[3]), .QN(n173) );
  DFF_X1 \f10_reg[2]  ( .D(n863), .CK(clk), .Q(f10[2]), .QN(n174) );
  DFF_X1 \f10_reg[1]  ( .D(n862), .CK(clk), .Q(f10[1]), .QN(n175) );
  DFF_X1 \f10_reg[0]  ( .D(n861), .CK(clk), .Q(f10[0]), .QN(n176) );
  DFF_X1 \f11_reg[14]  ( .D(n859), .CK(clk), .Q(f11[14]), .QN(n178) );
  DFF_X1 \f11_reg[13]  ( .D(n858), .CK(clk), .Q(f11[13]), .QN(n179) );
  DFF_X1 \f11_reg[12]  ( .D(n857), .CK(clk), .Q(f11[12]), .QN(n180) );
  DFF_X1 \f11_reg[11]  ( .D(n856), .CK(clk), .Q(f11[11]), .QN(n181) );
  DFF_X1 \f11_reg[10]  ( .D(n855), .CK(clk), .Q(f11[10]), .QN(n182) );
  DFF_X1 \f11_reg[9]  ( .D(n854), .CK(clk), .Q(f11[9]), .QN(n183) );
  DFF_X1 \f11_reg[8]  ( .D(n853), .CK(clk), .Q(f11[8]), .QN(n184) );
  DFF_X1 \f11_reg[7]  ( .D(n852), .CK(clk), .Q(f11[7]), .QN(n185) );
  DFF_X1 \f11_reg[6]  ( .D(n851), .CK(clk), .Q(f11[6]), .QN(n186) );
  DFF_X1 \f11_reg[5]  ( .D(n850), .CK(clk), .Q(f11[5]), .QN(n187) );
  DFF_X1 \f11_reg[4]  ( .D(n849), .CK(clk), .Q(f11[4]), .QN(n188) );
  DFF_X1 \f11_reg[3]  ( .D(n848), .CK(clk), .Q(f11[3]), .QN(n189) );
  DFF_X1 \f11_reg[2]  ( .D(n847), .CK(clk), .Q(f11[2]), .QN(n190) );
  DFF_X1 \f11_reg[1]  ( .D(n846), .CK(clk), .Q(f11[1]), .QN(n191) );
  DFF_X1 \f11_reg[0]  ( .D(n845), .CK(clk), .Q(f11[0]), .QN(n192) );
  DFF_X1 \f12_reg[14]  ( .D(n843), .CK(clk), .Q(f12[14]), .QN(n194) );
  DFF_X1 \f12_reg[13]  ( .D(n842), .CK(clk), .Q(f12[13]), .QN(n195) );
  DFF_X1 \f12_reg[12]  ( .D(n841), .CK(clk), .Q(f12[12]), .QN(n196) );
  DFF_X1 \f12_reg[11]  ( .D(n840), .CK(clk), .Q(f12[11]), .QN(n197) );
  DFF_X1 \f12_reg[10]  ( .D(n839), .CK(clk), .Q(f12[10]), .QN(n198) );
  DFF_X1 \f12_reg[9]  ( .D(n838), .CK(clk), .Q(f12[9]), .QN(n199) );
  DFF_X1 \f12_reg[8]  ( .D(n837), .CK(clk), .Q(f12[8]), .QN(n200) );
  DFF_X1 \f12_reg[7]  ( .D(n836), .CK(clk), .Q(f12[7]), .QN(n201) );
  DFF_X1 \f12_reg[6]  ( .D(n835), .CK(clk), .Q(f12[6]), .QN(n202) );
  DFF_X1 \f12_reg[5]  ( .D(n834), .CK(clk), .Q(f12[5]), .QN(n203) );
  DFF_X1 \f12_reg[4]  ( .D(n833), .CK(clk), .Q(f12[4]), .QN(n204) );
  DFF_X1 \f12_reg[3]  ( .D(n832), .CK(clk), .Q(f12[3]), .QN(n205) );
  DFF_X1 \f12_reg[2]  ( .D(n831), .CK(clk), .Q(f12[2]), .QN(n206) );
  DFF_X1 \f12_reg[1]  ( .D(n830), .CK(clk), .Q(f12[1]), .QN(n207) );
  DFF_X1 \f12_reg[0]  ( .D(n829), .CK(clk), .Q(f12[0]), .QN(n208) );
  DFF_X1 \f13_reg[14]  ( .D(n827), .CK(clk), .Q(f13[14]), .QN(n210) );
  DFF_X1 \f13_reg[13]  ( .D(n826), .CK(clk), .Q(f13[13]), .QN(n211) );
  DFF_X1 \f13_reg[12]  ( .D(n825), .CK(clk), .Q(f13[12]), .QN(n212) );
  DFF_X1 \f13_reg[11]  ( .D(n824), .CK(clk), .Q(f13[11]), .QN(n213) );
  DFF_X1 \f13_reg[10]  ( .D(n823), .CK(clk), .Q(f13[10]), .QN(n214) );
  DFF_X1 \f13_reg[9]  ( .D(n822), .CK(clk), .Q(f13[9]), .QN(n215) );
  DFF_X1 \f13_reg[8]  ( .D(n821), .CK(clk), .Q(f13[8]), .QN(n216) );
  DFF_X1 \f13_reg[7]  ( .D(n820), .CK(clk), .Q(f13[7]), .QN(n217) );
  DFF_X1 \f13_reg[6]  ( .D(n819), .CK(clk), .Q(f13[6]), .QN(n218) );
  DFF_X1 \f13_reg[5]  ( .D(n818), .CK(clk), .Q(f13[5]), .QN(n219) );
  DFF_X1 \f13_reg[4]  ( .D(n817), .CK(clk), .Q(f13[4]), .QN(n220) );
  DFF_X1 \f13_reg[3]  ( .D(n816), .CK(clk), .Q(f13[3]), .QN(n221) );
  DFF_X1 \f13_reg[2]  ( .D(n815), .CK(clk), .Q(f13[2]), .QN(n222) );
  DFF_X1 \f13_reg[1]  ( .D(n814), .CK(clk), .Q(f13[1]), .QN(n223) );
  DFF_X1 \f13_reg[0]  ( .D(n813), .CK(clk), .Q(f13[0]), .QN(n224) );
  DFF_X1 \f14_reg[14]  ( .D(n811), .CK(clk), .Q(f14[14]), .QN(n226) );
  DFF_X1 \f14_reg[13]  ( .D(n810), .CK(clk), .Q(f14[13]), .QN(n227) );
  DFF_X1 \f14_reg[12]  ( .D(n809), .CK(clk), .Q(f14[12]), .QN(n228) );
  DFF_X1 \f14_reg[11]  ( .D(n808), .CK(clk), .Q(f14[11]), .QN(n229) );
  DFF_X1 \f14_reg[10]  ( .D(n807), .CK(clk), .Q(f14[10]), .QN(n230) );
  DFF_X1 \f14_reg[9]  ( .D(n806), .CK(clk), .Q(f14[9]), .QN(n231) );
  DFF_X1 \f14_reg[8]  ( .D(n805), .CK(clk), .Q(f14[8]), .QN(n232) );
  DFF_X1 \f14_reg[7]  ( .D(n804), .CK(clk), .Q(f14[7]), .QN(n233) );
  DFF_X1 \f14_reg[6]  ( .D(n803), .CK(clk), .Q(f14[6]), .QN(n234) );
  DFF_X1 \f14_reg[5]  ( .D(n802), .CK(clk), .Q(f14[5]), .QN(n235) );
  DFF_X1 \f14_reg[4]  ( .D(n801), .CK(clk), .Q(f14[4]), .QN(n236) );
  DFF_X1 \f14_reg[3]  ( .D(n800), .CK(clk), .Q(f14[3]), .QN(n237) );
  DFF_X1 \f14_reg[2]  ( .D(n799), .CK(clk), .Q(f14[2]), .QN(n238) );
  DFF_X1 \f14_reg[1]  ( .D(n798), .CK(clk), .Q(f14[1]), .QN(n239) );
  DFF_X1 \f14_reg[0]  ( .D(n797), .CK(clk), .Q(f14[0]), .QN(n240) );
  DFF_X1 \f15_reg[15]  ( .D(n796), .CK(clk), .Q(f15[15]), .QN(n241) );
  DFF_X1 \f15_reg[14]  ( .D(n795), .CK(clk), .Q(f15[14]), .QN(n242) );
  DFF_X1 \f15_reg[13]  ( .D(n794), .CK(clk), .Q(f15[13]), .QN(n243) );
  DFF_X1 \f15_reg[12]  ( .D(n793), .CK(clk), .Q(f15[12]), .QN(n244) );
  DFF_X1 \f15_reg[11]  ( .D(n792), .CK(clk), .Q(f15[11]), .QN(n245) );
  DFF_X1 \f15_reg[10]  ( .D(n791), .CK(clk), .Q(f15[10]), .QN(n246) );
  DFF_X1 \f15_reg[9]  ( .D(n790), .CK(clk), .Q(f15[9]), .QN(n247) );
  DFF_X1 \f15_reg[8]  ( .D(n789), .CK(clk), .Q(f15[8]), .QN(n248) );
  DFF_X1 \f15_reg[7]  ( .D(n788), .CK(clk), .Q(f15[7]), .QN(n249) );
  DFF_X1 \f15_reg[6]  ( .D(n787), .CK(clk), .Q(f15[6]), .QN(n250) );
  DFF_X1 \f15_reg[5]  ( .D(n786), .CK(clk), .Q(f15[5]), .QN(n251) );
  DFF_X1 \f15_reg[4]  ( .D(n785), .CK(clk), .Q(f15[4]), .QN(n252) );
  DFF_X1 \f15_reg[3]  ( .D(n784), .CK(clk), .Q(f15[3]), .QN(n253) );
  DFF_X1 \f15_reg[2]  ( .D(n783), .CK(clk), .Q(f15[2]), .QN(n254) );
  DFF_X1 \f15_reg[1]  ( .D(n782), .CK(clk), .Q(f15[1]), .QN(n255) );
  DFF_X1 \f15_reg[0]  ( .D(n781), .CK(clk), .Q(f15[0]), .QN(n256) );
  DFF_X1 \f16_reg[15]  ( .D(n780), .CK(clk), .Q(f16[15]), .QN(n257) );
  DFF_X1 \f_reg[15]  ( .D(n749), .CK(clk), .Q(f[15]) );
  DFF_X1 \f16_reg[14]  ( .D(n779), .CK(clk), .Q(f16[14]), .QN(n258) );
  DFF_X1 \f_reg[14]  ( .D(n750), .CK(clk), .Q(f[14]) );
  DFF_X1 \f16_reg[13]  ( .D(n778), .CK(clk), .Q(f16[13]), .QN(n259) );
  DFF_X1 \f_reg[13]  ( .D(n751), .CK(clk), .Q(f[13]) );
  DFF_X1 \f16_reg[12]  ( .D(n777), .CK(clk), .Q(f16[12]), .QN(n260) );
  DFF_X1 \f_reg[12]  ( .D(n752), .CK(clk), .Q(f[12]) );
  DFF_X1 \f16_reg[11]  ( .D(n776), .CK(clk), .Q(f16[11]), .QN(n261) );
  DFF_X1 \f_reg[11]  ( .D(n753), .CK(clk), .Q(f[11]) );
  DFF_X1 \f16_reg[10]  ( .D(n775), .CK(clk), .Q(f16[10]), .QN(n262) );
  DFF_X1 \f_reg[10]  ( .D(n754), .CK(clk), .Q(f[10]) );
  DFF_X1 \f16_reg[9]  ( .D(n774), .CK(clk), .Q(f16[9]), .QN(n263) );
  DFF_X1 \f_reg[9]  ( .D(n755), .CK(clk), .Q(f[9]) );
  DFF_X1 \f16_reg[8]  ( .D(n773), .CK(clk), .Q(f16[8]), .QN(n264) );
  DFF_X1 \f_reg[8]  ( .D(n756), .CK(clk), .Q(f[8]) );
  DFF_X1 \f16_reg[7]  ( .D(n772), .CK(clk), .Q(f16[7]), .QN(n265) );
  DFF_X1 \f_reg[7]  ( .D(n757), .CK(clk), .Q(f[7]) );
  DFF_X1 \f16_reg[6]  ( .D(n771), .CK(clk), .Q(f16[6]), .QN(n266) );
  DFF_X1 \f_reg[6]  ( .D(n758), .CK(clk), .Q(f[6]) );
  DFF_X1 \f16_reg[5]  ( .D(n770), .CK(clk), .Q(f16[5]), .QN(n267) );
  DFF_X1 \f_reg[5]  ( .D(n759), .CK(clk), .Q(f[5]) );
  DFF_X1 \f16_reg[4]  ( .D(n769), .CK(clk), .Q(f16[4]), .QN(n268) );
  DFF_X1 \f_reg[4]  ( .D(n760), .CK(clk), .Q(f[4]) );
  DFF_X1 \f16_reg[3]  ( .D(n768), .CK(clk), .Q(f16[3]), .QN(n269) );
  DFF_X1 \f_reg[3]  ( .D(n761), .CK(clk), .Q(f[3]) );
  DFF_X1 \f16_reg[2]  ( .D(n767), .CK(clk), .Q(f16[2]), .QN(n270) );
  DFF_X1 \f_reg[2]  ( .D(n762), .CK(clk), .Q(f[2]) );
  DFF_X1 \f16_reg[1]  ( .D(n766), .CK(clk), .Q(f16[1]), .QN(n271) );
  DFF_X1 \f_reg[1]  ( .D(n763), .CK(clk), .Q(f[1]) );
  DFF_X1 \f16_reg[0]  ( .D(n765), .CK(clk), .Q(f16[0]), .QN(n272) );
  DFF_X1 \f_reg[0]  ( .D(n764), .CK(clk), .Q(f[0]) );
  NOR2_X2 U185 ( .A1(n1099), .A2(n293), .ZN(n290) );
  memory_WIDTH8_SIZE16_LOGSIZE4_0 mem_x ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_x), .addr(addr_x), .wr_en(wr_en_x) );
  memory_WIDTH8_SIZE16_LOGSIZE4_16 mem_a1 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a1), .addr(addr_a1), .wr_en(wr_en_a1) );
  memory_WIDTH8_SIZE16_LOGSIZE4_15 mem_a2 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a2), .addr(addr_a2), .wr_en(wr_en_a2) );
  memory_WIDTH8_SIZE16_LOGSIZE4_14 mem_a3 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a3), .addr(addr_a3), .wr_en(wr_en_a3) );
  memory_WIDTH8_SIZE16_LOGSIZE4_13 mem_a4 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a4), .addr(addr_a4), .wr_en(wr_en_a4) );
  memory_WIDTH8_SIZE16_LOGSIZE4_12 mem_a5 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a5), .addr(addr_a5), .wr_en(wr_en_a5) );
  memory_WIDTH8_SIZE16_LOGSIZE4_11 mem_a6 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a6), .addr(addr_a6), .wr_en(wr_en_a6) );
  memory_WIDTH8_SIZE16_LOGSIZE4_10 mem_a7 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a7), .addr(addr_a7), .wr_en(wr_en_a7) );
  memory_WIDTH8_SIZE16_LOGSIZE4_9 mem_a8 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a8), .addr(addr_a8), .wr_en(wr_en_a8) );
  memory_WIDTH8_SIZE16_LOGSIZE4_8 mem_a9 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a9), .addr(addr_a9), .wr_en(wr_en_a9) );
  memory_WIDTH8_SIZE16_LOGSIZE4_7 mem_a10 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a10), .addr(addr_a10), .wr_en(wr_en_a10) );
  memory_WIDTH8_SIZE16_LOGSIZE4_6 mem_a11 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a11), .addr(addr_a11), .wr_en(wr_en_a11) );
  memory_WIDTH8_SIZE16_LOGSIZE4_5 mem_a12 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a12), .addr(addr_a12), .wr_en(wr_en_a12) );
  memory_WIDTH8_SIZE16_LOGSIZE4_4 mem_a13 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a13), .addr(addr_a13), .wr_en(wr_en_a13) );
  memory_WIDTH8_SIZE16_LOGSIZE4_3 mem_a14 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a14), .addr(addr_a14), .wr_en(wr_en_a14) );
  memory_WIDTH8_SIZE16_LOGSIZE4_2 mem_a15 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a15), .addr(addr_a15), .wr_en(wr_en_a15) );
  memory_WIDTH8_SIZE16_LOGSIZE4_1 mem_a16 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a16), .addr(addr_a16), .wr_en(wr_en_a16) );
  memory_WIDTH16_SIZE16_LOGSIZE4 mem_y ( .clk(clk), .data_in(f), .data_out(
        data_out), .addr(addr_y), .wr_en(wr_en_y) );
  datapath_DW_mult_tc_15 mult_92 ( .a(data_out_a1), .b({n1087, n1085, n1082, 
        n4, n2, n1078, n283, n1073}), .product({\mul_out1[15] , \mul_out1[14] , 
        \mul_out1[13] , \mul_out1[12] , \mul_out1[11] , \mul_out1[10] , 
        \mul_out1[9] , \mul_out1[8] , \mul_out1[7] , \mul_out1[6] , 
        \mul_out1[5] , \mul_out1[4] , \mul_out1[3] , \mul_out1[2] , 
        \mul_out1[1] , \mul_out1[0] }) );
  datapath_DW01_add_15 add_93 ( .A(f1), .B({\mul_out1[15] , \mul_out1[14] , 
        \mul_out1[13] , \mul_out1[12] , \mul_out1[11] , \mul_out1[10] , 
        \mul_out1[9] , \mul_out1[8] , \mul_out1[7] , \mul_out1[6] , 
        \mul_out1[5] , \mul_out1[4] , \mul_out1[3] , \mul_out1[2] , 
        \mul_out1[1] , \mul_out1[0] }), .CI(1'b0), .SUM(add_r1) );
  datapath_DW_mult_tc_14 mult_94 ( .a(data_out_a2), .b({n1087, n1084, n1082, 
        n4, n3, n11, n284, n1073}), .product({\mul_out2[15] , \mul_out2[14] , 
        \mul_out2[13] , \mul_out2[12] , \mul_out2[11] , \mul_out2[10] , 
        \mul_out2[9] , \mul_out2[8] , \mul_out2[7] , \mul_out2[6] , 
        \mul_out2[5] , \mul_out2[4] , \mul_out2[3] , \mul_out2[2] , 
        \mul_out2[1] , \mul_out2[0] }) );
  datapath_DW01_add_14 add_95 ( .A(f2), .B({\mul_out2[15] , \mul_out2[14] , 
        \mul_out2[13] , \mul_out2[12] , \mul_out2[11] , \mul_out2[10] , 
        \mul_out2[9] , \mul_out2[8] , \mul_out2[7] , \mul_out2[6] , 
        \mul_out2[5] , \mul_out2[4] , \mul_out2[3] , \mul_out2[2] , 
        \mul_out2[1] , \mul_out2[0] }), .CI(1'b0), .SUM(add_r2) );
  datapath_DW_mult_tc_13 mult_96 ( .a(data_out_a3), .b({n1087, n1085, n1082, 
        n5, n2, n1078, n283, n1074}), .product({\mul_out3[15] , \mul_out3[14] , 
        \mul_out3[13] , \mul_out3[12] , \mul_out3[11] , \mul_out3[10] , 
        \mul_out3[9] , \mul_out3[8] , \mul_out3[7] , \mul_out3[6] , 
        \mul_out3[5] , \mul_out3[4] , \mul_out3[3] , \mul_out3[2] , 
        \mul_out3[1] , \mul_out3[0] }) );
  datapath_DW01_add_13 add_97 ( .A(f3), .B({\mul_out3[15] , \mul_out3[14] , 
        \mul_out3[13] , \mul_out3[12] , \mul_out3[11] , \mul_out3[10] , 
        \mul_out3[9] , \mul_out3[8] , \mul_out3[7] , \mul_out3[6] , 
        \mul_out3[5] , \mul_out3[4] , \mul_out3[3] , \mul_out3[2] , 
        \mul_out3[1] , \mul_out3[0] }), .CI(1'b0), .SUM(add_r3) );
  datapath_DW_mult_tc_12 mult_98 ( .a(data_out_a4), .b({n1087, n1084, n1082, 
        n5, n6, n1078, n284, n1074}), .product({\mul_out4[15] , \mul_out4[14] , 
        \mul_out4[13] , \mul_out4[12] , \mul_out4[11] , \mul_out4[10] , 
        \mul_out4[9] , \mul_out4[8] , \mul_out4[7] , \mul_out4[6] , 
        \mul_out4[5] , \mul_out4[4] , \mul_out4[3] , \mul_out4[2] , 
        \mul_out4[1] , \mul_out4[0] }) );
  datapath_DW01_add_12 add_99 ( .A(f4), .B({\mul_out4[15] , \mul_out4[14] , 
        \mul_out4[13] , \mul_out4[12] , \mul_out4[11] , \mul_out4[10] , 
        \mul_out4[9] , \mul_out4[8] , \mul_out4[7] , \mul_out4[6] , 
        \mul_out4[5] , \mul_out4[4] , \mul_out4[3] , \mul_out4[2] , 
        \mul_out4[1] , \mul_out4[0] }), .CI(1'b0), .SUM(add_r4) );
  datapath_DW_mult_tc_11 mult_100 ( .a(data_out_a5), .b({n1086, n1084, n1083, 
        n5, n1079, n10, n1022, n1074}), .product({\mul_out5[15] , 
        \mul_out5[14] , \mul_out5[13] , \mul_out5[12] , \mul_out5[11] , 
        \mul_out5[10] , \mul_out5[9] , \mul_out5[8] , \mul_out5[7] , 
        \mul_out5[6] , \mul_out5[5] , \mul_out5[4] , \mul_out5[3] , 
        \mul_out5[2] , \mul_out5[1] , \mul_out5[0] }) );
  datapath_DW01_add_11 add_101 ( .A(f5), .B({\mul_out5[15] , \mul_out5[14] , 
        \mul_out5[13] , \mul_out5[12] , \mul_out5[11] , \mul_out5[10] , 
        \mul_out5[9] , \mul_out5[8] , \mul_out5[7] , \mul_out5[6] , 
        \mul_out5[5] , \mul_out5[4] , \mul_out5[3] , \mul_out5[2] , 
        \mul_out5[1] , \mul_out5[0] }), .CI(1'b0), .SUM(add_r5) );
  datapath_DW_mult_tc_10 mult_102 ( .a(data_out_a6), .b({n1086, n1084, n1082, 
        n1081, n3, n11, n1075, n9}), .product({\mul_out6[15] , \mul_out6[14] , 
        \mul_out6[13] , \mul_out6[12] , \mul_out6[11] , \mul_out6[10] , 
        \mul_out6[9] , \mul_out6[8] , \mul_out6[7] , \mul_out6[6] , 
        \mul_out6[5] , \mul_out6[4] , \mul_out6[3] , \mul_out6[2] , 
        \mul_out6[1] , \mul_out6[0] }) );
  datapath_DW01_add_10 add_103 ( .A(f6), .B({\mul_out6[15] , \mul_out6[14] , 
        \mul_out6[13] , \mul_out6[12] , \mul_out6[11] , \mul_out6[10] , 
        \mul_out6[9] , \mul_out6[8] , \mul_out6[7] , \mul_out6[6] , 
        \mul_out6[5] , \mul_out6[4] , \mul_out6[3] , \mul_out6[2] , 
        \mul_out6[1] , \mul_out6[0] }), .CI(1'b0), .SUM(add_r6) );
  datapath_DW_mult_tc_9 mult_104 ( .a(data_out_a7), .b({n1086, n1084, n1082, 
        n4, n7, n10, n1076, n1073}), .product({\mul_out7[15] , \mul_out7[14] , 
        \mul_out7[13] , \mul_out7[12] , \mul_out7[11] , \mul_out7[10] , 
        \mul_out7[9] , \mul_out7[8] , \mul_out7[7] , \mul_out7[6] , 
        \mul_out7[5] , \mul_out7[4] , \mul_out7[3] , \mul_out7[2] , 
        \mul_out7[1] , \mul_out7[0] }) );
  datapath_DW01_add_9 add_105 ( .A(f7), .B({\mul_out7[15] , \mul_out7[14] , 
        \mul_out7[13] , \mul_out7[12] , \mul_out7[11] , \mul_out7[10] , 
        \mul_out7[9] , \mul_out7[8] , \mul_out7[7] , \mul_out7[6] , 
        \mul_out7[5] , \mul_out7[4] , \mul_out7[3] , \mul_out7[2] , 
        \mul_out7[1] , \mul_out7[0] }), .CI(1'b0), .SUM(add_r7) );
  datapath_DW_mult_tc_8 mult_106 ( .a(data_out_a8), .b({n1086, n1084, n1082, 
        n1081, n1080, n14, n1021, n1074}), .product({\mul_out8[15] , 
        \mul_out8[14] , \mul_out8[13] , \mul_out8[12] , \mul_out8[11] , 
        \mul_out8[10] , \mul_out8[9] , \mul_out8[8] , \mul_out8[7] , 
        \mul_out8[6] , \mul_out8[5] , \mul_out8[4] , \mul_out8[3] , 
        \mul_out8[2] , \mul_out8[1] , \mul_out8[0] }) );
  datapath_DW01_add_8 add_107 ( .A(f8), .B({\mul_out8[15] , \mul_out8[14] , 
        \mul_out8[13] , \mul_out8[12] , \mul_out8[11] , \mul_out8[10] , 
        \mul_out8[9] , \mul_out8[8] , \mul_out8[7] , \mul_out8[6] , 
        \mul_out8[5] , \mul_out8[4] , \mul_out8[3] , \mul_out8[2] , 
        \mul_out8[1] , \mul_out8[0] }), .CI(1'b0), .SUM(add_r8) );
  datapath_DW_mult_tc_7 mult_108 ( .a(data_out_a9), .b({n1086, n1085, n1083, 
        n1081, n3, n1078, n283, n1073}), .product({\mul_out9[15] , 
        \mul_out9[14] , \mul_out9[13] , \mul_out9[12] , \mul_out9[11] , 
        \mul_out9[10] , \mul_out9[9] , \mul_out9[8] , \mul_out9[7] , 
        \mul_out9[6] , \mul_out9[5] , \mul_out9[4] , \mul_out9[3] , 
        \mul_out9[2] , \mul_out9[1] , \mul_out9[0] }) );
  datapath_DW01_add_7 add_109 ( .A(f9), .B({\mul_out9[15] , \mul_out9[14] , 
        \mul_out9[13] , \mul_out9[12] , \mul_out9[11] , \mul_out9[10] , 
        \mul_out9[9] , \mul_out9[8] , \mul_out9[7] , \mul_out9[6] , 
        \mul_out9[5] , \mul_out9[4] , \mul_out9[3] , \mul_out9[2] , 
        \mul_out9[1] , \mul_out9[0] }), .CI(1'b0), .SUM(add_r9) );
  datapath_DW_mult_tc_6 mult_110 ( .a(data_out_a10), .b({n1086, n1085, n1083, 
        n5, n1080, n13, n284, n9}), .product({\mul_out10[15] , \mul_out10[14] , 
        \mul_out10[13] , \mul_out10[12] , \mul_out10[11] , \mul_out10[10] , 
        \mul_out10[9] , \mul_out10[8] , \mul_out10[7] , \mul_out10[6] , 
        \mul_out10[5] , \mul_out10[4] , \mul_out10[3] , \mul_out10[2] , 
        \mul_out10[1] , \mul_out10[0] }) );
  datapath_DW01_add_6 add_111 ( .A(f10), .B({\mul_out10[15] , \mul_out10[14] , 
        \mul_out10[13] , \mul_out10[12] , \mul_out10[11] , \mul_out10[10] , 
        \mul_out10[9] , \mul_out10[8] , \mul_out10[7] , \mul_out10[6] , 
        \mul_out10[5] , \mul_out10[4] , \mul_out10[3] , \mul_out10[2] , 
        \mul_out10[1] , \mul_out10[0] }), .CI(1'b0), .SUM(add_r10) );
  datapath_DW_mult_tc_5 mult_112 ( .a(data_out_a11), .b({n1086, n1084, n1083, 
        n4, n1079, n10, n1022, data_out_x[0]}), .product({\mul_out11[15] , 
        \mul_out11[14] , \mul_out11[13] , \mul_out11[12] , \mul_out11[11] , 
        \mul_out11[10] , \mul_out11[9] , \mul_out11[8] , \mul_out11[7] , 
        \mul_out11[6] , \mul_out11[5] , \mul_out11[4] , \mul_out11[3] , 
        \mul_out11[2] , \mul_out11[1] , \mul_out11[0] }) );
  datapath_DW01_add_5 add_113 ( .A(f11), .B({\mul_out11[15] , \mul_out11[14] , 
        \mul_out11[13] , \mul_out11[12] , \mul_out11[11] , \mul_out11[10] , 
        \mul_out11[9] , \mul_out11[8] , \mul_out11[7] , \mul_out11[6] , 
        \mul_out11[5] , \mul_out11[4] , \mul_out11[3] , \mul_out11[2] , 
        \mul_out11[1] , \mul_out11[0] }), .CI(1'b0), .SUM(add_r11) );
  datapath_DW_mult_tc_4 mult_114 ( .a(data_out_a12), .b({n1086, n1085, n1083, 
        n5, n1079, n13, n1022, n1074}), .product({\mul_out12[15] , 
        \mul_out12[14] , \mul_out12[13] , \mul_out12[12] , \mul_out12[11] , 
        \mul_out12[10] , \mul_out12[9] , \mul_out12[8] , \mul_out12[7] , 
        \mul_out12[6] , \mul_out12[5] , \mul_out12[4] , \mul_out12[3] , 
        \mul_out12[2] , \mul_out12[1] , \mul_out12[0] }) );
  datapath_DW01_add_4 add_115 ( .A(f12), .B({\mul_out12[15] , \mul_out12[14] , 
        \mul_out12[13] , \mul_out12[12] , \mul_out12[11] , \mul_out12[10] , 
        \mul_out12[9] , \mul_out12[8] , \mul_out12[7] , \mul_out12[6] , 
        \mul_out12[5] , \mul_out12[4] , \mul_out12[3] , \mul_out12[2] , 
        \mul_out12[1] , \mul_out12[0] }), .CI(1'b0), .SUM(add_r12) );
  datapath_DW_mult_tc_3 mult_116 ( .a(data_out_a13), .b({n1086, n1085, n1083, 
        n5, n7, n13, n1076, n1073}), .product({\mul_out13[15] , 
        \mul_out13[14] , \mul_out13[13] , \mul_out13[12] , \mul_out13[11] , 
        \mul_out13[10] , \mul_out13[9] , \mul_out13[8] , \mul_out13[7] , 
        \mul_out13[6] , \mul_out13[5] , \mul_out13[4] , \mul_out13[3] , 
        \mul_out13[2] , \mul_out13[1] , \mul_out13[0] }) );
  datapath_DW01_add_3 add_117 ( .A(f13), .B({\mul_out13[15] , \mul_out13[14] , 
        \mul_out13[13] , \mul_out13[12] , \mul_out13[11] , \mul_out13[10] , 
        \mul_out13[9] , \mul_out13[8] , \mul_out13[7] , \mul_out13[6] , 
        \mul_out13[5] , \mul_out13[4] , \mul_out13[3] , \mul_out13[2] , 
        \mul_out13[1] , \mul_out13[0] }), .CI(1'b0), .SUM(add_r13) );
  datapath_DW_mult_tc_2 mult_118 ( .a(data_out_a14), .b({n1086, n1085, n1082, 
        n4, n2, n14, n1076, n1073}), .product({\mul_out14[15] , 
        \mul_out14[14] , \mul_out14[13] , \mul_out14[12] , \mul_out14[11] , 
        \mul_out14[10] , \mul_out14[9] , \mul_out14[8] , \mul_out14[7] , 
        \mul_out14[6] , \mul_out14[5] , \mul_out14[4] , \mul_out14[3] , 
        \mul_out14[2] , \mul_out14[1] , \mul_out14[0] }) );
  datapath_DW01_add_2 add_119 ( .A(f14), .B({\mul_out14[15] , \mul_out14[14] , 
        \mul_out14[13] , \mul_out14[12] , \mul_out14[11] , \mul_out14[10] , 
        \mul_out14[9] , \mul_out14[8] , \mul_out14[7] , \mul_out14[6] , 
        \mul_out14[5] , \mul_out14[4] , \mul_out14[3] , \mul_out14[2] , 
        \mul_out14[1] , \mul_out14[0] }), .CI(1'b0), .SUM(add_r14) );
  datapath_DW_mult_tc_1 mult_120 ( .a(data_out_a15), .b({n1086, n1085, n1083, 
        n1081, n1080, n11, n1021, n9}), .product({\mul_out15[15] , 
        \mul_out15[14] , \mul_out15[13] , \mul_out15[12] , \mul_out15[11] , 
        \mul_out15[10] , \mul_out15[9] , \mul_out15[8] , \mul_out15[7] , 
        \mul_out15[6] , \mul_out15[5] , \mul_out15[4] , \mul_out15[3] , 
        \mul_out15[2] , \mul_out15[1] , \mul_out15[0] }) );
  datapath_DW01_add_1 add_121 ( .A(f15), .B({\mul_out15[15] , \mul_out15[14] , 
        \mul_out15[13] , \mul_out15[12] , \mul_out15[11] , \mul_out15[10] , 
        \mul_out15[9] , \mul_out15[8] , \mul_out15[7] , \mul_out15[6] , 
        \mul_out15[5] , \mul_out15[4] , \mul_out15[3] , \mul_out15[2] , 
        \mul_out15[1] , \mul_out15[0] }), .CI(1'b0), .SUM(add_r15) );
  datapath_DW_mult_tc_0 mult_122 ( .a(data_out_a16), .b({n1086, n1085, n1083, 
        n1081, n7, n14, n1021, n1073}), .product({\mul_out16[15] , 
        \mul_out16[14] , \mul_out16[13] , \mul_out16[12] , \mul_out16[11] , 
        \mul_out16[10] , \mul_out16[9] , \mul_out16[8] , \mul_out16[7] , 
        \mul_out16[6] , \mul_out16[5] , \mul_out16[4] , \mul_out16[3] , 
        \mul_out16[2] , \mul_out16[1] , \mul_out16[0] }) );
  datapath_DW01_add_0 add_123 ( .A(f16), .B({\mul_out16[15] , \mul_out16[14] , 
        \mul_out16[13] , \mul_out16[12] , \mul_out16[11] , \mul_out16[10] , 
        \mul_out16[9] , \mul_out16[8] , \mul_out16[7] , \mul_out16[6] , 
        \mul_out16[5] , \mul_out16[4] , \mul_out16[3] , \mul_out16[2] , 
        \mul_out16[1] , \mul_out16[0] }), .CI(1'b0), .SUM(add_r16) );
  DFF_X1 \f12_reg[15]  ( .D(n844), .CK(clk), .Q(f12[15]), .QN(n193) );
  DFF_X1 \f5_reg[15]  ( .D(n956), .CK(clk), .Q(f5[15]), .QN(n81) );
  DFF_X1 \f11_reg[15]  ( .D(n860), .CK(clk), .Q(f11[15]), .QN(n177) );
  DFF_X1 \f3_reg[15]  ( .D(n988), .CK(clk), .Q(f3[15]), .QN(n49) );
  DFF_X1 \f2_reg[15]  ( .D(n1004), .CK(clk), .Q(f2[15]), .QN(n33) );
  DFF_X1 \f4_reg[15]  ( .D(n972), .CK(clk), .Q(f4[15]), .QN(n65) );
  DFF_X1 \f13_reg[15]  ( .D(n828), .CK(clk), .Q(f13[15]), .QN(n209) );
  DFF_X1 \f14_reg[15]  ( .D(n812), .CK(clk), .Q(f14[15]), .QN(n225) );
  DFF_X1 \f7_reg[15]  ( .D(n924), .CK(clk), .Q(f7[15]), .QN(n113) );
  DFF_X1 \f6_reg[15]  ( .D(n940), .CK(clk), .Q(f6[15]), .QN(n97) );
  DFF_X1 \f8_reg[15]  ( .D(n908), .CK(clk), .Q(f8[15]), .QN(n129) );
  DFF_X1 \f10_reg[15]  ( .D(n876), .CK(clk), .Q(f10[15]), .QN(n161) );
  DFF_X1 \f1_reg[12]  ( .D(n1017), .CK(clk), .Q(f1[12]), .QN(n20) );
  DFF_X1 \f1_reg[13]  ( .D(n1018), .CK(clk), .Q(f1[13]), .QN(n19) );
  DFF_X1 \f6_reg[14]  ( .D(n939), .CK(clk), .Q(f6[14]), .QN(n98) );
  DFF_X1 \f4_reg[14]  ( .D(n971), .CK(clk), .Q(f4[14]), .QN(n66) );
  BUF_X2 U3 ( .A(n1077), .Z(n11) );
  BUF_X1 U4 ( .A(data_out_x[2]), .Z(n1077) );
  BUF_X1 U5 ( .A(data_out_x[3]), .Z(n6) );
  BUF_X1 U6 ( .A(data_out_x[1]), .Z(n1075) );
  BUF_X2 U7 ( .A(data_out_x[1]), .Z(n1076) );
  BUF_X2 U8 ( .A(data_out_x[1]), .Z(n1021) );
  BUF_X2 U9 ( .A(data_out_x[1]), .Z(n284) );
  BUF_X2 U10 ( .A(data_out_x[1]), .Z(n283) );
  BUF_X2 U11 ( .A(data_out_x[3]), .Z(n2) );
  BUF_X8 U12 ( .A(data_out_x[6]), .Z(n1085) );
  CLKBUF_X2 U13 ( .A(data_out_x[0]), .Z(n1074) );
  OR2_X1 U14 ( .A1(n1065), .A2(n146), .ZN(n1) );
  NAND2_X1 U15 ( .A1(n1), .A2(n619), .ZN(n891) );
  CLKBUF_X2 U16 ( .A(data_out_x[3]), .Z(n7) );
  CLKBUF_X2 U17 ( .A(data_out_x[3]), .Z(n1079) );
  CLKBUF_X2 U18 ( .A(data_out_x[3]), .Z(n1080) );
  BUF_X2 U19 ( .A(n1077), .Z(n10) );
  BUF_X4 U20 ( .A(data_out_x[5]), .Z(n1083) );
  BUF_X2 U21 ( .A(data_out_x[0]), .Z(n1073) );
  CLKBUF_X3 U22 ( .A(data_out_x[3]), .Z(n3) );
  BUF_X4 U23 ( .A(data_out_x[4]), .Z(n4) );
  BUF_X4 U24 ( .A(data_out_x[5]), .Z(n1082) );
  BUF_X4 U25 ( .A(data_out_x[6]), .Z(n1084) );
  BUF_X4 U26 ( .A(data_out_x[4]), .Z(n1081) );
  CLKBUF_X3 U27 ( .A(data_out_x[2]), .Z(n1078) );
  CLKBUF_X3 U28 ( .A(n1077), .Z(n13) );
  CLKBUF_X3 U29 ( .A(n1077), .Z(n14) );
  BUF_X4 U30 ( .A(data_out_x[4]), .Z(n5) );
  CLKBUF_X3 U31 ( .A(data_out_x[1]), .Z(n1022) );
  OR2_X1 U32 ( .A1(n1070), .A2(n50), .ZN(n8) );
  NAND2_X1 U33 ( .A1(n8), .A2(n715), .ZN(n987) );
  CLKBUF_X1 U34 ( .A(data_out_x[0]), .Z(n9) );
  OR2_X1 U35 ( .A1(n1064), .A2(n161), .ZN(n12) );
  NAND2_X1 U36 ( .A1(n604), .A2(n12), .ZN(n876) );
  OR2_X1 U37 ( .A1(n1057), .A2(n241), .ZN(n15) );
  NAND2_X1 U38 ( .A1(n524), .A2(n15), .ZN(n796) );
  OR2_X1 U39 ( .A1(n1066), .A2(n129), .ZN(n16) );
  NAND2_X1 U40 ( .A1(n636), .A2(n16), .ZN(n908) );
  OR2_X1 U41 ( .A1(n1067), .A2(n113), .ZN(n273) );
  NAND2_X1 U42 ( .A1(n652), .A2(n273), .ZN(n924) );
  OR2_X1 U43 ( .A1(n1069), .A2(n65), .ZN(n274) );
  NAND2_X1 U44 ( .A1(n700), .A2(n274), .ZN(n972) );
  OR2_X1 U45 ( .A1(n1071), .A2(n33), .ZN(n275) );
  NAND2_X1 U46 ( .A1(n732), .A2(n275), .ZN(n1004) );
  OR2_X1 U47 ( .A1(n1062), .A2(n177), .ZN(n276) );
  NAND2_X1 U48 ( .A1(n588), .A2(n276), .ZN(n860) );
  OR2_X1 U49 ( .A1(n1070), .A2(n97), .ZN(n277) );
  NAND2_X1 U50 ( .A1(n668), .A2(n277), .ZN(n940) );
  OR2_X1 U51 ( .A1(n1070), .A2(n49), .ZN(n278) );
  NAND2_X1 U52 ( .A1(n716), .A2(n278), .ZN(n988) );
  OR2_X1 U53 ( .A1(n1058), .A2(n225), .ZN(n279) );
  NAND2_X1 U54 ( .A1(n540), .A2(n279), .ZN(n812) );
  OR2_X1 U55 ( .A1(n1070), .A2(n81), .ZN(n280) );
  NAND2_X1 U56 ( .A1(n684), .A2(n280), .ZN(n956) );
  OR2_X1 U57 ( .A1(n1060), .A2(n209), .ZN(n281) );
  NAND2_X1 U58 ( .A1(n556), .A2(n281), .ZN(n828) );
  OR2_X1 U59 ( .A1(n1061), .A2(n193), .ZN(n282) );
  NAND2_X1 U60 ( .A1(n572), .A2(n282), .ZN(n844) );
  BUF_X4 U61 ( .A(data_out_x[7]), .Z(n1086) );
  BUF_X1 U62 ( .A(n1026), .Z(n1045) );
  BUF_X1 U63 ( .A(n1025), .Z(n1041) );
  BUF_X1 U64 ( .A(n1025), .Z(n1037) );
  BUF_X1 U65 ( .A(n1024), .Z(n1033) );
  BUF_X1 U66 ( .A(n1027), .Z(n1049) );
  BUF_X1 U67 ( .A(n1026), .Z(n1047) );
  BUF_X1 U68 ( .A(n1026), .Z(n1046) );
  BUF_X1 U69 ( .A(n1026), .Z(n1044) );
  BUF_X1 U70 ( .A(n1026), .Z(n1043) );
  BUF_X1 U71 ( .A(n1026), .Z(n1042) );
  BUF_X1 U72 ( .A(n1025), .Z(n1040) );
  BUF_X1 U73 ( .A(n1025), .Z(n1039) );
  BUF_X1 U74 ( .A(n1025), .Z(n1038) );
  BUF_X1 U75 ( .A(n1025), .Z(n1036) );
  BUF_X1 U76 ( .A(n1024), .Z(n1035) );
  BUF_X1 U77 ( .A(n1024), .Z(n1034) );
  BUF_X1 U78 ( .A(n1024), .Z(n1032) );
  BUF_X1 U79 ( .A(n1024), .Z(n1031) );
  BUF_X1 U80 ( .A(n1024), .Z(n1030) );
  BUF_X1 U81 ( .A(n1027), .Z(n1050) );
  BUF_X1 U82 ( .A(n1027), .Z(n1048) );
  BUF_X1 U83 ( .A(n1054), .Z(n1068) );
  BUF_X1 U84 ( .A(n1052), .Z(n1055) );
  BUF_X1 U85 ( .A(n1052), .Z(n1059) );
  BUF_X1 U86 ( .A(n1053), .Z(n1063) );
  BUF_X1 U87 ( .A(n491), .Z(n1072) );
  BUF_X1 U88 ( .A(n1054), .Z(n1067) );
  BUF_X1 U89 ( .A(n1054), .Z(n1069) );
  BUF_X1 U90 ( .A(n1052), .Z(n1057) );
  BUF_X1 U91 ( .A(n1052), .Z(n1058) );
  BUF_X1 U92 ( .A(n1052), .Z(n1060) );
  BUF_X1 U93 ( .A(n1053), .Z(n1061) );
  BUF_X1 U94 ( .A(n1053), .Z(n1062) );
  BUF_X1 U95 ( .A(n1053), .Z(n1064) );
  BUF_X1 U96 ( .A(n1053), .Z(n1066) );
  BUF_X1 U97 ( .A(n491), .Z(n1070) );
  BUF_X1 U98 ( .A(n491), .Z(n1071) );
  BUF_X1 U99 ( .A(n1028), .Z(n1026) );
  BUF_X1 U100 ( .A(n1029), .Z(n1025) );
  BUF_X1 U101 ( .A(n1029), .Z(n1024) );
  BUF_X1 U102 ( .A(n1028), .Z(n1027) );
  INV_X1 U103 ( .A(n488), .ZN(n1094) );
  INV_X1 U104 ( .A(n475), .ZN(n1096) );
  INV_X1 U105 ( .A(n487), .ZN(n1093) );
  INV_X1 U106 ( .A(n474), .ZN(n1090) );
  BUF_X1 U107 ( .A(n491), .Z(n1054) );
  BUF_X1 U108 ( .A(n491), .Z(n1052) );
  BUF_X1 U109 ( .A(n491), .Z(n1053) );
  NAND4_X1 U110 ( .A1(n488), .A2(n487), .A3(n310), .A4(n489), .ZN(n311) );
  NOR4_X1 U111 ( .A1(n309), .A2(n308), .A3(n1095), .A4(n1092), .ZN(n489) );
  INV_X1 U112 ( .A(n305), .ZN(n1092) );
  INV_X1 U113 ( .A(n306), .ZN(n1095) );
  NAND4_X1 U114 ( .A1(n475), .A2(n474), .A3(n299), .A4(n476), .ZN(n301) );
  NOR4_X1 U115 ( .A1(n298), .A2(n297), .A3(n1097), .A4(n1091), .ZN(n476) );
  INV_X1 U116 ( .A(n295), .ZN(n1097) );
  INV_X1 U117 ( .A(n294), .ZN(n1091) );
  BUF_X1 U118 ( .A(n493), .Z(n1028) );
  BUF_X1 U119 ( .A(n493), .Z(n1029) );
  NAND2_X1 U120 ( .A1(n490), .A2(n477), .ZN(n306) );
  NAND2_X1 U121 ( .A1(n490), .A2(n482), .ZN(n310) );
  NAND2_X1 U122 ( .A1(n482), .A2(n479), .ZN(n299) );
  NAND2_X1 U123 ( .A1(n481), .A2(n1088), .ZN(n305) );
  NAND2_X1 U124 ( .A1(n477), .A2(n478), .ZN(n294) );
  AND2_X1 U125 ( .A1(n477), .A2(n1088), .ZN(n308) );
  AND2_X1 U126 ( .A1(n480), .A2(n478), .ZN(n297) );
  AND2_X1 U127 ( .A1(n490), .A2(n481), .ZN(n309) );
  AND2_X1 U128 ( .A1(n481), .A2(n479), .ZN(n298) );
  NAND2_X1 U129 ( .A1(n477), .A2(n479), .ZN(n295) );
  NOR2_X1 U130 ( .A1(n1088), .A2(n1098), .ZN(n478) );
  NAND2_X1 U131 ( .A1(n490), .A2(n480), .ZN(n488) );
  NAND2_X1 U132 ( .A1(n480), .A2(n1088), .ZN(n487) );
  NAND2_X1 U133 ( .A1(n478), .A2(n482), .ZN(n474) );
  NAND2_X1 U134 ( .A1(n480), .A2(n479), .ZN(n475) );
  INV_X1 U135 ( .A(n287), .ZN(n1099) );
  AND2_X1 U136 ( .A1(n491), .A2(n1100), .ZN(n493) );
  NOR2_X2 U137 ( .A1(n1101), .A2(clear_acc), .ZN(n293) );
  NOR2_X1 U138 ( .A1(n1098), .A2(addr_y[0]), .ZN(n479) );
  NOR2_X1 U139 ( .A1(n1088), .A2(addr_y[3]), .ZN(n490) );
  NOR2_X1 U140 ( .A1(addr_y[2]), .A2(addr_y[1]), .ZN(n482) );
  OAI221_X1 U141 ( .B1(n310), .B2(n64), .C1(n311), .C2(n48), .A(n486), .ZN(
        n483) );
  AOI22_X1 U142 ( .A1(f5[0]), .A2(n1094), .B1(f4[0]), .B2(n1093), .ZN(n486) );
  OAI221_X1 U143 ( .B1(n310), .B2(n63), .C1(n311), .C2(n47), .A(n466), .ZN(
        n463) );
  AOI22_X1 U144 ( .A1(f5[1]), .A2(n1094), .B1(f4[1]), .B2(n1093), .ZN(n466) );
  OAI221_X1 U145 ( .B1(n310), .B2(n62), .C1(n311), .C2(n46), .A(n455), .ZN(
        n452) );
  AOI22_X1 U146 ( .A1(f5[2]), .A2(n1094), .B1(f4[2]), .B2(n1093), .ZN(n455) );
  OAI221_X1 U147 ( .B1(n310), .B2(n61), .C1(n311), .C2(n45), .A(n444), .ZN(
        n441) );
  AOI22_X1 U148 ( .A1(f5[3]), .A2(n1094), .B1(f4[3]), .B2(n1093), .ZN(n444) );
  OAI221_X1 U149 ( .B1(n310), .B2(n60), .C1(n311), .C2(n44), .A(n433), .ZN(
        n430) );
  AOI22_X1 U150 ( .A1(f5[4]), .A2(n1094), .B1(f4[4]), .B2(n1093), .ZN(n433) );
  OAI221_X1 U151 ( .B1(n310), .B2(n59), .C1(n311), .C2(n43), .A(n422), .ZN(
        n419) );
  AOI22_X1 U152 ( .A1(f5[5]), .A2(n1094), .B1(f4[5]), .B2(n1093), .ZN(n422) );
  OAI221_X1 U153 ( .B1(n310), .B2(n58), .C1(n311), .C2(n42), .A(n411), .ZN(
        n408) );
  AOI22_X1 U154 ( .A1(f5[6]), .A2(n1094), .B1(f4[6]), .B2(n1093), .ZN(n411) );
  OAI221_X1 U155 ( .B1(n310), .B2(n57), .C1(n311), .C2(n41), .A(n400), .ZN(
        n397) );
  AOI22_X1 U156 ( .A1(f5[7]), .A2(n1094), .B1(f4[7]), .B2(n1093), .ZN(n400) );
  OAI221_X1 U157 ( .B1(n310), .B2(n56), .C1(n311), .C2(n40), .A(n389), .ZN(
        n386) );
  AOI22_X1 U158 ( .A1(f5[8]), .A2(n1094), .B1(f4[8]), .B2(n1093), .ZN(n389) );
  OAI221_X1 U159 ( .B1(n310), .B2(n55), .C1(n311), .C2(n39), .A(n378), .ZN(
        n375) );
  AOI22_X1 U160 ( .A1(f5[9]), .A2(n1094), .B1(f4[9]), .B2(n1093), .ZN(n378) );
  OAI221_X1 U161 ( .B1(n310), .B2(n54), .C1(n311), .C2(n38), .A(n367), .ZN(
        n364) );
  AOI22_X1 U162 ( .A1(f5[10]), .A2(n1094), .B1(f4[10]), .B2(n1093), .ZN(n367)
         );
  OAI221_X1 U163 ( .B1(n310), .B2(n53), .C1(n311), .C2(n37), .A(n356), .ZN(
        n353) );
  AOI22_X1 U164 ( .A1(f5[11]), .A2(n1094), .B1(f4[11]), .B2(n1093), .ZN(n356)
         );
  OAI221_X1 U165 ( .B1(n310), .B2(n52), .C1(n311), .C2(n36), .A(n345), .ZN(
        n342) );
  AOI22_X1 U166 ( .A1(f5[12]), .A2(n1094), .B1(f4[12]), .B2(n1093), .ZN(n345)
         );
  OAI221_X1 U167 ( .B1(n310), .B2(n51), .C1(n311), .C2(n35), .A(n334), .ZN(
        n331) );
  AOI22_X1 U168 ( .A1(f5[13]), .A2(n1094), .B1(f4[13]), .B2(n1093), .ZN(n334)
         );
  OAI221_X1 U169 ( .B1(n310), .B2(n50), .C1(n311), .C2(n34), .A(n323), .ZN(
        n320) );
  AOI22_X1 U170 ( .A1(f5[14]), .A2(n1094), .B1(f4[14]), .B2(n1093), .ZN(n323)
         );
  OAI221_X1 U171 ( .B1(n310), .B2(n49), .C1(n311), .C2(n33), .A(n312), .ZN(
        n303) );
  AOI22_X1 U172 ( .A1(f5[15]), .A2(n1094), .B1(f4[15]), .B2(n1093), .ZN(n312)
         );
  NAND3_X1 U173 ( .A1(n1101), .A2(n1100), .A3(clc), .ZN(n287) );
  OAI221_X1 U174 ( .B1(n299), .B2(n176), .C1(n472), .C2(n301), .A(n473), .ZN(
        n469) );
  AOI22_X1 U175 ( .A1(f12[0]), .A2(n1096), .B1(f11[0]), .B2(n1090), .ZN(n473)
         );
  NOR2_X1 U176 ( .A1(n483), .A2(n484), .ZN(n472) );
  OAI221_X1 U177 ( .B1(n305), .B2(n144), .C1(n306), .C2(n128), .A(n485), .ZN(
        n484) );
  OAI221_X1 U178 ( .B1(n299), .B2(n175), .C1(n461), .C2(n301), .A(n462), .ZN(
        n458) );
  AOI22_X1 U179 ( .A1(f12[1]), .A2(n1096), .B1(f11[1]), .B2(n1090), .ZN(n462)
         );
  NOR2_X1 U180 ( .A1(n463), .A2(n464), .ZN(n461) );
  OAI221_X1 U181 ( .B1(n305), .B2(n143), .C1(n306), .C2(n127), .A(n465), .ZN(
        n464) );
  OAI221_X1 U182 ( .B1(n299), .B2(n174), .C1(n450), .C2(n301), .A(n451), .ZN(
        n447) );
  AOI22_X1 U183 ( .A1(f12[2]), .A2(n1096), .B1(f11[2]), .B2(n1090), .ZN(n451)
         );
  NOR2_X1 U184 ( .A1(n452), .A2(n453), .ZN(n450) );
  OAI221_X1 U186 ( .B1(n305), .B2(n142), .C1(n306), .C2(n126), .A(n454), .ZN(
        n453) );
  OAI221_X1 U187 ( .B1(n299), .B2(n173), .C1(n439), .C2(n301), .A(n440), .ZN(
        n436) );
  AOI22_X1 U188 ( .A1(f12[3]), .A2(n1096), .B1(f11[3]), .B2(n1090), .ZN(n440)
         );
  NOR2_X1 U189 ( .A1(n441), .A2(n442), .ZN(n439) );
  OAI221_X1 U190 ( .B1(n305), .B2(n141), .C1(n306), .C2(n125), .A(n443), .ZN(
        n442) );
  OAI221_X1 U191 ( .B1(n299), .B2(n172), .C1(n428), .C2(n301), .A(n429), .ZN(
        n425) );
  AOI22_X1 U192 ( .A1(f12[4]), .A2(n1096), .B1(f11[4]), .B2(n1090), .ZN(n429)
         );
  NOR2_X1 U193 ( .A1(n430), .A2(n431), .ZN(n428) );
  OAI221_X1 U194 ( .B1(n305), .B2(n140), .C1(n306), .C2(n124), .A(n432), .ZN(
        n431) );
  OAI221_X1 U195 ( .B1(n299), .B2(n171), .C1(n417), .C2(n301), .A(n418), .ZN(
        n414) );
  AOI22_X1 U196 ( .A1(f12[5]), .A2(n1096), .B1(f11[5]), .B2(n1090), .ZN(n418)
         );
  NOR2_X1 U197 ( .A1(n419), .A2(n420), .ZN(n417) );
  OAI221_X1 U198 ( .B1(n305), .B2(n139), .C1(n306), .C2(n123), .A(n421), .ZN(
        n420) );
  OAI221_X1 U199 ( .B1(n299), .B2(n170), .C1(n406), .C2(n301), .A(n407), .ZN(
        n403) );
  AOI22_X1 U200 ( .A1(f12[6]), .A2(n1096), .B1(f11[6]), .B2(n1090), .ZN(n407)
         );
  NOR2_X1 U201 ( .A1(n408), .A2(n409), .ZN(n406) );
  OAI221_X1 U202 ( .B1(n305), .B2(n138), .C1(n306), .C2(n122), .A(n410), .ZN(
        n409) );
  OAI221_X1 U203 ( .B1(n299), .B2(n169), .C1(n395), .C2(n301), .A(n396), .ZN(
        n392) );
  AOI22_X1 U204 ( .A1(f12[7]), .A2(n1096), .B1(f11[7]), .B2(n1090), .ZN(n396)
         );
  NOR2_X1 U205 ( .A1(n397), .A2(n398), .ZN(n395) );
  OAI221_X1 U206 ( .B1(n305), .B2(n137), .C1(n306), .C2(n121), .A(n399), .ZN(
        n398) );
  OAI221_X1 U207 ( .B1(n299), .B2(n168), .C1(n384), .C2(n301), .A(n385), .ZN(
        n381) );
  AOI22_X1 U208 ( .A1(f12[8]), .A2(n1096), .B1(f11[8]), .B2(n1090), .ZN(n385)
         );
  NOR2_X1 U209 ( .A1(n386), .A2(n387), .ZN(n384) );
  OAI221_X1 U210 ( .B1(n305), .B2(n136), .C1(n306), .C2(n120), .A(n388), .ZN(
        n387) );
  OAI221_X1 U211 ( .B1(n299), .B2(n167), .C1(n373), .C2(n301), .A(n374), .ZN(
        n370) );
  AOI22_X1 U212 ( .A1(f12[9]), .A2(n1096), .B1(f11[9]), .B2(n1090), .ZN(n374)
         );
  NOR2_X1 U213 ( .A1(n375), .A2(n376), .ZN(n373) );
  OAI221_X1 U214 ( .B1(n305), .B2(n135), .C1(n306), .C2(n119), .A(n377), .ZN(
        n376) );
  OAI221_X1 U215 ( .B1(n299), .B2(n166), .C1(n362), .C2(n301), .A(n363), .ZN(
        n359) );
  AOI22_X1 U216 ( .A1(f12[10]), .A2(n1096), .B1(f11[10]), .B2(n1090), .ZN(n363) );
  NOR2_X1 U217 ( .A1(n364), .A2(n365), .ZN(n362) );
  OAI221_X1 U218 ( .B1(n305), .B2(n134), .C1(n306), .C2(n118), .A(n366), .ZN(
        n365) );
  OAI221_X1 U219 ( .B1(n299), .B2(n165), .C1(n351), .C2(n301), .A(n352), .ZN(
        n348) );
  AOI22_X1 U220 ( .A1(f12[11]), .A2(n1096), .B1(f11[11]), .B2(n1090), .ZN(n352) );
  NOR2_X1 U221 ( .A1(n353), .A2(n354), .ZN(n351) );
  OAI221_X1 U222 ( .B1(n305), .B2(n133), .C1(n306), .C2(n117), .A(n355), .ZN(
        n354) );
  OAI221_X1 U223 ( .B1(n299), .B2(n164), .C1(n340), .C2(n301), .A(n341), .ZN(
        n337) );
  AOI22_X1 U224 ( .A1(f12[12]), .A2(n1096), .B1(f11[12]), .B2(n1090), .ZN(n341) );
  NOR2_X1 U225 ( .A1(n342), .A2(n343), .ZN(n340) );
  OAI221_X1 U226 ( .B1(n305), .B2(n132), .C1(n306), .C2(n116), .A(n344), .ZN(
        n343) );
  OAI221_X1 U227 ( .B1(n299), .B2(n163), .C1(n329), .C2(n301), .A(n330), .ZN(
        n326) );
  AOI22_X1 U228 ( .A1(f12[13]), .A2(n1096), .B1(f11[13]), .B2(n1090), .ZN(n330) );
  NOR2_X1 U229 ( .A1(n331), .A2(n332), .ZN(n329) );
  OAI221_X1 U230 ( .B1(n305), .B2(n131), .C1(n306), .C2(n115), .A(n333), .ZN(
        n332) );
  OAI221_X1 U231 ( .B1(n299), .B2(n162), .C1(n318), .C2(n301), .A(n319), .ZN(
        n315) );
  AOI22_X1 U232 ( .A1(f12[14]), .A2(n1096), .B1(f11[14]), .B2(n1090), .ZN(n319) );
  NOR2_X1 U233 ( .A1(n320), .A2(n321), .ZN(n318) );
  OAI221_X1 U234 ( .B1(n305), .B2(n130), .C1(n306), .C2(n114), .A(n322), .ZN(
        n321) );
  OAI221_X1 U235 ( .B1(n299), .B2(n161), .C1(n300), .C2(n301), .A(n302), .ZN(
        n291) );
  AOI22_X1 U236 ( .A1(f12[15]), .A2(n1096), .B1(f11[15]), .B2(n1090), .ZN(n302) );
  NOR2_X1 U237 ( .A1(n303), .A2(n304), .ZN(n300) );
  OAI221_X1 U238 ( .B1(n305), .B2(n129), .C1(n306), .C2(n113), .A(n307), .ZN(
        n304) );
  NOR2_X1 U239 ( .A1(n1089), .A2(addr_y[2]), .ZN(n480) );
  BUF_X2 U240 ( .A(data_out_x[7]), .Z(n1087) );
  INV_X1 U241 ( .A(addr_y[3]), .ZN(n1098) );
  AND2_X1 U242 ( .A1(addr_y[2]), .A2(n1089), .ZN(n477) );
  AOI22_X1 U243 ( .A1(f6[0]), .A2(n308), .B1(f9[0]), .B2(n309), .ZN(n485) );
  AOI22_X1 U244 ( .A1(f6[1]), .A2(n308), .B1(f9[1]), .B2(n309), .ZN(n465) );
  AOI22_X1 U245 ( .A1(f6[2]), .A2(n308), .B1(f9[2]), .B2(n309), .ZN(n454) );
  AOI22_X1 U246 ( .A1(f6[3]), .A2(n308), .B1(f9[3]), .B2(n309), .ZN(n443) );
  AOI22_X1 U247 ( .A1(f6[4]), .A2(n308), .B1(f9[4]), .B2(n309), .ZN(n432) );
  AOI22_X1 U248 ( .A1(f6[5]), .A2(n308), .B1(f9[5]), .B2(n309), .ZN(n421) );
  AOI22_X1 U249 ( .A1(f6[6]), .A2(n308), .B1(f9[6]), .B2(n309), .ZN(n410) );
  AOI22_X1 U250 ( .A1(f6[7]), .A2(n308), .B1(f9[7]), .B2(n309), .ZN(n399) );
  AOI22_X1 U251 ( .A1(f6[8]), .A2(n308), .B1(f9[8]), .B2(n309), .ZN(n388) );
  AOI22_X1 U252 ( .A1(f6[9]), .A2(n308), .B1(f9[9]), .B2(n309), .ZN(n377) );
  AOI22_X1 U253 ( .A1(f6[10]), .A2(n308), .B1(f9[10]), .B2(n309), .ZN(n366) );
  AOI22_X1 U254 ( .A1(f6[11]), .A2(n308), .B1(f9[11]), .B2(n309), .ZN(n355) );
  AOI22_X1 U255 ( .A1(f6[12]), .A2(n308), .B1(f9[12]), .B2(n309), .ZN(n344) );
  AOI22_X1 U256 ( .A1(f6[13]), .A2(n308), .B1(f9[13]), .B2(n309), .ZN(n333) );
  AOI22_X1 U257 ( .A1(f6[14]), .A2(n308), .B1(f9[14]), .B2(n309), .ZN(n322) );
  AOI22_X1 U258 ( .A1(f6[15]), .A2(n308), .B1(f9[15]), .B2(n309), .ZN(n307) );
  AOI22_X1 U259 ( .A1(f13[0]), .A2(n297), .B1(f16[0]), .B2(n298), .ZN(n471) );
  AOI22_X1 U260 ( .A1(f13[1]), .A2(n297), .B1(f16[1]), .B2(n298), .ZN(n460) );
  AOI22_X1 U261 ( .A1(f13[2]), .A2(n297), .B1(f16[2]), .B2(n298), .ZN(n449) );
  AOI22_X1 U262 ( .A1(f13[3]), .A2(n297), .B1(f16[3]), .B2(n298), .ZN(n438) );
  AOI22_X1 U263 ( .A1(f13[4]), .A2(n297), .B1(f16[4]), .B2(n298), .ZN(n427) );
  AOI22_X1 U264 ( .A1(f13[5]), .A2(n297), .B1(f16[5]), .B2(n298), .ZN(n416) );
  AOI22_X1 U265 ( .A1(f13[6]), .A2(n297), .B1(f16[6]), .B2(n298), .ZN(n405) );
  AOI22_X1 U266 ( .A1(f13[7]), .A2(n297), .B1(f16[7]), .B2(n298), .ZN(n394) );
  AOI22_X1 U267 ( .A1(f13[8]), .A2(n297), .B1(f16[8]), .B2(n298), .ZN(n383) );
  AOI22_X1 U268 ( .A1(f13[9]), .A2(n297), .B1(f16[9]), .B2(n298), .ZN(n372) );
  AOI22_X1 U269 ( .A1(f13[10]), .A2(n297), .B1(f16[10]), .B2(n298), .ZN(n361)
         );
  AOI22_X1 U270 ( .A1(f13[11]), .A2(n297), .B1(f16[11]), .B2(n298), .ZN(n350)
         );
  AOI22_X1 U271 ( .A1(f13[12]), .A2(n297), .B1(f16[12]), .B2(n298), .ZN(n339)
         );
  AOI22_X1 U272 ( .A1(f13[13]), .A2(n297), .B1(f16[13]), .B2(n298), .ZN(n328)
         );
  AOI22_X1 U273 ( .A1(f13[14]), .A2(n297), .B1(f16[14]), .B2(n298), .ZN(n317)
         );
  AOI22_X1 U274 ( .A1(f13[15]), .A2(n297), .B1(f16[15]), .B2(n298), .ZN(n296)
         );
  AOI21_X1 U275 ( .B1(n1100), .B2(clc1), .A(n1099), .ZN(n491) );
  OAI21_X1 U276 ( .B1(n1065), .B2(n151), .A(n614), .ZN(n886) );
  NAND2_X1 U277 ( .A1(add_r9[9]), .A2(n1041), .ZN(n614) );
  OAI21_X1 U278 ( .B1(n1065), .B2(n150), .A(n615), .ZN(n887) );
  NAND2_X1 U279 ( .A1(add_r9[10]), .A2(n1041), .ZN(n615) );
  OAI21_X1 U280 ( .B1(n1065), .B2(n149), .A(n616), .ZN(n888) );
  NAND2_X1 U281 ( .A1(add_r9[11]), .A2(n1041), .ZN(n616) );
  NAND2_X1 U282 ( .A1(add_r9[14]), .A2(n1040), .ZN(n619) );
  OAI21_X1 U283 ( .B1(n1056), .B2(n258), .A(n507), .ZN(n779) );
  NAND2_X1 U284 ( .A1(add_r16[14]), .A2(n1050), .ZN(n507) );
  OAI21_X1 U285 ( .B1(n1065), .B2(n147), .A(n618), .ZN(n890) );
  NAND2_X1 U286 ( .A1(add_r9[13]), .A2(n1040), .ZN(n618) );
  OAI21_X1 U287 ( .B1(n1056), .B2(n259), .A(n506), .ZN(n778) );
  NAND2_X1 U288 ( .A1(add_r16[13]), .A2(n1050), .ZN(n506) );
  OAI21_X1 U289 ( .B1(n1065), .B2(n148), .A(n617), .ZN(n889) );
  NAND2_X1 U290 ( .A1(add_r9[12]), .A2(n1040), .ZN(n617) );
  OAI21_X1 U291 ( .B1(n1056), .B2(n260), .A(n505), .ZN(n777) );
  NAND2_X1 U292 ( .A1(add_r16[12]), .A2(n1050), .ZN(n505) );
  OAI21_X1 U293 ( .B1(n1056), .B2(n256), .A(n509), .ZN(n781) );
  NAND2_X1 U294 ( .A1(add_r15[0]), .A2(n1049), .ZN(n509) );
  OAI21_X1 U295 ( .B1(n1056), .B2(n255), .A(n510), .ZN(n782) );
  NAND2_X1 U296 ( .A1(add_r15[1]), .A2(n1049), .ZN(n510) );
  OAI21_X1 U297 ( .B1(n1056), .B2(n254), .A(n511), .ZN(n783) );
  NAND2_X1 U298 ( .A1(add_r15[2]), .A2(n1049), .ZN(n511) );
  OAI21_X1 U299 ( .B1(n1056), .B2(n253), .A(n512), .ZN(n784) );
  NAND2_X1 U300 ( .A1(add_r15[3]), .A2(n1049), .ZN(n512) );
  OAI21_X1 U301 ( .B1(n1056), .B2(n252), .A(n513), .ZN(n785) );
  NAND2_X1 U302 ( .A1(add_r15[4]), .A2(n1049), .ZN(n513) );
  OAI21_X1 U303 ( .B1(n1056), .B2(n251), .A(n514), .ZN(n786) );
  NAND2_X1 U304 ( .A1(add_r15[5]), .A2(n1049), .ZN(n514) );
  OAI21_X1 U305 ( .B1(n1056), .B2(n250), .A(n515), .ZN(n787) );
  NAND2_X1 U306 ( .A1(add_r15[6]), .A2(n1049), .ZN(n515) );
  OAI21_X1 U307 ( .B1(n1056), .B2(n249), .A(n516), .ZN(n788) );
  NAND2_X1 U308 ( .A1(add_r15[7]), .A2(n1049), .ZN(n516) );
  OAI21_X1 U309 ( .B1(n1065), .B2(n152), .A(n613), .ZN(n885) );
  NAND2_X1 U310 ( .A1(add_r9[8]), .A2(n1041), .ZN(n613) );
  OAI211_X1 U311 ( .C1(n287), .C2(n32), .A(n467), .B(n468), .ZN(n764) );
  NAND2_X1 U312 ( .A1(f[0]), .A2(n290), .ZN(n468) );
  OAI21_X1 U313 ( .B1(n469), .B2(n470), .A(n293), .ZN(n467) );
  OAI221_X1 U314 ( .B1(n294), .B2(n256), .C1(n295), .C2(n240), .A(n471), .ZN(
        n470) );
  OAI211_X1 U315 ( .C1(n287), .C2(n31), .A(n456), .B(n457), .ZN(n763) );
  NAND2_X1 U316 ( .A1(f[1]), .A2(n290), .ZN(n457) );
  OAI21_X1 U317 ( .B1(n458), .B2(n459), .A(n293), .ZN(n456) );
  OAI221_X1 U318 ( .B1(n294), .B2(n255), .C1(n295), .C2(n239), .A(n460), .ZN(
        n459) );
  OAI211_X1 U319 ( .C1(n287), .C2(n30), .A(n445), .B(n446), .ZN(n762) );
  NAND2_X1 U320 ( .A1(f[2]), .A2(n290), .ZN(n446) );
  OAI21_X1 U321 ( .B1(n447), .B2(n448), .A(n293), .ZN(n445) );
  OAI221_X1 U322 ( .B1(n294), .B2(n254), .C1(n295), .C2(n238), .A(n449), .ZN(
        n448) );
  OAI211_X1 U323 ( .C1(n287), .C2(n29), .A(n434), .B(n435), .ZN(n761) );
  NAND2_X1 U324 ( .A1(f[3]), .A2(n290), .ZN(n435) );
  OAI21_X1 U325 ( .B1(n436), .B2(n437), .A(n293), .ZN(n434) );
  OAI221_X1 U326 ( .B1(n294), .B2(n253), .C1(n295), .C2(n237), .A(n438), .ZN(
        n437) );
  OAI211_X1 U327 ( .C1(n287), .C2(n28), .A(n423), .B(n424), .ZN(n760) );
  NAND2_X1 U328 ( .A1(f[4]), .A2(n290), .ZN(n424) );
  OAI21_X1 U329 ( .B1(n425), .B2(n426), .A(n293), .ZN(n423) );
  OAI221_X1 U330 ( .B1(n294), .B2(n252), .C1(n295), .C2(n236), .A(n427), .ZN(
        n426) );
  OAI211_X1 U331 ( .C1(n287), .C2(n27), .A(n412), .B(n413), .ZN(n759) );
  NAND2_X1 U332 ( .A1(f[5]), .A2(n290), .ZN(n413) );
  OAI21_X1 U333 ( .B1(n414), .B2(n415), .A(n293), .ZN(n412) );
  OAI221_X1 U334 ( .B1(n294), .B2(n251), .C1(n295), .C2(n235), .A(n416), .ZN(
        n415) );
  OAI211_X1 U335 ( .C1(n287), .C2(n26), .A(n401), .B(n402), .ZN(n758) );
  NAND2_X1 U336 ( .A1(f[6]), .A2(n290), .ZN(n402) );
  OAI21_X1 U337 ( .B1(n403), .B2(n404), .A(n293), .ZN(n401) );
  OAI221_X1 U338 ( .B1(n294), .B2(n250), .C1(n295), .C2(n234), .A(n405), .ZN(
        n404) );
  OAI211_X1 U339 ( .C1(n287), .C2(n25), .A(n390), .B(n391), .ZN(n757) );
  NAND2_X1 U340 ( .A1(f[7]), .A2(n290), .ZN(n391) );
  OAI21_X1 U341 ( .B1(n392), .B2(n393), .A(n293), .ZN(n390) );
  OAI221_X1 U342 ( .B1(n294), .B2(n249), .C1(n295), .C2(n233), .A(n394), .ZN(
        n393) );
  OAI211_X1 U343 ( .C1(n287), .C2(n24), .A(n379), .B(n380), .ZN(n756) );
  NAND2_X1 U344 ( .A1(f[8]), .A2(n290), .ZN(n380) );
  OAI21_X1 U345 ( .B1(n381), .B2(n382), .A(n293), .ZN(n379) );
  OAI221_X1 U346 ( .B1(n294), .B2(n248), .C1(n295), .C2(n232), .A(n383), .ZN(
        n382) );
  OAI211_X1 U347 ( .C1(n287), .C2(n23), .A(n368), .B(n369), .ZN(n755) );
  NAND2_X1 U348 ( .A1(f[9]), .A2(n290), .ZN(n369) );
  OAI21_X1 U349 ( .B1(n370), .B2(n371), .A(n293), .ZN(n368) );
  OAI221_X1 U350 ( .B1(n294), .B2(n247), .C1(n295), .C2(n231), .A(n372), .ZN(
        n371) );
  OAI211_X1 U351 ( .C1(n287), .C2(n22), .A(n357), .B(n358), .ZN(n754) );
  NAND2_X1 U352 ( .A1(f[10]), .A2(n290), .ZN(n358) );
  OAI21_X1 U353 ( .B1(n359), .B2(n360), .A(n293), .ZN(n357) );
  OAI221_X1 U354 ( .B1(n294), .B2(n246), .C1(n295), .C2(n230), .A(n361), .ZN(
        n360) );
  OAI211_X1 U355 ( .C1(n287), .C2(n21), .A(n346), .B(n347), .ZN(n753) );
  NAND2_X1 U356 ( .A1(f[11]), .A2(n290), .ZN(n347) );
  OAI21_X1 U357 ( .B1(n348), .B2(n349), .A(n293), .ZN(n346) );
  OAI221_X1 U358 ( .B1(n294), .B2(n245), .C1(n295), .C2(n229), .A(n350), .ZN(
        n349) );
  OAI211_X1 U359 ( .C1(n287), .C2(n20), .A(n335), .B(n336), .ZN(n752) );
  NAND2_X1 U360 ( .A1(f[12]), .A2(n290), .ZN(n336) );
  OAI21_X1 U361 ( .B1(n337), .B2(n338), .A(n293), .ZN(n335) );
  OAI221_X1 U362 ( .B1(n294), .B2(n244), .C1(n295), .C2(n228), .A(n339), .ZN(
        n338) );
  OAI211_X1 U363 ( .C1(n287), .C2(n19), .A(n324), .B(n325), .ZN(n751) );
  NAND2_X1 U364 ( .A1(f[13]), .A2(n290), .ZN(n325) );
  OAI21_X1 U365 ( .B1(n326), .B2(n327), .A(n293), .ZN(n324) );
  OAI221_X1 U366 ( .B1(n294), .B2(n243), .C1(n295), .C2(n227), .A(n328), .ZN(
        n327) );
  OAI211_X1 U367 ( .C1(n287), .C2(n18), .A(n313), .B(n314), .ZN(n750) );
  NAND2_X1 U368 ( .A1(f[14]), .A2(n290), .ZN(n314) );
  OAI21_X1 U369 ( .B1(n315), .B2(n316), .A(n293), .ZN(n313) );
  OAI221_X1 U370 ( .B1(n294), .B2(n242), .C1(n295), .C2(n226), .A(n317), .ZN(
        n316) );
  OAI211_X1 U371 ( .C1(n287), .C2(n17), .A(n288), .B(n289), .ZN(n749) );
  NAND2_X1 U372 ( .A1(f[15]), .A2(n290), .ZN(n289) );
  OAI21_X1 U373 ( .B1(n291), .B2(n292), .A(n293), .ZN(n288) );
  OAI221_X1 U374 ( .B1(n294), .B2(n241), .C1(n295), .C2(n225), .A(n296), .ZN(
        n292) );
  AND2_X1 U375 ( .A1(addr_y[2]), .A2(addr_y[1]), .ZN(n481) );
  INV_X1 U376 ( .A(clc1), .ZN(n1101) );
  INV_X1 U377 ( .A(clear_acc), .ZN(n1100) );
  OAI21_X1 U378 ( .B1(n1055), .B2(n18), .A(n747), .ZN(n1019) );
  NAND2_X1 U379 ( .A1(add_r1[14]), .A2(n1030), .ZN(n747) );
  OAI21_X1 U380 ( .B1(n1059), .B2(n19), .A(n746), .ZN(n1018) );
  NAND2_X1 U381 ( .A1(add_r1[13]), .A2(n1030), .ZN(n746) );
  OAI21_X1 U382 ( .B1(n1072), .B2(n20), .A(n745), .ZN(n1017) );
  NAND2_X1 U383 ( .A1(add_r1[12]), .A2(n1030), .ZN(n745) );
  OAI21_X1 U384 ( .B1(n1072), .B2(n118), .A(n647), .ZN(n919) );
  NAND2_X1 U385 ( .A1(add_r7[10]), .A2(n1038), .ZN(n647) );
  OAI21_X1 U386 ( .B1(n1063), .B2(n117), .A(n648), .ZN(n920) );
  NAND2_X1 U387 ( .A1(add_r7[11]), .A2(n1038), .ZN(n648) );
  OAI21_X1 U388 ( .B1(n1068), .B2(n71), .A(n694), .ZN(n966) );
  NAND2_X1 U389 ( .A1(add_r4[9]), .A2(n1034), .ZN(n694) );
  OAI21_X1 U390 ( .B1(n1068), .B2(n70), .A(n695), .ZN(n967) );
  NAND2_X1 U391 ( .A1(add_r4[10]), .A2(n1034), .ZN(n695) );
  OAI21_X1 U392 ( .B1(n1068), .B2(n69), .A(n696), .ZN(n968) );
  NAND2_X1 U393 ( .A1(add_r4[11]), .A2(n1034), .ZN(n696) );
  OAI21_X1 U394 ( .B1(n1055), .B2(n124), .A(n641), .ZN(n913) );
  NAND2_X1 U395 ( .A1(add_r7[4]), .A2(n1038), .ZN(n641) );
  OAI21_X1 U396 ( .B1(n1059), .B2(n123), .A(n642), .ZN(n914) );
  NAND2_X1 U397 ( .A1(add_r7[5]), .A2(n1038), .ZN(n642) );
  OAI21_X1 U398 ( .B1(n1071), .B2(n122), .A(n643), .ZN(n915) );
  NAND2_X1 U399 ( .A1(add_r7[6]), .A2(n1038), .ZN(n643) );
  OAI21_X1 U400 ( .B1(n1068), .B2(n121), .A(n644), .ZN(n916) );
  NAND2_X1 U401 ( .A1(add_r7[7]), .A2(n1038), .ZN(n644) );
  OAI21_X1 U402 ( .B1(n1070), .B2(n120), .A(n645), .ZN(n917) );
  NAND2_X1 U403 ( .A1(add_r7[8]), .A2(n1038), .ZN(n645) );
  OAI21_X1 U404 ( .B1(n491), .B2(n119), .A(n646), .ZN(n918) );
  NAND2_X1 U405 ( .A1(add_r7[9]), .A2(n1038), .ZN(n646) );
  OAI21_X1 U406 ( .B1(n1068), .B2(n75), .A(n690), .ZN(n962) );
  NAND2_X1 U407 ( .A1(add_r4[5]), .A2(n1034), .ZN(n690) );
  OAI21_X1 U408 ( .B1(n1068), .B2(n74), .A(n691), .ZN(n963) );
  NAND2_X1 U409 ( .A1(add_r4[6]), .A2(n1034), .ZN(n691) );
  OAI21_X1 U410 ( .B1(n1068), .B2(n73), .A(n692), .ZN(n964) );
  NAND2_X1 U411 ( .A1(add_r4[7]), .A2(n1034), .ZN(n692) );
  OAI21_X1 U412 ( .B1(n1068), .B2(n72), .A(n693), .ZN(n965) );
  NAND2_X1 U413 ( .A1(add_r4[8]), .A2(n1034), .ZN(n693) );
  OAI21_X1 U414 ( .B1(n1055), .B2(n263), .A(n502), .ZN(n774) );
  NAND2_X1 U415 ( .A1(add_r16[9]), .A2(n1050), .ZN(n502) );
  OAI21_X1 U416 ( .B1(n1055), .B2(n262), .A(n503), .ZN(n775) );
  NAND2_X1 U417 ( .A1(add_r16[10]), .A2(n1050), .ZN(n503) );
  OAI21_X1 U418 ( .B1(n1055), .B2(n261), .A(n504), .ZN(n776) );
  NAND2_X1 U419 ( .A1(add_r16[11]), .A2(n1050), .ZN(n504) );
  OAI21_X1 U420 ( .B1(n1059), .B2(n214), .A(n551), .ZN(n823) );
  NAND2_X1 U421 ( .A1(add_r13[10]), .A2(n1046), .ZN(n551) );
  OAI21_X1 U422 ( .B1(n1059), .B2(n213), .A(n552), .ZN(n824) );
  NAND2_X1 U423 ( .A1(add_r13[11]), .A2(n1046), .ZN(n552) );
  OAI21_X1 U424 ( .B1(n1063), .B2(n167), .A(n598), .ZN(n870) );
  NAND2_X1 U425 ( .A1(add_r10[9]), .A2(n1042), .ZN(n598) );
  OAI21_X1 U426 ( .B1(n1063), .B2(n166), .A(n599), .ZN(n871) );
  NAND2_X1 U427 ( .A1(add_r10[10]), .A2(n1042), .ZN(n599) );
  OAI21_X1 U428 ( .B1(n1063), .B2(n165), .A(n600), .ZN(n872) );
  NAND2_X1 U429 ( .A1(add_r10[11]), .A2(n1042), .ZN(n600) );
  OAI21_X1 U430 ( .B1(n1055), .B2(n272), .A(n492), .ZN(n765) );
  NAND2_X1 U431 ( .A1(add_r16[0]), .A2(n1051), .ZN(n492) );
  OAI21_X1 U432 ( .B1(n1055), .B2(n271), .A(n494), .ZN(n766) );
  NAND2_X1 U433 ( .A1(add_r16[1]), .A2(n1051), .ZN(n494) );
  OAI21_X1 U434 ( .B1(n1055), .B2(n270), .A(n495), .ZN(n767) );
  NAND2_X1 U435 ( .A1(add_r16[2]), .A2(n1051), .ZN(n495) );
  OAI21_X1 U436 ( .B1(n1055), .B2(n269), .A(n496), .ZN(n768) );
  NAND2_X1 U437 ( .A1(add_r16[3]), .A2(n1051), .ZN(n496) );
  OAI21_X1 U438 ( .B1(n1055), .B2(n268), .A(n497), .ZN(n769) );
  NAND2_X1 U439 ( .A1(add_r16[4]), .A2(n1050), .ZN(n497) );
  OAI21_X1 U440 ( .B1(n1055), .B2(n266), .A(n499), .ZN(n771) );
  NAND2_X1 U441 ( .A1(add_r16[6]), .A2(n1050), .ZN(n499) );
  OAI21_X1 U442 ( .B1(n1055), .B2(n265), .A(n500), .ZN(n772) );
  NAND2_X1 U443 ( .A1(add_r16[7]), .A2(n1050), .ZN(n500) );
  OAI21_X1 U444 ( .B1(n1055), .B2(n264), .A(n501), .ZN(n773) );
  NAND2_X1 U445 ( .A1(add_r16[8]), .A2(n1050), .ZN(n501) );
  OAI21_X1 U446 ( .B1(n1059), .B2(n220), .A(n545), .ZN(n817) );
  NAND2_X1 U447 ( .A1(add_r13[4]), .A2(n1046), .ZN(n545) );
  OAI21_X1 U448 ( .B1(n1059), .B2(n219), .A(n546), .ZN(n818) );
  NAND2_X1 U449 ( .A1(add_r13[5]), .A2(n1046), .ZN(n546) );
  OAI21_X1 U450 ( .B1(n1059), .B2(n218), .A(n547), .ZN(n819) );
  NAND2_X1 U451 ( .A1(add_r13[6]), .A2(n1046), .ZN(n547) );
  OAI21_X1 U452 ( .B1(n1059), .B2(n217), .A(n548), .ZN(n820) );
  NAND2_X1 U453 ( .A1(add_r13[7]), .A2(n1046), .ZN(n548) );
  OAI21_X1 U454 ( .B1(n1059), .B2(n216), .A(n549), .ZN(n821) );
  NAND2_X1 U455 ( .A1(add_r13[8]), .A2(n1046), .ZN(n549) );
  OAI21_X1 U456 ( .B1(n1059), .B2(n215), .A(n550), .ZN(n822) );
  NAND2_X1 U457 ( .A1(add_r13[9]), .A2(n1046), .ZN(n550) );
  OAI21_X1 U458 ( .B1(n1063), .B2(n170), .A(n595), .ZN(n867) );
  NAND2_X1 U459 ( .A1(add_r10[6]), .A2(n1042), .ZN(n595) );
  OAI21_X1 U460 ( .B1(n1063), .B2(n169), .A(n596), .ZN(n868) );
  NAND2_X1 U461 ( .A1(add_r10[7]), .A2(n1042), .ZN(n596) );
  OAI21_X1 U462 ( .B1(n1063), .B2(n168), .A(n597), .ZN(n869) );
  NAND2_X1 U463 ( .A1(add_r10[8]), .A2(n1042), .ZN(n597) );
  OAI21_X1 U464 ( .B1(n1072), .B2(n23), .A(n742), .ZN(n1014) );
  NAND2_X1 U465 ( .A1(add_r1[9]), .A2(n1030), .ZN(n742) );
  OAI21_X1 U466 ( .B1(n1072), .B2(n22), .A(n743), .ZN(n1015) );
  NAND2_X1 U467 ( .A1(add_r1[10]), .A2(n1030), .ZN(n743) );
  OAI21_X1 U468 ( .B1(n1072), .B2(n21), .A(n744), .ZN(n1016) );
  NAND2_X1 U469 ( .A1(add_r1[11]), .A2(n1030), .ZN(n744) );
  OAI21_X1 U470 ( .B1(n1072), .B2(n28), .A(n737), .ZN(n1009) );
  NAND2_X1 U471 ( .A1(add_r1[4]), .A2(n1030), .ZN(n737) );
  OAI21_X1 U472 ( .B1(n1072), .B2(n27), .A(n738), .ZN(n1010) );
  NAND2_X1 U473 ( .A1(add_r1[5]), .A2(n1030), .ZN(n738) );
  OAI21_X1 U474 ( .B1(n1072), .B2(n26), .A(n739), .ZN(n1011) );
  NAND2_X1 U475 ( .A1(add_r1[6]), .A2(n1030), .ZN(n739) );
  OAI21_X1 U476 ( .B1(n1072), .B2(n25), .A(n740), .ZN(n1012) );
  NAND2_X1 U477 ( .A1(add_r1[7]), .A2(n1030), .ZN(n740) );
  OAI21_X1 U478 ( .B1(n1072), .B2(n24), .A(n741), .ZN(n1013) );
  NAND2_X1 U479 ( .A1(add_r1[8]), .A2(n1030), .ZN(n741) );
  OAI21_X1 U480 ( .B1(n1071), .B2(n103), .A(n662), .ZN(n934) );
  NAND2_X1 U481 ( .A1(add_r6[9]), .A2(n1037), .ZN(n662) );
  OAI21_X1 U482 ( .B1(n1072), .B2(n102), .A(n663), .ZN(n935) );
  NAND2_X1 U483 ( .A1(add_r6[10]), .A2(n1037), .ZN(n663) );
  OAI21_X1 U484 ( .B1(n1070), .B2(n101), .A(n664), .ZN(n936) );
  NAND2_X1 U485 ( .A1(add_r6[11]), .A2(n1037), .ZN(n664) );
  OAI21_X1 U486 ( .B1(n1072), .B2(n86), .A(n679), .ZN(n951) );
  NAND2_X1 U487 ( .A1(add_r5[10]), .A2(n1035), .ZN(n679) );
  OAI21_X1 U488 ( .B1(n1068), .B2(n85), .A(n680), .ZN(n952) );
  NAND2_X1 U489 ( .A1(add_r5[11]), .A2(n1035), .ZN(n680) );
  OAI21_X1 U490 ( .B1(n1071), .B2(n98), .A(n667), .ZN(n939) );
  NAND2_X1 U491 ( .A1(add_r6[14]), .A2(n1036), .ZN(n667) );
  OAI21_X1 U492 ( .B1(n1069), .B2(n66), .A(n699), .ZN(n971) );
  NAND2_X1 U493 ( .A1(add_r4[14]), .A2(n1034), .ZN(n699) );
  OAI21_X1 U494 ( .B1(n1068), .B2(n82), .A(n683), .ZN(n955) );
  NAND2_X1 U495 ( .A1(add_r5[14]), .A2(n1035), .ZN(n683) );
  OAI21_X1 U496 ( .B1(n1067), .B2(n114), .A(n651), .ZN(n923) );
  NAND2_X1 U497 ( .A1(add_r7[14]), .A2(n1038), .ZN(n651) );
  OAI21_X1 U498 ( .B1(n1072), .B2(n99), .A(n666), .ZN(n938) );
  NAND2_X1 U499 ( .A1(add_r6[13]), .A2(n1036), .ZN(n666) );
  OAI21_X1 U500 ( .B1(n1069), .B2(n67), .A(n698), .ZN(n970) );
  NAND2_X1 U501 ( .A1(add_r4[13]), .A2(n1034), .ZN(n698) );
  OAI21_X1 U502 ( .B1(n1072), .B2(n83), .A(n682), .ZN(n954) );
  NAND2_X1 U503 ( .A1(add_r5[13]), .A2(n1035), .ZN(n682) );
  OAI21_X1 U504 ( .B1(n1067), .B2(n115), .A(n650), .ZN(n922) );
  NAND2_X1 U505 ( .A1(add_r7[13]), .A2(n1038), .ZN(n650) );
  OAI21_X1 U506 ( .B1(n1070), .B2(n100), .A(n665), .ZN(n937) );
  NAND2_X1 U507 ( .A1(add_r6[12]), .A2(n1036), .ZN(n665) );
  OAI21_X1 U508 ( .B1(n1069), .B2(n68), .A(n697), .ZN(n969) );
  NAND2_X1 U509 ( .A1(add_r4[12]), .A2(n1034), .ZN(n697) );
  OAI21_X1 U510 ( .B1(n1063), .B2(n84), .A(n681), .ZN(n953) );
  NAND2_X1 U511 ( .A1(add_r5[12]), .A2(n1035), .ZN(n681) );
  OAI21_X1 U512 ( .B1(n1067), .B2(n116), .A(n649), .ZN(n921) );
  NAND2_X1 U513 ( .A1(add_r7[12]), .A2(n1038), .ZN(n649) );
  OAI21_X1 U514 ( .B1(n1067), .B2(n112), .A(n653), .ZN(n925) );
  NAND2_X1 U515 ( .A1(add_r6[0]), .A2(n1037), .ZN(n653) );
  OAI21_X1 U516 ( .B1(n1067), .B2(n111), .A(n654), .ZN(n926) );
  NAND2_X1 U517 ( .A1(add_r6[1]), .A2(n1037), .ZN(n654) );
  OAI21_X1 U518 ( .B1(n1067), .B2(n110), .A(n655), .ZN(n927) );
  NAND2_X1 U519 ( .A1(add_r6[2]), .A2(n1037), .ZN(n655) );
  OAI21_X1 U520 ( .B1(n1067), .B2(n109), .A(n656), .ZN(n928) );
  NAND2_X1 U521 ( .A1(add_r6[3]), .A2(n1037), .ZN(n656) );
  OAI21_X1 U522 ( .B1(n1067), .B2(n108), .A(n657), .ZN(n929) );
  NAND2_X1 U523 ( .A1(add_r6[4]), .A2(n1037), .ZN(n657) );
  OAI21_X1 U524 ( .B1(n1067), .B2(n107), .A(n658), .ZN(n930) );
  NAND2_X1 U525 ( .A1(add_r6[5]), .A2(n1037), .ZN(n658) );
  OAI21_X1 U526 ( .B1(n1067), .B2(n106), .A(n659), .ZN(n931) );
  NAND2_X1 U527 ( .A1(add_r6[6]), .A2(n1037), .ZN(n659) );
  OAI21_X1 U528 ( .B1(n1067), .B2(n105), .A(n660), .ZN(n932) );
  NAND2_X1 U529 ( .A1(add_r6[7]), .A2(n1037), .ZN(n660) );
  OAI21_X1 U530 ( .B1(n1071), .B2(n104), .A(n661), .ZN(n933) );
  NAND2_X1 U531 ( .A1(add_r6[8]), .A2(n1037), .ZN(n661) );
  OAI21_X1 U532 ( .B1(n1055), .B2(n92), .A(n673), .ZN(n945) );
  NAND2_X1 U533 ( .A1(add_r5[4]), .A2(n1036), .ZN(n673) );
  OAI21_X1 U534 ( .B1(n1059), .B2(n91), .A(n674), .ZN(n946) );
  NAND2_X1 U535 ( .A1(add_r5[5]), .A2(n1036), .ZN(n674) );
  OAI21_X1 U536 ( .B1(n1068), .B2(n90), .A(n675), .ZN(n947) );
  NAND2_X1 U537 ( .A1(add_r5[6]), .A2(n1036), .ZN(n675) );
  OAI21_X1 U538 ( .B1(n1070), .B2(n89), .A(n676), .ZN(n948) );
  NAND2_X1 U539 ( .A1(add_r5[7]), .A2(n1036), .ZN(n676) );
  OAI21_X1 U540 ( .B1(n1072), .B2(n88), .A(n677), .ZN(n949) );
  NAND2_X1 U541 ( .A1(add_r5[8]), .A2(n1035), .ZN(n677) );
  OAI21_X1 U542 ( .B1(n1063), .B2(n87), .A(n678), .ZN(n950) );
  NAND2_X1 U543 ( .A1(add_r5[9]), .A2(n1035), .ZN(n678) );
  OAI21_X1 U544 ( .B1(n1069), .B2(n64), .A(n701), .ZN(n973) );
  NAND2_X1 U545 ( .A1(add_r3[0]), .A2(n1033), .ZN(n701) );
  OAI21_X1 U546 ( .B1(n1069), .B2(n63), .A(n702), .ZN(n974) );
  NAND2_X1 U547 ( .A1(add_r3[1]), .A2(n1033), .ZN(n702) );
  OAI21_X1 U548 ( .B1(n1069), .B2(n62), .A(n703), .ZN(n975) );
  NAND2_X1 U549 ( .A1(add_r3[2]), .A2(n1033), .ZN(n703) );
  OAI21_X1 U550 ( .B1(n1069), .B2(n61), .A(n704), .ZN(n976) );
  NAND2_X1 U551 ( .A1(add_r3[3]), .A2(n1033), .ZN(n704) );
  OAI21_X1 U552 ( .B1(n1069), .B2(n60), .A(n705), .ZN(n977) );
  NAND2_X1 U553 ( .A1(add_r3[4]), .A2(n1033), .ZN(n705) );
  OAI21_X1 U554 ( .B1(n1069), .B2(n59), .A(n706), .ZN(n978) );
  NAND2_X1 U555 ( .A1(add_r3[5]), .A2(n1033), .ZN(n706) );
  OAI21_X1 U556 ( .B1(n1069), .B2(n58), .A(n707), .ZN(n979) );
  NAND2_X1 U557 ( .A1(add_r3[6]), .A2(n1033), .ZN(n707) );
  OAI21_X1 U558 ( .B1(n1069), .B2(n57), .A(n708), .ZN(n980) );
  NAND2_X1 U559 ( .A1(add_r3[7]), .A2(n1033), .ZN(n708) );
  OAI21_X1 U560 ( .B1(n1057), .B2(n246), .A(n519), .ZN(n791) );
  NAND2_X1 U561 ( .A1(add_r15[10]), .A2(n1049), .ZN(n519) );
  OAI21_X1 U562 ( .B1(n1057), .B2(n245), .A(n520), .ZN(n792) );
  NAND2_X1 U563 ( .A1(add_r15[11]), .A2(n1049), .ZN(n520) );
  OAI21_X1 U564 ( .B1(n1058), .B2(n231), .A(n534), .ZN(n806) );
  NAND2_X1 U565 ( .A1(add_r14[9]), .A2(n1047), .ZN(n534) );
  OAI21_X1 U566 ( .B1(n1058), .B2(n230), .A(n535), .ZN(n807) );
  NAND2_X1 U567 ( .A1(add_r14[10]), .A2(n1047), .ZN(n535) );
  OAI21_X1 U568 ( .B1(n1058), .B2(n229), .A(n536), .ZN(n808) );
  NAND2_X1 U569 ( .A1(add_r14[11]), .A2(n1047), .ZN(n536) );
  OAI21_X1 U570 ( .B1(n1061), .B2(n199), .A(n566), .ZN(n838) );
  NAND2_X1 U571 ( .A1(add_r12[9]), .A2(n1045), .ZN(n566) );
  OAI21_X1 U572 ( .B1(n1061), .B2(n198), .A(n567), .ZN(n839) );
  NAND2_X1 U573 ( .A1(add_r12[10]), .A2(n1045), .ZN(n567) );
  OAI21_X1 U574 ( .B1(n1061), .B2(n197), .A(n568), .ZN(n840) );
  NAND2_X1 U575 ( .A1(add_r12[11]), .A2(n1045), .ZN(n568) );
  OAI21_X1 U576 ( .B1(n1062), .B2(n183), .A(n582), .ZN(n854) );
  NAND2_X1 U577 ( .A1(add_r11[9]), .A2(n1043), .ZN(n582) );
  OAI21_X1 U578 ( .B1(n1062), .B2(n182), .A(n583), .ZN(n855) );
  NAND2_X1 U579 ( .A1(add_r11[10]), .A2(n1043), .ZN(n583) );
  OAI21_X1 U580 ( .B1(n1062), .B2(n181), .A(n584), .ZN(n856) );
  NAND2_X1 U581 ( .A1(add_r11[11]), .A2(n1043), .ZN(n584) );
  OAI21_X1 U582 ( .B1(n1066), .B2(n134), .A(n631), .ZN(n903) );
  NAND2_X1 U583 ( .A1(add_r8[10]), .A2(n1039), .ZN(n631) );
  OAI21_X1 U584 ( .B1(n1066), .B2(n133), .A(n632), .ZN(n904) );
  NAND2_X1 U585 ( .A1(add_r8[11]), .A2(n1039), .ZN(n632) );
  OAI21_X1 U586 ( .B1(n1058), .B2(n226), .A(n539), .ZN(n811) );
  NAND2_X1 U587 ( .A1(add_r14[14]), .A2(n1047), .ZN(n539) );
  OAI21_X1 U588 ( .B1(n1062), .B2(n178), .A(n587), .ZN(n859) );
  NAND2_X1 U589 ( .A1(add_r11[14]), .A2(n1043), .ZN(n587) );
  OAI21_X1 U590 ( .B1(n1061), .B2(n194), .A(n571), .ZN(n843) );
  NAND2_X1 U591 ( .A1(add_r12[14]), .A2(n1044), .ZN(n571) );
  OAI21_X1 U592 ( .B1(n1064), .B2(n162), .A(n603), .ZN(n875) );
  NAND2_X1 U593 ( .A1(add_r10[14]), .A2(n1042), .ZN(n603) );
  OAI21_X1 U594 ( .B1(n1060), .B2(n210), .A(n555), .ZN(n827) );
  NAND2_X1 U595 ( .A1(add_r13[14]), .A2(n1046), .ZN(n555) );
  OAI21_X1 U596 ( .B1(n1066), .B2(n130), .A(n635), .ZN(n907) );
  NAND2_X1 U597 ( .A1(add_r8[14]), .A2(n1039), .ZN(n635) );
  OAI21_X1 U598 ( .B1(n1057), .B2(n242), .A(n523), .ZN(n795) );
  NAND2_X1 U599 ( .A1(add_r15[14]), .A2(n1048), .ZN(n523) );
  OAI21_X1 U600 ( .B1(n1058), .B2(n227), .A(n538), .ZN(n810) );
  NAND2_X1 U601 ( .A1(add_r14[13]), .A2(n1047), .ZN(n538) );
  OAI21_X1 U602 ( .B1(n1062), .B2(n179), .A(n586), .ZN(n858) );
  NAND2_X1 U603 ( .A1(add_r11[13]), .A2(n1043), .ZN(n586) );
  OAI21_X1 U604 ( .B1(n1061), .B2(n195), .A(n570), .ZN(n842) );
  NAND2_X1 U605 ( .A1(add_r12[13]), .A2(n1044), .ZN(n570) );
  OAI21_X1 U606 ( .B1(n1064), .B2(n163), .A(n602), .ZN(n874) );
  NAND2_X1 U607 ( .A1(add_r10[13]), .A2(n1042), .ZN(n602) );
  OAI21_X1 U608 ( .B1(n1060), .B2(n211), .A(n554), .ZN(n826) );
  NAND2_X1 U609 ( .A1(add_r13[13]), .A2(n1046), .ZN(n554) );
  OAI21_X1 U610 ( .B1(n1066), .B2(n131), .A(n634), .ZN(n906) );
  NAND2_X1 U611 ( .A1(add_r8[13]), .A2(n1039), .ZN(n634) );
  OAI21_X1 U612 ( .B1(n1057), .B2(n243), .A(n522), .ZN(n794) );
  NAND2_X1 U613 ( .A1(add_r15[13]), .A2(n1048), .ZN(n522) );
  OAI21_X1 U614 ( .B1(n1058), .B2(n228), .A(n537), .ZN(n809) );
  NAND2_X1 U615 ( .A1(add_r14[12]), .A2(n1047), .ZN(n537) );
  OAI21_X1 U616 ( .B1(n1062), .B2(n180), .A(n585), .ZN(n857) );
  NAND2_X1 U617 ( .A1(add_r11[12]), .A2(n1043), .ZN(n585) );
  OAI21_X1 U618 ( .B1(n1061), .B2(n196), .A(n569), .ZN(n841) );
  NAND2_X1 U619 ( .A1(add_r12[12]), .A2(n1044), .ZN(n569) );
  OAI21_X1 U620 ( .B1(n1064), .B2(n164), .A(n601), .ZN(n873) );
  NAND2_X1 U621 ( .A1(add_r10[12]), .A2(n1042), .ZN(n601) );
  OAI21_X1 U622 ( .B1(n1060), .B2(n212), .A(n553), .ZN(n825) );
  NAND2_X1 U623 ( .A1(add_r13[12]), .A2(n1046), .ZN(n553) );
  OAI21_X1 U624 ( .B1(n1066), .B2(n132), .A(n633), .ZN(n905) );
  NAND2_X1 U625 ( .A1(add_r8[12]), .A2(n1039), .ZN(n633) );
  OAI21_X1 U626 ( .B1(n1057), .B2(n244), .A(n521), .ZN(n793) );
  NAND2_X1 U627 ( .A1(add_r15[12]), .A2(n1048), .ZN(n521) );
  OAI21_X1 U628 ( .B1(n1057), .B2(n248), .A(n517), .ZN(n789) );
  NAND2_X1 U629 ( .A1(add_r15[8]), .A2(n1049), .ZN(n517) );
  OAI21_X1 U630 ( .B1(n1057), .B2(n247), .A(n518), .ZN(n790) );
  NAND2_X1 U631 ( .A1(add_r15[9]), .A2(n1049), .ZN(n518) );
  OAI21_X1 U632 ( .B1(n1057), .B2(n240), .A(n525), .ZN(n797) );
  NAND2_X1 U633 ( .A1(add_r14[0]), .A2(n1048), .ZN(n525) );
  OAI21_X1 U634 ( .B1(n1057), .B2(n239), .A(n526), .ZN(n798) );
  NAND2_X1 U635 ( .A1(add_r14[1]), .A2(n1048), .ZN(n526) );
  OAI21_X1 U636 ( .B1(n1057), .B2(n238), .A(n527), .ZN(n799) );
  NAND2_X1 U637 ( .A1(add_r14[2]), .A2(n1048), .ZN(n527) );
  OAI21_X1 U638 ( .B1(n1057), .B2(n237), .A(n528), .ZN(n800) );
  NAND2_X1 U639 ( .A1(add_r14[3]), .A2(n1048), .ZN(n528) );
  OAI21_X1 U640 ( .B1(n1058), .B2(n236), .A(n529), .ZN(n801) );
  NAND2_X1 U641 ( .A1(add_r14[4]), .A2(n1048), .ZN(n529) );
  OAI21_X1 U642 ( .B1(n1058), .B2(n234), .A(n531), .ZN(n803) );
  NAND2_X1 U643 ( .A1(add_r14[6]), .A2(n1048), .ZN(n531) );
  OAI21_X1 U644 ( .B1(n1058), .B2(n233), .A(n532), .ZN(n804) );
  NAND2_X1 U645 ( .A1(add_r14[7]), .A2(n1048), .ZN(n532) );
  OAI21_X1 U646 ( .B1(n1058), .B2(n232), .A(n533), .ZN(n805) );
  NAND2_X1 U647 ( .A1(add_r14[8]), .A2(n1047), .ZN(n533) );
  OAI21_X1 U648 ( .B1(n1060), .B2(n208), .A(n557), .ZN(n829) );
  NAND2_X1 U649 ( .A1(add_r12[0]), .A2(n1045), .ZN(n557) );
  OAI21_X1 U650 ( .B1(n1060), .B2(n207), .A(n558), .ZN(n830) );
  NAND2_X1 U651 ( .A1(add_r12[1]), .A2(n1045), .ZN(n558) );
  OAI21_X1 U652 ( .B1(n1060), .B2(n206), .A(n559), .ZN(n831) );
  NAND2_X1 U653 ( .A1(add_r12[2]), .A2(n1045), .ZN(n559) );
  OAI21_X1 U654 ( .B1(n1060), .B2(n205), .A(n560), .ZN(n832) );
  NAND2_X1 U655 ( .A1(add_r12[3]), .A2(n1045), .ZN(n560) );
  OAI21_X1 U656 ( .B1(n1060), .B2(n204), .A(n561), .ZN(n833) );
  NAND2_X1 U657 ( .A1(add_r12[4]), .A2(n1045), .ZN(n561) );
  OAI21_X1 U658 ( .B1(n1060), .B2(n203), .A(n562), .ZN(n834) );
  NAND2_X1 U659 ( .A1(add_r12[5]), .A2(n1045), .ZN(n562) );
  OAI21_X1 U660 ( .B1(n1060), .B2(n202), .A(n563), .ZN(n835) );
  NAND2_X1 U661 ( .A1(add_r12[6]), .A2(n1045), .ZN(n563) );
  OAI21_X1 U662 ( .B1(n1060), .B2(n201), .A(n564), .ZN(n836) );
  NAND2_X1 U663 ( .A1(add_r12[7]), .A2(n1045), .ZN(n564) );
  OAI21_X1 U664 ( .B1(n1061), .B2(n200), .A(n565), .ZN(n837) );
  NAND2_X1 U665 ( .A1(add_r12[8]), .A2(n1045), .ZN(n565) );
  OAI21_X1 U666 ( .B1(n1062), .B2(n186), .A(n579), .ZN(n851) );
  NAND2_X1 U667 ( .A1(add_r11[6]), .A2(n1044), .ZN(n579) );
  OAI21_X1 U668 ( .B1(n1062), .B2(n185), .A(n580), .ZN(n852) );
  NAND2_X1 U669 ( .A1(add_r11[7]), .A2(n1044), .ZN(n580) );
  OAI21_X1 U670 ( .B1(n1062), .B2(n184), .A(n581), .ZN(n853) );
  NAND2_X1 U671 ( .A1(add_r11[8]), .A2(n1043), .ZN(n581) );
  OAI21_X1 U672 ( .B1(n1064), .B2(n160), .A(n605), .ZN(n877) );
  NAND2_X1 U673 ( .A1(add_r9[0]), .A2(n1041), .ZN(n605) );
  OAI21_X1 U674 ( .B1(n1064), .B2(n159), .A(n606), .ZN(n878) );
  NAND2_X1 U675 ( .A1(add_r9[1]), .A2(n1041), .ZN(n606) );
  OAI21_X1 U676 ( .B1(n1064), .B2(n158), .A(n607), .ZN(n879) );
  NAND2_X1 U677 ( .A1(add_r9[2]), .A2(n1041), .ZN(n607) );
  OAI21_X1 U678 ( .B1(n1064), .B2(n157), .A(n608), .ZN(n880) );
  NAND2_X1 U679 ( .A1(add_r9[3]), .A2(n1041), .ZN(n608) );
  OAI21_X1 U680 ( .B1(n1064), .B2(n156), .A(n609), .ZN(n881) );
  NAND2_X1 U681 ( .A1(add_r9[4]), .A2(n1041), .ZN(n609) );
  OAI21_X1 U682 ( .B1(n1064), .B2(n155), .A(n610), .ZN(n882) );
  NAND2_X1 U683 ( .A1(add_r9[5]), .A2(n1041), .ZN(n610) );
  OAI21_X1 U684 ( .B1(n1064), .B2(n154), .A(n611), .ZN(n883) );
  NAND2_X1 U685 ( .A1(add_r9[6]), .A2(n1041), .ZN(n611) );
  OAI21_X1 U686 ( .B1(n1064), .B2(n153), .A(n612), .ZN(n884) );
  NAND2_X1 U687 ( .A1(add_r9[7]), .A2(n1041), .ZN(n612) );
  OAI21_X1 U688 ( .B1(n1066), .B2(n140), .A(n625), .ZN(n897) );
  NAND2_X1 U689 ( .A1(add_r8[4]), .A2(n1040), .ZN(n625) );
  OAI21_X1 U690 ( .B1(n1066), .B2(n139), .A(n626), .ZN(n898) );
  NAND2_X1 U691 ( .A1(add_r8[5]), .A2(n1040), .ZN(n626) );
  OAI21_X1 U692 ( .B1(n1066), .B2(n138), .A(n627), .ZN(n899) );
  NAND2_X1 U693 ( .A1(add_r8[6]), .A2(n1040), .ZN(n627) );
  OAI21_X1 U694 ( .B1(n1066), .B2(n137), .A(n628), .ZN(n900) );
  NAND2_X1 U695 ( .A1(add_r8[7]), .A2(n1040), .ZN(n628) );
  OAI21_X1 U696 ( .B1(n1066), .B2(n136), .A(n629), .ZN(n901) );
  NAND2_X1 U697 ( .A1(add_r8[8]), .A2(n1039), .ZN(n629) );
  OAI21_X1 U698 ( .B1(n1066), .B2(n135), .A(n630), .ZN(n902) );
  NAND2_X1 U699 ( .A1(add_r8[9]), .A2(n1039), .ZN(n630) );
  OAI21_X1 U700 ( .B1(n1070), .B2(n54), .A(n711), .ZN(n983) );
  NAND2_X1 U701 ( .A1(add_r3[10]), .A2(n1033), .ZN(n711) );
  OAI21_X1 U702 ( .B1(n1070), .B2(n53), .A(n712), .ZN(n984) );
  NAND2_X1 U703 ( .A1(add_r3[11]), .A2(n1033), .ZN(n712) );
  OAI21_X1 U704 ( .B1(n1071), .B2(n38), .A(n727), .ZN(n999) );
  NAND2_X1 U705 ( .A1(add_r2[10]), .A2(n1031), .ZN(n727) );
  OAI21_X1 U706 ( .B1(n1071), .B2(n37), .A(n728), .ZN(n1000) );
  NAND2_X1 U707 ( .A1(add_r2[11]), .A2(n1031), .ZN(n728) );
  OAI21_X1 U708 ( .B1(n1071), .B2(n34), .A(n731), .ZN(n1003) );
  NAND2_X1 U709 ( .A1(add_r2[14]), .A2(n1031), .ZN(n731) );
  NAND2_X1 U710 ( .A1(add_r3[14]), .A2(n1032), .ZN(n715) );
  OAI21_X1 U711 ( .B1(n1071), .B2(n35), .A(n730), .ZN(n1002) );
  NAND2_X1 U712 ( .A1(add_r2[13]), .A2(n1031), .ZN(n730) );
  OAI21_X1 U713 ( .B1(n1070), .B2(n51), .A(n714), .ZN(n986) );
  NAND2_X1 U714 ( .A1(add_r3[13]), .A2(n1032), .ZN(n714) );
  OAI21_X1 U715 ( .B1(n1071), .B2(n36), .A(n729), .ZN(n1001) );
  NAND2_X1 U716 ( .A1(add_r2[12]), .A2(n1031), .ZN(n729) );
  OAI21_X1 U717 ( .B1(n1070), .B2(n52), .A(n713), .ZN(n985) );
  NAND2_X1 U718 ( .A1(add_r3[12]), .A2(n1032), .ZN(n713) );
  OAI21_X1 U719 ( .B1(n1070), .B2(n56), .A(n709), .ZN(n981) );
  NAND2_X1 U720 ( .A1(add_r3[8]), .A2(n1033), .ZN(n709) );
  OAI21_X1 U721 ( .B1(n1070), .B2(n55), .A(n710), .ZN(n982) );
  NAND2_X1 U722 ( .A1(add_r3[9]), .A2(n1033), .ZN(n710) );
  OAI21_X1 U723 ( .B1(n1071), .B2(n42), .A(n723), .ZN(n995) );
  NAND2_X1 U724 ( .A1(add_r2[6]), .A2(n1032), .ZN(n723) );
  OAI21_X1 U725 ( .B1(n1071), .B2(n41), .A(n724), .ZN(n996) );
  NAND2_X1 U726 ( .A1(add_r2[7]), .A2(n1032), .ZN(n724) );
  OAI21_X1 U727 ( .B1(n1071), .B2(n40), .A(n725), .ZN(n997) );
  NAND2_X1 U728 ( .A1(add_r2[8]), .A2(n1031), .ZN(n725) );
  OAI21_X1 U729 ( .B1(n1071), .B2(n39), .A(n726), .ZN(n998) );
  NAND2_X1 U730 ( .A1(add_r2[9]), .A2(n1031), .ZN(n726) );
  OAI21_X1 U731 ( .B1(n1059), .B2(n224), .A(n541), .ZN(n813) );
  NAND2_X1 U732 ( .A1(add_r13[0]), .A2(n1047), .ZN(n541) );
  OAI21_X1 U733 ( .B1(n1059), .B2(n223), .A(n542), .ZN(n814) );
  NAND2_X1 U734 ( .A1(add_r13[1]), .A2(n1047), .ZN(n542) );
  OAI21_X1 U735 ( .B1(n1059), .B2(n222), .A(n543), .ZN(n815) );
  NAND2_X1 U736 ( .A1(add_r13[2]), .A2(n1047), .ZN(n543) );
  OAI21_X1 U737 ( .B1(n1059), .B2(n221), .A(n544), .ZN(n816) );
  NAND2_X1 U738 ( .A1(add_r13[3]), .A2(n1047), .ZN(n544) );
  OAI21_X1 U739 ( .B1(n1061), .B2(n192), .A(n573), .ZN(n845) );
  NAND2_X1 U740 ( .A1(add_r11[0]), .A2(n1044), .ZN(n573) );
  OAI21_X1 U741 ( .B1(n1061), .B2(n191), .A(n574), .ZN(n846) );
  NAND2_X1 U742 ( .A1(add_r11[1]), .A2(n1044), .ZN(n574) );
  OAI21_X1 U743 ( .B1(n1061), .B2(n190), .A(n575), .ZN(n847) );
  NAND2_X1 U744 ( .A1(add_r11[2]), .A2(n1044), .ZN(n575) );
  OAI21_X1 U745 ( .B1(n1061), .B2(n189), .A(n576), .ZN(n848) );
  NAND2_X1 U746 ( .A1(add_r11[3]), .A2(n1044), .ZN(n576) );
  OAI21_X1 U747 ( .B1(n1062), .B2(n188), .A(n577), .ZN(n849) );
  NAND2_X1 U748 ( .A1(add_r11[4]), .A2(n1044), .ZN(n577) );
  OAI21_X1 U749 ( .B1(n1062), .B2(n187), .A(n578), .ZN(n850) );
  NAND2_X1 U750 ( .A1(add_r11[5]), .A2(n1044), .ZN(n578) );
  OAI21_X1 U751 ( .B1(n1063), .B2(n176), .A(n589), .ZN(n861) );
  NAND2_X1 U752 ( .A1(add_r10[0]), .A2(n1043), .ZN(n589) );
  OAI21_X1 U753 ( .B1(n1063), .B2(n175), .A(n590), .ZN(n862) );
  NAND2_X1 U754 ( .A1(add_r10[1]), .A2(n1043), .ZN(n590) );
  OAI21_X1 U755 ( .B1(n1063), .B2(n174), .A(n591), .ZN(n863) );
  NAND2_X1 U756 ( .A1(add_r10[2]), .A2(n1043), .ZN(n591) );
  OAI21_X1 U757 ( .B1(n1063), .B2(n173), .A(n592), .ZN(n864) );
  NAND2_X1 U758 ( .A1(add_r10[3]), .A2(n1043), .ZN(n592) );
  OAI21_X1 U759 ( .B1(n1063), .B2(n172), .A(n593), .ZN(n865) );
  NAND2_X1 U760 ( .A1(add_r10[4]), .A2(n1042), .ZN(n593) );
  OAI21_X1 U761 ( .B1(n1063), .B2(n171), .A(n594), .ZN(n866) );
  NAND2_X1 U762 ( .A1(add_r10[5]), .A2(n1042), .ZN(n594) );
  OAI21_X1 U763 ( .B1(n1065), .B2(n144), .A(n621), .ZN(n893) );
  NAND2_X1 U764 ( .A1(add_r8[0]), .A2(n1040), .ZN(n621) );
  OAI21_X1 U765 ( .B1(n1065), .B2(n143), .A(n622), .ZN(n894) );
  NAND2_X1 U766 ( .A1(add_r8[1]), .A2(n1040), .ZN(n622) );
  OAI21_X1 U767 ( .B1(n1065), .B2(n142), .A(n623), .ZN(n895) );
  NAND2_X1 U768 ( .A1(add_r8[2]), .A2(n1040), .ZN(n623) );
  OAI21_X1 U769 ( .B1(n1065), .B2(n141), .A(n624), .ZN(n896) );
  NAND2_X1 U770 ( .A1(add_r8[3]), .A2(n1040), .ZN(n624) );
  OAI21_X1 U771 ( .B1(n1065), .B2(n128), .A(n637), .ZN(n909) );
  NAND2_X1 U772 ( .A1(add_r7[0]), .A2(n1039), .ZN(n637) );
  OAI21_X1 U773 ( .B1(n1063), .B2(n127), .A(n638), .ZN(n910) );
  NAND2_X1 U774 ( .A1(add_r7[1]), .A2(n1039), .ZN(n638) );
  OAI21_X1 U775 ( .B1(n1055), .B2(n126), .A(n639), .ZN(n911) );
  NAND2_X1 U776 ( .A1(add_r7[2]), .A2(n1039), .ZN(n639) );
  OAI21_X1 U777 ( .B1(n1059), .B2(n125), .A(n640), .ZN(n912) );
  NAND2_X1 U778 ( .A1(add_r7[3]), .A2(n1039), .ZN(n640) );
  OAI21_X1 U779 ( .B1(n1072), .B2(n96), .A(n669), .ZN(n941) );
  NAND2_X1 U780 ( .A1(add_r5[0]), .A2(n1036), .ZN(n669) );
  OAI21_X1 U781 ( .B1(n1070), .B2(n95), .A(n670), .ZN(n942) );
  NAND2_X1 U782 ( .A1(add_r5[1]), .A2(n1036), .ZN(n670) );
  OAI21_X1 U783 ( .B1(n1071), .B2(n94), .A(n671), .ZN(n943) );
  NAND2_X1 U784 ( .A1(add_r5[2]), .A2(n1036), .ZN(n671) );
  OAI21_X1 U785 ( .B1(n1072), .B2(n93), .A(n672), .ZN(n944) );
  NAND2_X1 U786 ( .A1(add_r5[3]), .A2(n1036), .ZN(n672) );
  OAI21_X1 U787 ( .B1(n1068), .B2(n80), .A(n685), .ZN(n957) );
  NAND2_X1 U788 ( .A1(add_r4[0]), .A2(n1035), .ZN(n685) );
  OAI21_X1 U789 ( .B1(n1068), .B2(n79), .A(n686), .ZN(n958) );
  NAND2_X1 U790 ( .A1(add_r4[1]), .A2(n1035), .ZN(n686) );
  OAI21_X1 U791 ( .B1(n1068), .B2(n78), .A(n687), .ZN(n959) );
  NAND2_X1 U792 ( .A1(add_r4[2]), .A2(n1035), .ZN(n687) );
  OAI21_X1 U793 ( .B1(n1068), .B2(n77), .A(n688), .ZN(n960) );
  NAND2_X1 U794 ( .A1(add_r4[3]), .A2(n1035), .ZN(n688) );
  OAI21_X1 U795 ( .B1(n1068), .B2(n76), .A(n689), .ZN(n961) );
  NAND2_X1 U796 ( .A1(add_r4[4]), .A2(n1034), .ZN(n689) );
  OAI21_X1 U797 ( .B1(n1070), .B2(n48), .A(n717), .ZN(n989) );
  NAND2_X1 U798 ( .A1(add_r2[0]), .A2(n1032), .ZN(n717) );
  OAI21_X1 U799 ( .B1(n1070), .B2(n47), .A(n718), .ZN(n990) );
  NAND2_X1 U800 ( .A1(add_r2[1]), .A2(n1032), .ZN(n718) );
  OAI21_X1 U801 ( .B1(n1070), .B2(n46), .A(n719), .ZN(n991) );
  NAND2_X1 U802 ( .A1(add_r2[2]), .A2(n1032), .ZN(n719) );
  OAI21_X1 U803 ( .B1(n1070), .B2(n45), .A(n720), .ZN(n992) );
  NAND2_X1 U804 ( .A1(add_r2[3]), .A2(n1032), .ZN(n720) );
  OAI21_X1 U805 ( .B1(n1071), .B2(n44), .A(n721), .ZN(n993) );
  NAND2_X1 U806 ( .A1(add_r2[4]), .A2(n1032), .ZN(n721) );
  OAI21_X1 U807 ( .B1(n1071), .B2(n43), .A(n722), .ZN(n994) );
  NAND2_X1 U808 ( .A1(add_r2[5]), .A2(n1032), .ZN(n722) );
  OAI21_X1 U809 ( .B1(n1072), .B2(n32), .A(n733), .ZN(n1005) );
  NAND2_X1 U810 ( .A1(add_r1[0]), .A2(n1031), .ZN(n733) );
  OAI21_X1 U811 ( .B1(n1072), .B2(n31), .A(n734), .ZN(n1006) );
  NAND2_X1 U812 ( .A1(add_r1[1]), .A2(n1031), .ZN(n734) );
  OAI21_X1 U813 ( .B1(n1072), .B2(n30), .A(n735), .ZN(n1007) );
  NAND2_X1 U814 ( .A1(add_r1[2]), .A2(n1031), .ZN(n735) );
  OAI21_X1 U815 ( .B1(n1072), .B2(n29), .A(n736), .ZN(n1008) );
  NAND2_X1 U816 ( .A1(add_r1[3]), .A2(n1031), .ZN(n736) );
  OAI21_X1 U817 ( .B1(n1055), .B2(n267), .A(n498), .ZN(n770) );
  NAND2_X1 U818 ( .A1(add_r16[5]), .A2(n1050), .ZN(n498) );
  OAI21_X1 U819 ( .B1(n1058), .B2(n235), .A(n530), .ZN(n802) );
  NAND2_X1 U820 ( .A1(add_r14[5]), .A2(n1048), .ZN(n530) );
  OR2_X1 U821 ( .A1(n1056), .A2(n257), .ZN(n285) );
  NAND2_X1 U822 ( .A1(n508), .A2(n285), .ZN(n780) );
  BUF_X1 U823 ( .A(n1052), .Z(n1056) );
  OR2_X1 U824 ( .A1(n1065), .A2(n145), .ZN(n286) );
  NAND2_X1 U825 ( .A1(n620), .A2(n286), .ZN(n892) );
  BUF_X1 U826 ( .A(n1053), .Z(n1065) );
  OR2_X1 U827 ( .A1(n1071), .A2(n17), .ZN(n1023) );
  NAND2_X1 U828 ( .A1(n748), .A2(n1023), .ZN(n1020) );
  NAND2_X1 U829 ( .A1(add_r15[15]), .A2(n1048), .ZN(n524) );
  NAND2_X1 U830 ( .A1(add_r16[15]), .A2(n1050), .ZN(n508) );
  NAND2_X1 U831 ( .A1(add_r2[15]), .A2(n1031), .ZN(n732) );
  NAND2_X1 U832 ( .A1(add_r3[15]), .A2(n1032), .ZN(n716) );
  NAND2_X1 U833 ( .A1(add_r4[15]), .A2(n1034), .ZN(n700) );
  NAND2_X1 U834 ( .A1(add_r5[15]), .A2(n1035), .ZN(n684) );
  NAND2_X1 U835 ( .A1(add_r6[15]), .A2(n1036), .ZN(n668) );
  NAND2_X1 U836 ( .A1(add_r7[15]), .A2(n1038), .ZN(n652) );
  NAND2_X1 U837 ( .A1(add_r8[15]), .A2(n1039), .ZN(n636) );
  NAND2_X1 U838 ( .A1(add_r9[15]), .A2(n1040), .ZN(n620) );
  NAND2_X1 U839 ( .A1(add_r10[15]), .A2(n1042), .ZN(n604) );
  NAND2_X1 U840 ( .A1(add_r11[15]), .A2(n1043), .ZN(n588) );
  NAND2_X1 U841 ( .A1(add_r12[15]), .A2(n1044), .ZN(n572) );
  NAND2_X1 U842 ( .A1(add_r13[15]), .A2(n1046), .ZN(n556) );
  NAND2_X1 U843 ( .A1(add_r14[15]), .A2(n1047), .ZN(n540) );
  NAND2_X1 U844 ( .A1(add_r1[15]), .A2(n1030), .ZN(n748) );
  CLKBUF_X1 U845 ( .A(n1027), .Z(n1051) );
  INV_X1 U846 ( .A(addr_y[0]), .ZN(n1088) );
  INV_X1 U847 ( .A(addr_y[1]), .ZN(n1089) );
endmodule


module ctrlpath ( clk, reset, start, addr_x, wr_en_x, addr_a1, addr_a2, 
        addr_a3, addr_a4, addr_a5, addr_a6, addr_a7, addr_a8, addr_a9, 
        addr_a10, addr_a11, addr_a12, addr_a13, addr_a14, addr_a15, addr_a16, 
        wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6, wr_en_a7, 
        wr_en_a8, wr_en_a9, wr_en_a10, wr_en_a11, wr_en_a12, wr_en_a13, 
        wr_en_a14, wr_en_a15, wr_en_a16, clear_acc, clc, clc1, addr_y, wr_en_y, 
        done, loadMatrix, loadVector );
  output [3:0] addr_x;
  output [3:0] addr_a1;
  output [3:0] addr_a2;
  output [3:0] addr_a3;
  output [3:0] addr_a4;
  output [3:0] addr_a5;
  output [3:0] addr_a6;
  output [3:0] addr_a7;
  output [3:0] addr_a8;
  output [3:0] addr_a9;
  output [3:0] addr_a10;
  output [3:0] addr_a11;
  output [3:0] addr_a12;
  output [3:0] addr_a13;
  output [3:0] addr_a14;
  output [3:0] addr_a15;
  output [3:0] addr_a16;
  output [3:0] addr_y;
  input clk, reset, start, loadMatrix, loadVector;
  output wr_en_x, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6,
         wr_en_a7, wr_en_a8, wr_en_a9, wr_en_a10, wr_en_a11, wr_en_a12,
         wr_en_a13, wr_en_a14, wr_en_a15, wr_en_a16, clear_acc, clc, clc1,
         wr_en_y, done;
  wire   N48, N49, N50, N51, N52, N53, N61, N62, N63, N64, N74, N75, N76, N77,
         N87, N88, N89, N90, N100, N101, N102, N103, N113, N114, N115, N116,
         N126, N127, N128, N129, N139, N140, N141, N142, N152, N153, N154,
         N155, N165, N166, N167, N168, N178, N179, N180, N181, N191, N192,
         N193, N194, N204, N205, N206, N207, N217, N218, N219, N220, N230,
         N231, N232, N233, N243, N244, N245, N246, N256, N257, N258, N259,
         N268, N269, N270, N271, N280, N281, N282, N283, N286, N287, N288,
         n140, n145, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n213, n214,
         n215, n216, n218, n219, n220, n222, n223, n224, n225, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75;
  wire   [4:0] state;

  DFF_X1 \addr_y_reg[0]  ( .D(N280), .CK(clk), .Q(addr_y[0]), .QN(n225) );
  DFF_X1 \addr_y_reg[2]  ( .D(N282), .CK(clk), .Q(addr_y[2]), .QN(n223) );
  DFF_X1 \addr_y_reg[3]  ( .D(N283), .CK(clk), .Q(addr_y[3]), .QN(n222) );
  DFF_X1 \state_reg[0]  ( .D(N48), .CK(clk), .Q(state[0]), .QN(n148) );
  DFF_X1 \addr_a16_reg[1]  ( .D(N257), .CK(clk), .Q(addr_a16[1]), .QN(n215) );
  DFF_X1 \addr_a16_reg[3]  ( .D(N259), .CK(clk), .Q(addr_a16[3]), .QN(n213) );
  DFF_X1 \state_reg[4]  ( .D(N52), .CK(clk), .Q(state[4]), .QN(n140) );
  DFF_X1 \addr_a15_reg[1]  ( .D(N244), .CK(clk), .Q(addr_a15[1]), .QN(n210) );
  DFF_X1 \addr_a15_reg[3]  ( .D(N246), .CK(clk), .Q(addr_a15[3]), .QN(n208) );
  DFF_X1 \state_reg[1]  ( .D(N49), .CK(clk), .Q(state[1]), .QN(n147) );
  DFF_X1 \addr_a13_reg[1]  ( .D(N218), .CK(clk), .Q(addr_a13[1]), .QN(n202) );
  DFF_X1 \addr_a13_reg[3]  ( .D(N220), .CK(clk), .Q(addr_a13[3]), .QN(n199) );
  DFF_X1 \state_reg[2]  ( .D(N50), .CK(clk), .Q(state[2]), .QN(n145) );
  DFF_X1 \addr_a5_reg[1]  ( .D(N114), .CK(clk), .Q(addr_a5[1]), .QN(n168) );
  DFF_X1 \addr_a5_reg[3]  ( .D(N116), .CK(clk), .Q(addr_a5[3]), .QN(n166) );
  DFF_X1 \state_reg[3]  ( .D(N51), .CK(clk), .Q(state[3]) );
  DFF_X1 \addr_y_reg[1]  ( .D(N281), .CK(clk), .Q(addr_y[1]), .QN(n224) );
  DFF_X1 done_reg ( .D(N53), .CK(clk), .Q(done) );
  DFF_X1 \addr_x_reg[0]  ( .D(N268), .CK(clk), .Q(addr_x[0]) );
  DFF_X1 \addr_x_reg[1]  ( .D(N269), .CK(clk), .Q(addr_x[1]), .QN(n220) );
  DFF_X1 \addr_x_reg[2]  ( .D(N270), .CK(clk), .Q(addr_x[2]), .QN(n219) );
  DFF_X1 \addr_x_reg[3]  ( .D(N271), .CK(clk), .Q(addr_x[3]), .QN(n218) );
  DFF_X1 \addr_a16_reg[0]  ( .D(N256), .CK(clk), .Q(addr_a16[0]), .QN(n216) );
  DFF_X1 \addr_a16_reg[2]  ( .D(N258), .CK(clk), .Q(addr_a16[2]), .QN(n214) );
  DFF_X1 \addr_a15_reg[0]  ( .D(N243), .CK(clk), .Q(addr_a15[0]), .QN(n211) );
  DFF_X1 \addr_a15_reg[2]  ( .D(N245), .CK(clk), .Q(addr_a15[2]), .QN(n209) );
  DFF_X1 \addr_a13_reg[0]  ( .D(N217), .CK(clk), .Q(addr_a13[0]), .QN(n203) );
  DFF_X1 \addr_a13_reg[2]  ( .D(N219), .CK(clk), .Q(addr_a13[2]), .QN(n201) );
  DFF_X1 \addr_a5_reg[0]  ( .D(N113), .CK(clk), .Q(addr_a5[0]), .QN(n169) );
  DFF_X1 \addr_a5_reg[2]  ( .D(N115), .CK(clk), .Q(addr_a5[2]), .QN(n167) );
  DFF_X1 \addr_a3_reg[0]  ( .D(N87), .CK(clk), .Q(addr_a3[0]), .QN(n161) );
  DFF_X1 \addr_a3_reg[1]  ( .D(N88), .CK(clk), .Q(addr_a3[1]), .QN(n160) );
  DFF_X1 \addr_a3_reg[2]  ( .D(N89), .CK(clk), .Q(addr_a3[2]), .QN(n159) );
  DFF_X1 \addr_a3_reg[3]  ( .D(N90), .CK(clk), .Q(addr_a3[3]), .QN(n157) );
  DFF_X1 \addr_a2_reg[0]  ( .D(N74), .CK(clk), .Q(addr_a2[0]), .QN(n156) );
  DFF_X1 \addr_a2_reg[1]  ( .D(N75), .CK(clk), .Q(addr_a2[1]), .QN(n155) );
  DFF_X1 \addr_a2_reg[2]  ( .D(N76), .CK(clk), .Q(addr_a2[2]), .QN(n154) );
  DFF_X1 \addr_a2_reg[3]  ( .D(N77), .CK(clk), .Q(addr_a2[3]), .QN(n153) );
  DFF_X1 \addr_a1_reg[0]  ( .D(N61), .CK(clk), .Q(addr_a1[0]), .QN(n152) );
  DFF_X1 \addr_a1_reg[1]  ( .D(N62), .CK(clk), .Q(addr_a1[1]), .QN(n151) );
  DFF_X1 \addr_a1_reg[2]  ( .D(N63), .CK(clk), .Q(addr_a1[2]), .QN(n150) );
  DFF_X1 \addr_a1_reg[3]  ( .D(N64), .CK(clk), .Q(addr_a1[3]), .QN(n149) );
  DFF_X1 \addr_a10_reg[0]  ( .D(N178), .CK(clk), .Q(addr_a10[0]), .QN(n189) );
  DFF_X1 \addr_a10_reg[1]  ( .D(N179), .CK(clk), .Q(addr_a10[1]), .QN(n188) );
  DFF_X1 \addr_a10_reg[2]  ( .D(N180), .CK(clk), .Q(addr_a10[2]), .QN(n187) );
  DFF_X1 \addr_a10_reg[3]  ( .D(N181), .CK(clk), .Q(addr_a10[3]), .QN(n186) );
  DFF_X1 \addr_a8_reg[0]  ( .D(N152), .CK(clk), .Q(addr_a8[0]), .QN(n181) );
  DFF_X1 \addr_a8_reg[1]  ( .D(N153), .CK(clk), .Q(addr_a8[1]), .QN(n180) );
  DFF_X1 \addr_a8_reg[2]  ( .D(N154), .CK(clk), .Q(addr_a8[2]), .QN(n179) );
  DFF_X1 \addr_a8_reg[3]  ( .D(N155), .CK(clk), .Q(addr_a8[3]), .QN(n178) );
  DFF_X1 \addr_a7_reg[0]  ( .D(N139), .CK(clk), .Q(addr_a7[0]), .QN(n177) );
  DFF_X1 \addr_a7_reg[1]  ( .D(N140), .CK(clk), .Q(addr_a7[1]), .QN(n176) );
  DFF_X1 \addr_a7_reg[2]  ( .D(N141), .CK(clk), .Q(addr_a7[2]), .QN(n175) );
  DFF_X1 \addr_a7_reg[3]  ( .D(N142), .CK(clk), .Q(addr_a7[3]), .QN(n174) );
  DFF_X1 \addr_a6_reg[0]  ( .D(N126), .CK(clk), .Q(addr_a6[0]), .QN(n173) );
  DFF_X1 \addr_a6_reg[1]  ( .D(N127), .CK(clk), .Q(addr_a6[1]), .QN(n172) );
  DFF_X1 \addr_a6_reg[2]  ( .D(N128), .CK(clk), .Q(addr_a6[2]), .QN(n171) );
  DFF_X1 \addr_a6_reg[3]  ( .D(N129), .CK(clk), .Q(addr_a6[3]), .QN(n170) );
  DFF_X1 \addr_a14_reg[0]  ( .D(N230), .CK(clk), .Q(addr_a14[0]), .QN(n207) );
  DFF_X1 \addr_a14_reg[1]  ( .D(N231), .CK(clk), .Q(addr_a14[1]), .QN(n206) );
  DFF_X1 \addr_a14_reg[2]  ( .D(N232), .CK(clk), .Q(addr_a14[2]), .QN(n205) );
  DFF_X1 \addr_a14_reg[3]  ( .D(N233), .CK(clk), .Q(addr_a14[3]), .QN(n204) );
  DFF_X1 \addr_a11_reg[0]  ( .D(N191), .CK(clk), .Q(addr_a11[0]), .QN(n194) );
  DFF_X1 \addr_a11_reg[1]  ( .D(N192), .CK(clk), .Q(addr_a11[1]), .QN(n193) );
  DFF_X1 \addr_a11_reg[2]  ( .D(N193), .CK(clk), .Q(addr_a11[2]), .QN(n192) );
  DFF_X1 \addr_a11_reg[3]  ( .D(N194), .CK(clk), .Q(addr_a11[3]), .QN(n191) );
  DFF_X1 \addr_a4_reg[0]  ( .D(N100), .CK(clk), .Q(addr_a4[0]), .QN(n165) );
  DFF_X1 \addr_a4_reg[1]  ( .D(N101), .CK(clk), .Q(addr_a4[1]), .QN(n164) );
  DFF_X1 \addr_a4_reg[2]  ( .D(N102), .CK(clk), .Q(addr_a4[2]), .QN(n163) );
  DFF_X1 \addr_a4_reg[3]  ( .D(N103), .CK(clk), .Q(addr_a4[3]), .QN(n162) );
  DFF_X1 \addr_a9_reg[0]  ( .D(N165), .CK(clk), .Q(addr_a9[0]), .QN(n185) );
  DFF_X1 \addr_a9_reg[1]  ( .D(N166), .CK(clk), .Q(addr_a9[1]), .QN(n184) );
  DFF_X1 \addr_a9_reg[2]  ( .D(N167), .CK(clk), .Q(addr_a9[2]), .QN(n183) );
  DFF_X1 \addr_a9_reg[3]  ( .D(N168), .CK(clk), .Q(addr_a9[3]), .QN(n182) );
  DFF_X1 \addr_a12_reg[0]  ( .D(N204), .CK(clk), .Q(addr_a12[0]), .QN(n198) );
  DFF_X1 \addr_a12_reg[1]  ( .D(N205), .CK(clk), .Q(addr_a12[1]), .QN(n197) );
  DFF_X1 \addr_a12_reg[2]  ( .D(N206), .CK(clk), .Q(addr_a12[2]), .QN(n196) );
  DFF_X1 \addr_a12_reg[3]  ( .D(N207), .CK(clk), .Q(addr_a12[3]), .QN(n195) );
  DFF_X1 clear_acc_reg ( .D(N286), .CK(clk), .Q(clear_acc) );
  DFF_X1 clc_reg ( .D(N287), .CK(clk), .Q(clc) );
  DFF_X1 clc1_reg ( .D(N288), .CK(clk), .Q(clc1) );
  NAND3_X1 U394 ( .A1(n247), .A2(n157), .A3(n248), .ZN(n246) );
  NAND3_X1 U395 ( .A1(n247), .A2(n160), .A3(addr_a3[0]), .ZN(n252) );
  NAND3_X1 U396 ( .A1(n256), .A2(n236), .A3(n257), .ZN(n255) );
  NAND3_X1 U397 ( .A1(n261), .A2(n155), .A3(addr_a2[0]), .ZN(n265) );
  NAND3_X1 U398 ( .A1(n256), .A2(n235), .A3(n257), .ZN(n266) );
  NAND3_X1 U399 ( .A1(n269), .A2(n149), .A3(n270), .ZN(n268) );
  NAND3_X1 U400 ( .A1(n269), .A2(n151), .A3(addr_a1[0]), .ZN(n274) );
  NAND3_X1 U401 ( .A1(n307), .A2(n75), .A3(loadVector), .ZN(n305) );
  OAI33_X1 U402 ( .A1(n170), .A2(n232), .A3(n321), .B1(n162), .B2(n234), .B3(
        n322), .ZN(n320) );
  OAI33_X1 U403 ( .A1(n195), .A2(n241), .A3(n324), .B1(n186), .B2(n243), .B3(
        n325), .ZN(n318) );
  OAI33_X1 U404 ( .A1(n153), .A2(n236), .A3(n260), .B1(n204), .B2(n239), .B3(
        n328), .ZN(n327) );
  NAND3_X1 U405 ( .A1(addr_a2[1]), .A2(addr_a2[0]), .A3(addr_a2[2]), .ZN(n260)
         );
  NAND3_X1 U406 ( .A1(n342), .A2(n222), .A3(n350), .ZN(n349) );
  NAND3_X1 U407 ( .A1(addr_y[0]), .A2(n224), .A3(n350), .ZN(n354) );
  NAND3_X1 U408 ( .A1(n355), .A2(n57), .A3(addr_y[0]), .ZN(n356) );
  NAND3_X1 U409 ( .A1(n366), .A2(n213), .A3(n343), .ZN(n365) );
  NAND3_X1 U410 ( .A1(n366), .A2(n215), .A3(addr_a16[0]), .ZN(n370) );
  NAND3_X1 U411 ( .A1(n375), .A2(n208), .A3(n376), .ZN(n374) );
  NAND3_X1 U412 ( .A1(n375), .A2(n210), .A3(addr_a15[0]), .ZN(n380) );
  NAND3_X1 U413 ( .A1(addr_a14[1]), .A2(addr_a14[0]), .A3(addr_a14[2]), .ZN(
        n328) );
  NAND3_X1 U414 ( .A1(n384), .A2(n206), .A3(addr_a14[0]), .ZN(n388) );
  NAND3_X1 U415 ( .A1(n51), .A2(n240), .A3(n39), .ZN(n389) );
  NAND3_X1 U416 ( .A1(n392), .A2(n199), .A3(n393), .ZN(n391) );
  NAND3_X1 U417 ( .A1(n392), .A2(n202), .A3(addr_a13[0]), .ZN(n397) );
  NAND3_X1 U418 ( .A1(addr_a12[1]), .A2(addr_a12[0]), .A3(addr_a12[2]), .ZN(
        n324) );
  NAND3_X1 U419 ( .A1(n402), .A2(n197), .A3(addr_a12[0]), .ZN(n406) );
  NAND3_X1 U420 ( .A1(n410), .A2(n191), .A3(n344), .ZN(n409) );
  NAND3_X1 U421 ( .A1(n410), .A2(n193), .A3(addr_a11[0]), .ZN(n414) );
  NAND3_X1 U422 ( .A1(addr_a10[1]), .A2(addr_a10[0]), .A3(addr_a10[2]), .ZN(
        n325) );
  NAND3_X1 U423 ( .A1(n418), .A2(n188), .A3(addr_a10[0]), .ZN(n422) );
  NAND3_X1 U424 ( .A1(n242), .A2(n232), .A3(n42), .ZN(n399) );
  NAND3_X1 U425 ( .A1(n427), .A2(n182), .A3(n335), .ZN(n426) );
  NAND3_X1 U426 ( .A1(n427), .A2(n184), .A3(addr_a9[0]), .ZN(n431) );
  NAND3_X1 U427 ( .A1(n436), .A2(n178), .A3(n323), .ZN(n435) );
  NAND3_X1 U428 ( .A1(n436), .A2(n180), .A3(addr_a8[0]), .ZN(n440) );
  NAND3_X1 U429 ( .A1(n444), .A2(n174), .A3(n333), .ZN(n443) );
  NAND3_X1 U430 ( .A1(n444), .A2(n176), .A3(addr_a7[0]), .ZN(n448) );
  NAND3_X1 U431 ( .A1(addr_a6[1]), .A2(addr_a6[0]), .A3(addr_a6[2]), .ZN(n321)
         );
  NAND3_X1 U432 ( .A1(n453), .A2(n172), .A3(addr_a6[0]), .ZN(n457) );
  NAND3_X1 U433 ( .A1(n461), .A2(n166), .A3(n462), .ZN(n460) );
  NAND3_X1 U434 ( .A1(n461), .A2(n168), .A3(addr_a5[0]), .ZN(n466) );
  NAND3_X1 U435 ( .A1(addr_a4[1]), .A2(addr_a4[0]), .A3(addr_a4[2]), .ZN(n322)
         );
  NAND3_X1 U436 ( .A1(n472), .A2(n164), .A3(addr_a4[0]), .ZN(n476) );
  NAND3_X1 U437 ( .A1(addr_x[1]), .A2(addr_x[0]), .A3(addr_x[2]), .ZN(n359) );
  NAND3_X1 U438 ( .A1(n276), .A2(n233), .A3(n449), .ZN(n371) );
  NAND3_X1 U439 ( .A1(n243), .A2(n242), .A3(n45), .ZN(n458) );
  NAND3_X1 U440 ( .A1(n240), .A2(n239), .A3(n241), .ZN(n423) );
  NOR2_X1 U3 ( .A1(n140), .A2(state[3]), .ZN(n488) );
  NOR2_X1 U4 ( .A1(state[4]), .A2(state[3]), .ZN(n358) );
  INV_X1 U5 ( .A(n418), .ZN(n17) );
  INV_X1 U6 ( .A(n472), .ZN(n11) );
  INV_X1 U7 ( .A(n453), .ZN(n15) );
  INV_X1 U8 ( .A(n468), .ZN(n58) );
  INV_X1 U9 ( .A(n444), .ZN(n5) );
  INV_X1 U10 ( .A(n269), .ZN(n32) );
  NOR3_X1 U11 ( .A1(n52), .A2(n67), .A3(n58), .ZN(n277) );
  OAI21_X1 U12 ( .B1(n53), .B2(n432), .A(n254), .ZN(n444) );
  INV_X1 U13 ( .A(n450), .ZN(n53) );
  OAI21_X1 U14 ( .B1(n423), .B2(n399), .A(n254), .ZN(n418) );
  OAI21_X1 U15 ( .B1(n58), .B2(n371), .A(n254), .ZN(n472) );
  OAI21_X1 U16 ( .B1(n458), .B2(n424), .A(n254), .ZN(n453) );
  NOR2_X1 U17 ( .A1(n66), .A2(n54), .ZN(n450) );
  NAND2_X1 U18 ( .A1(n254), .A2(n275), .ZN(n269) );
  NAND4_X1 U19 ( .A1(n43), .A2(n256), .A3(n276), .A4(n277), .ZN(n275) );
  NOR2_X1 U20 ( .A1(n59), .A2(n65), .ZN(n468) );
  INV_X1 U21 ( .A(n402), .ZN(n21) );
  INV_X1 U22 ( .A(n384), .ZN(n25) );
  INV_X1 U23 ( .A(n261), .ZN(n34) );
  INV_X1 U24 ( .A(n427), .ZN(n9) );
  INV_X1 U25 ( .A(n436), .ZN(n7) );
  INV_X1 U26 ( .A(n375), .ZN(n27) );
  INV_X1 U27 ( .A(n366), .ZN(n29) );
  INV_X1 U28 ( .A(n399), .ZN(n39) );
  INV_X1 U29 ( .A(n410), .ZN(n19) );
  INV_X1 U30 ( .A(n247), .ZN(n36) );
  INV_X1 U31 ( .A(n461), .ZN(n13) );
  INV_X1 U32 ( .A(n392), .ZN(n23) );
  INV_X1 U33 ( .A(n458), .ZN(n38) );
  INV_X1 U34 ( .A(n424), .ZN(n42) );
  INV_X1 U35 ( .A(n423), .ZN(n45) );
  INV_X1 U36 ( .A(n297), .ZN(n43) );
  INV_X1 U37 ( .A(n253), .ZN(n40) );
  NOR4_X1 U38 ( .A1(n286), .A2(n479), .A3(n56), .A4(N288), .ZN(n256) );
  NAND4_X1 U39 ( .A1(n46), .A2(n329), .A3(n257), .A4(n477), .ZN(n254) );
  INV_X1 U40 ( .A(n479), .ZN(n46) );
  NOR2_X1 U41 ( .A1(n297), .A2(n40), .ZN(n477) );
  OAI21_X1 U42 ( .B1(n432), .B2(n433), .A(n254), .ZN(n427) );
  NAND2_X1 U43 ( .A1(n231), .A2(n230), .ZN(n433) );
  OAI21_X1 U44 ( .B1(n432), .B2(n441), .A(n254), .ZN(n436) );
  NAND2_X1 U45 ( .A1(n231), .A2(n229), .ZN(n441) );
  OAI21_X1 U46 ( .B1(n371), .B2(n381), .A(n254), .ZN(n375) );
  NAND2_X1 U47 ( .A1(n313), .A2(n237), .ZN(n381) );
  OAI21_X1 U48 ( .B1(n371), .B2(n372), .A(n254), .ZN(n366) );
  NAND2_X1 U49 ( .A1(n238), .A2(n234), .ZN(n372) );
  NAND2_X1 U50 ( .A1(n254), .A2(n415), .ZN(n410) );
  NAND4_X1 U51 ( .A1(n42), .A2(n45), .A3(n243), .A4(n232), .ZN(n415) );
  NAND2_X1 U52 ( .A1(n254), .A2(n255), .ZN(n247) );
  NAND2_X1 U53 ( .A1(n254), .A2(n467), .ZN(n461) );
  NAND4_X1 U54 ( .A1(n449), .A2(n37), .A3(n468), .A4(n234), .ZN(n467) );
  NAND2_X1 U55 ( .A1(n254), .A2(n398), .ZN(n392) );
  OR3_X1 U56 ( .A1(n294), .A2(n287), .A3(n399), .ZN(n398) );
  NAND4_X1 U57 ( .A1(n449), .A2(n277), .A3(n38), .A4(n232), .ZN(n432) );
  NAND2_X1 U58 ( .A1(n254), .A2(n389), .ZN(n384) );
  INV_X1 U59 ( .A(n294), .ZN(n51) );
  NAND2_X1 U60 ( .A1(n254), .A2(n266), .ZN(n261) );
  NAND4_X1 U61 ( .A1(n449), .A2(n277), .A3(n450), .A4(n231), .ZN(n424) );
  AND3_X1 U62 ( .A1(n256), .A2(n244), .A3(n43), .ZN(n449) );
  NAND2_X1 U63 ( .A1(n243), .A2(n241), .ZN(n294) );
  INV_X1 U64 ( .A(n362), .ZN(n30) );
  AND3_X1 U65 ( .A1(n277), .A2(n244), .A3(n276), .ZN(n257) );
  NAND2_X1 U66 ( .A1(n236), .A2(n235), .ZN(n297) );
  NAND2_X1 U67 ( .A1(n254), .A2(n407), .ZN(n402) );
  NAND4_X1 U68 ( .A1(n39), .A2(n243), .A3(n240), .A4(n239), .ZN(n407) );
  NAND2_X1 U69 ( .A1(n329), .A2(n227), .ZN(N288) );
  INV_X1 U70 ( .A(n237), .ZN(n65) );
  INV_X1 U71 ( .A(n230), .ZN(n66) );
  NAND2_X1 U72 ( .A1(n336), .A2(n285), .ZN(n307) );
  INV_X1 U73 ( .A(n233), .ZN(n67) );
  INV_X1 U74 ( .A(n238), .ZN(n59) );
  NAND2_X1 U75 ( .A1(n228), .A2(n285), .ZN(N286) );
  INV_X1 U76 ( .A(n229), .ZN(n54) );
  INV_X1 U77 ( .A(n291), .ZN(n56) );
  AND4_X1 U78 ( .A1(n38), .A2(n450), .A3(n232), .A4(n231), .ZN(n276) );
  INV_X1 U79 ( .A(n234), .ZN(n52) );
  INV_X1 U80 ( .A(n227), .ZN(n41) );
  INV_X1 U81 ( .A(n231), .ZN(n60) );
  INV_X1 U82 ( .A(n329), .ZN(n49) );
  OAI221_X1 U83 ( .B1(n340), .B2(n238), .C1(n74), .C2(n242), .A(n341), .ZN(
        n330) );
  INV_X1 U84 ( .A(n311), .ZN(n74) );
  AOI222_X1 U85 ( .A1(n68), .A2(n65), .B1(n63), .B2(n299), .C1(n41), .C2(n303), 
        .ZN(n341) );
  INV_X1 U86 ( .A(n244), .ZN(n63) );
  OAI221_X1 U87 ( .B1(n47), .B2(n75), .C1(n73), .C2(n235), .A(n326), .ZN(n317)
         );
  INV_X1 U88 ( .A(n304), .ZN(n73) );
  INV_X1 U89 ( .A(n307), .ZN(n47) );
  NOR2_X1 U90 ( .A1(n49), .A2(n327), .ZN(n326) );
  OAI21_X1 U91 ( .B1(n312), .B2(n228), .A(n254), .ZN(n362) );
  NAND2_X1 U92 ( .A1(n482), .A2(n488), .ZN(n231) );
  OAI21_X1 U93 ( .B1(n64), .B2(n346), .A(n306), .ZN(n286) );
  INV_X1 U94 ( .A(n487), .ZN(n64) );
  NAND2_X1 U95 ( .A1(n488), .A2(n480), .ZN(n242) );
  NAND2_X1 U96 ( .A1(n487), .A2(n358), .ZN(n228) );
  OAI22_X1 U97 ( .A1(n291), .A2(n72), .B1(n229), .B2(n292), .ZN(n290) );
  AOI21_X1 U98 ( .B1(n59), .B2(n340), .A(n52), .ZN(n313) );
  NAND2_X1 U99 ( .A1(n478), .A2(n69), .ZN(n234) );
  NAND2_X1 U100 ( .A1(n357), .A2(n488), .ZN(n232) );
  NAND2_X1 U101 ( .A1(n488), .A2(n483), .ZN(n229) );
  OAI21_X1 U102 ( .B1(n240), .B2(n339), .A(n239), .ZN(n287) );
  NAND2_X1 U103 ( .A1(n481), .A2(n488), .ZN(n243) );
  NAND2_X1 U104 ( .A1(n486), .A2(n488), .ZN(n240) );
  INV_X1 U105 ( .A(n346), .ZN(n69) );
  NAND2_X1 U106 ( .A1(n488), .A2(n487), .ZN(n230) );
  INV_X1 U107 ( .A(n350), .ZN(n57) );
  NAND2_X1 U108 ( .A1(n69), .A2(n480), .ZN(n235) );
  NAND2_X1 U109 ( .A1(n478), .A2(n488), .ZN(n241) );
  NAND2_X1 U110 ( .A1(n485), .A2(n357), .ZN(n239) );
  NAND2_X1 U111 ( .A1(n482), .A2(n358), .ZN(n244) );
  NAND2_X1 U112 ( .A1(n358), .A2(n480), .ZN(n227) );
  NAND2_X1 U113 ( .A1(n485), .A2(n487), .ZN(n237) );
  OAI211_X1 U114 ( .C1(n312), .C2(n228), .A(n313), .B(n314), .ZN(n309) );
  NAND2_X1 U115 ( .A1(n485), .A2(n482), .ZN(n238) );
  NAND2_X1 U116 ( .A1(n69), .A2(n482), .ZN(n285) );
  NAND2_X1 U117 ( .A1(n69), .A2(n357), .ZN(n329) );
  NAND2_X1 U118 ( .A1(n69), .A2(n486), .ZN(n233) );
  INV_X1 U119 ( .A(n312), .ZN(n72) );
  NAND2_X1 U120 ( .A1(n481), .A2(n69), .ZN(n236) );
  NAND2_X1 U121 ( .A1(n483), .A2(n358), .ZN(n291) );
  NAND2_X1 U122 ( .A1(n478), .A2(n358), .ZN(n338) );
  NAND2_X1 U123 ( .A1(n481), .A2(n358), .ZN(n306) );
  NAND2_X1 U124 ( .A1(n357), .A2(n358), .ZN(n336) );
  INV_X1 U125 ( .A(n358), .ZN(n70) );
  OAI221_X1 U126 ( .B1(n2), .B2(n337), .C1(n71), .C2(n240), .A(n338), .ZN(n293) );
  INV_X1 U127 ( .A(n339), .ZN(n71) );
  INV_X1 U128 ( .A(n303), .ZN(n2) );
  NAND2_X1 U129 ( .A1(n486), .A2(n358), .ZN(n337) );
  INV_X1 U130 ( .A(n469), .ZN(n37) );
  OAI21_X1 U131 ( .B1(n233), .B2(n296), .A(n276), .ZN(n469) );
  INV_X1 U132 ( .A(n295), .ZN(n44) );
  AOI211_X1 U133 ( .C1(n296), .C2(n67), .A(n297), .B(n298), .ZN(n295) );
  OAI21_X1 U134 ( .B1(n299), .B2(n244), .A(n234), .ZN(n298) );
  NAND4_X1 U135 ( .A1(n336), .A2(n62), .A3(n338), .A4(n484), .ZN(n479) );
  AND2_X1 U136 ( .A1(n337), .A2(n283), .ZN(n484) );
  INV_X1 U137 ( .A(N286), .ZN(n62) );
  OAI22_X1 U138 ( .A1(n242), .A2(n311), .B1(n68), .B2(n237), .ZN(n310) );
  NOR2_X1 U139 ( .A1(n303), .A2(n227), .ZN(N53) );
  INV_X1 U140 ( .A(n279), .ZN(n68) );
  AOI211_X1 U141 ( .C1(n147), .C2(n148), .A(n145), .B(n70), .ZN(n350) );
  NOR3_X1 U142 ( .A1(state[0]), .A2(state[2]), .A3(n147), .ZN(n487) );
  NOR3_X1 U143 ( .A1(n148), .A2(state[2]), .A3(n147), .ZN(n483) );
  AOI211_X1 U144 ( .C1(n72), .C2(n56), .A(n293), .B(n48), .ZN(n314) );
  INV_X1 U145 ( .A(n334), .ZN(n48) );
  AOI222_X1 U146 ( .A1(n67), .A2(n296), .B1(start), .B2(n307), .C1(n54), .C2(
        n292), .ZN(n334) );
  NOR2_X1 U147 ( .A1(n218), .A2(n359), .ZN(n312) );
  AOI21_X1 U148 ( .B1(n300), .B2(n301), .A(reset), .ZN(N49) );
  NOR4_X1 U149 ( .A1(n302), .A2(n50), .A3(N53), .A4(n66), .ZN(n301) );
  AOI211_X1 U150 ( .C1(n308), .C2(n60), .A(n309), .B(n310), .ZN(n300) );
  INV_X1 U151 ( .A(n241), .ZN(n50) );
  NAND2_X1 U152 ( .A1(addr_y[3]), .A2(n342), .ZN(n303) );
  NOR3_X1 U153 ( .A1(n168), .A2(n169), .A3(n167), .ZN(n462) );
  NOR3_X1 U154 ( .A1(n202), .A2(n203), .A3(n201), .ZN(n393) );
  NOR3_X1 U155 ( .A1(n184), .A2(n185), .A3(n183), .ZN(n335) );
  NOR3_X1 U156 ( .A1(n224), .A2(n225), .A3(n223), .ZN(n342) );
  NOR2_X1 U157 ( .A1(n148), .A2(n345), .ZN(n480) );
  AOI22_X1 U158 ( .A1(n225), .A2(n350), .B1(n57), .B2(n355), .ZN(n353) );
  NOR2_X1 U159 ( .A1(n345), .A2(state[0]), .ZN(n481) );
  AOI22_X1 U160 ( .A1(n483), .A2(state[3]), .B1(state[2]), .B2(n485), .ZN(n283) );
  AOI21_X1 U161 ( .B1(n194), .B2(n410), .A(n40), .ZN(n413) );
  AOI21_X1 U162 ( .B1(n152), .B2(n269), .A(n40), .ZN(n273) );
  AOI21_X1 U163 ( .B1(n161), .B2(n247), .A(n40), .ZN(n251) );
  AOI21_X1 U164 ( .B1(n169), .B2(n461), .A(n40), .ZN(n465) );
  AOI21_X1 U165 ( .B1(n203), .B2(n392), .A(n40), .ZN(n396) );
  AOI21_X1 U166 ( .B1(n198), .B2(n402), .A(n40), .ZN(n405) );
  AOI21_X1 U167 ( .B1(n185), .B2(n427), .A(n40), .ZN(n430) );
  AOI21_X1 U168 ( .B1(n165), .B2(n472), .A(n40), .ZN(n475) );
  AOI21_X1 U169 ( .B1(n207), .B2(n384), .A(n40), .ZN(n387) );
  AOI21_X1 U170 ( .B1(n173), .B2(n453), .A(n40), .ZN(n456) );
  AOI21_X1 U171 ( .B1(n177), .B2(n444), .A(n40), .ZN(n447) );
  AOI21_X1 U172 ( .B1(n181), .B2(n436), .A(n40), .ZN(n439) );
  AOI21_X1 U173 ( .B1(n189), .B2(n418), .A(n40), .ZN(n421) );
  AOI21_X1 U174 ( .B1(n156), .B2(n261), .A(n40), .ZN(n264) );
  AOI21_X1 U175 ( .B1(n211), .B2(n375), .A(n40), .ZN(n379) );
  AOI21_X1 U176 ( .B1(n216), .B2(n366), .A(n40), .ZN(n369) );
  NOR3_X1 U177 ( .A1(n210), .A2(n211), .A3(n209), .ZN(n376) );
  AOI21_X1 U178 ( .B1(n288), .B2(n289), .A(reset), .ZN(N50) );
  NOR3_X1 U179 ( .A1(n293), .A2(n44), .A3(n294), .ZN(n288) );
  NOR3_X1 U180 ( .A1(n290), .A2(N288), .A3(n3), .ZN(n289) );
  INV_X1 U181 ( .A(n242), .ZN(n3) );
  OAI21_X1 U182 ( .B1(addr_y[1]), .B2(n57), .A(n353), .ZN(n351) );
  OAI21_X1 U183 ( .B1(addr_a12[1]), .B2(n21), .A(n405), .ZN(n403) );
  OAI21_X1 U184 ( .B1(addr_a9[1]), .B2(n9), .A(n430), .ZN(n428) );
  OAI21_X1 U185 ( .B1(addr_a11[1]), .B2(n19), .A(n413), .ZN(n411) );
  OAI21_X1 U186 ( .B1(addr_a4[1]), .B2(n11), .A(n475), .ZN(n473) );
  OAI21_X1 U187 ( .B1(addr_a14[1]), .B2(n25), .A(n387), .ZN(n385) );
  OAI21_X1 U188 ( .B1(addr_a6[1]), .B2(n15), .A(n456), .ZN(n454) );
  OAI21_X1 U189 ( .B1(addr_a7[1]), .B2(n5), .A(n447), .ZN(n445) );
  OAI21_X1 U190 ( .B1(addr_a8[1]), .B2(n7), .A(n439), .ZN(n437) );
  OAI21_X1 U191 ( .B1(addr_a1[1]), .B2(n32), .A(n273), .ZN(n271) );
  OAI21_X1 U192 ( .B1(addr_a5[1]), .B2(n13), .A(n465), .ZN(n463) );
  OAI21_X1 U193 ( .B1(addr_a13[1]), .B2(n23), .A(n396), .ZN(n394) );
  OAI21_X1 U194 ( .B1(addr_a10[1]), .B2(n17), .A(n421), .ZN(n419) );
  OAI21_X1 U195 ( .B1(addr_a2[1]), .B2(n34), .A(n264), .ZN(n262) );
  OAI21_X1 U196 ( .B1(addr_a3[1]), .B2(n36), .A(n251), .ZN(n249) );
  OAI21_X1 U197 ( .B1(addr_a15[1]), .B2(n27), .A(n379), .ZN(n377) );
  OAI21_X1 U198 ( .B1(addr_a16[1]), .B2(n29), .A(n369), .ZN(n367) );
  OAI22_X1 U199 ( .A1(n30), .A2(n218), .B1(n30), .B2(n359), .ZN(N271) );
  OAI22_X1 U200 ( .A1(addr_a9[0]), .A2(n9), .B1(n253), .B2(n185), .ZN(N165) );
  OAI22_X1 U201 ( .A1(addr_a11[0]), .A2(n19), .B1(n253), .B2(n194), .ZN(N191)
         );
  OAI22_X1 U202 ( .A1(addr_a7[0]), .A2(n5), .B1(n253), .B2(n177), .ZN(N139) );
  OAI22_X1 U203 ( .A1(addr_a8[0]), .A2(n7), .B1(n253), .B2(n181), .ZN(N152) );
  OAI22_X1 U204 ( .A1(addr_a1[0]), .A2(n32), .B1(n253), .B2(n152), .ZN(N61) );
  OAI22_X1 U205 ( .A1(addr_a3[0]), .A2(n36), .B1(n253), .B2(n161), .ZN(N87) );
  OAI22_X1 U206 ( .A1(addr_a5[0]), .A2(n13), .B1(n253), .B2(n169), .ZN(N113)
         );
  OAI22_X1 U207 ( .A1(addr_a13[0]), .A2(n23), .B1(n253), .B2(n203), .ZN(N217)
         );
  OAI22_X1 U208 ( .A1(addr_a15[0]), .A2(n27), .B1(n253), .B2(n211), .ZN(N243)
         );
  OAI22_X1 U209 ( .A1(addr_a16[0]), .A2(n29), .B1(n253), .B2(n216), .ZN(N256)
         );
  OAI22_X1 U210 ( .A1(addr_a12[0]), .A2(n21), .B1(n253), .B2(n198), .ZN(N204)
         );
  OAI22_X1 U211 ( .A1(addr_a4[0]), .A2(n11), .B1(n253), .B2(n165), .ZN(N100)
         );
  OAI22_X1 U212 ( .A1(addr_a14[0]), .A2(n25), .B1(n253), .B2(n207), .ZN(N230)
         );
  OAI22_X1 U213 ( .A1(addr_a6[0]), .A2(n15), .B1(n253), .B2(n173), .ZN(N126)
         );
  OAI22_X1 U214 ( .A1(addr_a10[0]), .A2(n17), .B1(n253), .B2(n189), .ZN(N178)
         );
  OAI22_X1 U215 ( .A1(addr_a2[0]), .A2(n34), .B1(n253), .B2(n156), .ZN(N74) );
  AND2_X1 U216 ( .A1(n490), .A2(n148), .ZN(n357) );
  NAND2_X1 U217 ( .A1(addr_a5[3]), .A2(n462), .ZN(n296) );
  NOR2_X1 U218 ( .A1(reset), .A2(n242), .ZN(wr_en_a11) );
  NOR2_X1 U219 ( .A1(reset), .A2(n228), .ZN(wr_en_x) );
  NOR2_X1 U220 ( .A1(reset), .A2(n231), .ZN(wr_en_a7) );
  OAI21_X1 U221 ( .B1(n470), .B2(n162), .A(n471), .ZN(N103) );
  OR3_X1 U222 ( .A1(n11), .A2(addr_a4[3]), .A3(n322), .ZN(n471) );
  AOI21_X1 U223 ( .B1(n472), .B2(n163), .A(n473), .ZN(n470) );
  NOR2_X1 U224 ( .A1(reset), .A2(n229), .ZN(wr_en_a9) );
  OAI21_X1 U225 ( .B1(n228), .B2(n72), .A(n284), .ZN(n282) );
  OR4_X1 U226 ( .A1(n285), .A2(loadMatrix), .A3(loadVector), .A4(start), .ZN(
        n284) );
  OAI211_X1 U227 ( .C1(loadVector), .C2(n285), .A(n314), .B(n61), .ZN(n331) );
  INV_X1 U228 ( .A(n332), .ZN(n61) );
  OAI22_X1 U229 ( .A1(n231), .A2(n308), .B1(n72), .B2(n228), .ZN(n332) );
  NOR2_X1 U230 ( .A1(reset), .A2(n232), .ZN(wr_en_a6) );
  NOR2_X1 U231 ( .A1(reset), .A2(n243), .ZN(wr_en_a10) );
  NOR2_X1 U232 ( .A1(reset), .A2(n240), .ZN(wr_en_a13) );
  NOR2_X1 U233 ( .A1(reset), .A2(n230), .ZN(wr_en_a8) );
  NAND2_X1 U234 ( .A1(addr_a9[3]), .A2(n335), .ZN(n292) );
  NOR2_X1 U235 ( .A1(reset), .A2(n241), .ZN(wr_en_a12) );
  NAND2_X1 U236 ( .A1(addr_a13[3]), .A2(n393), .ZN(n339) );
  NOR2_X1 U237 ( .A1(reset), .A2(n227), .ZN(wr_en_y) );
  NOR2_X1 U238 ( .A1(reset), .A2(n237), .ZN(wr_en_a16) );
  NOR2_X1 U239 ( .A1(reset), .A2(n234), .ZN(wr_en_a4) );
  NOR2_X1 U240 ( .A1(reset), .A2(n244), .ZN(wr_en_a1) );
  NOR2_X1 U241 ( .A1(reset), .A2(n235), .ZN(wr_en_a3) );
  NOR2_X1 U242 ( .A1(reset), .A2(n239), .ZN(wr_en_a14) );
  NOR2_X1 U243 ( .A1(reset), .A2(n236), .ZN(wr_en_a2) );
  NOR2_X1 U244 ( .A1(reset), .A2(n233), .ZN(wr_en_a5) );
  NOR2_X1 U245 ( .A1(reset), .A2(n238), .ZN(wr_en_a15) );
  AND2_X1 U246 ( .A1(n490), .A2(state[0]), .ZN(n482) );
  AND2_X1 U247 ( .A1(state[3]), .A2(state[4]), .ZN(n485) );
  NAND2_X1 U248 ( .A1(state[3]), .A2(n140), .ZN(n346) );
  NAND2_X1 U249 ( .A1(state[2]), .A2(n147), .ZN(n345) );
  NOR2_X1 U250 ( .A1(n30), .A2(addr_x[0]), .ZN(N268) );
  NOR2_X1 U251 ( .A1(n147), .A2(n145), .ZN(n489) );
  NOR2_X1 U252 ( .A1(state[2]), .A2(state[1]), .ZN(n490) );
  AOI21_X1 U253 ( .B1(n315), .B2(n316), .A(reset), .ZN(N48) );
  NOR4_X1 U254 ( .A1(n317), .A2(n318), .A3(n319), .A4(n320), .ZN(n316) );
  NOR2_X1 U255 ( .A1(n330), .A2(n331), .ZN(n315) );
  AND3_X1 U256 ( .A1(addr_a8[3]), .A2(n66), .A3(n323), .ZN(n319) );
  AOI21_X1 U257 ( .B1(n280), .B2(n281), .A(reset), .ZN(N51) );
  NOR3_X1 U258 ( .A1(n44), .A2(n286), .A3(n287), .ZN(n280) );
  NOR3_X1 U259 ( .A1(n282), .A2(n58), .A3(n55), .ZN(n281) );
  INV_X1 U260 ( .A(n283), .ZN(n55) );
  AOI21_X1 U261 ( .B1(n278), .B2(n37), .A(reset), .ZN(N52) );
  AOI21_X1 U262 ( .B1(n65), .B2(n279), .A(n59), .ZN(n278) );
  AND2_X1 U263 ( .A1(n489), .A2(state[0]), .ZN(n486) );
  AND2_X1 U264 ( .A1(n489), .A2(n148), .ZN(n478) );
  OAI21_X1 U265 ( .B1(n405), .B2(n197), .A(n406), .ZN(N205) );
  OAI21_X1 U266 ( .B1(n430), .B2(n184), .A(n431), .ZN(N166) );
  OAI21_X1 U267 ( .B1(n475), .B2(n164), .A(n476), .ZN(N101) );
  OAI21_X1 U268 ( .B1(n413), .B2(n193), .A(n414), .ZN(N192) );
  OAI21_X1 U269 ( .B1(n387), .B2(n206), .A(n388), .ZN(N231) );
  OAI21_X1 U270 ( .B1(n456), .B2(n172), .A(n457), .ZN(N127) );
  OAI21_X1 U271 ( .B1(n447), .B2(n176), .A(n448), .ZN(N140) );
  OAI21_X1 U272 ( .B1(n439), .B2(n180), .A(n440), .ZN(N153) );
  OAI21_X1 U273 ( .B1(n421), .B2(n188), .A(n422), .ZN(N179) );
  OAI21_X1 U274 ( .B1(n273), .B2(n151), .A(n274), .ZN(N62) );
  OAI21_X1 U275 ( .B1(n264), .B2(n155), .A(n265), .ZN(N75) );
  OAI21_X1 U276 ( .B1(n251), .B2(n160), .A(n252), .ZN(N88) );
  OAI21_X1 U277 ( .B1(n465), .B2(n168), .A(n466), .ZN(N114) );
  OAI21_X1 U278 ( .B1(n396), .B2(n202), .A(n397), .ZN(N218) );
  OAI21_X1 U279 ( .B1(n379), .B2(n210), .A(n380), .ZN(N244) );
  OAI21_X1 U280 ( .B1(n369), .B2(n215), .A(n370), .ZN(N257) );
  OAI21_X1 U281 ( .B1(n353), .B2(n224), .A(n354), .ZN(N281) );
  OAI21_X1 U282 ( .B1(n348), .B2(n222), .A(n349), .ZN(N283) );
  AOI21_X1 U283 ( .B1(n350), .B2(n223), .A(n351), .ZN(n348) );
  OAI21_X1 U284 ( .B1(addr_y[0]), .B2(n57), .A(n356), .ZN(N280) );
  OAI21_X1 U285 ( .B1(n8), .B2(n183), .A(n429), .ZN(N167) );
  NAND4_X1 U286 ( .A1(addr_a9[1]), .A2(addr_a9[0]), .A3(n427), .A4(n183), .ZN(
        n429) );
  INV_X1 U287 ( .A(n428), .ZN(n8) );
  OAI21_X1 U288 ( .B1(n18), .B2(n192), .A(n412), .ZN(N193) );
  NAND4_X1 U289 ( .A1(addr_a11[1]), .A2(addr_a11[0]), .A3(n410), .A4(n192), 
        .ZN(n412) );
  INV_X1 U290 ( .A(n411), .ZN(n18) );
  OAI21_X1 U291 ( .B1(n4), .B2(n175), .A(n446), .ZN(N141) );
  NAND4_X1 U292 ( .A1(addr_a7[1]), .A2(addr_a7[0]), .A3(n444), .A4(n175), .ZN(
        n446) );
  INV_X1 U293 ( .A(n445), .ZN(n4) );
  OAI21_X1 U294 ( .B1(n6), .B2(n179), .A(n438), .ZN(N154) );
  NAND4_X1 U295 ( .A1(addr_a8[1]), .A2(addr_a8[0]), .A3(n436), .A4(n179), .ZN(
        n438) );
  INV_X1 U296 ( .A(n437), .ZN(n6) );
  OAI21_X1 U297 ( .B1(n31), .B2(n150), .A(n272), .ZN(N63) );
  NAND4_X1 U298 ( .A1(addr_a1[1]), .A2(addr_a1[0]), .A3(n269), .A4(n150), .ZN(
        n272) );
  INV_X1 U299 ( .A(n271), .ZN(n31) );
  OAI21_X1 U300 ( .B1(n35), .B2(n159), .A(n250), .ZN(N89) );
  NAND4_X1 U301 ( .A1(addr_a3[1]), .A2(addr_a3[0]), .A3(n247), .A4(n159), .ZN(
        n250) );
  INV_X1 U302 ( .A(n249), .ZN(n35) );
  OAI21_X1 U303 ( .B1(n12), .B2(n167), .A(n464), .ZN(N115) );
  NAND4_X1 U304 ( .A1(addr_a5[1]), .A2(addr_a5[0]), .A3(n461), .A4(n167), .ZN(
        n464) );
  INV_X1 U305 ( .A(n463), .ZN(n12) );
  OAI21_X1 U306 ( .B1(n22), .B2(n201), .A(n395), .ZN(N219) );
  NAND4_X1 U307 ( .A1(addr_a13[1]), .A2(addr_a13[0]), .A3(n392), .A4(n201), 
        .ZN(n395) );
  INV_X1 U308 ( .A(n394), .ZN(n22) );
  OAI21_X1 U309 ( .B1(n26), .B2(n209), .A(n378), .ZN(N245) );
  NAND4_X1 U310 ( .A1(addr_a15[1]), .A2(addr_a15[0]), .A3(n375), .A4(n209), 
        .ZN(n378) );
  INV_X1 U311 ( .A(n377), .ZN(n26) );
  OAI21_X1 U312 ( .B1(n28), .B2(n214), .A(n368), .ZN(N258) );
  NAND4_X1 U313 ( .A1(addr_a16[1]), .A2(addr_a16[0]), .A3(n366), .A4(n214), 
        .ZN(n368) );
  INV_X1 U314 ( .A(n367), .ZN(n28) );
  OAI21_X1 U315 ( .B1(n1), .B2(n223), .A(n352), .ZN(N282) );
  NAND4_X1 U316 ( .A1(n350), .A2(addr_y[1]), .A3(addr_y[0]), .A4(n223), .ZN(
        n352) );
  INV_X1 U317 ( .A(n351), .ZN(n1) );
  OAI21_X1 U318 ( .B1(n20), .B2(n196), .A(n404), .ZN(N206) );
  NAND4_X1 U319 ( .A1(addr_a12[1]), .A2(addr_a12[0]), .A3(n402), .A4(n196), 
        .ZN(n404) );
  INV_X1 U320 ( .A(n403), .ZN(n20) );
  OAI21_X1 U321 ( .B1(n10), .B2(n163), .A(n474), .ZN(N102) );
  NAND4_X1 U322 ( .A1(addr_a4[1]), .A2(addr_a4[0]), .A3(n472), .A4(n163), .ZN(
        n474) );
  INV_X1 U323 ( .A(n473), .ZN(n10) );
  OAI21_X1 U324 ( .B1(n24), .B2(n205), .A(n386), .ZN(N232) );
  NAND4_X1 U325 ( .A1(addr_a14[1]), .A2(addr_a14[0]), .A3(n384), .A4(n205), 
        .ZN(n386) );
  INV_X1 U326 ( .A(n385), .ZN(n24) );
  OAI21_X1 U327 ( .B1(n14), .B2(n171), .A(n455), .ZN(N128) );
  NAND4_X1 U328 ( .A1(addr_a6[1]), .A2(addr_a6[0]), .A3(n453), .A4(n171), .ZN(
        n455) );
  INV_X1 U329 ( .A(n454), .ZN(n14) );
  OAI21_X1 U330 ( .B1(n16), .B2(n187), .A(n420), .ZN(N180) );
  NAND4_X1 U331 ( .A1(addr_a10[1]), .A2(addr_a10[0]), .A3(n418), .A4(n187), 
        .ZN(n420) );
  INV_X1 U332 ( .A(n419), .ZN(n16) );
  OAI21_X1 U333 ( .B1(n33), .B2(n154), .A(n263), .ZN(N76) );
  NAND4_X1 U334 ( .A1(addr_a2[1]), .A2(addr_a2[0]), .A3(n261), .A4(n154), .ZN(
        n263) );
  INV_X1 U335 ( .A(n262), .ZN(n33) );
  OAI21_X1 U336 ( .B1(n425), .B2(n182), .A(n426), .ZN(N168) );
  AOI21_X1 U337 ( .B1(n427), .B2(n183), .A(n428), .ZN(n425) );
  OAI21_X1 U338 ( .B1(n434), .B2(n178), .A(n435), .ZN(N155) );
  AOI21_X1 U339 ( .B1(n436), .B2(n179), .A(n437), .ZN(n434) );
  OAI21_X1 U340 ( .B1(n373), .B2(n208), .A(n374), .ZN(N246) );
  AOI21_X1 U341 ( .B1(n375), .B2(n209), .A(n377), .ZN(n373) );
  OAI21_X1 U342 ( .B1(n364), .B2(n213), .A(n365), .ZN(N259) );
  AOI21_X1 U343 ( .B1(n366), .B2(n214), .A(n367), .ZN(n364) );
  OAI21_X1 U344 ( .B1(n442), .B2(n174), .A(n443), .ZN(N142) );
  AOI21_X1 U345 ( .B1(n444), .B2(n175), .A(n445), .ZN(n442) );
  OAI21_X1 U346 ( .B1(n451), .B2(n170), .A(n452), .ZN(N129) );
  OR3_X1 U347 ( .A1(n15), .A2(addr_a6[3]), .A3(n321), .ZN(n452) );
  AOI21_X1 U348 ( .B1(n453), .B2(n171), .A(n454), .ZN(n451) );
  OAI21_X1 U349 ( .B1(n416), .B2(n186), .A(n417), .ZN(N181) );
  OR3_X1 U350 ( .A1(n17), .A2(addr_a10[3]), .A3(n325), .ZN(n417) );
  AOI21_X1 U351 ( .B1(n418), .B2(n187), .A(n419), .ZN(n416) );
  OAI21_X1 U352 ( .B1(n360), .B2(n219), .A(n361), .ZN(N270) );
  NAND4_X1 U353 ( .A1(addr_x[1]), .A2(addr_x[0]), .A3(n362), .A4(n219), .ZN(
        n361) );
  AOI21_X1 U354 ( .B1(n362), .B2(n220), .A(N268), .ZN(n360) );
  OAI21_X1 U355 ( .B1(n408), .B2(n191), .A(n409), .ZN(N194) );
  AOI21_X1 U356 ( .B1(n410), .B2(n192), .A(n411), .ZN(n408) );
  OAI21_X1 U357 ( .B1(n267), .B2(n149), .A(n268), .ZN(N64) );
  AOI21_X1 U358 ( .B1(n269), .B2(n150), .A(n271), .ZN(n267) );
  OAI21_X1 U359 ( .B1(n245), .B2(n157), .A(n246), .ZN(N90) );
  AOI21_X1 U360 ( .B1(n247), .B2(n159), .A(n249), .ZN(n245) );
  OAI21_X1 U361 ( .B1(n459), .B2(n166), .A(n460), .ZN(N116) );
  AOI21_X1 U362 ( .B1(n461), .B2(n167), .A(n463), .ZN(n459) );
  OAI21_X1 U363 ( .B1(n390), .B2(n199), .A(n391), .ZN(N220) );
  AOI21_X1 U364 ( .B1(n392), .B2(n201), .A(n394), .ZN(n390) );
  AND2_X1 U365 ( .A1(addr_a15[3]), .A2(n376), .ZN(n340) );
  OAI21_X1 U366 ( .B1(n400), .B2(n195), .A(n401), .ZN(N207) );
  OR3_X1 U367 ( .A1(n21), .A2(addr_a12[3]), .A3(n324), .ZN(n401) );
  AOI21_X1 U368 ( .B1(n402), .B2(n196), .A(n403), .ZN(n400) );
  OAI21_X1 U369 ( .B1(n382), .B2(n204), .A(n383), .ZN(N233) );
  OR3_X1 U370 ( .A1(n25), .A2(addr_a14[3]), .A3(n328), .ZN(n383) );
  AOI21_X1 U371 ( .B1(n384), .B2(n205), .A(n385), .ZN(n382) );
  OAI21_X1 U372 ( .B1(n258), .B2(n153), .A(n259), .ZN(N77) );
  OR3_X1 U373 ( .A1(n34), .A2(addr_a2[3]), .A3(n260), .ZN(n259) );
  AOI21_X1 U374 ( .B1(n261), .B2(n154), .A(n262), .ZN(n258) );
  NOR2_X1 U375 ( .A1(n30), .A2(n363), .ZN(N269) );
  XNOR2_X1 U376 ( .A(addr_x[0]), .B(addr_x[1]), .ZN(n363) );
  NOR3_X1 U377 ( .A1(n151), .A2(n152), .A3(n150), .ZN(n270) );
  NOR3_X1 U378 ( .A1(n215), .A2(n216), .A3(n214), .ZN(n343) );
  NOR3_X1 U379 ( .A1(n193), .A2(n194), .A3(n192), .ZN(n344) );
  NOR3_X1 U380 ( .A1(n160), .A2(n161), .A3(n159), .ZN(n248) );
  NOR3_X1 U381 ( .A1(n176), .A2(n177), .A3(n175), .ZN(n333) );
  NOR3_X1 U382 ( .A1(n180), .A2(n181), .A3(n179), .ZN(n323) );
  OAI22_X1 U383 ( .A1(n345), .A2(n70), .B1(n346), .B2(n347), .ZN(N287) );
  NAND2_X1 U384 ( .A1(n148), .A2(n145), .ZN(n347) );
  OAI211_X1 U385 ( .C1(n235), .C2(n304), .A(n305), .B(n306), .ZN(n302) );
  NAND2_X1 U386 ( .A1(addr_a11[3]), .A2(n344), .ZN(n311) );
  NAND2_X1 U387 ( .A1(addr_a3[3]), .A2(n248), .ZN(n304) );
  NAND2_X1 U388 ( .A1(addr_a16[3]), .A2(n343), .ZN(n279) );
  NAND2_X1 U389 ( .A1(addr_a1[3]), .A2(n270), .ZN(n299) );
  AND2_X1 U390 ( .A1(addr_a7[3]), .A2(n333), .ZN(n308) );
  NAND2_X1 U391 ( .A1(n357), .A2(n140), .ZN(n355) );
  INV_X1 U392 ( .A(loadMatrix), .ZN(n75) );
  AOI211_X4 U393 ( .C1(n56), .C2(n312), .A(n41), .B(n286), .ZN(n253) );
endmodule


module mvm_16_16_8_1 ( clk, reset, loadMatrix, loadVector, start, done, 
        data_in, data_out );
  input [7:0] data_in;
  output [15:0] data_out;
  input clk, reset, loadMatrix, loadVector, start;
  output done;
  wire   wr_en_x, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6,
         wr_en_a7, wr_en_a8, wr_en_a9, wr_en_a10, wr_en_a11, wr_en_a12,
         wr_en_a13, wr_en_a14, wr_en_a15, wr_en_a16, wr_en_y, clear_acc, clc,
         clc1;
  wire   [3:0] addr_x;
  wire   [3:0] addr_a1;
  wire   [3:0] addr_a2;
  wire   [3:0] addr_a3;
  wire   [3:0] addr_a4;
  wire   [3:0] addr_a5;
  wire   [3:0] addr_a6;
  wire   [3:0] addr_a7;
  wire   [3:0] addr_a8;
  wire   [3:0] addr_a9;
  wire   [3:0] addr_a10;
  wire   [3:0] addr_a11;
  wire   [3:0] addr_a12;
  wire   [3:0] addr_a13;
  wire   [3:0] addr_a14;
  wire   [3:0] addr_a15;
  wire   [3:0] addr_a16;
  wire   [3:0] addr_y;

  datapath d ( .clk(clk), .data_in(data_in), .addr_x(addr_x), .wr_en_x(wr_en_x), .addr_a1(addr_a1), .addr_a2(addr_a2), .addr_a3(addr_a3), .addr_a4(addr_a4), 
        .addr_a5(addr_a5), .addr_a6(addr_a6), .addr_a7(addr_a7), .addr_a8(
        addr_a8), .addr_a9(addr_a9), .addr_a10(addr_a10), .addr_a11(addr_a11), 
        .addr_a12(addr_a12), .addr_a13(addr_a13), .addr_a14(addr_a14), 
        .addr_a15(addr_a15), .addr_a16(addr_a16), .wr_en_a1(wr_en_a1), 
        .wr_en_a2(wr_en_a2), .wr_en_a3(wr_en_a3), .wr_en_a4(wr_en_a4), 
        .wr_en_a5(wr_en_a5), .wr_en_a6(wr_en_a6), .wr_en_a7(wr_en_a7), 
        .wr_en_a8(wr_en_a8), .wr_en_a9(wr_en_a9), .wr_en_a10(wr_en_a10), 
        .wr_en_a11(wr_en_a11), .wr_en_a12(wr_en_a12), .wr_en_a13(wr_en_a13), 
        .wr_en_a14(wr_en_a14), .wr_en_a15(wr_en_a15), .wr_en_a16(wr_en_a16), 
        .addr_y(addr_y), .wr_en_y(wr_en_y), .clear_acc(clear_acc), .clc(clc), 
        .clc1(clc1), .data_out(data_out) );
  ctrlpath c ( .clk(clk), .reset(reset), .start(start), .addr_x(addr_x), 
        .wr_en_x(wr_en_x), .addr_a1(addr_a1), .addr_a2(addr_a2), .addr_a3(
        addr_a3), .addr_a4(addr_a4), .addr_a5(addr_a5), .addr_a6(addr_a6), 
        .addr_a7(addr_a7), .addr_a8(addr_a8), .addr_a9(addr_a9), .addr_a10(
        addr_a10), .addr_a11(addr_a11), .addr_a12(addr_a12), .addr_a13(
        addr_a13), .addr_a14(addr_a14), .addr_a15(addr_a15), .addr_a16(
        addr_a16), .wr_en_a1(wr_en_a1), .wr_en_a2(wr_en_a2), .wr_en_a3(
        wr_en_a3), .wr_en_a4(wr_en_a4), .wr_en_a5(wr_en_a5), .wr_en_a6(
        wr_en_a6), .wr_en_a7(wr_en_a7), .wr_en_a8(wr_en_a8), .wr_en_a9(
        wr_en_a9), .wr_en_a10(wr_en_a10), .wr_en_a11(wr_en_a11), .wr_en_a12(
        wr_en_a12), .wr_en_a13(wr_en_a13), .wr_en_a14(wr_en_a14), .wr_en_a15(
        wr_en_a15), .wr_en_a16(wr_en_a16), .clear_acc(clear_acc), .clc(clc), 
        .clc1(clc1), .addr_y(addr_y), .wr_en_y(wr_en_y), .done(done), 
        .loadMatrix(loadMatrix), .loadVector(loadVector) );
endmodule

