
module memory_WIDTH12_SIZE8_LOGSIZE3_0 ( clk, data_in, data_out, addr, wr_en
 );
  input [11:0] data_in;
  output [11:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] ,
         \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] ,
         \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][11] , \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] ,
         \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] ,
         \mem[5][1] , \mem[5][0] , \mem[4][11] , \mem[4][10] , \mem[4][9] ,
         \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] ,
         \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] ,
         \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] ,
         \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][11] , \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] ,
         \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] ,
         \mem[0][1] , \mem[0][0] , n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \mem_reg[7][11]  ( .D(n217), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n216), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n215), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n214), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n213), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n212), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n211), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n210), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n209), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n208), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n207), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n206), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n205), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n204), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n203), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n202), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n201), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n200), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n199), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n198), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n197), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n196), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n195), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n194), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n193), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n192), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n191), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n190), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n189), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n188), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n187), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n186), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n185), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n184), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n183), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n182), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n181), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n180), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n179), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n178), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n177), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n176), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n175), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n174), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n173), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n172), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n171), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n170), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n169), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n168), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n167), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n166), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n165), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n164), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n163), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n162), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n161), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n160), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n159), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n158), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n157), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n156), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n155), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n154), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n153), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n152), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n151), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n150), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n149), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n148), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n147), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n146), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n145), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n144), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n143), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n142), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n141), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n140), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n139), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n138), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n137), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n136), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n135), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n134), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n133), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n132), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n131), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n130), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n129), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n128), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n127), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n126), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n125), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n124), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n123), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n122), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U212 ( .A1(n282), .A2(n283), .A3(n29), .ZN(n16) );
  NAND3_X1 U213 ( .A1(n29), .A2(n283), .A3(N10), .ZN(n30) );
  NAND3_X1 U214 ( .A1(n29), .A2(n282), .A3(N11), .ZN(n43) );
  NAND3_X1 U215 ( .A1(N10), .A2(n29), .A3(N11), .ZN(n56) );
  NAND3_X1 U216 ( .A1(n282), .A2(n283), .A3(n82), .ZN(n69) );
  NAND3_X1 U217 ( .A1(N10), .A2(n283), .A3(n82), .ZN(n83) );
  NAND3_X1 U218 ( .A1(N11), .A2(n282), .A3(n82), .ZN(n96) );
  NAND3_X1 U219 ( .A1(N11), .A2(N10), .A3(n82), .ZN(n109) );
  SDFF_X1 \data_out_reg[6]  ( .D(n248), .SI(n245), .SE(N12), .CK(clk), .Q(
        data_out[6]) );
  SDFF_X1 \data_out_reg[8]  ( .D(n260), .SI(n257), .SE(N12), .CK(clk), .Q(
        data_out[8]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n242), .SI(n239), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n266), .SI(n263), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[10]  ( .D(n272), .SI(n269), .SE(N12), .CK(clk), .Q(
        data_out[10]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n254), .SI(n251), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n230), .SI(n227), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[4]  ( .D(n236), .SI(n233), .SE(N12), .CK(clk), .Q(
        data_out[4]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n10), .SI(n7), .SE(N12), .CK(clk), .Q(
        data_out[0]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n218), .SI(n13), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n278), .SI(n275), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[2]  ( .D(n224), .SI(n221), .SE(N12), .CK(clk), .Q(
        data_out[2]) );
  BUF_X1 U3 ( .A(n281), .Z(n280) );
  BUF_X1 U4 ( .A(N11), .Z(n279) );
  BUF_X1 U5 ( .A(N10), .Z(n281) );
  NOR2_X1 U6 ( .A1(n284), .A2(N12), .ZN(n29) );
  INV_X1 U7 ( .A(wr_en), .ZN(n284) );
  AND2_X1 U8 ( .A1(N12), .A2(wr_en), .ZN(n82) );
  INV_X1 U9 ( .A(N10), .ZN(n282) );
  INV_X1 U10 ( .A(N11), .ZN(n283) );
  OAI21_X1 U11 ( .B1(n296), .B2(n30), .A(n31), .ZN(n134) );
  NAND2_X1 U12 ( .A1(\mem[1][0] ), .A2(n30), .ZN(n31) );
  OAI21_X1 U13 ( .B1(n295), .B2(n30), .A(n32), .ZN(n135) );
  NAND2_X1 U14 ( .A1(\mem[1][1] ), .A2(n30), .ZN(n32) );
  OAI21_X1 U15 ( .B1(n294), .B2(n30), .A(n33), .ZN(n136) );
  NAND2_X1 U16 ( .A1(\mem[1][2] ), .A2(n30), .ZN(n33) );
  OAI21_X1 U17 ( .B1(n293), .B2(n30), .A(n34), .ZN(n137) );
  NAND2_X1 U18 ( .A1(\mem[1][3] ), .A2(n30), .ZN(n34) );
  OAI21_X1 U19 ( .B1(n292), .B2(n30), .A(n35), .ZN(n138) );
  NAND2_X1 U20 ( .A1(\mem[1][4] ), .A2(n30), .ZN(n35) );
  OAI21_X1 U21 ( .B1(n291), .B2(n30), .A(n36), .ZN(n139) );
  NAND2_X1 U22 ( .A1(\mem[1][5] ), .A2(n30), .ZN(n36) );
  OAI21_X1 U23 ( .B1(n290), .B2(n30), .A(n37), .ZN(n140) );
  NAND2_X1 U24 ( .A1(\mem[1][6] ), .A2(n30), .ZN(n37) );
  OAI21_X1 U25 ( .B1(n289), .B2(n30), .A(n38), .ZN(n141) );
  NAND2_X1 U26 ( .A1(\mem[1][7] ), .A2(n30), .ZN(n38) );
  OAI21_X1 U27 ( .B1(n288), .B2(n30), .A(n39), .ZN(n142) );
  NAND2_X1 U28 ( .A1(\mem[1][8] ), .A2(n30), .ZN(n39) );
  OAI21_X1 U29 ( .B1(n287), .B2(n30), .A(n40), .ZN(n143) );
  NAND2_X1 U30 ( .A1(\mem[1][9] ), .A2(n30), .ZN(n40) );
  OAI21_X1 U31 ( .B1(n286), .B2(n30), .A(n41), .ZN(n144) );
  NAND2_X1 U32 ( .A1(\mem[1][10] ), .A2(n30), .ZN(n41) );
  OAI21_X1 U33 ( .B1(n285), .B2(n30), .A(n42), .ZN(n145) );
  NAND2_X1 U34 ( .A1(\mem[1][11] ), .A2(n30), .ZN(n42) );
  OAI21_X1 U35 ( .B1(n296), .B2(n43), .A(n44), .ZN(n146) );
  NAND2_X1 U36 ( .A1(\mem[2][0] ), .A2(n43), .ZN(n44) );
  OAI21_X1 U37 ( .B1(n295), .B2(n43), .A(n45), .ZN(n147) );
  NAND2_X1 U38 ( .A1(\mem[2][1] ), .A2(n43), .ZN(n45) );
  OAI21_X1 U39 ( .B1(n294), .B2(n43), .A(n46), .ZN(n148) );
  NAND2_X1 U40 ( .A1(\mem[2][2] ), .A2(n43), .ZN(n46) );
  OAI21_X1 U41 ( .B1(n293), .B2(n43), .A(n47), .ZN(n149) );
  NAND2_X1 U42 ( .A1(\mem[2][3] ), .A2(n43), .ZN(n47) );
  OAI21_X1 U43 ( .B1(n292), .B2(n43), .A(n48), .ZN(n150) );
  NAND2_X1 U44 ( .A1(\mem[2][4] ), .A2(n43), .ZN(n48) );
  OAI21_X1 U45 ( .B1(n291), .B2(n43), .A(n49), .ZN(n151) );
  NAND2_X1 U46 ( .A1(\mem[2][5] ), .A2(n43), .ZN(n49) );
  OAI21_X1 U47 ( .B1(n290), .B2(n43), .A(n50), .ZN(n152) );
  NAND2_X1 U48 ( .A1(\mem[2][6] ), .A2(n43), .ZN(n50) );
  OAI21_X1 U49 ( .B1(n289), .B2(n43), .A(n51), .ZN(n153) );
  NAND2_X1 U50 ( .A1(\mem[2][7] ), .A2(n43), .ZN(n51) );
  OAI21_X1 U51 ( .B1(n288), .B2(n43), .A(n52), .ZN(n154) );
  NAND2_X1 U52 ( .A1(\mem[2][8] ), .A2(n43), .ZN(n52) );
  OAI21_X1 U53 ( .B1(n287), .B2(n43), .A(n53), .ZN(n155) );
  NAND2_X1 U54 ( .A1(\mem[2][9] ), .A2(n43), .ZN(n53) );
  OAI21_X1 U55 ( .B1(n286), .B2(n43), .A(n54), .ZN(n156) );
  NAND2_X1 U56 ( .A1(\mem[2][10] ), .A2(n43), .ZN(n54) );
  OAI21_X1 U57 ( .B1(n285), .B2(n43), .A(n55), .ZN(n157) );
  NAND2_X1 U58 ( .A1(\mem[2][11] ), .A2(n43), .ZN(n55) );
  OAI21_X1 U59 ( .B1(n296), .B2(n56), .A(n57), .ZN(n158) );
  NAND2_X1 U60 ( .A1(\mem[3][0] ), .A2(n56), .ZN(n57) );
  OAI21_X1 U61 ( .B1(n295), .B2(n56), .A(n58), .ZN(n159) );
  NAND2_X1 U62 ( .A1(\mem[3][1] ), .A2(n56), .ZN(n58) );
  OAI21_X1 U63 ( .B1(n294), .B2(n56), .A(n59), .ZN(n160) );
  NAND2_X1 U64 ( .A1(\mem[3][2] ), .A2(n56), .ZN(n59) );
  OAI21_X1 U65 ( .B1(n293), .B2(n56), .A(n60), .ZN(n161) );
  NAND2_X1 U66 ( .A1(\mem[3][3] ), .A2(n56), .ZN(n60) );
  OAI21_X1 U67 ( .B1(n292), .B2(n56), .A(n61), .ZN(n162) );
  NAND2_X1 U68 ( .A1(\mem[3][4] ), .A2(n56), .ZN(n61) );
  OAI21_X1 U69 ( .B1(n291), .B2(n56), .A(n62), .ZN(n163) );
  NAND2_X1 U70 ( .A1(\mem[3][5] ), .A2(n56), .ZN(n62) );
  OAI21_X1 U71 ( .B1(n290), .B2(n56), .A(n63), .ZN(n164) );
  NAND2_X1 U72 ( .A1(\mem[3][6] ), .A2(n56), .ZN(n63) );
  OAI21_X1 U73 ( .B1(n289), .B2(n56), .A(n64), .ZN(n165) );
  NAND2_X1 U74 ( .A1(\mem[3][7] ), .A2(n56), .ZN(n64) );
  OAI21_X1 U75 ( .B1(n288), .B2(n56), .A(n65), .ZN(n166) );
  NAND2_X1 U76 ( .A1(\mem[3][8] ), .A2(n56), .ZN(n65) );
  OAI21_X1 U77 ( .B1(n287), .B2(n56), .A(n66), .ZN(n167) );
  NAND2_X1 U78 ( .A1(\mem[3][9] ), .A2(n56), .ZN(n66) );
  OAI21_X1 U79 ( .B1(n286), .B2(n56), .A(n67), .ZN(n168) );
  NAND2_X1 U80 ( .A1(\mem[3][10] ), .A2(n56), .ZN(n67) );
  OAI21_X1 U81 ( .B1(n285), .B2(n56), .A(n68), .ZN(n169) );
  NAND2_X1 U82 ( .A1(\mem[3][11] ), .A2(n56), .ZN(n68) );
  OAI21_X1 U83 ( .B1(n296), .B2(n69), .A(n70), .ZN(n170) );
  NAND2_X1 U84 ( .A1(\mem[4][0] ), .A2(n69), .ZN(n70) );
  OAI21_X1 U85 ( .B1(n295), .B2(n69), .A(n71), .ZN(n171) );
  NAND2_X1 U86 ( .A1(\mem[4][1] ), .A2(n69), .ZN(n71) );
  OAI21_X1 U87 ( .B1(n294), .B2(n69), .A(n72), .ZN(n172) );
  NAND2_X1 U88 ( .A1(\mem[4][2] ), .A2(n69), .ZN(n72) );
  OAI21_X1 U89 ( .B1(n293), .B2(n69), .A(n73), .ZN(n173) );
  NAND2_X1 U90 ( .A1(\mem[4][3] ), .A2(n69), .ZN(n73) );
  OAI21_X1 U91 ( .B1(n292), .B2(n69), .A(n74), .ZN(n174) );
  NAND2_X1 U92 ( .A1(\mem[4][4] ), .A2(n69), .ZN(n74) );
  OAI21_X1 U93 ( .B1(n291), .B2(n69), .A(n75), .ZN(n175) );
  NAND2_X1 U94 ( .A1(\mem[4][5] ), .A2(n69), .ZN(n75) );
  OAI21_X1 U95 ( .B1(n290), .B2(n69), .A(n76), .ZN(n176) );
  NAND2_X1 U96 ( .A1(\mem[4][6] ), .A2(n69), .ZN(n76) );
  OAI21_X1 U97 ( .B1(n289), .B2(n69), .A(n77), .ZN(n177) );
  NAND2_X1 U98 ( .A1(\mem[4][7] ), .A2(n69), .ZN(n77) );
  OAI21_X1 U99 ( .B1(n288), .B2(n69), .A(n78), .ZN(n178) );
  NAND2_X1 U100 ( .A1(\mem[4][8] ), .A2(n69), .ZN(n78) );
  OAI21_X1 U101 ( .B1(n287), .B2(n69), .A(n79), .ZN(n179) );
  NAND2_X1 U102 ( .A1(\mem[4][9] ), .A2(n69), .ZN(n79) );
  OAI21_X1 U103 ( .B1(n286), .B2(n69), .A(n80), .ZN(n180) );
  NAND2_X1 U104 ( .A1(\mem[4][10] ), .A2(n69), .ZN(n80) );
  OAI21_X1 U105 ( .B1(n285), .B2(n69), .A(n81), .ZN(n181) );
  NAND2_X1 U106 ( .A1(\mem[4][11] ), .A2(n69), .ZN(n81) );
  OAI21_X1 U107 ( .B1(n296), .B2(n83), .A(n84), .ZN(n182) );
  NAND2_X1 U108 ( .A1(\mem[5][0] ), .A2(n83), .ZN(n84) );
  OAI21_X1 U109 ( .B1(n295), .B2(n83), .A(n85), .ZN(n183) );
  NAND2_X1 U110 ( .A1(\mem[5][1] ), .A2(n83), .ZN(n85) );
  OAI21_X1 U111 ( .B1(n294), .B2(n83), .A(n86), .ZN(n184) );
  NAND2_X1 U112 ( .A1(\mem[5][2] ), .A2(n83), .ZN(n86) );
  OAI21_X1 U113 ( .B1(n293), .B2(n83), .A(n87), .ZN(n185) );
  NAND2_X1 U114 ( .A1(\mem[5][3] ), .A2(n83), .ZN(n87) );
  OAI21_X1 U115 ( .B1(n292), .B2(n83), .A(n88), .ZN(n186) );
  NAND2_X1 U116 ( .A1(\mem[5][4] ), .A2(n83), .ZN(n88) );
  OAI21_X1 U117 ( .B1(n291), .B2(n83), .A(n89), .ZN(n187) );
  NAND2_X1 U118 ( .A1(\mem[5][5] ), .A2(n83), .ZN(n89) );
  OAI21_X1 U119 ( .B1(n290), .B2(n83), .A(n90), .ZN(n188) );
  NAND2_X1 U120 ( .A1(\mem[5][6] ), .A2(n83), .ZN(n90) );
  OAI21_X1 U121 ( .B1(n289), .B2(n83), .A(n91), .ZN(n189) );
  NAND2_X1 U122 ( .A1(\mem[5][7] ), .A2(n83), .ZN(n91) );
  OAI21_X1 U123 ( .B1(n288), .B2(n83), .A(n92), .ZN(n190) );
  NAND2_X1 U124 ( .A1(\mem[5][8] ), .A2(n83), .ZN(n92) );
  OAI21_X1 U125 ( .B1(n287), .B2(n83), .A(n93), .ZN(n191) );
  NAND2_X1 U126 ( .A1(\mem[5][9] ), .A2(n83), .ZN(n93) );
  OAI21_X1 U127 ( .B1(n286), .B2(n83), .A(n94), .ZN(n192) );
  NAND2_X1 U128 ( .A1(\mem[5][10] ), .A2(n83), .ZN(n94) );
  OAI21_X1 U129 ( .B1(n285), .B2(n83), .A(n95), .ZN(n193) );
  NAND2_X1 U130 ( .A1(\mem[5][11] ), .A2(n83), .ZN(n95) );
  OAI21_X1 U131 ( .B1(n296), .B2(n96), .A(n97), .ZN(n194) );
  NAND2_X1 U132 ( .A1(\mem[6][0] ), .A2(n96), .ZN(n97) );
  OAI21_X1 U133 ( .B1(n295), .B2(n96), .A(n98), .ZN(n195) );
  NAND2_X1 U134 ( .A1(\mem[6][1] ), .A2(n96), .ZN(n98) );
  OAI21_X1 U135 ( .B1(n294), .B2(n96), .A(n99), .ZN(n196) );
  NAND2_X1 U136 ( .A1(\mem[6][2] ), .A2(n96), .ZN(n99) );
  OAI21_X1 U137 ( .B1(n293), .B2(n96), .A(n100), .ZN(n197) );
  NAND2_X1 U138 ( .A1(\mem[6][3] ), .A2(n96), .ZN(n100) );
  OAI21_X1 U139 ( .B1(n292), .B2(n96), .A(n101), .ZN(n198) );
  NAND2_X1 U140 ( .A1(\mem[6][4] ), .A2(n96), .ZN(n101) );
  OAI21_X1 U141 ( .B1(n291), .B2(n96), .A(n102), .ZN(n199) );
  NAND2_X1 U142 ( .A1(\mem[6][5] ), .A2(n96), .ZN(n102) );
  OAI21_X1 U143 ( .B1(n290), .B2(n96), .A(n103), .ZN(n200) );
  NAND2_X1 U144 ( .A1(\mem[6][6] ), .A2(n96), .ZN(n103) );
  OAI21_X1 U145 ( .B1(n289), .B2(n96), .A(n104), .ZN(n201) );
  NAND2_X1 U146 ( .A1(\mem[6][7] ), .A2(n96), .ZN(n104) );
  OAI21_X1 U147 ( .B1(n288), .B2(n96), .A(n105), .ZN(n202) );
  NAND2_X1 U148 ( .A1(\mem[6][8] ), .A2(n96), .ZN(n105) );
  OAI21_X1 U149 ( .B1(n287), .B2(n96), .A(n106), .ZN(n203) );
  NAND2_X1 U150 ( .A1(\mem[6][9] ), .A2(n96), .ZN(n106) );
  OAI21_X1 U151 ( .B1(n286), .B2(n96), .A(n107), .ZN(n204) );
  NAND2_X1 U152 ( .A1(\mem[6][10] ), .A2(n96), .ZN(n107) );
  OAI21_X1 U153 ( .B1(n285), .B2(n96), .A(n108), .ZN(n205) );
  NAND2_X1 U154 ( .A1(\mem[6][11] ), .A2(n96), .ZN(n108) );
  OAI21_X1 U155 ( .B1(n296), .B2(n109), .A(n110), .ZN(n206) );
  NAND2_X1 U156 ( .A1(\mem[7][0] ), .A2(n109), .ZN(n110) );
  OAI21_X1 U157 ( .B1(n295), .B2(n109), .A(n111), .ZN(n207) );
  NAND2_X1 U158 ( .A1(\mem[7][1] ), .A2(n109), .ZN(n111) );
  OAI21_X1 U159 ( .B1(n294), .B2(n109), .A(n112), .ZN(n208) );
  NAND2_X1 U160 ( .A1(\mem[7][2] ), .A2(n109), .ZN(n112) );
  OAI21_X1 U161 ( .B1(n293), .B2(n109), .A(n113), .ZN(n209) );
  NAND2_X1 U162 ( .A1(\mem[7][3] ), .A2(n109), .ZN(n113) );
  OAI21_X1 U163 ( .B1(n292), .B2(n109), .A(n114), .ZN(n210) );
  NAND2_X1 U164 ( .A1(\mem[7][4] ), .A2(n109), .ZN(n114) );
  OAI21_X1 U165 ( .B1(n291), .B2(n109), .A(n115), .ZN(n211) );
  NAND2_X1 U166 ( .A1(\mem[7][5] ), .A2(n109), .ZN(n115) );
  OAI21_X1 U167 ( .B1(n290), .B2(n109), .A(n116), .ZN(n212) );
  NAND2_X1 U168 ( .A1(\mem[7][6] ), .A2(n109), .ZN(n116) );
  OAI21_X1 U169 ( .B1(n289), .B2(n109), .A(n117), .ZN(n213) );
  NAND2_X1 U170 ( .A1(\mem[7][7] ), .A2(n109), .ZN(n117) );
  OAI21_X1 U171 ( .B1(n288), .B2(n109), .A(n118), .ZN(n214) );
  NAND2_X1 U172 ( .A1(\mem[7][8] ), .A2(n109), .ZN(n118) );
  OAI21_X1 U173 ( .B1(n287), .B2(n109), .A(n119), .ZN(n215) );
  NAND2_X1 U174 ( .A1(\mem[7][9] ), .A2(n109), .ZN(n119) );
  OAI21_X1 U175 ( .B1(n286), .B2(n109), .A(n120), .ZN(n216) );
  NAND2_X1 U176 ( .A1(\mem[7][10] ), .A2(n109), .ZN(n120) );
  OAI21_X1 U177 ( .B1(n285), .B2(n109), .A(n121), .ZN(n217) );
  NAND2_X1 U178 ( .A1(\mem[7][11] ), .A2(n109), .ZN(n121) );
  OAI21_X1 U179 ( .B1(n16), .B2(n296), .A(n17), .ZN(n122) );
  NAND2_X1 U180 ( .A1(\mem[0][0] ), .A2(n16), .ZN(n17) );
  OAI21_X1 U181 ( .B1(n16), .B2(n295), .A(n18), .ZN(n123) );
  NAND2_X1 U182 ( .A1(\mem[0][1] ), .A2(n16), .ZN(n18) );
  OAI21_X1 U183 ( .B1(n16), .B2(n294), .A(n19), .ZN(n124) );
  NAND2_X1 U184 ( .A1(\mem[0][2] ), .A2(n16), .ZN(n19) );
  OAI21_X1 U185 ( .B1(n16), .B2(n293), .A(n20), .ZN(n125) );
  NAND2_X1 U186 ( .A1(\mem[0][3] ), .A2(n16), .ZN(n20) );
  OAI21_X1 U187 ( .B1(n16), .B2(n292), .A(n21), .ZN(n126) );
  NAND2_X1 U188 ( .A1(\mem[0][4] ), .A2(n16), .ZN(n21) );
  OAI21_X1 U189 ( .B1(n16), .B2(n291), .A(n22), .ZN(n127) );
  NAND2_X1 U190 ( .A1(\mem[0][5] ), .A2(n16), .ZN(n22) );
  OAI21_X1 U191 ( .B1(n16), .B2(n290), .A(n23), .ZN(n128) );
  NAND2_X1 U192 ( .A1(\mem[0][6] ), .A2(n16), .ZN(n23) );
  OAI21_X1 U193 ( .B1(n16), .B2(n289), .A(n24), .ZN(n129) );
  NAND2_X1 U194 ( .A1(\mem[0][7] ), .A2(n16), .ZN(n24) );
  OAI21_X1 U195 ( .B1(n16), .B2(n288), .A(n25), .ZN(n130) );
  NAND2_X1 U196 ( .A1(\mem[0][8] ), .A2(n16), .ZN(n25) );
  OAI21_X1 U197 ( .B1(n16), .B2(n287), .A(n26), .ZN(n131) );
  NAND2_X1 U198 ( .A1(\mem[0][9] ), .A2(n16), .ZN(n26) );
  OAI21_X1 U199 ( .B1(n16), .B2(n286), .A(n27), .ZN(n132) );
  NAND2_X1 U200 ( .A1(\mem[0][10] ), .A2(n16), .ZN(n27) );
  OAI21_X1 U201 ( .B1(n16), .B2(n285), .A(n28), .ZN(n133) );
  NAND2_X1 U202 ( .A1(\mem[0][11] ), .A2(n16), .ZN(n28) );
  INV_X1 U203 ( .A(data_in[0]), .ZN(n296) );
  INV_X1 U204 ( .A(data_in[1]), .ZN(n295) );
  INV_X1 U205 ( .A(data_in[2]), .ZN(n294) );
  INV_X1 U206 ( .A(data_in[3]), .ZN(n293) );
  INV_X1 U207 ( .A(data_in[4]), .ZN(n292) );
  INV_X1 U208 ( .A(data_in[5]), .ZN(n291) );
  INV_X1 U209 ( .A(data_in[6]), .ZN(n290) );
  INV_X1 U210 ( .A(data_in[7]), .ZN(n289) );
  INV_X1 U211 ( .A(data_in[8]), .ZN(n288) );
  INV_X1 U220 ( .A(data_in[9]), .ZN(n287) );
  INV_X1 U221 ( .A(data_in[10]), .ZN(n286) );
  INV_X1 U222 ( .A(data_in[11]), .ZN(n285) );
  MUX2_X1 U223 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n280), .Z(n5) );
  MUX2_X1 U224 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n280), .Z(n6) );
  MUX2_X1 U225 ( .A(n6), .B(n5), .S(n279), .Z(n7) );
  MUX2_X1 U226 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n280), .Z(n8) );
  MUX2_X1 U227 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n280), .Z(n9) );
  MUX2_X1 U228 ( .A(n9), .B(n8), .S(n279), .Z(n10) );
  MUX2_X1 U229 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n280), .Z(n11) );
  MUX2_X1 U230 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n280), .Z(n12) );
  MUX2_X1 U231 ( .A(n12), .B(n11), .S(n279), .Z(n13) );
  MUX2_X1 U232 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n280), .Z(n14) );
  MUX2_X1 U233 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n280), .Z(n15) );
  MUX2_X1 U234 ( .A(n15), .B(n14), .S(n279), .Z(n218) );
  MUX2_X1 U235 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n280), .Z(n219) );
  MUX2_X1 U236 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n280), .Z(n220) );
  MUX2_X1 U237 ( .A(n220), .B(n219), .S(n279), .Z(n221) );
  MUX2_X1 U238 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n280), .Z(n222) );
  MUX2_X1 U239 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n280), .Z(n223) );
  MUX2_X1 U240 ( .A(n223), .B(n222), .S(n279), .Z(n224) );
  MUX2_X1 U241 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n281), .Z(n225) );
  MUX2_X1 U242 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n281), .Z(n226) );
  MUX2_X1 U243 ( .A(n226), .B(n225), .S(n279), .Z(n227) );
  MUX2_X1 U244 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n228) );
  MUX2_X1 U245 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n229) );
  MUX2_X1 U246 ( .A(n229), .B(n228), .S(n279), .Z(n230) );
  MUX2_X1 U247 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(N10), .Z(n231) );
  MUX2_X1 U248 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n281), .Z(n232) );
  MUX2_X1 U249 ( .A(n232), .B(n231), .S(n279), .Z(n233) );
  MUX2_X1 U250 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(N10), .Z(n234) );
  MUX2_X1 U251 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n235) );
  MUX2_X1 U252 ( .A(n235), .B(n234), .S(n279), .Z(n236) );
  MUX2_X1 U253 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n281), .Z(n237) );
  MUX2_X1 U254 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n281), .Z(n238) );
  MUX2_X1 U255 ( .A(n238), .B(n237), .S(n279), .Z(n239) );
  MUX2_X1 U256 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n240) );
  MUX2_X1 U257 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(N10), .Z(n241) );
  MUX2_X1 U258 ( .A(n241), .B(n240), .S(n279), .Z(n242) );
  MUX2_X1 U259 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n281), .Z(n243) );
  MUX2_X1 U260 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n281), .Z(n244) );
  MUX2_X1 U261 ( .A(n244), .B(n243), .S(n279), .Z(n245) );
  MUX2_X1 U262 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n281), .Z(n246) );
  MUX2_X1 U263 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n281), .Z(n247) );
  MUX2_X1 U264 ( .A(n247), .B(n246), .S(n279), .Z(n248) );
  MUX2_X1 U265 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n281), .Z(n249) );
  MUX2_X1 U266 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n281), .Z(n250) );
  MUX2_X1 U267 ( .A(n250), .B(n249), .S(n279), .Z(n251) );
  MUX2_X1 U268 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n281), .Z(n252) );
  MUX2_X1 U269 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n281), .Z(n253) );
  MUX2_X1 U270 ( .A(n253), .B(n252), .S(n279), .Z(n254) );
  MUX2_X1 U271 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n281), .Z(n255) );
  MUX2_X1 U272 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n281), .Z(n256) );
  MUX2_X1 U273 ( .A(n256), .B(n255), .S(n279), .Z(n257) );
  MUX2_X1 U274 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n281), .Z(n258) );
  MUX2_X1 U275 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n281), .Z(n259) );
  MUX2_X1 U276 ( .A(n259), .B(n258), .S(n279), .Z(n260) );
  MUX2_X1 U277 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n281), .Z(n261) );
  MUX2_X1 U278 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(N10), .Z(n262) );
  MUX2_X1 U279 ( .A(n262), .B(n261), .S(n279), .Z(n263) );
  MUX2_X1 U280 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(N10), .Z(n264) );
  MUX2_X1 U281 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n281), .Z(n265) );
  MUX2_X1 U282 ( .A(n265), .B(n264), .S(n279), .Z(n266) );
  MUX2_X1 U283 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n281), .Z(n267) );
  MUX2_X1 U284 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(N10), .Z(n268) );
  MUX2_X1 U285 ( .A(n268), .B(n267), .S(n279), .Z(n269) );
  MUX2_X1 U286 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(N10), .Z(n270) );
  MUX2_X1 U287 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n281), .Z(n271) );
  MUX2_X1 U288 ( .A(n271), .B(n270), .S(n279), .Z(n272) );
  MUX2_X1 U289 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(N10), .Z(n273) );
  MUX2_X1 U290 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(N10), .Z(n274) );
  MUX2_X1 U291 ( .A(n274), .B(n273), .S(n279), .Z(n275) );
  MUX2_X1 U292 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(N10), .Z(n276) );
  MUX2_X1 U293 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n281), .Z(n277) );
  MUX2_X1 U294 ( .A(n277), .B(n276), .S(N11), .Z(n278) );
endmodule


module memory_WIDTH12_SIZE8_LOGSIZE3_8 ( clk, data_in, data_out, addr, wr_en
 );
  input [11:0] data_in;
  output [11:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] ,
         \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] ,
         \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][11] , \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] ,
         \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] ,
         \mem[5][1] , \mem[5][0] , \mem[4][11] , \mem[4][10] , \mem[4][9] ,
         \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] ,
         \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] ,
         \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] ,
         \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][11] , \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] ,
         \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] ,
         \mem[0][1] , \mem[0][0] , N13, N18, N21, N22, N23, N24, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[11]  ( .D(N13), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[6]  ( .D(N18), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[3]  ( .D(N21), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N22), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N23), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N24), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][11]  ( .D(n293), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n294), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n295), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n296), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n297), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n298), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n299), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n300), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n301), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n302), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n303), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n304), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n305), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n306), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n307), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n308), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n309), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n310), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n311), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n312), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n313), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n314), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n315), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n316), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n317), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n318), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n319), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n320), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n321), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n322), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n323), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n324), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n325), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n326), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n327), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n328), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n329), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n330), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n331), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n332), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n333), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n334), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n335), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n336), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n337), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n338), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n339), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n340), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n341), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n342), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n343), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n344), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n345), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n346), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n347), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n348), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n349), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n350), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n351), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n352), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n353), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n354), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n355), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n356), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n357), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n358), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n359), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n360), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n361), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n362), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n363), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n364), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n365), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n366), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n367), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n368), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n369), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n370), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n371), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n372), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n373), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n374), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n375), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n376), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n377), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n378), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n379), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n380), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n381), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n382), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n383), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n384), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n385), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n386), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n387), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n388), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U212 ( .A1(n278), .A2(n279), .A3(n481), .ZN(n494) );
  NAND3_X1 U213 ( .A1(n481), .A2(n279), .A3(N10), .ZN(n480) );
  NAND3_X1 U214 ( .A1(n481), .A2(n278), .A3(N11), .ZN(n467) );
  NAND3_X1 U215 ( .A1(N10), .A2(n481), .A3(N11), .ZN(n454) );
  NAND3_X1 U216 ( .A1(n278), .A2(n279), .A3(n428), .ZN(n441) );
  NAND3_X1 U217 ( .A1(N10), .A2(n279), .A3(n428), .ZN(n427) );
  NAND3_X1 U218 ( .A1(N11), .A2(n278), .A3(n428), .ZN(n414) );
  NAND3_X1 U219 ( .A1(N11), .A2(N10), .A3(n428), .ZN(n401) );
  SDFF_X1 \data_out_reg[7]  ( .D(n250), .SI(n247), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n238), .SI(n235), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[4]  ( .D(n232), .SI(n229), .SE(N12), .CK(clk), .Q(
        data_out[4]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n262), .SI(n259), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[8]  ( .D(n256), .SI(n253), .SE(N12), .CK(clk), .Q(
        data_out[8]) );
  SDFF_X1 \data_out_reg[10]  ( .D(n268), .SI(n265), .SE(N12), .CK(clk), .Q(
        data_out[10]) );
  BUF_X1 U3 ( .A(n277), .Z(n276) );
  BUF_X1 U4 ( .A(N11), .Z(n275) );
  BUF_X1 U5 ( .A(N10), .Z(n277) );
  NOR2_X1 U6 ( .A1(n280), .A2(N12), .ZN(n481) );
  INV_X1 U7 ( .A(wr_en), .ZN(n280) );
  AND2_X1 U8 ( .A1(N12), .A2(wr_en), .ZN(n428) );
  INV_X1 U9 ( .A(N10), .ZN(n278) );
  INV_X1 U10 ( .A(N11), .ZN(n279) );
  OAI21_X1 U11 ( .B1(n292), .B2(n480), .A(n479), .ZN(n376) );
  NAND2_X1 U12 ( .A1(\mem[1][0] ), .A2(n480), .ZN(n479) );
  OAI21_X1 U13 ( .B1(n291), .B2(n480), .A(n478), .ZN(n375) );
  NAND2_X1 U14 ( .A1(\mem[1][1] ), .A2(n480), .ZN(n478) );
  OAI21_X1 U15 ( .B1(n290), .B2(n480), .A(n477), .ZN(n374) );
  NAND2_X1 U16 ( .A1(\mem[1][2] ), .A2(n480), .ZN(n477) );
  OAI21_X1 U17 ( .B1(n289), .B2(n480), .A(n476), .ZN(n373) );
  NAND2_X1 U18 ( .A1(\mem[1][3] ), .A2(n480), .ZN(n476) );
  OAI21_X1 U19 ( .B1(n288), .B2(n480), .A(n475), .ZN(n372) );
  NAND2_X1 U20 ( .A1(\mem[1][4] ), .A2(n480), .ZN(n475) );
  OAI21_X1 U21 ( .B1(n287), .B2(n480), .A(n474), .ZN(n371) );
  NAND2_X1 U22 ( .A1(\mem[1][5] ), .A2(n480), .ZN(n474) );
  OAI21_X1 U23 ( .B1(n286), .B2(n480), .A(n473), .ZN(n370) );
  NAND2_X1 U24 ( .A1(\mem[1][6] ), .A2(n480), .ZN(n473) );
  OAI21_X1 U25 ( .B1(n285), .B2(n480), .A(n472), .ZN(n369) );
  NAND2_X1 U26 ( .A1(\mem[1][7] ), .A2(n480), .ZN(n472) );
  OAI21_X1 U27 ( .B1(n284), .B2(n480), .A(n471), .ZN(n368) );
  NAND2_X1 U28 ( .A1(\mem[1][8] ), .A2(n480), .ZN(n471) );
  OAI21_X1 U29 ( .B1(n283), .B2(n480), .A(n470), .ZN(n367) );
  NAND2_X1 U30 ( .A1(\mem[1][9] ), .A2(n480), .ZN(n470) );
  OAI21_X1 U31 ( .B1(n282), .B2(n480), .A(n469), .ZN(n366) );
  NAND2_X1 U32 ( .A1(\mem[1][10] ), .A2(n480), .ZN(n469) );
  OAI21_X1 U33 ( .B1(n281), .B2(n480), .A(n468), .ZN(n365) );
  NAND2_X1 U34 ( .A1(\mem[1][11] ), .A2(n480), .ZN(n468) );
  OAI21_X1 U35 ( .B1(n292), .B2(n467), .A(n466), .ZN(n364) );
  NAND2_X1 U36 ( .A1(\mem[2][0] ), .A2(n467), .ZN(n466) );
  OAI21_X1 U37 ( .B1(n291), .B2(n467), .A(n465), .ZN(n363) );
  NAND2_X1 U38 ( .A1(\mem[2][1] ), .A2(n467), .ZN(n465) );
  OAI21_X1 U39 ( .B1(n290), .B2(n467), .A(n464), .ZN(n362) );
  NAND2_X1 U40 ( .A1(\mem[2][2] ), .A2(n467), .ZN(n464) );
  OAI21_X1 U41 ( .B1(n289), .B2(n467), .A(n463), .ZN(n361) );
  NAND2_X1 U42 ( .A1(\mem[2][3] ), .A2(n467), .ZN(n463) );
  OAI21_X1 U43 ( .B1(n288), .B2(n467), .A(n462), .ZN(n360) );
  NAND2_X1 U44 ( .A1(\mem[2][4] ), .A2(n467), .ZN(n462) );
  OAI21_X1 U45 ( .B1(n287), .B2(n467), .A(n461), .ZN(n359) );
  NAND2_X1 U46 ( .A1(\mem[2][5] ), .A2(n467), .ZN(n461) );
  OAI21_X1 U47 ( .B1(n286), .B2(n467), .A(n460), .ZN(n358) );
  NAND2_X1 U48 ( .A1(\mem[2][6] ), .A2(n467), .ZN(n460) );
  OAI21_X1 U49 ( .B1(n285), .B2(n467), .A(n459), .ZN(n357) );
  NAND2_X1 U50 ( .A1(\mem[2][7] ), .A2(n467), .ZN(n459) );
  OAI21_X1 U51 ( .B1(n284), .B2(n467), .A(n458), .ZN(n356) );
  NAND2_X1 U52 ( .A1(\mem[2][8] ), .A2(n467), .ZN(n458) );
  OAI21_X1 U53 ( .B1(n283), .B2(n467), .A(n457), .ZN(n355) );
  NAND2_X1 U54 ( .A1(\mem[2][9] ), .A2(n467), .ZN(n457) );
  OAI21_X1 U55 ( .B1(n282), .B2(n467), .A(n456), .ZN(n354) );
  NAND2_X1 U56 ( .A1(\mem[2][10] ), .A2(n467), .ZN(n456) );
  OAI21_X1 U57 ( .B1(n281), .B2(n467), .A(n455), .ZN(n353) );
  NAND2_X1 U58 ( .A1(\mem[2][11] ), .A2(n467), .ZN(n455) );
  OAI21_X1 U59 ( .B1(n292), .B2(n454), .A(n453), .ZN(n352) );
  NAND2_X1 U60 ( .A1(\mem[3][0] ), .A2(n454), .ZN(n453) );
  OAI21_X1 U61 ( .B1(n291), .B2(n454), .A(n452), .ZN(n351) );
  NAND2_X1 U62 ( .A1(\mem[3][1] ), .A2(n454), .ZN(n452) );
  OAI21_X1 U63 ( .B1(n290), .B2(n454), .A(n451), .ZN(n350) );
  NAND2_X1 U64 ( .A1(\mem[3][2] ), .A2(n454), .ZN(n451) );
  OAI21_X1 U65 ( .B1(n289), .B2(n454), .A(n450), .ZN(n349) );
  NAND2_X1 U66 ( .A1(\mem[3][3] ), .A2(n454), .ZN(n450) );
  OAI21_X1 U67 ( .B1(n288), .B2(n454), .A(n449), .ZN(n348) );
  NAND2_X1 U68 ( .A1(\mem[3][4] ), .A2(n454), .ZN(n449) );
  OAI21_X1 U69 ( .B1(n287), .B2(n454), .A(n448), .ZN(n347) );
  NAND2_X1 U70 ( .A1(\mem[3][5] ), .A2(n454), .ZN(n448) );
  OAI21_X1 U71 ( .B1(n286), .B2(n454), .A(n447), .ZN(n346) );
  NAND2_X1 U72 ( .A1(\mem[3][6] ), .A2(n454), .ZN(n447) );
  OAI21_X1 U73 ( .B1(n285), .B2(n454), .A(n446), .ZN(n345) );
  NAND2_X1 U74 ( .A1(\mem[3][7] ), .A2(n454), .ZN(n446) );
  OAI21_X1 U75 ( .B1(n284), .B2(n454), .A(n445), .ZN(n344) );
  NAND2_X1 U76 ( .A1(\mem[3][8] ), .A2(n454), .ZN(n445) );
  OAI21_X1 U77 ( .B1(n283), .B2(n454), .A(n444), .ZN(n343) );
  NAND2_X1 U78 ( .A1(\mem[3][9] ), .A2(n454), .ZN(n444) );
  OAI21_X1 U79 ( .B1(n282), .B2(n454), .A(n443), .ZN(n342) );
  NAND2_X1 U80 ( .A1(\mem[3][10] ), .A2(n454), .ZN(n443) );
  OAI21_X1 U81 ( .B1(n281), .B2(n454), .A(n442), .ZN(n341) );
  NAND2_X1 U82 ( .A1(\mem[3][11] ), .A2(n454), .ZN(n442) );
  OAI21_X1 U83 ( .B1(n292), .B2(n441), .A(n440), .ZN(n340) );
  NAND2_X1 U84 ( .A1(\mem[4][0] ), .A2(n441), .ZN(n440) );
  OAI21_X1 U85 ( .B1(n291), .B2(n441), .A(n439), .ZN(n339) );
  NAND2_X1 U86 ( .A1(\mem[4][1] ), .A2(n441), .ZN(n439) );
  OAI21_X1 U87 ( .B1(n290), .B2(n441), .A(n438), .ZN(n338) );
  NAND2_X1 U88 ( .A1(\mem[4][2] ), .A2(n441), .ZN(n438) );
  OAI21_X1 U89 ( .B1(n289), .B2(n441), .A(n437), .ZN(n337) );
  NAND2_X1 U90 ( .A1(\mem[4][3] ), .A2(n441), .ZN(n437) );
  OAI21_X1 U91 ( .B1(n288), .B2(n441), .A(n436), .ZN(n336) );
  NAND2_X1 U92 ( .A1(\mem[4][4] ), .A2(n441), .ZN(n436) );
  OAI21_X1 U93 ( .B1(n287), .B2(n441), .A(n435), .ZN(n335) );
  NAND2_X1 U94 ( .A1(\mem[4][5] ), .A2(n441), .ZN(n435) );
  OAI21_X1 U95 ( .B1(n286), .B2(n441), .A(n434), .ZN(n334) );
  NAND2_X1 U96 ( .A1(\mem[4][6] ), .A2(n441), .ZN(n434) );
  OAI21_X1 U97 ( .B1(n285), .B2(n441), .A(n433), .ZN(n333) );
  NAND2_X1 U98 ( .A1(\mem[4][7] ), .A2(n441), .ZN(n433) );
  OAI21_X1 U99 ( .B1(n284), .B2(n441), .A(n432), .ZN(n332) );
  NAND2_X1 U100 ( .A1(\mem[4][8] ), .A2(n441), .ZN(n432) );
  OAI21_X1 U101 ( .B1(n283), .B2(n441), .A(n431), .ZN(n331) );
  NAND2_X1 U102 ( .A1(\mem[4][9] ), .A2(n441), .ZN(n431) );
  OAI21_X1 U103 ( .B1(n282), .B2(n441), .A(n430), .ZN(n330) );
  NAND2_X1 U104 ( .A1(\mem[4][10] ), .A2(n441), .ZN(n430) );
  OAI21_X1 U105 ( .B1(n281), .B2(n441), .A(n429), .ZN(n329) );
  NAND2_X1 U106 ( .A1(\mem[4][11] ), .A2(n441), .ZN(n429) );
  OAI21_X1 U107 ( .B1(n292), .B2(n427), .A(n426), .ZN(n328) );
  NAND2_X1 U108 ( .A1(\mem[5][0] ), .A2(n427), .ZN(n426) );
  OAI21_X1 U109 ( .B1(n291), .B2(n427), .A(n425), .ZN(n327) );
  NAND2_X1 U110 ( .A1(\mem[5][1] ), .A2(n427), .ZN(n425) );
  OAI21_X1 U111 ( .B1(n290), .B2(n427), .A(n424), .ZN(n326) );
  NAND2_X1 U112 ( .A1(\mem[5][2] ), .A2(n427), .ZN(n424) );
  OAI21_X1 U113 ( .B1(n289), .B2(n427), .A(n423), .ZN(n325) );
  NAND2_X1 U114 ( .A1(\mem[5][3] ), .A2(n427), .ZN(n423) );
  OAI21_X1 U115 ( .B1(n288), .B2(n427), .A(n422), .ZN(n324) );
  NAND2_X1 U116 ( .A1(\mem[5][4] ), .A2(n427), .ZN(n422) );
  OAI21_X1 U117 ( .B1(n287), .B2(n427), .A(n421), .ZN(n323) );
  NAND2_X1 U118 ( .A1(\mem[5][5] ), .A2(n427), .ZN(n421) );
  OAI21_X1 U119 ( .B1(n286), .B2(n427), .A(n420), .ZN(n322) );
  NAND2_X1 U120 ( .A1(\mem[5][6] ), .A2(n427), .ZN(n420) );
  OAI21_X1 U121 ( .B1(n285), .B2(n427), .A(n419), .ZN(n321) );
  NAND2_X1 U122 ( .A1(\mem[5][7] ), .A2(n427), .ZN(n419) );
  OAI21_X1 U123 ( .B1(n284), .B2(n427), .A(n418), .ZN(n320) );
  NAND2_X1 U124 ( .A1(\mem[5][8] ), .A2(n427), .ZN(n418) );
  OAI21_X1 U125 ( .B1(n283), .B2(n427), .A(n417), .ZN(n319) );
  NAND2_X1 U126 ( .A1(\mem[5][9] ), .A2(n427), .ZN(n417) );
  OAI21_X1 U127 ( .B1(n282), .B2(n427), .A(n416), .ZN(n318) );
  NAND2_X1 U128 ( .A1(\mem[5][10] ), .A2(n427), .ZN(n416) );
  OAI21_X1 U129 ( .B1(n281), .B2(n427), .A(n415), .ZN(n317) );
  NAND2_X1 U130 ( .A1(\mem[5][11] ), .A2(n427), .ZN(n415) );
  OAI21_X1 U131 ( .B1(n292), .B2(n414), .A(n413), .ZN(n316) );
  NAND2_X1 U132 ( .A1(\mem[6][0] ), .A2(n414), .ZN(n413) );
  OAI21_X1 U133 ( .B1(n291), .B2(n414), .A(n412), .ZN(n315) );
  NAND2_X1 U134 ( .A1(\mem[6][1] ), .A2(n414), .ZN(n412) );
  OAI21_X1 U135 ( .B1(n290), .B2(n414), .A(n411), .ZN(n314) );
  NAND2_X1 U136 ( .A1(\mem[6][2] ), .A2(n414), .ZN(n411) );
  OAI21_X1 U137 ( .B1(n289), .B2(n414), .A(n410), .ZN(n313) );
  NAND2_X1 U138 ( .A1(\mem[6][3] ), .A2(n414), .ZN(n410) );
  OAI21_X1 U139 ( .B1(n288), .B2(n414), .A(n409), .ZN(n312) );
  NAND2_X1 U140 ( .A1(\mem[6][4] ), .A2(n414), .ZN(n409) );
  OAI21_X1 U141 ( .B1(n287), .B2(n414), .A(n408), .ZN(n311) );
  NAND2_X1 U142 ( .A1(\mem[6][5] ), .A2(n414), .ZN(n408) );
  OAI21_X1 U143 ( .B1(n286), .B2(n414), .A(n407), .ZN(n310) );
  NAND2_X1 U144 ( .A1(\mem[6][6] ), .A2(n414), .ZN(n407) );
  OAI21_X1 U145 ( .B1(n285), .B2(n414), .A(n406), .ZN(n309) );
  NAND2_X1 U146 ( .A1(\mem[6][7] ), .A2(n414), .ZN(n406) );
  OAI21_X1 U147 ( .B1(n284), .B2(n414), .A(n405), .ZN(n308) );
  NAND2_X1 U148 ( .A1(\mem[6][8] ), .A2(n414), .ZN(n405) );
  OAI21_X1 U149 ( .B1(n283), .B2(n414), .A(n404), .ZN(n307) );
  NAND2_X1 U150 ( .A1(\mem[6][9] ), .A2(n414), .ZN(n404) );
  OAI21_X1 U151 ( .B1(n282), .B2(n414), .A(n403), .ZN(n306) );
  NAND2_X1 U152 ( .A1(\mem[6][10] ), .A2(n414), .ZN(n403) );
  OAI21_X1 U153 ( .B1(n281), .B2(n414), .A(n402), .ZN(n305) );
  NAND2_X1 U154 ( .A1(\mem[6][11] ), .A2(n414), .ZN(n402) );
  OAI21_X1 U155 ( .B1(n292), .B2(n401), .A(n400), .ZN(n304) );
  NAND2_X1 U156 ( .A1(\mem[7][0] ), .A2(n401), .ZN(n400) );
  OAI21_X1 U157 ( .B1(n291), .B2(n401), .A(n399), .ZN(n303) );
  NAND2_X1 U158 ( .A1(\mem[7][1] ), .A2(n401), .ZN(n399) );
  OAI21_X1 U159 ( .B1(n290), .B2(n401), .A(n398), .ZN(n302) );
  NAND2_X1 U160 ( .A1(\mem[7][2] ), .A2(n401), .ZN(n398) );
  OAI21_X1 U161 ( .B1(n289), .B2(n401), .A(n397), .ZN(n301) );
  NAND2_X1 U162 ( .A1(\mem[7][3] ), .A2(n401), .ZN(n397) );
  OAI21_X1 U163 ( .B1(n288), .B2(n401), .A(n396), .ZN(n300) );
  NAND2_X1 U164 ( .A1(\mem[7][4] ), .A2(n401), .ZN(n396) );
  OAI21_X1 U165 ( .B1(n287), .B2(n401), .A(n395), .ZN(n299) );
  NAND2_X1 U166 ( .A1(\mem[7][5] ), .A2(n401), .ZN(n395) );
  OAI21_X1 U167 ( .B1(n286), .B2(n401), .A(n394), .ZN(n298) );
  NAND2_X1 U168 ( .A1(\mem[7][6] ), .A2(n401), .ZN(n394) );
  OAI21_X1 U169 ( .B1(n285), .B2(n401), .A(n393), .ZN(n297) );
  NAND2_X1 U170 ( .A1(\mem[7][7] ), .A2(n401), .ZN(n393) );
  OAI21_X1 U171 ( .B1(n284), .B2(n401), .A(n392), .ZN(n296) );
  NAND2_X1 U172 ( .A1(\mem[7][8] ), .A2(n401), .ZN(n392) );
  OAI21_X1 U173 ( .B1(n283), .B2(n401), .A(n391), .ZN(n295) );
  NAND2_X1 U174 ( .A1(\mem[7][9] ), .A2(n401), .ZN(n391) );
  OAI21_X1 U175 ( .B1(n282), .B2(n401), .A(n390), .ZN(n294) );
  NAND2_X1 U176 ( .A1(\mem[7][10] ), .A2(n401), .ZN(n390) );
  OAI21_X1 U177 ( .B1(n281), .B2(n401), .A(n389), .ZN(n293) );
  NAND2_X1 U178 ( .A1(\mem[7][11] ), .A2(n401), .ZN(n389) );
  OAI21_X1 U179 ( .B1(n494), .B2(n292), .A(n493), .ZN(n388) );
  NAND2_X1 U180 ( .A1(\mem[0][0] ), .A2(n494), .ZN(n493) );
  OAI21_X1 U181 ( .B1(n494), .B2(n291), .A(n492), .ZN(n387) );
  NAND2_X1 U182 ( .A1(\mem[0][1] ), .A2(n494), .ZN(n492) );
  OAI21_X1 U183 ( .B1(n494), .B2(n290), .A(n491), .ZN(n386) );
  NAND2_X1 U184 ( .A1(\mem[0][2] ), .A2(n494), .ZN(n491) );
  OAI21_X1 U185 ( .B1(n494), .B2(n289), .A(n490), .ZN(n385) );
  NAND2_X1 U186 ( .A1(\mem[0][3] ), .A2(n494), .ZN(n490) );
  OAI21_X1 U187 ( .B1(n494), .B2(n288), .A(n489), .ZN(n384) );
  NAND2_X1 U188 ( .A1(\mem[0][4] ), .A2(n494), .ZN(n489) );
  OAI21_X1 U189 ( .B1(n494), .B2(n287), .A(n488), .ZN(n383) );
  NAND2_X1 U190 ( .A1(\mem[0][5] ), .A2(n494), .ZN(n488) );
  OAI21_X1 U191 ( .B1(n494), .B2(n286), .A(n487), .ZN(n382) );
  NAND2_X1 U192 ( .A1(\mem[0][6] ), .A2(n494), .ZN(n487) );
  OAI21_X1 U193 ( .B1(n494), .B2(n285), .A(n486), .ZN(n381) );
  NAND2_X1 U194 ( .A1(\mem[0][7] ), .A2(n494), .ZN(n486) );
  OAI21_X1 U195 ( .B1(n494), .B2(n284), .A(n485), .ZN(n380) );
  NAND2_X1 U196 ( .A1(\mem[0][8] ), .A2(n494), .ZN(n485) );
  OAI21_X1 U197 ( .B1(n494), .B2(n283), .A(n484), .ZN(n379) );
  NAND2_X1 U198 ( .A1(\mem[0][9] ), .A2(n494), .ZN(n484) );
  OAI21_X1 U199 ( .B1(n494), .B2(n282), .A(n483), .ZN(n378) );
  NAND2_X1 U200 ( .A1(\mem[0][10] ), .A2(n494), .ZN(n483) );
  OAI21_X1 U201 ( .B1(n494), .B2(n281), .A(n482), .ZN(n377) );
  NAND2_X1 U202 ( .A1(\mem[0][11] ), .A2(n494), .ZN(n482) );
  INV_X1 U203 ( .A(data_in[0]), .ZN(n292) );
  INV_X1 U204 ( .A(data_in[1]), .ZN(n291) );
  INV_X1 U205 ( .A(data_in[2]), .ZN(n290) );
  INV_X1 U206 ( .A(data_in[3]), .ZN(n289) );
  INV_X1 U207 ( .A(data_in[4]), .ZN(n288) );
  INV_X1 U208 ( .A(data_in[5]), .ZN(n287) );
  INV_X1 U209 ( .A(data_in[6]), .ZN(n286) );
  INV_X1 U210 ( .A(data_in[7]), .ZN(n285) );
  INV_X1 U211 ( .A(data_in[8]), .ZN(n284) );
  INV_X1 U220 ( .A(data_in[9]), .ZN(n283) );
  INV_X1 U221 ( .A(data_in[10]), .ZN(n282) );
  INV_X1 U222 ( .A(data_in[11]), .ZN(n281) );
  MUX2_X1 U223 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n276), .Z(n1) );
  MUX2_X1 U224 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n276), .Z(n2) );
  MUX2_X1 U225 ( .A(n2), .B(n1), .S(n275), .Z(n3) );
  MUX2_X1 U226 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n276), .Z(n4) );
  MUX2_X1 U227 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n276), .Z(n5) );
  MUX2_X1 U228 ( .A(n5), .B(n4), .S(n275), .Z(n6) );
  MUX2_X1 U229 ( .A(n6), .B(n3), .S(N12), .Z(N24) );
  MUX2_X1 U230 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n276), .Z(n7) );
  MUX2_X1 U231 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n276), .Z(n8) );
  MUX2_X1 U232 ( .A(n8), .B(n7), .S(n275), .Z(n9) );
  MUX2_X1 U233 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n276), .Z(n10) );
  MUX2_X1 U234 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n276), .Z(n11) );
  MUX2_X1 U235 ( .A(n11), .B(n10), .S(n275), .Z(n12) );
  MUX2_X1 U236 ( .A(n12), .B(n9), .S(N12), .Z(N23) );
  MUX2_X1 U237 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n276), .Z(n13) );
  MUX2_X1 U238 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n276), .Z(n14) );
  MUX2_X1 U239 ( .A(n14), .B(n13), .S(n275), .Z(n15) );
  MUX2_X1 U240 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n276), .Z(n218) );
  MUX2_X1 U241 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n276), .Z(n219) );
  MUX2_X1 U242 ( .A(n219), .B(n218), .S(n275), .Z(n220) );
  MUX2_X1 U243 ( .A(n220), .B(n15), .S(N12), .Z(N22) );
  MUX2_X1 U244 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n277), .Z(n221) );
  MUX2_X1 U245 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n277), .Z(n222) );
  MUX2_X1 U246 ( .A(n222), .B(n221), .S(n275), .Z(n223) );
  MUX2_X1 U247 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n277), .Z(n224) );
  MUX2_X1 U248 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n277), .Z(n225) );
  MUX2_X1 U249 ( .A(n225), .B(n224), .S(n275), .Z(n226) );
  MUX2_X1 U250 ( .A(n226), .B(n223), .S(N12), .Z(N21) );
  MUX2_X1 U251 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n277), .Z(n227) );
  MUX2_X1 U252 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n277), .Z(n228) );
  MUX2_X1 U253 ( .A(n228), .B(n227), .S(n275), .Z(n229) );
  MUX2_X1 U254 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n277), .Z(n230) );
  MUX2_X1 U255 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n277), .Z(n231) );
  MUX2_X1 U256 ( .A(n231), .B(n230), .S(n275), .Z(n232) );
  MUX2_X1 U257 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n277), .Z(n233) );
  MUX2_X1 U258 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n277), .Z(n234) );
  MUX2_X1 U259 ( .A(n234), .B(n233), .S(n275), .Z(n235) );
  MUX2_X1 U260 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n277), .Z(n236) );
  MUX2_X1 U261 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n277), .Z(n237) );
  MUX2_X1 U262 ( .A(n237), .B(n236), .S(n275), .Z(n238) );
  MUX2_X1 U263 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n277), .Z(n239) );
  MUX2_X1 U264 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n240) );
  MUX2_X1 U265 ( .A(n240), .B(n239), .S(n275), .Z(n241) );
  MUX2_X1 U266 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n242) );
  MUX2_X1 U267 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n243) );
  MUX2_X1 U268 ( .A(n243), .B(n242), .S(n275), .Z(n244) );
  MUX2_X1 U269 ( .A(n244), .B(n241), .S(N12), .Z(N18) );
  MUX2_X1 U270 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n245) );
  MUX2_X1 U271 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n277), .Z(n246) );
  MUX2_X1 U272 ( .A(n246), .B(n245), .S(n275), .Z(n247) );
  MUX2_X1 U273 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n277), .Z(n248) );
  MUX2_X1 U274 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n277), .Z(n249) );
  MUX2_X1 U275 ( .A(n249), .B(n248), .S(n275), .Z(n250) );
  MUX2_X1 U276 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n277), .Z(n251) );
  MUX2_X1 U277 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n277), .Z(n252) );
  MUX2_X1 U278 ( .A(n252), .B(n251), .S(n275), .Z(n253) );
  MUX2_X1 U279 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n277), .Z(n254) );
  MUX2_X1 U280 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n277), .Z(n255) );
  MUX2_X1 U281 ( .A(n255), .B(n254), .S(n275), .Z(n256) );
  MUX2_X1 U282 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(N10), .Z(n257) );
  MUX2_X1 U283 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(N10), .Z(n258) );
  MUX2_X1 U284 ( .A(n258), .B(n257), .S(n275), .Z(n259) );
  MUX2_X1 U285 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(N10), .Z(n260) );
  MUX2_X1 U286 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(N10), .Z(n261) );
  MUX2_X1 U287 ( .A(n261), .B(n260), .S(N11), .Z(n262) );
  MUX2_X1 U288 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(N10), .Z(n263) );
  MUX2_X1 U289 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(N10), .Z(n264) );
  MUX2_X1 U290 ( .A(n264), .B(n263), .S(n275), .Z(n265) );
  MUX2_X1 U291 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(N10), .Z(n266) );
  MUX2_X1 U292 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(N10), .Z(n267) );
  MUX2_X1 U293 ( .A(n267), .B(n266), .S(N11), .Z(n268) );
  MUX2_X1 U294 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(N10), .Z(n269) );
  MUX2_X1 U295 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n277), .Z(n270) );
  MUX2_X1 U296 ( .A(n270), .B(n269), .S(n275), .Z(n271) );
  MUX2_X1 U297 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(N10), .Z(n272) );
  MUX2_X1 U298 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(N10), .Z(n273) );
  MUX2_X1 U299 ( .A(n273), .B(n272), .S(n275), .Z(n274) );
  MUX2_X1 U300 ( .A(n274), .B(n271), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH12_SIZE8_LOGSIZE3_7 ( clk, data_in, data_out, addr, wr_en
 );
  input [11:0] data_in;
  output [11:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] ,
         \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] ,
         \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][11] , \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] ,
         \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] ,
         \mem[5][1] , \mem[5][0] , \mem[4][11] , \mem[4][10] , \mem[4][9] ,
         \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] ,
         \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] ,
         \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] ,
         \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][11] , \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] ,
         \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] ,
         \mem[0][1] , \mem[0][0] , N13, N14, N15, N20, N21, N22, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[11]  ( .D(N13), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N14), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N15), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[4]  ( .D(N20), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N21), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N22), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \mem_reg[7][11]  ( .D(n293), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n294), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n295), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n296), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n297), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n298), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n299), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n300), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n301), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n302), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n303), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n304), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n305), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n306), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n307), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n308), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n309), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n310), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n311), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n312), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n313), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n314), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n315), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n316), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n317), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n318), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n319), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n320), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n321), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n322), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n323), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n324), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n325), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n326), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n327), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n328), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n329), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n330), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n331), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n332), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n333), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n334), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n335), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n336), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n337), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n338), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n339), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n340), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n341), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n342), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n343), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n344), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n345), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n346), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n347), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n348), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n349), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n350), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n351), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n352), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n353), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n354), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n355), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n356), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n357), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n358), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n359), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n360), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n361), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n362), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n363), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n364), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n365), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n366), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n367), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n368), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n369), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n370), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n371), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n372), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n373), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n374), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n375), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n376), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n377), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n378), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n379), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n380), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n381), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n382), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n383), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n384), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n385), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n386), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n387), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n388), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U212 ( .A1(n278), .A2(n279), .A3(n481), .ZN(n494) );
  NAND3_X1 U213 ( .A1(n481), .A2(n279), .A3(N10), .ZN(n480) );
  NAND3_X1 U214 ( .A1(n481), .A2(n278), .A3(N11), .ZN(n467) );
  NAND3_X1 U215 ( .A1(N10), .A2(n481), .A3(N11), .ZN(n454) );
  NAND3_X1 U216 ( .A1(n278), .A2(n279), .A3(n428), .ZN(n441) );
  NAND3_X1 U217 ( .A1(N10), .A2(n279), .A3(n428), .ZN(n427) );
  NAND3_X1 U218 ( .A1(N11), .A2(n278), .A3(n428), .ZN(n414) );
  NAND3_X1 U219 ( .A1(N11), .A2(N10), .A3(n428), .ZN(n401) );
  SDFF_X1 \data_out_reg[5]  ( .D(n238), .SI(n235), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n250), .SI(n247), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n12), .SI(n9), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[8]  ( .D(n256), .SI(n253), .SE(N12), .CK(clk), .Q(
        data_out[8]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n6), .SI(n3), .SE(N12), .CK(clk), .Q(
        data_out[0]) );
  SDFF_X1 \data_out_reg[6]  ( .D(n244), .SI(n241), .SE(N12), .CK(clk), .Q(
        data_out[6]) );
  BUF_X1 U3 ( .A(n277), .Z(n276) );
  BUF_X1 U4 ( .A(N11), .Z(n275) );
  BUF_X1 U5 ( .A(N10), .Z(n277) );
  AND2_X1 U6 ( .A1(N12), .A2(wr_en), .ZN(n428) );
  INV_X1 U7 ( .A(N10), .ZN(n278) );
  INV_X1 U8 ( .A(N11), .ZN(n279) );
  OAI21_X1 U9 ( .B1(n292), .B2(n480), .A(n479), .ZN(n376) );
  NAND2_X1 U10 ( .A1(\mem[1][0] ), .A2(n480), .ZN(n479) );
  OAI21_X1 U11 ( .B1(n291), .B2(n480), .A(n478), .ZN(n375) );
  NAND2_X1 U12 ( .A1(\mem[1][1] ), .A2(n480), .ZN(n478) );
  OAI21_X1 U13 ( .B1(n290), .B2(n480), .A(n477), .ZN(n374) );
  NAND2_X1 U14 ( .A1(\mem[1][2] ), .A2(n480), .ZN(n477) );
  OAI21_X1 U15 ( .B1(n289), .B2(n480), .A(n476), .ZN(n373) );
  NAND2_X1 U16 ( .A1(\mem[1][3] ), .A2(n480), .ZN(n476) );
  OAI21_X1 U17 ( .B1(n288), .B2(n480), .A(n475), .ZN(n372) );
  NAND2_X1 U18 ( .A1(\mem[1][4] ), .A2(n480), .ZN(n475) );
  OAI21_X1 U19 ( .B1(n287), .B2(n480), .A(n474), .ZN(n371) );
  NAND2_X1 U20 ( .A1(\mem[1][5] ), .A2(n480), .ZN(n474) );
  OAI21_X1 U21 ( .B1(n286), .B2(n480), .A(n473), .ZN(n370) );
  NAND2_X1 U22 ( .A1(\mem[1][6] ), .A2(n480), .ZN(n473) );
  OAI21_X1 U23 ( .B1(n285), .B2(n480), .A(n472), .ZN(n369) );
  NAND2_X1 U24 ( .A1(\mem[1][7] ), .A2(n480), .ZN(n472) );
  OAI21_X1 U25 ( .B1(n284), .B2(n480), .A(n471), .ZN(n368) );
  NAND2_X1 U26 ( .A1(\mem[1][8] ), .A2(n480), .ZN(n471) );
  OAI21_X1 U27 ( .B1(n283), .B2(n480), .A(n470), .ZN(n367) );
  NAND2_X1 U28 ( .A1(\mem[1][9] ), .A2(n480), .ZN(n470) );
  OAI21_X1 U29 ( .B1(n282), .B2(n480), .A(n469), .ZN(n366) );
  NAND2_X1 U30 ( .A1(\mem[1][10] ), .A2(n480), .ZN(n469) );
  OAI21_X1 U31 ( .B1(n281), .B2(n480), .A(n468), .ZN(n365) );
  NAND2_X1 U32 ( .A1(\mem[1][11] ), .A2(n480), .ZN(n468) );
  OAI21_X1 U33 ( .B1(n292), .B2(n467), .A(n466), .ZN(n364) );
  NAND2_X1 U34 ( .A1(\mem[2][0] ), .A2(n467), .ZN(n466) );
  OAI21_X1 U35 ( .B1(n291), .B2(n467), .A(n465), .ZN(n363) );
  NAND2_X1 U36 ( .A1(\mem[2][1] ), .A2(n467), .ZN(n465) );
  OAI21_X1 U37 ( .B1(n290), .B2(n467), .A(n464), .ZN(n362) );
  NAND2_X1 U38 ( .A1(\mem[2][2] ), .A2(n467), .ZN(n464) );
  OAI21_X1 U39 ( .B1(n289), .B2(n467), .A(n463), .ZN(n361) );
  NAND2_X1 U40 ( .A1(\mem[2][3] ), .A2(n467), .ZN(n463) );
  OAI21_X1 U41 ( .B1(n288), .B2(n467), .A(n462), .ZN(n360) );
  NAND2_X1 U42 ( .A1(\mem[2][4] ), .A2(n467), .ZN(n462) );
  OAI21_X1 U43 ( .B1(n287), .B2(n467), .A(n461), .ZN(n359) );
  NAND2_X1 U44 ( .A1(\mem[2][5] ), .A2(n467), .ZN(n461) );
  OAI21_X1 U45 ( .B1(n286), .B2(n467), .A(n460), .ZN(n358) );
  NAND2_X1 U46 ( .A1(\mem[2][6] ), .A2(n467), .ZN(n460) );
  OAI21_X1 U47 ( .B1(n285), .B2(n467), .A(n459), .ZN(n357) );
  NAND2_X1 U48 ( .A1(\mem[2][7] ), .A2(n467), .ZN(n459) );
  OAI21_X1 U49 ( .B1(n284), .B2(n467), .A(n458), .ZN(n356) );
  NAND2_X1 U50 ( .A1(\mem[2][8] ), .A2(n467), .ZN(n458) );
  OAI21_X1 U51 ( .B1(n283), .B2(n467), .A(n457), .ZN(n355) );
  NAND2_X1 U52 ( .A1(\mem[2][9] ), .A2(n467), .ZN(n457) );
  OAI21_X1 U53 ( .B1(n282), .B2(n467), .A(n456), .ZN(n354) );
  NAND2_X1 U54 ( .A1(\mem[2][10] ), .A2(n467), .ZN(n456) );
  OAI21_X1 U55 ( .B1(n281), .B2(n467), .A(n455), .ZN(n353) );
  NAND2_X1 U56 ( .A1(\mem[2][11] ), .A2(n467), .ZN(n455) );
  OAI21_X1 U57 ( .B1(n292), .B2(n454), .A(n453), .ZN(n352) );
  NAND2_X1 U58 ( .A1(\mem[3][0] ), .A2(n454), .ZN(n453) );
  OAI21_X1 U59 ( .B1(n291), .B2(n454), .A(n452), .ZN(n351) );
  NAND2_X1 U60 ( .A1(\mem[3][1] ), .A2(n454), .ZN(n452) );
  OAI21_X1 U61 ( .B1(n290), .B2(n454), .A(n451), .ZN(n350) );
  NAND2_X1 U62 ( .A1(\mem[3][2] ), .A2(n454), .ZN(n451) );
  OAI21_X1 U63 ( .B1(n289), .B2(n454), .A(n450), .ZN(n349) );
  NAND2_X1 U64 ( .A1(\mem[3][3] ), .A2(n454), .ZN(n450) );
  OAI21_X1 U65 ( .B1(n288), .B2(n454), .A(n449), .ZN(n348) );
  NAND2_X1 U66 ( .A1(\mem[3][4] ), .A2(n454), .ZN(n449) );
  OAI21_X1 U67 ( .B1(n287), .B2(n454), .A(n448), .ZN(n347) );
  NAND2_X1 U68 ( .A1(\mem[3][5] ), .A2(n454), .ZN(n448) );
  OAI21_X1 U69 ( .B1(n286), .B2(n454), .A(n447), .ZN(n346) );
  NAND2_X1 U70 ( .A1(\mem[3][6] ), .A2(n454), .ZN(n447) );
  OAI21_X1 U71 ( .B1(n285), .B2(n454), .A(n446), .ZN(n345) );
  NAND2_X1 U72 ( .A1(\mem[3][7] ), .A2(n454), .ZN(n446) );
  OAI21_X1 U73 ( .B1(n284), .B2(n454), .A(n445), .ZN(n344) );
  NAND2_X1 U74 ( .A1(\mem[3][8] ), .A2(n454), .ZN(n445) );
  OAI21_X1 U75 ( .B1(n283), .B2(n454), .A(n444), .ZN(n343) );
  NAND2_X1 U76 ( .A1(\mem[3][9] ), .A2(n454), .ZN(n444) );
  OAI21_X1 U77 ( .B1(n282), .B2(n454), .A(n443), .ZN(n342) );
  NAND2_X1 U78 ( .A1(\mem[3][10] ), .A2(n454), .ZN(n443) );
  OAI21_X1 U79 ( .B1(n281), .B2(n454), .A(n442), .ZN(n341) );
  NAND2_X1 U80 ( .A1(\mem[3][11] ), .A2(n454), .ZN(n442) );
  OAI21_X1 U81 ( .B1(n292), .B2(n441), .A(n440), .ZN(n340) );
  NAND2_X1 U82 ( .A1(\mem[4][0] ), .A2(n441), .ZN(n440) );
  OAI21_X1 U83 ( .B1(n291), .B2(n441), .A(n439), .ZN(n339) );
  NAND2_X1 U84 ( .A1(\mem[4][1] ), .A2(n441), .ZN(n439) );
  OAI21_X1 U85 ( .B1(n290), .B2(n441), .A(n438), .ZN(n338) );
  NAND2_X1 U86 ( .A1(\mem[4][2] ), .A2(n441), .ZN(n438) );
  OAI21_X1 U87 ( .B1(n289), .B2(n441), .A(n437), .ZN(n337) );
  NAND2_X1 U88 ( .A1(\mem[4][3] ), .A2(n441), .ZN(n437) );
  OAI21_X1 U89 ( .B1(n288), .B2(n441), .A(n436), .ZN(n336) );
  NAND2_X1 U90 ( .A1(\mem[4][4] ), .A2(n441), .ZN(n436) );
  OAI21_X1 U91 ( .B1(n287), .B2(n441), .A(n435), .ZN(n335) );
  NAND2_X1 U92 ( .A1(\mem[4][5] ), .A2(n441), .ZN(n435) );
  OAI21_X1 U93 ( .B1(n286), .B2(n441), .A(n434), .ZN(n334) );
  NAND2_X1 U94 ( .A1(\mem[4][6] ), .A2(n441), .ZN(n434) );
  OAI21_X1 U95 ( .B1(n285), .B2(n441), .A(n433), .ZN(n333) );
  NAND2_X1 U96 ( .A1(\mem[4][7] ), .A2(n441), .ZN(n433) );
  OAI21_X1 U97 ( .B1(n284), .B2(n441), .A(n432), .ZN(n332) );
  NAND2_X1 U98 ( .A1(\mem[4][8] ), .A2(n441), .ZN(n432) );
  OAI21_X1 U99 ( .B1(n283), .B2(n441), .A(n431), .ZN(n331) );
  NAND2_X1 U100 ( .A1(\mem[4][9] ), .A2(n441), .ZN(n431) );
  OAI21_X1 U101 ( .B1(n282), .B2(n441), .A(n430), .ZN(n330) );
  NAND2_X1 U102 ( .A1(\mem[4][10] ), .A2(n441), .ZN(n430) );
  OAI21_X1 U103 ( .B1(n281), .B2(n441), .A(n429), .ZN(n329) );
  NAND2_X1 U104 ( .A1(\mem[4][11] ), .A2(n441), .ZN(n429) );
  OAI21_X1 U105 ( .B1(n292), .B2(n427), .A(n426), .ZN(n328) );
  NAND2_X1 U106 ( .A1(\mem[5][0] ), .A2(n427), .ZN(n426) );
  OAI21_X1 U107 ( .B1(n291), .B2(n427), .A(n425), .ZN(n327) );
  NAND2_X1 U108 ( .A1(\mem[5][1] ), .A2(n427), .ZN(n425) );
  OAI21_X1 U109 ( .B1(n290), .B2(n427), .A(n424), .ZN(n326) );
  NAND2_X1 U110 ( .A1(\mem[5][2] ), .A2(n427), .ZN(n424) );
  OAI21_X1 U111 ( .B1(n289), .B2(n427), .A(n423), .ZN(n325) );
  NAND2_X1 U112 ( .A1(\mem[5][3] ), .A2(n427), .ZN(n423) );
  OAI21_X1 U113 ( .B1(n288), .B2(n427), .A(n422), .ZN(n324) );
  NAND2_X1 U114 ( .A1(\mem[5][4] ), .A2(n427), .ZN(n422) );
  OAI21_X1 U115 ( .B1(n287), .B2(n427), .A(n421), .ZN(n323) );
  NAND2_X1 U116 ( .A1(\mem[5][5] ), .A2(n427), .ZN(n421) );
  OAI21_X1 U117 ( .B1(n286), .B2(n427), .A(n420), .ZN(n322) );
  NAND2_X1 U118 ( .A1(\mem[5][6] ), .A2(n427), .ZN(n420) );
  OAI21_X1 U119 ( .B1(n285), .B2(n427), .A(n419), .ZN(n321) );
  NAND2_X1 U120 ( .A1(\mem[5][7] ), .A2(n427), .ZN(n419) );
  OAI21_X1 U121 ( .B1(n284), .B2(n427), .A(n418), .ZN(n320) );
  NAND2_X1 U122 ( .A1(\mem[5][8] ), .A2(n427), .ZN(n418) );
  OAI21_X1 U123 ( .B1(n283), .B2(n427), .A(n417), .ZN(n319) );
  NAND2_X1 U124 ( .A1(\mem[5][9] ), .A2(n427), .ZN(n417) );
  OAI21_X1 U125 ( .B1(n282), .B2(n427), .A(n416), .ZN(n318) );
  NAND2_X1 U126 ( .A1(\mem[5][10] ), .A2(n427), .ZN(n416) );
  OAI21_X1 U127 ( .B1(n281), .B2(n427), .A(n415), .ZN(n317) );
  NAND2_X1 U128 ( .A1(\mem[5][11] ), .A2(n427), .ZN(n415) );
  OAI21_X1 U129 ( .B1(n292), .B2(n414), .A(n413), .ZN(n316) );
  NAND2_X1 U130 ( .A1(\mem[6][0] ), .A2(n414), .ZN(n413) );
  OAI21_X1 U131 ( .B1(n291), .B2(n414), .A(n412), .ZN(n315) );
  NAND2_X1 U132 ( .A1(\mem[6][1] ), .A2(n414), .ZN(n412) );
  OAI21_X1 U133 ( .B1(n290), .B2(n414), .A(n411), .ZN(n314) );
  NAND2_X1 U134 ( .A1(\mem[6][2] ), .A2(n414), .ZN(n411) );
  OAI21_X1 U135 ( .B1(n289), .B2(n414), .A(n410), .ZN(n313) );
  NAND2_X1 U136 ( .A1(\mem[6][3] ), .A2(n414), .ZN(n410) );
  OAI21_X1 U137 ( .B1(n288), .B2(n414), .A(n409), .ZN(n312) );
  NAND2_X1 U138 ( .A1(\mem[6][4] ), .A2(n414), .ZN(n409) );
  OAI21_X1 U139 ( .B1(n287), .B2(n414), .A(n408), .ZN(n311) );
  NAND2_X1 U140 ( .A1(\mem[6][5] ), .A2(n414), .ZN(n408) );
  OAI21_X1 U141 ( .B1(n286), .B2(n414), .A(n407), .ZN(n310) );
  NAND2_X1 U142 ( .A1(\mem[6][6] ), .A2(n414), .ZN(n407) );
  OAI21_X1 U143 ( .B1(n285), .B2(n414), .A(n406), .ZN(n309) );
  NAND2_X1 U144 ( .A1(\mem[6][7] ), .A2(n414), .ZN(n406) );
  OAI21_X1 U145 ( .B1(n284), .B2(n414), .A(n405), .ZN(n308) );
  NAND2_X1 U146 ( .A1(\mem[6][8] ), .A2(n414), .ZN(n405) );
  OAI21_X1 U147 ( .B1(n283), .B2(n414), .A(n404), .ZN(n307) );
  NAND2_X1 U148 ( .A1(\mem[6][9] ), .A2(n414), .ZN(n404) );
  OAI21_X1 U149 ( .B1(n282), .B2(n414), .A(n403), .ZN(n306) );
  NAND2_X1 U150 ( .A1(\mem[6][10] ), .A2(n414), .ZN(n403) );
  OAI21_X1 U151 ( .B1(n281), .B2(n414), .A(n402), .ZN(n305) );
  NAND2_X1 U152 ( .A1(\mem[6][11] ), .A2(n414), .ZN(n402) );
  OAI21_X1 U153 ( .B1(n292), .B2(n401), .A(n400), .ZN(n304) );
  NAND2_X1 U154 ( .A1(\mem[7][0] ), .A2(n401), .ZN(n400) );
  OAI21_X1 U155 ( .B1(n291), .B2(n401), .A(n399), .ZN(n303) );
  NAND2_X1 U156 ( .A1(\mem[7][1] ), .A2(n401), .ZN(n399) );
  OAI21_X1 U157 ( .B1(n290), .B2(n401), .A(n398), .ZN(n302) );
  NAND2_X1 U158 ( .A1(\mem[7][2] ), .A2(n401), .ZN(n398) );
  OAI21_X1 U159 ( .B1(n289), .B2(n401), .A(n397), .ZN(n301) );
  NAND2_X1 U160 ( .A1(\mem[7][3] ), .A2(n401), .ZN(n397) );
  OAI21_X1 U161 ( .B1(n288), .B2(n401), .A(n396), .ZN(n300) );
  NAND2_X1 U162 ( .A1(\mem[7][4] ), .A2(n401), .ZN(n396) );
  OAI21_X1 U163 ( .B1(n287), .B2(n401), .A(n395), .ZN(n299) );
  NAND2_X1 U164 ( .A1(\mem[7][5] ), .A2(n401), .ZN(n395) );
  OAI21_X1 U165 ( .B1(n286), .B2(n401), .A(n394), .ZN(n298) );
  NAND2_X1 U166 ( .A1(\mem[7][6] ), .A2(n401), .ZN(n394) );
  OAI21_X1 U167 ( .B1(n285), .B2(n401), .A(n393), .ZN(n297) );
  NAND2_X1 U168 ( .A1(\mem[7][7] ), .A2(n401), .ZN(n393) );
  OAI21_X1 U169 ( .B1(n284), .B2(n401), .A(n392), .ZN(n296) );
  NAND2_X1 U170 ( .A1(\mem[7][8] ), .A2(n401), .ZN(n392) );
  OAI21_X1 U171 ( .B1(n283), .B2(n401), .A(n391), .ZN(n295) );
  NAND2_X1 U172 ( .A1(\mem[7][9] ), .A2(n401), .ZN(n391) );
  OAI21_X1 U173 ( .B1(n282), .B2(n401), .A(n390), .ZN(n294) );
  NAND2_X1 U174 ( .A1(\mem[7][10] ), .A2(n401), .ZN(n390) );
  OAI21_X1 U175 ( .B1(n281), .B2(n401), .A(n389), .ZN(n293) );
  NAND2_X1 U176 ( .A1(\mem[7][11] ), .A2(n401), .ZN(n389) );
  OAI21_X1 U177 ( .B1(n494), .B2(n292), .A(n493), .ZN(n388) );
  NAND2_X1 U178 ( .A1(\mem[0][0] ), .A2(n494), .ZN(n493) );
  OAI21_X1 U179 ( .B1(n494), .B2(n291), .A(n492), .ZN(n387) );
  NAND2_X1 U180 ( .A1(\mem[0][1] ), .A2(n494), .ZN(n492) );
  OAI21_X1 U181 ( .B1(n494), .B2(n290), .A(n491), .ZN(n386) );
  NAND2_X1 U182 ( .A1(\mem[0][2] ), .A2(n494), .ZN(n491) );
  OAI21_X1 U183 ( .B1(n494), .B2(n289), .A(n490), .ZN(n385) );
  NAND2_X1 U184 ( .A1(\mem[0][3] ), .A2(n494), .ZN(n490) );
  OAI21_X1 U185 ( .B1(n494), .B2(n288), .A(n489), .ZN(n384) );
  NAND2_X1 U186 ( .A1(\mem[0][4] ), .A2(n494), .ZN(n489) );
  OAI21_X1 U187 ( .B1(n494), .B2(n287), .A(n488), .ZN(n383) );
  NAND2_X1 U188 ( .A1(\mem[0][5] ), .A2(n494), .ZN(n488) );
  OAI21_X1 U189 ( .B1(n494), .B2(n286), .A(n487), .ZN(n382) );
  NAND2_X1 U190 ( .A1(\mem[0][6] ), .A2(n494), .ZN(n487) );
  OAI21_X1 U191 ( .B1(n494), .B2(n285), .A(n486), .ZN(n381) );
  NAND2_X1 U192 ( .A1(\mem[0][7] ), .A2(n494), .ZN(n486) );
  OAI21_X1 U193 ( .B1(n494), .B2(n284), .A(n485), .ZN(n380) );
  NAND2_X1 U194 ( .A1(\mem[0][8] ), .A2(n494), .ZN(n485) );
  OAI21_X1 U195 ( .B1(n494), .B2(n283), .A(n484), .ZN(n379) );
  NAND2_X1 U196 ( .A1(\mem[0][9] ), .A2(n494), .ZN(n484) );
  OAI21_X1 U197 ( .B1(n494), .B2(n282), .A(n483), .ZN(n378) );
  NAND2_X1 U198 ( .A1(\mem[0][10] ), .A2(n494), .ZN(n483) );
  OAI21_X1 U199 ( .B1(n494), .B2(n281), .A(n482), .ZN(n377) );
  NAND2_X1 U200 ( .A1(\mem[0][11] ), .A2(n494), .ZN(n482) );
  NOR2_X1 U201 ( .A1(n280), .A2(N12), .ZN(n481) );
  INV_X1 U202 ( .A(wr_en), .ZN(n280) );
  INV_X1 U203 ( .A(data_in[0]), .ZN(n292) );
  INV_X1 U204 ( .A(data_in[1]), .ZN(n291) );
  INV_X1 U205 ( .A(data_in[2]), .ZN(n290) );
  INV_X1 U206 ( .A(data_in[3]), .ZN(n289) );
  INV_X1 U207 ( .A(data_in[4]), .ZN(n288) );
  INV_X1 U208 ( .A(data_in[5]), .ZN(n287) );
  INV_X1 U209 ( .A(data_in[6]), .ZN(n286) );
  INV_X1 U210 ( .A(data_in[7]), .ZN(n285) );
  INV_X1 U211 ( .A(data_in[8]), .ZN(n284) );
  INV_X1 U220 ( .A(data_in[9]), .ZN(n283) );
  INV_X1 U221 ( .A(data_in[10]), .ZN(n282) );
  INV_X1 U222 ( .A(data_in[11]), .ZN(n281) );
  MUX2_X1 U223 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n276), .Z(n1) );
  MUX2_X1 U224 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n276), .Z(n2) );
  MUX2_X1 U225 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U226 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n276), .Z(n4) );
  MUX2_X1 U227 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n276), .Z(n5) );
  MUX2_X1 U228 ( .A(n5), .B(n4), .S(N11), .Z(n6) );
  MUX2_X1 U229 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n276), .Z(n7) );
  MUX2_X1 U230 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n276), .Z(n8) );
  MUX2_X1 U231 ( .A(n8), .B(n7), .S(N11), .Z(n9) );
  MUX2_X1 U232 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n276), .Z(n10) );
  MUX2_X1 U233 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n276), .Z(n11) );
  MUX2_X1 U234 ( .A(n11), .B(n10), .S(N11), .Z(n12) );
  MUX2_X1 U235 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n276), .Z(n13) );
  MUX2_X1 U236 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n276), .Z(n14) );
  MUX2_X1 U237 ( .A(n14), .B(n13), .S(N11), .Z(n15) );
  MUX2_X1 U238 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n276), .Z(n218) );
  MUX2_X1 U239 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n276), .Z(n219) );
  MUX2_X1 U240 ( .A(n219), .B(n218), .S(N11), .Z(n220) );
  MUX2_X1 U241 ( .A(n220), .B(n15), .S(N12), .Z(N22) );
  MUX2_X1 U242 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n277), .Z(n221) );
  MUX2_X1 U243 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n277), .Z(n222) );
  MUX2_X1 U244 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U245 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n277), .Z(n224) );
  MUX2_X1 U246 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n277), .Z(n225) );
  MUX2_X1 U247 ( .A(n225), .B(n224), .S(N11), .Z(n226) );
  MUX2_X1 U248 ( .A(n226), .B(n223), .S(N12), .Z(N21) );
  MUX2_X1 U249 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n277), .Z(n227) );
  MUX2_X1 U250 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n277), .Z(n228) );
  MUX2_X1 U251 ( .A(n228), .B(n227), .S(N11), .Z(n229) );
  MUX2_X1 U252 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n277), .Z(n230) );
  MUX2_X1 U253 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n277), .Z(n231) );
  MUX2_X1 U254 ( .A(n231), .B(n230), .S(N11), .Z(n232) );
  MUX2_X1 U255 ( .A(n232), .B(n229), .S(N12), .Z(N20) );
  MUX2_X1 U256 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n277), .Z(n233) );
  MUX2_X1 U257 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n277), .Z(n234) );
  MUX2_X1 U258 ( .A(n234), .B(n233), .S(N11), .Z(n235) );
  MUX2_X1 U259 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n277), .Z(n236) );
  MUX2_X1 U260 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n277), .Z(n237) );
  MUX2_X1 U261 ( .A(n237), .B(n236), .S(N11), .Z(n238) );
  MUX2_X1 U262 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n239) );
  MUX2_X1 U263 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n240) );
  MUX2_X1 U264 ( .A(n240), .B(n239), .S(n275), .Z(n241) );
  MUX2_X1 U265 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n277), .Z(n242) );
  MUX2_X1 U266 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n277), .Z(n243) );
  MUX2_X1 U267 ( .A(n243), .B(n242), .S(n275), .Z(n244) );
  MUX2_X1 U268 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n245) );
  MUX2_X1 U269 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n246) );
  MUX2_X1 U270 ( .A(n246), .B(n245), .S(n275), .Z(n247) );
  MUX2_X1 U271 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n277), .Z(n248) );
  MUX2_X1 U272 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n277), .Z(n249) );
  MUX2_X1 U273 ( .A(n249), .B(n248), .S(n275), .Z(n250) );
  MUX2_X1 U274 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(N10), .Z(n251) );
  MUX2_X1 U275 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n277), .Z(n252) );
  MUX2_X1 U276 ( .A(n252), .B(n251), .S(n275), .Z(n253) );
  MUX2_X1 U277 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n277), .Z(n254) );
  MUX2_X1 U278 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n277), .Z(n255) );
  MUX2_X1 U279 ( .A(n255), .B(n254), .S(n275), .Z(n256) );
  MUX2_X1 U280 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n277), .Z(n257) );
  MUX2_X1 U281 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(N10), .Z(n258) );
  MUX2_X1 U282 ( .A(n258), .B(n257), .S(n275), .Z(n259) );
  MUX2_X1 U283 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(N10), .Z(n260) );
  MUX2_X1 U284 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(N10), .Z(n261) );
  MUX2_X1 U285 ( .A(n261), .B(n260), .S(n275), .Z(n262) );
  MUX2_X1 U286 ( .A(n262), .B(n259), .S(N12), .Z(N15) );
  MUX2_X1 U287 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(N10), .Z(n263) );
  MUX2_X1 U288 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(N10), .Z(n264) );
  MUX2_X1 U289 ( .A(n264), .B(n263), .S(n275), .Z(n265) );
  MUX2_X1 U290 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(N10), .Z(n266) );
  MUX2_X1 U291 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(N10), .Z(n267) );
  MUX2_X1 U292 ( .A(n267), .B(n266), .S(n275), .Z(n268) );
  MUX2_X1 U293 ( .A(n268), .B(n265), .S(N12), .Z(N14) );
  MUX2_X1 U294 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(N10), .Z(n269) );
  MUX2_X1 U295 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(N10), .Z(n270) );
  MUX2_X1 U296 ( .A(n270), .B(n269), .S(n275), .Z(n271) );
  MUX2_X1 U297 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n277), .Z(n272) );
  MUX2_X1 U298 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(N10), .Z(n273) );
  MUX2_X1 U299 ( .A(n273), .B(n272), .S(n275), .Z(n274) );
  MUX2_X1 U300 ( .A(n274), .B(n271), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH12_SIZE8_LOGSIZE3_6 ( clk, data_in, data_out, addr, wr_en
 );
  input [11:0] data_in;
  output [11:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] ,
         \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] ,
         \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][11] , \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] ,
         \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] ,
         \mem[5][1] , \mem[5][0] , \mem[4][11] , \mem[4][10] , \mem[4][9] ,
         \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] ,
         \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] ,
         \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] ,
         \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][11] , \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] ,
         \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] ,
         \mem[0][1] , \mem[0][0] , N14, N18, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[10]  ( .D(N14), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[6]  ( .D(N18), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \mem_reg[7][11]  ( .D(n293), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n294), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n295), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n296), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n297), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n298), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n299), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n300), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n301), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n302), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n303), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n304), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n305), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n306), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n307), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n308), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n309), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n310), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n311), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n312), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n313), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n314), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n315), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n316), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n317), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n318), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n319), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n320), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n321), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n322), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n323), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n324), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n325), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n326), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n327), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n328), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n329), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n330), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n331), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n332), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n333), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n334), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n335), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n336), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n337), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n338), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n339), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n340), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n341), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n342), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n343), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n344), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n345), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n346), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n347), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n348), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n349), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n350), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n351), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n352), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n353), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n354), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n355), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n356), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n357), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n358), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n359), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n360), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n361), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n362), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n363), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n364), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n365), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n366), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n367), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n368), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n369), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n370), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n371), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n372), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n373), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n374), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n375), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n376), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n377), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n378), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n379), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n380), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n381), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n382), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n383), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n384), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n385), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n386), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n387), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n388), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U212 ( .A1(n278), .A2(n279), .A3(n481), .ZN(n494) );
  NAND3_X1 U213 ( .A1(n481), .A2(n279), .A3(N10), .ZN(n480) );
  NAND3_X1 U214 ( .A1(n481), .A2(n278), .A3(N11), .ZN(n467) );
  NAND3_X1 U215 ( .A1(N10), .A2(n481), .A3(N11), .ZN(n454) );
  NAND3_X1 U216 ( .A1(n278), .A2(n279), .A3(n428), .ZN(n441) );
  NAND3_X1 U217 ( .A1(N10), .A2(n279), .A3(n428), .ZN(n427) );
  NAND3_X1 U218 ( .A1(N11), .A2(n278), .A3(n428), .ZN(n414) );
  NAND3_X1 U219 ( .A1(N11), .A2(N10), .A3(n428), .ZN(n401) );
  SDFF_X1 \data_out_reg[5]  ( .D(n238), .SI(n235), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n262), .SI(n259), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n12), .SI(n9), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n250), .SI(n247), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n226), .SI(n223), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[4]  ( .D(n232), .SI(n229), .SE(N12), .CK(clk), .Q(
        data_out[4]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n274), .SI(n271), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[8]  ( .D(n256), .SI(n253), .SE(N12), .CK(clk), .Q(
        data_out[8]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n6), .SI(n3), .SE(N12), .CK(clk), .Q(
        data_out[0]) );
  SDFF_X1 \data_out_reg[2]  ( .D(n220), .SI(n15), .SE(N12), .CK(clk), .Q(
        data_out[2]) );
  BUF_X1 U3 ( .A(n277), .Z(n276) );
  BUF_X1 U4 ( .A(N11), .Z(n275) );
  BUF_X1 U5 ( .A(N10), .Z(n277) );
  NOR2_X1 U6 ( .A1(n280), .A2(N12), .ZN(n481) );
  INV_X1 U7 ( .A(wr_en), .ZN(n280) );
  AND2_X1 U8 ( .A1(N12), .A2(wr_en), .ZN(n428) );
  INV_X1 U9 ( .A(N10), .ZN(n278) );
  INV_X1 U10 ( .A(N11), .ZN(n279) );
  OAI21_X1 U11 ( .B1(n292), .B2(n480), .A(n479), .ZN(n376) );
  NAND2_X1 U12 ( .A1(\mem[1][0] ), .A2(n480), .ZN(n479) );
  OAI21_X1 U13 ( .B1(n291), .B2(n480), .A(n478), .ZN(n375) );
  NAND2_X1 U14 ( .A1(\mem[1][1] ), .A2(n480), .ZN(n478) );
  OAI21_X1 U15 ( .B1(n290), .B2(n480), .A(n477), .ZN(n374) );
  NAND2_X1 U16 ( .A1(\mem[1][2] ), .A2(n480), .ZN(n477) );
  OAI21_X1 U17 ( .B1(n289), .B2(n480), .A(n476), .ZN(n373) );
  NAND2_X1 U18 ( .A1(\mem[1][3] ), .A2(n480), .ZN(n476) );
  OAI21_X1 U19 ( .B1(n288), .B2(n480), .A(n475), .ZN(n372) );
  NAND2_X1 U20 ( .A1(\mem[1][4] ), .A2(n480), .ZN(n475) );
  OAI21_X1 U21 ( .B1(n287), .B2(n480), .A(n474), .ZN(n371) );
  NAND2_X1 U22 ( .A1(\mem[1][5] ), .A2(n480), .ZN(n474) );
  OAI21_X1 U23 ( .B1(n286), .B2(n480), .A(n473), .ZN(n370) );
  NAND2_X1 U24 ( .A1(\mem[1][6] ), .A2(n480), .ZN(n473) );
  OAI21_X1 U25 ( .B1(n285), .B2(n480), .A(n472), .ZN(n369) );
  NAND2_X1 U26 ( .A1(\mem[1][7] ), .A2(n480), .ZN(n472) );
  OAI21_X1 U27 ( .B1(n284), .B2(n480), .A(n471), .ZN(n368) );
  NAND2_X1 U28 ( .A1(\mem[1][8] ), .A2(n480), .ZN(n471) );
  OAI21_X1 U29 ( .B1(n283), .B2(n480), .A(n470), .ZN(n367) );
  NAND2_X1 U30 ( .A1(\mem[1][9] ), .A2(n480), .ZN(n470) );
  OAI21_X1 U31 ( .B1(n282), .B2(n480), .A(n469), .ZN(n366) );
  NAND2_X1 U32 ( .A1(\mem[1][10] ), .A2(n480), .ZN(n469) );
  OAI21_X1 U33 ( .B1(n281), .B2(n480), .A(n468), .ZN(n365) );
  NAND2_X1 U34 ( .A1(\mem[1][11] ), .A2(n480), .ZN(n468) );
  OAI21_X1 U35 ( .B1(n292), .B2(n467), .A(n466), .ZN(n364) );
  NAND2_X1 U36 ( .A1(\mem[2][0] ), .A2(n467), .ZN(n466) );
  OAI21_X1 U37 ( .B1(n291), .B2(n467), .A(n465), .ZN(n363) );
  NAND2_X1 U38 ( .A1(\mem[2][1] ), .A2(n467), .ZN(n465) );
  OAI21_X1 U39 ( .B1(n290), .B2(n467), .A(n464), .ZN(n362) );
  NAND2_X1 U40 ( .A1(\mem[2][2] ), .A2(n467), .ZN(n464) );
  OAI21_X1 U41 ( .B1(n289), .B2(n467), .A(n463), .ZN(n361) );
  NAND2_X1 U42 ( .A1(\mem[2][3] ), .A2(n467), .ZN(n463) );
  OAI21_X1 U43 ( .B1(n288), .B2(n467), .A(n462), .ZN(n360) );
  NAND2_X1 U44 ( .A1(\mem[2][4] ), .A2(n467), .ZN(n462) );
  OAI21_X1 U45 ( .B1(n287), .B2(n467), .A(n461), .ZN(n359) );
  NAND2_X1 U46 ( .A1(\mem[2][5] ), .A2(n467), .ZN(n461) );
  OAI21_X1 U47 ( .B1(n286), .B2(n467), .A(n460), .ZN(n358) );
  NAND2_X1 U48 ( .A1(\mem[2][6] ), .A2(n467), .ZN(n460) );
  OAI21_X1 U49 ( .B1(n285), .B2(n467), .A(n459), .ZN(n357) );
  NAND2_X1 U50 ( .A1(\mem[2][7] ), .A2(n467), .ZN(n459) );
  OAI21_X1 U51 ( .B1(n284), .B2(n467), .A(n458), .ZN(n356) );
  NAND2_X1 U52 ( .A1(\mem[2][8] ), .A2(n467), .ZN(n458) );
  OAI21_X1 U53 ( .B1(n283), .B2(n467), .A(n457), .ZN(n355) );
  NAND2_X1 U54 ( .A1(\mem[2][9] ), .A2(n467), .ZN(n457) );
  OAI21_X1 U55 ( .B1(n282), .B2(n467), .A(n456), .ZN(n354) );
  NAND2_X1 U56 ( .A1(\mem[2][10] ), .A2(n467), .ZN(n456) );
  OAI21_X1 U57 ( .B1(n281), .B2(n467), .A(n455), .ZN(n353) );
  NAND2_X1 U58 ( .A1(\mem[2][11] ), .A2(n467), .ZN(n455) );
  OAI21_X1 U59 ( .B1(n292), .B2(n454), .A(n453), .ZN(n352) );
  NAND2_X1 U60 ( .A1(\mem[3][0] ), .A2(n454), .ZN(n453) );
  OAI21_X1 U61 ( .B1(n291), .B2(n454), .A(n452), .ZN(n351) );
  NAND2_X1 U62 ( .A1(\mem[3][1] ), .A2(n454), .ZN(n452) );
  OAI21_X1 U63 ( .B1(n290), .B2(n454), .A(n451), .ZN(n350) );
  NAND2_X1 U64 ( .A1(\mem[3][2] ), .A2(n454), .ZN(n451) );
  OAI21_X1 U65 ( .B1(n289), .B2(n454), .A(n450), .ZN(n349) );
  NAND2_X1 U66 ( .A1(\mem[3][3] ), .A2(n454), .ZN(n450) );
  OAI21_X1 U67 ( .B1(n288), .B2(n454), .A(n449), .ZN(n348) );
  NAND2_X1 U68 ( .A1(\mem[3][4] ), .A2(n454), .ZN(n449) );
  OAI21_X1 U69 ( .B1(n287), .B2(n454), .A(n448), .ZN(n347) );
  NAND2_X1 U70 ( .A1(\mem[3][5] ), .A2(n454), .ZN(n448) );
  OAI21_X1 U71 ( .B1(n286), .B2(n454), .A(n447), .ZN(n346) );
  NAND2_X1 U72 ( .A1(\mem[3][6] ), .A2(n454), .ZN(n447) );
  OAI21_X1 U73 ( .B1(n285), .B2(n454), .A(n446), .ZN(n345) );
  NAND2_X1 U74 ( .A1(\mem[3][7] ), .A2(n454), .ZN(n446) );
  OAI21_X1 U75 ( .B1(n284), .B2(n454), .A(n445), .ZN(n344) );
  NAND2_X1 U76 ( .A1(\mem[3][8] ), .A2(n454), .ZN(n445) );
  OAI21_X1 U77 ( .B1(n283), .B2(n454), .A(n444), .ZN(n343) );
  NAND2_X1 U78 ( .A1(\mem[3][9] ), .A2(n454), .ZN(n444) );
  OAI21_X1 U79 ( .B1(n282), .B2(n454), .A(n443), .ZN(n342) );
  NAND2_X1 U80 ( .A1(\mem[3][10] ), .A2(n454), .ZN(n443) );
  OAI21_X1 U81 ( .B1(n281), .B2(n454), .A(n442), .ZN(n341) );
  NAND2_X1 U82 ( .A1(\mem[3][11] ), .A2(n454), .ZN(n442) );
  OAI21_X1 U83 ( .B1(n292), .B2(n441), .A(n440), .ZN(n340) );
  NAND2_X1 U84 ( .A1(\mem[4][0] ), .A2(n441), .ZN(n440) );
  OAI21_X1 U85 ( .B1(n291), .B2(n441), .A(n439), .ZN(n339) );
  NAND2_X1 U86 ( .A1(\mem[4][1] ), .A2(n441), .ZN(n439) );
  OAI21_X1 U87 ( .B1(n290), .B2(n441), .A(n438), .ZN(n338) );
  NAND2_X1 U88 ( .A1(\mem[4][2] ), .A2(n441), .ZN(n438) );
  OAI21_X1 U89 ( .B1(n289), .B2(n441), .A(n437), .ZN(n337) );
  NAND2_X1 U90 ( .A1(\mem[4][3] ), .A2(n441), .ZN(n437) );
  OAI21_X1 U91 ( .B1(n288), .B2(n441), .A(n436), .ZN(n336) );
  NAND2_X1 U92 ( .A1(\mem[4][4] ), .A2(n441), .ZN(n436) );
  OAI21_X1 U93 ( .B1(n287), .B2(n441), .A(n435), .ZN(n335) );
  NAND2_X1 U94 ( .A1(\mem[4][5] ), .A2(n441), .ZN(n435) );
  OAI21_X1 U95 ( .B1(n286), .B2(n441), .A(n434), .ZN(n334) );
  NAND2_X1 U96 ( .A1(\mem[4][6] ), .A2(n441), .ZN(n434) );
  OAI21_X1 U97 ( .B1(n285), .B2(n441), .A(n433), .ZN(n333) );
  NAND2_X1 U98 ( .A1(\mem[4][7] ), .A2(n441), .ZN(n433) );
  OAI21_X1 U99 ( .B1(n284), .B2(n441), .A(n432), .ZN(n332) );
  NAND2_X1 U100 ( .A1(\mem[4][8] ), .A2(n441), .ZN(n432) );
  OAI21_X1 U101 ( .B1(n283), .B2(n441), .A(n431), .ZN(n331) );
  NAND2_X1 U102 ( .A1(\mem[4][9] ), .A2(n441), .ZN(n431) );
  OAI21_X1 U103 ( .B1(n282), .B2(n441), .A(n430), .ZN(n330) );
  NAND2_X1 U104 ( .A1(\mem[4][10] ), .A2(n441), .ZN(n430) );
  OAI21_X1 U105 ( .B1(n281), .B2(n441), .A(n429), .ZN(n329) );
  NAND2_X1 U106 ( .A1(\mem[4][11] ), .A2(n441), .ZN(n429) );
  OAI21_X1 U107 ( .B1(n292), .B2(n427), .A(n426), .ZN(n328) );
  NAND2_X1 U108 ( .A1(\mem[5][0] ), .A2(n427), .ZN(n426) );
  OAI21_X1 U109 ( .B1(n291), .B2(n427), .A(n425), .ZN(n327) );
  NAND2_X1 U110 ( .A1(\mem[5][1] ), .A2(n427), .ZN(n425) );
  OAI21_X1 U111 ( .B1(n290), .B2(n427), .A(n424), .ZN(n326) );
  NAND2_X1 U112 ( .A1(\mem[5][2] ), .A2(n427), .ZN(n424) );
  OAI21_X1 U113 ( .B1(n289), .B2(n427), .A(n423), .ZN(n325) );
  NAND2_X1 U114 ( .A1(\mem[5][3] ), .A2(n427), .ZN(n423) );
  OAI21_X1 U115 ( .B1(n288), .B2(n427), .A(n422), .ZN(n324) );
  NAND2_X1 U116 ( .A1(\mem[5][4] ), .A2(n427), .ZN(n422) );
  OAI21_X1 U117 ( .B1(n287), .B2(n427), .A(n421), .ZN(n323) );
  NAND2_X1 U118 ( .A1(\mem[5][5] ), .A2(n427), .ZN(n421) );
  OAI21_X1 U119 ( .B1(n286), .B2(n427), .A(n420), .ZN(n322) );
  NAND2_X1 U120 ( .A1(\mem[5][6] ), .A2(n427), .ZN(n420) );
  OAI21_X1 U121 ( .B1(n285), .B2(n427), .A(n419), .ZN(n321) );
  NAND2_X1 U122 ( .A1(\mem[5][7] ), .A2(n427), .ZN(n419) );
  OAI21_X1 U123 ( .B1(n284), .B2(n427), .A(n418), .ZN(n320) );
  NAND2_X1 U124 ( .A1(\mem[5][8] ), .A2(n427), .ZN(n418) );
  OAI21_X1 U125 ( .B1(n283), .B2(n427), .A(n417), .ZN(n319) );
  NAND2_X1 U126 ( .A1(\mem[5][9] ), .A2(n427), .ZN(n417) );
  OAI21_X1 U127 ( .B1(n282), .B2(n427), .A(n416), .ZN(n318) );
  NAND2_X1 U128 ( .A1(\mem[5][10] ), .A2(n427), .ZN(n416) );
  OAI21_X1 U129 ( .B1(n281), .B2(n427), .A(n415), .ZN(n317) );
  NAND2_X1 U130 ( .A1(\mem[5][11] ), .A2(n427), .ZN(n415) );
  OAI21_X1 U131 ( .B1(n292), .B2(n414), .A(n413), .ZN(n316) );
  NAND2_X1 U132 ( .A1(\mem[6][0] ), .A2(n414), .ZN(n413) );
  OAI21_X1 U133 ( .B1(n291), .B2(n414), .A(n412), .ZN(n315) );
  NAND2_X1 U134 ( .A1(\mem[6][1] ), .A2(n414), .ZN(n412) );
  OAI21_X1 U135 ( .B1(n290), .B2(n414), .A(n411), .ZN(n314) );
  NAND2_X1 U136 ( .A1(\mem[6][2] ), .A2(n414), .ZN(n411) );
  OAI21_X1 U137 ( .B1(n289), .B2(n414), .A(n410), .ZN(n313) );
  NAND2_X1 U138 ( .A1(\mem[6][3] ), .A2(n414), .ZN(n410) );
  OAI21_X1 U139 ( .B1(n288), .B2(n414), .A(n409), .ZN(n312) );
  NAND2_X1 U140 ( .A1(\mem[6][4] ), .A2(n414), .ZN(n409) );
  OAI21_X1 U141 ( .B1(n287), .B2(n414), .A(n408), .ZN(n311) );
  NAND2_X1 U142 ( .A1(\mem[6][5] ), .A2(n414), .ZN(n408) );
  OAI21_X1 U143 ( .B1(n286), .B2(n414), .A(n407), .ZN(n310) );
  NAND2_X1 U144 ( .A1(\mem[6][6] ), .A2(n414), .ZN(n407) );
  OAI21_X1 U145 ( .B1(n285), .B2(n414), .A(n406), .ZN(n309) );
  NAND2_X1 U146 ( .A1(\mem[6][7] ), .A2(n414), .ZN(n406) );
  OAI21_X1 U147 ( .B1(n284), .B2(n414), .A(n405), .ZN(n308) );
  NAND2_X1 U148 ( .A1(\mem[6][8] ), .A2(n414), .ZN(n405) );
  OAI21_X1 U149 ( .B1(n283), .B2(n414), .A(n404), .ZN(n307) );
  NAND2_X1 U150 ( .A1(\mem[6][9] ), .A2(n414), .ZN(n404) );
  OAI21_X1 U151 ( .B1(n282), .B2(n414), .A(n403), .ZN(n306) );
  NAND2_X1 U152 ( .A1(\mem[6][10] ), .A2(n414), .ZN(n403) );
  OAI21_X1 U153 ( .B1(n281), .B2(n414), .A(n402), .ZN(n305) );
  NAND2_X1 U154 ( .A1(\mem[6][11] ), .A2(n414), .ZN(n402) );
  OAI21_X1 U155 ( .B1(n292), .B2(n401), .A(n400), .ZN(n304) );
  NAND2_X1 U156 ( .A1(\mem[7][0] ), .A2(n401), .ZN(n400) );
  OAI21_X1 U157 ( .B1(n291), .B2(n401), .A(n399), .ZN(n303) );
  NAND2_X1 U158 ( .A1(\mem[7][1] ), .A2(n401), .ZN(n399) );
  OAI21_X1 U159 ( .B1(n290), .B2(n401), .A(n398), .ZN(n302) );
  NAND2_X1 U160 ( .A1(\mem[7][2] ), .A2(n401), .ZN(n398) );
  OAI21_X1 U161 ( .B1(n289), .B2(n401), .A(n397), .ZN(n301) );
  NAND2_X1 U162 ( .A1(\mem[7][3] ), .A2(n401), .ZN(n397) );
  OAI21_X1 U163 ( .B1(n288), .B2(n401), .A(n396), .ZN(n300) );
  NAND2_X1 U164 ( .A1(\mem[7][4] ), .A2(n401), .ZN(n396) );
  OAI21_X1 U165 ( .B1(n287), .B2(n401), .A(n395), .ZN(n299) );
  NAND2_X1 U166 ( .A1(\mem[7][5] ), .A2(n401), .ZN(n395) );
  OAI21_X1 U167 ( .B1(n286), .B2(n401), .A(n394), .ZN(n298) );
  NAND2_X1 U168 ( .A1(\mem[7][6] ), .A2(n401), .ZN(n394) );
  OAI21_X1 U169 ( .B1(n285), .B2(n401), .A(n393), .ZN(n297) );
  NAND2_X1 U170 ( .A1(\mem[7][7] ), .A2(n401), .ZN(n393) );
  OAI21_X1 U171 ( .B1(n284), .B2(n401), .A(n392), .ZN(n296) );
  NAND2_X1 U172 ( .A1(\mem[7][8] ), .A2(n401), .ZN(n392) );
  OAI21_X1 U173 ( .B1(n283), .B2(n401), .A(n391), .ZN(n295) );
  NAND2_X1 U174 ( .A1(\mem[7][9] ), .A2(n401), .ZN(n391) );
  OAI21_X1 U175 ( .B1(n282), .B2(n401), .A(n390), .ZN(n294) );
  NAND2_X1 U176 ( .A1(\mem[7][10] ), .A2(n401), .ZN(n390) );
  OAI21_X1 U177 ( .B1(n281), .B2(n401), .A(n389), .ZN(n293) );
  NAND2_X1 U178 ( .A1(\mem[7][11] ), .A2(n401), .ZN(n389) );
  OAI21_X1 U179 ( .B1(n494), .B2(n292), .A(n493), .ZN(n388) );
  NAND2_X1 U180 ( .A1(\mem[0][0] ), .A2(n494), .ZN(n493) );
  OAI21_X1 U181 ( .B1(n494), .B2(n291), .A(n492), .ZN(n387) );
  NAND2_X1 U182 ( .A1(\mem[0][1] ), .A2(n494), .ZN(n492) );
  OAI21_X1 U183 ( .B1(n494), .B2(n290), .A(n491), .ZN(n386) );
  NAND2_X1 U184 ( .A1(\mem[0][2] ), .A2(n494), .ZN(n491) );
  OAI21_X1 U185 ( .B1(n494), .B2(n289), .A(n490), .ZN(n385) );
  NAND2_X1 U186 ( .A1(\mem[0][3] ), .A2(n494), .ZN(n490) );
  OAI21_X1 U187 ( .B1(n494), .B2(n288), .A(n489), .ZN(n384) );
  NAND2_X1 U188 ( .A1(\mem[0][4] ), .A2(n494), .ZN(n489) );
  OAI21_X1 U189 ( .B1(n494), .B2(n287), .A(n488), .ZN(n383) );
  NAND2_X1 U190 ( .A1(\mem[0][5] ), .A2(n494), .ZN(n488) );
  OAI21_X1 U191 ( .B1(n494), .B2(n286), .A(n487), .ZN(n382) );
  NAND2_X1 U192 ( .A1(\mem[0][6] ), .A2(n494), .ZN(n487) );
  OAI21_X1 U193 ( .B1(n494), .B2(n285), .A(n486), .ZN(n381) );
  NAND2_X1 U194 ( .A1(\mem[0][7] ), .A2(n494), .ZN(n486) );
  OAI21_X1 U195 ( .B1(n494), .B2(n284), .A(n485), .ZN(n380) );
  NAND2_X1 U196 ( .A1(\mem[0][8] ), .A2(n494), .ZN(n485) );
  OAI21_X1 U197 ( .B1(n494), .B2(n283), .A(n484), .ZN(n379) );
  NAND2_X1 U198 ( .A1(\mem[0][9] ), .A2(n494), .ZN(n484) );
  OAI21_X1 U199 ( .B1(n494), .B2(n282), .A(n483), .ZN(n378) );
  NAND2_X1 U200 ( .A1(\mem[0][10] ), .A2(n494), .ZN(n483) );
  OAI21_X1 U201 ( .B1(n494), .B2(n281), .A(n482), .ZN(n377) );
  NAND2_X1 U202 ( .A1(\mem[0][11] ), .A2(n494), .ZN(n482) );
  INV_X1 U203 ( .A(data_in[0]), .ZN(n292) );
  INV_X1 U204 ( .A(data_in[1]), .ZN(n291) );
  INV_X1 U205 ( .A(data_in[2]), .ZN(n290) );
  INV_X1 U206 ( .A(data_in[3]), .ZN(n289) );
  INV_X1 U207 ( .A(data_in[4]), .ZN(n288) );
  INV_X1 U208 ( .A(data_in[5]), .ZN(n287) );
  INV_X1 U209 ( .A(data_in[6]), .ZN(n286) );
  INV_X1 U210 ( .A(data_in[7]), .ZN(n285) );
  INV_X1 U211 ( .A(data_in[8]), .ZN(n284) );
  INV_X1 U220 ( .A(data_in[9]), .ZN(n283) );
  INV_X1 U221 ( .A(data_in[10]), .ZN(n282) );
  INV_X1 U222 ( .A(data_in[11]), .ZN(n281) );
  MUX2_X1 U223 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n276), .Z(n1) );
  MUX2_X1 U224 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n276), .Z(n2) );
  MUX2_X1 U225 ( .A(n2), .B(n1), .S(n275), .Z(n3) );
  MUX2_X1 U226 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n276), .Z(n4) );
  MUX2_X1 U227 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n276), .Z(n5) );
  MUX2_X1 U228 ( .A(n5), .B(n4), .S(n275), .Z(n6) );
  MUX2_X1 U229 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n276), .Z(n7) );
  MUX2_X1 U230 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n276), .Z(n8) );
  MUX2_X1 U231 ( .A(n8), .B(n7), .S(n275), .Z(n9) );
  MUX2_X1 U232 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n276), .Z(n10) );
  MUX2_X1 U233 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n276), .Z(n11) );
  MUX2_X1 U234 ( .A(n11), .B(n10), .S(n275), .Z(n12) );
  MUX2_X1 U235 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n276), .Z(n13) );
  MUX2_X1 U236 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n276), .Z(n14) );
  MUX2_X1 U237 ( .A(n14), .B(n13), .S(n275), .Z(n15) );
  MUX2_X1 U238 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n276), .Z(n218) );
  MUX2_X1 U239 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n276), .Z(n219) );
  MUX2_X1 U240 ( .A(n219), .B(n218), .S(n275), .Z(n220) );
  MUX2_X1 U241 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n277), .Z(n221) );
  MUX2_X1 U242 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n277), .Z(n222) );
  MUX2_X1 U243 ( .A(n222), .B(n221), .S(n275), .Z(n223) );
  MUX2_X1 U244 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n277), .Z(n224) );
  MUX2_X1 U245 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n277), .Z(n225) );
  MUX2_X1 U246 ( .A(n225), .B(n224), .S(n275), .Z(n226) );
  MUX2_X1 U247 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n277), .Z(n227) );
  MUX2_X1 U248 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n277), .Z(n228) );
  MUX2_X1 U249 ( .A(n228), .B(n227), .S(n275), .Z(n229) );
  MUX2_X1 U250 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n277), .Z(n230) );
  MUX2_X1 U251 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n277), .Z(n231) );
  MUX2_X1 U252 ( .A(n231), .B(n230), .S(n275), .Z(n232) );
  MUX2_X1 U253 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n277), .Z(n233) );
  MUX2_X1 U254 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n277), .Z(n234) );
  MUX2_X1 U255 ( .A(n234), .B(n233), .S(n275), .Z(n235) );
  MUX2_X1 U256 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n277), .Z(n236) );
  MUX2_X1 U257 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n277), .Z(n237) );
  MUX2_X1 U258 ( .A(n237), .B(n236), .S(n275), .Z(n238) );
  MUX2_X1 U259 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n277), .Z(n239) );
  MUX2_X1 U260 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n240) );
  MUX2_X1 U261 ( .A(n240), .B(n239), .S(n275), .Z(n241) );
  MUX2_X1 U262 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n242) );
  MUX2_X1 U263 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n243) );
  MUX2_X1 U264 ( .A(n243), .B(n242), .S(n275), .Z(n244) );
  MUX2_X1 U265 ( .A(n244), .B(n241), .S(N12), .Z(N18) );
  MUX2_X1 U266 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n245) );
  MUX2_X1 U267 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n246) );
  MUX2_X1 U268 ( .A(n246), .B(n245), .S(n275), .Z(n247) );
  MUX2_X1 U269 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n277), .Z(n248) );
  MUX2_X1 U270 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n277), .Z(n249) );
  MUX2_X1 U271 ( .A(n249), .B(n248), .S(n275), .Z(n250) );
  MUX2_X1 U272 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(N10), .Z(n251) );
  MUX2_X1 U273 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n277), .Z(n252) );
  MUX2_X1 U274 ( .A(n252), .B(n251), .S(n275), .Z(n253) );
  MUX2_X1 U275 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n277), .Z(n254) );
  MUX2_X1 U276 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n277), .Z(n255) );
  MUX2_X1 U277 ( .A(n255), .B(n254), .S(n275), .Z(n256) );
  MUX2_X1 U278 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(N10), .Z(n257) );
  MUX2_X1 U279 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(N10), .Z(n258) );
  MUX2_X1 U280 ( .A(n258), .B(n257), .S(n275), .Z(n259) );
  MUX2_X1 U281 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(N10), .Z(n260) );
  MUX2_X1 U282 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(N10), .Z(n261) );
  MUX2_X1 U283 ( .A(n261), .B(n260), .S(N11), .Z(n262) );
  MUX2_X1 U284 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n277), .Z(n263) );
  MUX2_X1 U285 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(N10), .Z(n264) );
  MUX2_X1 U286 ( .A(n264), .B(n263), .S(n275), .Z(n265) );
  MUX2_X1 U287 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n277), .Z(n266) );
  MUX2_X1 U288 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n277), .Z(n267) );
  MUX2_X1 U289 ( .A(n267), .B(n266), .S(n275), .Z(n268) );
  MUX2_X1 U290 ( .A(n268), .B(n265), .S(N12), .Z(N14) );
  MUX2_X1 U291 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(N10), .Z(n269) );
  MUX2_X1 U292 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(N10), .Z(n270) );
  MUX2_X1 U293 ( .A(n270), .B(n269), .S(n275), .Z(n271) );
  MUX2_X1 U294 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(N10), .Z(n272) );
  MUX2_X1 U295 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(N10), .Z(n273) );
  MUX2_X1 U296 ( .A(n273), .B(n272), .S(N11), .Z(n274) );
endmodule


module memory_WIDTH12_SIZE8_LOGSIZE3_5 ( clk, data_in, data_out, addr, wr_en
 );
  input [11:0] data_in;
  output [11:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] ,
         \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] ,
         \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][11] , \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] ,
         \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] ,
         \mem[5][1] , \mem[5][0] , \mem[4][11] , \mem[4][10] , \mem[4][9] ,
         \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] ,
         \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] ,
         \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] ,
         \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][11] , \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] ,
         \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] ,
         \mem[0][1] , \mem[0][0] , N17, N21, N23, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[7]  ( .D(N17), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[3]  ( .D(N21), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[1]  ( .D(N23), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[7][11]  ( .D(n293), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n294), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n295), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n296), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n297), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n298), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n299), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n300), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n301), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n302), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n303), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n304), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n305), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n306), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n307), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n308), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n309), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n310), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n311), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n312), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n313), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n314), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n315), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n316), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n317), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n318), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n319), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n320), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n321), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n322), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n323), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n324), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n325), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n326), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n327), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n328), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n329), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n330), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n331), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n332), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n333), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n334), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n335), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n336), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n337), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n338), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n339), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n340), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n341), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n342), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n343), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n344), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n345), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n346), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n347), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n348), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n349), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n350), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n351), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n352), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n353), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n354), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n355), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n356), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n357), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n358), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n359), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n360), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n361), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n362), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n363), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n364), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n365), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n366), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n367), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n368), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n369), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n370), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n371), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n372), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n373), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n374), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n375), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n376), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n377), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n378), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n379), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n380), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n381), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n382), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n383), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n384), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n385), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n386), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n387), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n388), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U212 ( .A1(n278), .A2(n279), .A3(n481), .ZN(n494) );
  NAND3_X1 U213 ( .A1(n481), .A2(n279), .A3(N10), .ZN(n480) );
  NAND3_X1 U214 ( .A1(n481), .A2(n278), .A3(N11), .ZN(n467) );
  NAND3_X1 U215 ( .A1(N10), .A2(n481), .A3(N11), .ZN(n454) );
  NAND3_X1 U216 ( .A1(n278), .A2(n279), .A3(n428), .ZN(n441) );
  NAND3_X1 U217 ( .A1(N10), .A2(n279), .A3(n428), .ZN(n427) );
  NAND3_X1 U218 ( .A1(N11), .A2(n278), .A3(n428), .ZN(n414) );
  NAND3_X1 U219 ( .A1(N11), .A2(N10), .A3(n428), .ZN(n401) );
  SDFF_X1 \data_out_reg[5]  ( .D(n238), .SI(n235), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n262), .SI(n259), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n274), .SI(n271), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[8]  ( .D(n256), .SI(n253), .SE(N12), .CK(clk), .Q(
        data_out[8]) );
  SDFF_X1 \data_out_reg[6]  ( .D(n244), .SI(n241), .SE(N12), .CK(clk), .Q(
        data_out[6]) );
  SDFF_X1 \data_out_reg[4]  ( .D(n232), .SI(n229), .SE(N12), .CK(clk), .Q(
        data_out[4]) );
  SDFF_X1 \data_out_reg[2]  ( .D(n220), .SI(n15), .SE(N12), .CK(clk), .Q(
        data_out[2]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n6), .SI(n3), .SE(N12), .CK(clk), .Q(
        data_out[0]) );
  SDFF_X1 \data_out_reg[10]  ( .D(n268), .SI(n265), .SE(N12), .CK(clk), .Q(
        data_out[10]) );
  BUF_X1 U3 ( .A(n277), .Z(n276) );
  BUF_X1 U4 ( .A(N11), .Z(n275) );
  BUF_X1 U5 ( .A(N10), .Z(n277) );
  NOR2_X1 U6 ( .A1(n280), .A2(N12), .ZN(n481) );
  INV_X1 U7 ( .A(wr_en), .ZN(n280) );
  AND2_X1 U8 ( .A1(N12), .A2(wr_en), .ZN(n428) );
  INV_X1 U9 ( .A(N10), .ZN(n278) );
  INV_X1 U10 ( .A(N11), .ZN(n279) );
  OAI21_X1 U11 ( .B1(n292), .B2(n480), .A(n479), .ZN(n376) );
  NAND2_X1 U12 ( .A1(\mem[1][0] ), .A2(n480), .ZN(n479) );
  OAI21_X1 U13 ( .B1(n291), .B2(n480), .A(n478), .ZN(n375) );
  NAND2_X1 U14 ( .A1(\mem[1][1] ), .A2(n480), .ZN(n478) );
  OAI21_X1 U15 ( .B1(n290), .B2(n480), .A(n477), .ZN(n374) );
  NAND2_X1 U16 ( .A1(\mem[1][2] ), .A2(n480), .ZN(n477) );
  OAI21_X1 U17 ( .B1(n289), .B2(n480), .A(n476), .ZN(n373) );
  NAND2_X1 U18 ( .A1(\mem[1][3] ), .A2(n480), .ZN(n476) );
  OAI21_X1 U19 ( .B1(n288), .B2(n480), .A(n475), .ZN(n372) );
  NAND2_X1 U20 ( .A1(\mem[1][4] ), .A2(n480), .ZN(n475) );
  OAI21_X1 U21 ( .B1(n287), .B2(n480), .A(n474), .ZN(n371) );
  NAND2_X1 U22 ( .A1(\mem[1][5] ), .A2(n480), .ZN(n474) );
  OAI21_X1 U23 ( .B1(n286), .B2(n480), .A(n473), .ZN(n370) );
  NAND2_X1 U24 ( .A1(\mem[1][6] ), .A2(n480), .ZN(n473) );
  OAI21_X1 U25 ( .B1(n285), .B2(n480), .A(n472), .ZN(n369) );
  NAND2_X1 U26 ( .A1(\mem[1][7] ), .A2(n480), .ZN(n472) );
  OAI21_X1 U27 ( .B1(n284), .B2(n480), .A(n471), .ZN(n368) );
  NAND2_X1 U28 ( .A1(\mem[1][8] ), .A2(n480), .ZN(n471) );
  OAI21_X1 U29 ( .B1(n283), .B2(n480), .A(n470), .ZN(n367) );
  NAND2_X1 U30 ( .A1(\mem[1][9] ), .A2(n480), .ZN(n470) );
  OAI21_X1 U31 ( .B1(n282), .B2(n480), .A(n469), .ZN(n366) );
  NAND2_X1 U32 ( .A1(\mem[1][10] ), .A2(n480), .ZN(n469) );
  OAI21_X1 U33 ( .B1(n281), .B2(n480), .A(n468), .ZN(n365) );
  NAND2_X1 U34 ( .A1(\mem[1][11] ), .A2(n480), .ZN(n468) );
  OAI21_X1 U35 ( .B1(n292), .B2(n467), .A(n466), .ZN(n364) );
  NAND2_X1 U36 ( .A1(\mem[2][0] ), .A2(n467), .ZN(n466) );
  OAI21_X1 U37 ( .B1(n291), .B2(n467), .A(n465), .ZN(n363) );
  NAND2_X1 U38 ( .A1(\mem[2][1] ), .A2(n467), .ZN(n465) );
  OAI21_X1 U39 ( .B1(n290), .B2(n467), .A(n464), .ZN(n362) );
  NAND2_X1 U40 ( .A1(\mem[2][2] ), .A2(n467), .ZN(n464) );
  OAI21_X1 U41 ( .B1(n289), .B2(n467), .A(n463), .ZN(n361) );
  NAND2_X1 U42 ( .A1(\mem[2][3] ), .A2(n467), .ZN(n463) );
  OAI21_X1 U43 ( .B1(n288), .B2(n467), .A(n462), .ZN(n360) );
  NAND2_X1 U44 ( .A1(\mem[2][4] ), .A2(n467), .ZN(n462) );
  OAI21_X1 U45 ( .B1(n287), .B2(n467), .A(n461), .ZN(n359) );
  NAND2_X1 U46 ( .A1(\mem[2][5] ), .A2(n467), .ZN(n461) );
  OAI21_X1 U47 ( .B1(n286), .B2(n467), .A(n460), .ZN(n358) );
  NAND2_X1 U48 ( .A1(\mem[2][6] ), .A2(n467), .ZN(n460) );
  OAI21_X1 U49 ( .B1(n285), .B2(n467), .A(n459), .ZN(n357) );
  NAND2_X1 U50 ( .A1(\mem[2][7] ), .A2(n467), .ZN(n459) );
  OAI21_X1 U51 ( .B1(n284), .B2(n467), .A(n458), .ZN(n356) );
  NAND2_X1 U52 ( .A1(\mem[2][8] ), .A2(n467), .ZN(n458) );
  OAI21_X1 U53 ( .B1(n283), .B2(n467), .A(n457), .ZN(n355) );
  NAND2_X1 U54 ( .A1(\mem[2][9] ), .A2(n467), .ZN(n457) );
  OAI21_X1 U55 ( .B1(n282), .B2(n467), .A(n456), .ZN(n354) );
  NAND2_X1 U56 ( .A1(\mem[2][10] ), .A2(n467), .ZN(n456) );
  OAI21_X1 U57 ( .B1(n281), .B2(n467), .A(n455), .ZN(n353) );
  NAND2_X1 U58 ( .A1(\mem[2][11] ), .A2(n467), .ZN(n455) );
  OAI21_X1 U59 ( .B1(n292), .B2(n454), .A(n453), .ZN(n352) );
  NAND2_X1 U60 ( .A1(\mem[3][0] ), .A2(n454), .ZN(n453) );
  OAI21_X1 U61 ( .B1(n291), .B2(n454), .A(n452), .ZN(n351) );
  NAND2_X1 U62 ( .A1(\mem[3][1] ), .A2(n454), .ZN(n452) );
  OAI21_X1 U63 ( .B1(n290), .B2(n454), .A(n451), .ZN(n350) );
  NAND2_X1 U64 ( .A1(\mem[3][2] ), .A2(n454), .ZN(n451) );
  OAI21_X1 U65 ( .B1(n289), .B2(n454), .A(n450), .ZN(n349) );
  NAND2_X1 U66 ( .A1(\mem[3][3] ), .A2(n454), .ZN(n450) );
  OAI21_X1 U67 ( .B1(n288), .B2(n454), .A(n449), .ZN(n348) );
  NAND2_X1 U68 ( .A1(\mem[3][4] ), .A2(n454), .ZN(n449) );
  OAI21_X1 U69 ( .B1(n287), .B2(n454), .A(n448), .ZN(n347) );
  NAND2_X1 U70 ( .A1(\mem[3][5] ), .A2(n454), .ZN(n448) );
  OAI21_X1 U71 ( .B1(n286), .B2(n454), .A(n447), .ZN(n346) );
  NAND2_X1 U72 ( .A1(\mem[3][6] ), .A2(n454), .ZN(n447) );
  OAI21_X1 U73 ( .B1(n285), .B2(n454), .A(n446), .ZN(n345) );
  NAND2_X1 U74 ( .A1(\mem[3][7] ), .A2(n454), .ZN(n446) );
  OAI21_X1 U75 ( .B1(n284), .B2(n454), .A(n445), .ZN(n344) );
  NAND2_X1 U76 ( .A1(\mem[3][8] ), .A2(n454), .ZN(n445) );
  OAI21_X1 U77 ( .B1(n283), .B2(n454), .A(n444), .ZN(n343) );
  NAND2_X1 U78 ( .A1(\mem[3][9] ), .A2(n454), .ZN(n444) );
  OAI21_X1 U79 ( .B1(n282), .B2(n454), .A(n443), .ZN(n342) );
  NAND2_X1 U80 ( .A1(\mem[3][10] ), .A2(n454), .ZN(n443) );
  OAI21_X1 U81 ( .B1(n281), .B2(n454), .A(n442), .ZN(n341) );
  NAND2_X1 U82 ( .A1(\mem[3][11] ), .A2(n454), .ZN(n442) );
  OAI21_X1 U83 ( .B1(n292), .B2(n441), .A(n440), .ZN(n340) );
  NAND2_X1 U84 ( .A1(\mem[4][0] ), .A2(n441), .ZN(n440) );
  OAI21_X1 U85 ( .B1(n291), .B2(n441), .A(n439), .ZN(n339) );
  NAND2_X1 U86 ( .A1(\mem[4][1] ), .A2(n441), .ZN(n439) );
  OAI21_X1 U87 ( .B1(n290), .B2(n441), .A(n438), .ZN(n338) );
  NAND2_X1 U88 ( .A1(\mem[4][2] ), .A2(n441), .ZN(n438) );
  OAI21_X1 U89 ( .B1(n289), .B2(n441), .A(n437), .ZN(n337) );
  NAND2_X1 U90 ( .A1(\mem[4][3] ), .A2(n441), .ZN(n437) );
  OAI21_X1 U91 ( .B1(n288), .B2(n441), .A(n436), .ZN(n336) );
  NAND2_X1 U92 ( .A1(\mem[4][4] ), .A2(n441), .ZN(n436) );
  OAI21_X1 U93 ( .B1(n287), .B2(n441), .A(n435), .ZN(n335) );
  NAND2_X1 U94 ( .A1(\mem[4][5] ), .A2(n441), .ZN(n435) );
  OAI21_X1 U95 ( .B1(n286), .B2(n441), .A(n434), .ZN(n334) );
  NAND2_X1 U96 ( .A1(\mem[4][6] ), .A2(n441), .ZN(n434) );
  OAI21_X1 U97 ( .B1(n285), .B2(n441), .A(n433), .ZN(n333) );
  NAND2_X1 U98 ( .A1(\mem[4][7] ), .A2(n441), .ZN(n433) );
  OAI21_X1 U99 ( .B1(n284), .B2(n441), .A(n432), .ZN(n332) );
  NAND2_X1 U100 ( .A1(\mem[4][8] ), .A2(n441), .ZN(n432) );
  OAI21_X1 U101 ( .B1(n283), .B2(n441), .A(n431), .ZN(n331) );
  NAND2_X1 U102 ( .A1(\mem[4][9] ), .A2(n441), .ZN(n431) );
  OAI21_X1 U103 ( .B1(n282), .B2(n441), .A(n430), .ZN(n330) );
  NAND2_X1 U104 ( .A1(\mem[4][10] ), .A2(n441), .ZN(n430) );
  OAI21_X1 U105 ( .B1(n281), .B2(n441), .A(n429), .ZN(n329) );
  NAND2_X1 U106 ( .A1(\mem[4][11] ), .A2(n441), .ZN(n429) );
  OAI21_X1 U107 ( .B1(n292), .B2(n427), .A(n426), .ZN(n328) );
  NAND2_X1 U108 ( .A1(\mem[5][0] ), .A2(n427), .ZN(n426) );
  OAI21_X1 U109 ( .B1(n291), .B2(n427), .A(n425), .ZN(n327) );
  NAND2_X1 U110 ( .A1(\mem[5][1] ), .A2(n427), .ZN(n425) );
  OAI21_X1 U111 ( .B1(n290), .B2(n427), .A(n424), .ZN(n326) );
  NAND2_X1 U112 ( .A1(\mem[5][2] ), .A2(n427), .ZN(n424) );
  OAI21_X1 U113 ( .B1(n289), .B2(n427), .A(n423), .ZN(n325) );
  NAND2_X1 U114 ( .A1(\mem[5][3] ), .A2(n427), .ZN(n423) );
  OAI21_X1 U115 ( .B1(n288), .B2(n427), .A(n422), .ZN(n324) );
  NAND2_X1 U116 ( .A1(\mem[5][4] ), .A2(n427), .ZN(n422) );
  OAI21_X1 U117 ( .B1(n287), .B2(n427), .A(n421), .ZN(n323) );
  NAND2_X1 U118 ( .A1(\mem[5][5] ), .A2(n427), .ZN(n421) );
  OAI21_X1 U119 ( .B1(n286), .B2(n427), .A(n420), .ZN(n322) );
  NAND2_X1 U120 ( .A1(\mem[5][6] ), .A2(n427), .ZN(n420) );
  OAI21_X1 U121 ( .B1(n285), .B2(n427), .A(n419), .ZN(n321) );
  NAND2_X1 U122 ( .A1(\mem[5][7] ), .A2(n427), .ZN(n419) );
  OAI21_X1 U123 ( .B1(n284), .B2(n427), .A(n418), .ZN(n320) );
  NAND2_X1 U124 ( .A1(\mem[5][8] ), .A2(n427), .ZN(n418) );
  OAI21_X1 U125 ( .B1(n283), .B2(n427), .A(n417), .ZN(n319) );
  NAND2_X1 U126 ( .A1(\mem[5][9] ), .A2(n427), .ZN(n417) );
  OAI21_X1 U127 ( .B1(n282), .B2(n427), .A(n416), .ZN(n318) );
  NAND2_X1 U128 ( .A1(\mem[5][10] ), .A2(n427), .ZN(n416) );
  OAI21_X1 U129 ( .B1(n281), .B2(n427), .A(n415), .ZN(n317) );
  NAND2_X1 U130 ( .A1(\mem[5][11] ), .A2(n427), .ZN(n415) );
  OAI21_X1 U131 ( .B1(n292), .B2(n414), .A(n413), .ZN(n316) );
  NAND2_X1 U132 ( .A1(\mem[6][0] ), .A2(n414), .ZN(n413) );
  OAI21_X1 U133 ( .B1(n291), .B2(n414), .A(n412), .ZN(n315) );
  NAND2_X1 U134 ( .A1(\mem[6][1] ), .A2(n414), .ZN(n412) );
  OAI21_X1 U135 ( .B1(n290), .B2(n414), .A(n411), .ZN(n314) );
  NAND2_X1 U136 ( .A1(\mem[6][2] ), .A2(n414), .ZN(n411) );
  OAI21_X1 U137 ( .B1(n289), .B2(n414), .A(n410), .ZN(n313) );
  NAND2_X1 U138 ( .A1(\mem[6][3] ), .A2(n414), .ZN(n410) );
  OAI21_X1 U139 ( .B1(n288), .B2(n414), .A(n409), .ZN(n312) );
  NAND2_X1 U140 ( .A1(\mem[6][4] ), .A2(n414), .ZN(n409) );
  OAI21_X1 U141 ( .B1(n287), .B2(n414), .A(n408), .ZN(n311) );
  NAND2_X1 U142 ( .A1(\mem[6][5] ), .A2(n414), .ZN(n408) );
  OAI21_X1 U143 ( .B1(n286), .B2(n414), .A(n407), .ZN(n310) );
  NAND2_X1 U144 ( .A1(\mem[6][6] ), .A2(n414), .ZN(n407) );
  OAI21_X1 U145 ( .B1(n285), .B2(n414), .A(n406), .ZN(n309) );
  NAND2_X1 U146 ( .A1(\mem[6][7] ), .A2(n414), .ZN(n406) );
  OAI21_X1 U147 ( .B1(n284), .B2(n414), .A(n405), .ZN(n308) );
  NAND2_X1 U148 ( .A1(\mem[6][8] ), .A2(n414), .ZN(n405) );
  OAI21_X1 U149 ( .B1(n283), .B2(n414), .A(n404), .ZN(n307) );
  NAND2_X1 U150 ( .A1(\mem[6][9] ), .A2(n414), .ZN(n404) );
  OAI21_X1 U151 ( .B1(n282), .B2(n414), .A(n403), .ZN(n306) );
  NAND2_X1 U152 ( .A1(\mem[6][10] ), .A2(n414), .ZN(n403) );
  OAI21_X1 U153 ( .B1(n281), .B2(n414), .A(n402), .ZN(n305) );
  NAND2_X1 U154 ( .A1(\mem[6][11] ), .A2(n414), .ZN(n402) );
  OAI21_X1 U155 ( .B1(n292), .B2(n401), .A(n400), .ZN(n304) );
  NAND2_X1 U156 ( .A1(\mem[7][0] ), .A2(n401), .ZN(n400) );
  OAI21_X1 U157 ( .B1(n291), .B2(n401), .A(n399), .ZN(n303) );
  NAND2_X1 U158 ( .A1(\mem[7][1] ), .A2(n401), .ZN(n399) );
  OAI21_X1 U159 ( .B1(n290), .B2(n401), .A(n398), .ZN(n302) );
  NAND2_X1 U160 ( .A1(\mem[7][2] ), .A2(n401), .ZN(n398) );
  OAI21_X1 U161 ( .B1(n289), .B2(n401), .A(n397), .ZN(n301) );
  NAND2_X1 U162 ( .A1(\mem[7][3] ), .A2(n401), .ZN(n397) );
  OAI21_X1 U163 ( .B1(n288), .B2(n401), .A(n396), .ZN(n300) );
  NAND2_X1 U164 ( .A1(\mem[7][4] ), .A2(n401), .ZN(n396) );
  OAI21_X1 U165 ( .B1(n287), .B2(n401), .A(n395), .ZN(n299) );
  NAND2_X1 U166 ( .A1(\mem[7][5] ), .A2(n401), .ZN(n395) );
  OAI21_X1 U167 ( .B1(n286), .B2(n401), .A(n394), .ZN(n298) );
  NAND2_X1 U168 ( .A1(\mem[7][6] ), .A2(n401), .ZN(n394) );
  OAI21_X1 U169 ( .B1(n285), .B2(n401), .A(n393), .ZN(n297) );
  NAND2_X1 U170 ( .A1(\mem[7][7] ), .A2(n401), .ZN(n393) );
  OAI21_X1 U171 ( .B1(n284), .B2(n401), .A(n392), .ZN(n296) );
  NAND2_X1 U172 ( .A1(\mem[7][8] ), .A2(n401), .ZN(n392) );
  OAI21_X1 U173 ( .B1(n283), .B2(n401), .A(n391), .ZN(n295) );
  NAND2_X1 U174 ( .A1(\mem[7][9] ), .A2(n401), .ZN(n391) );
  OAI21_X1 U175 ( .B1(n282), .B2(n401), .A(n390), .ZN(n294) );
  NAND2_X1 U176 ( .A1(\mem[7][10] ), .A2(n401), .ZN(n390) );
  OAI21_X1 U177 ( .B1(n281), .B2(n401), .A(n389), .ZN(n293) );
  NAND2_X1 U178 ( .A1(\mem[7][11] ), .A2(n401), .ZN(n389) );
  OAI21_X1 U179 ( .B1(n494), .B2(n292), .A(n493), .ZN(n388) );
  NAND2_X1 U180 ( .A1(\mem[0][0] ), .A2(n494), .ZN(n493) );
  OAI21_X1 U181 ( .B1(n494), .B2(n291), .A(n492), .ZN(n387) );
  NAND2_X1 U182 ( .A1(\mem[0][1] ), .A2(n494), .ZN(n492) );
  OAI21_X1 U183 ( .B1(n494), .B2(n290), .A(n491), .ZN(n386) );
  NAND2_X1 U184 ( .A1(\mem[0][2] ), .A2(n494), .ZN(n491) );
  OAI21_X1 U185 ( .B1(n494), .B2(n289), .A(n490), .ZN(n385) );
  NAND2_X1 U186 ( .A1(\mem[0][3] ), .A2(n494), .ZN(n490) );
  OAI21_X1 U187 ( .B1(n494), .B2(n288), .A(n489), .ZN(n384) );
  NAND2_X1 U188 ( .A1(\mem[0][4] ), .A2(n494), .ZN(n489) );
  OAI21_X1 U189 ( .B1(n494), .B2(n287), .A(n488), .ZN(n383) );
  NAND2_X1 U190 ( .A1(\mem[0][5] ), .A2(n494), .ZN(n488) );
  OAI21_X1 U191 ( .B1(n494), .B2(n286), .A(n487), .ZN(n382) );
  NAND2_X1 U192 ( .A1(\mem[0][6] ), .A2(n494), .ZN(n487) );
  OAI21_X1 U193 ( .B1(n494), .B2(n285), .A(n486), .ZN(n381) );
  NAND2_X1 U194 ( .A1(\mem[0][7] ), .A2(n494), .ZN(n486) );
  OAI21_X1 U195 ( .B1(n494), .B2(n284), .A(n485), .ZN(n380) );
  NAND2_X1 U196 ( .A1(\mem[0][8] ), .A2(n494), .ZN(n485) );
  OAI21_X1 U197 ( .B1(n494), .B2(n283), .A(n484), .ZN(n379) );
  NAND2_X1 U198 ( .A1(\mem[0][9] ), .A2(n494), .ZN(n484) );
  OAI21_X1 U199 ( .B1(n494), .B2(n282), .A(n483), .ZN(n378) );
  NAND2_X1 U200 ( .A1(\mem[0][10] ), .A2(n494), .ZN(n483) );
  OAI21_X1 U201 ( .B1(n494), .B2(n281), .A(n482), .ZN(n377) );
  NAND2_X1 U202 ( .A1(\mem[0][11] ), .A2(n494), .ZN(n482) );
  INV_X1 U203 ( .A(data_in[0]), .ZN(n292) );
  INV_X1 U204 ( .A(data_in[1]), .ZN(n291) );
  INV_X1 U205 ( .A(data_in[2]), .ZN(n290) );
  INV_X1 U206 ( .A(data_in[3]), .ZN(n289) );
  INV_X1 U207 ( .A(data_in[4]), .ZN(n288) );
  INV_X1 U208 ( .A(data_in[5]), .ZN(n287) );
  INV_X1 U209 ( .A(data_in[6]), .ZN(n286) );
  INV_X1 U210 ( .A(data_in[7]), .ZN(n285) );
  INV_X1 U211 ( .A(data_in[8]), .ZN(n284) );
  INV_X1 U220 ( .A(data_in[9]), .ZN(n283) );
  INV_X1 U221 ( .A(data_in[10]), .ZN(n282) );
  INV_X1 U222 ( .A(data_in[11]), .ZN(n281) );
  MUX2_X1 U223 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n276), .Z(n1) );
  MUX2_X1 U224 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n276), .Z(n2) );
  MUX2_X1 U225 ( .A(n2), .B(n1), .S(n275), .Z(n3) );
  MUX2_X1 U226 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n276), .Z(n4) );
  MUX2_X1 U227 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n276), .Z(n5) );
  MUX2_X1 U228 ( .A(n5), .B(n4), .S(n275), .Z(n6) );
  MUX2_X1 U229 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n276), .Z(n7) );
  MUX2_X1 U230 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n276), .Z(n8) );
  MUX2_X1 U231 ( .A(n8), .B(n7), .S(n275), .Z(n9) );
  MUX2_X1 U232 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n276), .Z(n10) );
  MUX2_X1 U233 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n276), .Z(n11) );
  MUX2_X1 U234 ( .A(n11), .B(n10), .S(n275), .Z(n12) );
  MUX2_X1 U235 ( .A(n12), .B(n9), .S(N12), .Z(N23) );
  MUX2_X1 U236 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n276), .Z(n13) );
  MUX2_X1 U237 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n276), .Z(n14) );
  MUX2_X1 U238 ( .A(n14), .B(n13), .S(n275), .Z(n15) );
  MUX2_X1 U239 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n276), .Z(n218) );
  MUX2_X1 U240 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n276), .Z(n219) );
  MUX2_X1 U241 ( .A(n219), .B(n218), .S(n275), .Z(n220) );
  MUX2_X1 U242 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n277), .Z(n221) );
  MUX2_X1 U243 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n277), .Z(n222) );
  MUX2_X1 U244 ( .A(n222), .B(n221), .S(n275), .Z(n223) );
  MUX2_X1 U245 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n277), .Z(n224) );
  MUX2_X1 U246 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n277), .Z(n225) );
  MUX2_X1 U247 ( .A(n225), .B(n224), .S(n275), .Z(n226) );
  MUX2_X1 U248 ( .A(n226), .B(n223), .S(N12), .Z(N21) );
  MUX2_X1 U249 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n277), .Z(n227) );
  MUX2_X1 U250 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n277), .Z(n228) );
  MUX2_X1 U251 ( .A(n228), .B(n227), .S(n275), .Z(n229) );
  MUX2_X1 U252 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n277), .Z(n230) );
  MUX2_X1 U253 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n277), .Z(n231) );
  MUX2_X1 U254 ( .A(n231), .B(n230), .S(n275), .Z(n232) );
  MUX2_X1 U255 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n277), .Z(n233) );
  MUX2_X1 U256 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n277), .Z(n234) );
  MUX2_X1 U257 ( .A(n234), .B(n233), .S(n275), .Z(n235) );
  MUX2_X1 U258 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n277), .Z(n236) );
  MUX2_X1 U259 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n277), .Z(n237) );
  MUX2_X1 U260 ( .A(n237), .B(n236), .S(n275), .Z(n238) );
  MUX2_X1 U261 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n239) );
  MUX2_X1 U262 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n277), .Z(n240) );
  MUX2_X1 U263 ( .A(n240), .B(n239), .S(n275), .Z(n241) );
  MUX2_X1 U264 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n277), .Z(n242) );
  MUX2_X1 U265 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n277), .Z(n243) );
  MUX2_X1 U266 ( .A(n243), .B(n242), .S(n275), .Z(n244) );
  MUX2_X1 U267 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n277), .Z(n245) );
  MUX2_X1 U268 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n246) );
  MUX2_X1 U269 ( .A(n246), .B(n245), .S(n275), .Z(n247) );
  MUX2_X1 U270 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n248) );
  MUX2_X1 U271 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n249) );
  MUX2_X1 U272 ( .A(n249), .B(n248), .S(n275), .Z(n250) );
  MUX2_X1 U273 ( .A(n250), .B(n247), .S(N12), .Z(N17) );
  MUX2_X1 U274 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(N10), .Z(n251) );
  MUX2_X1 U275 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n277), .Z(n252) );
  MUX2_X1 U276 ( .A(n252), .B(n251), .S(n275), .Z(n253) );
  MUX2_X1 U277 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n277), .Z(n254) );
  MUX2_X1 U278 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n277), .Z(n255) );
  MUX2_X1 U279 ( .A(n255), .B(n254), .S(n275), .Z(n256) );
  MUX2_X1 U280 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n277), .Z(n257) );
  MUX2_X1 U281 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(N10), .Z(n258) );
  MUX2_X1 U282 ( .A(n258), .B(n257), .S(n275), .Z(n259) );
  MUX2_X1 U283 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(N10), .Z(n260) );
  MUX2_X1 U284 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(N10), .Z(n261) );
  MUX2_X1 U285 ( .A(n261), .B(n260), .S(n275), .Z(n262) );
  MUX2_X1 U286 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(N10), .Z(n263) );
  MUX2_X1 U287 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(N10), .Z(n264) );
  MUX2_X1 U288 ( .A(n264), .B(n263), .S(n275), .Z(n265) );
  MUX2_X1 U289 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(N10), .Z(n266) );
  MUX2_X1 U290 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(N10), .Z(n267) );
  MUX2_X1 U291 ( .A(n267), .B(n266), .S(N11), .Z(n268) );
  MUX2_X1 U292 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n277), .Z(n269) );
  MUX2_X1 U293 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(N10), .Z(n270) );
  MUX2_X1 U294 ( .A(n270), .B(n269), .S(n275), .Z(n271) );
  MUX2_X1 U295 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(N10), .Z(n272) );
  MUX2_X1 U296 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(N10), .Z(n273) );
  MUX2_X1 U297 ( .A(n273), .B(n272), .S(N11), .Z(n274) );
endmodule


module memory_WIDTH12_SIZE8_LOGSIZE3_4 ( clk, data_in, data_out, addr, wr_en
 );
  input [11:0] data_in;
  output [11:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] ,
         \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] ,
         \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][11] , \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] ,
         \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] ,
         \mem[5][1] , \mem[5][0] , \mem[4][11] , \mem[4][10] , \mem[4][9] ,
         \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] ,
         \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] ,
         \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] ,
         \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][11] , \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] ,
         \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] ,
         \mem[0][1] , \mem[0][0] , N13, N14, N15, N17, N19, N20, N22, N23, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[11]  ( .D(N13), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N14), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N15), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[7]  ( .D(N17), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[5]  ( .D(N19), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N20), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N22), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N23), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \mem_reg[7][11]  ( .D(n293), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n294), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n295), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n296), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n297), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n298), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n299), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n300), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n301), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n302), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n303), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n304), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n305), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n306), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n307), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n308), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n309), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n310), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n311), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n312), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n313), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n314), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n315), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n316), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n317), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n318), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n319), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n320), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n321), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n322), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n323), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n324), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n325), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n326), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n327), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n328), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n329), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n330), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n331), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n332), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n333), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n334), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n335), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n336), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n337), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n338), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n339), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n340), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n341), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n342), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n343), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n344), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n345), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n346), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n347), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n348), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n349), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n350), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n351), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n352), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n353), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n354), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n355), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n356), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n357), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n358), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n359), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n360), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n361), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n362), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n363), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n364), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n365), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n366), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n367), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n368), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n369), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n370), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n371), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n372), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n373), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n374), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n375), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n376), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n377), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n378), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n379), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n380), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n381), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n382), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n383), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n384), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n385), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n386), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n387), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n388), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U212 ( .A1(n278), .A2(n279), .A3(n481), .ZN(n494) );
  NAND3_X1 U213 ( .A1(n481), .A2(n279), .A3(N10), .ZN(n480) );
  NAND3_X1 U214 ( .A1(n481), .A2(n278), .A3(N11), .ZN(n467) );
  NAND3_X1 U215 ( .A1(N10), .A2(n481), .A3(N11), .ZN(n454) );
  NAND3_X1 U216 ( .A1(n278), .A2(n279), .A3(n428), .ZN(n441) );
  NAND3_X1 U217 ( .A1(N10), .A2(n279), .A3(n428), .ZN(n427) );
  NAND3_X1 U218 ( .A1(N11), .A2(n278), .A3(n428), .ZN(n414) );
  NAND3_X1 U219 ( .A1(N11), .A2(N10), .A3(n428), .ZN(n401) );
  SDFF_X1 \data_out_reg[3]  ( .D(n226), .SI(n223), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[8]  ( .D(n256), .SI(n253), .SE(N12), .CK(clk), .Q(
        data_out[8]) );
  SDFF_X1 \data_out_reg[6]  ( .D(n244), .SI(n241), .SE(N12), .CK(clk), .Q(
        data_out[6]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n6), .SI(n3), .SE(N12), .CK(clk), .Q(
        data_out[0]) );
  BUF_X1 U3 ( .A(n277), .Z(n276) );
  BUF_X1 U4 ( .A(N11), .Z(n275) );
  BUF_X1 U5 ( .A(N10), .Z(n277) );
  NOR2_X1 U6 ( .A1(n280), .A2(N12), .ZN(n481) );
  INV_X1 U7 ( .A(wr_en), .ZN(n280) );
  AND2_X1 U8 ( .A1(N12), .A2(wr_en), .ZN(n428) );
  INV_X1 U9 ( .A(N10), .ZN(n278) );
  INV_X1 U10 ( .A(N11), .ZN(n279) );
  OAI21_X1 U11 ( .B1(n292), .B2(n480), .A(n479), .ZN(n376) );
  NAND2_X1 U12 ( .A1(\mem[1][0] ), .A2(n480), .ZN(n479) );
  OAI21_X1 U13 ( .B1(n291), .B2(n480), .A(n478), .ZN(n375) );
  NAND2_X1 U14 ( .A1(\mem[1][1] ), .A2(n480), .ZN(n478) );
  OAI21_X1 U15 ( .B1(n290), .B2(n480), .A(n477), .ZN(n374) );
  NAND2_X1 U16 ( .A1(\mem[1][2] ), .A2(n480), .ZN(n477) );
  OAI21_X1 U17 ( .B1(n289), .B2(n480), .A(n476), .ZN(n373) );
  NAND2_X1 U18 ( .A1(\mem[1][3] ), .A2(n480), .ZN(n476) );
  OAI21_X1 U19 ( .B1(n288), .B2(n480), .A(n475), .ZN(n372) );
  NAND2_X1 U20 ( .A1(\mem[1][4] ), .A2(n480), .ZN(n475) );
  OAI21_X1 U21 ( .B1(n287), .B2(n480), .A(n474), .ZN(n371) );
  NAND2_X1 U22 ( .A1(\mem[1][5] ), .A2(n480), .ZN(n474) );
  OAI21_X1 U23 ( .B1(n286), .B2(n480), .A(n473), .ZN(n370) );
  NAND2_X1 U24 ( .A1(\mem[1][6] ), .A2(n480), .ZN(n473) );
  OAI21_X1 U25 ( .B1(n285), .B2(n480), .A(n472), .ZN(n369) );
  NAND2_X1 U26 ( .A1(\mem[1][7] ), .A2(n480), .ZN(n472) );
  OAI21_X1 U27 ( .B1(n284), .B2(n480), .A(n471), .ZN(n368) );
  NAND2_X1 U28 ( .A1(\mem[1][8] ), .A2(n480), .ZN(n471) );
  OAI21_X1 U29 ( .B1(n283), .B2(n480), .A(n470), .ZN(n367) );
  NAND2_X1 U30 ( .A1(\mem[1][9] ), .A2(n480), .ZN(n470) );
  OAI21_X1 U31 ( .B1(n282), .B2(n480), .A(n469), .ZN(n366) );
  NAND2_X1 U32 ( .A1(\mem[1][10] ), .A2(n480), .ZN(n469) );
  OAI21_X1 U33 ( .B1(n281), .B2(n480), .A(n468), .ZN(n365) );
  NAND2_X1 U34 ( .A1(\mem[1][11] ), .A2(n480), .ZN(n468) );
  OAI21_X1 U35 ( .B1(n292), .B2(n467), .A(n466), .ZN(n364) );
  NAND2_X1 U36 ( .A1(\mem[2][0] ), .A2(n467), .ZN(n466) );
  OAI21_X1 U37 ( .B1(n291), .B2(n467), .A(n465), .ZN(n363) );
  NAND2_X1 U38 ( .A1(\mem[2][1] ), .A2(n467), .ZN(n465) );
  OAI21_X1 U39 ( .B1(n290), .B2(n467), .A(n464), .ZN(n362) );
  NAND2_X1 U40 ( .A1(\mem[2][2] ), .A2(n467), .ZN(n464) );
  OAI21_X1 U41 ( .B1(n289), .B2(n467), .A(n463), .ZN(n361) );
  NAND2_X1 U42 ( .A1(\mem[2][3] ), .A2(n467), .ZN(n463) );
  OAI21_X1 U43 ( .B1(n288), .B2(n467), .A(n462), .ZN(n360) );
  NAND2_X1 U44 ( .A1(\mem[2][4] ), .A2(n467), .ZN(n462) );
  OAI21_X1 U45 ( .B1(n287), .B2(n467), .A(n461), .ZN(n359) );
  NAND2_X1 U46 ( .A1(\mem[2][5] ), .A2(n467), .ZN(n461) );
  OAI21_X1 U47 ( .B1(n286), .B2(n467), .A(n460), .ZN(n358) );
  NAND2_X1 U48 ( .A1(\mem[2][6] ), .A2(n467), .ZN(n460) );
  OAI21_X1 U49 ( .B1(n285), .B2(n467), .A(n459), .ZN(n357) );
  NAND2_X1 U50 ( .A1(\mem[2][7] ), .A2(n467), .ZN(n459) );
  OAI21_X1 U51 ( .B1(n284), .B2(n467), .A(n458), .ZN(n356) );
  NAND2_X1 U52 ( .A1(\mem[2][8] ), .A2(n467), .ZN(n458) );
  OAI21_X1 U53 ( .B1(n283), .B2(n467), .A(n457), .ZN(n355) );
  NAND2_X1 U54 ( .A1(\mem[2][9] ), .A2(n467), .ZN(n457) );
  OAI21_X1 U55 ( .B1(n282), .B2(n467), .A(n456), .ZN(n354) );
  NAND2_X1 U56 ( .A1(\mem[2][10] ), .A2(n467), .ZN(n456) );
  OAI21_X1 U57 ( .B1(n281), .B2(n467), .A(n455), .ZN(n353) );
  NAND2_X1 U58 ( .A1(\mem[2][11] ), .A2(n467), .ZN(n455) );
  OAI21_X1 U59 ( .B1(n292), .B2(n454), .A(n453), .ZN(n352) );
  NAND2_X1 U60 ( .A1(\mem[3][0] ), .A2(n454), .ZN(n453) );
  OAI21_X1 U61 ( .B1(n291), .B2(n454), .A(n452), .ZN(n351) );
  NAND2_X1 U62 ( .A1(\mem[3][1] ), .A2(n454), .ZN(n452) );
  OAI21_X1 U63 ( .B1(n290), .B2(n454), .A(n451), .ZN(n350) );
  NAND2_X1 U64 ( .A1(\mem[3][2] ), .A2(n454), .ZN(n451) );
  OAI21_X1 U65 ( .B1(n289), .B2(n454), .A(n450), .ZN(n349) );
  NAND2_X1 U66 ( .A1(\mem[3][3] ), .A2(n454), .ZN(n450) );
  OAI21_X1 U67 ( .B1(n288), .B2(n454), .A(n449), .ZN(n348) );
  NAND2_X1 U68 ( .A1(\mem[3][4] ), .A2(n454), .ZN(n449) );
  OAI21_X1 U69 ( .B1(n287), .B2(n454), .A(n448), .ZN(n347) );
  NAND2_X1 U70 ( .A1(\mem[3][5] ), .A2(n454), .ZN(n448) );
  OAI21_X1 U71 ( .B1(n286), .B2(n454), .A(n447), .ZN(n346) );
  NAND2_X1 U72 ( .A1(\mem[3][6] ), .A2(n454), .ZN(n447) );
  OAI21_X1 U73 ( .B1(n285), .B2(n454), .A(n446), .ZN(n345) );
  NAND2_X1 U74 ( .A1(\mem[3][7] ), .A2(n454), .ZN(n446) );
  OAI21_X1 U75 ( .B1(n284), .B2(n454), .A(n445), .ZN(n344) );
  NAND2_X1 U76 ( .A1(\mem[3][8] ), .A2(n454), .ZN(n445) );
  OAI21_X1 U77 ( .B1(n283), .B2(n454), .A(n444), .ZN(n343) );
  NAND2_X1 U78 ( .A1(\mem[3][9] ), .A2(n454), .ZN(n444) );
  OAI21_X1 U79 ( .B1(n282), .B2(n454), .A(n443), .ZN(n342) );
  NAND2_X1 U80 ( .A1(\mem[3][10] ), .A2(n454), .ZN(n443) );
  OAI21_X1 U81 ( .B1(n281), .B2(n454), .A(n442), .ZN(n341) );
  NAND2_X1 U82 ( .A1(\mem[3][11] ), .A2(n454), .ZN(n442) );
  OAI21_X1 U83 ( .B1(n292), .B2(n441), .A(n440), .ZN(n340) );
  NAND2_X1 U84 ( .A1(\mem[4][0] ), .A2(n441), .ZN(n440) );
  OAI21_X1 U85 ( .B1(n291), .B2(n441), .A(n439), .ZN(n339) );
  NAND2_X1 U86 ( .A1(\mem[4][1] ), .A2(n441), .ZN(n439) );
  OAI21_X1 U87 ( .B1(n290), .B2(n441), .A(n438), .ZN(n338) );
  NAND2_X1 U88 ( .A1(\mem[4][2] ), .A2(n441), .ZN(n438) );
  OAI21_X1 U89 ( .B1(n289), .B2(n441), .A(n437), .ZN(n337) );
  NAND2_X1 U90 ( .A1(\mem[4][3] ), .A2(n441), .ZN(n437) );
  OAI21_X1 U91 ( .B1(n288), .B2(n441), .A(n436), .ZN(n336) );
  NAND2_X1 U92 ( .A1(\mem[4][4] ), .A2(n441), .ZN(n436) );
  OAI21_X1 U93 ( .B1(n287), .B2(n441), .A(n435), .ZN(n335) );
  NAND2_X1 U94 ( .A1(\mem[4][5] ), .A2(n441), .ZN(n435) );
  OAI21_X1 U95 ( .B1(n286), .B2(n441), .A(n434), .ZN(n334) );
  NAND2_X1 U96 ( .A1(\mem[4][6] ), .A2(n441), .ZN(n434) );
  OAI21_X1 U97 ( .B1(n285), .B2(n441), .A(n433), .ZN(n333) );
  NAND2_X1 U98 ( .A1(\mem[4][7] ), .A2(n441), .ZN(n433) );
  OAI21_X1 U99 ( .B1(n284), .B2(n441), .A(n432), .ZN(n332) );
  NAND2_X1 U100 ( .A1(\mem[4][8] ), .A2(n441), .ZN(n432) );
  OAI21_X1 U101 ( .B1(n283), .B2(n441), .A(n431), .ZN(n331) );
  NAND2_X1 U102 ( .A1(\mem[4][9] ), .A2(n441), .ZN(n431) );
  OAI21_X1 U103 ( .B1(n282), .B2(n441), .A(n430), .ZN(n330) );
  NAND2_X1 U104 ( .A1(\mem[4][10] ), .A2(n441), .ZN(n430) );
  OAI21_X1 U105 ( .B1(n281), .B2(n441), .A(n429), .ZN(n329) );
  NAND2_X1 U106 ( .A1(\mem[4][11] ), .A2(n441), .ZN(n429) );
  OAI21_X1 U107 ( .B1(n292), .B2(n427), .A(n426), .ZN(n328) );
  NAND2_X1 U108 ( .A1(\mem[5][0] ), .A2(n427), .ZN(n426) );
  OAI21_X1 U109 ( .B1(n291), .B2(n427), .A(n425), .ZN(n327) );
  NAND2_X1 U110 ( .A1(\mem[5][1] ), .A2(n427), .ZN(n425) );
  OAI21_X1 U111 ( .B1(n290), .B2(n427), .A(n424), .ZN(n326) );
  NAND2_X1 U112 ( .A1(\mem[5][2] ), .A2(n427), .ZN(n424) );
  OAI21_X1 U113 ( .B1(n289), .B2(n427), .A(n423), .ZN(n325) );
  NAND2_X1 U114 ( .A1(\mem[5][3] ), .A2(n427), .ZN(n423) );
  OAI21_X1 U115 ( .B1(n288), .B2(n427), .A(n422), .ZN(n324) );
  NAND2_X1 U116 ( .A1(\mem[5][4] ), .A2(n427), .ZN(n422) );
  OAI21_X1 U117 ( .B1(n287), .B2(n427), .A(n421), .ZN(n323) );
  NAND2_X1 U118 ( .A1(\mem[5][5] ), .A2(n427), .ZN(n421) );
  OAI21_X1 U119 ( .B1(n286), .B2(n427), .A(n420), .ZN(n322) );
  NAND2_X1 U120 ( .A1(\mem[5][6] ), .A2(n427), .ZN(n420) );
  OAI21_X1 U121 ( .B1(n285), .B2(n427), .A(n419), .ZN(n321) );
  NAND2_X1 U122 ( .A1(\mem[5][7] ), .A2(n427), .ZN(n419) );
  OAI21_X1 U123 ( .B1(n284), .B2(n427), .A(n418), .ZN(n320) );
  NAND2_X1 U124 ( .A1(\mem[5][8] ), .A2(n427), .ZN(n418) );
  OAI21_X1 U125 ( .B1(n283), .B2(n427), .A(n417), .ZN(n319) );
  NAND2_X1 U126 ( .A1(\mem[5][9] ), .A2(n427), .ZN(n417) );
  OAI21_X1 U127 ( .B1(n282), .B2(n427), .A(n416), .ZN(n318) );
  NAND2_X1 U128 ( .A1(\mem[5][10] ), .A2(n427), .ZN(n416) );
  OAI21_X1 U129 ( .B1(n281), .B2(n427), .A(n415), .ZN(n317) );
  NAND2_X1 U130 ( .A1(\mem[5][11] ), .A2(n427), .ZN(n415) );
  OAI21_X1 U131 ( .B1(n292), .B2(n414), .A(n413), .ZN(n316) );
  NAND2_X1 U132 ( .A1(\mem[6][0] ), .A2(n414), .ZN(n413) );
  OAI21_X1 U133 ( .B1(n291), .B2(n414), .A(n412), .ZN(n315) );
  NAND2_X1 U134 ( .A1(\mem[6][1] ), .A2(n414), .ZN(n412) );
  OAI21_X1 U135 ( .B1(n290), .B2(n414), .A(n411), .ZN(n314) );
  NAND2_X1 U136 ( .A1(\mem[6][2] ), .A2(n414), .ZN(n411) );
  OAI21_X1 U137 ( .B1(n289), .B2(n414), .A(n410), .ZN(n313) );
  NAND2_X1 U138 ( .A1(\mem[6][3] ), .A2(n414), .ZN(n410) );
  OAI21_X1 U139 ( .B1(n288), .B2(n414), .A(n409), .ZN(n312) );
  NAND2_X1 U140 ( .A1(\mem[6][4] ), .A2(n414), .ZN(n409) );
  OAI21_X1 U141 ( .B1(n287), .B2(n414), .A(n408), .ZN(n311) );
  NAND2_X1 U142 ( .A1(\mem[6][5] ), .A2(n414), .ZN(n408) );
  OAI21_X1 U143 ( .B1(n286), .B2(n414), .A(n407), .ZN(n310) );
  NAND2_X1 U144 ( .A1(\mem[6][6] ), .A2(n414), .ZN(n407) );
  OAI21_X1 U145 ( .B1(n285), .B2(n414), .A(n406), .ZN(n309) );
  NAND2_X1 U146 ( .A1(\mem[6][7] ), .A2(n414), .ZN(n406) );
  OAI21_X1 U147 ( .B1(n284), .B2(n414), .A(n405), .ZN(n308) );
  NAND2_X1 U148 ( .A1(\mem[6][8] ), .A2(n414), .ZN(n405) );
  OAI21_X1 U149 ( .B1(n283), .B2(n414), .A(n404), .ZN(n307) );
  NAND2_X1 U150 ( .A1(\mem[6][9] ), .A2(n414), .ZN(n404) );
  OAI21_X1 U151 ( .B1(n282), .B2(n414), .A(n403), .ZN(n306) );
  NAND2_X1 U152 ( .A1(\mem[6][10] ), .A2(n414), .ZN(n403) );
  OAI21_X1 U153 ( .B1(n281), .B2(n414), .A(n402), .ZN(n305) );
  NAND2_X1 U154 ( .A1(\mem[6][11] ), .A2(n414), .ZN(n402) );
  OAI21_X1 U155 ( .B1(n292), .B2(n401), .A(n400), .ZN(n304) );
  NAND2_X1 U156 ( .A1(\mem[7][0] ), .A2(n401), .ZN(n400) );
  OAI21_X1 U157 ( .B1(n291), .B2(n401), .A(n399), .ZN(n303) );
  NAND2_X1 U158 ( .A1(\mem[7][1] ), .A2(n401), .ZN(n399) );
  OAI21_X1 U159 ( .B1(n290), .B2(n401), .A(n398), .ZN(n302) );
  NAND2_X1 U160 ( .A1(\mem[7][2] ), .A2(n401), .ZN(n398) );
  OAI21_X1 U161 ( .B1(n289), .B2(n401), .A(n397), .ZN(n301) );
  NAND2_X1 U162 ( .A1(\mem[7][3] ), .A2(n401), .ZN(n397) );
  OAI21_X1 U163 ( .B1(n288), .B2(n401), .A(n396), .ZN(n300) );
  NAND2_X1 U164 ( .A1(\mem[7][4] ), .A2(n401), .ZN(n396) );
  OAI21_X1 U165 ( .B1(n287), .B2(n401), .A(n395), .ZN(n299) );
  NAND2_X1 U166 ( .A1(\mem[7][5] ), .A2(n401), .ZN(n395) );
  OAI21_X1 U167 ( .B1(n286), .B2(n401), .A(n394), .ZN(n298) );
  NAND2_X1 U168 ( .A1(\mem[7][6] ), .A2(n401), .ZN(n394) );
  OAI21_X1 U169 ( .B1(n285), .B2(n401), .A(n393), .ZN(n297) );
  NAND2_X1 U170 ( .A1(\mem[7][7] ), .A2(n401), .ZN(n393) );
  OAI21_X1 U171 ( .B1(n284), .B2(n401), .A(n392), .ZN(n296) );
  NAND2_X1 U172 ( .A1(\mem[7][8] ), .A2(n401), .ZN(n392) );
  OAI21_X1 U173 ( .B1(n283), .B2(n401), .A(n391), .ZN(n295) );
  NAND2_X1 U174 ( .A1(\mem[7][9] ), .A2(n401), .ZN(n391) );
  OAI21_X1 U175 ( .B1(n282), .B2(n401), .A(n390), .ZN(n294) );
  NAND2_X1 U176 ( .A1(\mem[7][10] ), .A2(n401), .ZN(n390) );
  OAI21_X1 U177 ( .B1(n281), .B2(n401), .A(n389), .ZN(n293) );
  NAND2_X1 U178 ( .A1(\mem[7][11] ), .A2(n401), .ZN(n389) );
  OAI21_X1 U179 ( .B1(n494), .B2(n292), .A(n493), .ZN(n388) );
  NAND2_X1 U180 ( .A1(\mem[0][0] ), .A2(n494), .ZN(n493) );
  OAI21_X1 U181 ( .B1(n494), .B2(n291), .A(n492), .ZN(n387) );
  NAND2_X1 U182 ( .A1(\mem[0][1] ), .A2(n494), .ZN(n492) );
  OAI21_X1 U183 ( .B1(n494), .B2(n290), .A(n491), .ZN(n386) );
  NAND2_X1 U184 ( .A1(\mem[0][2] ), .A2(n494), .ZN(n491) );
  OAI21_X1 U185 ( .B1(n494), .B2(n289), .A(n490), .ZN(n385) );
  NAND2_X1 U186 ( .A1(\mem[0][3] ), .A2(n494), .ZN(n490) );
  OAI21_X1 U187 ( .B1(n494), .B2(n288), .A(n489), .ZN(n384) );
  NAND2_X1 U188 ( .A1(\mem[0][4] ), .A2(n494), .ZN(n489) );
  OAI21_X1 U189 ( .B1(n494), .B2(n287), .A(n488), .ZN(n383) );
  NAND2_X1 U190 ( .A1(\mem[0][5] ), .A2(n494), .ZN(n488) );
  OAI21_X1 U191 ( .B1(n494), .B2(n286), .A(n487), .ZN(n382) );
  NAND2_X1 U192 ( .A1(\mem[0][6] ), .A2(n494), .ZN(n487) );
  OAI21_X1 U193 ( .B1(n494), .B2(n285), .A(n486), .ZN(n381) );
  NAND2_X1 U194 ( .A1(\mem[0][7] ), .A2(n494), .ZN(n486) );
  OAI21_X1 U195 ( .B1(n494), .B2(n284), .A(n485), .ZN(n380) );
  NAND2_X1 U196 ( .A1(\mem[0][8] ), .A2(n494), .ZN(n485) );
  OAI21_X1 U197 ( .B1(n494), .B2(n283), .A(n484), .ZN(n379) );
  NAND2_X1 U198 ( .A1(\mem[0][9] ), .A2(n494), .ZN(n484) );
  OAI21_X1 U199 ( .B1(n494), .B2(n282), .A(n483), .ZN(n378) );
  NAND2_X1 U200 ( .A1(\mem[0][10] ), .A2(n494), .ZN(n483) );
  OAI21_X1 U201 ( .B1(n494), .B2(n281), .A(n482), .ZN(n377) );
  NAND2_X1 U202 ( .A1(\mem[0][11] ), .A2(n494), .ZN(n482) );
  INV_X1 U203 ( .A(data_in[0]), .ZN(n292) );
  INV_X1 U204 ( .A(data_in[1]), .ZN(n291) );
  INV_X1 U205 ( .A(data_in[2]), .ZN(n290) );
  INV_X1 U206 ( .A(data_in[3]), .ZN(n289) );
  INV_X1 U207 ( .A(data_in[4]), .ZN(n288) );
  INV_X1 U208 ( .A(data_in[5]), .ZN(n287) );
  INV_X1 U209 ( .A(data_in[6]), .ZN(n286) );
  INV_X1 U210 ( .A(data_in[7]), .ZN(n285) );
  INV_X1 U211 ( .A(data_in[8]), .ZN(n284) );
  INV_X1 U220 ( .A(data_in[9]), .ZN(n283) );
  INV_X1 U221 ( .A(data_in[10]), .ZN(n282) );
  INV_X1 U222 ( .A(data_in[11]), .ZN(n281) );
  MUX2_X1 U223 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n276), .Z(n1) );
  MUX2_X1 U224 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n276), .Z(n2) );
  MUX2_X1 U225 ( .A(n2), .B(n1), .S(n275), .Z(n3) );
  MUX2_X1 U226 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n276), .Z(n4) );
  MUX2_X1 U227 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n276), .Z(n5) );
  MUX2_X1 U228 ( .A(n5), .B(n4), .S(n275), .Z(n6) );
  MUX2_X1 U229 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n276), .Z(n7) );
  MUX2_X1 U230 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n276), .Z(n8) );
  MUX2_X1 U231 ( .A(n8), .B(n7), .S(n275), .Z(n9) );
  MUX2_X1 U232 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n276), .Z(n10) );
  MUX2_X1 U233 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n276), .Z(n11) );
  MUX2_X1 U234 ( .A(n11), .B(n10), .S(n275), .Z(n12) );
  MUX2_X1 U235 ( .A(n12), .B(n9), .S(N12), .Z(N23) );
  MUX2_X1 U236 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n276), .Z(n13) );
  MUX2_X1 U237 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n276), .Z(n14) );
  MUX2_X1 U238 ( .A(n14), .B(n13), .S(n275), .Z(n15) );
  MUX2_X1 U239 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n276), .Z(n218) );
  MUX2_X1 U240 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n276), .Z(n219) );
  MUX2_X1 U241 ( .A(n219), .B(n218), .S(n275), .Z(n220) );
  MUX2_X1 U242 ( .A(n220), .B(n15), .S(N12), .Z(N22) );
  MUX2_X1 U243 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n277), .Z(n221) );
  MUX2_X1 U244 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n277), .Z(n222) );
  MUX2_X1 U245 ( .A(n222), .B(n221), .S(n275), .Z(n223) );
  MUX2_X1 U246 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n277), .Z(n224) );
  MUX2_X1 U247 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n277), .Z(n225) );
  MUX2_X1 U248 ( .A(n225), .B(n224), .S(n275), .Z(n226) );
  MUX2_X1 U249 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n277), .Z(n227) );
  MUX2_X1 U250 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n277), .Z(n228) );
  MUX2_X1 U251 ( .A(n228), .B(n227), .S(n275), .Z(n229) );
  MUX2_X1 U252 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n277), .Z(n230) );
  MUX2_X1 U253 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n277), .Z(n231) );
  MUX2_X1 U254 ( .A(n231), .B(n230), .S(n275), .Z(n232) );
  MUX2_X1 U255 ( .A(n232), .B(n229), .S(N12), .Z(N20) );
  MUX2_X1 U256 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n277), .Z(n233) );
  MUX2_X1 U257 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n277), .Z(n234) );
  MUX2_X1 U258 ( .A(n234), .B(n233), .S(n275), .Z(n235) );
  MUX2_X1 U259 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n277), .Z(n236) );
  MUX2_X1 U260 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n277), .Z(n237) );
  MUX2_X1 U261 ( .A(n237), .B(n236), .S(n275), .Z(n238) );
  MUX2_X1 U262 ( .A(n238), .B(n235), .S(N12), .Z(N19) );
  MUX2_X1 U263 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n239) );
  MUX2_X1 U264 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n277), .Z(n240) );
  MUX2_X1 U265 ( .A(n240), .B(n239), .S(n275), .Z(n241) );
  MUX2_X1 U266 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n277), .Z(n242) );
  MUX2_X1 U267 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n277), .Z(n243) );
  MUX2_X1 U268 ( .A(n243), .B(n242), .S(N11), .Z(n244) );
  MUX2_X1 U269 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n277), .Z(n245) );
  MUX2_X1 U270 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n246) );
  MUX2_X1 U271 ( .A(n246), .B(n245), .S(n275), .Z(n247) );
  MUX2_X1 U272 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n248) );
  MUX2_X1 U273 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n249) );
  MUX2_X1 U274 ( .A(n249), .B(n248), .S(n275), .Z(n250) );
  MUX2_X1 U275 ( .A(n250), .B(n247), .S(N12), .Z(N17) );
  MUX2_X1 U276 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n277), .Z(n251) );
  MUX2_X1 U277 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n277), .Z(n252) );
  MUX2_X1 U278 ( .A(n252), .B(n251), .S(n275), .Z(n253) );
  MUX2_X1 U279 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n277), .Z(n254) );
  MUX2_X1 U280 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n277), .Z(n255) );
  MUX2_X1 U281 ( .A(n255), .B(n254), .S(N11), .Z(n256) );
  MUX2_X1 U282 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(N10), .Z(n257) );
  MUX2_X1 U283 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(N10), .Z(n258) );
  MUX2_X1 U284 ( .A(n258), .B(n257), .S(n275), .Z(n259) );
  MUX2_X1 U285 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(N10), .Z(n260) );
  MUX2_X1 U286 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(N10), .Z(n261) );
  MUX2_X1 U287 ( .A(n261), .B(n260), .S(n275), .Z(n262) );
  MUX2_X1 U288 ( .A(n262), .B(n259), .S(N12), .Z(N15) );
  MUX2_X1 U289 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(N10), .Z(n263) );
  MUX2_X1 U290 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(N10), .Z(n264) );
  MUX2_X1 U291 ( .A(n264), .B(n263), .S(n275), .Z(n265) );
  MUX2_X1 U292 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(N10), .Z(n266) );
  MUX2_X1 U293 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(N10), .Z(n267) );
  MUX2_X1 U294 ( .A(n267), .B(n266), .S(n275), .Z(n268) );
  MUX2_X1 U295 ( .A(n268), .B(n265), .S(N12), .Z(N14) );
  MUX2_X1 U296 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n277), .Z(n269) );
  MUX2_X1 U297 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(N10), .Z(n270) );
  MUX2_X1 U298 ( .A(n270), .B(n269), .S(n275), .Z(n271) );
  MUX2_X1 U299 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(N10), .Z(n272) );
  MUX2_X1 U300 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(N10), .Z(n273) );
  MUX2_X1 U301 ( .A(n273), .B(n272), .S(n275), .Z(n274) );
  MUX2_X1 U302 ( .A(n274), .B(n271), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH12_SIZE8_LOGSIZE3_3 ( clk, data_in, data_out, addr, wr_en
 );
  input [11:0] data_in;
  output [11:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] ,
         \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] ,
         \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][11] , \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] ,
         \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] ,
         \mem[5][1] , \mem[5][0] , \mem[4][11] , \mem[4][10] , \mem[4][9] ,
         \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] ,
         \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] ,
         \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] ,
         \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][11] , \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] ,
         \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] ,
         \mem[0][1] , \mem[0][0] , N13, N17, N19, N21, N24, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[11]  ( .D(N13), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[7]  ( .D(N17), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[5]  ( .D(N19), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[3]  ( .D(N21), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[0]  ( .D(N24), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][11]  ( .D(n293), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n294), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n295), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n296), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n297), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n298), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n299), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n300), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n301), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n302), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n303), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n304), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n305), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n306), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n307), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n308), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n309), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n310), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n311), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n312), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n313), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n314), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n315), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n316), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n317), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n318), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n319), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n320), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n321), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n322), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n323), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n324), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n325), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n326), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n327), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n328), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n329), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n330), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n331), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n332), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n333), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n334), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n335), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n336), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n337), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n338), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n339), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n340), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n341), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n342), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n343), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n344), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n345), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n346), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n347), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n348), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n349), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n350), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n351), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n352), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n353), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n354), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n355), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n356), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n357), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n358), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n359), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n360), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n361), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n362), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n363), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n364), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n365), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n366), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n367), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n368), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n369), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n370), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n371), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n372), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n373), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n374), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n375), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n376), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n377), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n378), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n379), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n380), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n381), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n382), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n383), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n384), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n385), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n386), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n387), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n388), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U212 ( .A1(n278), .A2(n279), .A3(n481), .ZN(n494) );
  NAND3_X1 U213 ( .A1(n481), .A2(n279), .A3(N10), .ZN(n480) );
  NAND3_X1 U214 ( .A1(n481), .A2(n278), .A3(N11), .ZN(n467) );
  NAND3_X1 U215 ( .A1(N10), .A2(n481), .A3(N11), .ZN(n454) );
  NAND3_X1 U216 ( .A1(n278), .A2(n279), .A3(n428), .ZN(n441) );
  NAND3_X1 U217 ( .A1(N10), .A2(n279), .A3(n428), .ZN(n427) );
  NAND3_X1 U218 ( .A1(N11), .A2(n278), .A3(n428), .ZN(n414) );
  NAND3_X1 U219 ( .A1(N11), .A2(N10), .A3(n428), .ZN(n401) );
  SDFF_X1 \data_out_reg[1]  ( .D(n12), .SI(n9), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[10]  ( .D(n268), .SI(n265), .SE(N12), .CK(clk), .Q(
        data_out[10]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n262), .SI(n259), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[8]  ( .D(n256), .SI(n253), .SE(N12), .CK(clk), .Q(
        data_out[8]) );
  SDFF_X1 \data_out_reg[4]  ( .D(n232), .SI(n229), .SE(N12), .CK(clk), .Q(
        data_out[4]) );
  SDFF_X1 \data_out_reg[2]  ( .D(n220), .SI(n15), .SE(N12), .CK(clk), .Q(
        data_out[2]) );
  SDFF_X1 \data_out_reg[6]  ( .D(n244), .SI(n241), .SE(N12), .CK(clk), .Q(
        data_out[6]) );
  BUF_X1 U3 ( .A(n277), .Z(n276) );
  BUF_X1 U4 ( .A(N11), .Z(n275) );
  BUF_X1 U5 ( .A(N10), .Z(n277) );
  NOR2_X1 U6 ( .A1(n280), .A2(N12), .ZN(n481) );
  INV_X1 U7 ( .A(wr_en), .ZN(n280) );
  AND2_X1 U8 ( .A1(N12), .A2(wr_en), .ZN(n428) );
  INV_X1 U9 ( .A(N10), .ZN(n278) );
  INV_X1 U10 ( .A(N11), .ZN(n279) );
  OAI21_X1 U11 ( .B1(n292), .B2(n480), .A(n479), .ZN(n376) );
  NAND2_X1 U12 ( .A1(\mem[1][0] ), .A2(n480), .ZN(n479) );
  OAI21_X1 U13 ( .B1(n291), .B2(n480), .A(n478), .ZN(n375) );
  NAND2_X1 U14 ( .A1(\mem[1][1] ), .A2(n480), .ZN(n478) );
  OAI21_X1 U15 ( .B1(n290), .B2(n480), .A(n477), .ZN(n374) );
  NAND2_X1 U16 ( .A1(\mem[1][2] ), .A2(n480), .ZN(n477) );
  OAI21_X1 U17 ( .B1(n289), .B2(n480), .A(n476), .ZN(n373) );
  NAND2_X1 U18 ( .A1(\mem[1][3] ), .A2(n480), .ZN(n476) );
  OAI21_X1 U19 ( .B1(n288), .B2(n480), .A(n475), .ZN(n372) );
  NAND2_X1 U20 ( .A1(\mem[1][4] ), .A2(n480), .ZN(n475) );
  OAI21_X1 U21 ( .B1(n287), .B2(n480), .A(n474), .ZN(n371) );
  NAND2_X1 U22 ( .A1(\mem[1][5] ), .A2(n480), .ZN(n474) );
  OAI21_X1 U23 ( .B1(n286), .B2(n480), .A(n473), .ZN(n370) );
  NAND2_X1 U24 ( .A1(\mem[1][6] ), .A2(n480), .ZN(n473) );
  OAI21_X1 U25 ( .B1(n285), .B2(n480), .A(n472), .ZN(n369) );
  NAND2_X1 U26 ( .A1(\mem[1][7] ), .A2(n480), .ZN(n472) );
  OAI21_X1 U27 ( .B1(n284), .B2(n480), .A(n471), .ZN(n368) );
  NAND2_X1 U28 ( .A1(\mem[1][8] ), .A2(n480), .ZN(n471) );
  OAI21_X1 U29 ( .B1(n283), .B2(n480), .A(n470), .ZN(n367) );
  NAND2_X1 U30 ( .A1(\mem[1][9] ), .A2(n480), .ZN(n470) );
  OAI21_X1 U31 ( .B1(n282), .B2(n480), .A(n469), .ZN(n366) );
  NAND2_X1 U32 ( .A1(\mem[1][10] ), .A2(n480), .ZN(n469) );
  OAI21_X1 U33 ( .B1(n281), .B2(n480), .A(n468), .ZN(n365) );
  NAND2_X1 U34 ( .A1(\mem[1][11] ), .A2(n480), .ZN(n468) );
  OAI21_X1 U35 ( .B1(n292), .B2(n467), .A(n466), .ZN(n364) );
  NAND2_X1 U36 ( .A1(\mem[2][0] ), .A2(n467), .ZN(n466) );
  OAI21_X1 U37 ( .B1(n291), .B2(n467), .A(n465), .ZN(n363) );
  NAND2_X1 U38 ( .A1(\mem[2][1] ), .A2(n467), .ZN(n465) );
  OAI21_X1 U39 ( .B1(n290), .B2(n467), .A(n464), .ZN(n362) );
  NAND2_X1 U40 ( .A1(\mem[2][2] ), .A2(n467), .ZN(n464) );
  OAI21_X1 U41 ( .B1(n289), .B2(n467), .A(n463), .ZN(n361) );
  NAND2_X1 U42 ( .A1(\mem[2][3] ), .A2(n467), .ZN(n463) );
  OAI21_X1 U43 ( .B1(n288), .B2(n467), .A(n462), .ZN(n360) );
  NAND2_X1 U44 ( .A1(\mem[2][4] ), .A2(n467), .ZN(n462) );
  OAI21_X1 U45 ( .B1(n287), .B2(n467), .A(n461), .ZN(n359) );
  NAND2_X1 U46 ( .A1(\mem[2][5] ), .A2(n467), .ZN(n461) );
  OAI21_X1 U47 ( .B1(n286), .B2(n467), .A(n460), .ZN(n358) );
  NAND2_X1 U48 ( .A1(\mem[2][6] ), .A2(n467), .ZN(n460) );
  OAI21_X1 U49 ( .B1(n285), .B2(n467), .A(n459), .ZN(n357) );
  NAND2_X1 U50 ( .A1(\mem[2][7] ), .A2(n467), .ZN(n459) );
  OAI21_X1 U51 ( .B1(n284), .B2(n467), .A(n458), .ZN(n356) );
  NAND2_X1 U52 ( .A1(\mem[2][8] ), .A2(n467), .ZN(n458) );
  OAI21_X1 U53 ( .B1(n283), .B2(n467), .A(n457), .ZN(n355) );
  NAND2_X1 U54 ( .A1(\mem[2][9] ), .A2(n467), .ZN(n457) );
  OAI21_X1 U55 ( .B1(n282), .B2(n467), .A(n456), .ZN(n354) );
  NAND2_X1 U56 ( .A1(\mem[2][10] ), .A2(n467), .ZN(n456) );
  OAI21_X1 U57 ( .B1(n281), .B2(n467), .A(n455), .ZN(n353) );
  NAND2_X1 U58 ( .A1(\mem[2][11] ), .A2(n467), .ZN(n455) );
  OAI21_X1 U59 ( .B1(n292), .B2(n454), .A(n453), .ZN(n352) );
  NAND2_X1 U60 ( .A1(\mem[3][0] ), .A2(n454), .ZN(n453) );
  OAI21_X1 U61 ( .B1(n291), .B2(n454), .A(n452), .ZN(n351) );
  NAND2_X1 U62 ( .A1(\mem[3][1] ), .A2(n454), .ZN(n452) );
  OAI21_X1 U63 ( .B1(n290), .B2(n454), .A(n451), .ZN(n350) );
  NAND2_X1 U64 ( .A1(\mem[3][2] ), .A2(n454), .ZN(n451) );
  OAI21_X1 U65 ( .B1(n289), .B2(n454), .A(n450), .ZN(n349) );
  NAND2_X1 U66 ( .A1(\mem[3][3] ), .A2(n454), .ZN(n450) );
  OAI21_X1 U67 ( .B1(n288), .B2(n454), .A(n449), .ZN(n348) );
  NAND2_X1 U68 ( .A1(\mem[3][4] ), .A2(n454), .ZN(n449) );
  OAI21_X1 U69 ( .B1(n287), .B2(n454), .A(n448), .ZN(n347) );
  NAND2_X1 U70 ( .A1(\mem[3][5] ), .A2(n454), .ZN(n448) );
  OAI21_X1 U71 ( .B1(n286), .B2(n454), .A(n447), .ZN(n346) );
  NAND2_X1 U72 ( .A1(\mem[3][6] ), .A2(n454), .ZN(n447) );
  OAI21_X1 U73 ( .B1(n285), .B2(n454), .A(n446), .ZN(n345) );
  NAND2_X1 U74 ( .A1(\mem[3][7] ), .A2(n454), .ZN(n446) );
  OAI21_X1 U75 ( .B1(n284), .B2(n454), .A(n445), .ZN(n344) );
  NAND2_X1 U76 ( .A1(\mem[3][8] ), .A2(n454), .ZN(n445) );
  OAI21_X1 U77 ( .B1(n283), .B2(n454), .A(n444), .ZN(n343) );
  NAND2_X1 U78 ( .A1(\mem[3][9] ), .A2(n454), .ZN(n444) );
  OAI21_X1 U79 ( .B1(n282), .B2(n454), .A(n443), .ZN(n342) );
  NAND2_X1 U80 ( .A1(\mem[3][10] ), .A2(n454), .ZN(n443) );
  OAI21_X1 U81 ( .B1(n281), .B2(n454), .A(n442), .ZN(n341) );
  NAND2_X1 U82 ( .A1(\mem[3][11] ), .A2(n454), .ZN(n442) );
  OAI21_X1 U83 ( .B1(n292), .B2(n441), .A(n440), .ZN(n340) );
  NAND2_X1 U84 ( .A1(\mem[4][0] ), .A2(n441), .ZN(n440) );
  OAI21_X1 U85 ( .B1(n291), .B2(n441), .A(n439), .ZN(n339) );
  NAND2_X1 U86 ( .A1(\mem[4][1] ), .A2(n441), .ZN(n439) );
  OAI21_X1 U87 ( .B1(n290), .B2(n441), .A(n438), .ZN(n338) );
  NAND2_X1 U88 ( .A1(\mem[4][2] ), .A2(n441), .ZN(n438) );
  OAI21_X1 U89 ( .B1(n289), .B2(n441), .A(n437), .ZN(n337) );
  NAND2_X1 U90 ( .A1(\mem[4][3] ), .A2(n441), .ZN(n437) );
  OAI21_X1 U91 ( .B1(n288), .B2(n441), .A(n436), .ZN(n336) );
  NAND2_X1 U92 ( .A1(\mem[4][4] ), .A2(n441), .ZN(n436) );
  OAI21_X1 U93 ( .B1(n287), .B2(n441), .A(n435), .ZN(n335) );
  NAND2_X1 U94 ( .A1(\mem[4][5] ), .A2(n441), .ZN(n435) );
  OAI21_X1 U95 ( .B1(n286), .B2(n441), .A(n434), .ZN(n334) );
  NAND2_X1 U96 ( .A1(\mem[4][6] ), .A2(n441), .ZN(n434) );
  OAI21_X1 U97 ( .B1(n285), .B2(n441), .A(n433), .ZN(n333) );
  NAND2_X1 U98 ( .A1(\mem[4][7] ), .A2(n441), .ZN(n433) );
  OAI21_X1 U99 ( .B1(n284), .B2(n441), .A(n432), .ZN(n332) );
  NAND2_X1 U100 ( .A1(\mem[4][8] ), .A2(n441), .ZN(n432) );
  OAI21_X1 U101 ( .B1(n283), .B2(n441), .A(n431), .ZN(n331) );
  NAND2_X1 U102 ( .A1(\mem[4][9] ), .A2(n441), .ZN(n431) );
  OAI21_X1 U103 ( .B1(n282), .B2(n441), .A(n430), .ZN(n330) );
  NAND2_X1 U104 ( .A1(\mem[4][10] ), .A2(n441), .ZN(n430) );
  OAI21_X1 U105 ( .B1(n281), .B2(n441), .A(n429), .ZN(n329) );
  NAND2_X1 U106 ( .A1(\mem[4][11] ), .A2(n441), .ZN(n429) );
  OAI21_X1 U107 ( .B1(n292), .B2(n427), .A(n426), .ZN(n328) );
  NAND2_X1 U108 ( .A1(\mem[5][0] ), .A2(n427), .ZN(n426) );
  OAI21_X1 U109 ( .B1(n291), .B2(n427), .A(n425), .ZN(n327) );
  NAND2_X1 U110 ( .A1(\mem[5][1] ), .A2(n427), .ZN(n425) );
  OAI21_X1 U111 ( .B1(n290), .B2(n427), .A(n424), .ZN(n326) );
  NAND2_X1 U112 ( .A1(\mem[5][2] ), .A2(n427), .ZN(n424) );
  OAI21_X1 U113 ( .B1(n289), .B2(n427), .A(n423), .ZN(n325) );
  NAND2_X1 U114 ( .A1(\mem[5][3] ), .A2(n427), .ZN(n423) );
  OAI21_X1 U115 ( .B1(n288), .B2(n427), .A(n422), .ZN(n324) );
  NAND2_X1 U116 ( .A1(\mem[5][4] ), .A2(n427), .ZN(n422) );
  OAI21_X1 U117 ( .B1(n287), .B2(n427), .A(n421), .ZN(n323) );
  NAND2_X1 U118 ( .A1(\mem[5][5] ), .A2(n427), .ZN(n421) );
  OAI21_X1 U119 ( .B1(n286), .B2(n427), .A(n420), .ZN(n322) );
  NAND2_X1 U120 ( .A1(\mem[5][6] ), .A2(n427), .ZN(n420) );
  OAI21_X1 U121 ( .B1(n285), .B2(n427), .A(n419), .ZN(n321) );
  NAND2_X1 U122 ( .A1(\mem[5][7] ), .A2(n427), .ZN(n419) );
  OAI21_X1 U123 ( .B1(n284), .B2(n427), .A(n418), .ZN(n320) );
  NAND2_X1 U124 ( .A1(\mem[5][8] ), .A2(n427), .ZN(n418) );
  OAI21_X1 U125 ( .B1(n283), .B2(n427), .A(n417), .ZN(n319) );
  NAND2_X1 U126 ( .A1(\mem[5][9] ), .A2(n427), .ZN(n417) );
  OAI21_X1 U127 ( .B1(n282), .B2(n427), .A(n416), .ZN(n318) );
  NAND2_X1 U128 ( .A1(\mem[5][10] ), .A2(n427), .ZN(n416) );
  OAI21_X1 U129 ( .B1(n281), .B2(n427), .A(n415), .ZN(n317) );
  NAND2_X1 U130 ( .A1(\mem[5][11] ), .A2(n427), .ZN(n415) );
  OAI21_X1 U131 ( .B1(n292), .B2(n414), .A(n413), .ZN(n316) );
  NAND2_X1 U132 ( .A1(\mem[6][0] ), .A2(n414), .ZN(n413) );
  OAI21_X1 U133 ( .B1(n291), .B2(n414), .A(n412), .ZN(n315) );
  NAND2_X1 U134 ( .A1(\mem[6][1] ), .A2(n414), .ZN(n412) );
  OAI21_X1 U135 ( .B1(n290), .B2(n414), .A(n411), .ZN(n314) );
  NAND2_X1 U136 ( .A1(\mem[6][2] ), .A2(n414), .ZN(n411) );
  OAI21_X1 U137 ( .B1(n289), .B2(n414), .A(n410), .ZN(n313) );
  NAND2_X1 U138 ( .A1(\mem[6][3] ), .A2(n414), .ZN(n410) );
  OAI21_X1 U139 ( .B1(n288), .B2(n414), .A(n409), .ZN(n312) );
  NAND2_X1 U140 ( .A1(\mem[6][4] ), .A2(n414), .ZN(n409) );
  OAI21_X1 U141 ( .B1(n287), .B2(n414), .A(n408), .ZN(n311) );
  NAND2_X1 U142 ( .A1(\mem[6][5] ), .A2(n414), .ZN(n408) );
  OAI21_X1 U143 ( .B1(n286), .B2(n414), .A(n407), .ZN(n310) );
  NAND2_X1 U144 ( .A1(\mem[6][6] ), .A2(n414), .ZN(n407) );
  OAI21_X1 U145 ( .B1(n285), .B2(n414), .A(n406), .ZN(n309) );
  NAND2_X1 U146 ( .A1(\mem[6][7] ), .A2(n414), .ZN(n406) );
  OAI21_X1 U147 ( .B1(n284), .B2(n414), .A(n405), .ZN(n308) );
  NAND2_X1 U148 ( .A1(\mem[6][8] ), .A2(n414), .ZN(n405) );
  OAI21_X1 U149 ( .B1(n283), .B2(n414), .A(n404), .ZN(n307) );
  NAND2_X1 U150 ( .A1(\mem[6][9] ), .A2(n414), .ZN(n404) );
  OAI21_X1 U151 ( .B1(n282), .B2(n414), .A(n403), .ZN(n306) );
  NAND2_X1 U152 ( .A1(\mem[6][10] ), .A2(n414), .ZN(n403) );
  OAI21_X1 U153 ( .B1(n281), .B2(n414), .A(n402), .ZN(n305) );
  NAND2_X1 U154 ( .A1(\mem[6][11] ), .A2(n414), .ZN(n402) );
  OAI21_X1 U155 ( .B1(n292), .B2(n401), .A(n400), .ZN(n304) );
  NAND2_X1 U156 ( .A1(\mem[7][0] ), .A2(n401), .ZN(n400) );
  OAI21_X1 U157 ( .B1(n291), .B2(n401), .A(n399), .ZN(n303) );
  NAND2_X1 U158 ( .A1(\mem[7][1] ), .A2(n401), .ZN(n399) );
  OAI21_X1 U159 ( .B1(n290), .B2(n401), .A(n398), .ZN(n302) );
  NAND2_X1 U160 ( .A1(\mem[7][2] ), .A2(n401), .ZN(n398) );
  OAI21_X1 U161 ( .B1(n289), .B2(n401), .A(n397), .ZN(n301) );
  NAND2_X1 U162 ( .A1(\mem[7][3] ), .A2(n401), .ZN(n397) );
  OAI21_X1 U163 ( .B1(n288), .B2(n401), .A(n396), .ZN(n300) );
  NAND2_X1 U164 ( .A1(\mem[7][4] ), .A2(n401), .ZN(n396) );
  OAI21_X1 U165 ( .B1(n287), .B2(n401), .A(n395), .ZN(n299) );
  NAND2_X1 U166 ( .A1(\mem[7][5] ), .A2(n401), .ZN(n395) );
  OAI21_X1 U167 ( .B1(n286), .B2(n401), .A(n394), .ZN(n298) );
  NAND2_X1 U168 ( .A1(\mem[7][6] ), .A2(n401), .ZN(n394) );
  OAI21_X1 U169 ( .B1(n285), .B2(n401), .A(n393), .ZN(n297) );
  NAND2_X1 U170 ( .A1(\mem[7][7] ), .A2(n401), .ZN(n393) );
  OAI21_X1 U171 ( .B1(n284), .B2(n401), .A(n392), .ZN(n296) );
  NAND2_X1 U172 ( .A1(\mem[7][8] ), .A2(n401), .ZN(n392) );
  OAI21_X1 U173 ( .B1(n283), .B2(n401), .A(n391), .ZN(n295) );
  NAND2_X1 U174 ( .A1(\mem[7][9] ), .A2(n401), .ZN(n391) );
  OAI21_X1 U175 ( .B1(n282), .B2(n401), .A(n390), .ZN(n294) );
  NAND2_X1 U176 ( .A1(\mem[7][10] ), .A2(n401), .ZN(n390) );
  OAI21_X1 U177 ( .B1(n281), .B2(n401), .A(n389), .ZN(n293) );
  NAND2_X1 U178 ( .A1(\mem[7][11] ), .A2(n401), .ZN(n389) );
  OAI21_X1 U179 ( .B1(n494), .B2(n292), .A(n493), .ZN(n388) );
  NAND2_X1 U180 ( .A1(\mem[0][0] ), .A2(n494), .ZN(n493) );
  OAI21_X1 U181 ( .B1(n494), .B2(n291), .A(n492), .ZN(n387) );
  NAND2_X1 U182 ( .A1(\mem[0][1] ), .A2(n494), .ZN(n492) );
  OAI21_X1 U183 ( .B1(n494), .B2(n290), .A(n491), .ZN(n386) );
  NAND2_X1 U184 ( .A1(\mem[0][2] ), .A2(n494), .ZN(n491) );
  OAI21_X1 U185 ( .B1(n494), .B2(n289), .A(n490), .ZN(n385) );
  NAND2_X1 U186 ( .A1(\mem[0][3] ), .A2(n494), .ZN(n490) );
  OAI21_X1 U187 ( .B1(n494), .B2(n288), .A(n489), .ZN(n384) );
  NAND2_X1 U188 ( .A1(\mem[0][4] ), .A2(n494), .ZN(n489) );
  OAI21_X1 U189 ( .B1(n494), .B2(n287), .A(n488), .ZN(n383) );
  NAND2_X1 U190 ( .A1(\mem[0][5] ), .A2(n494), .ZN(n488) );
  OAI21_X1 U191 ( .B1(n494), .B2(n286), .A(n487), .ZN(n382) );
  NAND2_X1 U192 ( .A1(\mem[0][6] ), .A2(n494), .ZN(n487) );
  OAI21_X1 U193 ( .B1(n494), .B2(n285), .A(n486), .ZN(n381) );
  NAND2_X1 U194 ( .A1(\mem[0][7] ), .A2(n494), .ZN(n486) );
  OAI21_X1 U195 ( .B1(n494), .B2(n284), .A(n485), .ZN(n380) );
  NAND2_X1 U196 ( .A1(\mem[0][8] ), .A2(n494), .ZN(n485) );
  OAI21_X1 U197 ( .B1(n494), .B2(n283), .A(n484), .ZN(n379) );
  NAND2_X1 U198 ( .A1(\mem[0][9] ), .A2(n494), .ZN(n484) );
  OAI21_X1 U199 ( .B1(n494), .B2(n282), .A(n483), .ZN(n378) );
  NAND2_X1 U200 ( .A1(\mem[0][10] ), .A2(n494), .ZN(n483) );
  OAI21_X1 U201 ( .B1(n494), .B2(n281), .A(n482), .ZN(n377) );
  NAND2_X1 U202 ( .A1(\mem[0][11] ), .A2(n494), .ZN(n482) );
  INV_X1 U203 ( .A(data_in[0]), .ZN(n292) );
  INV_X1 U204 ( .A(data_in[1]), .ZN(n291) );
  INV_X1 U205 ( .A(data_in[2]), .ZN(n290) );
  INV_X1 U206 ( .A(data_in[3]), .ZN(n289) );
  INV_X1 U207 ( .A(data_in[4]), .ZN(n288) );
  INV_X1 U208 ( .A(data_in[5]), .ZN(n287) );
  INV_X1 U209 ( .A(data_in[6]), .ZN(n286) );
  INV_X1 U210 ( .A(data_in[7]), .ZN(n285) );
  INV_X1 U211 ( .A(data_in[8]), .ZN(n284) );
  INV_X1 U220 ( .A(data_in[9]), .ZN(n283) );
  INV_X1 U221 ( .A(data_in[10]), .ZN(n282) );
  INV_X1 U222 ( .A(data_in[11]), .ZN(n281) );
  MUX2_X1 U223 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n277), .Z(n1) );
  MUX2_X1 U224 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(N10), .Z(n2) );
  MUX2_X1 U225 ( .A(n2), .B(n1), .S(n275), .Z(n3) );
  MUX2_X1 U226 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(N10), .Z(n4) );
  MUX2_X1 U227 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n5) );
  MUX2_X1 U228 ( .A(n5), .B(n4), .S(n275), .Z(n6) );
  MUX2_X1 U229 ( .A(n6), .B(n3), .S(N12), .Z(N24) );
  MUX2_X1 U230 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(N10), .Z(n7) );
  MUX2_X1 U231 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n277), .Z(n8) );
  MUX2_X1 U232 ( .A(n8), .B(n7), .S(n275), .Z(n9) );
  MUX2_X1 U233 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n277), .Z(n10) );
  MUX2_X1 U234 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n277), .Z(n11) );
  MUX2_X1 U235 ( .A(n11), .B(n10), .S(n275), .Z(n12) );
  MUX2_X1 U236 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n277), .Z(n13) );
  MUX2_X1 U237 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n277), .Z(n14) );
  MUX2_X1 U238 ( .A(n14), .B(n13), .S(n275), .Z(n15) );
  MUX2_X1 U239 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n277), .Z(n218) );
  MUX2_X1 U240 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n277), .Z(n219) );
  MUX2_X1 U241 ( .A(n219), .B(n218), .S(n275), .Z(n220) );
  MUX2_X1 U242 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(N10), .Z(n221) );
  MUX2_X1 U243 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n222) );
  MUX2_X1 U244 ( .A(n222), .B(n221), .S(n275), .Z(n223) );
  MUX2_X1 U245 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n277), .Z(n224) );
  MUX2_X1 U246 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n225) );
  MUX2_X1 U247 ( .A(n225), .B(n224), .S(n275), .Z(n226) );
  MUX2_X1 U248 ( .A(n226), .B(n223), .S(N12), .Z(N21) );
  MUX2_X1 U249 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(N10), .Z(n227) );
  MUX2_X1 U250 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(N10), .Z(n228) );
  MUX2_X1 U251 ( .A(n228), .B(n227), .S(n275), .Z(n229) );
  MUX2_X1 U252 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(N10), .Z(n230) );
  MUX2_X1 U253 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n231) );
  MUX2_X1 U254 ( .A(n231), .B(n230), .S(n275), .Z(n232) );
  MUX2_X1 U255 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(N10), .Z(n233) );
  MUX2_X1 U256 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(N10), .Z(n234) );
  MUX2_X1 U257 ( .A(n234), .B(n233), .S(n275), .Z(n235) );
  MUX2_X1 U258 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n236) );
  MUX2_X1 U259 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(N10), .Z(n237) );
  MUX2_X1 U260 ( .A(n237), .B(n236), .S(n275), .Z(n238) );
  MUX2_X1 U261 ( .A(n238), .B(n235), .S(N12), .Z(N19) );
  MUX2_X1 U262 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n276), .Z(n239) );
  MUX2_X1 U263 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n276), .Z(n240) );
  MUX2_X1 U264 ( .A(n240), .B(n239), .S(n275), .Z(n241) );
  MUX2_X1 U265 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n276), .Z(n242) );
  MUX2_X1 U266 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n276), .Z(n243) );
  MUX2_X1 U267 ( .A(n243), .B(n242), .S(n275), .Z(n244) );
  MUX2_X1 U268 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n276), .Z(n245) );
  MUX2_X1 U269 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n276), .Z(n246) );
  MUX2_X1 U270 ( .A(n246), .B(n245), .S(n275), .Z(n247) );
  MUX2_X1 U271 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n276), .Z(n248) );
  MUX2_X1 U272 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n276), .Z(n249) );
  MUX2_X1 U273 ( .A(n249), .B(n248), .S(n275), .Z(n250) );
  MUX2_X1 U274 ( .A(n250), .B(n247), .S(N12), .Z(N17) );
  MUX2_X1 U275 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n276), .Z(n251) );
  MUX2_X1 U276 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n276), .Z(n252) );
  MUX2_X1 U277 ( .A(n252), .B(n251), .S(n275), .Z(n253) );
  MUX2_X1 U278 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n276), .Z(n254) );
  MUX2_X1 U279 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n276), .Z(n255) );
  MUX2_X1 U280 ( .A(n255), .B(n254), .S(n275), .Z(n256) );
  MUX2_X1 U281 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n277), .Z(n257) );
  MUX2_X1 U282 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n277), .Z(n258) );
  MUX2_X1 U283 ( .A(n258), .B(n257), .S(n275), .Z(n259) );
  MUX2_X1 U284 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n277), .Z(n260) );
  MUX2_X1 U285 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n277), .Z(n261) );
  MUX2_X1 U286 ( .A(n261), .B(n260), .S(N11), .Z(n262) );
  MUX2_X1 U287 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n277), .Z(n263) );
  MUX2_X1 U288 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n277), .Z(n264) );
  MUX2_X1 U289 ( .A(n264), .B(n263), .S(n275), .Z(n265) );
  MUX2_X1 U290 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n277), .Z(n266) );
  MUX2_X1 U291 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n277), .Z(n267) );
  MUX2_X1 U292 ( .A(n267), .B(n266), .S(N11), .Z(n268) );
  MUX2_X1 U293 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n277), .Z(n269) );
  MUX2_X1 U294 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n277), .Z(n270) );
  MUX2_X1 U295 ( .A(n270), .B(n269), .S(n275), .Z(n271) );
  MUX2_X1 U296 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n277), .Z(n272) );
  MUX2_X1 U297 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n277), .Z(n273) );
  MUX2_X1 U298 ( .A(n273), .B(n272), .S(n275), .Z(n274) );
  MUX2_X1 U299 ( .A(n274), .B(n271), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH12_SIZE8_LOGSIZE3_2 ( clk, data_in, data_out, addr, wr_en
 );
  input [11:0] data_in;
  output [11:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] ,
         \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] ,
         \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][11] , \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] ,
         \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] ,
         \mem[5][1] , \mem[5][0] , \mem[4][11] , \mem[4][10] , \mem[4][9] ,
         \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] ,
         \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] ,
         \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] ,
         \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][11] , \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] ,
         \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] ,
         \mem[0][1] , \mem[0][0] , N13, N14, n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[11]  ( .D(N13), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N14), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \mem_reg[7][11]  ( .D(n293), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n294), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n295), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n296), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n297), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n298), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n299), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n300), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n301), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n302), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n303), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n304), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n305), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n306), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n307), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n308), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n309), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n310), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n311), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n312), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n313), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n314), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n315), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n316), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n317), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n318), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n319), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n320), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n321), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n322), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n323), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n324), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n325), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n326), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n327), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n328), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n329), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n330), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n331), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n332), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n333), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n334), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n335), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n336), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n337), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n338), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n339), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n340), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n341), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n342), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n343), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n344), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n345), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n346), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n347), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n348), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n349), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n350), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n351), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n352), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n353), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n354), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n355), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n356), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n357), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n358), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n359), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n360), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n361), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n362), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n363), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n364), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n365), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n366), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n367), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n368), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n369), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n370), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n371), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n372), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n373), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n374), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n375), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n376), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n377), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n378), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n379), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n380), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n381), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n382), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n383), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n384), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n385), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n386), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n387), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n388), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U212 ( .A1(n278), .A2(n279), .A3(n481), .ZN(n494) );
  NAND3_X1 U213 ( .A1(n481), .A2(n279), .A3(N10), .ZN(n480) );
  NAND3_X1 U214 ( .A1(n481), .A2(n278), .A3(N11), .ZN(n467) );
  NAND3_X1 U215 ( .A1(N10), .A2(n481), .A3(N11), .ZN(n454) );
  NAND3_X1 U216 ( .A1(n278), .A2(n279), .A3(n428), .ZN(n441) );
  NAND3_X1 U217 ( .A1(N10), .A2(n279), .A3(n428), .ZN(n427) );
  NAND3_X1 U218 ( .A1(N11), .A2(n278), .A3(n428), .ZN(n414) );
  NAND3_X1 U219 ( .A1(N11), .A2(N10), .A3(n428), .ZN(n401) );
  SDFF_X1 \data_out_reg[7]  ( .D(n250), .SI(n247), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n238), .SI(n235), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[6]  ( .D(n244), .SI(n241), .SE(N12), .CK(clk), .Q(
        data_out[6]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n262), .SI(n259), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[4]  ( .D(n232), .SI(n229), .SE(N12), .CK(clk), .Q(
        data_out[4]) );
  SDFF_X1 \data_out_reg[2]  ( .D(n220), .SI(n15), .SE(N12), .CK(clk), .Q(
        data_out[2]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n6), .SI(n3), .SE(N12), .CK(clk), .Q(
        data_out[0]) );
  SDFF_X1 \data_out_reg[8]  ( .D(n256), .SI(n253), .SE(N12), .CK(clk), .Q(
        data_out[8]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n12), .SI(n9), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n226), .SI(n223), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  BUF_X1 U3 ( .A(N10), .Z(n276) );
  BUF_X1 U4 ( .A(N11), .Z(n275) );
  BUF_X1 U5 ( .A(N10), .Z(n277) );
  AND2_X1 U6 ( .A1(N12), .A2(wr_en), .ZN(n428) );
  INV_X1 U7 ( .A(N10), .ZN(n278) );
  INV_X1 U8 ( .A(N11), .ZN(n279) );
  OAI21_X1 U9 ( .B1(n292), .B2(n480), .A(n479), .ZN(n376) );
  NAND2_X1 U10 ( .A1(\mem[1][0] ), .A2(n480), .ZN(n479) );
  OAI21_X1 U11 ( .B1(n291), .B2(n480), .A(n478), .ZN(n375) );
  NAND2_X1 U12 ( .A1(\mem[1][1] ), .A2(n480), .ZN(n478) );
  OAI21_X1 U13 ( .B1(n290), .B2(n480), .A(n477), .ZN(n374) );
  NAND2_X1 U14 ( .A1(\mem[1][2] ), .A2(n480), .ZN(n477) );
  OAI21_X1 U15 ( .B1(n289), .B2(n480), .A(n476), .ZN(n373) );
  NAND2_X1 U16 ( .A1(\mem[1][3] ), .A2(n480), .ZN(n476) );
  OAI21_X1 U17 ( .B1(n288), .B2(n480), .A(n475), .ZN(n372) );
  NAND2_X1 U18 ( .A1(\mem[1][4] ), .A2(n480), .ZN(n475) );
  OAI21_X1 U19 ( .B1(n287), .B2(n480), .A(n474), .ZN(n371) );
  NAND2_X1 U20 ( .A1(\mem[1][5] ), .A2(n480), .ZN(n474) );
  OAI21_X1 U21 ( .B1(n286), .B2(n480), .A(n473), .ZN(n370) );
  NAND2_X1 U22 ( .A1(\mem[1][6] ), .A2(n480), .ZN(n473) );
  OAI21_X1 U23 ( .B1(n285), .B2(n480), .A(n472), .ZN(n369) );
  NAND2_X1 U24 ( .A1(\mem[1][7] ), .A2(n480), .ZN(n472) );
  OAI21_X1 U25 ( .B1(n284), .B2(n480), .A(n471), .ZN(n368) );
  NAND2_X1 U26 ( .A1(\mem[1][8] ), .A2(n480), .ZN(n471) );
  OAI21_X1 U27 ( .B1(n283), .B2(n480), .A(n470), .ZN(n367) );
  NAND2_X1 U28 ( .A1(\mem[1][9] ), .A2(n480), .ZN(n470) );
  OAI21_X1 U29 ( .B1(n282), .B2(n480), .A(n469), .ZN(n366) );
  NAND2_X1 U30 ( .A1(\mem[1][10] ), .A2(n480), .ZN(n469) );
  OAI21_X1 U31 ( .B1(n281), .B2(n480), .A(n468), .ZN(n365) );
  NAND2_X1 U32 ( .A1(\mem[1][11] ), .A2(n480), .ZN(n468) );
  OAI21_X1 U33 ( .B1(n292), .B2(n467), .A(n466), .ZN(n364) );
  NAND2_X1 U34 ( .A1(\mem[2][0] ), .A2(n467), .ZN(n466) );
  OAI21_X1 U35 ( .B1(n291), .B2(n467), .A(n465), .ZN(n363) );
  NAND2_X1 U36 ( .A1(\mem[2][1] ), .A2(n467), .ZN(n465) );
  OAI21_X1 U37 ( .B1(n290), .B2(n467), .A(n464), .ZN(n362) );
  NAND2_X1 U38 ( .A1(\mem[2][2] ), .A2(n467), .ZN(n464) );
  OAI21_X1 U39 ( .B1(n289), .B2(n467), .A(n463), .ZN(n361) );
  NAND2_X1 U40 ( .A1(\mem[2][3] ), .A2(n467), .ZN(n463) );
  OAI21_X1 U41 ( .B1(n288), .B2(n467), .A(n462), .ZN(n360) );
  NAND2_X1 U42 ( .A1(\mem[2][4] ), .A2(n467), .ZN(n462) );
  OAI21_X1 U43 ( .B1(n287), .B2(n467), .A(n461), .ZN(n359) );
  NAND2_X1 U44 ( .A1(\mem[2][5] ), .A2(n467), .ZN(n461) );
  OAI21_X1 U45 ( .B1(n286), .B2(n467), .A(n460), .ZN(n358) );
  NAND2_X1 U46 ( .A1(\mem[2][6] ), .A2(n467), .ZN(n460) );
  OAI21_X1 U47 ( .B1(n285), .B2(n467), .A(n459), .ZN(n357) );
  NAND2_X1 U48 ( .A1(\mem[2][7] ), .A2(n467), .ZN(n459) );
  OAI21_X1 U49 ( .B1(n284), .B2(n467), .A(n458), .ZN(n356) );
  NAND2_X1 U50 ( .A1(\mem[2][8] ), .A2(n467), .ZN(n458) );
  OAI21_X1 U51 ( .B1(n283), .B2(n467), .A(n457), .ZN(n355) );
  NAND2_X1 U52 ( .A1(\mem[2][9] ), .A2(n467), .ZN(n457) );
  OAI21_X1 U53 ( .B1(n282), .B2(n467), .A(n456), .ZN(n354) );
  NAND2_X1 U54 ( .A1(\mem[2][10] ), .A2(n467), .ZN(n456) );
  OAI21_X1 U55 ( .B1(n281), .B2(n467), .A(n455), .ZN(n353) );
  NAND2_X1 U56 ( .A1(\mem[2][11] ), .A2(n467), .ZN(n455) );
  OAI21_X1 U57 ( .B1(n292), .B2(n454), .A(n453), .ZN(n352) );
  NAND2_X1 U58 ( .A1(\mem[3][0] ), .A2(n454), .ZN(n453) );
  OAI21_X1 U59 ( .B1(n291), .B2(n454), .A(n452), .ZN(n351) );
  NAND2_X1 U60 ( .A1(\mem[3][1] ), .A2(n454), .ZN(n452) );
  OAI21_X1 U61 ( .B1(n290), .B2(n454), .A(n451), .ZN(n350) );
  NAND2_X1 U62 ( .A1(\mem[3][2] ), .A2(n454), .ZN(n451) );
  OAI21_X1 U63 ( .B1(n289), .B2(n454), .A(n450), .ZN(n349) );
  NAND2_X1 U64 ( .A1(\mem[3][3] ), .A2(n454), .ZN(n450) );
  OAI21_X1 U65 ( .B1(n288), .B2(n454), .A(n449), .ZN(n348) );
  NAND2_X1 U66 ( .A1(\mem[3][4] ), .A2(n454), .ZN(n449) );
  OAI21_X1 U67 ( .B1(n287), .B2(n454), .A(n448), .ZN(n347) );
  NAND2_X1 U68 ( .A1(\mem[3][5] ), .A2(n454), .ZN(n448) );
  OAI21_X1 U69 ( .B1(n286), .B2(n454), .A(n447), .ZN(n346) );
  NAND2_X1 U70 ( .A1(\mem[3][6] ), .A2(n454), .ZN(n447) );
  OAI21_X1 U71 ( .B1(n285), .B2(n454), .A(n446), .ZN(n345) );
  NAND2_X1 U72 ( .A1(\mem[3][7] ), .A2(n454), .ZN(n446) );
  OAI21_X1 U73 ( .B1(n284), .B2(n454), .A(n445), .ZN(n344) );
  NAND2_X1 U74 ( .A1(\mem[3][8] ), .A2(n454), .ZN(n445) );
  OAI21_X1 U75 ( .B1(n283), .B2(n454), .A(n444), .ZN(n343) );
  NAND2_X1 U76 ( .A1(\mem[3][9] ), .A2(n454), .ZN(n444) );
  OAI21_X1 U77 ( .B1(n282), .B2(n454), .A(n443), .ZN(n342) );
  NAND2_X1 U78 ( .A1(\mem[3][10] ), .A2(n454), .ZN(n443) );
  OAI21_X1 U79 ( .B1(n281), .B2(n454), .A(n442), .ZN(n341) );
  NAND2_X1 U80 ( .A1(\mem[3][11] ), .A2(n454), .ZN(n442) );
  OAI21_X1 U81 ( .B1(n292), .B2(n441), .A(n440), .ZN(n340) );
  NAND2_X1 U82 ( .A1(\mem[4][0] ), .A2(n441), .ZN(n440) );
  OAI21_X1 U83 ( .B1(n291), .B2(n441), .A(n439), .ZN(n339) );
  NAND2_X1 U84 ( .A1(\mem[4][1] ), .A2(n441), .ZN(n439) );
  OAI21_X1 U85 ( .B1(n290), .B2(n441), .A(n438), .ZN(n338) );
  NAND2_X1 U86 ( .A1(\mem[4][2] ), .A2(n441), .ZN(n438) );
  OAI21_X1 U87 ( .B1(n289), .B2(n441), .A(n437), .ZN(n337) );
  NAND2_X1 U88 ( .A1(\mem[4][3] ), .A2(n441), .ZN(n437) );
  OAI21_X1 U89 ( .B1(n288), .B2(n441), .A(n436), .ZN(n336) );
  NAND2_X1 U90 ( .A1(\mem[4][4] ), .A2(n441), .ZN(n436) );
  OAI21_X1 U91 ( .B1(n287), .B2(n441), .A(n435), .ZN(n335) );
  NAND2_X1 U92 ( .A1(\mem[4][5] ), .A2(n441), .ZN(n435) );
  OAI21_X1 U93 ( .B1(n286), .B2(n441), .A(n434), .ZN(n334) );
  NAND2_X1 U94 ( .A1(\mem[4][6] ), .A2(n441), .ZN(n434) );
  OAI21_X1 U95 ( .B1(n285), .B2(n441), .A(n433), .ZN(n333) );
  NAND2_X1 U96 ( .A1(\mem[4][7] ), .A2(n441), .ZN(n433) );
  OAI21_X1 U97 ( .B1(n284), .B2(n441), .A(n432), .ZN(n332) );
  NAND2_X1 U98 ( .A1(\mem[4][8] ), .A2(n441), .ZN(n432) );
  OAI21_X1 U99 ( .B1(n283), .B2(n441), .A(n431), .ZN(n331) );
  NAND2_X1 U100 ( .A1(\mem[4][9] ), .A2(n441), .ZN(n431) );
  OAI21_X1 U101 ( .B1(n282), .B2(n441), .A(n430), .ZN(n330) );
  NAND2_X1 U102 ( .A1(\mem[4][10] ), .A2(n441), .ZN(n430) );
  OAI21_X1 U103 ( .B1(n281), .B2(n441), .A(n429), .ZN(n329) );
  NAND2_X1 U104 ( .A1(\mem[4][11] ), .A2(n441), .ZN(n429) );
  OAI21_X1 U105 ( .B1(n292), .B2(n427), .A(n426), .ZN(n328) );
  NAND2_X1 U106 ( .A1(\mem[5][0] ), .A2(n427), .ZN(n426) );
  OAI21_X1 U107 ( .B1(n291), .B2(n427), .A(n425), .ZN(n327) );
  NAND2_X1 U108 ( .A1(\mem[5][1] ), .A2(n427), .ZN(n425) );
  OAI21_X1 U109 ( .B1(n290), .B2(n427), .A(n424), .ZN(n326) );
  NAND2_X1 U110 ( .A1(\mem[5][2] ), .A2(n427), .ZN(n424) );
  OAI21_X1 U111 ( .B1(n289), .B2(n427), .A(n423), .ZN(n325) );
  NAND2_X1 U112 ( .A1(\mem[5][3] ), .A2(n427), .ZN(n423) );
  OAI21_X1 U113 ( .B1(n288), .B2(n427), .A(n422), .ZN(n324) );
  NAND2_X1 U114 ( .A1(\mem[5][4] ), .A2(n427), .ZN(n422) );
  OAI21_X1 U115 ( .B1(n287), .B2(n427), .A(n421), .ZN(n323) );
  NAND2_X1 U116 ( .A1(\mem[5][5] ), .A2(n427), .ZN(n421) );
  OAI21_X1 U117 ( .B1(n286), .B2(n427), .A(n420), .ZN(n322) );
  NAND2_X1 U118 ( .A1(\mem[5][6] ), .A2(n427), .ZN(n420) );
  OAI21_X1 U119 ( .B1(n285), .B2(n427), .A(n419), .ZN(n321) );
  NAND2_X1 U120 ( .A1(\mem[5][7] ), .A2(n427), .ZN(n419) );
  OAI21_X1 U121 ( .B1(n284), .B2(n427), .A(n418), .ZN(n320) );
  NAND2_X1 U122 ( .A1(\mem[5][8] ), .A2(n427), .ZN(n418) );
  OAI21_X1 U123 ( .B1(n283), .B2(n427), .A(n417), .ZN(n319) );
  NAND2_X1 U124 ( .A1(\mem[5][9] ), .A2(n427), .ZN(n417) );
  OAI21_X1 U125 ( .B1(n282), .B2(n427), .A(n416), .ZN(n318) );
  NAND2_X1 U126 ( .A1(\mem[5][10] ), .A2(n427), .ZN(n416) );
  OAI21_X1 U127 ( .B1(n281), .B2(n427), .A(n415), .ZN(n317) );
  NAND2_X1 U128 ( .A1(\mem[5][11] ), .A2(n427), .ZN(n415) );
  OAI21_X1 U129 ( .B1(n292), .B2(n414), .A(n413), .ZN(n316) );
  NAND2_X1 U130 ( .A1(\mem[6][0] ), .A2(n414), .ZN(n413) );
  OAI21_X1 U131 ( .B1(n291), .B2(n414), .A(n412), .ZN(n315) );
  NAND2_X1 U132 ( .A1(\mem[6][1] ), .A2(n414), .ZN(n412) );
  OAI21_X1 U133 ( .B1(n290), .B2(n414), .A(n411), .ZN(n314) );
  NAND2_X1 U134 ( .A1(\mem[6][2] ), .A2(n414), .ZN(n411) );
  OAI21_X1 U135 ( .B1(n289), .B2(n414), .A(n410), .ZN(n313) );
  NAND2_X1 U136 ( .A1(\mem[6][3] ), .A2(n414), .ZN(n410) );
  OAI21_X1 U137 ( .B1(n288), .B2(n414), .A(n409), .ZN(n312) );
  NAND2_X1 U138 ( .A1(\mem[6][4] ), .A2(n414), .ZN(n409) );
  OAI21_X1 U139 ( .B1(n287), .B2(n414), .A(n408), .ZN(n311) );
  NAND2_X1 U140 ( .A1(\mem[6][5] ), .A2(n414), .ZN(n408) );
  OAI21_X1 U141 ( .B1(n286), .B2(n414), .A(n407), .ZN(n310) );
  NAND2_X1 U142 ( .A1(\mem[6][6] ), .A2(n414), .ZN(n407) );
  OAI21_X1 U143 ( .B1(n285), .B2(n414), .A(n406), .ZN(n309) );
  NAND2_X1 U144 ( .A1(\mem[6][7] ), .A2(n414), .ZN(n406) );
  OAI21_X1 U145 ( .B1(n284), .B2(n414), .A(n405), .ZN(n308) );
  NAND2_X1 U146 ( .A1(\mem[6][8] ), .A2(n414), .ZN(n405) );
  OAI21_X1 U147 ( .B1(n283), .B2(n414), .A(n404), .ZN(n307) );
  NAND2_X1 U148 ( .A1(\mem[6][9] ), .A2(n414), .ZN(n404) );
  OAI21_X1 U149 ( .B1(n282), .B2(n414), .A(n403), .ZN(n306) );
  NAND2_X1 U150 ( .A1(\mem[6][10] ), .A2(n414), .ZN(n403) );
  OAI21_X1 U151 ( .B1(n281), .B2(n414), .A(n402), .ZN(n305) );
  NAND2_X1 U152 ( .A1(\mem[6][11] ), .A2(n414), .ZN(n402) );
  OAI21_X1 U153 ( .B1(n292), .B2(n401), .A(n400), .ZN(n304) );
  NAND2_X1 U154 ( .A1(\mem[7][0] ), .A2(n401), .ZN(n400) );
  OAI21_X1 U155 ( .B1(n291), .B2(n401), .A(n399), .ZN(n303) );
  NAND2_X1 U156 ( .A1(\mem[7][1] ), .A2(n401), .ZN(n399) );
  OAI21_X1 U157 ( .B1(n290), .B2(n401), .A(n398), .ZN(n302) );
  NAND2_X1 U158 ( .A1(\mem[7][2] ), .A2(n401), .ZN(n398) );
  OAI21_X1 U159 ( .B1(n289), .B2(n401), .A(n397), .ZN(n301) );
  NAND2_X1 U160 ( .A1(\mem[7][3] ), .A2(n401), .ZN(n397) );
  OAI21_X1 U161 ( .B1(n288), .B2(n401), .A(n396), .ZN(n300) );
  NAND2_X1 U162 ( .A1(\mem[7][4] ), .A2(n401), .ZN(n396) );
  OAI21_X1 U163 ( .B1(n287), .B2(n401), .A(n395), .ZN(n299) );
  NAND2_X1 U164 ( .A1(\mem[7][5] ), .A2(n401), .ZN(n395) );
  OAI21_X1 U165 ( .B1(n286), .B2(n401), .A(n394), .ZN(n298) );
  NAND2_X1 U166 ( .A1(\mem[7][6] ), .A2(n401), .ZN(n394) );
  OAI21_X1 U167 ( .B1(n285), .B2(n401), .A(n393), .ZN(n297) );
  NAND2_X1 U168 ( .A1(\mem[7][7] ), .A2(n401), .ZN(n393) );
  OAI21_X1 U169 ( .B1(n284), .B2(n401), .A(n392), .ZN(n296) );
  NAND2_X1 U170 ( .A1(\mem[7][8] ), .A2(n401), .ZN(n392) );
  OAI21_X1 U171 ( .B1(n283), .B2(n401), .A(n391), .ZN(n295) );
  NAND2_X1 U172 ( .A1(\mem[7][9] ), .A2(n401), .ZN(n391) );
  OAI21_X1 U173 ( .B1(n282), .B2(n401), .A(n390), .ZN(n294) );
  NAND2_X1 U174 ( .A1(\mem[7][10] ), .A2(n401), .ZN(n390) );
  OAI21_X1 U175 ( .B1(n281), .B2(n401), .A(n389), .ZN(n293) );
  NAND2_X1 U176 ( .A1(\mem[7][11] ), .A2(n401), .ZN(n389) );
  OAI21_X1 U177 ( .B1(n494), .B2(n292), .A(n493), .ZN(n388) );
  NAND2_X1 U178 ( .A1(\mem[0][0] ), .A2(n494), .ZN(n493) );
  OAI21_X1 U179 ( .B1(n494), .B2(n291), .A(n492), .ZN(n387) );
  NAND2_X1 U180 ( .A1(\mem[0][1] ), .A2(n494), .ZN(n492) );
  OAI21_X1 U181 ( .B1(n494), .B2(n290), .A(n491), .ZN(n386) );
  NAND2_X1 U182 ( .A1(\mem[0][2] ), .A2(n494), .ZN(n491) );
  OAI21_X1 U183 ( .B1(n494), .B2(n289), .A(n490), .ZN(n385) );
  NAND2_X1 U184 ( .A1(\mem[0][3] ), .A2(n494), .ZN(n490) );
  OAI21_X1 U185 ( .B1(n494), .B2(n288), .A(n489), .ZN(n384) );
  NAND2_X1 U186 ( .A1(\mem[0][4] ), .A2(n494), .ZN(n489) );
  OAI21_X1 U187 ( .B1(n494), .B2(n287), .A(n488), .ZN(n383) );
  NAND2_X1 U188 ( .A1(\mem[0][5] ), .A2(n494), .ZN(n488) );
  OAI21_X1 U189 ( .B1(n494), .B2(n286), .A(n487), .ZN(n382) );
  NAND2_X1 U190 ( .A1(\mem[0][6] ), .A2(n494), .ZN(n487) );
  OAI21_X1 U191 ( .B1(n494), .B2(n285), .A(n486), .ZN(n381) );
  NAND2_X1 U192 ( .A1(\mem[0][7] ), .A2(n494), .ZN(n486) );
  OAI21_X1 U193 ( .B1(n494), .B2(n284), .A(n485), .ZN(n380) );
  NAND2_X1 U194 ( .A1(\mem[0][8] ), .A2(n494), .ZN(n485) );
  OAI21_X1 U195 ( .B1(n494), .B2(n283), .A(n484), .ZN(n379) );
  NAND2_X1 U196 ( .A1(\mem[0][9] ), .A2(n494), .ZN(n484) );
  OAI21_X1 U197 ( .B1(n494), .B2(n282), .A(n483), .ZN(n378) );
  NAND2_X1 U198 ( .A1(\mem[0][10] ), .A2(n494), .ZN(n483) );
  OAI21_X1 U199 ( .B1(n494), .B2(n281), .A(n482), .ZN(n377) );
  NAND2_X1 U200 ( .A1(\mem[0][11] ), .A2(n494), .ZN(n482) );
  NOR2_X1 U201 ( .A1(n280), .A2(N12), .ZN(n481) );
  INV_X1 U202 ( .A(wr_en), .ZN(n280) );
  INV_X1 U203 ( .A(data_in[0]), .ZN(n292) );
  INV_X1 U204 ( .A(data_in[1]), .ZN(n291) );
  INV_X1 U205 ( .A(data_in[2]), .ZN(n290) );
  INV_X1 U206 ( .A(data_in[3]), .ZN(n289) );
  INV_X1 U207 ( .A(data_in[4]), .ZN(n288) );
  INV_X1 U208 ( .A(data_in[5]), .ZN(n287) );
  INV_X1 U209 ( .A(data_in[6]), .ZN(n286) );
  INV_X1 U210 ( .A(data_in[7]), .ZN(n285) );
  INV_X1 U211 ( .A(data_in[8]), .ZN(n284) );
  INV_X1 U220 ( .A(data_in[9]), .ZN(n283) );
  INV_X1 U221 ( .A(data_in[10]), .ZN(n282) );
  INV_X1 U222 ( .A(data_in[11]), .ZN(n281) );
  MUX2_X1 U223 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n277), .Z(n1) );
  MUX2_X1 U224 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n277), .Z(n2) );
  MUX2_X1 U225 ( .A(n2), .B(n1), .S(n275), .Z(n3) );
  MUX2_X1 U226 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n277), .Z(n4) );
  MUX2_X1 U227 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n277), .Z(n5) );
  MUX2_X1 U228 ( .A(n5), .B(n4), .S(n275), .Z(n6) );
  MUX2_X1 U229 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n277), .Z(n7) );
  MUX2_X1 U230 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n277), .Z(n8) );
  MUX2_X1 U231 ( .A(n8), .B(n7), .S(n275), .Z(n9) );
  MUX2_X1 U232 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n277), .Z(n10) );
  MUX2_X1 U233 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n277), .Z(n11) );
  MUX2_X1 U234 ( .A(n11), .B(n10), .S(n275), .Z(n12) );
  MUX2_X1 U235 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n277), .Z(n13) );
  MUX2_X1 U236 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n277), .Z(n14) );
  MUX2_X1 U237 ( .A(n14), .B(n13), .S(n275), .Z(n15) );
  MUX2_X1 U238 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n277), .Z(n218) );
  MUX2_X1 U239 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n277), .Z(n219) );
  MUX2_X1 U240 ( .A(n219), .B(n218), .S(n275), .Z(n220) );
  MUX2_X1 U241 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n276), .Z(n221) );
  MUX2_X1 U242 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n276), .Z(n222) );
  MUX2_X1 U243 ( .A(n222), .B(n221), .S(n275), .Z(n223) );
  MUX2_X1 U244 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n276), .Z(n224) );
  MUX2_X1 U245 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n225) );
  MUX2_X1 U246 ( .A(n225), .B(n224), .S(n275), .Z(n226) );
  MUX2_X1 U247 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n276), .Z(n227) );
  MUX2_X1 U248 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n276), .Z(n228) );
  MUX2_X1 U249 ( .A(n228), .B(n227), .S(n275), .Z(n229) );
  MUX2_X1 U250 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(N10), .Z(n230) );
  MUX2_X1 U251 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n231) );
  MUX2_X1 U252 ( .A(n231), .B(n230), .S(n275), .Z(n232) );
  MUX2_X1 U253 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n276), .Z(n233) );
  MUX2_X1 U254 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n277), .Z(n234) );
  MUX2_X1 U255 ( .A(n234), .B(n233), .S(n275), .Z(n235) );
  MUX2_X1 U256 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n236) );
  MUX2_X1 U257 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(N10), .Z(n237) );
  MUX2_X1 U258 ( .A(n237), .B(n236), .S(n275), .Z(n238) );
  MUX2_X1 U259 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n277), .Z(n239) );
  MUX2_X1 U260 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n277), .Z(n240) );
  MUX2_X1 U261 ( .A(n240), .B(n239), .S(n275), .Z(n241) );
  MUX2_X1 U262 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n242) );
  MUX2_X1 U263 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n243) );
  MUX2_X1 U264 ( .A(n243), .B(n242), .S(n275), .Z(n244) );
  MUX2_X1 U265 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n277), .Z(n245) );
  MUX2_X1 U266 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n246) );
  MUX2_X1 U267 ( .A(n246), .B(n245), .S(n275), .Z(n247) );
  MUX2_X1 U268 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n248) );
  MUX2_X1 U269 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n249) );
  MUX2_X1 U270 ( .A(n249), .B(n248), .S(n275), .Z(n250) );
  MUX2_X1 U271 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n277), .Z(n251) );
  MUX2_X1 U272 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(N10), .Z(n252) );
  MUX2_X1 U273 ( .A(n252), .B(n251), .S(n275), .Z(n253) );
  MUX2_X1 U274 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(N10), .Z(n254) );
  MUX2_X1 U275 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(N10), .Z(n255) );
  MUX2_X1 U276 ( .A(n255), .B(n254), .S(N11), .Z(n256) );
  MUX2_X1 U277 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n276), .Z(n257) );
  MUX2_X1 U278 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n276), .Z(n258) );
  MUX2_X1 U279 ( .A(n258), .B(n257), .S(n275), .Z(n259) );
  MUX2_X1 U280 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n276), .Z(n260) );
  MUX2_X1 U281 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n276), .Z(n261) );
  MUX2_X1 U282 ( .A(n261), .B(n260), .S(N11), .Z(n262) );
  MUX2_X1 U283 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n276), .Z(n263) );
  MUX2_X1 U284 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n276), .Z(n264) );
  MUX2_X1 U285 ( .A(n264), .B(n263), .S(n275), .Z(n265) );
  MUX2_X1 U286 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n276), .Z(n266) );
  MUX2_X1 U287 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n276), .Z(n267) );
  MUX2_X1 U288 ( .A(n267), .B(n266), .S(n275), .Z(n268) );
  MUX2_X1 U289 ( .A(n268), .B(n265), .S(N12), .Z(N14) );
  MUX2_X1 U290 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n276), .Z(n269) );
  MUX2_X1 U291 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n276), .Z(n270) );
  MUX2_X1 U292 ( .A(n270), .B(n269), .S(n275), .Z(n271) );
  MUX2_X1 U293 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n276), .Z(n272) );
  MUX2_X1 U294 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n276), .Z(n273) );
  MUX2_X1 U295 ( .A(n273), .B(n272), .S(n275), .Z(n274) );
  MUX2_X1 U296 ( .A(n274), .B(n271), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH12_SIZE8_LOGSIZE3_1 ( clk, data_in, data_out, addr, wr_en
 );
  input [11:0] data_in;
  output [11:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] ,
         \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] ,
         \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][11] , \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] ,
         \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] ,
         \mem[5][1] , \mem[5][0] , \mem[4][11] , \mem[4][10] , \mem[4][9] ,
         \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] ,
         \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] ,
         \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] ,
         \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][11] , \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] ,
         \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] ,
         \mem[0][1] , \mem[0][0] , N20, N23, N24, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[4]  ( .D(N20), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[1]  ( .D(N23), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N24), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][11]  ( .D(n293), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n294), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n295), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n296), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n297), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n298), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n299), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n300), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n301), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n302), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n303), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n304), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n305), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n306), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n307), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n308), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n309), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n310), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n311), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n312), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n313), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n314), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n315), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n316), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n317), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n318), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n319), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n320), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n321), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n322), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n323), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n324), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n325), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n326), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n327), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n328), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n329), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n330), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n331), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n332), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n333), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n334), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n335), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n336), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n337), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n338), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n339), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n340), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n341), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n342), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n343), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n344), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n345), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n346), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n347), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n348), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n349), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n350), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n351), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n352), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n353), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n354), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n355), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n356), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n357), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n358), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n359), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n360), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n361), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n362), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n363), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n364), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n365), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n366), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n367), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n368), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n369), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n370), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n371), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n372), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n373), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n374), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n375), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n376), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n377), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n378), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n379), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n380), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n381), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n382), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n383), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n384), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n385), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n386), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n387), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n388), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U212 ( .A1(n278), .A2(n279), .A3(n481), .ZN(n494) );
  NAND3_X1 U213 ( .A1(n481), .A2(n279), .A3(N10), .ZN(n480) );
  NAND3_X1 U214 ( .A1(n481), .A2(n278), .A3(N11), .ZN(n467) );
  NAND3_X1 U215 ( .A1(N10), .A2(n481), .A3(N11), .ZN(n454) );
  NAND3_X1 U216 ( .A1(n278), .A2(n279), .A3(n428), .ZN(n441) );
  NAND3_X1 U217 ( .A1(N10), .A2(n279), .A3(n428), .ZN(n427) );
  NAND3_X1 U218 ( .A1(N11), .A2(n278), .A3(n428), .ZN(n414) );
  NAND3_X1 U219 ( .A1(N11), .A2(N10), .A3(n428), .ZN(n401) );
  SDFF_X1 \data_out_reg[3]  ( .D(n226), .SI(n223), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n238), .SI(n235), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[10]  ( .D(n268), .SI(n265), .SE(N12), .CK(clk), .Q(
        data_out[10]) );
  SDFF_X1 \data_out_reg[8]  ( .D(n256), .SI(n253), .SE(N12), .CK(clk), .Q(
        data_out[8]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n250), .SI(n247), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[2]  ( .D(n220), .SI(n15), .SE(N12), .CK(clk), .Q(
        data_out[2]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n262), .SI(n259), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[6]  ( .D(n244), .SI(n241), .SE(N12), .CK(clk), .Q(
        data_out[6]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n274), .SI(n271), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  BUF_X1 U3 ( .A(N10), .Z(n276) );
  BUF_X1 U4 ( .A(N11), .Z(n275) );
  BUF_X1 U5 ( .A(N10), .Z(n277) );
  NOR2_X1 U6 ( .A1(n280), .A2(N12), .ZN(n481) );
  INV_X1 U7 ( .A(wr_en), .ZN(n280) );
  AND2_X1 U8 ( .A1(N12), .A2(wr_en), .ZN(n428) );
  INV_X1 U9 ( .A(N10), .ZN(n278) );
  INV_X1 U10 ( .A(N11), .ZN(n279) );
  OAI21_X1 U11 ( .B1(n292), .B2(n480), .A(n479), .ZN(n376) );
  NAND2_X1 U12 ( .A1(\mem[1][0] ), .A2(n480), .ZN(n479) );
  OAI21_X1 U13 ( .B1(n291), .B2(n480), .A(n478), .ZN(n375) );
  NAND2_X1 U14 ( .A1(\mem[1][1] ), .A2(n480), .ZN(n478) );
  OAI21_X1 U15 ( .B1(n290), .B2(n480), .A(n477), .ZN(n374) );
  NAND2_X1 U16 ( .A1(\mem[1][2] ), .A2(n480), .ZN(n477) );
  OAI21_X1 U17 ( .B1(n289), .B2(n480), .A(n476), .ZN(n373) );
  NAND2_X1 U18 ( .A1(\mem[1][3] ), .A2(n480), .ZN(n476) );
  OAI21_X1 U19 ( .B1(n288), .B2(n480), .A(n475), .ZN(n372) );
  NAND2_X1 U20 ( .A1(\mem[1][4] ), .A2(n480), .ZN(n475) );
  OAI21_X1 U21 ( .B1(n287), .B2(n480), .A(n474), .ZN(n371) );
  NAND2_X1 U22 ( .A1(\mem[1][5] ), .A2(n480), .ZN(n474) );
  OAI21_X1 U23 ( .B1(n286), .B2(n480), .A(n473), .ZN(n370) );
  NAND2_X1 U24 ( .A1(\mem[1][6] ), .A2(n480), .ZN(n473) );
  OAI21_X1 U25 ( .B1(n285), .B2(n480), .A(n472), .ZN(n369) );
  NAND2_X1 U26 ( .A1(\mem[1][7] ), .A2(n480), .ZN(n472) );
  OAI21_X1 U27 ( .B1(n284), .B2(n480), .A(n471), .ZN(n368) );
  NAND2_X1 U28 ( .A1(\mem[1][8] ), .A2(n480), .ZN(n471) );
  OAI21_X1 U29 ( .B1(n283), .B2(n480), .A(n470), .ZN(n367) );
  NAND2_X1 U30 ( .A1(\mem[1][9] ), .A2(n480), .ZN(n470) );
  OAI21_X1 U31 ( .B1(n282), .B2(n480), .A(n469), .ZN(n366) );
  NAND2_X1 U32 ( .A1(\mem[1][10] ), .A2(n480), .ZN(n469) );
  OAI21_X1 U33 ( .B1(n281), .B2(n480), .A(n468), .ZN(n365) );
  NAND2_X1 U34 ( .A1(\mem[1][11] ), .A2(n480), .ZN(n468) );
  OAI21_X1 U35 ( .B1(n292), .B2(n467), .A(n466), .ZN(n364) );
  NAND2_X1 U36 ( .A1(\mem[2][0] ), .A2(n467), .ZN(n466) );
  OAI21_X1 U37 ( .B1(n291), .B2(n467), .A(n465), .ZN(n363) );
  NAND2_X1 U38 ( .A1(\mem[2][1] ), .A2(n467), .ZN(n465) );
  OAI21_X1 U39 ( .B1(n290), .B2(n467), .A(n464), .ZN(n362) );
  NAND2_X1 U40 ( .A1(\mem[2][2] ), .A2(n467), .ZN(n464) );
  OAI21_X1 U41 ( .B1(n289), .B2(n467), .A(n463), .ZN(n361) );
  NAND2_X1 U42 ( .A1(\mem[2][3] ), .A2(n467), .ZN(n463) );
  OAI21_X1 U43 ( .B1(n288), .B2(n467), .A(n462), .ZN(n360) );
  NAND2_X1 U44 ( .A1(\mem[2][4] ), .A2(n467), .ZN(n462) );
  OAI21_X1 U45 ( .B1(n287), .B2(n467), .A(n461), .ZN(n359) );
  NAND2_X1 U46 ( .A1(\mem[2][5] ), .A2(n467), .ZN(n461) );
  OAI21_X1 U47 ( .B1(n286), .B2(n467), .A(n460), .ZN(n358) );
  NAND2_X1 U48 ( .A1(\mem[2][6] ), .A2(n467), .ZN(n460) );
  OAI21_X1 U49 ( .B1(n285), .B2(n467), .A(n459), .ZN(n357) );
  NAND2_X1 U50 ( .A1(\mem[2][7] ), .A2(n467), .ZN(n459) );
  OAI21_X1 U51 ( .B1(n284), .B2(n467), .A(n458), .ZN(n356) );
  NAND2_X1 U52 ( .A1(\mem[2][8] ), .A2(n467), .ZN(n458) );
  OAI21_X1 U53 ( .B1(n283), .B2(n467), .A(n457), .ZN(n355) );
  NAND2_X1 U54 ( .A1(\mem[2][9] ), .A2(n467), .ZN(n457) );
  OAI21_X1 U55 ( .B1(n282), .B2(n467), .A(n456), .ZN(n354) );
  NAND2_X1 U56 ( .A1(\mem[2][10] ), .A2(n467), .ZN(n456) );
  OAI21_X1 U57 ( .B1(n281), .B2(n467), .A(n455), .ZN(n353) );
  NAND2_X1 U58 ( .A1(\mem[2][11] ), .A2(n467), .ZN(n455) );
  OAI21_X1 U59 ( .B1(n292), .B2(n454), .A(n453), .ZN(n352) );
  NAND2_X1 U60 ( .A1(\mem[3][0] ), .A2(n454), .ZN(n453) );
  OAI21_X1 U61 ( .B1(n291), .B2(n454), .A(n452), .ZN(n351) );
  NAND2_X1 U62 ( .A1(\mem[3][1] ), .A2(n454), .ZN(n452) );
  OAI21_X1 U63 ( .B1(n290), .B2(n454), .A(n451), .ZN(n350) );
  NAND2_X1 U64 ( .A1(\mem[3][2] ), .A2(n454), .ZN(n451) );
  OAI21_X1 U65 ( .B1(n289), .B2(n454), .A(n450), .ZN(n349) );
  NAND2_X1 U66 ( .A1(\mem[3][3] ), .A2(n454), .ZN(n450) );
  OAI21_X1 U67 ( .B1(n288), .B2(n454), .A(n449), .ZN(n348) );
  NAND2_X1 U68 ( .A1(\mem[3][4] ), .A2(n454), .ZN(n449) );
  OAI21_X1 U69 ( .B1(n287), .B2(n454), .A(n448), .ZN(n347) );
  NAND2_X1 U70 ( .A1(\mem[3][5] ), .A2(n454), .ZN(n448) );
  OAI21_X1 U71 ( .B1(n286), .B2(n454), .A(n447), .ZN(n346) );
  NAND2_X1 U72 ( .A1(\mem[3][6] ), .A2(n454), .ZN(n447) );
  OAI21_X1 U73 ( .B1(n285), .B2(n454), .A(n446), .ZN(n345) );
  NAND2_X1 U74 ( .A1(\mem[3][7] ), .A2(n454), .ZN(n446) );
  OAI21_X1 U75 ( .B1(n284), .B2(n454), .A(n445), .ZN(n344) );
  NAND2_X1 U76 ( .A1(\mem[3][8] ), .A2(n454), .ZN(n445) );
  OAI21_X1 U77 ( .B1(n283), .B2(n454), .A(n444), .ZN(n343) );
  NAND2_X1 U78 ( .A1(\mem[3][9] ), .A2(n454), .ZN(n444) );
  OAI21_X1 U79 ( .B1(n282), .B2(n454), .A(n443), .ZN(n342) );
  NAND2_X1 U80 ( .A1(\mem[3][10] ), .A2(n454), .ZN(n443) );
  OAI21_X1 U81 ( .B1(n281), .B2(n454), .A(n442), .ZN(n341) );
  NAND2_X1 U82 ( .A1(\mem[3][11] ), .A2(n454), .ZN(n442) );
  OAI21_X1 U83 ( .B1(n292), .B2(n441), .A(n440), .ZN(n340) );
  NAND2_X1 U84 ( .A1(\mem[4][0] ), .A2(n441), .ZN(n440) );
  OAI21_X1 U85 ( .B1(n291), .B2(n441), .A(n439), .ZN(n339) );
  NAND2_X1 U86 ( .A1(\mem[4][1] ), .A2(n441), .ZN(n439) );
  OAI21_X1 U87 ( .B1(n290), .B2(n441), .A(n438), .ZN(n338) );
  NAND2_X1 U88 ( .A1(\mem[4][2] ), .A2(n441), .ZN(n438) );
  OAI21_X1 U89 ( .B1(n289), .B2(n441), .A(n437), .ZN(n337) );
  NAND2_X1 U90 ( .A1(\mem[4][3] ), .A2(n441), .ZN(n437) );
  OAI21_X1 U91 ( .B1(n288), .B2(n441), .A(n436), .ZN(n336) );
  NAND2_X1 U92 ( .A1(\mem[4][4] ), .A2(n441), .ZN(n436) );
  OAI21_X1 U93 ( .B1(n287), .B2(n441), .A(n435), .ZN(n335) );
  NAND2_X1 U94 ( .A1(\mem[4][5] ), .A2(n441), .ZN(n435) );
  OAI21_X1 U95 ( .B1(n286), .B2(n441), .A(n434), .ZN(n334) );
  NAND2_X1 U96 ( .A1(\mem[4][6] ), .A2(n441), .ZN(n434) );
  OAI21_X1 U97 ( .B1(n285), .B2(n441), .A(n433), .ZN(n333) );
  NAND2_X1 U98 ( .A1(\mem[4][7] ), .A2(n441), .ZN(n433) );
  OAI21_X1 U99 ( .B1(n284), .B2(n441), .A(n432), .ZN(n332) );
  NAND2_X1 U100 ( .A1(\mem[4][8] ), .A2(n441), .ZN(n432) );
  OAI21_X1 U101 ( .B1(n283), .B2(n441), .A(n431), .ZN(n331) );
  NAND2_X1 U102 ( .A1(\mem[4][9] ), .A2(n441), .ZN(n431) );
  OAI21_X1 U103 ( .B1(n282), .B2(n441), .A(n430), .ZN(n330) );
  NAND2_X1 U104 ( .A1(\mem[4][10] ), .A2(n441), .ZN(n430) );
  OAI21_X1 U105 ( .B1(n281), .B2(n441), .A(n429), .ZN(n329) );
  NAND2_X1 U106 ( .A1(\mem[4][11] ), .A2(n441), .ZN(n429) );
  OAI21_X1 U107 ( .B1(n292), .B2(n427), .A(n426), .ZN(n328) );
  NAND2_X1 U108 ( .A1(\mem[5][0] ), .A2(n427), .ZN(n426) );
  OAI21_X1 U109 ( .B1(n291), .B2(n427), .A(n425), .ZN(n327) );
  NAND2_X1 U110 ( .A1(\mem[5][1] ), .A2(n427), .ZN(n425) );
  OAI21_X1 U111 ( .B1(n290), .B2(n427), .A(n424), .ZN(n326) );
  NAND2_X1 U112 ( .A1(\mem[5][2] ), .A2(n427), .ZN(n424) );
  OAI21_X1 U113 ( .B1(n289), .B2(n427), .A(n423), .ZN(n325) );
  NAND2_X1 U114 ( .A1(\mem[5][3] ), .A2(n427), .ZN(n423) );
  OAI21_X1 U115 ( .B1(n288), .B2(n427), .A(n422), .ZN(n324) );
  NAND2_X1 U116 ( .A1(\mem[5][4] ), .A2(n427), .ZN(n422) );
  OAI21_X1 U117 ( .B1(n287), .B2(n427), .A(n421), .ZN(n323) );
  NAND2_X1 U118 ( .A1(\mem[5][5] ), .A2(n427), .ZN(n421) );
  OAI21_X1 U119 ( .B1(n286), .B2(n427), .A(n420), .ZN(n322) );
  NAND2_X1 U120 ( .A1(\mem[5][6] ), .A2(n427), .ZN(n420) );
  OAI21_X1 U121 ( .B1(n285), .B2(n427), .A(n419), .ZN(n321) );
  NAND2_X1 U122 ( .A1(\mem[5][7] ), .A2(n427), .ZN(n419) );
  OAI21_X1 U123 ( .B1(n284), .B2(n427), .A(n418), .ZN(n320) );
  NAND2_X1 U124 ( .A1(\mem[5][8] ), .A2(n427), .ZN(n418) );
  OAI21_X1 U125 ( .B1(n283), .B2(n427), .A(n417), .ZN(n319) );
  NAND2_X1 U126 ( .A1(\mem[5][9] ), .A2(n427), .ZN(n417) );
  OAI21_X1 U127 ( .B1(n282), .B2(n427), .A(n416), .ZN(n318) );
  NAND2_X1 U128 ( .A1(\mem[5][10] ), .A2(n427), .ZN(n416) );
  OAI21_X1 U129 ( .B1(n281), .B2(n427), .A(n415), .ZN(n317) );
  NAND2_X1 U130 ( .A1(\mem[5][11] ), .A2(n427), .ZN(n415) );
  OAI21_X1 U131 ( .B1(n292), .B2(n414), .A(n413), .ZN(n316) );
  NAND2_X1 U132 ( .A1(\mem[6][0] ), .A2(n414), .ZN(n413) );
  OAI21_X1 U133 ( .B1(n291), .B2(n414), .A(n412), .ZN(n315) );
  NAND2_X1 U134 ( .A1(\mem[6][1] ), .A2(n414), .ZN(n412) );
  OAI21_X1 U135 ( .B1(n290), .B2(n414), .A(n411), .ZN(n314) );
  NAND2_X1 U136 ( .A1(\mem[6][2] ), .A2(n414), .ZN(n411) );
  OAI21_X1 U137 ( .B1(n289), .B2(n414), .A(n410), .ZN(n313) );
  NAND2_X1 U138 ( .A1(\mem[6][3] ), .A2(n414), .ZN(n410) );
  OAI21_X1 U139 ( .B1(n288), .B2(n414), .A(n409), .ZN(n312) );
  NAND2_X1 U140 ( .A1(\mem[6][4] ), .A2(n414), .ZN(n409) );
  OAI21_X1 U141 ( .B1(n287), .B2(n414), .A(n408), .ZN(n311) );
  NAND2_X1 U142 ( .A1(\mem[6][5] ), .A2(n414), .ZN(n408) );
  OAI21_X1 U143 ( .B1(n286), .B2(n414), .A(n407), .ZN(n310) );
  NAND2_X1 U144 ( .A1(\mem[6][6] ), .A2(n414), .ZN(n407) );
  OAI21_X1 U145 ( .B1(n285), .B2(n414), .A(n406), .ZN(n309) );
  NAND2_X1 U146 ( .A1(\mem[6][7] ), .A2(n414), .ZN(n406) );
  OAI21_X1 U147 ( .B1(n284), .B2(n414), .A(n405), .ZN(n308) );
  NAND2_X1 U148 ( .A1(\mem[6][8] ), .A2(n414), .ZN(n405) );
  OAI21_X1 U149 ( .B1(n283), .B2(n414), .A(n404), .ZN(n307) );
  NAND2_X1 U150 ( .A1(\mem[6][9] ), .A2(n414), .ZN(n404) );
  OAI21_X1 U151 ( .B1(n282), .B2(n414), .A(n403), .ZN(n306) );
  NAND2_X1 U152 ( .A1(\mem[6][10] ), .A2(n414), .ZN(n403) );
  OAI21_X1 U153 ( .B1(n281), .B2(n414), .A(n402), .ZN(n305) );
  NAND2_X1 U154 ( .A1(\mem[6][11] ), .A2(n414), .ZN(n402) );
  OAI21_X1 U155 ( .B1(n292), .B2(n401), .A(n400), .ZN(n304) );
  NAND2_X1 U156 ( .A1(\mem[7][0] ), .A2(n401), .ZN(n400) );
  OAI21_X1 U157 ( .B1(n291), .B2(n401), .A(n399), .ZN(n303) );
  NAND2_X1 U158 ( .A1(\mem[7][1] ), .A2(n401), .ZN(n399) );
  OAI21_X1 U159 ( .B1(n290), .B2(n401), .A(n398), .ZN(n302) );
  NAND2_X1 U160 ( .A1(\mem[7][2] ), .A2(n401), .ZN(n398) );
  OAI21_X1 U161 ( .B1(n289), .B2(n401), .A(n397), .ZN(n301) );
  NAND2_X1 U162 ( .A1(\mem[7][3] ), .A2(n401), .ZN(n397) );
  OAI21_X1 U163 ( .B1(n288), .B2(n401), .A(n396), .ZN(n300) );
  NAND2_X1 U164 ( .A1(\mem[7][4] ), .A2(n401), .ZN(n396) );
  OAI21_X1 U165 ( .B1(n287), .B2(n401), .A(n395), .ZN(n299) );
  NAND2_X1 U166 ( .A1(\mem[7][5] ), .A2(n401), .ZN(n395) );
  OAI21_X1 U167 ( .B1(n286), .B2(n401), .A(n394), .ZN(n298) );
  NAND2_X1 U168 ( .A1(\mem[7][6] ), .A2(n401), .ZN(n394) );
  OAI21_X1 U169 ( .B1(n285), .B2(n401), .A(n393), .ZN(n297) );
  NAND2_X1 U170 ( .A1(\mem[7][7] ), .A2(n401), .ZN(n393) );
  OAI21_X1 U171 ( .B1(n284), .B2(n401), .A(n392), .ZN(n296) );
  NAND2_X1 U172 ( .A1(\mem[7][8] ), .A2(n401), .ZN(n392) );
  OAI21_X1 U173 ( .B1(n283), .B2(n401), .A(n391), .ZN(n295) );
  NAND2_X1 U174 ( .A1(\mem[7][9] ), .A2(n401), .ZN(n391) );
  OAI21_X1 U175 ( .B1(n282), .B2(n401), .A(n390), .ZN(n294) );
  NAND2_X1 U176 ( .A1(\mem[7][10] ), .A2(n401), .ZN(n390) );
  OAI21_X1 U177 ( .B1(n281), .B2(n401), .A(n389), .ZN(n293) );
  NAND2_X1 U178 ( .A1(\mem[7][11] ), .A2(n401), .ZN(n389) );
  OAI21_X1 U179 ( .B1(n494), .B2(n292), .A(n493), .ZN(n388) );
  NAND2_X1 U180 ( .A1(\mem[0][0] ), .A2(n494), .ZN(n493) );
  OAI21_X1 U181 ( .B1(n494), .B2(n291), .A(n492), .ZN(n387) );
  NAND2_X1 U182 ( .A1(\mem[0][1] ), .A2(n494), .ZN(n492) );
  OAI21_X1 U183 ( .B1(n494), .B2(n290), .A(n491), .ZN(n386) );
  NAND2_X1 U184 ( .A1(\mem[0][2] ), .A2(n494), .ZN(n491) );
  OAI21_X1 U185 ( .B1(n494), .B2(n289), .A(n490), .ZN(n385) );
  NAND2_X1 U186 ( .A1(\mem[0][3] ), .A2(n494), .ZN(n490) );
  OAI21_X1 U187 ( .B1(n494), .B2(n288), .A(n489), .ZN(n384) );
  NAND2_X1 U188 ( .A1(\mem[0][4] ), .A2(n494), .ZN(n489) );
  OAI21_X1 U189 ( .B1(n494), .B2(n287), .A(n488), .ZN(n383) );
  NAND2_X1 U190 ( .A1(\mem[0][5] ), .A2(n494), .ZN(n488) );
  OAI21_X1 U191 ( .B1(n494), .B2(n286), .A(n487), .ZN(n382) );
  NAND2_X1 U192 ( .A1(\mem[0][6] ), .A2(n494), .ZN(n487) );
  OAI21_X1 U193 ( .B1(n494), .B2(n285), .A(n486), .ZN(n381) );
  NAND2_X1 U194 ( .A1(\mem[0][7] ), .A2(n494), .ZN(n486) );
  OAI21_X1 U195 ( .B1(n494), .B2(n284), .A(n485), .ZN(n380) );
  NAND2_X1 U196 ( .A1(\mem[0][8] ), .A2(n494), .ZN(n485) );
  OAI21_X1 U197 ( .B1(n494), .B2(n283), .A(n484), .ZN(n379) );
  NAND2_X1 U198 ( .A1(\mem[0][9] ), .A2(n494), .ZN(n484) );
  OAI21_X1 U199 ( .B1(n494), .B2(n282), .A(n483), .ZN(n378) );
  NAND2_X1 U200 ( .A1(\mem[0][10] ), .A2(n494), .ZN(n483) );
  OAI21_X1 U201 ( .B1(n494), .B2(n281), .A(n482), .ZN(n377) );
  NAND2_X1 U202 ( .A1(\mem[0][11] ), .A2(n494), .ZN(n482) );
  INV_X1 U203 ( .A(data_in[0]), .ZN(n292) );
  INV_X1 U204 ( .A(data_in[1]), .ZN(n291) );
  INV_X1 U205 ( .A(data_in[2]), .ZN(n290) );
  INV_X1 U206 ( .A(data_in[3]), .ZN(n289) );
  INV_X1 U207 ( .A(data_in[4]), .ZN(n288) );
  INV_X1 U208 ( .A(data_in[5]), .ZN(n287) );
  INV_X1 U209 ( .A(data_in[6]), .ZN(n286) );
  INV_X1 U210 ( .A(data_in[7]), .ZN(n285) );
  INV_X1 U211 ( .A(data_in[8]), .ZN(n284) );
  INV_X1 U220 ( .A(data_in[9]), .ZN(n283) );
  INV_X1 U221 ( .A(data_in[10]), .ZN(n282) );
  INV_X1 U222 ( .A(data_in[11]), .ZN(n281) );
  MUX2_X1 U223 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n277), .Z(n1) );
  MUX2_X1 U224 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(N10), .Z(n2) );
  MUX2_X1 U225 ( .A(n2), .B(n1), .S(n275), .Z(n3) );
  MUX2_X1 U226 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n277), .Z(n4) );
  MUX2_X1 U227 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n5) );
  MUX2_X1 U228 ( .A(n5), .B(n4), .S(n275), .Z(n6) );
  MUX2_X1 U229 ( .A(n6), .B(n3), .S(N12), .Z(N24) );
  MUX2_X1 U230 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n277), .Z(n7) );
  MUX2_X1 U231 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(N10), .Z(n8) );
  MUX2_X1 U232 ( .A(n8), .B(n7), .S(n275), .Z(n9) );
  MUX2_X1 U233 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n277), .Z(n10) );
  MUX2_X1 U234 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(N10), .Z(n11) );
  MUX2_X1 U235 ( .A(n11), .B(n10), .S(n275), .Z(n12) );
  MUX2_X1 U236 ( .A(n12), .B(n9), .S(N12), .Z(N23) );
  MUX2_X1 U237 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(N10), .Z(n13) );
  MUX2_X1 U238 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(N10), .Z(n14) );
  MUX2_X1 U239 ( .A(n14), .B(n13), .S(n275), .Z(n15) );
  MUX2_X1 U240 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(N10), .Z(n218) );
  MUX2_X1 U241 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(N10), .Z(n219) );
  MUX2_X1 U242 ( .A(n219), .B(n218), .S(n275), .Z(n220) );
  MUX2_X1 U243 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n276), .Z(n221) );
  MUX2_X1 U244 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n276), .Z(n222) );
  MUX2_X1 U245 ( .A(n222), .B(n221), .S(n275), .Z(n223) );
  MUX2_X1 U246 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n276), .Z(n224) );
  MUX2_X1 U247 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n276), .Z(n225) );
  MUX2_X1 U248 ( .A(n225), .B(n224), .S(n275), .Z(n226) );
  MUX2_X1 U249 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n276), .Z(n227) );
  MUX2_X1 U250 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n276), .Z(n228) );
  MUX2_X1 U251 ( .A(n228), .B(n227), .S(n275), .Z(n229) );
  MUX2_X1 U252 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n276), .Z(n230) );
  MUX2_X1 U253 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n276), .Z(n231) );
  MUX2_X1 U254 ( .A(n231), .B(n230), .S(n275), .Z(n232) );
  MUX2_X1 U255 ( .A(n232), .B(n229), .S(N12), .Z(N20) );
  MUX2_X1 U256 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n276), .Z(n233) );
  MUX2_X1 U257 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n276), .Z(n234) );
  MUX2_X1 U258 ( .A(n234), .B(n233), .S(n275), .Z(n235) );
  MUX2_X1 U259 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n276), .Z(n236) );
  MUX2_X1 U260 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n276), .Z(n237) );
  MUX2_X1 U261 ( .A(n237), .B(n236), .S(n275), .Z(n238) );
  MUX2_X1 U262 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n277), .Z(n239) );
  MUX2_X1 U263 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n277), .Z(n240) );
  MUX2_X1 U264 ( .A(n240), .B(n239), .S(n275), .Z(n241) );
  MUX2_X1 U265 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n277), .Z(n242) );
  MUX2_X1 U266 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n277), .Z(n243) );
  MUX2_X1 U267 ( .A(n243), .B(n242), .S(n275), .Z(n244) );
  MUX2_X1 U268 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n277), .Z(n245) );
  MUX2_X1 U269 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n277), .Z(n246) );
  MUX2_X1 U270 ( .A(n246), .B(n245), .S(n275), .Z(n247) );
  MUX2_X1 U271 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n277), .Z(n248) );
  MUX2_X1 U272 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n277), .Z(n249) );
  MUX2_X1 U273 ( .A(n249), .B(n248), .S(n275), .Z(n250) );
  MUX2_X1 U274 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n277), .Z(n251) );
  MUX2_X1 U275 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n277), .Z(n252) );
  MUX2_X1 U276 ( .A(n252), .B(n251), .S(n275), .Z(n253) );
  MUX2_X1 U277 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n277), .Z(n254) );
  MUX2_X1 U278 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n277), .Z(n255) );
  MUX2_X1 U279 ( .A(n255), .B(n254), .S(n275), .Z(n256) );
  MUX2_X1 U280 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n276), .Z(n257) );
  MUX2_X1 U281 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n276), .Z(n258) );
  MUX2_X1 U282 ( .A(n258), .B(n257), .S(n275), .Z(n259) );
  MUX2_X1 U283 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n276), .Z(n260) );
  MUX2_X1 U284 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(N10), .Z(n261) );
  MUX2_X1 U285 ( .A(n261), .B(n260), .S(n275), .Z(n262) );
  MUX2_X1 U286 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n276), .Z(n263) );
  MUX2_X1 U287 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n276), .Z(n264) );
  MUX2_X1 U288 ( .A(n264), .B(n263), .S(n275), .Z(n265) );
  MUX2_X1 U289 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(N10), .Z(n266) );
  MUX2_X1 U290 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(N10), .Z(n267) );
  MUX2_X1 U291 ( .A(n267), .B(n266), .S(n275), .Z(n268) );
  MUX2_X1 U292 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n276), .Z(n269) );
  MUX2_X1 U293 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n277), .Z(n270) );
  MUX2_X1 U294 ( .A(n270), .B(n269), .S(n275), .Z(n271) );
  MUX2_X1 U295 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(N10), .Z(n272) );
  MUX2_X1 U296 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(N10), .Z(n273) );
  MUX2_X1 U297 ( .A(n273), .B(n272), .S(N11), .Z(n274) );
endmodule


module memory_WIDTH24_SIZE8_LOGSIZE3 ( clk, data_in, data_out, addr, wr_en );
  input [23:0] data_in;
  output [23:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][23] , \mem[7][22] , \mem[7][21] , \mem[7][20] ,
         \mem[7][19] , \mem[7][18] , \mem[7][17] , \mem[7][16] , \mem[7][15] ,
         \mem[7][14] , \mem[7][13] , \mem[7][12] , \mem[7][11] , \mem[7][10] ,
         \mem[7][9] , \mem[7][8] , \mem[7][7] , \mem[7][6] , \mem[7][5] ,
         \mem[7][4] , \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] ,
         \mem[6][23] , \mem[6][22] , \mem[6][21] , \mem[6][20] , \mem[6][19] ,
         \mem[6][18] , \mem[6][17] , \mem[6][16] , \mem[6][15] , \mem[6][14] ,
         \mem[6][13] , \mem[6][12] , \mem[6][11] , \mem[6][10] , \mem[6][9] ,
         \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] ,
         \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[5][23] ,
         \mem[5][22] , \mem[5][21] , \mem[5][20] , \mem[5][19] , \mem[5][18] ,
         \mem[5][17] , \mem[5][16] , \mem[5][15] , \mem[5][14] , \mem[5][13] ,
         \mem[5][12] , \mem[5][11] , \mem[5][10] , \mem[5][9] , \mem[5][8] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][23] , \mem[4][22] ,
         \mem[4][21] , \mem[4][20] , \mem[4][19] , \mem[4][18] , \mem[4][17] ,
         \mem[4][16] , \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] ,
         \mem[4][11] , \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] ,
         \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] ,
         \mem[4][1] , \mem[4][0] , \mem[3][23] , \mem[3][22] , \mem[3][21] ,
         \mem[3][20] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][23] , \mem[2][22] , \mem[2][21] , \mem[2][20] ,
         \mem[2][19] , \mem[2][18] , \mem[2][17] , \mem[2][16] , \mem[2][15] ,
         \mem[2][14] , \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] ,
         \mem[2][9] , \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] ,
         \mem[2][4] , \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] ,
         \mem[1][23] , \mem[1][22] , \mem[1][21] , \mem[1][20] , \mem[1][19] ,
         \mem[1][18] , \mem[1][17] , \mem[1][16] , \mem[1][15] , \mem[1][14] ,
         \mem[1][13] , \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] ,
         \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] ,
         \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][23] ,
         \mem[0][22] , \mem[0][21] , \mem[0][20] , \mem[0][19] , \mem[0][18] ,
         \mem[0][17] , \mem[0][16] , \mem[0][15] , \mem[0][14] , \mem[0][13] ,
         \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] , \mem[0][8] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[23]  ( .D(N13), .CK(clk), .Q(data_out[23]) );
  DFF_X1 \data_out_reg[22]  ( .D(N14), .CK(clk), .Q(data_out[22]) );
  DFF_X1 \data_out_reg[21]  ( .D(N15), .CK(clk), .Q(data_out[21]) );
  DFF_X1 \data_out_reg[20]  ( .D(N16), .CK(clk), .Q(data_out[20]) );
  DFF_X1 \data_out_reg[19]  ( .D(N17), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \data_out_reg[18]  ( .D(N18), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[17]  ( .D(N19), .CK(clk), .Q(data_out[17]) );
  DFF_X1 \data_out_reg[16]  ( .D(N20), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[15]  ( .D(N21), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N22), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(N23), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(N24), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(N25), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N26), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N27), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N28), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N29), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N30), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N31), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N32), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N33), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N34), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N35), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N36), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][23]  ( .D(n421), .CK(clk), .Q(\mem[7][23] ) );
  DFF_X1 \mem_reg[7][22]  ( .D(n420), .CK(clk), .Q(\mem[7][22] ) );
  DFF_X1 \mem_reg[7][21]  ( .D(n419), .CK(clk), .Q(\mem[7][21] ) );
  DFF_X1 \mem_reg[7][20]  ( .D(n418), .CK(clk), .Q(\mem[7][20] ) );
  DFF_X1 \mem_reg[7][19]  ( .D(n417), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n416), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n415), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n414), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n413), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n412), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n411), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n410), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n409), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n408), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n407), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n406), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n405), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n404), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n403), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n402), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n401), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n400), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n399), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n398), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][23]  ( .D(n397), .CK(clk), .Q(\mem[6][23] ) );
  DFF_X1 \mem_reg[6][22]  ( .D(n396), .CK(clk), .Q(\mem[6][22] ) );
  DFF_X1 \mem_reg[6][21]  ( .D(n395), .CK(clk), .Q(\mem[6][21] ) );
  DFF_X1 \mem_reg[6][20]  ( .D(n394), .CK(clk), .Q(\mem[6][20] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n393), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n392), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n391), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n390), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n389), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n388), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n387), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n386), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n385), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n384), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n383), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n382), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n381), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n380), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n379), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n378), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n377), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n376), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n375), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n374), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][23]  ( .D(n373), .CK(clk), .Q(\mem[5][23] ) );
  DFF_X1 \mem_reg[5][22]  ( .D(n372), .CK(clk), .Q(\mem[5][22] ) );
  DFF_X1 \mem_reg[5][21]  ( .D(n371), .CK(clk), .Q(\mem[5][21] ) );
  DFF_X1 \mem_reg[5][20]  ( .D(n370), .CK(clk), .Q(\mem[5][20] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n369), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n368), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n367), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n366), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n365), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n364), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n363), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n362), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n361), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n360), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n359), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n358), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n357), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n356), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n355), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n354), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n353), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n352), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n351), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n350), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][23]  ( .D(n349), .CK(clk), .Q(\mem[4][23] ) );
  DFF_X1 \mem_reg[4][22]  ( .D(n348), .CK(clk), .Q(\mem[4][22] ) );
  DFF_X1 \mem_reg[4][21]  ( .D(n347), .CK(clk), .Q(\mem[4][21] ) );
  DFF_X1 \mem_reg[4][20]  ( .D(n346), .CK(clk), .Q(\mem[4][20] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n345), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n344), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n343), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n342), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n341), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n340), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n339), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n338), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n337), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n336), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n335), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n334), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n333), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n332), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n331), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n330), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n329), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n328), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n327), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n326), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][23]  ( .D(n325), .CK(clk), .Q(\mem[3][23] ) );
  DFF_X1 \mem_reg[3][22]  ( .D(n324), .CK(clk), .Q(\mem[3][22] ) );
  DFF_X1 \mem_reg[3][21]  ( .D(n323), .CK(clk), .Q(\mem[3][21] ) );
  DFF_X1 \mem_reg[3][20]  ( .D(n322), .CK(clk), .Q(\mem[3][20] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n321), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n320), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n319), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n318), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n317), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n316), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n315), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n314), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n313), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n312), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n311), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n310), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n309), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n308), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n307), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n306), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n305), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n304), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n303), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n302), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][23]  ( .D(n301), .CK(clk), .Q(\mem[2][23] ) );
  DFF_X1 \mem_reg[2][22]  ( .D(n300), .CK(clk), .Q(\mem[2][22] ) );
  DFF_X1 \mem_reg[2][21]  ( .D(n299), .CK(clk), .Q(\mem[2][21] ) );
  DFF_X1 \mem_reg[2][20]  ( .D(n298), .CK(clk), .Q(\mem[2][20] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n297), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n296), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n295), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n294), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n293), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n292), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n291), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n290), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n289), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n288), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n287), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n286), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n285), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n284), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n283), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n282), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n281), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n280), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n279), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n278), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][23]  ( .D(n277), .CK(clk), .Q(\mem[1][23] ) );
  DFF_X1 \mem_reg[1][22]  ( .D(n276), .CK(clk), .Q(\mem[1][22] ) );
  DFF_X1 \mem_reg[1][21]  ( .D(n275), .CK(clk), .Q(\mem[1][21] ) );
  DFF_X1 \mem_reg[1][20]  ( .D(n274), .CK(clk), .Q(\mem[1][20] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n273), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n272), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n271), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n270), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n269), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n268), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n267), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n266), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n265), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n264), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n263), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n262), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n261), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n260), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n259), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n258), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n257), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n256), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n255), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n254), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][23]  ( .D(n253), .CK(clk), .Q(\mem[0][23] ) );
  DFF_X1 \mem_reg[0][22]  ( .D(n252), .CK(clk), .Q(\mem[0][22] ) );
  DFF_X1 \mem_reg[0][21]  ( .D(n251), .CK(clk), .Q(\mem[0][21] ) );
  DFF_X1 \mem_reg[0][20]  ( .D(n250), .CK(clk), .Q(\mem[0][20] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n249), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n248), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n247), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n246), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n245), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n244), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n243), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n242), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n241), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n240), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n239), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n238), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n237), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n236), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n235), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n234), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n233), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n232), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n231), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n230), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U416 ( .A1(n554), .A2(n555), .A3(n53), .ZN(n28) );
  NAND3_X1 U417 ( .A1(n53), .A2(n555), .A3(N10), .ZN(n54) );
  NAND3_X1 U418 ( .A1(n53), .A2(n554), .A3(N11), .ZN(n79) );
  NAND3_X1 U419 ( .A1(N10), .A2(n53), .A3(N11), .ZN(n104) );
  NAND3_X1 U420 ( .A1(n554), .A2(n555), .A3(n154), .ZN(n129) );
  NAND3_X1 U421 ( .A1(N10), .A2(n555), .A3(n154), .ZN(n155) );
  NAND3_X1 U422 ( .A1(N11), .A2(n554), .A3(n154), .ZN(n180) );
  NAND3_X1 U423 ( .A1(N11), .A2(N10), .A3(n154), .ZN(n205) );
  BUF_X1 U3 ( .A(n545), .Z(n542) );
  BUF_X1 U4 ( .A(n545), .Z(n543) );
  BUF_X1 U5 ( .A(n545), .Z(n544) );
  BUF_X1 U6 ( .A(n541), .Z(n540) );
  BUF_X1 U7 ( .A(n155), .Z(n548) );
  BUF_X1 U8 ( .A(n205), .Z(n546) );
  BUF_X1 U9 ( .A(n129), .Z(n549) );
  BUF_X1 U10 ( .A(N11), .Z(n541) );
  BUF_X1 U11 ( .A(n28), .Z(n553) );
  BUF_X1 U12 ( .A(n54), .Z(n552) );
  BUF_X1 U13 ( .A(n104), .Z(n550) );
  BUF_X1 U14 ( .A(n180), .Z(n547) );
  BUF_X1 U15 ( .A(n79), .Z(n551) );
  INV_X1 U16 ( .A(N10), .ZN(n554) );
  INV_X1 U17 ( .A(N11), .ZN(n555) );
  BUF_X1 U18 ( .A(N12), .Z(n539) );
  NOR2_X1 U19 ( .A1(n556), .A2(N12), .ZN(n53) );
  INV_X1 U20 ( .A(wr_en), .ZN(n556) );
  AND2_X1 U21 ( .A1(N12), .A2(wr_en), .ZN(n154) );
  OAI21_X1 U22 ( .B1(n576), .B2(n54), .A(n59), .ZN(n258) );
  NAND2_X1 U23 ( .A1(\mem[1][4] ), .A2(n552), .ZN(n59) );
  OAI21_X1 U24 ( .B1(n575), .B2(n54), .A(n60), .ZN(n259) );
  NAND2_X1 U25 ( .A1(\mem[1][5] ), .A2(n552), .ZN(n60) );
  OAI21_X1 U26 ( .B1(n574), .B2(n54), .A(n61), .ZN(n260) );
  NAND2_X1 U27 ( .A1(\mem[1][6] ), .A2(n552), .ZN(n61) );
  OAI21_X1 U28 ( .B1(n573), .B2(n54), .A(n62), .ZN(n261) );
  NAND2_X1 U29 ( .A1(\mem[1][7] ), .A2(n552), .ZN(n62) );
  OAI21_X1 U30 ( .B1(n572), .B2(n54), .A(n63), .ZN(n262) );
  NAND2_X1 U31 ( .A1(\mem[1][8] ), .A2(n552), .ZN(n63) );
  OAI21_X1 U32 ( .B1(n571), .B2(n54), .A(n64), .ZN(n263) );
  NAND2_X1 U33 ( .A1(\mem[1][9] ), .A2(n552), .ZN(n64) );
  OAI21_X1 U34 ( .B1(n570), .B2(n54), .A(n65), .ZN(n264) );
  NAND2_X1 U35 ( .A1(\mem[1][10] ), .A2(n552), .ZN(n65) );
  OAI21_X1 U36 ( .B1(n569), .B2(n552), .A(n66), .ZN(n265) );
  NAND2_X1 U37 ( .A1(\mem[1][11] ), .A2(n552), .ZN(n66) );
  OAI21_X1 U38 ( .B1(n568), .B2(n552), .A(n67), .ZN(n266) );
  NAND2_X1 U39 ( .A1(\mem[1][12] ), .A2(n552), .ZN(n67) );
  OAI21_X1 U40 ( .B1(n567), .B2(n54), .A(n68), .ZN(n267) );
  NAND2_X1 U41 ( .A1(\mem[1][13] ), .A2(n552), .ZN(n68) );
  OAI21_X1 U42 ( .B1(n566), .B2(n54), .A(n69), .ZN(n268) );
  NAND2_X1 U43 ( .A1(\mem[1][14] ), .A2(n552), .ZN(n69) );
  OAI21_X1 U44 ( .B1(n565), .B2(n54), .A(n70), .ZN(n269) );
  NAND2_X1 U45 ( .A1(\mem[1][15] ), .A2(n552), .ZN(n70) );
  OAI21_X1 U46 ( .B1(n564), .B2(n54), .A(n71), .ZN(n270) );
  NAND2_X1 U47 ( .A1(\mem[1][16] ), .A2(n552), .ZN(n71) );
  OAI21_X1 U48 ( .B1(n563), .B2(n54), .A(n72), .ZN(n271) );
  NAND2_X1 U49 ( .A1(\mem[1][17] ), .A2(n552), .ZN(n72) );
  OAI21_X1 U50 ( .B1(n576), .B2(n551), .A(n84), .ZN(n282) );
  NAND2_X1 U51 ( .A1(\mem[2][4] ), .A2(n551), .ZN(n84) );
  OAI21_X1 U52 ( .B1(n575), .B2(n551), .A(n85), .ZN(n283) );
  NAND2_X1 U53 ( .A1(\mem[2][5] ), .A2(n551), .ZN(n85) );
  OAI21_X1 U54 ( .B1(n574), .B2(n79), .A(n86), .ZN(n284) );
  NAND2_X1 U55 ( .A1(\mem[2][6] ), .A2(n551), .ZN(n86) );
  OAI21_X1 U56 ( .B1(n573), .B2(n79), .A(n87), .ZN(n285) );
  NAND2_X1 U57 ( .A1(\mem[2][7] ), .A2(n551), .ZN(n87) );
  OAI21_X1 U58 ( .B1(n572), .B2(n79), .A(n88), .ZN(n286) );
  NAND2_X1 U59 ( .A1(\mem[2][8] ), .A2(n79), .ZN(n88) );
  OAI21_X1 U60 ( .B1(n571), .B2(n79), .A(n89), .ZN(n287) );
  NAND2_X1 U61 ( .A1(\mem[2][9] ), .A2(n79), .ZN(n89) );
  OAI21_X1 U62 ( .B1(n570), .B2(n79), .A(n90), .ZN(n288) );
  NAND2_X1 U63 ( .A1(\mem[2][10] ), .A2(n79), .ZN(n90) );
  OAI21_X1 U64 ( .B1(n569), .B2(n551), .A(n91), .ZN(n289) );
  NAND2_X1 U65 ( .A1(\mem[2][11] ), .A2(n79), .ZN(n91) );
  OAI21_X1 U66 ( .B1(n568), .B2(n551), .A(n92), .ZN(n290) );
  NAND2_X1 U67 ( .A1(\mem[2][12] ), .A2(n79), .ZN(n92) );
  OAI21_X1 U68 ( .B1(n567), .B2(n551), .A(n93), .ZN(n291) );
  NAND2_X1 U69 ( .A1(\mem[2][13] ), .A2(n79), .ZN(n93) );
  OAI21_X1 U70 ( .B1(n566), .B2(n551), .A(n94), .ZN(n292) );
  NAND2_X1 U71 ( .A1(\mem[2][14] ), .A2(n79), .ZN(n94) );
  OAI21_X1 U72 ( .B1(n565), .B2(n551), .A(n95), .ZN(n293) );
  NAND2_X1 U73 ( .A1(\mem[2][15] ), .A2(n79), .ZN(n95) );
  OAI21_X1 U74 ( .B1(n564), .B2(n551), .A(n96), .ZN(n294) );
  NAND2_X1 U75 ( .A1(\mem[2][16] ), .A2(n79), .ZN(n96) );
  OAI21_X1 U76 ( .B1(n563), .B2(n551), .A(n97), .ZN(n295) );
  NAND2_X1 U77 ( .A1(\mem[2][17] ), .A2(n79), .ZN(n97) );
  OAI21_X1 U78 ( .B1(n576), .B2(n104), .A(n109), .ZN(n306) );
  NAND2_X1 U79 ( .A1(\mem[3][4] ), .A2(n550), .ZN(n109) );
  OAI21_X1 U80 ( .B1(n575), .B2(n104), .A(n110), .ZN(n307) );
  NAND2_X1 U81 ( .A1(\mem[3][5] ), .A2(n550), .ZN(n110) );
  OAI21_X1 U82 ( .B1(n574), .B2(n104), .A(n111), .ZN(n308) );
  NAND2_X1 U83 ( .A1(\mem[3][6] ), .A2(n550), .ZN(n111) );
  OAI21_X1 U84 ( .B1(n573), .B2(n104), .A(n112), .ZN(n309) );
  NAND2_X1 U85 ( .A1(\mem[3][7] ), .A2(n550), .ZN(n112) );
  OAI21_X1 U86 ( .B1(n572), .B2(n104), .A(n113), .ZN(n310) );
  NAND2_X1 U87 ( .A1(\mem[3][8] ), .A2(n550), .ZN(n113) );
  OAI21_X1 U88 ( .B1(n571), .B2(n104), .A(n114), .ZN(n311) );
  NAND2_X1 U89 ( .A1(\mem[3][9] ), .A2(n550), .ZN(n114) );
  OAI21_X1 U90 ( .B1(n570), .B2(n104), .A(n115), .ZN(n312) );
  NAND2_X1 U91 ( .A1(\mem[3][10] ), .A2(n550), .ZN(n115) );
  OAI21_X1 U92 ( .B1(n569), .B2(n550), .A(n116), .ZN(n313) );
  NAND2_X1 U93 ( .A1(\mem[3][11] ), .A2(n550), .ZN(n116) );
  OAI21_X1 U94 ( .B1(n568), .B2(n550), .A(n117), .ZN(n314) );
  NAND2_X1 U95 ( .A1(\mem[3][12] ), .A2(n550), .ZN(n117) );
  OAI21_X1 U96 ( .B1(n567), .B2(n104), .A(n118), .ZN(n315) );
  NAND2_X1 U97 ( .A1(\mem[3][13] ), .A2(n550), .ZN(n118) );
  OAI21_X1 U98 ( .B1(n566), .B2(n104), .A(n119), .ZN(n316) );
  NAND2_X1 U99 ( .A1(\mem[3][14] ), .A2(n550), .ZN(n119) );
  OAI21_X1 U100 ( .B1(n565), .B2(n104), .A(n120), .ZN(n317) );
  NAND2_X1 U101 ( .A1(\mem[3][15] ), .A2(n550), .ZN(n120) );
  OAI21_X1 U102 ( .B1(n564), .B2(n104), .A(n121), .ZN(n318) );
  NAND2_X1 U103 ( .A1(\mem[3][16] ), .A2(n550), .ZN(n121) );
  OAI21_X1 U104 ( .B1(n563), .B2(n104), .A(n122), .ZN(n319) );
  NAND2_X1 U105 ( .A1(\mem[3][17] ), .A2(n550), .ZN(n122) );
  OAI21_X1 U106 ( .B1(n576), .B2(n129), .A(n134), .ZN(n330) );
  NAND2_X1 U107 ( .A1(\mem[4][4] ), .A2(n129), .ZN(n134) );
  OAI21_X1 U108 ( .B1(n575), .B2(n549), .A(n135), .ZN(n331) );
  NAND2_X1 U109 ( .A1(\mem[4][5] ), .A2(n129), .ZN(n135) );
  OAI21_X1 U110 ( .B1(n574), .B2(n549), .A(n136), .ZN(n332) );
  NAND2_X1 U111 ( .A1(\mem[4][6] ), .A2(n129), .ZN(n136) );
  OAI21_X1 U112 ( .B1(n573), .B2(n549), .A(n137), .ZN(n333) );
  NAND2_X1 U113 ( .A1(\mem[4][7] ), .A2(n129), .ZN(n137) );
  OAI21_X1 U114 ( .B1(n572), .B2(n549), .A(n138), .ZN(n334) );
  NAND2_X1 U115 ( .A1(\mem[4][8] ), .A2(n129), .ZN(n138) );
  OAI21_X1 U116 ( .B1(n571), .B2(n549), .A(n139), .ZN(n335) );
  NAND2_X1 U117 ( .A1(\mem[4][9] ), .A2(n129), .ZN(n139) );
  OAI21_X1 U118 ( .B1(n570), .B2(n549), .A(n140), .ZN(n336) );
  NAND2_X1 U119 ( .A1(\mem[4][10] ), .A2(n129), .ZN(n140) );
  OAI21_X1 U120 ( .B1(n569), .B2(n549), .A(n141), .ZN(n337) );
  NAND2_X1 U121 ( .A1(\mem[4][11] ), .A2(n129), .ZN(n141) );
  OAI21_X1 U122 ( .B1(n568), .B2(n549), .A(n142), .ZN(n338) );
  NAND2_X1 U123 ( .A1(\mem[4][12] ), .A2(n129), .ZN(n142) );
  OAI21_X1 U124 ( .B1(n567), .B2(n549), .A(n143), .ZN(n339) );
  NAND2_X1 U125 ( .A1(\mem[4][13] ), .A2(n129), .ZN(n143) );
  OAI21_X1 U126 ( .B1(n566), .B2(n549), .A(n144), .ZN(n340) );
  NAND2_X1 U127 ( .A1(\mem[4][14] ), .A2(n129), .ZN(n144) );
  OAI21_X1 U128 ( .B1(n565), .B2(n549), .A(n145), .ZN(n341) );
  NAND2_X1 U129 ( .A1(\mem[4][15] ), .A2(n129), .ZN(n145) );
  OAI21_X1 U130 ( .B1(n564), .B2(n549), .A(n146), .ZN(n342) );
  NAND2_X1 U131 ( .A1(\mem[4][16] ), .A2(n129), .ZN(n146) );
  OAI21_X1 U132 ( .B1(n563), .B2(n549), .A(n147), .ZN(n343) );
  NAND2_X1 U133 ( .A1(\mem[4][17] ), .A2(n129), .ZN(n147) );
  OAI21_X1 U134 ( .B1(n576), .B2(n155), .A(n160), .ZN(n354) );
  NAND2_X1 U135 ( .A1(\mem[5][4] ), .A2(n548), .ZN(n160) );
  OAI21_X1 U136 ( .B1(n575), .B2(n548), .A(n161), .ZN(n355) );
  NAND2_X1 U137 ( .A1(\mem[5][5] ), .A2(n548), .ZN(n161) );
  OAI21_X1 U138 ( .B1(n574), .B2(n548), .A(n162), .ZN(n356) );
  NAND2_X1 U139 ( .A1(\mem[5][6] ), .A2(n548), .ZN(n162) );
  OAI21_X1 U140 ( .B1(n573), .B2(n155), .A(n163), .ZN(n357) );
  NAND2_X1 U141 ( .A1(\mem[5][7] ), .A2(n155), .ZN(n163) );
  OAI21_X1 U142 ( .B1(n572), .B2(n155), .A(n164), .ZN(n358) );
  NAND2_X1 U143 ( .A1(\mem[5][8] ), .A2(n548), .ZN(n164) );
  OAI21_X1 U144 ( .B1(n571), .B2(n155), .A(n165), .ZN(n359) );
  NAND2_X1 U145 ( .A1(\mem[5][9] ), .A2(n548), .ZN(n165) );
  OAI21_X1 U146 ( .B1(n570), .B2(n155), .A(n166), .ZN(n360) );
  NAND2_X1 U147 ( .A1(\mem[5][10] ), .A2(n548), .ZN(n166) );
  OAI21_X1 U148 ( .B1(n569), .B2(n155), .A(n167), .ZN(n361) );
  NAND2_X1 U149 ( .A1(\mem[5][11] ), .A2(n548), .ZN(n167) );
  OAI21_X1 U150 ( .B1(n568), .B2(n548), .A(n168), .ZN(n362) );
  NAND2_X1 U151 ( .A1(\mem[5][12] ), .A2(n548), .ZN(n168) );
  OAI21_X1 U152 ( .B1(n567), .B2(n548), .A(n169), .ZN(n363) );
  NAND2_X1 U153 ( .A1(\mem[5][13] ), .A2(n548), .ZN(n169) );
  OAI21_X1 U154 ( .B1(n566), .B2(n155), .A(n170), .ZN(n364) );
  NAND2_X1 U155 ( .A1(\mem[5][14] ), .A2(n548), .ZN(n170) );
  OAI21_X1 U156 ( .B1(n565), .B2(n155), .A(n171), .ZN(n365) );
  NAND2_X1 U157 ( .A1(\mem[5][15] ), .A2(n548), .ZN(n171) );
  OAI21_X1 U158 ( .B1(n564), .B2(n155), .A(n172), .ZN(n366) );
  NAND2_X1 U159 ( .A1(\mem[5][16] ), .A2(n548), .ZN(n172) );
  OAI21_X1 U160 ( .B1(n563), .B2(n155), .A(n173), .ZN(n367) );
  NAND2_X1 U161 ( .A1(\mem[5][17] ), .A2(n548), .ZN(n173) );
  OAI21_X1 U162 ( .B1(n576), .B2(n547), .A(n185), .ZN(n378) );
  NAND2_X1 U163 ( .A1(\mem[6][4] ), .A2(n180), .ZN(n185) );
  OAI21_X1 U164 ( .B1(n575), .B2(n547), .A(n186), .ZN(n379) );
  NAND2_X1 U165 ( .A1(\mem[6][5] ), .A2(n547), .ZN(n186) );
  OAI21_X1 U166 ( .B1(n574), .B2(n547), .A(n187), .ZN(n380) );
  NAND2_X1 U167 ( .A1(\mem[6][6] ), .A2(n547), .ZN(n187) );
  OAI21_X1 U168 ( .B1(n573), .B2(n547), .A(n188), .ZN(n381) );
  NAND2_X1 U169 ( .A1(\mem[6][7] ), .A2(n180), .ZN(n188) );
  OAI21_X1 U170 ( .B1(n572), .B2(n547), .A(n189), .ZN(n382) );
  NAND2_X1 U171 ( .A1(\mem[6][8] ), .A2(n547), .ZN(n189) );
  OAI21_X1 U172 ( .B1(n571), .B2(n547), .A(n190), .ZN(n383) );
  NAND2_X1 U173 ( .A1(\mem[6][9] ), .A2(n547), .ZN(n190) );
  OAI21_X1 U174 ( .B1(n570), .B2(n547), .A(n191), .ZN(n384) );
  NAND2_X1 U175 ( .A1(\mem[6][10] ), .A2(n547), .ZN(n191) );
  OAI21_X1 U176 ( .B1(n569), .B2(n547), .A(n192), .ZN(n385) );
  NAND2_X1 U177 ( .A1(\mem[6][11] ), .A2(n547), .ZN(n192) );
  OAI21_X1 U178 ( .B1(n568), .B2(n180), .A(n193), .ZN(n386) );
  NAND2_X1 U179 ( .A1(\mem[6][12] ), .A2(n547), .ZN(n193) );
  OAI21_X1 U180 ( .B1(n567), .B2(n180), .A(n194), .ZN(n387) );
  NAND2_X1 U181 ( .A1(\mem[6][13] ), .A2(n180), .ZN(n194) );
  OAI21_X1 U182 ( .B1(n566), .B2(n180), .A(n195), .ZN(n388) );
  NAND2_X1 U183 ( .A1(\mem[6][14] ), .A2(n180), .ZN(n195) );
  OAI21_X1 U184 ( .B1(n565), .B2(n180), .A(n196), .ZN(n389) );
  NAND2_X1 U185 ( .A1(\mem[6][15] ), .A2(n180), .ZN(n196) );
  OAI21_X1 U186 ( .B1(n564), .B2(n180), .A(n197), .ZN(n390) );
  NAND2_X1 U187 ( .A1(\mem[6][16] ), .A2(n547), .ZN(n197) );
  OAI21_X1 U188 ( .B1(n563), .B2(n180), .A(n198), .ZN(n391) );
  NAND2_X1 U189 ( .A1(\mem[6][17] ), .A2(n547), .ZN(n198) );
  OAI21_X1 U190 ( .B1(n576), .B2(n205), .A(n210), .ZN(n402) );
  NAND2_X1 U191 ( .A1(\mem[7][4] ), .A2(n546), .ZN(n210) );
  OAI21_X1 U192 ( .B1(n575), .B2(n546), .A(n211), .ZN(n403) );
  NAND2_X1 U193 ( .A1(\mem[7][5] ), .A2(n546), .ZN(n211) );
  OAI21_X1 U194 ( .B1(n574), .B2(n546), .A(n212), .ZN(n404) );
  NAND2_X1 U195 ( .A1(\mem[7][6] ), .A2(n546), .ZN(n212) );
  OAI21_X1 U196 ( .B1(n573), .B2(n205), .A(n213), .ZN(n405) );
  NAND2_X1 U197 ( .A1(\mem[7][7] ), .A2(n205), .ZN(n213) );
  OAI21_X1 U198 ( .B1(n572), .B2(n205), .A(n214), .ZN(n406) );
  NAND2_X1 U199 ( .A1(\mem[7][8] ), .A2(n546), .ZN(n214) );
  OAI21_X1 U200 ( .B1(n571), .B2(n205), .A(n215), .ZN(n407) );
  NAND2_X1 U201 ( .A1(\mem[7][9] ), .A2(n546), .ZN(n215) );
  OAI21_X1 U202 ( .B1(n570), .B2(n205), .A(n216), .ZN(n408) );
  NAND2_X1 U203 ( .A1(\mem[7][10] ), .A2(n546), .ZN(n216) );
  OAI21_X1 U204 ( .B1(n569), .B2(n205), .A(n217), .ZN(n409) );
  NAND2_X1 U205 ( .A1(\mem[7][11] ), .A2(n546), .ZN(n217) );
  OAI21_X1 U206 ( .B1(n568), .B2(n546), .A(n218), .ZN(n410) );
  NAND2_X1 U207 ( .A1(\mem[7][12] ), .A2(n546), .ZN(n218) );
  OAI21_X1 U208 ( .B1(n567), .B2(n546), .A(n219), .ZN(n411) );
  NAND2_X1 U209 ( .A1(\mem[7][13] ), .A2(n546), .ZN(n219) );
  OAI21_X1 U210 ( .B1(n566), .B2(n205), .A(n220), .ZN(n412) );
  NAND2_X1 U211 ( .A1(\mem[7][14] ), .A2(n546), .ZN(n220) );
  OAI21_X1 U212 ( .B1(n565), .B2(n205), .A(n221), .ZN(n413) );
  NAND2_X1 U213 ( .A1(\mem[7][15] ), .A2(n546), .ZN(n221) );
  OAI21_X1 U214 ( .B1(n564), .B2(n205), .A(n222), .ZN(n414) );
  NAND2_X1 U215 ( .A1(\mem[7][16] ), .A2(n546), .ZN(n222) );
  OAI21_X1 U216 ( .B1(n563), .B2(n205), .A(n223), .ZN(n415) );
  NAND2_X1 U217 ( .A1(\mem[7][17] ), .A2(n546), .ZN(n223) );
  OAI21_X1 U218 ( .B1(n580), .B2(n54), .A(n55), .ZN(n254) );
  NAND2_X1 U219 ( .A1(\mem[1][0] ), .A2(n54), .ZN(n55) );
  OAI21_X1 U220 ( .B1(n579), .B2(n54), .A(n56), .ZN(n255) );
  NAND2_X1 U221 ( .A1(\mem[1][1] ), .A2(n54), .ZN(n56) );
  OAI21_X1 U222 ( .B1(n578), .B2(n54), .A(n57), .ZN(n256) );
  NAND2_X1 U223 ( .A1(\mem[1][2] ), .A2(n552), .ZN(n57) );
  OAI21_X1 U224 ( .B1(n577), .B2(n54), .A(n58), .ZN(n257) );
  NAND2_X1 U225 ( .A1(\mem[1][3] ), .A2(n552), .ZN(n58) );
  OAI21_X1 U226 ( .B1(n562), .B2(n54), .A(n73), .ZN(n272) );
  NAND2_X1 U227 ( .A1(\mem[1][18] ), .A2(n552), .ZN(n73) );
  OAI21_X1 U228 ( .B1(n561), .B2(n54), .A(n74), .ZN(n273) );
  NAND2_X1 U229 ( .A1(\mem[1][19] ), .A2(n552), .ZN(n74) );
  OAI21_X1 U230 ( .B1(n560), .B2(n54), .A(n75), .ZN(n274) );
  NAND2_X1 U231 ( .A1(\mem[1][20] ), .A2(n552), .ZN(n75) );
  OAI21_X1 U232 ( .B1(n559), .B2(n54), .A(n76), .ZN(n275) );
  NAND2_X1 U233 ( .A1(\mem[1][21] ), .A2(n552), .ZN(n76) );
  OAI21_X1 U234 ( .B1(n558), .B2(n54), .A(n77), .ZN(n276) );
  NAND2_X1 U235 ( .A1(\mem[1][22] ), .A2(n552), .ZN(n77) );
  OAI21_X1 U236 ( .B1(n557), .B2(n54), .A(n78), .ZN(n277) );
  NAND2_X1 U237 ( .A1(\mem[1][23] ), .A2(n552), .ZN(n78) );
  OAI21_X1 U238 ( .B1(n580), .B2(n79), .A(n80), .ZN(n278) );
  NAND2_X1 U239 ( .A1(\mem[2][0] ), .A2(n551), .ZN(n80) );
  OAI21_X1 U240 ( .B1(n579), .B2(n79), .A(n81), .ZN(n279) );
  NAND2_X1 U241 ( .A1(\mem[2][1] ), .A2(n551), .ZN(n81) );
  OAI21_X1 U242 ( .B1(n578), .B2(n79), .A(n82), .ZN(n280) );
  NAND2_X1 U243 ( .A1(\mem[2][2] ), .A2(n551), .ZN(n82) );
  OAI21_X1 U244 ( .B1(n577), .B2(n79), .A(n83), .ZN(n281) );
  NAND2_X1 U245 ( .A1(\mem[2][3] ), .A2(n551), .ZN(n83) );
  OAI21_X1 U246 ( .B1(n562), .B2(n551), .A(n98), .ZN(n296) );
  NAND2_X1 U247 ( .A1(\mem[2][18] ), .A2(n551), .ZN(n98) );
  OAI21_X1 U248 ( .B1(n561), .B2(n79), .A(n99), .ZN(n297) );
  NAND2_X1 U249 ( .A1(\mem[2][19] ), .A2(n551), .ZN(n99) );
  OAI21_X1 U250 ( .B1(n560), .B2(n79), .A(n100), .ZN(n298) );
  NAND2_X1 U251 ( .A1(\mem[2][20] ), .A2(n551), .ZN(n100) );
  OAI21_X1 U252 ( .B1(n559), .B2(n551), .A(n101), .ZN(n299) );
  NAND2_X1 U253 ( .A1(\mem[2][21] ), .A2(n79), .ZN(n101) );
  OAI21_X1 U254 ( .B1(n558), .B2(n551), .A(n102), .ZN(n300) );
  NAND2_X1 U255 ( .A1(\mem[2][22] ), .A2(n79), .ZN(n102) );
  OAI21_X1 U256 ( .B1(n557), .B2(n79), .A(n103), .ZN(n301) );
  NAND2_X1 U257 ( .A1(\mem[2][23] ), .A2(n551), .ZN(n103) );
  OAI21_X1 U258 ( .B1(n580), .B2(n104), .A(n105), .ZN(n302) );
  NAND2_X1 U259 ( .A1(\mem[3][0] ), .A2(n104), .ZN(n105) );
  OAI21_X1 U260 ( .B1(n579), .B2(n104), .A(n106), .ZN(n303) );
  NAND2_X1 U261 ( .A1(\mem[3][1] ), .A2(n104), .ZN(n106) );
  OAI21_X1 U262 ( .B1(n578), .B2(n104), .A(n107), .ZN(n304) );
  NAND2_X1 U263 ( .A1(\mem[3][2] ), .A2(n550), .ZN(n107) );
  OAI21_X1 U264 ( .B1(n577), .B2(n104), .A(n108), .ZN(n305) );
  NAND2_X1 U265 ( .A1(\mem[3][3] ), .A2(n550), .ZN(n108) );
  OAI21_X1 U266 ( .B1(n562), .B2(n104), .A(n123), .ZN(n320) );
  NAND2_X1 U267 ( .A1(\mem[3][18] ), .A2(n550), .ZN(n123) );
  OAI21_X1 U268 ( .B1(n561), .B2(n104), .A(n124), .ZN(n321) );
  NAND2_X1 U269 ( .A1(\mem[3][19] ), .A2(n550), .ZN(n124) );
  OAI21_X1 U270 ( .B1(n560), .B2(n104), .A(n125), .ZN(n322) );
  NAND2_X1 U271 ( .A1(\mem[3][20] ), .A2(n550), .ZN(n125) );
  OAI21_X1 U272 ( .B1(n559), .B2(n104), .A(n126), .ZN(n323) );
  NAND2_X1 U273 ( .A1(\mem[3][21] ), .A2(n550), .ZN(n126) );
  OAI21_X1 U274 ( .B1(n558), .B2(n104), .A(n127), .ZN(n324) );
  NAND2_X1 U275 ( .A1(\mem[3][22] ), .A2(n550), .ZN(n127) );
  OAI21_X1 U276 ( .B1(n557), .B2(n104), .A(n128), .ZN(n325) );
  NAND2_X1 U277 ( .A1(\mem[3][23] ), .A2(n550), .ZN(n128) );
  OAI21_X1 U278 ( .B1(n580), .B2(n549), .A(n130), .ZN(n326) );
  NAND2_X1 U279 ( .A1(\mem[4][0] ), .A2(n129), .ZN(n130) );
  OAI21_X1 U280 ( .B1(n579), .B2(n549), .A(n131), .ZN(n327) );
  NAND2_X1 U281 ( .A1(\mem[4][1] ), .A2(n129), .ZN(n131) );
  OAI21_X1 U282 ( .B1(n578), .B2(n549), .A(n132), .ZN(n328) );
  NAND2_X1 U283 ( .A1(\mem[4][2] ), .A2(n129), .ZN(n132) );
  OAI21_X1 U284 ( .B1(n577), .B2(n549), .A(n133), .ZN(n329) );
  NAND2_X1 U285 ( .A1(\mem[4][3] ), .A2(n129), .ZN(n133) );
  OAI21_X1 U286 ( .B1(n562), .B2(n549), .A(n148), .ZN(n344) );
  NAND2_X1 U287 ( .A1(\mem[4][18] ), .A2(n129), .ZN(n148) );
  OAI21_X1 U288 ( .B1(n561), .B2(n549), .A(n149), .ZN(n345) );
  NAND2_X1 U289 ( .A1(\mem[4][19] ), .A2(n129), .ZN(n149) );
  OAI21_X1 U290 ( .B1(n560), .B2(n549), .A(n150), .ZN(n346) );
  NAND2_X1 U291 ( .A1(\mem[4][20] ), .A2(n129), .ZN(n150) );
  OAI21_X1 U292 ( .B1(n559), .B2(n549), .A(n151), .ZN(n347) );
  NAND2_X1 U293 ( .A1(\mem[4][21] ), .A2(n549), .ZN(n151) );
  OAI21_X1 U294 ( .B1(n558), .B2(n549), .A(n152), .ZN(n348) );
  NAND2_X1 U295 ( .A1(\mem[4][22] ), .A2(n129), .ZN(n152) );
  OAI21_X1 U296 ( .B1(n557), .B2(n549), .A(n153), .ZN(n349) );
  NAND2_X1 U297 ( .A1(\mem[4][23] ), .A2(n129), .ZN(n153) );
  OAI21_X1 U298 ( .B1(n580), .B2(n155), .A(n156), .ZN(n350) );
  NAND2_X1 U299 ( .A1(\mem[5][0] ), .A2(n155), .ZN(n156) );
  OAI21_X1 U300 ( .B1(n579), .B2(n155), .A(n157), .ZN(n351) );
  NAND2_X1 U301 ( .A1(\mem[5][1] ), .A2(n155), .ZN(n157) );
  OAI21_X1 U302 ( .B1(n578), .B2(n155), .A(n158), .ZN(n352) );
  NAND2_X1 U303 ( .A1(\mem[5][2] ), .A2(n155), .ZN(n158) );
  OAI21_X1 U304 ( .B1(n577), .B2(n155), .A(n159), .ZN(n353) );
  NAND2_X1 U305 ( .A1(\mem[5][3] ), .A2(n548), .ZN(n159) );
  OAI21_X1 U306 ( .B1(n562), .B2(n155), .A(n174), .ZN(n368) );
  NAND2_X1 U307 ( .A1(\mem[5][18] ), .A2(n548), .ZN(n174) );
  OAI21_X1 U308 ( .B1(n561), .B2(n155), .A(n175), .ZN(n369) );
  NAND2_X1 U309 ( .A1(\mem[5][19] ), .A2(n548), .ZN(n175) );
  OAI21_X1 U310 ( .B1(n560), .B2(n155), .A(n176), .ZN(n370) );
  NAND2_X1 U311 ( .A1(\mem[5][20] ), .A2(n548), .ZN(n176) );
  OAI21_X1 U312 ( .B1(n559), .B2(n155), .A(n177), .ZN(n371) );
  NAND2_X1 U313 ( .A1(\mem[5][21] ), .A2(n548), .ZN(n177) );
  OAI21_X1 U314 ( .B1(n558), .B2(n155), .A(n178), .ZN(n372) );
  NAND2_X1 U315 ( .A1(\mem[5][22] ), .A2(n548), .ZN(n178) );
  OAI21_X1 U316 ( .B1(n557), .B2(n155), .A(n179), .ZN(n373) );
  NAND2_X1 U317 ( .A1(\mem[5][23] ), .A2(n548), .ZN(n179) );
  OAI21_X1 U318 ( .B1(n580), .B2(n547), .A(n181), .ZN(n374) );
  NAND2_X1 U319 ( .A1(\mem[6][0] ), .A2(n180), .ZN(n181) );
  OAI21_X1 U320 ( .B1(n579), .B2(n547), .A(n182), .ZN(n375) );
  NAND2_X1 U321 ( .A1(\mem[6][1] ), .A2(n180), .ZN(n182) );
  OAI21_X1 U322 ( .B1(n578), .B2(n547), .A(n183), .ZN(n376) );
  NAND2_X1 U323 ( .A1(\mem[6][2] ), .A2(n180), .ZN(n183) );
  OAI21_X1 U324 ( .B1(n577), .B2(n547), .A(n184), .ZN(n377) );
  NAND2_X1 U325 ( .A1(\mem[6][3] ), .A2(n180), .ZN(n184) );
  OAI21_X1 U326 ( .B1(n562), .B2(n180), .A(n199), .ZN(n392) );
  NAND2_X1 U327 ( .A1(\mem[6][18] ), .A2(n547), .ZN(n199) );
  OAI21_X1 U328 ( .B1(n561), .B2(n180), .A(n200), .ZN(n393) );
  NAND2_X1 U329 ( .A1(\mem[6][19] ), .A2(n547), .ZN(n200) );
  OAI21_X1 U330 ( .B1(n560), .B2(n180), .A(n201), .ZN(n394) );
  NAND2_X1 U331 ( .A1(\mem[6][20] ), .A2(n180), .ZN(n201) );
  OAI21_X1 U332 ( .B1(n559), .B2(n180), .A(n202), .ZN(n395) );
  NAND2_X1 U333 ( .A1(\mem[6][21] ), .A2(n180), .ZN(n202) );
  OAI21_X1 U334 ( .B1(n558), .B2(n180), .A(n203), .ZN(n396) );
  NAND2_X1 U335 ( .A1(\mem[6][22] ), .A2(n180), .ZN(n203) );
  OAI21_X1 U336 ( .B1(n557), .B2(n547), .A(n204), .ZN(n397) );
  NAND2_X1 U337 ( .A1(\mem[6][23] ), .A2(n180), .ZN(n204) );
  OAI21_X1 U338 ( .B1(n580), .B2(n205), .A(n206), .ZN(n398) );
  NAND2_X1 U339 ( .A1(\mem[7][0] ), .A2(n205), .ZN(n206) );
  OAI21_X1 U340 ( .B1(n579), .B2(n205), .A(n207), .ZN(n399) );
  NAND2_X1 U341 ( .A1(\mem[7][1] ), .A2(n205), .ZN(n207) );
  OAI21_X1 U342 ( .B1(n578), .B2(n205), .A(n208), .ZN(n400) );
  NAND2_X1 U343 ( .A1(\mem[7][2] ), .A2(n205), .ZN(n208) );
  OAI21_X1 U344 ( .B1(n577), .B2(n205), .A(n209), .ZN(n401) );
  NAND2_X1 U345 ( .A1(\mem[7][3] ), .A2(n546), .ZN(n209) );
  OAI21_X1 U346 ( .B1(n562), .B2(n205), .A(n224), .ZN(n416) );
  NAND2_X1 U347 ( .A1(\mem[7][18] ), .A2(n546), .ZN(n224) );
  OAI21_X1 U348 ( .B1(n561), .B2(n205), .A(n225), .ZN(n417) );
  NAND2_X1 U349 ( .A1(\mem[7][19] ), .A2(n546), .ZN(n225) );
  OAI21_X1 U350 ( .B1(n560), .B2(n205), .A(n226), .ZN(n418) );
  NAND2_X1 U351 ( .A1(\mem[7][20] ), .A2(n546), .ZN(n226) );
  OAI21_X1 U352 ( .B1(n559), .B2(n205), .A(n227), .ZN(n419) );
  NAND2_X1 U353 ( .A1(\mem[7][21] ), .A2(n546), .ZN(n227) );
  OAI21_X1 U354 ( .B1(n558), .B2(n205), .A(n228), .ZN(n420) );
  NAND2_X1 U355 ( .A1(\mem[7][22] ), .A2(n546), .ZN(n228) );
  OAI21_X1 U356 ( .B1(n557), .B2(n205), .A(n229), .ZN(n421) );
  NAND2_X1 U357 ( .A1(\mem[7][23] ), .A2(n546), .ZN(n229) );
  OAI21_X1 U358 ( .B1(n28), .B2(n580), .A(n29), .ZN(n230) );
  NAND2_X1 U359 ( .A1(\mem[0][0] ), .A2(n553), .ZN(n29) );
  OAI21_X1 U360 ( .B1(n28), .B2(n579), .A(n30), .ZN(n231) );
  NAND2_X1 U361 ( .A1(\mem[0][1] ), .A2(n553), .ZN(n30) );
  OAI21_X1 U362 ( .B1(n28), .B2(n578), .A(n31), .ZN(n232) );
  NAND2_X1 U363 ( .A1(\mem[0][2] ), .A2(n553), .ZN(n31) );
  OAI21_X1 U364 ( .B1(n28), .B2(n577), .A(n32), .ZN(n233) );
  NAND2_X1 U365 ( .A1(\mem[0][3] ), .A2(n553), .ZN(n32) );
  OAI21_X1 U366 ( .B1(n28), .B2(n576), .A(n33), .ZN(n234) );
  NAND2_X1 U367 ( .A1(\mem[0][4] ), .A2(n553), .ZN(n33) );
  OAI21_X1 U368 ( .B1(n28), .B2(n575), .A(n34), .ZN(n235) );
  NAND2_X1 U369 ( .A1(\mem[0][5] ), .A2(n553), .ZN(n34) );
  OAI21_X1 U370 ( .B1(n28), .B2(n574), .A(n35), .ZN(n236) );
  NAND2_X1 U371 ( .A1(\mem[0][6] ), .A2(n553), .ZN(n35) );
  OAI21_X1 U372 ( .B1(n28), .B2(n573), .A(n36), .ZN(n237) );
  NAND2_X1 U373 ( .A1(\mem[0][7] ), .A2(n553), .ZN(n36) );
  OAI21_X1 U374 ( .B1(n28), .B2(n572), .A(n37), .ZN(n238) );
  NAND2_X1 U375 ( .A1(\mem[0][8] ), .A2(n553), .ZN(n37) );
  OAI21_X1 U376 ( .B1(n28), .B2(n571), .A(n38), .ZN(n239) );
  NAND2_X1 U377 ( .A1(\mem[0][9] ), .A2(n553), .ZN(n38) );
  OAI21_X1 U378 ( .B1(n28), .B2(n570), .A(n39), .ZN(n240) );
  NAND2_X1 U379 ( .A1(\mem[0][10] ), .A2(n553), .ZN(n39) );
  OAI21_X1 U380 ( .B1(n28), .B2(n569), .A(n40), .ZN(n241) );
  NAND2_X1 U381 ( .A1(\mem[0][11] ), .A2(n553), .ZN(n40) );
  OAI21_X1 U382 ( .B1(n28), .B2(n557), .A(n52), .ZN(n253) );
  NAND2_X1 U383 ( .A1(\mem[0][23] ), .A2(n553), .ZN(n52) );
  OAI21_X1 U384 ( .B1(n553), .B2(n568), .A(n41), .ZN(n242) );
  NAND2_X1 U385 ( .A1(\mem[0][12] ), .A2(n553), .ZN(n41) );
  OAI21_X1 U386 ( .B1(n28), .B2(n567), .A(n42), .ZN(n243) );
  NAND2_X1 U387 ( .A1(\mem[0][13] ), .A2(n553), .ZN(n42) );
  OAI21_X1 U388 ( .B1(n28), .B2(n566), .A(n43), .ZN(n244) );
  NAND2_X1 U389 ( .A1(\mem[0][14] ), .A2(n553), .ZN(n43) );
  OAI21_X1 U390 ( .B1(n28), .B2(n565), .A(n44), .ZN(n245) );
  NAND2_X1 U391 ( .A1(\mem[0][15] ), .A2(n553), .ZN(n44) );
  OAI21_X1 U392 ( .B1(n28), .B2(n564), .A(n45), .ZN(n246) );
  NAND2_X1 U393 ( .A1(\mem[0][16] ), .A2(n553), .ZN(n45) );
  OAI21_X1 U394 ( .B1(n28), .B2(n563), .A(n46), .ZN(n247) );
  NAND2_X1 U395 ( .A1(\mem[0][17] ), .A2(n553), .ZN(n46) );
  OAI21_X1 U396 ( .B1(n28), .B2(n562), .A(n47), .ZN(n248) );
  NAND2_X1 U397 ( .A1(\mem[0][18] ), .A2(n553), .ZN(n47) );
  OAI21_X1 U398 ( .B1(n28), .B2(n561), .A(n48), .ZN(n249) );
  NAND2_X1 U399 ( .A1(\mem[0][19] ), .A2(n553), .ZN(n48) );
  OAI21_X1 U400 ( .B1(n28), .B2(n560), .A(n49), .ZN(n250) );
  NAND2_X1 U401 ( .A1(\mem[0][20] ), .A2(n28), .ZN(n49) );
  OAI21_X1 U402 ( .B1(n28), .B2(n559), .A(n50), .ZN(n251) );
  NAND2_X1 U403 ( .A1(\mem[0][21] ), .A2(n553), .ZN(n50) );
  OAI21_X1 U404 ( .B1(n28), .B2(n558), .A(n51), .ZN(n252) );
  NAND2_X1 U405 ( .A1(\mem[0][22] ), .A2(n553), .ZN(n51) );
  INV_X1 U406 ( .A(data_in[0]), .ZN(n580) );
  INV_X1 U407 ( .A(data_in[1]), .ZN(n579) );
  INV_X1 U408 ( .A(data_in[2]), .ZN(n578) );
  INV_X1 U409 ( .A(data_in[3]), .ZN(n577) );
  INV_X1 U410 ( .A(data_in[4]), .ZN(n576) );
  INV_X1 U411 ( .A(data_in[5]), .ZN(n575) );
  INV_X1 U412 ( .A(data_in[6]), .ZN(n574) );
  INV_X1 U413 ( .A(data_in[7]), .ZN(n573) );
  INV_X1 U414 ( .A(data_in[8]), .ZN(n572) );
  INV_X1 U415 ( .A(data_in[9]), .ZN(n571) );
  INV_X1 U424 ( .A(data_in[10]), .ZN(n570) );
  INV_X1 U425 ( .A(data_in[11]), .ZN(n569) );
  INV_X1 U426 ( .A(data_in[12]), .ZN(n568) );
  INV_X1 U427 ( .A(data_in[13]), .ZN(n567) );
  INV_X1 U428 ( .A(data_in[14]), .ZN(n566) );
  INV_X1 U429 ( .A(data_in[15]), .ZN(n565) );
  INV_X1 U430 ( .A(data_in[16]), .ZN(n564) );
  INV_X1 U431 ( .A(data_in[17]), .ZN(n563) );
  INV_X1 U432 ( .A(data_in[18]), .ZN(n562) );
  INV_X1 U433 ( .A(data_in[19]), .ZN(n561) );
  INV_X1 U434 ( .A(data_in[20]), .ZN(n560) );
  INV_X1 U435 ( .A(data_in[21]), .ZN(n559) );
  INV_X1 U436 ( .A(data_in[22]), .ZN(n558) );
  INV_X1 U437 ( .A(data_in[23]), .ZN(n557) );
  MUX2_X1 U438 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n544), .Z(n1) );
  MUX2_X1 U439 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n542), .Z(n2) );
  MUX2_X1 U440 ( .A(n2), .B(n1), .S(n540), .Z(n3) );
  MUX2_X1 U441 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n545), .Z(n4) );
  MUX2_X1 U442 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n542), .Z(n5) );
  MUX2_X1 U443 ( .A(n5), .B(n4), .S(n540), .Z(n6) );
  MUX2_X1 U444 ( .A(n6), .B(n3), .S(n539), .Z(N36) );
  MUX2_X1 U445 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n542), .Z(n7) );
  MUX2_X1 U446 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n543), .Z(n8) );
  MUX2_X1 U447 ( .A(n8), .B(n7), .S(n540), .Z(n9) );
  MUX2_X1 U448 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n545), .Z(n10) );
  MUX2_X1 U449 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n543), .Z(n11) );
  MUX2_X1 U450 ( .A(n11), .B(n10), .S(n540), .Z(n12) );
  MUX2_X1 U451 ( .A(n12), .B(n9), .S(n539), .Z(N35) );
  MUX2_X1 U452 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n543), .Z(n13) );
  MUX2_X1 U453 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n544), .Z(n14) );
  MUX2_X1 U454 ( .A(n14), .B(n13), .S(n540), .Z(n15) );
  MUX2_X1 U455 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n545), .Z(n16) );
  MUX2_X1 U456 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n544), .Z(n17) );
  MUX2_X1 U457 ( .A(n17), .B(n16), .S(n540), .Z(n18) );
  MUX2_X1 U458 ( .A(n18), .B(n15), .S(n539), .Z(N34) );
  MUX2_X1 U459 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n544), .Z(n19) );
  MUX2_X1 U460 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n20) );
  MUX2_X1 U461 ( .A(n20), .B(n19), .S(n540), .Z(n21) );
  MUX2_X1 U462 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n22) );
  MUX2_X1 U463 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n23) );
  MUX2_X1 U464 ( .A(n23), .B(n22), .S(n540), .Z(n24) );
  MUX2_X1 U465 ( .A(n24), .B(n21), .S(n539), .Z(N33) );
  MUX2_X1 U466 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n542), .Z(n25) );
  MUX2_X1 U467 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(N10), .Z(n26) );
  MUX2_X1 U468 ( .A(n26), .B(n25), .S(n540), .Z(n27) );
  MUX2_X1 U469 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(N10), .Z(n422) );
  MUX2_X1 U470 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n423) );
  MUX2_X1 U471 ( .A(n423), .B(n422), .S(n540), .Z(n424) );
  MUX2_X1 U472 ( .A(n424), .B(n27), .S(n539), .Z(N32) );
  MUX2_X1 U473 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n545), .Z(n425) );
  MUX2_X1 U474 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(N10), .Z(n426) );
  MUX2_X1 U475 ( .A(n426), .B(n425), .S(n540), .Z(n427) );
  MUX2_X1 U476 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n428) );
  MUX2_X1 U477 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n543), .Z(n429) );
  MUX2_X1 U478 ( .A(n429), .B(n428), .S(n540), .Z(n430) );
  MUX2_X1 U479 ( .A(n430), .B(n427), .S(n539), .Z(N31) );
  MUX2_X1 U480 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n542), .Z(n431) );
  MUX2_X1 U481 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n542), .Z(n432) );
  MUX2_X1 U482 ( .A(n432), .B(n431), .S(n541), .Z(n433) );
  MUX2_X1 U483 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n542), .Z(n434) );
  MUX2_X1 U484 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n542), .Z(n435) );
  MUX2_X1 U485 ( .A(n435), .B(n434), .S(n541), .Z(n436) );
  MUX2_X1 U486 ( .A(n436), .B(n433), .S(n539), .Z(N30) );
  MUX2_X1 U487 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n542), .Z(n437) );
  MUX2_X1 U488 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n542), .Z(n438) );
  MUX2_X1 U489 ( .A(n438), .B(n437), .S(n541), .Z(n439) );
  MUX2_X1 U490 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n542), .Z(n440) );
  MUX2_X1 U491 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n542), .Z(n441) );
  MUX2_X1 U492 ( .A(n441), .B(n440), .S(n541), .Z(n442) );
  MUX2_X1 U493 ( .A(n442), .B(n439), .S(n539), .Z(N29) );
  MUX2_X1 U494 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n542), .Z(n443) );
  MUX2_X1 U495 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n542), .Z(n444) );
  MUX2_X1 U496 ( .A(n444), .B(n443), .S(n541), .Z(n445) );
  MUX2_X1 U497 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n542), .Z(n446) );
  MUX2_X1 U498 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n542), .Z(n447) );
  MUX2_X1 U499 ( .A(n447), .B(n446), .S(n541), .Z(n448) );
  MUX2_X1 U500 ( .A(n448), .B(n445), .S(n539), .Z(N28) );
  MUX2_X1 U501 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n543), .Z(n449) );
  MUX2_X1 U502 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n543), .Z(n450) );
  MUX2_X1 U503 ( .A(n450), .B(n449), .S(n541), .Z(n451) );
  MUX2_X1 U504 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n543), .Z(n452) );
  MUX2_X1 U505 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n543), .Z(n453) );
  MUX2_X1 U506 ( .A(n453), .B(n452), .S(n541), .Z(n454) );
  MUX2_X1 U507 ( .A(n454), .B(n451), .S(n539), .Z(N27) );
  MUX2_X1 U508 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n543), .Z(n455) );
  MUX2_X1 U509 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n543), .Z(n456) );
  MUX2_X1 U510 ( .A(n456), .B(n455), .S(n541), .Z(n457) );
  MUX2_X1 U511 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n543), .Z(n458) );
  MUX2_X1 U512 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n543), .Z(n459) );
  MUX2_X1 U513 ( .A(n459), .B(n458), .S(n541), .Z(n460) );
  MUX2_X1 U514 ( .A(n460), .B(n457), .S(n539), .Z(N26) );
  MUX2_X1 U515 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n543), .Z(n461) );
  MUX2_X1 U516 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n543), .Z(n462) );
  MUX2_X1 U517 ( .A(n462), .B(n461), .S(n541), .Z(n463) );
  MUX2_X1 U518 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n543), .Z(n464) );
  MUX2_X1 U519 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n543), .Z(n465) );
  MUX2_X1 U520 ( .A(n465), .B(n464), .S(n541), .Z(n466) );
  MUX2_X1 U521 ( .A(n466), .B(n463), .S(n539), .Z(N25) );
  MUX2_X1 U522 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n544), .Z(n467) );
  MUX2_X1 U523 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n544), .Z(n468) );
  MUX2_X1 U524 ( .A(n468), .B(n467), .S(n541), .Z(n469) );
  MUX2_X1 U525 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n544), .Z(n470) );
  MUX2_X1 U526 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n544), .Z(n471) );
  MUX2_X1 U527 ( .A(n471), .B(n470), .S(n541), .Z(n472) );
  MUX2_X1 U528 ( .A(n472), .B(n469), .S(n539), .Z(N24) );
  MUX2_X1 U529 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n544), .Z(n473) );
  MUX2_X1 U530 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n544), .Z(n474) );
  MUX2_X1 U531 ( .A(n474), .B(n473), .S(N11), .Z(n475) );
  MUX2_X1 U532 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n544), .Z(n476) );
  MUX2_X1 U533 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n544), .Z(n477) );
  MUX2_X1 U534 ( .A(n477), .B(n476), .S(n541), .Z(n478) );
  MUX2_X1 U535 ( .A(n478), .B(n475), .S(n539), .Z(N23) );
  MUX2_X1 U536 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n544), .Z(n479) );
  MUX2_X1 U537 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n544), .Z(n480) );
  MUX2_X1 U538 ( .A(n480), .B(n479), .S(N11), .Z(n481) );
  MUX2_X1 U539 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n544), .Z(n482) );
  MUX2_X1 U540 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n544), .Z(n483) );
  MUX2_X1 U541 ( .A(n483), .B(n482), .S(n541), .Z(n484) );
  MUX2_X1 U542 ( .A(n484), .B(n481), .S(n539), .Z(N22) );
  MUX2_X1 U543 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n545), .Z(n485) );
  MUX2_X1 U544 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n542), .Z(n486) );
  MUX2_X1 U545 ( .A(n486), .B(n485), .S(N11), .Z(n487) );
  MUX2_X1 U546 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n545), .Z(n488) );
  MUX2_X1 U547 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n545), .Z(n489) );
  MUX2_X1 U548 ( .A(n489), .B(n488), .S(n541), .Z(n490) );
  MUX2_X1 U549 ( .A(n490), .B(n487), .S(n539), .Z(N21) );
  MUX2_X1 U550 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(N10), .Z(n491) );
  MUX2_X1 U551 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(n545), .Z(n492) );
  MUX2_X1 U552 ( .A(n492), .B(n491), .S(N11), .Z(n493) );
  MUX2_X1 U553 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(n544), .Z(n494) );
  MUX2_X1 U554 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(N10), .Z(n495) );
  MUX2_X1 U555 ( .A(n495), .B(n494), .S(n541), .Z(n496) );
  MUX2_X1 U556 ( .A(n496), .B(n493), .S(n539), .Z(N20) );
  MUX2_X1 U557 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n545), .Z(n497) );
  MUX2_X1 U558 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n545), .Z(n498) );
  MUX2_X1 U559 ( .A(n498), .B(n497), .S(n541), .Z(n499) );
  MUX2_X1 U560 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n545), .Z(n500) );
  MUX2_X1 U561 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(N10), .Z(n501) );
  MUX2_X1 U562 ( .A(n501), .B(n500), .S(n541), .Z(n502) );
  MUX2_X1 U563 ( .A(n502), .B(n499), .S(n539), .Z(N19) );
  MUX2_X1 U564 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n543), .Z(n503) );
  MUX2_X1 U565 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n542), .Z(n504) );
  MUX2_X1 U566 ( .A(n504), .B(n503), .S(n541), .Z(n505) );
  MUX2_X1 U567 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n545), .Z(n506) );
  MUX2_X1 U568 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n543), .Z(n507) );
  MUX2_X1 U569 ( .A(n507), .B(n506), .S(N11), .Z(n508) );
  MUX2_X1 U570 ( .A(n508), .B(n505), .S(n539), .Z(N18) );
  MUX2_X1 U571 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(n543), .Z(n509) );
  MUX2_X1 U572 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n545), .Z(n510) );
  MUX2_X1 U573 ( .A(n510), .B(n509), .S(n541), .Z(n511) );
  MUX2_X1 U574 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n544), .Z(n512) );
  MUX2_X1 U575 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(n544), .Z(n513) );
  MUX2_X1 U576 ( .A(n513), .B(n512), .S(N11), .Z(n514) );
  MUX2_X1 U577 ( .A(n514), .B(n511), .S(n539), .Z(N17) );
  MUX2_X1 U578 ( .A(\mem[6][20] ), .B(\mem[7][20] ), .S(n545), .Z(n515) );
  MUX2_X1 U579 ( .A(\mem[4][20] ), .B(\mem[5][20] ), .S(n545), .Z(n516) );
  MUX2_X1 U580 ( .A(n516), .B(n515), .S(N11), .Z(n517) );
  MUX2_X1 U581 ( .A(\mem[2][20] ), .B(\mem[3][20] ), .S(n545), .Z(n518) );
  MUX2_X1 U582 ( .A(\mem[0][20] ), .B(\mem[1][20] ), .S(n545), .Z(n519) );
  MUX2_X1 U583 ( .A(n519), .B(n518), .S(N11), .Z(n520) );
  MUX2_X1 U584 ( .A(n520), .B(n517), .S(n539), .Z(N16) );
  MUX2_X1 U585 ( .A(\mem[6][21] ), .B(\mem[7][21] ), .S(n544), .Z(n521) );
  MUX2_X1 U586 ( .A(\mem[4][21] ), .B(\mem[5][21] ), .S(n543), .Z(n522) );
  MUX2_X1 U587 ( .A(n522), .B(n521), .S(N11), .Z(n523) );
  MUX2_X1 U588 ( .A(\mem[2][21] ), .B(\mem[3][21] ), .S(n542), .Z(n524) );
  MUX2_X1 U589 ( .A(\mem[0][21] ), .B(\mem[1][21] ), .S(n542), .Z(n525) );
  MUX2_X1 U590 ( .A(n525), .B(n524), .S(N11), .Z(n526) );
  MUX2_X1 U591 ( .A(n526), .B(n523), .S(n539), .Z(N15) );
  MUX2_X1 U592 ( .A(\mem[6][22] ), .B(\mem[7][22] ), .S(n542), .Z(n527) );
  MUX2_X1 U593 ( .A(\mem[4][22] ), .B(\mem[5][22] ), .S(n544), .Z(n528) );
  MUX2_X1 U594 ( .A(n528), .B(n527), .S(N11), .Z(n529) );
  MUX2_X1 U595 ( .A(\mem[2][22] ), .B(\mem[3][22] ), .S(n543), .Z(n530) );
  MUX2_X1 U596 ( .A(\mem[0][22] ), .B(\mem[1][22] ), .S(n543), .Z(n531) );
  MUX2_X1 U597 ( .A(n531), .B(n530), .S(N11), .Z(n532) );
  MUX2_X1 U598 ( .A(n532), .B(n529), .S(n539), .Z(N14) );
  MUX2_X1 U599 ( .A(\mem[6][23] ), .B(\mem[7][23] ), .S(n545), .Z(n533) );
  MUX2_X1 U600 ( .A(\mem[4][23] ), .B(\mem[5][23] ), .S(n545), .Z(n534) );
  MUX2_X1 U601 ( .A(n534), .B(n533), .S(N11), .Z(n535) );
  MUX2_X1 U602 ( .A(\mem[2][23] ), .B(\mem[3][23] ), .S(n545), .Z(n536) );
  MUX2_X1 U603 ( .A(\mem[0][23] ), .B(\mem[1][23] ), .S(n545), .Z(n537) );
  MUX2_X1 U604 ( .A(n537), .B(n536), .S(N11), .Z(n538) );
  MUX2_X1 U605 ( .A(n538), .B(n535), .S(N12), .Z(N13) );
  CLKBUF_X1 U606 ( .A(N10), .Z(n545) );
endmodule


module datapath_DW_mult_tc_16 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n1, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n34, n36, n37, n38, n39, n40, n41, n42, n43, n45, n47, n48, n49, n52,
         n54, n55, n56, n57, n58, n59, n61, n63, n64, n66, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n112,
         n114, n115, n117, n119, n120, n121, n123, n125, n126, n127, n128,
         n129, n131, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n143, n145, n146, n148, n149, n150, n156, n157, n158, n160, n161,
         n165, n167, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n284, n285, n286, n287, n288, n290, n291,
         n293, n294, n296, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n467, n468, n469, n470, n471, n472, n479, n480,
         n481, n482, n483, n484, n485, n487, n488, n489, n490, n491, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594;

  FA_X1 U4 ( .A(n305), .B(n171), .CI(n149), .CO(n24), .S(product[22]) );
  FA_X1 U194 ( .A(n306), .B(n177), .CI(n313), .CO(n173), .S(n174) );
  FA_X1 U195 ( .A(n178), .B(n314), .CI(n181), .CO(n175), .S(n176) );
  FA_X1 U197 ( .A(n185), .B(n326), .CI(n182), .CO(n179), .S(n180) );
  FA_X1 U198 ( .A(n307), .B(n187), .CI(n315), .CO(n181), .S(n182) );
  FA_X1 U199 ( .A(n186), .B(n193), .CI(n191), .CO(n183), .S(n184) );
  FA_X1 U200 ( .A(n327), .B(n316), .CI(n188), .CO(n185), .S(n186) );
  FA_X1 U202 ( .A(n197), .B(n194), .CI(n192), .CO(n189), .S(n190) );
  FA_X1 U203 ( .A(n317), .B(n308), .CI(n199), .CO(n191), .S(n192) );
  FA_X1 U204 ( .A(n328), .B(n201), .CI(n339), .CO(n193), .S(n194) );
  FA_X1 U205 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U206 ( .A(n209), .B(n202), .CI(n207), .CO(n197), .S(n198) );
  FA_X1 U207 ( .A(n329), .B(n340), .CI(n318), .CO(n199), .S(n200) );
  FA_X1 U209 ( .A(n213), .B(n208), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U210 ( .A(n215), .B(n217), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U211 ( .A(n341), .B(n309), .CI(n352), .CO(n207), .S(n208) );
  FA_X1 U212 ( .A(n319), .B(n330), .CI(n219), .CO(n209), .S(n210) );
  FA_X1 U213 ( .A(n223), .B(n216), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U214 ( .A(n218), .B(n227), .CI(n225), .CO(n213), .S(n214) );
  FA_X1 U215 ( .A(n220), .B(n320), .CI(n229), .CO(n215), .S(n216) );
  FA_X1 U216 ( .A(n331), .B(n342), .CI(n353), .CO(n217), .S(n218) );
  FA_X1 U218 ( .A(n233), .B(n226), .CI(n224), .CO(n221), .S(n222) );
  FA_X1 U219 ( .A(n228), .B(n237), .CI(n235), .CO(n223), .S(n224) );
  FA_X1 U220 ( .A(n239), .B(n365), .CI(n230), .CO(n225), .S(n226) );
  FA_X1 U221 ( .A(n332), .B(n354), .CI(n321), .CO(n227), .S(n228) );
  FA_X1 U224 ( .A(n243), .B(n236), .CI(n234), .CO(n231), .S(n232) );
  FA_X1 U225 ( .A(n245), .B(n247), .CI(n238), .CO(n233), .S(n234) );
  FA_X1 U226 ( .A(n333), .B(n322), .CI(n240), .CO(n235), .S(n236) );
  FA_X1 U227 ( .A(n366), .B(n344), .CI(n355), .CO(n237), .S(n238) );
  HA_X1 U228 ( .A(n311), .B(n299), .CO(n239), .S(n240) );
  FA_X1 U229 ( .A(n251), .B(n246), .CI(n244), .CO(n241), .S(n242) );
  FA_X1 U230 ( .A(n253), .B(n255), .CI(n248), .CO(n243), .S(n244) );
  FA_X1 U231 ( .A(n334), .B(n356), .CI(n367), .CO(n245), .S(n246) );
  FA_X1 U232 ( .A(n323), .B(n312), .CI(n345), .CO(n247), .S(n248) );
  FA_X1 U235 ( .A(n335), .B(n324), .CI(n368), .CO(n253), .S(n254) );
  HA_X1 U236 ( .A(n346), .B(n300), .CO(n255), .S(n256) );
  FA_X1 U237 ( .A(n262), .B(n265), .CI(n260), .CO(n257), .S(n258) );
  FA_X1 U238 ( .A(n369), .B(n336), .CI(n267), .CO(n259), .S(n260) );
  FA_X1 U239 ( .A(n347), .B(n325), .CI(n358), .CO(n261), .S(n262) );
  FA_X1 U240 ( .A(n271), .B(n268), .CI(n266), .CO(n263), .S(n264) );
  FA_X1 U241 ( .A(n337), .B(n359), .CI(n370), .CO(n265), .S(n266) );
  HA_X1 U242 ( .A(n301), .B(n348), .CO(n267), .S(n268) );
  FA_X1 U243 ( .A(n275), .B(n371), .CI(n272), .CO(n269), .S(n270) );
  FA_X1 U244 ( .A(n349), .B(n338), .CI(n360), .CO(n271), .S(n272) );
  FA_X1 U245 ( .A(n372), .B(n361), .CI(n276), .CO(n273), .S(n274) );
  HA_X1 U246 ( .A(n350), .B(n302), .CO(n275), .S(n276) );
  FA_X1 U247 ( .A(n362), .B(n351), .CI(n373), .CO(n277), .S(n278) );
  HA_X1 U248 ( .A(n363), .B(n303), .CO(n279), .S(n280) );
  CLKBUF_X1 U484 ( .A(b[6]), .Z(n460) );
  BUF_X1 U485 ( .A(a[9]), .Z(n594) );
  BUF_X1 U486 ( .A(b[5]), .Z(n461) );
  BUF_X2 U487 ( .A(a[7]), .Z(n493) );
  BUF_X2 U488 ( .A(n504), .Z(n480) );
  AOI21_X1 U489 ( .B1(n66), .B2(n581), .A(n61), .ZN(n59) );
  AND2_X1 U490 ( .A1(n588), .A2(n148), .ZN(product[1]) );
  BUF_X2 U491 ( .A(a[11]), .Z(n491) );
  CLKBUF_X1 U492 ( .A(n41), .Z(n561) );
  CLKBUF_X1 U493 ( .A(n69), .Z(n562) );
  BUF_X1 U494 ( .A(b[7]), .Z(n459) );
  CLKBUF_X1 U495 ( .A(n497), .Z(n563) );
  NAND2_X1 U496 ( .A1(n467), .A2(n503), .ZN(n497) );
  BUF_X1 U497 ( .A(b[9]), .Z(n457) );
  AOI21_X1 U498 ( .B1(n100), .B2(n108), .A(n101), .ZN(n564) );
  XNOR2_X1 U499 ( .A(n565), .B(n261), .ZN(n252) );
  XNOR2_X1 U500 ( .A(n256), .B(n357), .ZN(n565) );
  AOI21_X1 U501 ( .B1(n578), .B2(n56), .A(n57), .ZN(n566) );
  BUF_X4 U502 ( .A(n503), .Z(n479) );
  NOR2_X2 U503 ( .A1(n232), .A2(n241), .ZN(n102) );
  CLKBUF_X1 U504 ( .A(b[4]), .Z(n462) );
  AOI21_X1 U505 ( .B1(n561), .B2(n584), .A(n34), .ZN(n567) );
  NOR2_X2 U506 ( .A1(n212), .A2(n221), .ZN(n91) );
  BUF_X1 U507 ( .A(b[8]), .Z(n458) );
  XOR2_X1 U508 ( .A(n254), .B(n259), .Z(n568) );
  XOR2_X1 U509 ( .A(n568), .B(n252), .Z(n250) );
  NAND2_X1 U510 ( .A1(n256), .A2(n357), .ZN(n569) );
  NAND2_X1 U511 ( .A1(n256), .A2(n261), .ZN(n570) );
  NAND2_X1 U512 ( .A1(n357), .A2(n261), .ZN(n571) );
  NAND3_X1 U513 ( .A1(n569), .A2(n570), .A3(n571), .ZN(n251) );
  NAND2_X1 U514 ( .A1(n254), .A2(n259), .ZN(n572) );
  NAND2_X1 U515 ( .A1(n254), .A2(n252), .ZN(n573) );
  NAND2_X1 U516 ( .A1(n259), .A2(n252), .ZN(n574) );
  NAND3_X1 U517 ( .A1(n572), .A2(n573), .A3(n574), .ZN(n249) );
  CLKBUF_X3 U518 ( .A(n506), .Z(n482) );
  BUF_X2 U519 ( .A(b[3]), .Z(n463) );
  OR2_X1 U520 ( .A1(n280), .A2(n374), .ZN(n575) );
  CLKBUF_X1 U521 ( .A(b[0]), .Z(n576) );
  AOI21_X1 U522 ( .B1(n100), .B2(n108), .A(n101), .ZN(n99) );
  AOI21_X1 U523 ( .B1(n590), .B2(n134), .A(n131), .ZN(n577) );
  OAI21_X1 U524 ( .B1(n564), .B2(n71), .A(n72), .ZN(n578) );
  XNOR2_X1 U525 ( .A(n69), .B(n579), .ZN(product[16]) );
  AND2_X1 U526 ( .A1(n582), .A2(n68), .ZN(n579) );
  OR2_X1 U527 ( .A1(n258), .A2(n263), .ZN(n580) );
  OR2_X1 U528 ( .A1(n184), .A2(n189), .ZN(n581) );
  OR2_X1 U529 ( .A1(n190), .A2(n195), .ZN(n582) );
  OR2_X1 U530 ( .A1(n250), .A2(n257), .ZN(n583) );
  OR2_X1 U531 ( .A1(n175), .A2(n174), .ZN(n584) );
  OR2_X1 U532 ( .A1(n176), .A2(n179), .ZN(n585) );
  OR2_X1 U533 ( .A1(n180), .A2(n183), .ZN(n586) );
  OR2_X1 U534 ( .A1(n375), .A2(n364), .ZN(n587) );
  OR2_X1 U535 ( .A1(n376), .A2(n304), .ZN(n588) );
  OR2_X1 U536 ( .A1(n264), .A2(n269), .ZN(n589) );
  OR2_X1 U537 ( .A1(n274), .A2(n277), .ZN(n590) );
  BUF_X2 U538 ( .A(n507), .Z(n483) );
  BUF_X1 U539 ( .A(a[9]), .Z(n593) );
  CLKBUF_X3 U540 ( .A(a[3]), .Z(n495) );
  CLKBUF_X3 U541 ( .A(a[1]), .Z(n496) );
  INV_X1 U542 ( .A(n281), .ZN(n305) );
  NAND2_X1 U543 ( .A1(n150), .A2(n29), .ZN(n3) );
  NOR2_X1 U544 ( .A1(n173), .A2(n172), .ZN(n28) );
  INV_X1 U545 ( .A(n28), .ZN(n150) );
  NAND2_X1 U546 ( .A1(n173), .A2(n172), .ZN(n29) );
  INV_X1 U547 ( .A(n287), .ZN(n326) );
  NAND2_X1 U548 ( .A1(n584), .A2(n36), .ZN(n4) );
  INV_X1 U549 ( .A(n36), .ZN(n34) );
  NAND2_X1 U550 ( .A1(n175), .A2(n174), .ZN(n36) );
  INV_X1 U551 ( .A(n171), .ZN(n172) );
  NAND2_X1 U552 ( .A1(n585), .A2(n47), .ZN(n5) );
  BUF_X2 U553 ( .A(n508), .Z(n484) );
  NAND2_X1 U554 ( .A1(n176), .A2(n179), .ZN(n47) );
  INV_X1 U555 ( .A(n586), .ZN(n49) );
  NAND2_X1 U556 ( .A1(n586), .A2(n54), .ZN(n6) );
  INV_X1 U557 ( .A(n157), .ZN(n80) );
  INV_X1 U558 ( .A(n290), .ZN(n339) );
  INV_X1 U559 ( .A(n47), .ZN(n45) );
  NAND2_X2 U560 ( .A1(n469), .A2(n505), .ZN(n499) );
  NOR2_X1 U561 ( .A1(n58), .A2(n42), .ZN(n40) );
  NAND2_X1 U562 ( .A1(n180), .A2(n183), .ZN(n54) );
  NAND2_X1 U563 ( .A1(n375), .A2(n364), .ZN(n145) );
  CLKBUF_X3 U564 ( .A(a[5]), .Z(n494) );
  NAND2_X2 U565 ( .A1(n472), .A2(n508), .ZN(n502) );
  NOR2_X1 U566 ( .A1(n196), .A2(n203), .ZN(n75) );
  INV_X1 U567 ( .A(n40), .ZN(n38) );
  NAND2_X1 U568 ( .A1(n161), .A2(n106), .ZN(n14) );
  INV_X1 U569 ( .A(n54), .ZN(n52) );
  NOR2_X1 U570 ( .A1(n280), .A2(n374), .ZN(n139) );
  INV_X1 U571 ( .A(n135), .ZN(n167) );
  NOR2_X1 U572 ( .A1(n278), .A2(n279), .ZN(n135) );
  INV_X1 U573 ( .A(n58), .ZN(n56) );
  NOR2_X1 U574 ( .A1(n222), .A2(n231), .ZN(n96) );
  NAND2_X1 U575 ( .A1(n278), .A2(n279), .ZN(n136) );
  XNOR2_X1 U576 ( .A(n496), .B(n461), .ZN(n448) );
  XNOR2_X1 U577 ( .A(n496), .B(n460), .ZN(n447) );
  OAI21_X1 U578 ( .B1(n564), .B2(n71), .A(n72), .ZN(n70) );
  INV_X1 U579 ( .A(n88), .ZN(n86) );
  NAND2_X1 U580 ( .A1(n582), .A2(n581), .ZN(n58) );
  INV_X1 U581 ( .A(n87), .ZN(n85) );
  NOR2_X1 U582 ( .A1(n87), .A2(n80), .ZN(n78) );
  INV_X1 U583 ( .A(n89), .ZN(n87) );
  XNOR2_X1 U584 ( .A(n495), .B(n460), .ZN(n434) );
  XNOR2_X1 U585 ( .A(n495), .B(n461), .ZN(n435) );
  INV_X1 U586 ( .A(n145), .ZN(n143) );
  INV_X1 U587 ( .A(n102), .ZN(n160) );
  NAND2_X1 U588 ( .A1(n580), .A2(n119), .ZN(n16) );
  INV_X1 U589 ( .A(n119), .ZN(n117) );
  AOI21_X1 U590 ( .B1(n499), .B2(n481), .A(n403), .ZN(n287) );
  OAI22_X1 U591 ( .A1(n499), .A2(n410), .B1(n409), .B2(n481), .ZN(n333) );
  OAI22_X1 U592 ( .A1(n499), .A2(n405), .B1(n404), .B2(n481), .ZN(n328) );
  OAI22_X1 U593 ( .A1(n499), .A2(n413), .B1(n412), .B2(n481), .ZN(n336) );
  INV_X1 U594 ( .A(n481), .ZN(n288) );
  OAI22_X1 U595 ( .A1(n499), .A2(n404), .B1(n403), .B2(n481), .ZN(n327) );
  OAI22_X1 U596 ( .A1(n499), .A2(n407), .B1(n406), .B2(n481), .ZN(n330) );
  OAI22_X1 U597 ( .A1(n499), .A2(n408), .B1(n407), .B2(n481), .ZN(n331) );
  OAI22_X1 U598 ( .A1(n499), .A2(n409), .B1(n408), .B2(n481), .ZN(n332) );
  OAI22_X1 U599 ( .A1(n499), .A2(n406), .B1(n405), .B2(n481), .ZN(n329) );
  NAND2_X1 U600 ( .A1(n583), .A2(n114), .ZN(n15) );
  INV_X1 U601 ( .A(n82), .ZN(n157) );
  NAND2_X1 U602 ( .A1(n270), .A2(n273), .ZN(n128) );
  NAND2_X1 U603 ( .A1(n258), .A2(n263), .ZN(n119) );
  AOI21_X1 U604 ( .B1(n587), .B2(n146), .A(n143), .ZN(n141) );
  CLKBUF_X3 U605 ( .A(n505), .Z(n481) );
  NAND2_X1 U606 ( .A1(n250), .A2(n257), .ZN(n114) );
  INV_X1 U607 ( .A(n133), .ZN(n131) );
  INV_X1 U608 ( .A(n482), .ZN(n291) );
  INV_X1 U609 ( .A(n75), .ZN(n156) );
  NAND2_X1 U610 ( .A1(n156), .A2(n76), .ZN(n9) );
  INV_X1 U611 ( .A(n125), .ZN(n123) );
  NAND2_X1 U612 ( .A1(n280), .A2(n374), .ZN(n140) );
  NAND2_X1 U613 ( .A1(n196), .A2(n203), .ZN(n76) );
  NAND2_X1 U614 ( .A1(n274), .A2(n277), .ZN(n133) );
  NAND2_X1 U615 ( .A1(n264), .A2(n269), .ZN(n125) );
  INV_X1 U616 ( .A(n293), .ZN(n352) );
  INV_X1 U617 ( .A(n91), .ZN(n158) );
  NOR2_X1 U618 ( .A1(n91), .A2(n96), .ZN(n89) );
  NAND2_X1 U619 ( .A1(n158), .A2(n92), .ZN(n11) );
  INV_X1 U620 ( .A(n127), .ZN(n165) );
  NOR2_X1 U621 ( .A1(n270), .A2(n273), .ZN(n127) );
  OAI22_X1 U622 ( .A1(n499), .A2(n414), .B1(n413), .B2(n481), .ZN(n337) );
  INV_X1 U623 ( .A(n284), .ZN(n313) );
  INV_X1 U624 ( .A(n114), .ZN(n112) );
  NAND2_X1 U625 ( .A1(n212), .A2(n221), .ZN(n92) );
  INV_X1 U626 ( .A(n105), .ZN(n161) );
  NOR2_X1 U627 ( .A1(n242), .A2(n249), .ZN(n105) );
  XNOR2_X1 U628 ( .A(a[7]), .B(a[8]), .ZN(n504) );
  XNOR2_X1 U629 ( .A(n496), .B(n463), .ZN(n450) );
  XNOR2_X1 U630 ( .A(n463), .B(n495), .ZN(n437) );
  XNOR2_X1 U631 ( .A(n463), .B(n494), .ZN(n424) );
  XNOR2_X1 U632 ( .A(n496), .B(n457), .ZN(n444) );
  XNOR2_X1 U633 ( .A(n494), .B(n457), .ZN(n418) );
  XNOR2_X1 U634 ( .A(n593), .B(n457), .ZN(n392) );
  XNOR2_X1 U635 ( .A(n496), .B(n462), .ZN(n449) );
  XNOR2_X1 U636 ( .A(n462), .B(n495), .ZN(n436) );
  XNOR2_X1 U637 ( .A(n462), .B(n494), .ZN(n423) );
  XNOR2_X1 U638 ( .A(n462), .B(n593), .ZN(n397) );
  NAND2_X1 U639 ( .A1(n242), .A2(n249), .ZN(n106) );
  XNOR2_X1 U640 ( .A(n494), .B(n461), .ZN(n422) );
  INV_X1 U641 ( .A(n296), .ZN(n365) );
  XNOR2_X1 U642 ( .A(n594), .B(n461), .ZN(n396) );
  XNOR2_X1 U643 ( .A(n594), .B(n460), .ZN(n395) );
  BUF_X1 U644 ( .A(n498), .Z(n591) );
  BUF_X1 U645 ( .A(n498), .Z(n592) );
  NAND2_X1 U646 ( .A1(n468), .A2(n504), .ZN(n498) );
  XNOR2_X1 U647 ( .A(n310), .B(n343), .ZN(n230) );
  INV_X1 U648 ( .A(n483), .ZN(n294) );
  NOR2_X1 U649 ( .A1(n82), .A2(n75), .ZN(n73) );
  NAND2_X1 U650 ( .A1(n157), .A2(n83), .ZN(n10) );
  OAI21_X1 U651 ( .B1(n88), .B2(n80), .A(n83), .ZN(n79) );
  NOR2_X1 U652 ( .A1(n204), .A2(n211), .ZN(n82) );
  XNOR2_X1 U653 ( .A(n496), .B(b[2]), .ZN(n451) );
  XNOR2_X1 U654 ( .A(n495), .B(b[2]), .ZN(n438) );
  XNOR2_X1 U655 ( .A(n494), .B(b[2]), .ZN(n425) );
  INV_X1 U656 ( .A(n96), .ZN(n94) );
  NAND2_X1 U657 ( .A1(n94), .A2(n97), .ZN(n12) );
  OAI21_X1 U658 ( .B1(n91), .B2(n97), .A(n92), .ZN(n90) );
  INV_X1 U659 ( .A(n97), .ZN(n95) );
  NAND2_X1 U660 ( .A1(n89), .A2(n73), .ZN(n71) );
  INV_X1 U661 ( .A(n90), .ZN(n88) );
  NAND2_X1 U662 ( .A1(n204), .A2(n211), .ZN(n83) );
  NAND2_X1 U663 ( .A1(n222), .A2(n231), .ZN(n97) );
  OAI21_X1 U664 ( .B1(n102), .B2(n106), .A(n103), .ZN(n101) );
  NOR2_X1 U665 ( .A1(n102), .A2(n105), .ZN(n100) );
  NAND2_X1 U666 ( .A1(n160), .A2(n103), .ZN(n13) );
  OAI22_X1 U667 ( .A1(n502), .A2(n448), .B1(n447), .B2(n484), .ZN(n371) );
  OAI22_X1 U668 ( .A1(n502), .A2(n451), .B1(n450), .B2(n484), .ZN(n374) );
  OAI22_X1 U669 ( .A1(n502), .A2(n449), .B1(n448), .B2(n484), .ZN(n372) );
  OAI22_X1 U670 ( .A1(n502), .A2(n450), .B1(n449), .B2(n484), .ZN(n373) );
  OAI22_X1 U671 ( .A1(n502), .A2(n490), .B1(n454), .B2(n484), .ZN(n304) );
  OAI22_X1 U672 ( .A1(n502), .A2(n453), .B1(n452), .B2(n484), .ZN(n376) );
  OAI22_X1 U673 ( .A1(n502), .A2(n446), .B1(n445), .B2(n484), .ZN(n369) );
  OAI22_X1 U674 ( .A1(n502), .A2(n447), .B1(n446), .B2(n484), .ZN(n370) );
  OAI22_X1 U675 ( .A1(n502), .A2(n452), .B1(n451), .B2(n484), .ZN(n375) );
  OAI22_X1 U676 ( .A1(n502), .A2(n445), .B1(n444), .B2(n484), .ZN(n368) );
  OAI22_X1 U677 ( .A1(n502), .A2(n444), .B1(n443), .B2(n484), .ZN(n367) );
  AOI21_X1 U678 ( .B1(n502), .B2(n484), .A(n442), .ZN(n296) );
  OR2_X1 U679 ( .A1(n310), .A2(n343), .ZN(n229) );
  NAND2_X2 U680 ( .A1(n470), .A2(n506), .ZN(n500) );
  NAND2_X2 U681 ( .A1(n471), .A2(n507), .ZN(n501) );
  XNOR2_X1 U682 ( .A(n496), .B(n456), .ZN(n443) );
  XNOR2_X1 U683 ( .A(n495), .B(n456), .ZN(n430) );
  XNOR2_X1 U684 ( .A(n494), .B(n456), .ZN(n417) );
  XNOR2_X1 U685 ( .A(n594), .B(n456), .ZN(n391) );
  BUF_X2 U686 ( .A(b[10]), .Z(n456) );
  AOI21_X1 U687 ( .B1(n591), .B2(n480), .A(n390), .ZN(n284) );
  OAI22_X1 U688 ( .A1(n498), .A2(n391), .B1(n480), .B2(n390), .ZN(n314) );
  OAI22_X1 U689 ( .A1(n592), .A2(n394), .B1(n480), .B2(n393), .ZN(n317) );
  OAI22_X1 U690 ( .A1(n591), .A2(n393), .B1(n480), .B2(n392), .ZN(n316) );
  OAI22_X1 U691 ( .A1(n591), .A2(n392), .B1(n480), .B2(n391), .ZN(n315) );
  OAI22_X1 U692 ( .A1(n592), .A2(n395), .B1(n480), .B2(n394), .ZN(n318) );
  OAI22_X1 U693 ( .A1(n591), .A2(n397), .B1(n480), .B2(n396), .ZN(n320) );
  OAI22_X1 U694 ( .A1(n591), .A2(n286), .B1(n402), .B2(n480), .ZN(n300) );
  OAI22_X1 U695 ( .A1(n592), .A2(n396), .B1(n480), .B2(n395), .ZN(n319) );
  INV_X1 U696 ( .A(n480), .ZN(n285) );
  OAI22_X1 U697 ( .A1(n592), .A2(n401), .B1(n480), .B2(n400), .ZN(n324) );
  XNOR2_X1 U698 ( .A(n496), .B(b[1]), .ZN(n452) );
  XNOR2_X1 U699 ( .A(n495), .B(b[1]), .ZN(n439) );
  XNOR2_X1 U700 ( .A(n494), .B(b[1]), .ZN(n426) );
  OAI22_X1 U701 ( .A1(n499), .A2(n412), .B1(n411), .B2(n481), .ZN(n335) );
  OAI22_X1 U702 ( .A1(n499), .A2(n411), .B1(n410), .B2(n481), .ZN(n334) );
  OAI22_X1 U703 ( .A1(n501), .A2(n438), .B1(n437), .B2(n483), .ZN(n361) );
  OAI22_X1 U704 ( .A1(n501), .A2(n434), .B1(n483), .B2(n433), .ZN(n357) );
  OAI22_X1 U705 ( .A1(n501), .A2(n439), .B1(n483), .B2(n438), .ZN(n362) );
  OAI22_X1 U706 ( .A1(n501), .A2(n437), .B1(n436), .B2(n483), .ZN(n360) );
  OAI22_X1 U707 ( .A1(n501), .A2(n436), .B1(n483), .B2(n435), .ZN(n359) );
  OAI22_X1 U708 ( .A1(n501), .A2(n440), .B1(n483), .B2(n439), .ZN(n363) );
  OAI22_X1 U709 ( .A1(n501), .A2(n435), .B1(n483), .B2(n434), .ZN(n358) );
  AOI21_X1 U710 ( .B1(n501), .B2(n483), .A(n429), .ZN(n293) );
  OAI22_X1 U711 ( .A1(n501), .A2(n430), .B1(n429), .B2(n483), .ZN(n353) );
  OAI22_X1 U712 ( .A1(n501), .A2(n433), .B1(n483), .B2(n432), .ZN(n356) );
  XNOR2_X1 U713 ( .A(a[5]), .B(a[6]), .ZN(n505) );
  XNOR2_X1 U714 ( .A(n496), .B(n455), .ZN(n442) );
  XNOR2_X1 U715 ( .A(n495), .B(n455), .ZN(n429) );
  XNOR2_X1 U716 ( .A(n494), .B(n455), .ZN(n416) );
  XNOR2_X1 U717 ( .A(n593), .B(n455), .ZN(n390) );
  BUF_X2 U718 ( .A(b[11]), .Z(n455) );
  OAI22_X1 U719 ( .A1(n592), .A2(n399), .B1(n398), .B2(n480), .ZN(n322) );
  OAI22_X1 U720 ( .A1(n592), .A2(n398), .B1(n397), .B2(n480), .ZN(n321) );
  XNOR2_X1 U721 ( .A(n463), .B(n594), .ZN(n398) );
  XNOR2_X1 U722 ( .A(n593), .B(b[2]), .ZN(n399) );
  AOI21_X1 U723 ( .B1(n500), .B2(n482), .A(n416), .ZN(n290) );
  OAI22_X1 U724 ( .A1(n500), .A2(n426), .B1(n482), .B2(n425), .ZN(n349) );
  OAI22_X1 U725 ( .A1(n500), .A2(n417), .B1(n482), .B2(n416), .ZN(n340) );
  OAI22_X1 U726 ( .A1(n500), .A2(n418), .B1(n482), .B2(n417), .ZN(n341) );
  OAI22_X1 U727 ( .A1(n500), .A2(n425), .B1(n424), .B2(n482), .ZN(n348) );
  OAI22_X1 U728 ( .A1(n500), .A2(n427), .B1(n482), .B2(n426), .ZN(n350) );
  OAI22_X1 U729 ( .A1(n500), .A2(n423), .B1(n482), .B2(n422), .ZN(n346) );
  OAI22_X1 U730 ( .A1(n500), .A2(n424), .B1(n423), .B2(n482), .ZN(n347) );
  OAI22_X1 U731 ( .A1(n500), .A2(n419), .B1(n482), .B2(n418), .ZN(n342) );
  OAI22_X1 U732 ( .A1(n500), .A2(n422), .B1(n482), .B2(n421), .ZN(n345) );
  OAI22_X1 U733 ( .A1(n500), .A2(n420), .B1(n482), .B2(n419), .ZN(n343) );
  XOR2_X1 U734 ( .A(a[1]), .B(a[0]), .Z(n472) );
  BUF_X1 U735 ( .A(b[0]), .Z(n1) );
  OAI22_X1 U736 ( .A1(n502), .A2(n443), .B1(n442), .B2(n484), .ZN(n366) );
  XNOR2_X1 U737 ( .A(n493), .B(n456), .ZN(n404) );
  XNOR2_X1 U738 ( .A(n493), .B(n455), .ZN(n403) );
  XNOR2_X1 U739 ( .A(n493), .B(n457), .ZN(n405) );
  XNOR2_X1 U740 ( .A(n493), .B(b[1]), .ZN(n413) );
  XNOR2_X1 U741 ( .A(n493), .B(b[2]), .ZN(n412) );
  XNOR2_X1 U742 ( .A(n493), .B(n461), .ZN(n409) );
  XNOR2_X1 U743 ( .A(n493), .B(n460), .ZN(n408) );
  XNOR2_X1 U744 ( .A(n462), .B(n493), .ZN(n410) );
  XNOR2_X1 U745 ( .A(n463), .B(n493), .ZN(n411) );
  XNOR2_X1 U746 ( .A(a[3]), .B(a[4]), .ZN(n506) );
  OAI22_X1 U747 ( .A1(n498), .A2(n400), .B1(n480), .B2(n399), .ZN(n323) );
  XNOR2_X1 U748 ( .A(n594), .B(b[1]), .ZN(n400) );
  OAI22_X1 U749 ( .A1(n500), .A2(n421), .B1(n482), .B2(n420), .ZN(n344) );
  XNOR2_X1 U750 ( .A(n494), .B(n460), .ZN(n421) );
  XNOR2_X1 U751 ( .A(a[1]), .B(a[2]), .ZN(n507) );
  OAI22_X1 U752 ( .A1(n501), .A2(n432), .B1(n483), .B2(n431), .ZN(n355) );
  OAI22_X1 U753 ( .A1(n501), .A2(n431), .B1(n483), .B2(n430), .ZN(n354) );
  XNOR2_X1 U754 ( .A(n495), .B(n457), .ZN(n431) );
  XNOR2_X1 U755 ( .A(n496), .B(n458), .ZN(n445) );
  XNOR2_X1 U756 ( .A(n495), .B(n458), .ZN(n432) );
  XNOR2_X1 U757 ( .A(n494), .B(n458), .ZN(n419) );
  XNOR2_X1 U758 ( .A(n493), .B(n458), .ZN(n406) );
  XNOR2_X1 U759 ( .A(n594), .B(n458), .ZN(n393) );
  INV_X1 U760 ( .A(n479), .ZN(n282) );
  AND2_X1 U761 ( .A1(n1), .A2(n291), .ZN(n351) );
  AND2_X1 U762 ( .A1(n1), .A2(n288), .ZN(n338) );
  AND2_X1 U763 ( .A1(n576), .A2(n294), .ZN(n364) );
  XNOR2_X1 U764 ( .A(n1), .B(n496), .ZN(n453) );
  OR2_X1 U765 ( .A1(n1), .A2(n490), .ZN(n454) );
  AND2_X1 U766 ( .A1(n1), .A2(n285), .ZN(n325) );
  XNOR2_X1 U767 ( .A(n576), .B(n493), .ZN(n414) );
  XNOR2_X1 U768 ( .A(n1), .B(n495), .ZN(n440) );
  OR2_X1 U769 ( .A1(n1), .A2(n487), .ZN(n415) );
  OR2_X1 U770 ( .A1(n1), .A2(n489), .ZN(n441) );
  XNOR2_X1 U771 ( .A(n1), .B(n494), .ZN(n427) );
  OR2_X1 U772 ( .A1(n1), .A2(n488), .ZN(n428) );
  AND2_X1 U773 ( .A1(n1), .A2(n282), .ZN(n312) );
  OR2_X1 U774 ( .A1(n1), .A2(n286), .ZN(n402) );
  XNOR2_X1 U775 ( .A(n576), .B(n593), .ZN(n401) );
  OR2_X1 U776 ( .A1(b[0]), .A2(n485), .ZN(n389) );
  INV_X1 U777 ( .A(n177), .ZN(n178) );
  XOR2_X1 U778 ( .A(a[7]), .B(a[6]), .Z(n469) );
  XOR2_X1 U779 ( .A(a[9]), .B(a[8]), .Z(n468) );
  XOR2_X1 U780 ( .A(a[3]), .B(a[2]), .Z(n471) );
  OAI22_X1 U781 ( .A1(n497), .A2(n382), .B1(n479), .B2(n381), .ZN(n187) );
  INV_X1 U782 ( .A(n187), .ZN(n188) );
  XOR2_X1 U783 ( .A(a[5]), .B(a[4]), .Z(n470) );
  OAI22_X1 U784 ( .A1(n497), .A2(n384), .B1(n479), .B2(n383), .ZN(n201) );
  INV_X1 U785 ( .A(n201), .ZN(n202) );
  NAND2_X1 U786 ( .A1(n232), .A2(n241), .ZN(n103) );
  NAND2_X1 U787 ( .A1(n581), .A2(n63), .ZN(n7) );
  INV_X1 U788 ( .A(n63), .ZN(n61) );
  NAND2_X1 U789 ( .A1(n184), .A2(n189), .ZN(n63) );
  INV_X1 U790 ( .A(a[9]), .ZN(n286) );
  OAI22_X1 U791 ( .A1(n497), .A2(n485), .B1(n389), .B2(n479), .ZN(n299) );
  OAI22_X1 U792 ( .A1(n497), .A2(n387), .B1(n479), .B2(n386), .ZN(n310) );
  OAI22_X1 U793 ( .A1(n497), .A2(n386), .B1(n385), .B2(n479), .ZN(n219) );
  OAI22_X1 U794 ( .A1(n563), .A2(n381), .B1(n479), .B2(n380), .ZN(n307) );
  OAI22_X1 U795 ( .A1(n563), .A2(n378), .B1(n479), .B2(n377), .ZN(n171) );
  AOI21_X1 U796 ( .B1(n563), .B2(n479), .A(n377), .ZN(n281) );
  OAI22_X1 U797 ( .A1(n563), .A2(n379), .B1(n479), .B2(n378), .ZN(n306) );
  OAI22_X1 U798 ( .A1(n563), .A2(n383), .B1(n479), .B2(n382), .ZN(n308) );
  OAI22_X1 U799 ( .A1(n497), .A2(n385), .B1(n384), .B2(n479), .ZN(n309) );
  OAI22_X1 U800 ( .A1(n563), .A2(n380), .B1(n479), .B2(n379), .ZN(n177) );
  OAI22_X1 U801 ( .A1(n497), .A2(n388), .B1(n479), .B2(n387), .ZN(n311) );
  INV_X1 U802 ( .A(n496), .ZN(n490) );
  XNOR2_X1 U803 ( .A(n496), .B(n459), .ZN(n446) );
  XNOR2_X1 U804 ( .A(n495), .B(n459), .ZN(n433) );
  XNOR2_X1 U805 ( .A(n494), .B(n459), .ZN(n420) );
  XNOR2_X1 U806 ( .A(n493), .B(n459), .ZN(n407) );
  XNOR2_X1 U807 ( .A(n593), .B(n459), .ZN(n394) );
  NAND2_X1 U808 ( .A1(n586), .A2(n585), .ZN(n42) );
  AOI21_X1 U809 ( .B1(n41), .B2(n584), .A(n34), .ZN(n32) );
  AOI21_X1 U810 ( .B1(n90), .B2(n73), .A(n74), .ZN(n72) );
  OAI21_X1 U811 ( .B1(n83), .B2(n75), .A(n76), .ZN(n74) );
  XOR2_X1 U812 ( .A(a[11]), .B(a[10]), .Z(n467) );
  AOI21_X1 U813 ( .B1(n583), .B2(n117), .A(n112), .ZN(n110) );
  NAND2_X1 U814 ( .A1(n40), .A2(n584), .ZN(n31) );
  OAI22_X1 U815 ( .A1(n501), .A2(n489), .B1(n441), .B2(n483), .ZN(n303) );
  INV_X1 U816 ( .A(n495), .ZN(n489) );
  INV_X1 U817 ( .A(n148), .ZN(n146) );
  NAND2_X1 U818 ( .A1(n376), .A2(n304), .ZN(n148) );
  OAI22_X1 U819 ( .A1(n500), .A2(n488), .B1(n428), .B2(n482), .ZN(n302) );
  INV_X1 U820 ( .A(n494), .ZN(n488) );
  OAI21_X1 U821 ( .B1(n32), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X1 U822 ( .B1(n52), .B2(n585), .A(n45), .ZN(n43) );
  AOI21_X1 U823 ( .B1(n590), .B2(n134), .A(n131), .ZN(n129) );
  OAI21_X1 U824 ( .B1(n135), .B2(n137), .A(n136), .ZN(n134) );
  OAI22_X1 U825 ( .A1(n499), .A2(n487), .B1(n415), .B2(n481), .ZN(n301) );
  INV_X1 U826 ( .A(n493), .ZN(n487) );
  AOI21_X1 U827 ( .B1(n126), .B2(n589), .A(n123), .ZN(n121) );
  XNOR2_X1 U828 ( .A(a[9]), .B(a[10]), .ZN(n503) );
  XNOR2_X1 U829 ( .A(n491), .B(n456), .ZN(n378) );
  XNOR2_X1 U830 ( .A(n455), .B(n491), .ZN(n377) );
  INV_X1 U831 ( .A(n491), .ZN(n485) );
  XNOR2_X1 U832 ( .A(n463), .B(n491), .ZN(n385) );
  XNOR2_X1 U833 ( .A(n576), .B(n491), .ZN(n388) );
  XNOR2_X1 U834 ( .A(n491), .B(b[1]), .ZN(n387) );
  XNOR2_X1 U835 ( .A(n491), .B(b[2]), .ZN(n386) );
  XNOR2_X1 U836 ( .A(n491), .B(n458), .ZN(n380) );
  XNOR2_X1 U837 ( .A(n491), .B(n457), .ZN(n379) );
  XNOR2_X1 U838 ( .A(n462), .B(n491), .ZN(n384) );
  XNOR2_X1 U839 ( .A(n491), .B(n461), .ZN(n383) );
  XNOR2_X1 U840 ( .A(n491), .B(n460), .ZN(n382) );
  XNOR2_X1 U841 ( .A(n491), .B(n459), .ZN(n381) );
  NOR2_X1 U842 ( .A1(n31), .A2(n28), .ZN(n26) );
  INV_X1 U843 ( .A(a[0]), .ZN(n508) );
  OAI21_X1 U844 ( .B1(n127), .B2(n129), .A(n128), .ZN(n126) );
  NAND2_X1 U845 ( .A1(n583), .A2(n580), .ZN(n109) );
  INV_X1 U846 ( .A(n561), .ZN(n39) );
  INV_X1 U847 ( .A(n138), .ZN(n137) );
  OAI21_X1 U848 ( .B1(n139), .B2(n141), .A(n140), .ZN(n138) );
  OAI21_X1 U849 ( .B1(n59), .B2(n42), .A(n43), .ZN(n41) );
  INV_X1 U850 ( .A(n59), .ZN(n57) );
  OAI21_X1 U851 ( .B1(n121), .B2(n109), .A(n110), .ZN(n108) );
  INV_X1 U852 ( .A(n219), .ZN(n220) );
  INV_X1 U853 ( .A(n68), .ZN(n66) );
  NAND2_X1 U854 ( .A1(n190), .A2(n195), .ZN(n68) );
  AOI21_X1 U855 ( .B1(n578), .B2(n26), .A(n27), .ZN(n25) );
  AND2_X1 U856 ( .A1(n576), .A2(a[0]), .ZN(product[0]) );
  XNOR2_X1 U857 ( .A(n22), .B(n146), .ZN(product[2]) );
  NAND2_X1 U858 ( .A1(n587), .A2(n145), .ZN(n22) );
  XOR2_X1 U859 ( .A(n20), .B(n137), .Z(product[4]) );
  NAND2_X1 U860 ( .A1(n167), .A2(n136), .ZN(n20) );
  XOR2_X1 U861 ( .A(n18), .B(n577), .Z(product[6]) );
  NAND2_X1 U862 ( .A1(n165), .A2(n128), .ZN(n18) );
  XOR2_X1 U863 ( .A(n21), .B(n141), .Z(product[3]) );
  NAND2_X1 U864 ( .A1(n575), .A2(n140), .ZN(n21) );
  XNOR2_X1 U865 ( .A(n19), .B(n134), .ZN(product[5]) );
  NAND2_X1 U866 ( .A1(n590), .A2(n133), .ZN(n19) );
  XNOR2_X1 U867 ( .A(n126), .B(n17), .ZN(product[7]) );
  NAND2_X1 U868 ( .A1(n589), .A2(n125), .ZN(n17) );
  XNOR2_X1 U869 ( .A(n120), .B(n16), .ZN(product[8]) );
  INV_X1 U870 ( .A(n121), .ZN(n120) );
  XOR2_X1 U871 ( .A(n115), .B(n15), .Z(product[9]) );
  AOI21_X1 U872 ( .B1(n120), .B2(n580), .A(n117), .ZN(n115) );
  XOR2_X1 U873 ( .A(n14), .B(n107), .Z(product[10]) );
  INV_X1 U874 ( .A(n108), .ZN(n107) );
  XNOR2_X1 U875 ( .A(n98), .B(n12), .ZN(product[12]) );
  INV_X1 U876 ( .A(n99), .ZN(n98) );
  XNOR2_X1 U877 ( .A(n37), .B(n4), .ZN(product[20]) );
  OAI21_X1 U878 ( .B1(n69), .B2(n38), .A(n39), .ZN(n37) );
  XNOR2_X1 U879 ( .A(n104), .B(n13), .ZN(product[11]) );
  OAI21_X1 U880 ( .B1(n107), .B2(n105), .A(n106), .ZN(n104) );
  XOR2_X1 U881 ( .A(n566), .B(n6), .Z(product[18]) );
  AOI21_X1 U882 ( .B1(n70), .B2(n56), .A(n57), .ZN(n55) );
  XOR2_X1 U883 ( .A(n77), .B(n9), .Z(product[15]) );
  AOI21_X1 U884 ( .B1(n78), .B2(n98), .A(n79), .ZN(n77) );
  INV_X1 U885 ( .A(n70), .ZN(n69) );
  XNOR2_X1 U886 ( .A(n30), .B(n3), .ZN(product[21]) );
  OAI21_X1 U887 ( .B1(n562), .B2(n31), .A(n567), .ZN(n30) );
  XOR2_X1 U888 ( .A(n84), .B(n10), .Z(product[14]) );
  AOI21_X1 U889 ( .B1(n98), .B2(n85), .A(n86), .ZN(n84) );
  XOR2_X1 U890 ( .A(n64), .B(n7), .Z(product[17]) );
  AOI21_X1 U891 ( .B1(n578), .B2(n582), .A(n66), .ZN(n64) );
  XNOR2_X1 U892 ( .A(n48), .B(n5), .ZN(product[19]) );
  OAI21_X1 U893 ( .B1(n55), .B2(n49), .A(n54), .ZN(n48) );
  XOR2_X1 U894 ( .A(n93), .B(n11), .Z(product[13]) );
  AOI21_X1 U895 ( .B1(n98), .B2(n94), .A(n95), .ZN(n93) );
  INV_X1 U896 ( .A(n25), .ZN(n149) );
  INV_X1 U897 ( .A(n24), .ZN(product[23]) );
endmodule


module datapath_DW_mult_tc_17 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n1, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n40, n41, n42, n43, n44, n48, n50, n51, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n66, n68, n69, n71, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n87, n88, n89,
         n90, n91, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n130, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n142, n144, n145, n147, n148, n149, n150, n152, n156,
         n157, n160, n161, n162, n163, n164, n166, n167, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n286, n287, n288, n289, n290, n291, n292, n293, n295,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n466, n467, n468, n469, n470, n471, n476, n479,
         n480, n481, n482, n483, n485, n488, n491, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n600, n601, n602, n603,
         n604, n605, n606;

  FA_X1 U5 ( .A(n304), .B(n170), .CI(n148), .CO(n25), .S(product[22]) );
  FA_X1 U193 ( .A(n305), .B(n176), .CI(n313), .CO(n172), .S(n173) );
  FA_X1 U194 ( .A(n177), .B(n314), .CI(n180), .CO(n174), .S(n175) );
  FA_X1 U196 ( .A(n184), .B(n306), .CI(n181), .CO(n178), .S(n179) );
  FA_X1 U197 ( .A(n315), .B(n186), .CI(n326), .CO(n180), .S(n181) );
  FA_X1 U198 ( .A(n185), .B(n192), .CI(n190), .CO(n182), .S(n183) );
  FA_X1 U199 ( .A(n316), .B(n327), .CI(n187), .CO(n184), .S(n185) );
  FA_X1 U201 ( .A(n196), .B(n193), .CI(n191), .CO(n188), .S(n189) );
  FA_X1 U202 ( .A(n338), .B(n307), .CI(n198), .CO(n190), .S(n191) );
  FA_X1 U203 ( .A(n317), .B(n200), .CI(n328), .CO(n192), .S(n193) );
  FA_X1 U204 ( .A(n204), .B(n199), .CI(n197), .CO(n194), .S(n195) );
  FA_X1 U205 ( .A(n208), .B(n201), .CI(n206), .CO(n196), .S(n197) );
  FA_X1 U206 ( .A(n329), .B(n318), .CI(n339), .CO(n198), .S(n199) );
  FA_X1 U208 ( .A(n212), .B(n207), .CI(n205), .CO(n202), .S(n203) );
  FA_X1 U209 ( .A(n214), .B(n216), .CI(n209), .CO(n204), .S(n205) );
  FA_X1 U210 ( .A(n218), .B(n319), .CI(n351), .CO(n206), .S(n207) );
  FA_X1 U211 ( .A(n330), .B(n340), .CI(n308), .CO(n208), .S(n209) );
  FA_X1 U212 ( .A(n222), .B(n215), .CI(n213), .CO(n210), .S(n211) );
  FA_X1 U213 ( .A(n217), .B(n226), .CI(n224), .CO(n212), .S(n213) );
  FA_X1 U215 ( .A(n352), .B(n320), .CI(n341), .CO(n216), .S(n217) );
  FA_X1 U217 ( .A(n232), .B(n225), .CI(n223), .CO(n220), .S(n221) );
  FA_X1 U218 ( .A(n227), .B(n236), .CI(n234), .CO(n222), .S(n223) );
  FA_X1 U219 ( .A(n238), .B(n310), .CI(n229), .CO(n224), .S(n225) );
  FA_X1 U220 ( .A(n364), .B(n353), .CI(n342), .CO(n226), .S(n227) );
  FA_X1 U223 ( .A(n242), .B(n235), .CI(n233), .CO(n230), .S(n231) );
  FA_X1 U224 ( .A(n244), .B(n246), .CI(n237), .CO(n232), .S(n233) );
  FA_X1 U225 ( .A(n311), .B(n354), .CI(n239), .CO(n234), .S(n235) );
  FA_X1 U226 ( .A(n322), .B(n343), .CI(n365), .CO(n236), .S(n237) );
  HA_X1 U227 ( .A(n298), .B(n332), .CO(n238), .S(n239) );
  FA_X1 U228 ( .A(n250), .B(n245), .CI(n243), .CO(n240), .S(n241) );
  FA_X1 U229 ( .A(n252), .B(n254), .CI(n247), .CO(n242), .S(n243) );
  FA_X1 U230 ( .A(n344), .B(n355), .CI(n323), .CO(n244), .S(n245) );
  FA_X1 U231 ( .A(n366), .B(n312), .CI(n333), .CO(n246), .S(n247) );
  FA_X1 U232 ( .A(n253), .B(n258), .CI(n251), .CO(n248), .S(n249) );
  FA_X1 U233 ( .A(n255), .B(n334), .CI(n260), .CO(n250), .S(n251) );
  FA_X1 U234 ( .A(n345), .B(n356), .CI(n324), .CO(n252), .S(n253) );
  HA_X1 U235 ( .A(n367), .B(n299), .CO(n254), .S(n255) );
  FA_X1 U236 ( .A(n261), .B(n264), .CI(n259), .CO(n256), .S(n257) );
  FA_X1 U238 ( .A(n368), .B(n325), .CI(n357), .CO(n260), .S(n261) );
  FA_X1 U239 ( .A(n270), .B(n267), .CI(n265), .CO(n262), .S(n263) );
  FA_X1 U240 ( .A(n336), .B(n358), .CI(n347), .CO(n264), .S(n265) );
  HA_X1 U241 ( .A(n300), .B(n369), .CO(n266), .S(n267) );
  FA_X1 U242 ( .A(n274), .B(n348), .CI(n271), .CO(n268), .S(n269) );
  FA_X1 U243 ( .A(n370), .B(n337), .CI(n359), .CO(n270), .S(n271) );
  FA_X1 U244 ( .A(n349), .B(n360), .CI(n275), .CO(n272), .S(n273) );
  HA_X1 U245 ( .A(n301), .B(n371), .CO(n274), .S(n275) );
  FA_X1 U246 ( .A(n372), .B(n350), .CI(n361), .CO(n276), .S(n277) );
  HA_X1 U247 ( .A(n373), .B(n302), .CO(n278), .S(n279) );
  BUF_X2 U483 ( .A(b[3]), .Z(n462) );
  INV_X1 U484 ( .A(n160), .ZN(n559) );
  AOI21_X2 U485 ( .B1(n117), .B2(n125), .A(n118), .ZN(n116) );
  BUF_X2 U486 ( .A(a[5]), .Z(n493) );
  BUF_X2 U487 ( .A(b[2]), .Z(n463) );
  BUF_X2 U488 ( .A(n505), .Z(n481) );
  BUF_X2 U489 ( .A(n503), .Z(n479) );
  BUF_X1 U490 ( .A(b[10]), .Z(n455) );
  BUF_X2 U491 ( .A(b[11]), .Z(n454) );
  BUF_X2 U492 ( .A(a[1]), .Z(n495) );
  CLKBUF_X1 U493 ( .A(n499), .Z(n560) );
  BUF_X2 U494 ( .A(n499), .Z(n561) );
  NAND2_X1 U495 ( .A1(n505), .A2(n469), .ZN(n499) );
  CLKBUF_X1 U496 ( .A(n108), .Z(n562) );
  OR2_X1 U497 ( .A1(n101), .A2(n96), .ZN(n563) );
  BUF_X1 U498 ( .A(b[8]), .Z(n457) );
  AOI21_X1 U499 ( .B1(n596), .B2(n133), .A(n130), .ZN(n564) );
  OAI21_X2 U500 ( .B1(n134), .B2(n136), .A(n135), .ZN(n133) );
  OR2_X1 U501 ( .A1(n331), .A2(n321), .ZN(n228) );
  NAND2_X2 U502 ( .A1(n467), .A2(n503), .ZN(n497) );
  INV_X1 U503 ( .A(n100), .ZN(n565) );
  CLKBUF_X1 U504 ( .A(n111), .Z(n566) );
  CLKBUF_X1 U505 ( .A(n502), .Z(n567) );
  BUF_X2 U506 ( .A(n502), .Z(n568) );
  XNOR2_X1 U507 ( .A(a[5]), .B(a[6]), .ZN(n569) );
  CLKBUF_X1 U508 ( .A(n335), .Z(n570) );
  CLKBUF_X1 U509 ( .A(n591), .Z(n571) );
  CLKBUF_X1 U510 ( .A(n1), .Z(n572) );
  CLKBUF_X3 U511 ( .A(b[0]), .Z(n1) );
  NOR2_X1 U512 ( .A1(n231), .A2(n240), .ZN(n573) );
  BUF_X1 U513 ( .A(b[4]), .Z(n461) );
  CLKBUF_X1 U514 ( .A(n96), .Z(n574) );
  BUF_X1 U515 ( .A(b[6]), .Z(n459) );
  BUF_X2 U516 ( .A(n504), .Z(n480) );
  CLKBUF_X1 U517 ( .A(b[1]), .Z(n464) );
  BUF_X1 U518 ( .A(b[1]), .Z(n575) );
  BUF_X1 U519 ( .A(b[7]), .Z(n458) );
  XOR2_X1 U520 ( .A(n219), .B(n309), .Z(n576) );
  XOR2_X1 U521 ( .A(n228), .B(n576), .Z(n215) );
  NAND2_X1 U522 ( .A1(n228), .A2(n219), .ZN(n577) );
  NAND2_X1 U523 ( .A1(n228), .A2(n309), .ZN(n578) );
  NAND2_X1 U524 ( .A1(n219), .A2(n309), .ZN(n579) );
  NAND3_X1 U525 ( .A1(n577), .A2(n578), .A3(n579), .ZN(n214) );
  XOR2_X1 U526 ( .A(n335), .B(n346), .Z(n580) );
  XOR2_X1 U527 ( .A(n266), .B(n580), .Z(n259) );
  NAND2_X1 U528 ( .A1(n266), .A2(n570), .ZN(n581) );
  NAND2_X1 U529 ( .A1(n266), .A2(n346), .ZN(n582) );
  NAND2_X1 U530 ( .A1(n570), .A2(n346), .ZN(n583) );
  NAND3_X1 U531 ( .A1(n581), .A2(n582), .A3(n583), .ZN(n258) );
  OAI21_X1 U532 ( .B1(n116), .B2(n114), .A(n115), .ZN(n584) );
  BUF_X1 U533 ( .A(b[9]), .Z(n456) );
  NOR2_X1 U534 ( .A1(n257), .A2(n262), .ZN(n585) );
  NOR2_X1 U535 ( .A1(n257), .A2(n262), .ZN(n119) );
  OR2_X1 U536 ( .A1(n231), .A2(n240), .ZN(n586) );
  OR2_X1 U537 ( .A1(n195), .A2(n202), .ZN(n587) );
  XNOR2_X1 U538 ( .A(n51), .B(n588), .ZN(product[19]) );
  AND2_X1 U539 ( .A1(n595), .A2(n50), .ZN(n588) );
  NOR2_X1 U540 ( .A1(n211), .A2(n220), .ZN(n589) );
  AOI21_X1 U541 ( .B1(n105), .B2(n584), .A(n106), .ZN(n590) );
  OAI21_X1 U542 ( .B1(n590), .B2(n76), .A(n77), .ZN(n591) );
  XNOR2_X1 U543 ( .A(n60), .B(n592), .ZN(product[18]) );
  AND2_X1 U544 ( .A1(n152), .A2(n59), .ZN(n592) );
  XOR2_X1 U545 ( .A(n124), .B(n18), .Z(product[7]) );
  OR2_X1 U546 ( .A1(n183), .A2(n188), .ZN(n593) );
  OR2_X1 U547 ( .A1(n189), .A2(n194), .ZN(n594) );
  OR2_X1 U548 ( .A1(n175), .A2(n178), .ZN(n595) );
  OR2_X1 U549 ( .A1(n273), .A2(n276), .ZN(n596) );
  OR2_X1 U550 ( .A1(n374), .A2(n363), .ZN(n597) );
  OR2_X1 U551 ( .A1(n375), .A2(n303), .ZN(n598) );
  BUF_X2 U552 ( .A(n506), .Z(n482) );
  BUF_X2 U553 ( .A(n491), .Z(n602) );
  BUF_X2 U554 ( .A(a[11]), .Z(n604) );
  BUF_X2 U555 ( .A(a[11]), .Z(n603) );
  AND2_X1 U556 ( .A1(n598), .A2(n147), .ZN(product[1]) );
  NOR2_X1 U557 ( .A1(n174), .A2(n173), .ZN(n40) );
  NAND2_X1 U558 ( .A1(n149), .A2(n34), .ZN(n4) );
  NOR2_X1 U559 ( .A1(n172), .A2(n171), .ZN(n33) );
  INV_X1 U560 ( .A(n33), .ZN(n149) );
  NAND2_X1 U561 ( .A1(n172), .A2(n171), .ZN(n34) );
  AOI21_X1 U562 ( .B1(n31), .B2(n48), .A(n32), .ZN(n30) );
  NAND2_X1 U563 ( .A1(n595), .A2(n31), .ZN(n29) );
  INV_X1 U564 ( .A(n40), .ZN(n150) );
  NOR2_X1 U565 ( .A1(n40), .A2(n33), .ZN(n31) );
  NAND2_X1 U566 ( .A1(n150), .A2(n41), .ZN(n5) );
  OAI21_X1 U567 ( .B1(n41), .B2(n33), .A(n34), .ZN(n32) );
  INV_X1 U568 ( .A(n50), .ZN(n48) );
  NAND2_X1 U569 ( .A1(n174), .A2(n173), .ZN(n41) );
  NAND2_X1 U570 ( .A1(n175), .A2(n178), .ZN(n50) );
  NOR2_X1 U571 ( .A1(n43), .A2(n40), .ZN(n36) );
  INV_X1 U572 ( .A(n58), .ZN(n152) );
  NOR2_X1 U573 ( .A1(n179), .A2(n182), .ZN(n58) );
  NAND2_X1 U574 ( .A1(n179), .A2(n182), .ZN(n59) );
  BUF_X2 U575 ( .A(n507), .Z(n483) );
  INV_X1 U576 ( .A(n289), .ZN(n338) );
  INV_X1 U577 ( .A(n156), .ZN(n85) );
  CLKBUF_X3 U578 ( .A(a[3]), .Z(n494) );
  NAND2_X1 U579 ( .A1(n593), .A2(n68), .ZN(n8) );
  NOR2_X1 U580 ( .A1(n269), .A2(n272), .ZN(n126) );
  BUF_X2 U581 ( .A(n491), .Z(n601) );
  NAND2_X1 U582 ( .A1(n183), .A2(n188), .ZN(n68) );
  XNOR2_X1 U583 ( .A(n602), .B(n457), .ZN(n392) );
  XNOR2_X1 U584 ( .A(n603), .B(n457), .ZN(n379) );
  INV_X1 U585 ( .A(n283), .ZN(n313) );
  BUF_X1 U586 ( .A(a[9]), .Z(n491) );
  XNOR2_X1 U587 ( .A(n495), .B(n456), .ZN(n443) );
  XNOR2_X1 U588 ( .A(n495), .B(n455), .ZN(n442) );
  NAND2_X1 U589 ( .A1(n157), .A2(n97), .ZN(n12) );
  OAI21_X1 U590 ( .B1(n44), .B2(n40), .A(n41), .ZN(n37) );
  XNOR2_X1 U591 ( .A(n602), .B(n459), .ZN(n394) );
  XNOR2_X1 U592 ( .A(n604), .B(n459), .ZN(n381) );
  INV_X1 U593 ( .A(n93), .ZN(n91) );
  INV_X1 U594 ( .A(n563), .ZN(n90) );
  NOR2_X1 U595 ( .A1(n563), .A2(n85), .ZN(n83) );
  OAI22_X1 U596 ( .A1(n497), .A2(n392), .B1(n391), .B2(n479), .ZN(n316) );
  OAI22_X1 U597 ( .A1(n497), .A2(n391), .B1(n390), .B2(n479), .ZN(n315) );
  OAI22_X1 U598 ( .A1(n497), .A2(n390), .B1(n389), .B2(n479), .ZN(n314) );
  AOI21_X1 U599 ( .B1(n497), .B2(n479), .A(n389), .ZN(n283) );
  OAI22_X1 U600 ( .A1(n497), .A2(n485), .B1(n401), .B2(n479), .ZN(n299) );
  NAND2_X1 U601 ( .A1(n277), .A2(n278), .ZN(n135) );
  BUF_X1 U602 ( .A(n491), .Z(n600) );
  NOR2_X1 U603 ( .A1(n241), .A2(n248), .ZN(n110) );
  NOR2_X1 U604 ( .A1(n263), .A2(n268), .ZN(n122) );
  NAND2_X2 U605 ( .A1(n468), .A2(n569), .ZN(n498) );
  NOR2_X1 U606 ( .A1(n195), .A2(n202), .ZN(n80) );
  INV_X1 U607 ( .A(n481), .ZN(n290) );
  INV_X1 U608 ( .A(n144), .ZN(n142) );
  INV_X1 U609 ( .A(n126), .ZN(n164) );
  XNOR2_X1 U610 ( .A(n495), .B(n459), .ZN(n446) );
  NAND2_X1 U611 ( .A1(n99), .A2(n565), .ZN(n13) );
  INV_X1 U612 ( .A(n102), .ZN(n100) );
  NAND2_X1 U613 ( .A1(n211), .A2(n220), .ZN(n97) );
  NAND2_X1 U614 ( .A1(n162), .A2(n120), .ZN(n17) );
  NAND2_X1 U615 ( .A1(n263), .A2(n268), .ZN(n123) );
  INV_X1 U616 ( .A(n495), .ZN(n297) );
  OAI22_X1 U617 ( .A1(n501), .A2(n297), .B1(n453), .B2(n483), .ZN(n303) );
  INV_X1 U618 ( .A(n87), .ZN(n156) );
  AOI21_X1 U619 ( .B1(n476), .B2(n482), .A(n428), .ZN(n292) );
  INV_X1 U620 ( .A(n114), .ZN(n161) );
  NOR2_X1 U621 ( .A1(n249), .A2(n256), .ZN(n114) );
  NAND2_X1 U622 ( .A1(n221), .A2(n230), .ZN(n102) );
  XNOR2_X1 U623 ( .A(n495), .B(n454), .ZN(n441) );
  NAND2_X1 U624 ( .A1(n269), .A2(n272), .ZN(n127) );
  XNOR2_X1 U625 ( .A(n495), .B(n457), .ZN(n444) );
  OAI22_X1 U626 ( .A1(n497), .A2(n394), .B1(n393), .B2(n479), .ZN(n318) );
  OAI22_X1 U627 ( .A1(n497), .A2(n393), .B1(n392), .B2(n479), .ZN(n317) );
  INV_X1 U628 ( .A(n138), .ZN(n167) );
  NOR2_X1 U629 ( .A1(n279), .A2(n362), .ZN(n138) );
  XNOR2_X1 U630 ( .A(n462), .B(n495), .ZN(n449) );
  INV_X1 U631 ( .A(n122), .ZN(n163) );
  NAND2_X1 U632 ( .A1(n249), .A2(n256), .ZN(n115) );
  NAND2_X1 U633 ( .A1(n257), .A2(n262), .ZN(n120) );
  INV_X1 U634 ( .A(n132), .ZN(n130) );
  OAI22_X1 U635 ( .A1(n561), .A2(n425), .B1(n424), .B2(n481), .ZN(n348) );
  OAI22_X1 U636 ( .A1(n561), .A2(n426), .B1(n425), .B2(n481), .ZN(n349) );
  OAI22_X1 U637 ( .A1(n561), .A2(n422), .B1(n421), .B2(n481), .ZN(n345) );
  OAI22_X1 U638 ( .A1(n560), .A2(n423), .B1(n422), .B2(n481), .ZN(n346) );
  AOI21_X1 U639 ( .B1(n561), .B2(n481), .A(n415), .ZN(n289) );
  OAI22_X1 U640 ( .A1(n561), .A2(n418), .B1(n417), .B2(n481), .ZN(n341) );
  OAI22_X1 U641 ( .A1(n561), .A2(n421), .B1(n420), .B2(n481), .ZN(n344) );
  OAI22_X1 U642 ( .A1(n561), .A2(n416), .B1(n415), .B2(n481), .ZN(n339) );
  OAI22_X1 U643 ( .A1(n561), .A2(n419), .B1(n418), .B2(n481), .ZN(n342) );
  OAI22_X1 U644 ( .A1(n560), .A2(n420), .B1(n419), .B2(n481), .ZN(n343) );
  OAI22_X1 U645 ( .A1(n561), .A2(n417), .B1(n416), .B2(n481), .ZN(n340) );
  OAI22_X1 U646 ( .A1(n561), .A2(n291), .B1(n427), .B2(n481), .ZN(n301) );
  OAI22_X1 U647 ( .A1(n561), .A2(n424), .B1(n423), .B2(n481), .ZN(n347) );
  INV_X1 U648 ( .A(n95), .ZN(n93) );
  NAND2_X1 U649 ( .A1(n587), .A2(n81), .ZN(n10) );
  INV_X1 U650 ( .A(n479), .ZN(n284) );
  NAND2_X1 U651 ( .A1(n273), .A2(n276), .ZN(n132) );
  NAND2_X2 U652 ( .A1(n502), .A2(n466), .ZN(n496) );
  XOR2_X1 U653 ( .A(a[11]), .B(a[10]), .Z(n466) );
  NAND2_X1 U654 ( .A1(n160), .A2(n566), .ZN(n15) );
  INV_X1 U655 ( .A(n110), .ZN(n160) );
  INV_X1 U656 ( .A(n134), .ZN(n166) );
  NOR2_X1 U657 ( .A1(n277), .A2(n278), .ZN(n134) );
  XNOR2_X1 U658 ( .A(n493), .B(n454), .ZN(n415) );
  XNOR2_X1 U659 ( .A(n493), .B(n462), .ZN(n423) );
  XNOR2_X1 U660 ( .A(n493), .B(n459), .ZN(n420) );
  XNOR2_X1 U661 ( .A(n493), .B(n456), .ZN(n417) );
  XNOR2_X1 U662 ( .A(n493), .B(n455), .ZN(n416) );
  XNOR2_X1 U663 ( .A(n493), .B(n457), .ZN(n418) );
  OAI22_X1 U664 ( .A1(n399), .A2(n479), .B1(n497), .B2(n400), .ZN(n324) );
  INV_X1 U665 ( .A(n482), .ZN(n293) );
  OAI22_X1 U666 ( .A1(n438), .A2(n482), .B1(n476), .B2(n439), .ZN(n362) );
  OAI22_X1 U667 ( .A1(n438), .A2(n476), .B1(n437), .B2(n482), .ZN(n361) );
  OAI22_X1 U668 ( .A1(n437), .A2(n476), .B1(n436), .B2(n482), .ZN(n360) );
  OAI22_X1 U669 ( .A1(n476), .A2(n436), .B1(n435), .B2(n482), .ZN(n359) );
  OAI22_X1 U670 ( .A1(n476), .A2(n435), .B1(n434), .B2(n482), .ZN(n358) );
  OAI22_X1 U671 ( .A1(n476), .A2(n434), .B1(n433), .B2(n482), .ZN(n357) );
  OAI22_X1 U672 ( .A1(n476), .A2(n433), .B1(n432), .B2(n482), .ZN(n356) );
  OAI22_X1 U673 ( .A1(n476), .A2(n431), .B1(n430), .B2(n482), .ZN(n354) );
  OAI22_X1 U674 ( .A1(n476), .A2(n430), .B1(n429), .B2(n482), .ZN(n353) );
  OAI22_X1 U675 ( .A1(n476), .A2(n429), .B1(n428), .B2(n482), .ZN(n352) );
  BUF_X2 U676 ( .A(n500), .Z(n476) );
  AND2_X1 U677 ( .A1(n572), .A2(n293), .ZN(n363) );
  NAND2_X1 U678 ( .A1(n279), .A2(n362), .ZN(n139) );
  INV_X1 U679 ( .A(n292), .ZN(n351) );
  XNOR2_X1 U680 ( .A(n495), .B(n460), .ZN(n447) );
  XNOR2_X1 U681 ( .A(n493), .B(n460), .ZN(n421) );
  BUF_X2 U682 ( .A(b[5]), .Z(n460) );
  AOI21_X1 U683 ( .B1(n57), .B2(n595), .A(n48), .ZN(n44) );
  AOI21_X1 U684 ( .B1(n501), .B2(n483), .A(n441), .ZN(n295) );
  OAI22_X1 U685 ( .A1(n501), .A2(n445), .B1(n444), .B2(n483), .ZN(n368) );
  OAI22_X1 U686 ( .A1(n501), .A2(n447), .B1(n446), .B2(n483), .ZN(n370) );
  OAI22_X1 U687 ( .A1(n450), .A2(n501), .B1(n449), .B2(n483), .ZN(n373) );
  OAI22_X1 U688 ( .A1(n501), .A2(n444), .B1(n443), .B2(n483), .ZN(n367) );
  OAI22_X1 U689 ( .A1(n501), .A2(n449), .B1(n448), .B2(n483), .ZN(n372) );
  OAI22_X1 U690 ( .A1(n451), .A2(n483), .B1(n501), .B2(n452), .ZN(n375) );
  OAI22_X1 U691 ( .A1(n501), .A2(n448), .B1(n447), .B2(n483), .ZN(n371) );
  OAI22_X1 U692 ( .A1(n451), .A2(n501), .B1(n450), .B2(n483), .ZN(n374) );
  NAND2_X1 U693 ( .A1(n375), .A2(n303), .ZN(n147) );
  NAND2_X1 U694 ( .A1(n374), .A2(n363), .ZN(n144) );
  NAND2_X1 U695 ( .A1(n195), .A2(n202), .ZN(n81) );
  NAND2_X1 U696 ( .A1(n241), .A2(n248), .ZN(n111) );
  XNOR2_X1 U697 ( .A(n461), .B(n495), .ZN(n448) );
  XNOR2_X1 U698 ( .A(n493), .B(n461), .ZN(n422) );
  INV_X1 U699 ( .A(n574), .ZN(n157) );
  NOR2_X1 U700 ( .A1(n211), .A2(n220), .ZN(n96) );
  OAI22_X1 U701 ( .A1(n496), .A2(n377), .B1(n568), .B2(n376), .ZN(n170) );
  XOR2_X1 U702 ( .A(a[5]), .B(a[4]), .Z(n469) );
  BUF_X2 U703 ( .A(a[7]), .Z(n606) );
  INV_X1 U704 ( .A(n585), .ZN(n162) );
  NOR2_X1 U705 ( .A1(n101), .A2(n96), .ZN(n94) );
  BUF_X2 U706 ( .A(a[7]), .Z(n605) );
  NOR2_X1 U707 ( .A1(n54), .A2(n29), .ZN(n27) );
  INV_X1 U708 ( .A(n56), .ZN(n54) );
  OAI22_X1 U709 ( .A1(n497), .A2(n395), .B1(n394), .B2(n479), .ZN(n319) );
  OAI22_X1 U710 ( .A1(n497), .A2(n396), .B1(n395), .B2(n479), .ZN(n320) );
  XNOR2_X1 U711 ( .A(a[1]), .B(a[2]), .ZN(n506) );
  OR2_X1 U712 ( .A1(n1), .A2(n488), .ZN(n440) );
  XNOR2_X1 U713 ( .A(n1), .B(n602), .ZN(n400) );
  AND2_X1 U714 ( .A1(n572), .A2(n284), .ZN(n325) );
  AND2_X1 U715 ( .A1(n572), .A2(n290), .ZN(n350) );
  XNOR2_X1 U716 ( .A(n1), .B(n493), .ZN(n426) );
  OR2_X1 U717 ( .A1(n1), .A2(n297), .ZN(n453) );
  OR2_X1 U718 ( .A1(n1), .A2(n485), .ZN(n401) );
  OR2_X1 U719 ( .A1(n291), .A2(n1), .ZN(n427) );
  OR2_X1 U720 ( .A1(n1), .A2(n288), .ZN(n414) );
  XNOR2_X1 U721 ( .A(n575), .B(n495), .ZN(n451) );
  XNOR2_X1 U722 ( .A(n575), .B(n493), .ZN(n425) );
  XNOR2_X1 U723 ( .A(n575), .B(n602), .ZN(n399) );
  OAI21_X1 U724 ( .B1(n589), .B2(n102), .A(n97), .ZN(n95) );
  OAI22_X1 U725 ( .A1(n501), .A2(n443), .B1(n442), .B2(n483), .ZN(n366) );
  XNOR2_X1 U726 ( .A(n464), .B(n605), .ZN(n412) );
  XNOR2_X1 U727 ( .A(n605), .B(n457), .ZN(n405) );
  XNOR2_X1 U728 ( .A(n605), .B(n454), .ZN(n402) );
  XNOR2_X1 U729 ( .A(n461), .B(n600), .ZN(n396) );
  OAI22_X1 U730 ( .A1(n498), .A2(n407), .B1(n480), .B2(n406), .ZN(n218) );
  OR2_X1 U731 ( .A1(n1), .A2(n282), .ZN(n388) );
  OAI22_X1 U732 ( .A1(n497), .A2(n397), .B1(n396), .B2(n479), .ZN(n321) );
  OAI21_X1 U733 ( .B1(n107), .B2(n111), .A(n108), .ZN(n106) );
  NOR2_X1 U734 ( .A1(n573), .A2(n110), .ZN(n105) );
  NAND2_X1 U735 ( .A1(n586), .A2(n562), .ZN(n14) );
  NOR2_X1 U736 ( .A1(n231), .A2(n240), .ZN(n107) );
  XNOR2_X1 U737 ( .A(n462), .B(n600), .ZN(n397) );
  XOR2_X1 U738 ( .A(a[9]), .B(a[8]), .Z(n467) );
  OAI22_X1 U739 ( .A1(n501), .A2(n442), .B1(n441), .B2(n483), .ZN(n365) );
  XNOR2_X1 U740 ( .A(n572), .B(n494), .ZN(n439) );
  XNOR2_X1 U741 ( .A(n464), .B(n494), .ZN(n438) );
  XNOR2_X1 U742 ( .A(n494), .B(n462), .ZN(n436) );
  XNOR2_X1 U743 ( .A(n494), .B(n461), .ZN(n435) );
  XNOR2_X1 U744 ( .A(n494), .B(n460), .ZN(n434) );
  XNOR2_X1 U745 ( .A(n494), .B(n456), .ZN(n430) );
  XNOR2_X1 U746 ( .A(n494), .B(n459), .ZN(n433) );
  XNOR2_X1 U747 ( .A(n494), .B(n457), .ZN(n431) );
  XNOR2_X1 U748 ( .A(n494), .B(n455), .ZN(n429) );
  XNOR2_X1 U749 ( .A(n494), .B(n454), .ZN(n428) );
  XNOR2_X1 U750 ( .A(n461), .B(n606), .ZN(n409) );
  INV_X1 U751 ( .A(n295), .ZN(n364) );
  XNOR2_X1 U752 ( .A(n601), .B(n454), .ZN(n389) );
  XNOR2_X1 U753 ( .A(n601), .B(n456), .ZN(n391) );
  XNOR2_X1 U754 ( .A(n601), .B(n460), .ZN(n395) );
  XNOR2_X1 U755 ( .A(n463), .B(n495), .ZN(n450) );
  XNOR2_X1 U756 ( .A(n463), .B(n494), .ZN(n437) );
  XNOR2_X1 U757 ( .A(n463), .B(n493), .ZN(n424) );
  NAND2_X1 U758 ( .A1(n470), .A2(n506), .ZN(n500) );
  XOR2_X1 U759 ( .A(a[3]), .B(a[2]), .Z(n470) );
  OAI22_X1 U760 ( .A1(n476), .A2(n432), .B1(n431), .B2(n482), .ZN(n355) );
  OAI22_X1 U761 ( .A1(n399), .A2(n497), .B1(n398), .B2(n479), .ZN(n323) );
  XOR2_X1 U762 ( .A(a[1]), .B(a[0]), .Z(n471) );
  XNOR2_X1 U763 ( .A(n463), .B(n602), .ZN(n398) );
  INV_X1 U764 ( .A(n567), .ZN(n281) );
  OAI22_X1 U765 ( .A1(n386), .A2(n568), .B1(n496), .B2(n387), .ZN(n311) );
  OAI22_X1 U766 ( .A1(n386), .A2(n496), .B1(n385), .B2(n568), .ZN(n310) );
  OAI22_X1 U767 ( .A1(n385), .A2(n496), .B1(n384), .B2(n568), .ZN(n309) );
  OAI22_X1 U768 ( .A1(n496), .A2(n384), .B1(n383), .B2(n568), .ZN(n308) );
  OAI22_X1 U769 ( .A1(n496), .A2(n380), .B1(n568), .B2(n379), .ZN(n306) );
  OAI22_X1 U770 ( .A1(n496), .A2(n378), .B1(n568), .B2(n377), .ZN(n305) );
  AOI21_X1 U771 ( .B1(n496), .B2(n568), .A(n376), .ZN(n280) );
  OAI22_X1 U772 ( .A1(n496), .A2(n282), .B1(n388), .B2(n567), .ZN(n298) );
  AND2_X1 U773 ( .A1(n1), .A2(n281), .ZN(n312) );
  INV_X1 U774 ( .A(n170), .ZN(n171) );
  INV_X1 U775 ( .A(n280), .ZN(n304) );
  XNOR2_X1 U776 ( .A(a[3]), .B(a[4]), .ZN(n505) );
  XNOR2_X1 U777 ( .A(a[7]), .B(a[8]), .ZN(n503) );
  NOR2_X1 U778 ( .A1(n87), .A2(n80), .ZN(n78) );
  NAND2_X1 U779 ( .A1(n156), .A2(n88), .ZN(n11) );
  OAI21_X1 U780 ( .B1(n93), .B2(n85), .A(n88), .ZN(n84) );
  NOR2_X1 U781 ( .A1(n203), .A2(n210), .ZN(n87) );
  OAI22_X1 U782 ( .A1(n398), .A2(n497), .B1(n397), .B2(n479), .ZN(n322) );
  XNOR2_X1 U783 ( .A(n606), .B(n460), .ZN(n408) );
  XNOR2_X1 U784 ( .A(n605), .B(n455), .ZN(n403) );
  XNOR2_X1 U785 ( .A(n462), .B(n605), .ZN(n410) );
  XNOR2_X1 U786 ( .A(n463), .B(n605), .ZN(n411) );
  INV_X1 U787 ( .A(n606), .ZN(n288) );
  INV_X1 U788 ( .A(n601), .ZN(n485) );
  XNOR2_X1 U789 ( .A(n601), .B(n455), .ZN(n390) );
  INV_X1 U790 ( .A(n603), .ZN(n282) );
  XNOR2_X1 U791 ( .A(n462), .B(n603), .ZN(n384) );
  XNOR2_X1 U792 ( .A(n463), .B(n603), .ZN(n385) );
  XNOR2_X1 U793 ( .A(n464), .B(n603), .ZN(n386) );
  XNOR2_X1 U794 ( .A(n603), .B(n455), .ZN(n377) );
  XNOR2_X1 U795 ( .A(n603), .B(n456), .ZN(n378) );
  OAI22_X1 U796 ( .A1(n496), .A2(n383), .B1(n568), .B2(n382), .ZN(n200) );
  INV_X1 U797 ( .A(n200), .ZN(n201) );
  OAI22_X1 U798 ( .A1(n496), .A2(n382), .B1(n568), .B2(n381), .ZN(n307) );
  OAI22_X1 U799 ( .A1(n496), .A2(n379), .B1(n568), .B2(n378), .ZN(n176) );
  INV_X1 U800 ( .A(n176), .ZN(n177) );
  OAI22_X1 U801 ( .A1(n496), .A2(n381), .B1(n568), .B2(n380), .ZN(n186) );
  INV_X1 U802 ( .A(n186), .ZN(n187) );
  XNOR2_X1 U803 ( .A(n461), .B(n604), .ZN(n383) );
  XNOR2_X1 U804 ( .A(n454), .B(n604), .ZN(n376) );
  XNOR2_X1 U805 ( .A(n1), .B(n604), .ZN(n387) );
  XNOR2_X1 U806 ( .A(n604), .B(n460), .ZN(n382) );
  AOI21_X1 U807 ( .B1(n597), .B2(n145), .A(n142), .ZN(n140) );
  NOR2_X1 U808 ( .A1(n585), .A2(n122), .ZN(n117) );
  NAND2_X2 U809 ( .A1(n471), .A2(n507), .ZN(n501) );
  INV_X1 U810 ( .A(a[0]), .ZN(n507) );
  OAI21_X1 U811 ( .B1(n119), .B2(n123), .A(n120), .ZN(n118) );
  NAND2_X1 U812 ( .A1(n231), .A2(n240), .ZN(n108) );
  NAND2_X1 U813 ( .A1(n56), .A2(n595), .ZN(n43) );
  AOI21_X1 U814 ( .B1(n596), .B2(n133), .A(n130), .ZN(n128) );
  OAI21_X1 U815 ( .B1(n55), .B2(n29), .A(n30), .ZN(n28) );
  INV_X1 U816 ( .A(n101), .ZN(n99) );
  NOR2_X1 U817 ( .A1(n221), .A2(n230), .ZN(n101) );
  INV_X1 U818 ( .A(n57), .ZN(n55) );
  INV_X1 U819 ( .A(n68), .ZN(n66) );
  OAI21_X1 U820 ( .B1(n116), .B2(n114), .A(n115), .ZN(n113) );
  INV_X1 U821 ( .A(n504), .ZN(n287) );
  OAI22_X1 U822 ( .A1(n412), .A2(n480), .B1(n498), .B2(n413), .ZN(n336) );
  OAI22_X1 U823 ( .A1(n412), .A2(n498), .B1(n411), .B2(n480), .ZN(n335) );
  OAI22_X1 U824 ( .A1(n411), .A2(n498), .B1(n480), .B2(n410), .ZN(n334) );
  OAI22_X1 U825 ( .A1(n498), .A2(n410), .B1(n480), .B2(n409), .ZN(n333) );
  OAI22_X1 U826 ( .A1(n409), .A2(n498), .B1(n480), .B2(n408), .ZN(n332) );
  OAI22_X1 U827 ( .A1(n498), .A2(n406), .B1(n480), .B2(n405), .ZN(n330) );
  OAI22_X1 U828 ( .A1(n498), .A2(n405), .B1(n480), .B2(n404), .ZN(n329) );
  OAI22_X1 U829 ( .A1(n498), .A2(n404), .B1(n480), .B2(n403), .ZN(n328) );
  OAI22_X1 U830 ( .A1(n498), .A2(n403), .B1(n480), .B2(n402), .ZN(n327) );
  AOI21_X1 U831 ( .B1(n498), .B2(n480), .A(n402), .ZN(n286) );
  OAI22_X1 U832 ( .A1(n498), .A2(n288), .B1(n414), .B2(n480), .ZN(n300) );
  AND2_X1 U833 ( .A1(n1), .A2(n287), .ZN(n337) );
  INV_X1 U834 ( .A(n218), .ZN(n219) );
  INV_X1 U835 ( .A(n286), .ZN(n326) );
  XNOR2_X1 U836 ( .A(n321), .B(n331), .ZN(n229) );
  OAI22_X1 U837 ( .A1(n498), .A2(n408), .B1(n407), .B2(n480), .ZN(n331) );
  XNOR2_X1 U838 ( .A(n606), .B(n459), .ZN(n407) );
  OAI21_X1 U839 ( .B1(n590), .B2(n76), .A(n77), .ZN(n75) );
  NAND2_X1 U840 ( .A1(n94), .A2(n78), .ZN(n76) );
  AOI21_X1 U841 ( .B1(n105), .B2(n113), .A(n106), .ZN(n104) );
  XOR2_X1 U842 ( .A(a[7]), .B(a[6]), .Z(n468) );
  XNOR2_X1 U843 ( .A(n495), .B(n458), .ZN(n445) );
  XNOR2_X1 U844 ( .A(n494), .B(n458), .ZN(n432) );
  XNOR2_X1 U845 ( .A(n493), .B(n458), .ZN(n419) );
  XNOR2_X1 U846 ( .A(n605), .B(n458), .ZN(n406) );
  XNOR2_X1 U847 ( .A(n601), .B(n458), .ZN(n393) );
  XNOR2_X1 U848 ( .A(n604), .B(n458), .ZN(n380) );
  OAI22_X1 U849 ( .A1(n501), .A2(n446), .B1(n445), .B2(n483), .ZN(n369) );
  INV_X1 U850 ( .A(n137), .ZN(n136) );
  OAI21_X1 U851 ( .B1(n64), .B2(n58), .A(n59), .ZN(n57) );
  INV_X1 U852 ( .A(n64), .ZN(n62) );
  AOI21_X1 U853 ( .B1(n71), .B2(n593), .A(n66), .ZN(n64) );
  INV_X1 U854 ( .A(n493), .ZN(n291) );
  XNOR2_X1 U855 ( .A(a[5]), .B(a[6]), .ZN(n504) );
  AOI21_X1 U856 ( .B1(n95), .B2(n78), .A(n79), .ZN(n77) );
  OAI21_X1 U857 ( .B1(n88), .B2(n80), .A(n81), .ZN(n79) );
  XNOR2_X1 U858 ( .A(n605), .B(n456), .ZN(n404) );
  XNOR2_X1 U859 ( .A(n1), .B(n605), .ZN(n413) );
  NAND2_X1 U860 ( .A1(n203), .A2(n210), .ZN(n88) );
  XNOR2_X1 U861 ( .A(a[9]), .B(a[10]), .ZN(n502) );
  NAND2_X1 U862 ( .A1(n594), .A2(n73), .ZN(n9) );
  INV_X1 U863 ( .A(n73), .ZN(n71) );
  NAND2_X1 U864 ( .A1(n189), .A2(n194), .ZN(n73) );
  NOR2_X1 U865 ( .A1(n63), .A2(n58), .ZN(n56) );
  INV_X1 U866 ( .A(n63), .ZN(n61) );
  NAND2_X1 U867 ( .A1(n594), .A2(n593), .ZN(n63) );
  AOI21_X1 U868 ( .B1(n591), .B2(n27), .A(n28), .ZN(n26) );
  OAI21_X1 U869 ( .B1(n138), .B2(n140), .A(n139), .ZN(n137) );
  OAI22_X1 U870 ( .A1(n476), .A2(n488), .B1(n440), .B2(n482), .ZN(n302) );
  INV_X1 U871 ( .A(n494), .ZN(n488) );
  OAI21_X1 U872 ( .B1(n126), .B2(n128), .A(n127), .ZN(n125) );
  INV_X1 U873 ( .A(n147), .ZN(n145) );
  XNOR2_X1 U874 ( .A(n1), .B(n495), .ZN(n452) );
  AND2_X1 U875 ( .A1(n572), .A2(a[0]), .ZN(product[0]) );
  XNOR2_X1 U876 ( .A(n23), .B(n145), .ZN(product[2]) );
  NAND2_X1 U877 ( .A1(n597), .A2(n144), .ZN(n23) );
  XOR2_X1 U878 ( .A(n21), .B(n136), .Z(product[4]) );
  NAND2_X1 U879 ( .A1(n166), .A2(n135), .ZN(n21) );
  XOR2_X1 U880 ( .A(n22), .B(n140), .Z(product[3]) );
  NAND2_X1 U881 ( .A1(n167), .A2(n139), .ZN(n22) );
  XOR2_X1 U882 ( .A(n19), .B(n564), .Z(product[6]) );
  NAND2_X1 U883 ( .A1(n164), .A2(n127), .ZN(n19) );
  XNOR2_X1 U884 ( .A(n20), .B(n133), .ZN(product[5]) );
  NAND2_X1 U885 ( .A1(n596), .A2(n132), .ZN(n20) );
  NAND2_X1 U886 ( .A1(n163), .A2(n123), .ZN(n18) );
  XOR2_X1 U887 ( .A(n116), .B(n16), .Z(product[9]) );
  NAND2_X1 U888 ( .A1(n161), .A2(n115), .ZN(n16) );
  INV_X1 U889 ( .A(n125), .ZN(n124) );
  XNOR2_X1 U890 ( .A(n121), .B(n17), .ZN(product[8]) );
  OAI21_X1 U891 ( .B1(n124), .B2(n122), .A(n123), .ZN(n121) );
  XOR2_X1 U892 ( .A(n112), .B(n15), .Z(product[10]) );
  INV_X1 U893 ( .A(n584), .ZN(n112) );
  XNOR2_X1 U894 ( .A(n103), .B(n13), .ZN(product[12]) );
  INV_X1 U895 ( .A(n104), .ZN(n103) );
  XNOR2_X1 U896 ( .A(n109), .B(n14), .ZN(product[11]) );
  OAI21_X1 U897 ( .B1(n112), .B2(n559), .A(n566), .ZN(n109) );
  XOR2_X1 U898 ( .A(n89), .B(n11), .Z(product[14]) );
  AOI21_X1 U899 ( .B1(n103), .B2(n90), .A(n91), .ZN(n89) );
  XOR2_X1 U900 ( .A(n98), .B(n12), .Z(product[13]) );
  AOI21_X1 U901 ( .B1(n103), .B2(n99), .A(n100), .ZN(n98) );
  XOR2_X1 U902 ( .A(n82), .B(n10), .Z(product[15]) );
  AOI21_X1 U903 ( .B1(n83), .B2(n103), .A(n84), .ZN(n82) );
  XOR2_X1 U904 ( .A(n35), .B(n4), .Z(product[21]) );
  AOI21_X1 U905 ( .B1(n571), .B2(n36), .A(n37), .ZN(n35) );
  AOI21_X1 U906 ( .B1(n591), .B2(n61), .A(n62), .ZN(n60) );
  XOR2_X1 U907 ( .A(n74), .B(n9), .Z(product[16]) );
  INV_X1 U908 ( .A(n75), .ZN(n74) );
  AOI21_X1 U909 ( .B1(n591), .B2(n56), .A(n57), .ZN(n51) );
  XOR2_X1 U910 ( .A(n69), .B(n8), .Z(product[17]) );
  AOI21_X1 U911 ( .B1(n75), .B2(n594), .A(n71), .ZN(n69) );
  XNOR2_X1 U912 ( .A(n42), .B(n5), .ZN(product[20]) );
  OAI21_X1 U913 ( .B1(n74), .B2(n43), .A(n44), .ZN(n42) );
  INV_X1 U914 ( .A(n26), .ZN(n148) );
  INV_X1 U915 ( .A(n25), .ZN(product[23]) );
endmodule


module datapath_DW_mult_tc_18 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n1, n4, n5, n6, n7, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n26, n28, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n43, n45, n46, n47, n48, n49, n50, n51, n52, n55,
         n56, n57, n58, n59, n60, n61, n65, n67, n68, n70, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n86, n87, n88, n89, n90,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n129, n131, n132, n133, n134, n135, n136, n137, n138, n139, n141,
         n143, n144, n146, n148, n149, n150, n151, n154, n159, n160, n161,
         n162, n163, n165, n166, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n285, n286,
         n288, n289, n290, n291, n292, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n465,
         n466, n467, n468, n469, n470, n472, n474, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n487, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n594, n595, n596;
  assign product[23] = n26;

  FA_X1 U193 ( .A(n304), .B(n175), .CI(n314), .CO(n171), .S(n172) );
  FA_X1 U194 ( .A(n176), .B(n315), .CI(n179), .CO(n173), .S(n174) );
  FA_X1 U196 ( .A(n183), .B(n327), .CI(n180), .CO(n177), .S(n178) );
  FA_X1 U197 ( .A(n305), .B(n185), .CI(n316), .CO(n179), .S(n180) );
  FA_X1 U198 ( .A(n184), .B(n191), .CI(n189), .CO(n181), .S(n182) );
  FA_X1 U199 ( .A(n317), .B(n306), .CI(n186), .CO(n183), .S(n184) );
  FA_X1 U201 ( .A(n195), .B(n192), .CI(n190), .CO(n187), .S(n188) );
  FA_X1 U202 ( .A(n338), .B(n328), .CI(n197), .CO(n189), .S(n190) );
  FA_X1 U203 ( .A(n307), .B(n199), .CI(n318), .CO(n191), .S(n192) );
  FA_X1 U204 ( .A(n203), .B(n198), .CI(n196), .CO(n193), .S(n194) );
  FA_X1 U205 ( .A(n207), .B(n200), .CI(n205), .CO(n195), .S(n196) );
  FA_X1 U206 ( .A(n339), .B(n308), .CI(n319), .CO(n197), .S(n198) );
  FA_X1 U208 ( .A(n211), .B(n206), .CI(n204), .CO(n201), .S(n202) );
  FA_X1 U209 ( .A(n213), .B(n215), .CI(n208), .CO(n203), .S(n204) );
  FA_X1 U210 ( .A(n351), .B(n329), .CI(n340), .CO(n205), .S(n206) );
  FA_X1 U211 ( .A(n309), .B(n217), .CI(n320), .CO(n207), .S(n208) );
  FA_X1 U212 ( .A(n221), .B(n214), .CI(n212), .CO(n209), .S(n210) );
  FA_X1 U213 ( .A(n216), .B(n225), .CI(n223), .CO(n211), .S(n212) );
  FA_X1 U214 ( .A(n218), .B(n341), .CI(n227), .CO(n213), .S(n214) );
  FA_X1 U215 ( .A(n310), .B(n330), .CI(n321), .CO(n215), .S(n216) );
  FA_X1 U217 ( .A(n231), .B(n224), .CI(n222), .CO(n219), .S(n220) );
  FA_X1 U218 ( .A(n226), .B(n235), .CI(n233), .CO(n221), .S(n222) );
  FA_X1 U219 ( .A(n237), .B(n311), .CI(n228), .CO(n223), .S(n224) );
  FA_X1 U220 ( .A(n342), .B(n363), .CI(n322), .CO(n225), .S(n226) );
  FA_X1 U223 ( .A(n241), .B(n234), .CI(n232), .CO(n229), .S(n230) );
  FA_X1 U224 ( .A(n243), .B(n245), .CI(n236), .CO(n231), .S(n232) );
  FA_X1 U225 ( .A(n323), .B(n312), .CI(n238), .CO(n233), .S(n234) );
  FA_X1 U226 ( .A(n297), .B(n353), .CI(n343), .CO(n235), .S(n236) );
  HA_X1 U227 ( .A(n332), .B(n364), .CO(n237), .S(n238) );
  FA_X1 U228 ( .A(n249), .B(n244), .CI(n242), .CO(n239), .S(n240) );
  FA_X1 U229 ( .A(n251), .B(n253), .CI(n246), .CO(n241), .S(n242) );
  FA_X1 U230 ( .A(n344), .B(n354), .CI(n324), .CO(n243), .S(n244) );
  FA_X1 U231 ( .A(n365), .B(n313), .CI(n333), .CO(n245), .S(n246) );
  FA_X1 U232 ( .A(n252), .B(n257), .CI(n250), .CO(n247), .S(n248) );
  FA_X1 U233 ( .A(n254), .B(n345), .CI(n259), .CO(n249), .S(n250) );
  FA_X1 U234 ( .A(n298), .B(n334), .CI(n325), .CO(n251), .S(n252) );
  HA_X1 U235 ( .A(n355), .B(n366), .CO(n253), .S(n254) );
  FA_X1 U237 ( .A(n335), .B(n346), .CI(n265), .CO(n257), .S(n258) );
  FA_X1 U238 ( .A(n367), .B(n326), .CI(n356), .CO(n259), .S(n260) );
  FA_X1 U239 ( .A(n269), .B(n266), .CI(n264), .CO(n261), .S(n262) );
  FA_X1 U240 ( .A(n336), .B(n299), .CI(n347), .CO(n263), .S(n264) );
  HA_X1 U241 ( .A(n357), .B(n368), .CO(n265), .S(n266) );
  FA_X1 U242 ( .A(n273), .B(n348), .CI(n270), .CO(n267), .S(n268) );
  FA_X1 U243 ( .A(n369), .B(n337), .CI(n358), .CO(n269), .S(n270) );
  FA_X1 U244 ( .A(n349), .B(n300), .CI(n274), .CO(n271), .S(n272) );
  HA_X1 U245 ( .A(n359), .B(n370), .CO(n273), .S(n274) );
  FA_X1 U246 ( .A(n371), .B(n350), .CI(n360), .CO(n275), .S(n276) );
  HA_X1 U247 ( .A(n301), .B(n372), .CO(n277), .S(n278) );
  CLKBUF_X3 U483 ( .A(a[7]), .Z(n491) );
  CLKBUF_X3 U484 ( .A(a[11]), .Z(n489) );
  OR2_X1 U485 ( .A1(n303), .A2(n169), .ZN(n558) );
  XNOR2_X1 U486 ( .A(n559), .B(n258), .ZN(n256) );
  XNOR2_X1 U487 ( .A(n260), .B(n263), .ZN(n559) );
  XNOR2_X1 U488 ( .A(n596), .B(n454), .ZN(n560) );
  BUF_X1 U489 ( .A(b[9]), .Z(n455) );
  OR2_X1 U490 ( .A1(n210), .A2(n219), .ZN(n561) );
  CLKBUF_X3 U491 ( .A(n502), .Z(n478) );
  BUF_X1 U492 ( .A(b[3]), .Z(n461) );
  INV_X1 U493 ( .A(n99), .ZN(n562) );
  BUF_X1 U494 ( .A(b[6]), .Z(n458) );
  OR2_X1 U495 ( .A1(n230), .A2(n239), .ZN(n563) );
  BUF_X1 U496 ( .A(n494), .Z(n594) );
  XNOR2_X1 U497 ( .A(a[9]), .B(a[10]), .ZN(n564) );
  BUF_X1 U498 ( .A(b[2]), .Z(n462) );
  CLKBUF_X3 U499 ( .A(b[0]), .Z(n1) );
  NOR2_X1 U500 ( .A1(n86), .A2(n79), .ZN(n565) );
  NOR2_X1 U501 ( .A1(n194), .A2(n201), .ZN(n566) );
  CLKBUF_X1 U502 ( .A(b[4]), .Z(n460) );
  CLKBUF_X1 U503 ( .A(n74), .Z(n567) );
  NAND2_X1 U504 ( .A1(n258), .A2(n260), .ZN(n568) );
  NAND2_X1 U505 ( .A1(n258), .A2(n263), .ZN(n569) );
  NAND2_X1 U506 ( .A1(n260), .A2(n263), .ZN(n570) );
  NAND3_X1 U507 ( .A1(n568), .A2(n569), .A3(n570), .ZN(n255) );
  OR2_X1 U508 ( .A1(n500), .A2(n445), .ZN(n571) );
  OR2_X1 U509 ( .A1(n444), .A2(n482), .ZN(n572) );
  NAND2_X1 U510 ( .A1(n571), .A2(n572), .ZN(n368) );
  BUF_X1 U511 ( .A(b[7]), .Z(n457) );
  BUF_X1 U512 ( .A(n87), .Z(n573) );
  OR2_X1 U513 ( .A1(n100), .A2(n582), .ZN(n574) );
  OR2_X1 U514 ( .A1(n202), .A2(n209), .ZN(n575) );
  INV_X1 U515 ( .A(n123), .ZN(n576) );
  OAI21_X1 U516 ( .B1(n115), .B2(n113), .A(n114), .ZN(n577) );
  CLKBUF_X3 U517 ( .A(b[10]), .Z(n454) );
  CLKBUF_X2 U518 ( .A(b[1]), .Z(n463) );
  CLKBUF_X3 U519 ( .A(b[5]), .Z(n459) );
  XNOR2_X1 U520 ( .A(n57), .B(n578), .ZN(product[18]) );
  AND2_X1 U521 ( .A1(n151), .A2(n56), .ZN(n578) );
  AOI21_X1 U522 ( .B1(n116), .B2(n576), .A(n117), .ZN(n579) );
  AOI21_X1 U523 ( .B1(n104), .B2(n577), .A(n105), .ZN(n580) );
  XNOR2_X1 U524 ( .A(n68), .B(n581), .ZN(product[17]) );
  AND2_X1 U525 ( .A1(n588), .A2(n67), .ZN(n581) );
  NOR2_X1 U526 ( .A1(n210), .A2(n219), .ZN(n582) );
  AOI21_X1 U527 ( .B1(n104), .B2(n577), .A(n105), .ZN(n583) );
  OAI21_X1 U528 ( .B1(n583), .B2(n75), .A(n76), .ZN(n584) );
  NOR2_X1 U529 ( .A1(n256), .A2(n261), .ZN(n585) );
  OR2_X1 U530 ( .A1(n188), .A2(n193), .ZN(n589) );
  XNOR2_X1 U531 ( .A(n73), .B(n586), .ZN(product[16]) );
  AND2_X1 U532 ( .A1(n589), .A2(n72), .ZN(n586) );
  AND2_X1 U533 ( .A1(n588), .A2(n46), .ZN(n587) );
  XOR2_X1 U534 ( .A(n123), .B(n19), .Z(product[7]) );
  NOR2_X1 U535 ( .A1(n256), .A2(n261), .ZN(n118) );
  OR2_X1 U536 ( .A1(n187), .A2(n182), .ZN(n588) );
  OR2_X1 U537 ( .A1(n373), .A2(n362), .ZN(n590) );
  OR2_X1 U538 ( .A1(n272), .A2(n275), .ZN(n591) );
  OR2_X1 U539 ( .A1(n374), .A2(n302), .ZN(n592) );
  BUF_X2 U540 ( .A(n501), .Z(n477) );
  BUF_X2 U541 ( .A(a[5]), .Z(n492) );
  BUF_X2 U542 ( .A(a[9]), .Z(n490) );
  AND2_X1 U543 ( .A1(n592), .A2(n146), .ZN(product[1]) );
  NOR2_X1 U544 ( .A1(n171), .A2(n170), .ZN(n32) );
  NAND2_X1 U545 ( .A1(n148), .A2(n33), .ZN(n5) );
  NAND2_X1 U546 ( .A1(n558), .A2(n30), .ZN(n4) );
  INV_X1 U547 ( .A(n30), .ZN(n28) );
  NAND2_X1 U548 ( .A1(n149), .A2(n38), .ZN(n6) );
  NAND2_X1 U549 ( .A1(n173), .A2(n172), .ZN(n38) );
  INV_X1 U550 ( .A(n32), .ZN(n148) );
  NAND2_X1 U551 ( .A1(n171), .A2(n170), .ZN(n33) );
  INV_X1 U552 ( .A(n37), .ZN(n149) );
  NOR2_X1 U553 ( .A1(n173), .A2(n172), .ZN(n37) );
  NAND2_X1 U554 ( .A1(n150), .A2(n49), .ZN(n7) );
  OR2_X1 U555 ( .A1(n1), .A2(n290), .ZN(n426) );
  NOR2_X1 U556 ( .A1(n60), .A2(n55), .ZN(n51) );
  NAND2_X1 U557 ( .A1(n589), .A2(n588), .ZN(n60) );
  NAND2_X1 U558 ( .A1(n174), .A2(n177), .ZN(n49) );
  BUF_X2 U559 ( .A(n506), .Z(n482) );
  OR2_X1 U560 ( .A1(n1), .A2(n484), .ZN(n400) );
  AND2_X1 U561 ( .A1(n1), .A2(n292), .ZN(n362) );
  OR2_X1 U562 ( .A1(n1), .A2(n485), .ZN(n413) );
  CLKBUF_X3 U563 ( .A(a[3]), .Z(n493) );
  OR2_X1 U564 ( .A1(n1), .A2(n487), .ZN(n439) );
  XNOR2_X1 U565 ( .A(n1), .B(n492), .ZN(n425) );
  NOR2_X1 U566 ( .A1(n178), .A2(n181), .ZN(n55) );
  AOI21_X1 U567 ( .B1(n70), .B2(n588), .A(n65), .ZN(n61) );
  BUF_X2 U568 ( .A(n496), .Z(n472) );
  INV_X1 U569 ( .A(n282), .ZN(n314) );
  AND2_X1 U570 ( .A1(n1), .A2(n283), .ZN(n326) );
  NOR2_X1 U571 ( .A1(n278), .A2(n361), .ZN(n137) );
  XNOR2_X1 U572 ( .A(n492), .B(n461), .ZN(n422) );
  BUF_X2 U573 ( .A(n504), .Z(n480) );
  XOR2_X1 U574 ( .A(a[10]), .B(a[11]), .Z(n465) );
  INV_X1 U575 ( .A(n575), .ZN(n84) );
  OAI22_X1 U576 ( .A1(n495), .A2(n376), .B1(n477), .B2(n375), .ZN(n169) );
  INV_X1 U577 ( .A(n279), .ZN(n303) );
  NAND2_X1 U578 ( .A1(n303), .A2(n169), .ZN(n30) );
  INV_X1 U579 ( .A(n169), .ZN(n170) );
  XNOR2_X1 U580 ( .A(a[7]), .B(a[8]), .ZN(n502) );
  OAI22_X1 U581 ( .A1(n495), .A2(n378), .B1(n477), .B2(n377), .ZN(n175) );
  AND2_X1 U582 ( .A1(n1), .A2(n280), .ZN(n313) );
  NAND2_X1 U583 ( .A1(n276), .A2(n277), .ZN(n134) );
  XNOR2_X1 U584 ( .A(n463), .B(n492), .ZN(n424) );
  NAND2_X1 U585 ( .A1(n154), .A2(n80), .ZN(n11) );
  BUF_X2 U586 ( .A(n505), .Z(n481) );
  NAND2_X2 U587 ( .A1(n467), .A2(n503), .ZN(n497) );
  XNOR2_X1 U588 ( .A(n492), .B(n456), .ZN(n417) );
  CLKBUF_X1 U589 ( .A(b[8]), .Z(n456) );
  XNOR2_X1 U590 ( .A(n492), .B(n460), .ZN(n421) );
  NAND2_X2 U591 ( .A1(n469), .A2(n505), .ZN(n499) );
  XNOR2_X1 U592 ( .A(n492), .B(n455), .ZN(n416) );
  XNOR2_X1 U593 ( .A(n492), .B(n458), .ZN(n419) );
  NAND2_X2 U594 ( .A1(n470), .A2(n506), .ZN(n500) );
  OR2_X1 U595 ( .A1(n1), .A2(n296), .ZN(n452) );
  OAI22_X1 U596 ( .A1(n500), .A2(n296), .B1(n452), .B2(n482), .ZN(n302) );
  NAND2_X1 U597 ( .A1(n561), .A2(n96), .ZN(n13) );
  INV_X1 U598 ( .A(n72), .ZN(n70) );
  NAND2_X1 U599 ( .A1(n188), .A2(n193), .ZN(n72) );
  INV_X1 U600 ( .A(n92), .ZN(n90) );
  NAND2_X1 U601 ( .A1(n248), .A2(n255), .ZN(n114) );
  NOR2_X1 U602 ( .A1(n248), .A2(n255), .ZN(n113) );
  XNOR2_X1 U603 ( .A(n492), .B(n457), .ZN(n418) );
  AOI21_X1 U604 ( .B1(n500), .B2(n482), .A(n440), .ZN(n294) );
  INV_X1 U605 ( .A(n143), .ZN(n141) );
  NAND2_X1 U606 ( .A1(n262), .A2(n267), .ZN(n122) );
  NOR2_X1 U607 ( .A1(n262), .A2(n267), .ZN(n121) );
  INV_X1 U608 ( .A(n133), .ZN(n165) );
  NOR2_X1 U609 ( .A1(n276), .A2(n277), .ZN(n133) );
  OAI22_X1 U610 ( .A1(n429), .A2(n499), .B1(n428), .B2(n481), .ZN(n352) );
  INV_X1 U611 ( .A(n61), .ZN(n59) );
  INV_X1 U612 ( .A(n60), .ZN(n58) );
  INV_X1 U613 ( .A(n55), .ZN(n151) );
  OAI21_X1 U614 ( .B1(n61), .B2(n55), .A(n56), .ZN(n52) );
  NAND2_X1 U615 ( .A1(n178), .A2(n181), .ZN(n56) );
  XNOR2_X1 U616 ( .A(n492), .B(n459), .ZN(n420) );
  NAND2_X1 U617 ( .A1(n161), .A2(n119), .ZN(n18) );
  INV_X1 U618 ( .A(n125), .ZN(n163) );
  NOR2_X1 U619 ( .A1(n268), .A2(n271), .ZN(n125) );
  BUF_X1 U620 ( .A(n494), .Z(n595) );
  OR2_X1 U621 ( .A1(n1), .A2(n281), .ZN(n387) );
  NAND2_X1 U622 ( .A1(n210), .A2(n219), .ZN(n96) );
  NOR2_X1 U623 ( .A1(n240), .A2(n247), .ZN(n109) );
  NOR2_X1 U624 ( .A1(n210), .A2(n219), .ZN(n95) );
  INV_X1 U625 ( .A(n574), .ZN(n89) );
  NOR2_X1 U626 ( .A1(n574), .A2(n84), .ZN(n82) );
  OAI22_X1 U627 ( .A1(n500), .A2(n446), .B1(n445), .B2(n482), .ZN(n369) );
  NAND2_X1 U628 ( .A1(n256), .A2(n261), .ZN(n119) );
  INV_X1 U629 ( .A(n146), .ZN(n144) );
  INV_X1 U630 ( .A(n94), .ZN(n92) );
  OAI21_X1 U631 ( .B1(n95), .B2(n101), .A(n96), .ZN(n94) );
  NAND2_X1 U632 ( .A1(n268), .A2(n271), .ZN(n126) );
  INV_X1 U633 ( .A(n480), .ZN(n289) );
  OAI22_X1 U634 ( .A1(n474), .A2(n425), .B1(n424), .B2(n480), .ZN(n349) );
  OAI22_X1 U635 ( .A1(n474), .A2(n424), .B1(n423), .B2(n480), .ZN(n348) );
  OAI22_X1 U636 ( .A1(n474), .A2(n423), .B1(n422), .B2(n480), .ZN(n347) );
  OAI22_X1 U637 ( .A1(n474), .A2(n422), .B1(n421), .B2(n480), .ZN(n346) );
  OAI22_X1 U638 ( .A1(n474), .A2(n421), .B1(n420), .B2(n480), .ZN(n345) );
  OAI22_X1 U639 ( .A1(n474), .A2(n418), .B1(n417), .B2(n480), .ZN(n342) );
  OAI22_X1 U640 ( .A1(n474), .A2(n417), .B1(n416), .B2(n480), .ZN(n341) );
  OAI22_X1 U641 ( .A1(n474), .A2(n416), .B1(n415), .B2(n480), .ZN(n340) );
  AOI21_X1 U642 ( .B1(n474), .B2(n480), .A(n414), .ZN(n288) );
  OAI22_X1 U643 ( .A1(n474), .A2(n290), .B1(n426), .B2(n480), .ZN(n300) );
  BUF_X2 U644 ( .A(n498), .Z(n474) );
  AND2_X1 U645 ( .A1(n1), .A2(n289), .ZN(n350) );
  INV_X1 U646 ( .A(n288), .ZN(n338) );
  NOR2_X1 U647 ( .A1(n100), .A2(n582), .ZN(n93) );
  BUF_X2 U648 ( .A(n494), .Z(n596) );
  XNOR2_X1 U649 ( .A(n594), .B(n458), .ZN(n445) );
  XNOR2_X1 U650 ( .A(n461), .B(n595), .ZN(n448) );
  XNOR2_X1 U651 ( .A(n457), .B(n596), .ZN(n444) );
  XNOR2_X1 U652 ( .A(n459), .B(n596), .ZN(n446) );
  OAI22_X1 U653 ( .A1(n500), .A2(n444), .B1(n443), .B2(n482), .ZN(n367) );
  OAI22_X1 U654 ( .A1(n500), .A2(n448), .B1(n447), .B2(n482), .ZN(n371) );
  OAI22_X1 U655 ( .A1(n500), .A2(n447), .B1(n446), .B2(n482), .ZN(n370) );
  XNOR2_X1 U656 ( .A(n456), .B(n494), .ZN(n443) );
  XNOR2_X1 U657 ( .A(n460), .B(n494), .ZN(n447) );
  BUF_X2 U658 ( .A(a[1]), .Z(n494) );
  INV_X1 U659 ( .A(n175), .ZN(n176) );
  INV_X1 U660 ( .A(n479), .ZN(n286) );
  OAI22_X1 U661 ( .A1(n411), .A2(n479), .B1(n497), .B2(n412), .ZN(n336) );
  OAI22_X1 U662 ( .A1(n497), .A2(n409), .B1(n479), .B2(n408), .ZN(n333) );
  OAI22_X1 U663 ( .A1(n497), .A2(n406), .B1(n479), .B2(n405), .ZN(n330) );
  OAI22_X1 U664 ( .A1(n497), .A2(n405), .B1(n479), .B2(n404), .ZN(n329) );
  OAI22_X1 U665 ( .A1(n497), .A2(n403), .B1(n479), .B2(n402), .ZN(n328) );
  AOI21_X1 U666 ( .B1(n497), .B2(n479), .A(n401), .ZN(n285) );
  OAI22_X1 U667 ( .A1(n497), .A2(n485), .B1(n413), .B2(n479), .ZN(n299) );
  CLKBUF_X3 U668 ( .A(n503), .Z(n479) );
  AND2_X1 U669 ( .A1(n1), .A2(n286), .ZN(n337) );
  INV_X1 U670 ( .A(n285), .ZN(n327) );
  INV_X1 U671 ( .A(n131), .ZN(n129) );
  OAI21_X1 U672 ( .B1(n133), .B2(n135), .A(n134), .ZN(n132) );
  NOR2_X1 U673 ( .A1(n40), .A2(n37), .ZN(n35) );
  NAND2_X1 U674 ( .A1(n589), .A2(n587), .ZN(n40) );
  INV_X1 U675 ( .A(n79), .ZN(n154) );
  NOR2_X1 U676 ( .A1(n194), .A2(n201), .ZN(n79) );
  INV_X1 U677 ( .A(n136), .ZN(n135) );
  INV_X1 U678 ( .A(n67), .ZN(n65) );
  INV_X1 U679 ( .A(n137), .ZN(n166) );
  NAND2_X1 U680 ( .A1(n187), .A2(n182), .ZN(n67) );
  NAND2_X1 U681 ( .A1(n272), .A2(n275), .ZN(n131) );
  INV_X1 U682 ( .A(n121), .ZN(n162) );
  OAI22_X1 U683 ( .A1(n474), .A2(n415), .B1(n414), .B2(n480), .ZN(n339) );
  NOR2_X1 U684 ( .A1(n86), .A2(n79), .ZN(n77) );
  NAND2_X1 U685 ( .A1(n575), .A2(n573), .ZN(n12) );
  OAI21_X1 U686 ( .B1(n87), .B2(n566), .A(n80), .ZN(n78) );
  OAI21_X1 U687 ( .B1(n92), .B2(n84), .A(n573), .ZN(n83) );
  NOR2_X1 U688 ( .A1(n202), .A2(n209), .ZN(n86) );
  NAND2_X1 U689 ( .A1(n373), .A2(n362), .ZN(n143) );
  OAI22_X1 U690 ( .A1(n449), .A2(n482), .B1(n450), .B2(n500), .ZN(n373) );
  OAI22_X1 U691 ( .A1(n449), .A2(n500), .B1(n448), .B2(n482), .ZN(n372) );
  NAND2_X1 U692 ( .A1(n194), .A2(n201), .ZN(n80) );
  INV_X1 U693 ( .A(n48), .ZN(n150) );
  NOR2_X1 U694 ( .A1(n174), .A2(n177), .ZN(n48) );
  XNOR2_X1 U695 ( .A(n463), .B(n596), .ZN(n450) );
  NAND2_X1 U696 ( .A1(n202), .A2(n209), .ZN(n87) );
  AOI21_X1 U697 ( .B1(n591), .B2(n132), .A(n129), .ZN(n127) );
  OAI21_X1 U698 ( .B1(n34), .B2(n32), .A(n33), .ZN(n31) );
  OAI21_X1 U699 ( .B1(n106), .B2(n110), .A(n107), .ZN(n105) );
  NOR2_X1 U700 ( .A1(n106), .A2(n109), .ZN(n104) );
  NAND2_X1 U701 ( .A1(n563), .A2(n107), .ZN(n15) );
  NOR2_X1 U702 ( .A1(n230), .A2(n239), .ZN(n106) );
  OAI21_X1 U703 ( .B1(n583), .B2(n75), .A(n76), .ZN(n74) );
  NAND2_X1 U704 ( .A1(n77), .A2(n93), .ZN(n75) );
  AOI21_X1 U705 ( .B1(n94), .B2(n565), .A(n78), .ZN(n76) );
  NAND2_X1 U706 ( .A1(n230), .A2(n239), .ZN(n107) );
  OAI22_X1 U707 ( .A1(n474), .A2(n420), .B1(n419), .B2(n480), .ZN(n344) );
  XNOR2_X1 U708 ( .A(a[3]), .B(a[4]), .ZN(n504) );
  INV_X1 U709 ( .A(n100), .ZN(n98) );
  NAND2_X1 U710 ( .A1(n98), .A2(n562), .ZN(n14) );
  INV_X1 U711 ( .A(n101), .ZN(n99) );
  NOR2_X1 U712 ( .A1(n220), .A2(n229), .ZN(n100) );
  NAND2_X1 U713 ( .A1(n159), .A2(n110), .ZN(n16) );
  INV_X1 U714 ( .A(n109), .ZN(n159) );
  OAI21_X1 U715 ( .B1(n115), .B2(n113), .A(n114), .ZN(n112) );
  AOI21_X1 U716 ( .B1(n116), .B2(n124), .A(n117), .ZN(n115) );
  NAND2_X1 U717 ( .A1(n220), .A2(n229), .ZN(n101) );
  OAI22_X1 U718 ( .A1(n500), .A2(n443), .B1(n442), .B2(n482), .ZN(n366) );
  OAI21_X1 U719 ( .B1(n41), .B2(n37), .A(n38), .ZN(n36) );
  AOI21_X1 U720 ( .B1(n587), .B2(n70), .A(n43), .ZN(n41) );
  OAI22_X1 U721 ( .A1(n497), .A2(n407), .B1(n479), .B2(n406), .ZN(n331) );
  NAND2_X1 U722 ( .A1(n240), .A2(n247), .ZN(n110) );
  XNOR2_X1 U723 ( .A(n462), .B(n596), .ZN(n449) );
  XNOR2_X1 U724 ( .A(n462), .B(n492), .ZN(n423) );
  AOI21_X1 U725 ( .B1(n472), .B2(n478), .A(n388), .ZN(n282) );
  OAI22_X1 U726 ( .A1(n472), .A2(n389), .B1(n388), .B2(n478), .ZN(n315) );
  OAI22_X1 U727 ( .A1(n472), .A2(n390), .B1(n389), .B2(n478), .ZN(n316) );
  OAI22_X1 U728 ( .A1(n472), .A2(n392), .B1(n391), .B2(n478), .ZN(n318) );
  OAI22_X1 U729 ( .A1(n472), .A2(n391), .B1(n390), .B2(n478), .ZN(n317) );
  OAI22_X1 U730 ( .A1(n472), .A2(n397), .B1(n396), .B2(n478), .ZN(n323) );
  OAI22_X1 U731 ( .A1(n472), .A2(n394), .B1(n393), .B2(n478), .ZN(n320) );
  OAI22_X1 U732 ( .A1(n472), .A2(n393), .B1(n392), .B2(n478), .ZN(n319) );
  OAI22_X1 U733 ( .A1(n472), .A2(n395), .B1(n394), .B2(n478), .ZN(n321) );
  INV_X1 U734 ( .A(n478), .ZN(n283) );
  OAI22_X1 U735 ( .A1(n472), .A2(n484), .B1(n400), .B2(n478), .ZN(n298) );
  OAI22_X1 U736 ( .A1(n472), .A2(n396), .B1(n395), .B2(n478), .ZN(n322) );
  INV_X1 U737 ( .A(n585), .ZN(n161) );
  OAI22_X1 U738 ( .A1(n472), .A2(n399), .B1(n398), .B2(n478), .ZN(n325) );
  OAI22_X1 U739 ( .A1(n472), .A2(n398), .B1(n397), .B2(n478), .ZN(n324) );
  OAI22_X1 U740 ( .A1(n500), .A2(n441), .B1(n440), .B2(n482), .ZN(n364) );
  XNOR2_X1 U741 ( .A(n453), .B(n594), .ZN(n440) );
  XNOR2_X1 U742 ( .A(n492), .B(n453), .ZN(n414) );
  BUF_X2 U743 ( .A(b[11]), .Z(n453) );
  OAI22_X1 U744 ( .A1(n497), .A2(n408), .B1(n479), .B2(n407), .ZN(n332) );
  NAND2_X1 U745 ( .A1(n468), .A2(n504), .ZN(n498) );
  XOR2_X1 U746 ( .A(a[5]), .B(a[4]), .Z(n468) );
  XNOR2_X1 U747 ( .A(n596), .B(n454), .ZN(n441) );
  XNOR2_X1 U748 ( .A(n492), .B(n454), .ZN(n415) );
  XOR2_X1 U749 ( .A(a[1]), .B(a[0]), .Z(n470) );
  OAI22_X1 U750 ( .A1(n474), .A2(n419), .B1(n418), .B2(n480), .ZN(n343) );
  NAND2_X1 U751 ( .A1(n466), .A2(n502), .ZN(n496) );
  XOR2_X1 U752 ( .A(a[9]), .B(a[8]), .Z(n466) );
  OAI22_X1 U753 ( .A1(n410), .A2(n479), .B1(n411), .B2(n497), .ZN(n335) );
  OAI22_X1 U754 ( .A1(n410), .A2(n497), .B1(n479), .B2(n409), .ZN(n334) );
  INV_X1 U755 ( .A(n113), .ZN(n160) );
  OAI22_X1 U756 ( .A1(n500), .A2(n442), .B1(n560), .B2(n482), .ZN(n365) );
  XNOR2_X1 U757 ( .A(n595), .B(n455), .ZN(n442) );
  INV_X1 U758 ( .A(n294), .ZN(n363) );
  OAI22_X1 U759 ( .A1(n495), .A2(n483), .B1(n387), .B2(n477), .ZN(n297) );
  OAI22_X1 U760 ( .A1(n495), .A2(n382), .B1(n477), .B2(n381), .ZN(n308) );
  OAI22_X1 U761 ( .A1(n495), .A2(n380), .B1(n477), .B2(n379), .ZN(n306) );
  OAI22_X1 U762 ( .A1(n384), .A2(n477), .B1(n385), .B2(n495), .ZN(n311) );
  OAI22_X1 U763 ( .A1(n495), .A2(n379), .B1(n477), .B2(n378), .ZN(n305) );
  OAI22_X1 U764 ( .A1(n495), .A2(n377), .B1(n477), .B2(n376), .ZN(n304) );
  AOI21_X1 U765 ( .B1(n495), .B2(n477), .A(n375), .ZN(n279) );
  OAI22_X1 U766 ( .A1(n495), .A2(n381), .B1(n477), .B2(n380), .ZN(n307) );
  OAI22_X1 U767 ( .A1(n385), .A2(n477), .B1(n495), .B2(n386), .ZN(n312) );
  OAI22_X1 U768 ( .A1(n495), .A2(n383), .B1(n477), .B2(n382), .ZN(n309) );
  OAI22_X1 U769 ( .A1(n384), .A2(n495), .B1(n477), .B2(n383), .ZN(n310) );
  INV_X1 U770 ( .A(n501), .ZN(n280) );
  XNOR2_X1 U771 ( .A(a[9]), .B(a[10]), .ZN(n501) );
  NAND2_X2 U772 ( .A1(n465), .A2(n564), .ZN(n495) );
  AOI21_X1 U773 ( .B1(n46), .B2(n65), .A(n47), .ZN(n45) );
  OAI21_X1 U774 ( .B1(n56), .B2(n48), .A(n49), .ZN(n47) );
  NOR2_X1 U775 ( .A1(n55), .A2(n48), .ZN(n46) );
  INV_X1 U776 ( .A(n45), .ZN(n43) );
  OAI22_X1 U777 ( .A1(n497), .A2(n402), .B1(n479), .B2(n401), .ZN(n185) );
  INV_X1 U778 ( .A(n185), .ZN(n186) );
  OAI21_X1 U779 ( .B1(n139), .B2(n137), .A(n138), .ZN(n136) );
  AOI21_X1 U780 ( .B1(n590), .B2(n144), .A(n141), .ZN(n139) );
  INV_X1 U781 ( .A(n481), .ZN(n292) );
  OAI22_X1 U782 ( .A1(n437), .A2(n481), .B1(n499), .B2(n438), .ZN(n361) );
  OAI22_X1 U783 ( .A1(n436), .A2(n481), .B1(n437), .B2(n499), .ZN(n360) );
  OAI22_X1 U784 ( .A1(n436), .A2(n499), .B1(n435), .B2(n481), .ZN(n359) );
  OAI22_X1 U785 ( .A1(n499), .A2(n435), .B1(n434), .B2(n481), .ZN(n358) );
  OAI22_X1 U786 ( .A1(n499), .A2(n434), .B1(n433), .B2(n481), .ZN(n357) );
  OAI22_X1 U787 ( .A1(n499), .A2(n433), .B1(n432), .B2(n481), .ZN(n356) );
  OAI22_X1 U788 ( .A1(n499), .A2(n432), .B1(n431), .B2(n481), .ZN(n355) );
  OAI22_X1 U789 ( .A1(n499), .A2(n431), .B1(n430), .B2(n481), .ZN(n354) );
  OAI22_X1 U790 ( .A1(n499), .A2(n430), .B1(n429), .B2(n481), .ZN(n353) );
  AOI21_X1 U791 ( .B1(n499), .B2(n481), .A(n427), .ZN(n291) );
  NAND2_X1 U792 ( .A1(n278), .A2(n361), .ZN(n138) );
  OR2_X1 U793 ( .A1(n352), .A2(n331), .ZN(n227) );
  XNOR2_X1 U794 ( .A(n331), .B(n352), .ZN(n228) );
  INV_X1 U795 ( .A(n291), .ZN(n351) );
  XNOR2_X1 U796 ( .A(n463), .B(n493), .ZN(n437) );
  XNOR2_X1 U797 ( .A(n1), .B(n493), .ZN(n438) );
  XNOR2_X1 U798 ( .A(n493), .B(n458), .ZN(n432) );
  XNOR2_X1 U799 ( .A(n493), .B(n457), .ZN(n431) );
  XNOR2_X1 U800 ( .A(n460), .B(n493), .ZN(n434) );
  XNOR2_X1 U801 ( .A(n493), .B(n459), .ZN(n433) );
  XNOR2_X1 U802 ( .A(n462), .B(n493), .ZN(n436) );
  XNOR2_X1 U803 ( .A(n493), .B(n456), .ZN(n430) );
  XNOR2_X1 U804 ( .A(n461), .B(n493), .ZN(n435) );
  XNOR2_X1 U805 ( .A(n493), .B(n455), .ZN(n429) );
  XNOR2_X1 U806 ( .A(n493), .B(n454), .ZN(n428) );
  XNOR2_X1 U807 ( .A(n493), .B(n453), .ZN(n427) );
  INV_X1 U808 ( .A(n492), .ZN(n290) );
  OAI22_X1 U809 ( .A1(n497), .A2(n404), .B1(n479), .B2(n403), .ZN(n199) );
  INV_X1 U810 ( .A(n199), .ZN(n200) );
  XNOR2_X1 U811 ( .A(a[5]), .B(a[6]), .ZN(n503) );
  XNOR2_X1 U812 ( .A(n490), .B(n453), .ZN(n388) );
  XNOR2_X1 U813 ( .A(n490), .B(n456), .ZN(n391) );
  XNOR2_X1 U814 ( .A(n490), .B(n454), .ZN(n389) );
  XNOR2_X1 U815 ( .A(n490), .B(n455), .ZN(n390) );
  XNOR2_X1 U816 ( .A(n490), .B(n457), .ZN(n392) );
  INV_X1 U817 ( .A(n490), .ZN(n484) );
  XNOR2_X1 U818 ( .A(n1), .B(n490), .ZN(n399) );
  XNOR2_X1 U819 ( .A(n462), .B(n490), .ZN(n397) );
  XNOR2_X1 U820 ( .A(n463), .B(n490), .ZN(n398) );
  XNOR2_X1 U821 ( .A(n490), .B(n461), .ZN(n396) );
  XNOR2_X1 U822 ( .A(n490), .B(n458), .ZN(n393) );
  XNOR2_X1 U823 ( .A(n490), .B(n460), .ZN(n395) );
  XNOR2_X1 U824 ( .A(n490), .B(n459), .ZN(n394) );
  INV_X1 U825 ( .A(n491), .ZN(n485) );
  XNOR2_X1 U826 ( .A(n1), .B(n491), .ZN(n412) );
  XNOR2_X1 U827 ( .A(n463), .B(n491), .ZN(n411) );
  XNOR2_X1 U828 ( .A(n462), .B(n491), .ZN(n410) );
  XNOR2_X1 U829 ( .A(n461), .B(n491), .ZN(n409) );
  XNOR2_X1 U830 ( .A(n491), .B(n457), .ZN(n405) );
  XNOR2_X1 U831 ( .A(n460), .B(n491), .ZN(n408) );
  XNOR2_X1 U832 ( .A(n491), .B(n459), .ZN(n407) );
  XNOR2_X1 U833 ( .A(n491), .B(n458), .ZN(n406) );
  XNOR2_X1 U834 ( .A(n491), .B(n454), .ZN(n402) );
  XNOR2_X1 U835 ( .A(n491), .B(n453), .ZN(n401) );
  XNOR2_X1 U836 ( .A(n491), .B(n456), .ZN(n404) );
  XNOR2_X1 U837 ( .A(n491), .B(n455), .ZN(n403) );
  XOR2_X1 U838 ( .A(a[7]), .B(a[6]), .Z(n467) );
  OAI21_X1 U839 ( .B1(n118), .B2(n122), .A(n119), .ZN(n117) );
  NOR2_X1 U840 ( .A1(n585), .A2(n121), .ZN(n116) );
  XNOR2_X1 U841 ( .A(n489), .B(n454), .ZN(n376) );
  XNOR2_X1 U842 ( .A(n453), .B(n489), .ZN(n375) );
  XNOR2_X1 U843 ( .A(n489), .B(n458), .ZN(n380) );
  XNOR2_X1 U844 ( .A(n489), .B(n457), .ZN(n379) );
  XNOR2_X1 U845 ( .A(n489), .B(n459), .ZN(n381) );
  XNOR2_X1 U846 ( .A(n1), .B(n489), .ZN(n386) );
  INV_X1 U847 ( .A(n489), .ZN(n483) );
  XNOR2_X1 U848 ( .A(n463), .B(n489), .ZN(n385) );
  XNOR2_X1 U849 ( .A(n489), .B(n456), .ZN(n378) );
  XNOR2_X1 U850 ( .A(n489), .B(n455), .ZN(n377) );
  XNOR2_X1 U851 ( .A(n462), .B(n489), .ZN(n384) );
  XNOR2_X1 U852 ( .A(n460), .B(n489), .ZN(n382) );
  INV_X1 U853 ( .A(n489), .ZN(n281) );
  XNOR2_X1 U854 ( .A(n461), .B(n489), .ZN(n383) );
  INV_X1 U855 ( .A(n595), .ZN(n296) );
  OAI22_X1 U856 ( .A1(n499), .A2(n428), .B1(n427), .B2(n481), .ZN(n217) );
  INV_X1 U857 ( .A(n217), .ZN(n218) );
  XNOR2_X1 U858 ( .A(a[1]), .B(a[2]), .ZN(n505) );
  INV_X1 U859 ( .A(a[0]), .ZN(n506) );
  OAI22_X1 U860 ( .A1(n499), .A2(n487), .B1(n439), .B2(n481), .ZN(n301) );
  INV_X1 U861 ( .A(n493), .ZN(n487) );
  XNOR2_X1 U862 ( .A(n1), .B(n595), .ZN(n451) );
  XOR2_X1 U863 ( .A(a[3]), .B(a[2]), .Z(n469) );
  NAND2_X1 U864 ( .A1(n302), .A2(n374), .ZN(n146) );
  OAI22_X1 U865 ( .A1(n450), .A2(n482), .B1(n500), .B2(n451), .ZN(n374) );
  OAI21_X1 U866 ( .B1(n125), .B2(n127), .A(n126), .ZN(n124) );
  AND2_X1 U867 ( .A1(n1), .A2(n295), .ZN(product[0]) );
  INV_X1 U868 ( .A(n482), .ZN(n295) );
  XNOR2_X1 U869 ( .A(n24), .B(n144), .ZN(product[2]) );
  NAND2_X1 U870 ( .A1(n590), .A2(n143), .ZN(n24) );
  XOR2_X1 U871 ( .A(n22), .B(n135), .Z(product[4]) );
  NAND2_X1 U872 ( .A1(n165), .A2(n134), .ZN(n22) );
  XOR2_X1 U873 ( .A(n23), .B(n139), .Z(product[3]) );
  NAND2_X1 U874 ( .A1(n166), .A2(n138), .ZN(n23) );
  XNOR2_X1 U875 ( .A(n21), .B(n132), .ZN(product[5]) );
  NAND2_X1 U876 ( .A1(n591), .A2(n131), .ZN(n21) );
  XOR2_X1 U877 ( .A(n20), .B(n127), .Z(product[6]) );
  NAND2_X1 U878 ( .A1(n163), .A2(n126), .ZN(n20) );
  XOR2_X1 U879 ( .A(n579), .B(n17), .Z(product[9]) );
  NAND2_X1 U880 ( .A1(n160), .A2(n114), .ZN(n17) );
  NAND2_X1 U881 ( .A1(n162), .A2(n122), .ZN(n19) );
  INV_X1 U882 ( .A(n124), .ZN(n123) );
  XNOR2_X1 U883 ( .A(n120), .B(n18), .ZN(product[8]) );
  OAI21_X1 U884 ( .B1(n123), .B2(n121), .A(n122), .ZN(n120) );
  XOR2_X1 U885 ( .A(n111), .B(n16), .Z(product[10]) );
  INV_X1 U886 ( .A(n112), .ZN(n111) );
  XNOR2_X1 U887 ( .A(n102), .B(n14), .ZN(product[12]) );
  INV_X1 U888 ( .A(n580), .ZN(n102) );
  XNOR2_X1 U889 ( .A(n108), .B(n15), .ZN(product[11]) );
  OAI21_X1 U890 ( .B1(n111), .B2(n109), .A(n110), .ZN(n108) );
  XOR2_X1 U891 ( .A(n88), .B(n12), .Z(product[14]) );
  AOI21_X1 U892 ( .B1(n102), .B2(n89), .A(n90), .ZN(n88) );
  XOR2_X1 U893 ( .A(n97), .B(n13), .Z(product[13]) );
  AOI21_X1 U894 ( .B1(n102), .B2(n98), .A(n99), .ZN(n97) );
  XOR2_X1 U895 ( .A(n81), .B(n11), .Z(product[15]) );
  AOI21_X1 U896 ( .B1(n82), .B2(n102), .A(n83), .ZN(n81) );
  AOI21_X1 U897 ( .B1(n31), .B2(n558), .A(n28), .ZN(n26) );
  XOR2_X1 U898 ( .A(n34), .B(n5), .Z(product[21]) );
  AOI21_X1 U899 ( .B1(n74), .B2(n35), .A(n36), .ZN(n34) );
  AOI21_X1 U900 ( .B1(n584), .B2(n58), .A(n59), .ZN(n57) );
  XOR2_X1 U901 ( .A(n50), .B(n7), .Z(product[19]) );
  AOI21_X1 U902 ( .B1(n567), .B2(n51), .A(n52), .ZN(n50) );
  INV_X1 U903 ( .A(n584), .ZN(n73) );
  AOI21_X1 U904 ( .B1(n74), .B2(n589), .A(n70), .ZN(n68) );
  XNOR2_X1 U905 ( .A(n39), .B(n6), .ZN(product[20]) );
  OAI21_X1 U906 ( .B1(n73), .B2(n40), .A(n41), .ZN(n39) );
  XNOR2_X1 U907 ( .A(n31), .B(n4), .ZN(product[22]) );
endmodule


module datapath_DW_mult_tc_19 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n1, n4, n5, n6, n10, n11, n12, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n25, n26, n27, n28, n29, n30, n31, n32, n33, n35, n37, n38,
         n39, n40, n41, n42, n43, n44, n46, n48, n49, n50, n51, n52, n55, n57,
         n58, n62, n63, n64, n65, n66, n68, n70, n71, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n89, n90, n91, n93, n94,
         n95, n96, n97, n98, n99, n100, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n132, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n144, n146, n147, n149, n150, n151, n157, n158, n159, n160, n162,
         n163, n164, n165, n166, n168, n169, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n285, n286, n287,
         n288, n289, n291, n292, n294, n295, n297, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n464, n465, n466, n468, n469, n470,
         n471, n472, n473, n480, n481, n482, n483, n484, n485, n486, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n561,
         n562, n563, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601;

  FA_X1 U5 ( .A(n306), .B(n172), .CI(n150), .CO(n25), .S(product[22]) );
  FA_X1 U195 ( .A(n307), .B(n178), .CI(n315), .CO(n174), .S(n175) );
  FA_X1 U196 ( .A(n179), .B(n316), .CI(n182), .CO(n176), .S(n177) );
  FA_X1 U198 ( .A(n186), .B(n328), .CI(n183), .CO(n180), .S(n181) );
  FA_X1 U199 ( .A(n308), .B(n188), .CI(n317), .CO(n182), .S(n183) );
  FA_X1 U200 ( .A(n187), .B(n194), .CI(n192), .CO(n184), .S(n185) );
  FA_X1 U201 ( .A(n329), .B(n318), .CI(n189), .CO(n186), .S(n187) );
  FA_X1 U203 ( .A(n198), .B(n195), .CI(n193), .CO(n190), .S(n191) );
  FA_X1 U204 ( .A(n341), .B(n309), .CI(n200), .CO(n192), .S(n193) );
  FA_X1 U205 ( .A(n319), .B(n202), .CI(n330), .CO(n194), .S(n195) );
  FA_X1 U206 ( .A(n206), .B(n201), .CI(n199), .CO(n196), .S(n197) );
  FA_X1 U207 ( .A(n208), .B(n203), .CI(n210), .CO(n198), .S(n199) );
  FA_X1 U208 ( .A(n331), .B(n320), .CI(n342), .CO(n200), .S(n201) );
  FA_X1 U210 ( .A(n214), .B(n209), .CI(n207), .CO(n204), .S(n205) );
  FA_X1 U211 ( .A(n211), .B(n218), .CI(n216), .CO(n206), .S(n207) );
  FA_X1 U212 ( .A(n220), .B(n321), .CI(n354), .CO(n208), .S(n209) );
  FA_X1 U213 ( .A(n332), .B(n310), .CI(n343), .CO(n210), .S(n211) );
  FA_X1 U214 ( .A(n224), .B(n217), .CI(n215), .CO(n212), .S(n213) );
  FA_X1 U215 ( .A(n219), .B(n228), .CI(n226), .CO(n214), .S(n215) );
  FA_X1 U216 ( .A(n221), .B(n311), .CI(n230), .CO(n216), .S(n217) );
  FA_X1 U217 ( .A(n333), .B(n344), .CI(n322), .CO(n218), .S(n219) );
  FA_X1 U220 ( .A(n229), .B(n238), .CI(n236), .CO(n224), .S(n225) );
  FA_X1 U221 ( .A(n240), .B(n366), .CI(n231), .CO(n226), .S(n227) );
  FA_X1 U222 ( .A(n345), .B(n334), .CI(n312), .CO(n228), .S(n229) );
  FA_X1 U225 ( .A(n244), .B(n237), .CI(n235), .CO(n232), .S(n233) );
  FA_X1 U226 ( .A(n246), .B(n248), .CI(n239), .CO(n234), .S(n235) );
  FA_X1 U227 ( .A(n324), .B(n367), .CI(n241), .CO(n236), .S(n237) );
  FA_X1 U228 ( .A(n346), .B(n335), .CI(n313), .CO(n238), .S(n239) );
  HA_X1 U229 ( .A(n300), .B(n356), .CO(n240), .S(n241) );
  FA_X1 U231 ( .A(n254), .B(n256), .CI(n249), .CO(n244), .S(n245) );
  FA_X1 U232 ( .A(n347), .B(n368), .CI(n325), .CO(n246), .S(n247) );
  FA_X1 U233 ( .A(n357), .B(n314), .CI(n336), .CO(n248), .S(n249) );
  FA_X1 U234 ( .A(n255), .B(n260), .CI(n253), .CO(n250), .S(n251) );
  FA_X1 U235 ( .A(n257), .B(n348), .CI(n262), .CO(n252), .S(n253) );
  FA_X1 U236 ( .A(n326), .B(n369), .CI(n337), .CO(n254), .S(n255) );
  HA_X1 U237 ( .A(n301), .B(n358), .CO(n256), .S(n257) );
  FA_X1 U239 ( .A(n338), .B(n349), .CI(n268), .CO(n260), .S(n261) );
  FA_X1 U240 ( .A(n359), .B(n327), .CI(n370), .CO(n262), .S(n263) );
  FA_X1 U241 ( .A(n272), .B(n269), .CI(n267), .CO(n264), .S(n265) );
  FA_X1 U242 ( .A(n339), .B(n371), .CI(n350), .CO(n266), .S(n267) );
  HA_X1 U243 ( .A(n302), .B(n360), .CO(n268), .S(n269) );
  FA_X1 U244 ( .A(n276), .B(n351), .CI(n273), .CO(n270), .S(n271) );
  FA_X1 U245 ( .A(n372), .B(n340), .CI(n361), .CO(n272), .S(n273) );
  FA_X1 U246 ( .A(n352), .B(n303), .CI(n277), .CO(n274), .S(n275) );
  HA_X1 U247 ( .A(n362), .B(n373), .CO(n276), .S(n277) );
  FA_X1 U248 ( .A(n374), .B(n353), .CI(n363), .CO(n278), .S(n279) );
  HA_X1 U249 ( .A(n364), .B(n304), .CO(n280), .S(n281) );
  OR2_X1 U485 ( .A1(n233), .A2(n242), .ZN(n561) );
  INV_X1 U486 ( .A(n488), .ZN(n562) );
  INV_X1 U487 ( .A(n486), .ZN(n563) );
  BUF_X1 U488 ( .A(b[5]), .Z(n462) );
  BUF_X2 U489 ( .A(a[5]), .Z(n495) );
  BUF_X2 U490 ( .A(a[7]), .Z(n494) );
  BUF_X2 U491 ( .A(n505), .Z(n481) );
  NOR2_X1 U492 ( .A1(n233), .A2(n242), .ZN(n109) );
  AND2_X1 U493 ( .A1(n599), .A2(n149), .ZN(product[1]) );
  CLKBUF_X1 U494 ( .A(n583), .Z(n565) );
  CLKBUF_X2 U495 ( .A(b[9]), .Z(n458) );
  XNOR2_X1 U496 ( .A(n71), .B(n566), .ZN(product[17]) );
  AND2_X1 U497 ( .A1(n593), .A2(n70), .ZN(n566) );
  BUF_X1 U498 ( .A(b[7]), .Z(n460) );
  BUF_X1 U499 ( .A(b[3]), .Z(n464) );
  CLKBUF_X1 U500 ( .A(b[0]), .Z(n1) );
  BUF_X1 U501 ( .A(n1), .Z(n567) );
  XNOR2_X1 U502 ( .A(n261), .B(n568), .ZN(n259) );
  XNOR2_X1 U503 ( .A(n263), .B(n266), .ZN(n568) );
  NAND2_X1 U504 ( .A1(n261), .A2(n263), .ZN(n569) );
  NAND2_X1 U505 ( .A1(n261), .A2(n266), .ZN(n570) );
  NAND2_X1 U506 ( .A1(n263), .A2(n266), .ZN(n571) );
  NAND3_X1 U507 ( .A1(n569), .A2(n570), .A3(n571), .ZN(n258) );
  CLKBUF_X1 U508 ( .A(b[0]), .Z(n572) );
  CLKBUF_X1 U509 ( .A(b[2]), .Z(n465) );
  XOR2_X1 U510 ( .A(n252), .B(n247), .Z(n573) );
  XOR2_X1 U511 ( .A(n245), .B(n573), .Z(n243) );
  NAND2_X1 U512 ( .A1(n245), .A2(n252), .ZN(n574) );
  NAND2_X1 U513 ( .A1(n245), .A2(n247), .ZN(n575) );
  NAND2_X1 U514 ( .A1(n252), .A2(n247), .ZN(n576) );
  NAND3_X1 U515 ( .A1(n574), .A2(n575), .A3(n576), .ZN(n242) );
  BUF_X1 U516 ( .A(b[8]), .Z(n459) );
  CLKBUF_X1 U517 ( .A(b[4]), .Z(n577) );
  XOR2_X1 U518 ( .A(n234), .B(n227), .Z(n578) );
  XOR2_X1 U519 ( .A(n225), .B(n578), .Z(n223) );
  NAND2_X1 U520 ( .A1(n225), .A2(n234), .ZN(n579) );
  NAND2_X1 U521 ( .A1(n225), .A2(n227), .ZN(n580) );
  NAND2_X1 U522 ( .A1(n234), .A2(n227), .ZN(n581) );
  NAND3_X1 U523 ( .A1(n579), .A2(n580), .A3(n581), .ZN(n222) );
  CLKBUF_X3 U524 ( .A(a[9]), .Z(n493) );
  OAI21_X1 U525 ( .B1(n118), .B2(n116), .A(n117), .ZN(n582) );
  BUF_X1 U526 ( .A(b[6]), .Z(n461) );
  NOR2_X1 U527 ( .A1(n213), .A2(n222), .ZN(n583) );
  CLKBUF_X3 U528 ( .A(n504), .Z(n480) );
  NOR2_X1 U529 ( .A1(n89), .A2(n82), .ZN(n584) );
  NOR2_X2 U530 ( .A1(n197), .A2(n204), .ZN(n82) );
  NOR2_X1 U531 ( .A1(n82), .A2(n89), .ZN(n80) );
  XNOR2_X1 U532 ( .A(n106), .B(n585), .ZN(product[12]) );
  AND2_X1 U533 ( .A1(n160), .A2(n104), .ZN(n585) );
  XNOR2_X1 U534 ( .A(n58), .B(n586), .ZN(product[18]) );
  AND2_X1 U535 ( .A1(n597), .A2(n57), .ZN(n586) );
  CLKBUF_X1 U536 ( .A(n118), .Z(n587) );
  OAI21_X1 U537 ( .B1(n590), .B2(n78), .A(n79), .ZN(n588) );
  INV_X1 U538 ( .A(n94), .ZN(n589) );
  OAI21_X1 U539 ( .B1(n590), .B2(n78), .A(n79), .ZN(n77) );
  AOI21_X1 U540 ( .B1(n107), .B2(n115), .A(n108), .ZN(n590) );
  NOR2_X1 U541 ( .A1(n259), .A2(n264), .ZN(n591) );
  BUF_X2 U542 ( .A(a[1]), .Z(n497) );
  XNOR2_X1 U543 ( .A(n76), .B(n592), .ZN(product[16]) );
  AND2_X1 U544 ( .A1(n594), .A2(n75), .ZN(n592) );
  OR2_X1 U545 ( .A1(n185), .A2(n190), .ZN(n593) );
  OR2_X1 U546 ( .A1(n191), .A2(n196), .ZN(n594) );
  OR2_X1 U547 ( .A1(n176), .A2(n175), .ZN(n595) );
  OR2_X1 U548 ( .A1(n177), .A2(n180), .ZN(n596) );
  OR2_X1 U549 ( .A1(n181), .A2(n184), .ZN(n597) );
  OR2_X1 U550 ( .A1(n376), .A2(n365), .ZN(n598) );
  OR2_X1 U551 ( .A1(n377), .A2(n305), .ZN(n599) );
  OR2_X1 U552 ( .A1(n275), .A2(n278), .ZN(n600) );
  CLKBUF_X3 U553 ( .A(a[11]), .Z(n492) );
  NAND2_X1 U554 ( .A1(n151), .A2(n30), .ZN(n4) );
  NOR2_X1 U555 ( .A1(n174), .A2(n173), .ZN(n29) );
  INV_X1 U556 ( .A(n29), .ZN(n151) );
  NAND2_X1 U557 ( .A1(n174), .A2(n173), .ZN(n30) );
  NAND2_X1 U558 ( .A1(n595), .A2(n37), .ZN(n5) );
  INV_X1 U559 ( .A(n37), .ZN(n35) );
  NAND2_X1 U560 ( .A1(n176), .A2(n175), .ZN(n37) );
  BUF_X2 U561 ( .A(n509), .Z(n485) );
  NAND2_X1 U562 ( .A1(n596), .A2(n48), .ZN(n6) );
  INV_X1 U563 ( .A(n48), .ZN(n46) );
  INV_X1 U564 ( .A(n291), .ZN(n341) );
  NAND2_X1 U565 ( .A1(n597), .A2(n596), .ZN(n43) );
  INV_X1 U566 ( .A(n597), .ZN(n52) );
  NOR2_X1 U567 ( .A1(n65), .A2(n52), .ZN(n50) );
  OAI21_X1 U568 ( .B1(n62), .B2(n52), .A(n57), .ZN(n51) );
  CLKBUF_X3 U569 ( .A(a[3]), .Z(n496) );
  NAND2_X2 U570 ( .A1(n473), .A2(n509), .ZN(n503) );
  OAI22_X1 U571 ( .A1(n503), .A2(n451), .B1(n450), .B2(n485), .ZN(n374) );
  OAI22_X1 U572 ( .A1(n503), .A2(n448), .B1(n447), .B2(n485), .ZN(n371) );
  OAI22_X1 U573 ( .A1(n503), .A2(n447), .B1(n446), .B2(n485), .ZN(n370) );
  OAI22_X1 U574 ( .A1(n503), .A2(n444), .B1(n443), .B2(n485), .ZN(n367) );
  OAI22_X1 U575 ( .A1(n503), .A2(n446), .B1(n445), .B2(n485), .ZN(n369) );
  INV_X1 U576 ( .A(n41), .ZN(n39) );
  NOR2_X1 U577 ( .A1(n65), .A2(n43), .ZN(n41) );
  OAI22_X1 U578 ( .A1(n503), .A2(n445), .B1(n444), .B2(n485), .ZN(n368) );
  INV_X1 U579 ( .A(n64), .ZN(n62) );
  NAND2_X1 U580 ( .A1(n251), .A2(n258), .ZN(n117) );
  OAI22_X1 U581 ( .A1(n503), .A2(n449), .B1(n448), .B2(n485), .ZN(n372) );
  NOR2_X1 U582 ( .A1(n265), .A2(n270), .ZN(n124) );
  NOR2_X1 U583 ( .A1(n94), .A2(n87), .ZN(n85) );
  NAND2_X1 U584 ( .A1(n279), .A2(n280), .ZN(n137) );
  NAND2_X1 U585 ( .A1(n271), .A2(n274), .ZN(n129) );
  NAND2_X1 U586 ( .A1(n177), .A2(n180), .ZN(n48) );
  INV_X1 U587 ( .A(n158), .ZN(n87) );
  INV_X1 U588 ( .A(n65), .ZN(n63) );
  NAND2_X2 U589 ( .A1(n469), .A2(n505), .ZN(n499) );
  NAND2_X2 U590 ( .A1(n470), .A2(n506), .ZN(n500) );
  INV_X1 U591 ( .A(n66), .ZN(n64) );
  AOI21_X1 U592 ( .B1(n73), .B2(n593), .A(n68), .ZN(n66) );
  NAND2_X1 U593 ( .A1(n162), .A2(n113), .ZN(n15) );
  BUF_X2 U594 ( .A(n507), .Z(n483) );
  NAND2_X1 U595 ( .A1(n594), .A2(n593), .ZN(n65) );
  XNOR2_X1 U596 ( .A(a[3]), .B(a[4]), .ZN(n507) );
  INV_X1 U597 ( .A(n89), .ZN(n158) );
  NAND2_X1 U598 ( .A1(n164), .A2(n122), .ZN(n17) );
  INV_X1 U599 ( .A(n136), .ZN(n168) );
  OAI21_X1 U600 ( .B1(n136), .B2(n138), .A(n137), .ZN(n135) );
  NOR2_X1 U601 ( .A1(n279), .A2(n280), .ZN(n136) );
  INV_X1 U602 ( .A(n128), .ZN(n166) );
  NOR2_X1 U603 ( .A1(n271), .A2(n274), .ZN(n128) );
  NAND2_X2 U604 ( .A1(n471), .A2(n507), .ZN(n501) );
  OAI22_X1 U605 ( .A1(n498), .A2(n379), .B1(n480), .B2(n378), .ZN(n172) );
  INV_X1 U606 ( .A(n97), .ZN(n95) );
  XNOR2_X1 U607 ( .A(n497), .B(n457), .ZN(n444) );
  XNOR2_X1 U608 ( .A(b[4]), .B(n497), .ZN(n450) );
  XNOR2_X1 U609 ( .A(n497), .B(n461), .ZN(n448) );
  OAI22_X1 U610 ( .A1(n503), .A2(n491), .B1(n455), .B2(n485), .ZN(n305) );
  INV_X1 U611 ( .A(n146), .ZN(n144) );
  INV_X1 U612 ( .A(n42), .ZN(n40) );
  INV_X1 U613 ( .A(n95), .ZN(n93) );
  INV_X1 U614 ( .A(n124), .ZN(n165) );
  INV_X1 U615 ( .A(n134), .ZN(n132) );
  AOI21_X1 U616 ( .B1(n55), .B2(n596), .A(n46), .ZN(n44) );
  OAI21_X1 U617 ( .B1(n66), .B2(n43), .A(n44), .ZN(n42) );
  INV_X1 U618 ( .A(n140), .ZN(n169) );
  NOR2_X1 U619 ( .A1(n281), .A2(n375), .ZN(n140) );
  NAND2_X1 U620 ( .A1(n265), .A2(n270), .ZN(n125) );
  NAND2_X2 U621 ( .A1(n468), .A2(n504), .ZN(n498) );
  NOR2_X1 U622 ( .A1(n98), .A2(n103), .ZN(n96) );
  NOR2_X1 U623 ( .A1(n213), .A2(n222), .ZN(n98) );
  NOR2_X1 U624 ( .A1(n223), .A2(n232), .ZN(n103) );
  NAND2_X1 U625 ( .A1(n259), .A2(n264), .ZN(n122) );
  NOR2_X1 U626 ( .A1(n259), .A2(n264), .ZN(n121) );
  OAI22_X1 U627 ( .A1(n503), .A2(n454), .B1(n453), .B2(n485), .ZN(n377) );
  OAI22_X1 U628 ( .A1(n452), .A2(n503), .B1(n451), .B2(n485), .ZN(n375) );
  AOI21_X1 U629 ( .B1(n598), .B2(n147), .A(n144), .ZN(n142) );
  NAND2_X1 U630 ( .A1(n376), .A2(n365), .ZN(n146) );
  OAI22_X1 U631 ( .A1(n503), .A2(n453), .B1(n452), .B2(n485), .ZN(n376) );
  NAND2_X1 U632 ( .A1(n157), .A2(n83), .ZN(n10) );
  INV_X1 U633 ( .A(n82), .ZN(n157) );
  INV_X1 U634 ( .A(n482), .ZN(n289) );
  OAI22_X1 U635 ( .A1(n500), .A2(n415), .B1(n414), .B2(n482), .ZN(n339) );
  OAI22_X1 U636 ( .A1(n500), .A2(n410), .B1(n482), .B2(n409), .ZN(n334) );
  OAI22_X1 U637 ( .A1(n500), .A2(n405), .B1(n482), .B2(n404), .ZN(n329) );
  AOI21_X1 U638 ( .B1(n500), .B2(n482), .A(n404), .ZN(n288) );
  OAI22_X1 U639 ( .A1(n500), .A2(n409), .B1(n482), .B2(n408), .ZN(n333) );
  CLKBUF_X3 U640 ( .A(n506), .Z(n482) );
  INV_X1 U641 ( .A(n288), .ZN(n328) );
  OAI21_X1 U642 ( .B1(n583), .B2(n104), .A(n99), .ZN(n97) );
  INV_X1 U643 ( .A(n104), .ZN(n102) );
  NAND2_X1 U644 ( .A1(n275), .A2(n278), .ZN(n134) );
  OAI22_X1 U645 ( .A1(n503), .A2(n450), .B1(n449), .B2(n485), .ZN(n373) );
  XNOR2_X1 U646 ( .A(n497), .B(n462), .ZN(n449) );
  NOR2_X1 U647 ( .A1(n32), .A2(n29), .ZN(n27) );
  NAND2_X1 U648 ( .A1(n41), .A2(n595), .ZN(n32) );
  NAND2_X1 U649 ( .A1(n281), .A2(n375), .ZN(n141) );
  INV_X1 U650 ( .A(n57), .ZN(n55) );
  NAND2_X1 U651 ( .A1(n197), .A2(n204), .ZN(n83) );
  INV_X1 U652 ( .A(n591), .ZN(n164) );
  XNOR2_X1 U653 ( .A(n497), .B(n464), .ZN(n451) );
  NAND2_X1 U654 ( .A1(n181), .A2(n184), .ZN(n57) );
  OAI22_X1 U655 ( .A1(n500), .A2(n406), .B1(n482), .B2(n405), .ZN(n330) );
  INV_X1 U656 ( .A(n103), .ZN(n160) );
  OAI22_X1 U657 ( .A1(n500), .A2(n408), .B1(n482), .B2(n407), .ZN(n332) );
  INV_X1 U658 ( .A(n112), .ZN(n162) );
  NOR2_X1 U659 ( .A1(n243), .A2(n250), .ZN(n112) );
  OAI22_X1 U660 ( .A1(n500), .A2(n488), .B1(n416), .B2(n482), .ZN(n302) );
  NAND2_X1 U661 ( .A1(n159), .A2(n99), .ZN(n12) );
  INV_X1 U662 ( .A(n565), .ZN(n159) );
  BUF_X2 U663 ( .A(b[10]), .Z(n457) );
  NAND2_X1 U664 ( .A1(n223), .A2(n232), .ZN(n104) );
  XNOR2_X1 U665 ( .A(n497), .B(n458), .ZN(n445) );
  OAI22_X1 U666 ( .A1(n387), .A2(n480), .B1(n388), .B2(n498), .ZN(n312) );
  OAI22_X1 U667 ( .A1(n387), .A2(n498), .B1(n386), .B2(n480), .ZN(n311) );
  OAI22_X1 U668 ( .A1(n498), .A2(n386), .B1(n385), .B2(n480), .ZN(n310) );
  OAI22_X1 U669 ( .A1(n498), .A2(n384), .B1(n480), .B2(n383), .ZN(n309) );
  OAI22_X1 U670 ( .A1(n498), .A2(n382), .B1(n480), .B2(n381), .ZN(n308) );
  OAI22_X1 U671 ( .A1(n498), .A2(n380), .B1(n480), .B2(n379), .ZN(n307) );
  AOI21_X1 U672 ( .B1(n498), .B2(n480), .A(n378), .ZN(n282) );
  INV_X1 U673 ( .A(n172), .ZN(n173) );
  INV_X1 U674 ( .A(n282), .ZN(n306) );
  BUF_X1 U675 ( .A(n1), .Z(n601) );
  NAND2_X1 U676 ( .A1(n243), .A2(n250), .ZN(n113) );
  OAI22_X1 U677 ( .A1(n501), .A2(n427), .B1(n426), .B2(n483), .ZN(n351) );
  OAI22_X1 U678 ( .A1(n501), .A2(n424), .B1(n423), .B2(n483), .ZN(n348) );
  OAI22_X1 U679 ( .A1(n501), .A2(n426), .B1(n425), .B2(n483), .ZN(n350) );
  OAI22_X1 U680 ( .A1(n501), .A2(n428), .B1(n427), .B2(n483), .ZN(n352) );
  OAI22_X1 U681 ( .A1(n501), .A2(n489), .B1(n429), .B2(n483), .ZN(n303) );
  INV_X1 U682 ( .A(n483), .ZN(n292) );
  OAI22_X1 U683 ( .A1(n501), .A2(n425), .B1(n424), .B2(n483), .ZN(n349) );
  OAI22_X1 U684 ( .A1(n501), .A2(n423), .B1(n422), .B2(n483), .ZN(n347) );
  OAI22_X1 U685 ( .A1(n501), .A2(n422), .B1(n421), .B2(n483), .ZN(n346) );
  AOI21_X1 U686 ( .B1(n501), .B2(n483), .A(n417), .ZN(n291) );
  OAI22_X1 U687 ( .A1(n501), .A2(n419), .B1(n418), .B2(n483), .ZN(n343) );
  OAI22_X1 U688 ( .A1(n501), .A2(n418), .B1(n417), .B2(n483), .ZN(n342) );
  OAI22_X1 U689 ( .A1(n501), .A2(n421), .B1(n420), .B2(n483), .ZN(n345) );
  OAI22_X1 U690 ( .A1(n501), .A2(n420), .B1(n419), .B2(n483), .ZN(n344) );
  INV_X1 U691 ( .A(n96), .ZN(n94) );
  XNOR2_X1 U692 ( .A(a[5]), .B(a[6]), .ZN(n506) );
  XNOR2_X1 U693 ( .A(n497), .B(n459), .ZN(n446) );
  NAND2_X2 U694 ( .A1(n508), .A2(n472), .ZN(n502) );
  XNOR2_X1 U695 ( .A(n497), .B(n460), .ZN(n447) );
  OAI22_X1 U696 ( .A1(n500), .A2(n414), .B1(n413), .B2(n482), .ZN(n338) );
  OAI22_X1 U697 ( .A1(n413), .A2(n500), .B1(n482), .B2(n412), .ZN(n337) );
  OAI22_X1 U698 ( .A1(n500), .A2(n412), .B1(n482), .B2(n411), .ZN(n336) );
  OAI22_X1 U699 ( .A1(n498), .A2(n486), .B1(n390), .B2(n480), .ZN(n300) );
  AND2_X1 U700 ( .A1(n601), .A2(n295), .ZN(n365) );
  NAND2_X1 U701 ( .A1(n158), .A2(n90), .ZN(n11) );
  OAI21_X1 U702 ( .B1(n90), .B2(n82), .A(n83), .ZN(n81) );
  OAI21_X1 U703 ( .B1(n95), .B2(n87), .A(n90), .ZN(n86) );
  NOR2_X1 U704 ( .A1(n205), .A2(n212), .ZN(n89) );
  OAI22_X1 U705 ( .A1(n500), .A2(n407), .B1(n482), .B2(n406), .ZN(n331) );
  INV_X1 U706 ( .A(n297), .ZN(n366) );
  AOI21_X1 U707 ( .B1(n503), .B2(n485), .A(n443), .ZN(n297) );
  AOI21_X1 U708 ( .B1(n97), .B2(n584), .A(n81), .ZN(n79) );
  NAND2_X1 U709 ( .A1(n205), .A2(n212), .ZN(n90) );
  INV_X1 U710 ( .A(n481), .ZN(n286) );
  OAI22_X1 U711 ( .A1(n401), .A2(n481), .B1(n499), .B2(n402), .ZN(n326) );
  OAI22_X1 U712 ( .A1(n400), .A2(n481), .B1(n401), .B2(n499), .ZN(n325) );
  OAI22_X1 U713 ( .A1(n499), .A2(n398), .B1(n481), .B2(n397), .ZN(n322) );
  OAI22_X1 U714 ( .A1(n499), .A2(n397), .B1(n481), .B2(n396), .ZN(n321) );
  OAI22_X1 U715 ( .A1(n499), .A2(n396), .B1(n481), .B2(n395), .ZN(n320) );
  OAI22_X1 U716 ( .A1(n499), .A2(n395), .B1(n481), .B2(n394), .ZN(n319) );
  OAI22_X1 U717 ( .A1(n499), .A2(n394), .B1(n481), .B2(n393), .ZN(n318) );
  OAI22_X1 U718 ( .A1(n499), .A2(n393), .B1(n481), .B2(n392), .ZN(n317) );
  OAI22_X1 U719 ( .A1(n499), .A2(n392), .B1(n481), .B2(n391), .ZN(n316) );
  AOI21_X1 U720 ( .B1(n499), .B2(n481), .A(n391), .ZN(n285) );
  OAI22_X1 U721 ( .A1(n499), .A2(n287), .B1(n403), .B2(n481), .ZN(n301) );
  INV_X1 U722 ( .A(n285), .ZN(n315) );
  XNOR2_X1 U723 ( .A(n497), .B(n456), .ZN(n443) );
  BUF_X2 U724 ( .A(b[11]), .Z(n456) );
  OAI22_X1 U725 ( .A1(n400), .A2(n499), .B1(n481), .B2(n399), .ZN(n324) );
  XOR2_X1 U726 ( .A(a[11]), .B(a[10]), .Z(n468) );
  OAI21_X1 U727 ( .B1(n33), .B2(n29), .A(n30), .ZN(n28) );
  AOI21_X1 U728 ( .B1(n42), .B2(n595), .A(n35), .ZN(n33) );
  NAND2_X1 U729 ( .A1(n213), .A2(n222), .ZN(n99) );
  OR2_X1 U730 ( .A1(n323), .A2(n355), .ZN(n230) );
  OAI22_X1 U731 ( .A1(n499), .A2(n399), .B1(n398), .B2(n481), .ZN(n323) );
  XOR2_X1 U732 ( .A(a[1]), .B(a[0]), .Z(n473) );
  OAI21_X1 U733 ( .B1(n109), .B2(n113), .A(n110), .ZN(n108) );
  NOR2_X1 U734 ( .A1(n109), .A2(n112), .ZN(n107) );
  NAND2_X1 U735 ( .A1(n561), .A2(n110), .ZN(n14) );
  NAND2_X1 U736 ( .A1(n233), .A2(n242), .ZN(n110) );
  OAI22_X1 U737 ( .A1(n500), .A2(n411), .B1(n482), .B2(n410), .ZN(n335) );
  INV_X1 U738 ( .A(n70), .ZN(n68) );
  OAI22_X1 U739 ( .A1(n388), .A2(n480), .B1(n498), .B2(n389), .ZN(n313) );
  XNOR2_X1 U740 ( .A(a[7]), .B(a[8]), .ZN(n505) );
  XNOR2_X1 U741 ( .A(n493), .B(n456), .ZN(n391) );
  XNOR2_X1 U742 ( .A(n493), .B(n457), .ZN(n392) );
  XNOR2_X1 U743 ( .A(n493), .B(n459), .ZN(n394) );
  XNOR2_X1 U744 ( .A(n493), .B(n458), .ZN(n393) );
  XNOR2_X1 U745 ( .A(n466), .B(n493), .ZN(n401) );
  XNOR2_X1 U746 ( .A(n493), .B(n460), .ZN(n395) );
  XNOR2_X1 U747 ( .A(n493), .B(n462), .ZN(n397) );
  XNOR2_X1 U748 ( .A(n493), .B(n461), .ZN(n396) );
  XNOR2_X1 U749 ( .A(n464), .B(n493), .ZN(n399) );
  XNOR2_X1 U750 ( .A(b[4]), .B(n493), .ZN(n398) );
  NAND2_X1 U751 ( .A1(n191), .A2(n196), .ZN(n75) );
  INV_X1 U752 ( .A(n75), .ZN(n73) );
  NAND2_X1 U753 ( .A1(n185), .A2(n190), .ZN(n70) );
  OAI22_X1 U754 ( .A1(n498), .A2(n381), .B1(n480), .B2(n380), .ZN(n178) );
  INV_X1 U755 ( .A(n178), .ZN(n179) );
  INV_X1 U756 ( .A(n480), .ZN(n283) );
  NAND2_X1 U757 ( .A1(n96), .A2(n80), .ZN(n78) );
  OAI21_X1 U758 ( .B1(n121), .B2(n125), .A(n122), .ZN(n120) );
  NOR2_X1 U759 ( .A1(n591), .A2(n124), .ZN(n119) );
  AOI21_X1 U760 ( .B1(n582), .B2(n107), .A(n108), .ZN(n106) );
  CLKBUF_X3 U761 ( .A(n508), .Z(n484) );
  INV_X1 U762 ( .A(n139), .ZN(n138) );
  OAI21_X1 U763 ( .B1(n140), .B2(n142), .A(n141), .ZN(n139) );
  XNOR2_X1 U764 ( .A(n466), .B(n497), .ZN(n453) );
  BUF_X2 U765 ( .A(b[1]), .Z(n466) );
  XOR2_X1 U766 ( .A(a[5]), .B(a[4]), .Z(n471) );
  XNOR2_X1 U767 ( .A(n465), .B(n497), .ZN(n452) );
  XNOR2_X1 U768 ( .A(n465), .B(n493), .ZN(n400) );
  INV_X1 U769 ( .A(n484), .ZN(n295) );
  OAI22_X1 U770 ( .A1(n439), .A2(n484), .B1(n440), .B2(n502), .ZN(n363) );
  OAI22_X1 U771 ( .A1(n439), .A2(n502), .B1(n484), .B2(n438), .ZN(n362) );
  OAI22_X1 U772 ( .A1(n502), .A2(n438), .B1(n484), .B2(n437), .ZN(n361) );
  OAI22_X1 U773 ( .A1(n502), .A2(n437), .B1(n484), .B2(n436), .ZN(n360) );
  OAI22_X1 U774 ( .A1(n502), .A2(n436), .B1(n484), .B2(n435), .ZN(n359) );
  OAI22_X1 U775 ( .A1(n502), .A2(n435), .B1(n484), .B2(n434), .ZN(n358) );
  OAI22_X1 U776 ( .A1(n502), .A2(n434), .B1(n484), .B2(n433), .ZN(n357) );
  OAI22_X1 U777 ( .A1(n433), .A2(n502), .B1(n484), .B2(n432), .ZN(n356) );
  OAI22_X1 U778 ( .A1(n502), .A2(n432), .B1(n484), .B2(n431), .ZN(n355) );
  OAI22_X1 U779 ( .A1(n502), .A2(n431), .B1(n484), .B2(n430), .ZN(n220) );
  AOI21_X1 U780 ( .B1(n502), .B2(n484), .A(n430), .ZN(n294) );
  XNOR2_X1 U781 ( .A(n323), .B(n355), .ZN(n231) );
  INV_X1 U782 ( .A(n294), .ZN(n354) );
  OAI22_X1 U783 ( .A1(n498), .A2(n383), .B1(n480), .B2(n382), .ZN(n188) );
  INV_X1 U784 ( .A(n188), .ZN(n189) );
  OR2_X1 U785 ( .A1(n567), .A2(n491), .ZN(n455) );
  OR2_X1 U786 ( .A1(n567), .A2(n287), .ZN(n403) );
  AND2_X1 U787 ( .A1(n567), .A2(n286), .ZN(n327) );
  AND2_X1 U788 ( .A1(n572), .A2(n289), .ZN(n340) );
  OR2_X1 U789 ( .A1(n572), .A2(n490), .ZN(n442) );
  OR2_X1 U790 ( .A1(n567), .A2(n488), .ZN(n416) );
  OR2_X1 U791 ( .A1(n1), .A2(n486), .ZN(n390) );
  AND2_X1 U792 ( .A1(n572), .A2(n292), .ZN(n353) );
  OR2_X1 U793 ( .A1(n567), .A2(n489), .ZN(n429) );
  AND2_X1 U794 ( .A1(n567), .A2(n283), .ZN(n314) );
  XNOR2_X1 U795 ( .A(n601), .B(n493), .ZN(n402) );
  XNOR2_X1 U796 ( .A(n601), .B(n497), .ZN(n454) );
  OAI22_X1 U797 ( .A1(n440), .A2(n484), .B1(n502), .B2(n441), .ZN(n364) );
  XOR2_X1 U798 ( .A(a[7]), .B(a[6]), .Z(n470) );
  XNOR2_X1 U799 ( .A(a[1]), .B(a[2]), .ZN(n508) );
  XOR2_X1 U800 ( .A(a[9]), .B(a[8]), .Z(n469) );
  XNOR2_X1 U801 ( .A(n496), .B(n460), .ZN(n434) );
  XNOR2_X1 U802 ( .A(n496), .B(n461), .ZN(n435) );
  XNOR2_X1 U803 ( .A(n465), .B(n496), .ZN(n439) );
  XNOR2_X1 U804 ( .A(n464), .B(n496), .ZN(n438) );
  XNOR2_X1 U805 ( .A(b[4]), .B(n496), .ZN(n437) );
  XNOR2_X1 U806 ( .A(n496), .B(n457), .ZN(n431) );
  XNOR2_X1 U807 ( .A(n496), .B(n459), .ZN(n433) );
  XNOR2_X1 U808 ( .A(n496), .B(n458), .ZN(n432) );
  XNOR2_X1 U809 ( .A(n496), .B(n462), .ZN(n436) );
  XNOR2_X1 U810 ( .A(n496), .B(n456), .ZN(n430) );
  XNOR2_X1 U811 ( .A(n466), .B(n496), .ZN(n440) );
  XNOR2_X1 U812 ( .A(n1), .B(n496), .ZN(n441) );
  INV_X1 U813 ( .A(n495), .ZN(n489) );
  XNOR2_X1 U814 ( .A(n495), .B(n456), .ZN(n417) );
  XNOR2_X1 U815 ( .A(n601), .B(n495), .ZN(n428) );
  XNOR2_X1 U816 ( .A(n466), .B(n495), .ZN(n427) );
  XNOR2_X1 U817 ( .A(n495), .B(n462), .ZN(n423) );
  XNOR2_X1 U818 ( .A(n465), .B(n495), .ZN(n426) );
  XNOR2_X1 U819 ( .A(n495), .B(n461), .ZN(n422) );
  XNOR2_X1 U820 ( .A(n495), .B(n577), .ZN(n424) );
  XNOR2_X1 U821 ( .A(n495), .B(n464), .ZN(n425) );
  XNOR2_X1 U822 ( .A(n495), .B(n457), .ZN(n418) );
  XNOR2_X1 U823 ( .A(n495), .B(n458), .ZN(n419) );
  XNOR2_X1 U824 ( .A(n495), .B(n460), .ZN(n421) );
  XNOR2_X1 U825 ( .A(n495), .B(n459), .ZN(n420) );
  OAI22_X1 U826 ( .A1(n498), .A2(n385), .B1(n480), .B2(n384), .ZN(n202) );
  INV_X1 U827 ( .A(n202), .ZN(n203) );
  INV_X1 U828 ( .A(n493), .ZN(n287) );
  XNOR2_X1 U829 ( .A(a[9]), .B(a[10]), .ZN(n504) );
  INV_X1 U830 ( .A(n116), .ZN(n163) );
  OAI21_X1 U831 ( .B1(n116), .B2(n118), .A(n117), .ZN(n115) );
  NOR2_X1 U832 ( .A1(n251), .A2(n258), .ZN(n116) );
  XNOR2_X1 U833 ( .A(n563), .B(n457), .ZN(n379) );
  XNOR2_X1 U834 ( .A(n456), .B(n563), .ZN(n378) );
  XNOR2_X1 U835 ( .A(n563), .B(n459), .ZN(n381) );
  XNOR2_X1 U836 ( .A(n563), .B(n458), .ZN(n380) );
  INV_X1 U837 ( .A(n492), .ZN(n486) );
  XNOR2_X1 U838 ( .A(n572), .B(n492), .ZN(n389) );
  XNOR2_X1 U839 ( .A(n465), .B(n492), .ZN(n387) );
  XNOR2_X1 U840 ( .A(n464), .B(n492), .ZN(n386) );
  XNOR2_X1 U841 ( .A(n466), .B(n492), .ZN(n388) );
  XNOR2_X1 U842 ( .A(n492), .B(n461), .ZN(n383) );
  XNOR2_X1 U843 ( .A(n492), .B(n460), .ZN(n382) );
  XNOR2_X1 U844 ( .A(b[4]), .B(n492), .ZN(n385) );
  XNOR2_X1 U845 ( .A(n563), .B(n462), .ZN(n384) );
  INV_X1 U846 ( .A(n497), .ZN(n491) );
  INV_X1 U847 ( .A(n220), .ZN(n221) );
  OAI22_X1 U848 ( .A1(n502), .A2(n490), .B1(n442), .B2(n484), .ZN(n304) );
  INV_X1 U849 ( .A(n496), .ZN(n490) );
  XNOR2_X1 U850 ( .A(n562), .B(n457), .ZN(n405) );
  XNOR2_X1 U851 ( .A(n562), .B(n456), .ZN(n404) );
  XNOR2_X1 U852 ( .A(n494), .B(n458), .ZN(n406) );
  XNOR2_X1 U853 ( .A(n494), .B(n464), .ZN(n412) );
  XNOR2_X1 U854 ( .A(b[4]), .B(n494), .ZN(n411) );
  XNOR2_X1 U855 ( .A(n572), .B(n494), .ZN(n415) );
  XNOR2_X1 U856 ( .A(n494), .B(n459), .ZN(n407) );
  INV_X1 U857 ( .A(n494), .ZN(n488) );
  XNOR2_X1 U858 ( .A(n494), .B(n460), .ZN(n408) );
  XNOR2_X1 U859 ( .A(n465), .B(n494), .ZN(n413) );
  XNOR2_X1 U860 ( .A(n466), .B(n494), .ZN(n414) );
  XNOR2_X1 U861 ( .A(n494), .B(n462), .ZN(n410) );
  XNOR2_X1 U862 ( .A(n494), .B(n461), .ZN(n409) );
  XOR2_X1 U863 ( .A(a[3]), .B(a[2]), .Z(n472) );
  INV_X1 U864 ( .A(n149), .ZN(n147) );
  NAND2_X1 U865 ( .A1(n377), .A2(n305), .ZN(n149) );
  OAI21_X1 U866 ( .B1(n130), .B2(n128), .A(n129), .ZN(n127) );
  INV_X1 U867 ( .A(a[0]), .ZN(n509) );
  AOI21_X1 U868 ( .B1(n588), .B2(n27), .A(n28), .ZN(n26) );
  AND2_X1 U869 ( .A1(n567), .A2(a[0]), .ZN(product[0]) );
  XNOR2_X1 U870 ( .A(n23), .B(n147), .ZN(product[2]) );
  NAND2_X1 U871 ( .A1(n598), .A2(n146), .ZN(n23) );
  XOR2_X1 U872 ( .A(n21), .B(n138), .Z(product[4]) );
  NAND2_X1 U873 ( .A1(n168), .A2(n137), .ZN(n21) );
  AOI21_X1 U874 ( .B1(n600), .B2(n135), .A(n132), .ZN(n130) );
  XOR2_X1 U875 ( .A(n22), .B(n142), .Z(product[3]) );
  NAND2_X1 U876 ( .A1(n169), .A2(n141), .ZN(n22) );
  XOR2_X1 U877 ( .A(n19), .B(n130), .Z(product[6]) );
  NAND2_X1 U878 ( .A1(n166), .A2(n129), .ZN(n19) );
  XNOR2_X1 U879 ( .A(n20), .B(n135), .ZN(product[5]) );
  NAND2_X1 U880 ( .A1(n600), .A2(n134), .ZN(n20) );
  NAND2_X1 U881 ( .A1(n165), .A2(n125), .ZN(n18) );
  XOR2_X1 U882 ( .A(n587), .B(n16), .Z(product[9]) );
  NAND2_X1 U883 ( .A1(n163), .A2(n117), .ZN(n16) );
  AOI21_X1 U884 ( .B1(n127), .B2(n119), .A(n120), .ZN(n118) );
  XOR2_X1 U885 ( .A(n18), .B(n126), .Z(product[7]) );
  INV_X1 U886 ( .A(n127), .ZN(n126) );
  XNOR2_X1 U887 ( .A(n123), .B(n17), .ZN(product[8]) );
  OAI21_X1 U888 ( .B1(n126), .B2(n124), .A(n125), .ZN(n123) );
  XOR2_X1 U889 ( .A(n114), .B(n15), .Z(product[10]) );
  INV_X1 U890 ( .A(n582), .ZN(n114) );
  INV_X1 U891 ( .A(n106), .ZN(n105) );
  XNOR2_X1 U892 ( .A(n111), .B(n14), .ZN(product[11]) );
  OAI21_X1 U893 ( .B1(n114), .B2(n112), .A(n113), .ZN(n111) );
  XOR2_X1 U894 ( .A(n91), .B(n11), .Z(product[14]) );
  AOI21_X1 U895 ( .B1(n105), .B2(n589), .A(n93), .ZN(n91) );
  XOR2_X1 U896 ( .A(n84), .B(n10), .Z(product[15]) );
  AOI21_X1 U897 ( .B1(n85), .B2(n105), .A(n86), .ZN(n84) );
  XOR2_X1 U898 ( .A(n100), .B(n12), .Z(product[13]) );
  AOI21_X1 U899 ( .B1(n105), .B2(n160), .A(n102), .ZN(n100) );
  AOI21_X1 U900 ( .B1(n588), .B2(n63), .A(n64), .ZN(n58) );
  XNOR2_X1 U901 ( .A(n31), .B(n4), .ZN(product[21]) );
  OAI21_X1 U902 ( .B1(n76), .B2(n32), .A(n33), .ZN(n31) );
  XOR2_X1 U903 ( .A(n49), .B(n6), .Z(product[19]) );
  AOI21_X1 U904 ( .B1(n77), .B2(n50), .A(n51), .ZN(n49) );
  XNOR2_X1 U905 ( .A(n38), .B(n5), .ZN(product[20]) );
  OAI21_X1 U906 ( .B1(n39), .B2(n76), .A(n40), .ZN(n38) );
  AOI21_X1 U907 ( .B1(n77), .B2(n594), .A(n73), .ZN(n71) );
  INV_X1 U908 ( .A(n588), .ZN(n76) );
  INV_X1 U909 ( .A(n26), .ZN(n150) );
  INV_X1 U910 ( .A(n25), .ZN(product[23]) );
endmodule


module datapath_DW_mult_tc_20 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n1, n3, n4, n6, n7, n9, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n25, n26, n27, n28, n30, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n45, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n73, n74, n75, n76, n77, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n103, n105, n106, n108, n110, n111, n112, n114,
         n116, n117, n118, n119, n120, n124, n125, n126, n127, n128, n130,
         n132, n133, n134, n136, n138, n141, n142, n144, n145, n147, n150,
         n153, n154, n158, n160, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n277, n278, n279, n280, n281,
         n283, n284, n285, n286, n287, n289, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n450, n451, n452,
         n453, n456, n457, n458, n460, n461, n462, n463, n464, n465, n472,
         n473, n474, n475, n476, n477, n478, n480, n482, n483, n484, n485,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597;

  FA_X1 U188 ( .A(n299), .B(n170), .CI(n307), .CO(n166), .S(n167) );
  FA_X1 U189 ( .A(n171), .B(n308), .CI(n174), .CO(n168), .S(n169) );
  FA_X1 U191 ( .A(n178), .B(n300), .CI(n175), .CO(n172), .S(n173) );
  FA_X1 U192 ( .A(n309), .B(n180), .CI(n320), .CO(n174), .S(n175) );
  FA_X1 U193 ( .A(n179), .B(n186), .CI(n184), .CO(n176), .S(n177) );
  FA_X1 U194 ( .A(n310), .B(n321), .CI(n181), .CO(n178), .S(n179) );
  FA_X1 U196 ( .A(n190), .B(n187), .CI(n185), .CO(n182), .S(n183) );
  FA_X1 U197 ( .A(n332), .B(n301), .CI(n192), .CO(n184), .S(n185) );
  FA_X1 U198 ( .A(n311), .B(n194), .CI(n322), .CO(n186), .S(n187) );
  FA_X1 U199 ( .A(n191), .B(n193), .CI(n198), .CO(n188), .S(n189) );
  FA_X1 U200 ( .A(n202), .B(n195), .CI(n200), .CO(n190), .S(n191) );
  FA_X1 U201 ( .A(n323), .B(n312), .CI(n333), .CO(n192), .S(n193) );
  FA_X1 U203 ( .A(n206), .B(n201), .CI(n199), .CO(n196), .S(n197) );
  FA_X1 U204 ( .A(n208), .B(n210), .CI(n203), .CO(n198), .S(n199) );
  FA_X1 U205 ( .A(n313), .B(n324), .CI(n345), .CO(n200), .S(n201) );
  FA_X1 U206 ( .A(n302), .B(n334), .CI(n212), .CO(n202), .S(n203) );
  FA_X1 U207 ( .A(n216), .B(n209), .CI(n207), .CO(n204), .S(n205) );
  FA_X1 U208 ( .A(n211), .B(n220), .CI(n218), .CO(n206), .S(n207) );
  FA_X1 U209 ( .A(n213), .B(n303), .CI(n222), .CO(n208), .S(n209) );
  FA_X1 U210 ( .A(n335), .B(n314), .CI(n346), .CO(n210), .S(n211) );
  FA_X1 U213 ( .A(n221), .B(n230), .CI(n228), .CO(n216), .S(n217) );
  FA_X1 U214 ( .A(n232), .B(n358), .CI(n223), .CO(n218), .S(n219) );
  FA_X1 U215 ( .A(n347), .B(n336), .CI(n304), .CO(n220), .S(n221) );
  FA_X1 U218 ( .A(n236), .B(n229), .CI(n227), .CO(n224), .S(n225) );
  FA_X1 U219 ( .A(n238), .B(n240), .CI(n231), .CO(n226), .S(n227) );
  FA_X1 U220 ( .A(n316), .B(n305), .CI(n233), .CO(n228), .S(n229) );
  FA_X1 U221 ( .A(n337), .B(n348), .CI(n292), .CO(n230), .S(n231) );
  HA_X1 U222 ( .A(n359), .B(n326), .CO(n232), .S(n233) );
  FA_X1 U223 ( .A(n244), .B(n239), .CI(n237), .CO(n234), .S(n235) );
  FA_X1 U224 ( .A(n246), .B(n248), .CI(n241), .CO(n236), .S(n237) );
  FA_X1 U225 ( .A(n349), .B(n338), .CI(n317), .CO(n238), .S(n239) );
  FA_X1 U226 ( .A(n327), .B(n306), .CI(n360), .CO(n240), .S(n241) );
  FA_X1 U228 ( .A(n249), .B(n328), .CI(n254), .CO(n244), .S(n245) );
  FA_X1 U229 ( .A(n350), .B(n339), .CI(n318), .CO(n246), .S(n247) );
  HA_X1 U230 ( .A(n293), .B(n361), .CO(n248), .S(n249) );
  FA_X1 U231 ( .A(n255), .B(n258), .CI(n253), .CO(n250), .S(n251) );
  FA_X1 U232 ( .A(n329), .B(n351), .CI(n260), .CO(n252), .S(n253) );
  FA_X1 U233 ( .A(n362), .B(n319), .CI(n340), .CO(n254), .S(n255) );
  FA_X1 U234 ( .A(n264), .B(n261), .CI(n259), .CO(n256), .S(n257) );
  FA_X1 U235 ( .A(n330), .B(n352), .CI(n341), .CO(n258), .S(n259) );
  HA_X1 U236 ( .A(n294), .B(n363), .CO(n260), .S(n261) );
  FA_X1 U237 ( .A(n268), .B(n342), .CI(n265), .CO(n262), .S(n263) );
  FA_X1 U238 ( .A(n364), .B(n331), .CI(n353), .CO(n264), .S(n265) );
  FA_X1 U239 ( .A(n354), .B(n343), .CI(n269), .CO(n266), .S(n267) );
  HA_X1 U240 ( .A(n295), .B(n365), .CO(n268), .S(n269) );
  FA_X1 U241 ( .A(n366), .B(n344), .CI(n355), .CO(n270), .S(n271) );
  HA_X1 U242 ( .A(n367), .B(n296), .CO(n272), .S(n273) );
  CLKBUF_X3 U478 ( .A(a[7]), .Z(n597) );
  CLKBUF_X3 U479 ( .A(a[5]), .Z(n487) );
  AOI21_X1 U480 ( .B1(n591), .B2(n133), .A(n130), .ZN(n128) );
  BUF_X1 U481 ( .A(b[0]), .Z(n1) );
  AND2_X1 U482 ( .A1(n595), .A2(n141), .ZN(product[1]) );
  OR2_X1 U483 ( .A1(n166), .A2(n165), .ZN(n554) );
  CLKBUF_X1 U484 ( .A(n73), .Z(n573) );
  OR2_X1 U485 ( .A1(n576), .A2(n214), .ZN(n555) );
  INV_X1 U486 ( .A(n586), .ZN(n556) );
  NOR2_X1 U487 ( .A1(n225), .A2(n234), .ZN(n557) );
  NOR2_X1 U488 ( .A1(n225), .A2(n234), .ZN(n93) );
  OR2_X1 U489 ( .A1(n189), .A2(n196), .ZN(n558) );
  BUF_X1 U490 ( .A(n36), .Z(n585) );
  BUF_X1 U491 ( .A(b[3]), .Z(n456) );
  CLKBUF_X3 U492 ( .A(a[1]), .Z(n489) );
  BUF_X2 U493 ( .A(n488), .Z(n562) );
  CLKBUF_X1 U494 ( .A(n28), .Z(n559) );
  NAND2_X1 U495 ( .A1(n460), .A2(n496), .ZN(n490) );
  CLKBUF_X3 U496 ( .A(n496), .Z(n472) );
  CLKBUF_X1 U497 ( .A(n492), .Z(n560) );
  NAND2_X1 U498 ( .A1(n498), .A2(n462), .ZN(n492) );
  NAND2_X2 U499 ( .A1(n464), .A2(n500), .ZN(n494) );
  CLKBUF_X1 U500 ( .A(n488), .Z(n561) );
  BUF_X2 U501 ( .A(n488), .Z(n563) );
  BUF_X1 U502 ( .A(a[3]), .Z(n488) );
  CLKBUF_X1 U503 ( .A(n1), .Z(n564) );
  AND2_X1 U504 ( .A1(n369), .A2(n297), .ZN(n565) );
  CLKBUF_X1 U505 ( .A(b[2]), .Z(n457) );
  AND2_X1 U506 ( .A1(n267), .A2(n270), .ZN(n566) );
  CLKBUF_X3 U507 ( .A(a[11]), .Z(n484) );
  CLKBUF_X1 U508 ( .A(n74), .Z(n567) );
  CLKBUF_X1 U509 ( .A(b[8]), .Z(n451) );
  NAND2_X2 U510 ( .A1(n497), .A2(n461), .ZN(n491) );
  XOR2_X1 U511 ( .A(n247), .B(n252), .Z(n568) );
  XOR2_X1 U512 ( .A(n245), .B(n568), .Z(n243) );
  NAND2_X1 U513 ( .A1(n245), .A2(n247), .ZN(n569) );
  NAND2_X1 U514 ( .A1(n245), .A2(n252), .ZN(n570) );
  NAND2_X1 U515 ( .A1(n247), .A2(n252), .ZN(n571) );
  NAND3_X1 U516 ( .A1(n569), .A2(n570), .A3(n571), .ZN(n242) );
  BUF_X1 U517 ( .A(b[6]), .Z(n453) );
  OR2_X1 U518 ( .A1(n82), .A2(n87), .ZN(n572) );
  BUF_X4 U519 ( .A(n498), .Z(n474) );
  NAND2_X2 U520 ( .A1(n463), .A2(n499), .ZN(n493) );
  BUF_X1 U521 ( .A(b[1]), .Z(n458) );
  CLKBUF_X3 U522 ( .A(n497), .Z(n473) );
  BUF_X1 U523 ( .A(b[9]), .Z(n450) );
  CLKBUF_X1 U524 ( .A(n83), .Z(n574) );
  XNOR2_X1 U525 ( .A(n36), .B(n575), .ZN(product[20]) );
  AND2_X1 U526 ( .A1(n144), .A2(n35), .ZN(n575) );
  CLKBUF_X1 U527 ( .A(n205), .Z(n576) );
  XOR2_X1 U528 ( .A(n226), .B(n219), .Z(n577) );
  XOR2_X1 U529 ( .A(n217), .B(n577), .Z(n215) );
  NAND2_X1 U530 ( .A1(n217), .A2(n226), .ZN(n578) );
  NAND2_X1 U531 ( .A1(n217), .A2(n219), .ZN(n579) );
  NAND2_X1 U532 ( .A1(n226), .A2(n219), .ZN(n580) );
  NAND3_X1 U533 ( .A1(n578), .A2(n579), .A3(n580), .ZN(n214) );
  AOI21_X1 U534 ( .B1(n91), .B2(n99), .A(n92), .ZN(n581) );
  AOI21_X1 U535 ( .B1(n99), .B2(n91), .A(n92), .ZN(n90) );
  NOR2_X1 U536 ( .A1(n205), .A2(n214), .ZN(n582) );
  NOR2_X1 U537 ( .A1(n205), .A2(n214), .ZN(n82) );
  XNOR2_X1 U538 ( .A(n55), .B(n583), .ZN(product[17]) );
  AND2_X1 U539 ( .A1(n147), .A2(n54), .ZN(n583) );
  XNOR2_X1 U540 ( .A(n68), .B(n584), .ZN(product[15]) );
  AND2_X1 U541 ( .A1(n558), .A2(n67), .ZN(n584) );
  NAND2_X2 U542 ( .A1(n465), .A2(n501), .ZN(n495) );
  OAI21_X1 U543 ( .B1(n581), .B2(n62), .A(n63), .ZN(n586) );
  CLKBUF_X1 U544 ( .A(n451), .Z(n587) );
  XOR2_X1 U545 ( .A(n98), .B(n15), .Z(product[10]) );
  XNOR2_X1 U546 ( .A(n111), .B(n17), .ZN(product[8]) );
  OR2_X1 U547 ( .A1(n251), .A2(n256), .ZN(n588) );
  OR2_X1 U548 ( .A1(n243), .A2(n250), .ZN(n589) );
  OR2_X1 U549 ( .A1(n173), .A2(n176), .ZN(n590) );
  OR2_X1 U550 ( .A1(n273), .A2(n356), .ZN(n591) );
  OR2_X1 U551 ( .A1(n368), .A2(n357), .ZN(n592) );
  OR2_X1 U552 ( .A1(n257), .A2(n262), .ZN(n593) );
  OR2_X1 U553 ( .A1(n267), .A2(n270), .ZN(n594) );
  OR2_X1 U554 ( .A1(n369), .A2(n297), .ZN(n595) );
  BUF_X1 U555 ( .A(n501), .Z(n477) );
  BUF_X2 U556 ( .A(n499), .Z(n475) );
  BUF_X2 U557 ( .A(a[9]), .Z(n485) );
  BUF_X1 U558 ( .A(b[7]), .Z(n452) );
  NOR2_X1 U559 ( .A1(n298), .A2(n164), .ZN(n26) );
  NOR2_X1 U560 ( .A1(n168), .A2(n167), .ZN(n34) );
  NAND2_X1 U561 ( .A1(n142), .A2(n27), .ZN(n3) );
  INV_X1 U562 ( .A(n26), .ZN(n142) );
  INV_X1 U563 ( .A(n274), .ZN(n298) );
  NAND2_X1 U564 ( .A1(n554), .A2(n32), .ZN(n4) );
  INV_X1 U565 ( .A(n32), .ZN(n30) );
  NAND2_X1 U566 ( .A1(n166), .A2(n165), .ZN(n32) );
  INV_X1 U567 ( .A(n39), .ZN(n145) );
  INV_X1 U568 ( .A(n34), .ZN(n144) );
  NAND2_X1 U569 ( .A1(n168), .A2(n167), .ZN(n35) );
  INV_X1 U570 ( .A(n283), .ZN(n332) );
  NAND2_X1 U571 ( .A1(n298), .A2(n164), .ZN(n27) );
  INV_X1 U572 ( .A(n164), .ZN(n165) );
  OAI22_X1 U573 ( .A1(n490), .A2(n371), .B1(n472), .B2(n370), .ZN(n164) );
  NOR2_X1 U574 ( .A1(n169), .A2(n172), .ZN(n39) );
  NAND2_X1 U575 ( .A1(n145), .A2(n40), .ZN(n6) );
  NAND2_X1 U576 ( .A1(n169), .A2(n172), .ZN(n40) );
  NAND2_X1 U577 ( .A1(n590), .A2(n47), .ZN(n7) );
  INV_X1 U578 ( .A(n47), .ZN(n45) );
  NAND2_X1 U579 ( .A1(n173), .A2(n176), .ZN(n47) );
  NOR2_X1 U580 ( .A1(n177), .A2(n182), .ZN(n53) );
  AND2_X1 U581 ( .A1(n1), .A2(n284), .ZN(n344) );
  AOI21_X1 U582 ( .B1(n52), .B2(n590), .A(n45), .ZN(n43) );
  OR2_X1 U583 ( .A1(n1), .A2(n483), .ZN(n447) );
  NOR2_X1 U584 ( .A1(n42), .A2(n39), .ZN(n37) );
  OR2_X1 U585 ( .A1(n1), .A2(n482), .ZN(n434) );
  OR2_X1 U586 ( .A1(n1), .A2(n480), .ZN(n408) );
  INV_X1 U587 ( .A(n280), .ZN(n320) );
  BUF_X2 U588 ( .A(n500), .Z(n476) );
  AND2_X1 U589 ( .A1(n1), .A2(n275), .ZN(n306) );
  INV_X1 U590 ( .A(n476), .ZN(n287) );
  AND2_X1 U591 ( .A1(n564), .A2(n287), .ZN(n357) );
  INV_X1 U592 ( .A(n286), .ZN(n345) );
  AOI21_X1 U593 ( .B1(n494), .B2(n476), .A(n422), .ZN(n286) );
  OR2_X1 U594 ( .A1(n1), .A2(n279), .ZN(n395) );
  INV_X1 U595 ( .A(n96), .ZN(n154) );
  INV_X1 U596 ( .A(n79), .ZN(n77) );
  NAND2_X1 U597 ( .A1(n263), .A2(n266), .ZN(n119) );
  NOR2_X1 U598 ( .A1(n263), .A2(n266), .ZN(n118) );
  NAND2_X1 U599 ( .A1(n51), .A2(n590), .ZN(n42) );
  INV_X1 U600 ( .A(n51), .ZN(n49) );
  NOR2_X1 U601 ( .A1(n58), .A2(n53), .ZN(n51) );
  INV_X1 U602 ( .A(n572), .ZN(n76) );
  NOR2_X1 U603 ( .A1(n572), .A2(n573), .ZN(n69) );
  NAND2_X1 U604 ( .A1(n189), .A2(n196), .ZN(n67) );
  NAND2_X1 U605 ( .A1(n589), .A2(n105), .ZN(n16) );
  INV_X1 U606 ( .A(n118), .ZN(n158) );
  AND2_X1 U607 ( .A1(n1), .A2(n281), .ZN(n331) );
  OAI21_X1 U608 ( .B1(n43), .B2(n39), .A(n40), .ZN(n38) );
  INV_X1 U609 ( .A(n573), .ZN(n150) );
  INV_X1 U610 ( .A(n52), .ZN(n50) );
  OAI21_X1 U611 ( .B1(n59), .B2(n53), .A(n54), .ZN(n52) );
  INV_X1 U612 ( .A(n81), .ZN(n79) );
  NAND2_X1 U613 ( .A1(n368), .A2(n357), .ZN(n138) );
  INV_X1 U614 ( .A(n126), .ZN(n160) );
  NOR2_X1 U615 ( .A1(n271), .A2(n272), .ZN(n126) );
  INV_X1 U616 ( .A(n116), .ZN(n114) );
  NAND2_X1 U617 ( .A1(n257), .A2(n262), .ZN(n116) );
  NAND2_X1 U618 ( .A1(n243), .A2(n250), .ZN(n105) );
  NOR2_X1 U619 ( .A1(n215), .A2(n224), .ZN(n87) );
  NAND2_X1 U620 ( .A1(n267), .A2(n270), .ZN(n124) );
  OR2_X1 U621 ( .A1(n1), .A2(n285), .ZN(n421) );
  NAND2_X1 U622 ( .A1(n271), .A2(n272), .ZN(n127) );
  NAND2_X1 U623 ( .A1(n588), .A2(n110), .ZN(n17) );
  INV_X1 U624 ( .A(n110), .ZN(n108) );
  NAND2_X1 U625 ( .A1(n251), .A2(n256), .ZN(n110) );
  INV_X1 U626 ( .A(n138), .ZN(n136) );
  NAND2_X1 U627 ( .A1(n273), .A2(n356), .ZN(n132) );
  NAND2_X1 U628 ( .A1(n153), .A2(n94), .ZN(n14) );
  INV_X1 U629 ( .A(n557), .ZN(n153) );
  OR2_X1 U630 ( .A1(n1), .A2(n478), .ZN(n382) );
  INV_X1 U631 ( .A(n105), .ZN(n103) );
  OAI22_X1 U632 ( .A1(n419), .A2(n493), .B1(n418), .B2(n475), .ZN(n342) );
  OAI22_X1 U633 ( .A1(n419), .A2(n475), .B1(n493), .B2(n420), .ZN(n343) );
  OAI22_X1 U634 ( .A1(n493), .A2(n411), .B1(n475), .B2(n410), .ZN(n334) );
  AOI21_X1 U635 ( .B1(n493), .B2(n475), .A(n409), .ZN(n283) );
  OAI22_X1 U636 ( .A1(n493), .A2(n410), .B1(n475), .B2(n409), .ZN(n333) );
  OAI22_X1 U637 ( .A1(n418), .A2(n493), .B1(n475), .B2(n417), .ZN(n341) );
  INV_X1 U638 ( .A(n475), .ZN(n284) );
  OAI22_X1 U639 ( .A1(n493), .A2(n416), .B1(n475), .B2(n415), .ZN(n339) );
  OAI22_X1 U640 ( .A1(n493), .A2(n415), .B1(n475), .B2(n414), .ZN(n338) );
  OAI22_X1 U641 ( .A1(n493), .A2(n414), .B1(n475), .B2(n413), .ZN(n337) );
  XOR2_X1 U642 ( .A(a[9]), .B(a[8]), .Z(n461) );
  NOR2_X1 U643 ( .A1(n189), .A2(n196), .ZN(n66) );
  OAI22_X1 U644 ( .A1(n493), .A2(n417), .B1(n416), .B2(n475), .ZN(n340) );
  NOR2_X1 U645 ( .A1(n183), .A2(n188), .ZN(n58) );
  INV_X1 U646 ( .A(n58), .ZN(n56) );
  NAND2_X1 U647 ( .A1(n56), .A2(n59), .ZN(n9) );
  INV_X1 U648 ( .A(n59), .ZN(n57) );
  INV_X1 U649 ( .A(n53), .ZN(n147) );
  XNOR2_X1 U650 ( .A(n1), .B(n487), .ZN(n420) );
  XNOR2_X1 U651 ( .A(n458), .B(n487), .ZN(n419) );
  XNOR2_X1 U652 ( .A(n457), .B(n487), .ZN(n418) );
  INV_X1 U653 ( .A(n487), .ZN(n285) );
  XNOR2_X1 U654 ( .A(n487), .B(n456), .ZN(n417) );
  XNOR2_X1 U655 ( .A(n487), .B(n453), .ZN(n414) );
  NAND2_X1 U656 ( .A1(n225), .A2(n234), .ZN(n94) );
  NAND2_X1 U657 ( .A1(n183), .A2(n188), .ZN(n59) );
  INV_X1 U658 ( .A(n170), .ZN(n171) );
  NAND2_X1 U659 ( .A1(n177), .A2(n182), .ZN(n54) );
  NOR2_X1 U660 ( .A1(n82), .A2(n87), .ZN(n80) );
  OAI21_X1 U661 ( .B1(n582), .B2(n88), .A(n83), .ZN(n81) );
  NAND2_X1 U662 ( .A1(n555), .A2(n574), .ZN(n12) );
  NOR2_X1 U663 ( .A1(n73), .A2(n66), .ZN(n64) );
  NAND2_X1 U664 ( .A1(n150), .A2(n567), .ZN(n11) );
  OAI21_X1 U665 ( .B1(n74), .B2(n66), .A(n67), .ZN(n65) );
  OAI21_X1 U666 ( .B1(n79), .B2(n573), .A(n567), .ZN(n70) );
  NOR2_X1 U667 ( .A1(n197), .A2(n204), .ZN(n73) );
  INV_X1 U668 ( .A(n474), .ZN(n281) );
  OAI21_X1 U669 ( .B1(n585), .B2(n34), .A(n35), .ZN(n33) );
  NAND2_X1 U670 ( .A1(n205), .A2(n214), .ZN(n83) );
  OAI22_X1 U671 ( .A1(n493), .A2(n412), .B1(n475), .B2(n411), .ZN(n335) );
  OAI22_X1 U672 ( .A1(n494), .A2(n423), .B1(n422), .B2(n476), .ZN(n346) );
  OAI22_X1 U673 ( .A1(n494), .A2(n426), .B1(n425), .B2(n476), .ZN(n349) );
  OAI22_X1 U674 ( .A1(n494), .A2(n427), .B1(n426), .B2(n476), .ZN(n350) );
  OAI22_X1 U675 ( .A1(n494), .A2(n428), .B1(n427), .B2(n476), .ZN(n351) );
  OAI22_X1 U676 ( .A1(n494), .A2(n432), .B1(n431), .B2(n476), .ZN(n355) );
  OAI22_X1 U677 ( .A1(n494), .A2(n433), .B1(n432), .B2(n476), .ZN(n356) );
  OAI22_X1 U678 ( .A1(n494), .A2(n431), .B1(n430), .B2(n476), .ZN(n354) );
  OAI22_X1 U679 ( .A1(n494), .A2(n430), .B1(n429), .B2(n476), .ZN(n353) );
  OAI22_X1 U680 ( .A1(n494), .A2(n429), .B1(n428), .B2(n476), .ZN(n352) );
  OAI22_X1 U681 ( .A1(n494), .A2(n482), .B1(n434), .B2(n476), .ZN(n296) );
  INV_X1 U682 ( .A(n289), .ZN(n358) );
  XNOR2_X1 U683 ( .A(n487), .B(n450), .ZN(n411) );
  NOR2_X1 U684 ( .A1(n557), .A2(n96), .ZN(n91) );
  NAND2_X1 U685 ( .A1(n154), .A2(n97), .ZN(n15) );
  OAI21_X1 U686 ( .B1(n93), .B2(n97), .A(n94), .ZN(n92) );
  NOR2_X1 U687 ( .A1(n235), .A2(n242), .ZN(n96) );
  OAI22_X1 U688 ( .A1(n495), .A2(n483), .B1(n447), .B2(n477), .ZN(n297) );
  OAI22_X1 U689 ( .A1(n445), .A2(n477), .B1(n495), .B2(n446), .ZN(n369) );
  OAI22_X1 U690 ( .A1(n495), .A2(n441), .B1(n440), .B2(n477), .ZN(n364) );
  OAI22_X1 U691 ( .A1(n495), .A2(n443), .B1(n442), .B2(n477), .ZN(n366) );
  OAI22_X1 U692 ( .A1(n495), .A2(n442), .B1(n441), .B2(n477), .ZN(n365) );
  OAI22_X1 U693 ( .A1(n495), .A2(n440), .B1(n439), .B2(n477), .ZN(n363) );
  OAI22_X1 U694 ( .A1(n444), .A2(n477), .B1(n445), .B2(n495), .ZN(n368) );
  OAI22_X1 U695 ( .A1(n444), .A2(n495), .B1(n443), .B2(n477), .ZN(n367) );
  XNOR2_X1 U696 ( .A(n484), .B(n453), .ZN(n375) );
  XNOR2_X1 U697 ( .A(n456), .B(n484), .ZN(n378) );
  XNOR2_X1 U698 ( .A(n484), .B(n450), .ZN(n372) );
  NAND2_X1 U699 ( .A1(n589), .A2(n588), .ZN(n100) );
  AOI21_X1 U700 ( .B1(n589), .B2(n108), .A(n103), .ZN(n101) );
  NAND2_X1 U701 ( .A1(n235), .A2(n242), .ZN(n97) );
  OAI21_X1 U702 ( .B1(n581), .B2(n62), .A(n63), .ZN(n61) );
  INV_X1 U703 ( .A(n87), .ZN(n85) );
  NAND2_X1 U704 ( .A1(n85), .A2(n88), .ZN(n13) );
  INV_X1 U705 ( .A(n88), .ZN(n86) );
  NAND2_X1 U706 ( .A1(n64), .A2(n80), .ZN(n62) );
  AOI21_X1 U707 ( .B1(n81), .B2(n64), .A(n65), .ZN(n63) );
  XNOR2_X1 U708 ( .A(n1), .B(n484), .ZN(n381) );
  BUF_X1 U709 ( .A(a[7]), .Z(n596) );
  XNOR2_X1 U710 ( .A(n487), .B(n451), .ZN(n412) );
  XNOR2_X1 U711 ( .A(n484), .B(n587), .ZN(n373) );
  OAI22_X1 U712 ( .A1(n494), .A2(n425), .B1(n424), .B2(n476), .ZN(n348) );
  OAI22_X1 U713 ( .A1(n494), .A2(n424), .B1(n423), .B2(n476), .ZN(n347) );
  XNOR2_X1 U714 ( .A(a[3]), .B(a[4]), .ZN(n499) );
  XNOR2_X1 U715 ( .A(a[1]), .B(a[2]), .ZN(n500) );
  OAI22_X1 U716 ( .A1(n495), .A2(n439), .B1(n438), .B2(n477), .ZN(n362) );
  OAI22_X1 U717 ( .A1(n495), .A2(n438), .B1(n437), .B2(n477), .ZN(n361) );
  XNOR2_X1 U718 ( .A(n487), .B(b[11]), .ZN(n409) );
  XNOR2_X1 U719 ( .A(b[11]), .B(n484), .ZN(n370) );
  XNOR2_X1 U720 ( .A(n458), .B(n484), .ZN(n380) );
  XNOR2_X1 U721 ( .A(n457), .B(n484), .ZN(n379) );
  NAND2_X1 U722 ( .A1(n215), .A2(n224), .ZN(n88) );
  XNOR2_X1 U723 ( .A(n487), .B(b[10]), .ZN(n410) );
  XNOR2_X1 U724 ( .A(n484), .B(b[10]), .ZN(n371) );
  OAI22_X1 U725 ( .A1(n560), .A2(n398), .B1(n474), .B2(n397), .ZN(n322) );
  OAI22_X1 U726 ( .A1(n560), .A2(n397), .B1(n474), .B2(n396), .ZN(n321) );
  AOI21_X1 U727 ( .B1(n560), .B2(n474), .A(n396), .ZN(n280) );
  OAI22_X1 U728 ( .A1(n406), .A2(n474), .B1(n492), .B2(n407), .ZN(n330) );
  OAI22_X1 U729 ( .A1(n405), .A2(n474), .B1(n406), .B2(n560), .ZN(n329) );
  OAI22_X1 U730 ( .A1(n405), .A2(n560), .B1(n474), .B2(n404), .ZN(n328) );
  OAI22_X1 U731 ( .A1(n492), .A2(n399), .B1(n474), .B2(n398), .ZN(n323) );
  OAI22_X1 U732 ( .A1(n492), .A2(n400), .B1(n474), .B2(n399), .ZN(n324) );
  OAI22_X1 U733 ( .A1(n492), .A2(n480), .B1(n408), .B2(n474), .ZN(n294) );
  OAI22_X1 U734 ( .A1(n492), .A2(n402), .B1(n401), .B2(n474), .ZN(n325) );
  XOR2_X1 U735 ( .A(a[1]), .B(a[0]), .Z(n465) );
  INV_X1 U736 ( .A(n472), .ZN(n275) );
  INV_X1 U737 ( .A(n489), .ZN(n483) );
  XNOR2_X1 U738 ( .A(n1), .B(n489), .ZN(n446) );
  XNOR2_X1 U739 ( .A(n458), .B(n489), .ZN(n445) );
  XNOR2_X1 U740 ( .A(n457), .B(n489), .ZN(n444) );
  XNOR2_X1 U741 ( .A(n456), .B(n489), .ZN(n443) );
  XNOR2_X1 U742 ( .A(n489), .B(n453), .ZN(n440) );
  XNOR2_X1 U743 ( .A(n489), .B(n450), .ZN(n437) );
  XNOR2_X1 U744 ( .A(n489), .B(n451), .ZN(n438) );
  XOR2_X1 U745 ( .A(a[5]), .B(a[4]), .Z(n463) );
  OAI22_X1 U746 ( .A1(n493), .A2(n413), .B1(n475), .B2(n412), .ZN(n336) );
  INV_X1 U747 ( .A(n473), .ZN(n278) );
  OAI22_X1 U748 ( .A1(n393), .A2(n473), .B1(n491), .B2(n394), .ZN(n318) );
  OAI22_X1 U749 ( .A1(n392), .A2(n473), .B1(n393), .B2(n491), .ZN(n317) );
  OAI22_X1 U750 ( .A1(n392), .A2(n491), .B1(n391), .B2(n473), .ZN(n316) );
  OAI22_X1 U751 ( .A1(n491), .A2(n391), .B1(n390), .B2(n473), .ZN(n315) );
  OAI22_X1 U752 ( .A1(n390), .A2(n491), .B1(n389), .B2(n473), .ZN(n314) );
  OAI22_X1 U753 ( .A1(n491), .A2(n389), .B1(n388), .B2(n473), .ZN(n313) );
  OAI22_X1 U754 ( .A1(n491), .A2(n388), .B1(n387), .B2(n473), .ZN(n312) );
  OAI22_X1 U755 ( .A1(n491), .A2(n387), .B1(n386), .B2(n473), .ZN(n311) );
  OAI22_X1 U756 ( .A1(n491), .A2(n386), .B1(n385), .B2(n473), .ZN(n310) );
  OAI22_X1 U757 ( .A1(n491), .A2(n385), .B1(n384), .B2(n473), .ZN(n309) );
  OAI22_X1 U758 ( .A1(n491), .A2(n384), .B1(n383), .B2(n473), .ZN(n308) );
  AOI21_X1 U759 ( .B1(n491), .B2(n473), .A(n383), .ZN(n277) );
  OAI22_X1 U760 ( .A1(n491), .A2(n279), .B1(n395), .B2(n473), .ZN(n293) );
  AND2_X1 U761 ( .A1(n1), .A2(n278), .ZN(n319) );
  OR2_X1 U762 ( .A1(n315), .A2(n325), .ZN(n222) );
  XNOR2_X1 U763 ( .A(n315), .B(n325), .ZN(n223) );
  INV_X1 U764 ( .A(n277), .ZN(n307) );
  AOI21_X1 U765 ( .B1(n495), .B2(n477), .A(n435), .ZN(n289) );
  XOR2_X1 U766 ( .A(a[3]), .B(a[2]), .Z(n464) );
  OAI22_X1 U767 ( .A1(n492), .A2(n404), .B1(n403), .B2(n474), .ZN(n327) );
  OAI22_X1 U768 ( .A1(n403), .A2(n492), .B1(n474), .B2(n402), .ZN(n326) );
  XNOR2_X1 U769 ( .A(n489), .B(b[11]), .ZN(n435) );
  OAI22_X1 U770 ( .A1(n495), .A2(n437), .B1(n436), .B2(n477), .ZN(n360) );
  OAI22_X1 U771 ( .A1(n495), .A2(n436), .B1(n435), .B2(n477), .ZN(n359) );
  XNOR2_X1 U772 ( .A(n489), .B(b[10]), .ZN(n436) );
  OAI21_X1 U773 ( .B1(n100), .B2(n112), .A(n101), .ZN(n99) );
  OAI22_X1 U774 ( .A1(n490), .A2(n377), .B1(n472), .B2(n376), .ZN(n194) );
  INV_X1 U775 ( .A(n194), .ZN(n195) );
  XNOR2_X1 U776 ( .A(a[7]), .B(a[8]), .ZN(n497) );
  XNOR2_X1 U777 ( .A(n489), .B(b[5]), .ZN(n441) );
  XNOR2_X1 U778 ( .A(n487), .B(b[5]), .ZN(n415) );
  XNOR2_X1 U779 ( .A(n484), .B(b[5]), .ZN(n376) );
  XNOR2_X1 U780 ( .A(b[4]), .B(n489), .ZN(n442) );
  XNOR2_X1 U781 ( .A(b[4]), .B(n487), .ZN(n416) );
  XNOR2_X1 U782 ( .A(b[4]), .B(n484), .ZN(n377) );
  INV_X1 U783 ( .A(n180), .ZN(n181) );
  OAI22_X1 U784 ( .A1(n490), .A2(n375), .B1(n472), .B2(n374), .ZN(n180) );
  XOR2_X1 U785 ( .A(a[11]), .B(a[10]), .Z(n460) );
  OAI22_X1 U786 ( .A1(n379), .A2(n472), .B1(n380), .B2(n490), .ZN(n304) );
  OAI22_X1 U787 ( .A1(n380), .A2(n472), .B1(n490), .B2(n381), .ZN(n305) );
  OAI22_X1 U788 ( .A1(n379), .A2(n490), .B1(n378), .B2(n472), .ZN(n303) );
  OAI22_X1 U789 ( .A1(n490), .A2(n376), .B1(n472), .B2(n375), .ZN(n301) );
  OAI22_X1 U790 ( .A1(n490), .A2(n374), .B1(n472), .B2(n373), .ZN(n300) );
  AOI21_X1 U791 ( .B1(n490), .B2(n472), .A(n370), .ZN(n274) );
  OAI22_X1 U792 ( .A1(n490), .A2(n372), .B1(n472), .B2(n371), .ZN(n299) );
  OAI22_X1 U793 ( .A1(n490), .A2(n373), .B1(n472), .B2(n372), .ZN(n170) );
  OAI22_X1 U794 ( .A1(n490), .A2(n378), .B1(n377), .B2(n472), .ZN(n302) );
  XNOR2_X1 U795 ( .A(n489), .B(n452), .ZN(n439) );
  XNOR2_X1 U796 ( .A(n487), .B(n452), .ZN(n413) );
  XNOR2_X1 U797 ( .A(n484), .B(n452), .ZN(n374) );
  NAND2_X1 U798 ( .A1(n369), .A2(n297), .ZN(n141) );
  XNOR2_X1 U799 ( .A(n564), .B(n562), .ZN(n433) );
  INV_X1 U800 ( .A(n561), .ZN(n482) );
  XNOR2_X1 U801 ( .A(n458), .B(n562), .ZN(n432) );
  XNOR2_X1 U802 ( .A(n457), .B(n563), .ZN(n431) );
  XNOR2_X1 U803 ( .A(n563), .B(n456), .ZN(n430) );
  XNOR2_X1 U804 ( .A(n563), .B(b[5]), .ZN(n428) );
  XNOR2_X1 U805 ( .A(b[4]), .B(n563), .ZN(n429) );
  XNOR2_X1 U806 ( .A(n562), .B(n451), .ZN(n425) );
  XNOR2_X1 U807 ( .A(n562), .B(n452), .ZN(n426) );
  XNOR2_X1 U808 ( .A(n563), .B(n453), .ZN(n427) );
  XNOR2_X1 U809 ( .A(n562), .B(b[11]), .ZN(n422) );
  XNOR2_X1 U810 ( .A(n562), .B(n450), .ZN(n424) );
  XNOR2_X1 U811 ( .A(n563), .B(b[10]), .ZN(n423) );
  XNOR2_X1 U812 ( .A(a[9]), .B(a[10]), .ZN(n496) );
  OAI22_X1 U813 ( .A1(n493), .A2(n285), .B1(n421), .B2(n475), .ZN(n295) );
  OAI22_X1 U814 ( .A1(n490), .A2(n478), .B1(n382), .B2(n472), .ZN(n292) );
  INV_X1 U815 ( .A(n484), .ZN(n478) );
  INV_X1 U816 ( .A(n212), .ZN(n213) );
  OAI22_X1 U817 ( .A1(n492), .A2(n401), .B1(n474), .B2(n400), .ZN(n212) );
  INV_X1 U818 ( .A(n134), .ZN(n133) );
  AOI21_X1 U819 ( .B1(n592), .B2(n565), .A(n136), .ZN(n134) );
  INV_X1 U820 ( .A(a[0]), .ZN(n501) );
  INV_X1 U821 ( .A(n132), .ZN(n130) );
  XNOR2_X1 U822 ( .A(a[5]), .B(a[6]), .ZN(n498) );
  XNOR2_X1 U823 ( .A(n597), .B(b[10]), .ZN(n397) );
  XNOR2_X1 U824 ( .A(n597), .B(b[11]), .ZN(n396) );
  INV_X1 U825 ( .A(n597), .ZN(n480) );
  XNOR2_X1 U826 ( .A(n597), .B(n451), .ZN(n399) );
  XNOR2_X1 U827 ( .A(n597), .B(n450), .ZN(n398) );
  XNOR2_X1 U828 ( .A(n457), .B(n597), .ZN(n405) );
  XNOR2_X1 U829 ( .A(n1), .B(n597), .ZN(n407) );
  XNOR2_X1 U830 ( .A(n458), .B(n597), .ZN(n406) );
  XNOR2_X1 U831 ( .A(n456), .B(n597), .ZN(n404) );
  XNOR2_X1 U832 ( .A(b[4]), .B(n596), .ZN(n403) );
  XNOR2_X1 U833 ( .A(n596), .B(b[5]), .ZN(n402) );
  XNOR2_X1 U834 ( .A(n597), .B(n453), .ZN(n401) );
  XNOR2_X1 U835 ( .A(n597), .B(n452), .ZN(n400) );
  XOR2_X1 U836 ( .A(a[7]), .B(a[6]), .Z(n462) );
  NAND2_X1 U837 ( .A1(n197), .A2(n204), .ZN(n74) );
  XNOR2_X1 U838 ( .A(n485), .B(b[11]), .ZN(n383) );
  XNOR2_X1 U839 ( .A(n485), .B(b[10]), .ZN(n384) );
  XNOR2_X1 U840 ( .A(n485), .B(n587), .ZN(n386) );
  XNOR2_X1 U841 ( .A(n485), .B(n450), .ZN(n385) );
  XNOR2_X1 U842 ( .A(n485), .B(n452), .ZN(n387) );
  XNOR2_X1 U843 ( .A(n485), .B(n453), .ZN(n388) );
  XNOR2_X1 U844 ( .A(n1), .B(n485), .ZN(n394) );
  XNOR2_X1 U845 ( .A(n458), .B(n485), .ZN(n393) );
  XNOR2_X1 U846 ( .A(n457), .B(n485), .ZN(n392) );
  XNOR2_X1 U847 ( .A(n485), .B(b[5]), .ZN(n389) );
  XNOR2_X1 U848 ( .A(n456), .B(n485), .ZN(n391) );
  XNOR2_X1 U849 ( .A(b[4]), .B(n485), .ZN(n390) );
  INV_X1 U850 ( .A(n485), .ZN(n279) );
  OAI21_X1 U851 ( .B1(n126), .B2(n128), .A(n127), .ZN(n125) );
  AOI21_X1 U852 ( .B1(n117), .B2(n593), .A(n114), .ZN(n112) );
  OAI21_X1 U853 ( .B1(n118), .B2(n120), .A(n119), .ZN(n117) );
  AND2_X1 U854 ( .A1(n564), .A2(a[0]), .ZN(product[0]) );
  XNOR2_X1 U855 ( .A(n23), .B(n565), .ZN(product[2]) );
  NAND2_X1 U856 ( .A1(n592), .A2(n138), .ZN(n23) );
  XOR2_X1 U857 ( .A(n21), .B(n128), .Z(product[4]) );
  NAND2_X1 U858 ( .A1(n160), .A2(n127), .ZN(n21) );
  XNOR2_X1 U859 ( .A(n22), .B(n133), .ZN(product[3]) );
  NAND2_X1 U860 ( .A1(n591), .A2(n132), .ZN(n22) );
  XOR2_X1 U861 ( .A(n19), .B(n120), .Z(product[6]) );
  NAND2_X1 U862 ( .A1(n158), .A2(n119), .ZN(n19) );
  AOI21_X1 U863 ( .B1(n594), .B2(n125), .A(n566), .ZN(n120) );
  XNOR2_X1 U864 ( .A(n20), .B(n125), .ZN(product[5]) );
  NAND2_X1 U865 ( .A1(n594), .A2(n124), .ZN(n20) );
  XNOR2_X1 U866 ( .A(n117), .B(n18), .ZN(product[7]) );
  NAND2_X1 U867 ( .A1(n593), .A2(n116), .ZN(n18) );
  INV_X1 U868 ( .A(n112), .ZN(n111) );
  XOR2_X1 U869 ( .A(n106), .B(n16), .Z(product[9]) );
  AOI21_X1 U870 ( .B1(n111), .B2(n588), .A(n108), .ZN(n106) );
  INV_X1 U871 ( .A(n99), .ZN(n98) );
  XNOR2_X1 U872 ( .A(n95), .B(n14), .ZN(product[11]) );
  OAI21_X1 U873 ( .B1(n98), .B2(n96), .A(n97), .ZN(n95) );
  AOI21_X1 U874 ( .B1(n586), .B2(n37), .A(n38), .ZN(n36) );
  XNOR2_X1 U875 ( .A(n89), .B(n13), .ZN(product[12]) );
  INV_X1 U876 ( .A(n90), .ZN(n89) );
  AOI21_X1 U877 ( .B1(n61), .B2(n56), .A(n57), .ZN(n55) );
  XNOR2_X1 U878 ( .A(n33), .B(n4), .ZN(product[21]) );
  XOR2_X1 U879 ( .A(n75), .B(n11), .Z(product[14]) );
  AOI21_X1 U880 ( .B1(n89), .B2(n76), .A(n77), .ZN(n75) );
  XNOR2_X1 U881 ( .A(n48), .B(n7), .ZN(product[18]) );
  OAI21_X1 U882 ( .B1(n60), .B2(n49), .A(n50), .ZN(n48) );
  AOI21_X1 U883 ( .B1(n69), .B2(n89), .A(n70), .ZN(n68) );
  XNOR2_X1 U884 ( .A(n41), .B(n6), .ZN(product[19]) );
  OAI21_X1 U885 ( .B1(n556), .B2(n42), .A(n43), .ZN(n41) );
  XOR2_X1 U886 ( .A(n84), .B(n12), .Z(product[13]) );
  AOI21_X1 U887 ( .B1(n89), .B2(n85), .A(n86), .ZN(n84) );
  XOR2_X1 U888 ( .A(n60), .B(n9), .Z(product[16]) );
  INV_X1 U889 ( .A(n61), .ZN(n60) );
  XOR2_X1 U890 ( .A(n28), .B(n3), .Z(product[22]) );
  AOI21_X1 U891 ( .B1(n33), .B2(n554), .A(n30), .ZN(n28) );
  INV_X1 U892 ( .A(n25), .ZN(product[23]) );
  OAI21_X1 U893 ( .B1(n559), .B2(n26), .A(n27), .ZN(n25) );
endmodule


module datapath_DW_mult_tc_21 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n1, n3, n4, n6, n7, n8, n9, n10, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n25, n26, n27, n28, n30, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n45, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n95, n96,
         n98, n100, n101, n102, n104, n106, n107, n108, n109, n110, n112, n114,
         n115, n116, n117, n118, n120, n122, n123, n124, n126, n128, n129,
         n131, n132, n134, n135, n137, n138, n139, n140, n141, n143, n144,
         n148, n150, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n259, n260, n261, n262, n263,
         n264, n265, n267, n268, n269, n270, n271, n273, n274, n275, n276,
         n277, n278, n279, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n450, n451, n452, n453, n454, n455,
         n458, n460, n462, n463, n464, n465, n466, n467, n468, n470, n473,
         n476, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n602, n603, n604, n605;

  FA_X1 U178 ( .A(n289), .B(n160), .CI(n298), .CO(n156), .S(n157) );
  FA_X1 U179 ( .A(n161), .B(n299), .CI(n164), .CO(n158), .S(n159) );
  FA_X1 U181 ( .A(n168), .B(n311), .CI(n165), .CO(n162), .S(n163) );
  FA_X1 U182 ( .A(n290), .B(n170), .CI(n300), .CO(n164), .S(n165) );
  FA_X1 U183 ( .A(n169), .B(n176), .CI(n174), .CO(n166), .S(n167) );
  FA_X1 U184 ( .A(n312), .B(n301), .CI(n171), .CO(n168), .S(n169) );
  FA_X1 U186 ( .A(n180), .B(n177), .CI(n175), .CO(n172), .S(n173) );
  FA_X1 U187 ( .A(n323), .B(n302), .CI(n182), .CO(n174), .S(n175) );
  FA_X1 U188 ( .A(n291), .B(n184), .CI(n313), .CO(n176), .S(n177) );
  FA_X1 U189 ( .A(n188), .B(n183), .CI(n181), .CO(n178), .S(n179) );
  FA_X1 U190 ( .A(n192), .B(n324), .CI(n190), .CO(n180), .S(n181) );
  FA_X1 U191 ( .A(n292), .B(n303), .CI(n185), .CO(n182), .S(n183) );
  FA_X1 U193 ( .A(n196), .B(n191), .CI(n189), .CO(n186), .S(n187) );
  FA_X1 U194 ( .A(n193), .B(n200), .CI(n198), .CO(n188), .S(n189) );
  FA_X1 U195 ( .A(n304), .B(n293), .CI(n335), .CO(n190), .S(n191) );
  FA_X1 U196 ( .A(n314), .B(n570), .CI(n325), .CO(n192), .S(n193) );
  FA_X1 U197 ( .A(n206), .B(n199), .CI(n197), .CO(n194), .S(n195) );
  FA_X1 U198 ( .A(n201), .B(n210), .CI(n208), .CO(n196), .S(n197) );
  FA_X1 U199 ( .A(n336), .B(n305), .CI(n212), .CO(n198), .S(n199) );
  FA_X1 U200 ( .A(n315), .B(n294), .CI(n203), .CO(n200), .S(n201) );
  FA_X1 U202 ( .A(n216), .B(n209), .CI(n207), .CO(n204), .S(n205) );
  FA_X1 U203 ( .A(n211), .B(n220), .CI(n218), .CO(n206), .S(n207) );
  FA_X1 U204 ( .A(n545), .B(n348), .CI(n213), .CO(n208), .S(n209) );
  FA_X1 U205 ( .A(n295), .B(n306), .CI(n337), .CO(n210), .S(n211) );
  FA_X1 U209 ( .A(n228), .B(n230), .CI(n221), .CO(n216), .S(n217) );
  FA_X1 U210 ( .A(n349), .B(n307), .CI(n223), .CO(n218), .S(n219) );
  FA_X1 U211 ( .A(n317), .B(n282), .CI(n296), .CO(n220), .S(n221) );
  FA_X1 U213 ( .A(n234), .B(n229), .CI(n227), .CO(n224), .S(n225) );
  FA_X1 U214 ( .A(n236), .B(n238), .CI(n231), .CO(n226), .S(n227) );
  FA_X1 U215 ( .A(n308), .B(n350), .CI(n318), .CO(n228), .S(n229) );
  FA_X1 U216 ( .A(n339), .B(n297), .CI(n328), .CO(n230), .S(n231) );
  FA_X1 U218 ( .A(n239), .B(n283), .CI(n244), .CO(n234), .S(n235) );
  FA_X1 U219 ( .A(n329), .B(n319), .CI(n309), .CO(n236), .S(n237) );
  HA_X1 U220 ( .A(n351), .B(n340), .CO(n238), .S(n239) );
  FA_X1 U221 ( .A(n245), .B(n248), .CI(n243), .CO(n240), .S(n241) );
  FA_X1 U222 ( .A(n320), .B(n330), .CI(n250), .CO(n242), .S(n243) );
  FA_X1 U223 ( .A(n341), .B(n310), .CI(n352), .CO(n244), .S(n245) );
  FA_X1 U224 ( .A(n254), .B(n251), .CI(n249), .CO(n246), .S(n247) );
  FA_X1 U225 ( .A(n321), .B(n331), .CI(n342), .CO(n248), .S(n249) );
  HA_X1 U226 ( .A(n284), .B(n353), .CO(n250), .S(n251) );
  FA_X1 U227 ( .A(n543), .B(n332), .CI(n255), .CO(n252), .S(n253) );
  FA_X1 U228 ( .A(n354), .B(n322), .CI(n343), .CO(n254), .S(n255) );
  FA_X1 U229 ( .A(n355), .B(n333), .CI(n259), .CO(n256), .S(n257) );
  FA_X1 U231 ( .A(n345), .B(n334), .CI(n356), .CO(n260), .S(n261) );
  HA_X1 U232 ( .A(n357), .B(n286), .CO(n262), .S(n263) );
  CLKBUF_X3 U468 ( .A(n488), .Z(n464) );
  BUF_X2 U469 ( .A(n482), .Z(n458) );
  BUF_X2 U470 ( .A(a[1]), .Z(n479) );
  BUF_X1 U471 ( .A(a[9]), .Z(n603) );
  BUF_X1 U472 ( .A(n480), .Z(n566) );
  BUF_X2 U473 ( .A(n490), .Z(n466) );
  OR2_X2 U474 ( .A1(n233), .A2(n240), .ZN(n574) );
  BUF_X2 U475 ( .A(a[3]), .Z(n478) );
  BUF_X1 U476 ( .A(b[10]), .Z(n439) );
  BUF_X2 U477 ( .A(a[11]), .Z(n564) );
  BUF_X1 U478 ( .A(n484), .Z(n460) );
  BUF_X2 U479 ( .A(n486), .Z(n462) );
  AOI21_X1 U480 ( .B1(n598), .B2(n115), .A(n112), .ZN(n110) );
  AND2_X1 U481 ( .A1(n344), .A2(n285), .ZN(n543) );
  AND2_X1 U482 ( .A1(n451), .A2(n487), .ZN(n600) );
  OR2_X1 U483 ( .A1(n163), .A2(n166), .ZN(n544) );
  AND2_X1 U484 ( .A1(n338), .A2(n327), .ZN(n545) );
  OR2_X1 U485 ( .A1(n156), .A2(n155), .ZN(n546) );
  BUF_X2 U486 ( .A(n487), .Z(n463) );
  CLKBUF_X1 U487 ( .A(n68), .Z(n547) );
  BUF_X2 U488 ( .A(n489), .Z(n465) );
  XOR2_X1 U489 ( .A(n226), .B(n219), .Z(n548) );
  XOR2_X1 U490 ( .A(n217), .B(n548), .Z(n215) );
  NAND2_X1 U491 ( .A1(n217), .A2(n226), .ZN(n549) );
  NAND2_X1 U492 ( .A1(n217), .A2(n219), .ZN(n550) );
  NAND2_X1 U493 ( .A1(n226), .A2(n219), .ZN(n551) );
  NAND3_X1 U494 ( .A1(n549), .A2(n550), .A3(n551), .ZN(n214) );
  CLKBUF_X3 U495 ( .A(n482), .Z(n578) );
  BUF_X2 U496 ( .A(b[8]), .Z(n441) );
  BUF_X2 U497 ( .A(a[5]), .Z(n604) );
  CLKBUF_X1 U498 ( .A(b[11]), .Z(n552) );
  CLKBUF_X1 U499 ( .A(b[11]), .Z(n553) );
  BUF_X2 U500 ( .A(b[7]), .Z(n442) );
  CLKBUF_X1 U501 ( .A(n483), .Z(n554) );
  XOR2_X1 U502 ( .A(n344), .B(n285), .Z(n259) );
  BUF_X2 U503 ( .A(b[0]), .Z(n1) );
  BUF_X2 U504 ( .A(b[9]), .Z(n440) );
  XOR2_X1 U505 ( .A(n237), .B(n242), .Z(n555) );
  XOR2_X1 U506 ( .A(n235), .B(n555), .Z(n233) );
  NAND2_X1 U507 ( .A1(n235), .A2(n237), .ZN(n556) );
  NAND2_X1 U508 ( .A1(n235), .A2(n242), .ZN(n557) );
  NAND2_X1 U509 ( .A1(n237), .A2(n242), .ZN(n558) );
  NAND3_X1 U510 ( .A1(n556), .A2(n557), .A3(n558), .ZN(n232) );
  INV_X1 U511 ( .A(n271), .ZN(n559) );
  INV_X1 U512 ( .A(n470), .ZN(n560) );
  CLKBUF_X1 U513 ( .A(n478), .Z(n561) );
  CLKBUF_X1 U514 ( .A(n107), .Z(n562) );
  CLKBUF_X1 U515 ( .A(n77), .Z(n563) );
  INV_X1 U516 ( .A(n600), .ZN(n565) );
  INV_X1 U517 ( .A(n600), .ZN(n481) );
  CLKBUF_X1 U518 ( .A(n1), .Z(n567) );
  AOI21_X1 U519 ( .B1(n107), .B2(n597), .A(n104), .ZN(n568) );
  CLKBUF_X1 U520 ( .A(n115), .Z(n569) );
  OAI22_X1 U521 ( .A1(n483), .A2(n402), .B1(n401), .B2(n465), .ZN(n570) );
  INV_X1 U522 ( .A(n278), .ZN(n571) );
  CLKBUF_X1 U523 ( .A(n465), .Z(n572) );
  CLKBUF_X1 U524 ( .A(n483), .Z(n573) );
  BUF_X2 U525 ( .A(n484), .Z(n584) );
  BUF_X1 U526 ( .A(a[5]), .Z(n605) );
  BUF_X2 U527 ( .A(b[1]), .Z(n448) );
  INV_X1 U528 ( .A(n579), .ZN(n95) );
  XNOR2_X1 U529 ( .A(n442), .B(n604), .ZN(n575) );
  CLKBUF_X1 U530 ( .A(b[4]), .Z(n445) );
  CLKBUF_X1 U531 ( .A(b[2]), .Z(n576) );
  CLKBUF_X1 U532 ( .A(b[2]), .Z(n447) );
  BUF_X2 U533 ( .A(b[3]), .Z(n446) );
  XOR2_X1 U534 ( .A(n338), .B(n327), .Z(n223) );
  CLKBUF_X3 U535 ( .A(b[6]), .Z(n443) );
  XNOR2_X1 U536 ( .A(n69), .B(n577), .ZN(product[14]) );
  AND2_X1 U537 ( .A1(n140), .A2(n547), .ZN(n577) );
  AND2_X1 U538 ( .A1(n233), .A2(n240), .ZN(n579) );
  CLKBUF_X1 U539 ( .A(n73), .Z(n580) );
  NAND2_X1 U540 ( .A1(n450), .A2(n486), .ZN(n480) );
  CLKBUF_X1 U541 ( .A(n59), .Z(n588) );
  NOR2_X1 U542 ( .A1(n563), .A2(n585), .ZN(n581) );
  NOR2_X1 U543 ( .A1(n195), .A2(n204), .ZN(n582) );
  CLKBUF_X1 U544 ( .A(n78), .Z(n583) );
  CLKBUF_X1 U545 ( .A(n72), .Z(n585) );
  NOR2_X1 U546 ( .A1(n195), .A2(n204), .ZN(n72) );
  CLKBUF_X1 U547 ( .A(n67), .Z(n586) );
  NOR2_X1 U548 ( .A1(n187), .A2(n194), .ZN(n67) );
  CLKBUF_X1 U549 ( .A(n71), .Z(n587) );
  AOI21_X1 U550 ( .B1(n89), .B2(n81), .A(n82), .ZN(n589) );
  BUF_X2 U551 ( .A(n445), .Z(n590) );
  NOR2_X1 U552 ( .A1(n179), .A2(n186), .ZN(n591) );
  NOR2_X1 U553 ( .A1(n215), .A2(n224), .ZN(n592) );
  XNOR2_X1 U554 ( .A(n85), .B(n14), .ZN(product[11]) );
  XNOR2_X1 U555 ( .A(n101), .B(n17), .ZN(product[8]) );
  XNOR2_X1 U556 ( .A(n36), .B(n593), .ZN(product[20]) );
  AND2_X1 U557 ( .A1(n134), .A2(n35), .ZN(n593) );
  OR2_X1 U558 ( .A1(n241), .A2(n246), .ZN(n594) );
  OR2_X1 U559 ( .A1(n263), .A2(n346), .ZN(n595) );
  OR2_X1 U560 ( .A1(n358), .A2(n347), .ZN(n596) );
  OR2_X1 U561 ( .A1(n247), .A2(n252), .ZN(n597) );
  OR2_X1 U562 ( .A1(n257), .A2(n260), .ZN(n598) );
  OR2_X1 U563 ( .A1(n359), .A2(n287), .ZN(n599) );
  BUF_X1 U564 ( .A(a[9]), .Z(n602) );
  AND2_X1 U565 ( .A1(n599), .A2(n131), .ZN(product[1]) );
  NOR2_X1 U566 ( .A1(n288), .A2(n154), .ZN(n26) );
  NAND2_X1 U567 ( .A1(n546), .A2(n32), .ZN(n4) );
  INV_X1 U568 ( .A(n32), .ZN(n30) );
  NOR2_X1 U569 ( .A1(n158), .A2(n157), .ZN(n34) );
  NAND2_X1 U570 ( .A1(n132), .A2(n27), .ZN(n3) );
  INV_X1 U571 ( .A(n26), .ZN(n132) );
  NAND2_X1 U572 ( .A1(n156), .A2(n155), .ZN(n32) );
  INV_X1 U573 ( .A(n39), .ZN(n135) );
  INV_X1 U574 ( .A(n34), .ZN(n134) );
  NAND2_X1 U575 ( .A1(n158), .A2(n157), .ZN(n35) );
  NOR2_X1 U576 ( .A1(n159), .A2(n162), .ZN(n39) );
  NAND2_X1 U577 ( .A1(n135), .A2(n40), .ZN(n6) );
  NAND2_X1 U578 ( .A1(n159), .A2(n162), .ZN(n40) );
  BUF_X2 U579 ( .A(n491), .Z(n467) );
  INV_X1 U580 ( .A(n602), .ZN(n269) );
  INV_X1 U581 ( .A(n273), .ZN(n323) );
  AOI21_X1 U582 ( .B1(n565), .B2(n463), .A(n373), .ZN(n267) );
  XNOR2_X1 U583 ( .A(n602), .B(n446), .ZN(n381) );
  CLKBUF_X3 U584 ( .A(a[7]), .Z(n476) );
  NAND2_X1 U585 ( .A1(n594), .A2(n100), .ZN(n17) );
  XNOR2_X1 U586 ( .A(n552), .B(n602), .ZN(n373) );
  CLKBUF_X1 U587 ( .A(b[11]), .Z(n438) );
  XOR2_X1 U588 ( .A(a[9]), .B(a[8]), .Z(n451) );
  XOR2_X1 U589 ( .A(a[10]), .B(a[11]), .Z(n450) );
  NAND2_X2 U590 ( .A1(n455), .A2(n491), .ZN(n485) );
  OAI22_X1 U591 ( .A1(n485), .A2(n473), .B1(n437), .B2(n467), .ZN(n287) );
  AND2_X1 U592 ( .A1(n567), .A2(n277), .ZN(n347) );
  OAI22_X1 U593 ( .A1(n422), .A2(n466), .B1(n584), .B2(n423), .ZN(n346) );
  OAI22_X1 U594 ( .A1(n424), .A2(n466), .B1(n460), .B2(n278), .ZN(n286) );
  NAND2_X1 U595 ( .A1(n241), .A2(n246), .ZN(n100) );
  XNOR2_X1 U596 ( .A(n602), .B(n441), .ZN(n376) );
  XNOR2_X1 U597 ( .A(n448), .B(n603), .ZN(n383) );
  OAI22_X1 U598 ( .A1(n481), .A2(n377), .B1(n376), .B2(n463), .ZN(n302) );
  OAI22_X1 U599 ( .A1(n565), .A2(n376), .B1(n375), .B2(n463), .ZN(n301) );
  OAI22_X1 U600 ( .A1(n565), .A2(n375), .B1(n374), .B2(n463), .ZN(n300) );
  OAI22_X1 U601 ( .A1(n565), .A2(n374), .B1(n373), .B2(n463), .ZN(n299) );
  OAI22_X1 U602 ( .A1(n481), .A2(n269), .B1(n385), .B2(n463), .ZN(n283) );
  INV_X1 U603 ( .A(n267), .ZN(n298) );
  INV_X1 U604 ( .A(n53), .ZN(n137) );
  OAI22_X1 U605 ( .A1(n481), .A2(n379), .B1(n378), .B2(n463), .ZN(n304) );
  NOR2_X1 U606 ( .A1(n173), .A2(n178), .ZN(n56) );
  OAI22_X1 U607 ( .A1(n485), .A2(n428), .B1(n427), .B2(n467), .ZN(n351) );
  XNOR2_X1 U608 ( .A(n603), .B(n440), .ZN(n375) );
  NAND2_X1 U609 ( .A1(n253), .A2(n256), .ZN(n109) );
  INV_X1 U610 ( .A(n465), .ZN(n274) );
  NAND2_X2 U611 ( .A1(n489), .A2(n453), .ZN(n483) );
  OAI22_X1 U612 ( .A1(n413), .A2(n584), .B1(n412), .B2(n466), .ZN(n336) );
  XNOR2_X1 U613 ( .A(n439), .B(n603), .ZN(n374) );
  NOR2_X1 U614 ( .A1(n225), .A2(n232), .ZN(n86) );
  NAND2_X1 U615 ( .A1(n261), .A2(n262), .ZN(n117) );
  OAI21_X1 U616 ( .B1(n88), .B2(n86), .A(n87), .ZN(n85) );
  NAND2_X1 U617 ( .A1(n141), .A2(n580), .ZN(n12) );
  INV_X1 U618 ( .A(n106), .ZN(n104) );
  OAI22_X1 U619 ( .A1(n380), .A2(n565), .B1(n379), .B2(n463), .ZN(n305) );
  OAI22_X1 U620 ( .A1(n432), .A2(n467), .B1(n485), .B2(n433), .ZN(n356) );
  NAND2_X1 U621 ( .A1(n544), .A2(n47), .ZN(n7) );
  INV_X1 U622 ( .A(n47), .ZN(n45) );
  INV_X1 U623 ( .A(n279), .ZN(n348) );
  AOI21_X1 U624 ( .B1(n485), .B2(n467), .A(n425), .ZN(n279) );
  NAND2_X1 U625 ( .A1(n263), .A2(n346), .ZN(n122) );
  OAI22_X1 U626 ( .A1(n565), .A2(n384), .B1(n383), .B2(n463), .ZN(n309) );
  INV_X1 U627 ( .A(n114), .ZN(n112) );
  OAI22_X1 U628 ( .A1(n421), .A2(n466), .B1(n422), .B2(n584), .ZN(n345) );
  NAND2_X1 U629 ( .A1(n247), .A2(n252), .ZN(n106) );
  INV_X1 U630 ( .A(n100), .ZN(n98) );
  OAI22_X1 U631 ( .A1(n380), .A2(n463), .B1(n481), .B2(n381), .ZN(n306) );
  NAND2_X1 U632 ( .A1(n137), .A2(n54), .ZN(n8) );
  NOR2_X1 U633 ( .A1(n167), .A2(n172), .ZN(n53) );
  NOR2_X1 U634 ( .A1(n253), .A2(n256), .ZN(n108) );
  NAND2_X1 U635 ( .A1(n163), .A2(n166), .ZN(n47) );
  NAND2_X1 U636 ( .A1(n167), .A2(n172), .ZN(n54) );
  OAI22_X1 U637 ( .A1(n419), .A2(n466), .B1(n584), .B2(n420), .ZN(n343) );
  NOR2_X1 U638 ( .A1(n42), .A2(n39), .ZN(n37) );
  XNOR2_X1 U639 ( .A(n590), .B(n602), .ZN(n380) );
  NOR2_X1 U640 ( .A1(n56), .A2(n53), .ZN(n51) );
  INV_X1 U641 ( .A(n64), .ZN(n139) );
  OAI22_X1 U642 ( .A1(n408), .A2(n572), .B1(n409), .B2(n573), .ZN(n332) );
  OAI22_X1 U643 ( .A1(n400), .A2(n573), .B1(n399), .B2(n572), .ZN(n324) );
  OAI22_X1 U644 ( .A1(n409), .A2(n465), .B1(n573), .B2(n410), .ZN(n333) );
  AOI21_X1 U645 ( .B1(n554), .B2(n572), .A(n399), .ZN(n273) );
  OAI22_X1 U646 ( .A1(n406), .A2(n483), .B1(n405), .B2(n465), .ZN(n329) );
  OAI22_X1 U647 ( .A1(n408), .A2(n554), .B1(n407), .B2(n465), .ZN(n331) );
  OAI22_X1 U648 ( .A1(n405), .A2(n483), .B1(n465), .B2(n404), .ZN(n328) );
  OAI22_X1 U649 ( .A1(n411), .A2(n465), .B1(n483), .B2(n275), .ZN(n285) );
  OAI22_X1 U650 ( .A1(n404), .A2(n483), .B1(n465), .B2(n575), .ZN(n327) );
  XNOR2_X1 U651 ( .A(n443), .B(n604), .ZN(n404) );
  OAI22_X1 U652 ( .A1(n432), .A2(n485), .B1(n431), .B2(n467), .ZN(n355) );
  OAI22_X1 U653 ( .A1(n431), .A2(n485), .B1(n430), .B2(n467), .ZN(n354) );
  INV_X1 U654 ( .A(n592), .ZN(n143) );
  INV_X1 U655 ( .A(n464), .ZN(n271) );
  OAI22_X1 U656 ( .A1(n396), .A2(n464), .B1(n578), .B2(n397), .ZN(n321) );
  OAI22_X1 U657 ( .A1(n395), .A2(n464), .B1(n396), .B2(n578), .ZN(n320) );
  OAI22_X1 U658 ( .A1(n395), .A2(n578), .B1(n394), .B2(n464), .ZN(n319) );
  OAI22_X1 U659 ( .A1(n458), .A2(n391), .B1(n390), .B2(n464), .ZN(n315) );
  OAI22_X1 U660 ( .A1(n458), .A2(n390), .B1(n389), .B2(n464), .ZN(n314) );
  OAI22_X1 U661 ( .A1(n387), .A2(n559), .B1(n578), .B2(n388), .ZN(n313) );
  OAI22_X1 U662 ( .A1(n387), .A2(n578), .B1(n386), .B2(n559), .ZN(n312) );
  AOI21_X1 U663 ( .B1(n578), .B2(n559), .A(n386), .ZN(n270) );
  OAI22_X1 U664 ( .A1(n578), .A2(n470), .B1(n398), .B2(n464), .ZN(n284) );
  INV_X1 U665 ( .A(n270), .ZN(n311) );
  NAND2_X1 U666 ( .A1(n195), .A2(n204), .ZN(n73) );
  OAI22_X1 U667 ( .A1(n361), .A2(n566), .B1(n360), .B2(n462), .ZN(n154) );
  OAI22_X1 U668 ( .A1(n566), .A2(n363), .B1(n462), .B2(n362), .ZN(n160) );
  INV_X1 U669 ( .A(n128), .ZN(n126) );
  INV_X1 U670 ( .A(n131), .ZN(n129) );
  XNOR2_X1 U671 ( .A(a[4]), .B(a[3]), .ZN(n489) );
  OAI22_X1 U672 ( .A1(n421), .A2(n584), .B1(n420), .B2(n466), .ZN(n344) );
  OAI22_X1 U673 ( .A1(n400), .A2(n465), .B1(n483), .B2(n401), .ZN(n325) );
  NAND2_X1 U674 ( .A1(n359), .A2(n287), .ZN(n131) );
  OAI22_X1 U675 ( .A1(n435), .A2(n467), .B1(n485), .B2(n436), .ZN(n359) );
  NAND2_X1 U676 ( .A1(n358), .A2(n347), .ZN(n128) );
  OAI22_X1 U677 ( .A1(n434), .A2(n467), .B1(n435), .B2(n485), .ZN(n358) );
  INV_X1 U678 ( .A(n122), .ZN(n120) );
  NAND2_X1 U679 ( .A1(n139), .A2(n65), .ZN(n10) );
  NOR2_X1 U680 ( .A1(n179), .A2(n186), .ZN(n64) );
  XOR2_X1 U681 ( .A(a[3]), .B(a[2]), .Z(n454) );
  AOI21_X1 U682 ( .B1(n574), .B2(n98), .A(n579), .ZN(n91) );
  NAND2_X1 U683 ( .A1(n574), .A2(n594), .ZN(n90) );
  INV_X1 U684 ( .A(n466), .ZN(n277) );
  NAND2_X1 U685 ( .A1(n179), .A2(n186), .ZN(n65) );
  INV_X1 U686 ( .A(n116), .ZN(n150) );
  NOR2_X1 U687 ( .A1(n261), .A2(n262), .ZN(n116) );
  OAI21_X1 U688 ( .B1(n43), .B2(n39), .A(n40), .ZN(n38) );
  AOI21_X1 U689 ( .B1(n52), .B2(n544), .A(n45), .ZN(n43) );
  INV_X1 U690 ( .A(n586), .ZN(n140) );
  NAND2_X1 U691 ( .A1(n574), .A2(n95), .ZN(n16) );
  OAI22_X1 U692 ( .A1(n406), .A2(n572), .B1(n573), .B2(n407), .ZN(n330) );
  NAND2_X1 U693 ( .A1(n257), .A2(n260), .ZN(n114) );
  OAI22_X1 U694 ( .A1(n485), .A2(n430), .B1(n429), .B2(n467), .ZN(n353) );
  NAND2_X1 U695 ( .A1(n187), .A2(n194), .ZN(n68) );
  XNOR2_X1 U696 ( .A(n444), .B(n602), .ZN(n379) );
  OAI22_X1 U697 ( .A1(n485), .A2(n429), .B1(n428), .B2(n467), .ZN(n352) );
  BUF_X2 U698 ( .A(b[5]), .Z(n444) );
  XNOR2_X1 U699 ( .A(n442), .B(n604), .ZN(n403) );
  INV_X1 U700 ( .A(n56), .ZN(n138) );
  NAND2_X1 U701 ( .A1(n138), .A2(n57), .ZN(n9) );
  NAND2_X1 U702 ( .A1(n51), .A2(n544), .ZN(n42) );
  INV_X1 U703 ( .A(n51), .ZN(n49) );
  OAI22_X1 U704 ( .A1(n403), .A2(n483), .B1(n402), .B2(n465), .ZN(n326) );
  XOR2_X1 U705 ( .A(a[1]), .B(a[0]), .Z(n455) );
  OAI21_X1 U706 ( .B1(n68), .B2(n591), .A(n65), .ZN(n63) );
  OAI22_X1 U707 ( .A1(n584), .A2(n417), .B1(n466), .B2(n416), .ZN(n340) );
  INV_X1 U708 ( .A(n108), .ZN(n148) );
  INV_X1 U709 ( .A(n585), .ZN(n141) );
  OAI22_X1 U710 ( .A1(n419), .A2(n584), .B1(n418), .B2(n466), .ZN(n342) );
  OAI22_X1 U711 ( .A1(n418), .A2(n584), .B1(n417), .B2(n466), .ZN(n341) );
  NAND2_X1 U712 ( .A1(n173), .A2(n178), .ZN(n57) );
  OAI22_X1 U713 ( .A1(n565), .A2(n378), .B1(n377), .B2(n463), .ZN(n303) );
  XNOR2_X1 U714 ( .A(n603), .B(n442), .ZN(n377) );
  XNOR2_X1 U715 ( .A(n443), .B(n603), .ZN(n378) );
  OAI21_X1 U716 ( .B1(n83), .B2(n87), .A(n84), .ZN(n82) );
  NOR2_X1 U717 ( .A1(n592), .A2(n86), .ZN(n81) );
  NAND2_X1 U718 ( .A1(n143), .A2(n84), .ZN(n14) );
  NOR2_X1 U719 ( .A1(n215), .A2(n224), .ZN(n83) );
  AOI21_X1 U720 ( .B1(n71), .B2(n62), .A(n63), .ZN(n61) );
  NOR2_X1 U721 ( .A1(n67), .A2(n64), .ZN(n62) );
  NAND2_X1 U722 ( .A1(n215), .A2(n224), .ZN(n84) );
  INV_X1 U723 ( .A(n463), .ZN(n268) );
  NAND2_X1 U724 ( .A1(n70), .A2(n62), .ZN(n60) );
  OAI22_X1 U725 ( .A1(n426), .A2(n467), .B1(n485), .B2(n427), .ZN(n350) );
  OAI22_X1 U726 ( .A1(n426), .A2(n485), .B1(n425), .B2(n467), .ZN(n349) );
  INV_X1 U727 ( .A(n276), .ZN(n335) );
  AOI21_X1 U728 ( .B1(n584), .B2(n466), .A(n412), .ZN(n276) );
  OAI22_X1 U729 ( .A1(n393), .A2(n464), .B1(n578), .B2(n394), .ZN(n318) );
  AND2_X1 U730 ( .A1(n567), .A2(n274), .ZN(n334) );
  OR2_X1 U731 ( .A1(n567), .A2(n269), .ZN(n385) );
  AND2_X1 U732 ( .A1(n567), .A2(n271), .ZN(n322) );
  OR2_X1 U733 ( .A1(n1), .A2(n278), .ZN(n424) );
  AND2_X1 U734 ( .A1(n567), .A2(n268), .ZN(n310) );
  OR2_X1 U735 ( .A1(n1), .A2(n473), .ZN(n437) );
  OR2_X1 U736 ( .A1(n1), .A2(n275), .ZN(n411) );
  XNOR2_X1 U737 ( .A(n1), .B(n603), .ZN(n384) );
  OR2_X1 U738 ( .A1(n1), .A2(n470), .ZN(n398) );
  OR2_X1 U739 ( .A1(n1), .A2(n468), .ZN(n372) );
  OAI22_X1 U740 ( .A1(n565), .A2(n383), .B1(n382), .B2(n463), .ZN(n308) );
  OAI22_X1 U741 ( .A1(n481), .A2(n382), .B1(n381), .B2(n463), .ZN(n307) );
  XNOR2_X1 U742 ( .A(n576), .B(n603), .ZN(n382) );
  INV_X1 U743 ( .A(n486), .ZN(n265) );
  OAI22_X1 U744 ( .A1(n369), .A2(n462), .B1(n370), .B2(n480), .ZN(n295) );
  OAI22_X1 U745 ( .A1(n369), .A2(n480), .B1(n462), .B2(n368), .ZN(n294) );
  OAI22_X1 U746 ( .A1(n367), .A2(n462), .B1(n480), .B2(n368), .ZN(n293) );
  OAI22_X1 U747 ( .A1(n367), .A2(n566), .B1(n366), .B2(n462), .ZN(n292) );
  OAI22_X1 U748 ( .A1(n366), .A2(n566), .B1(n462), .B2(n365), .ZN(n291) );
  OAI22_X1 U749 ( .A1(n566), .A2(n364), .B1(n462), .B2(n363), .ZN(n290) );
  OAI22_X1 U750 ( .A1(n361), .A2(n462), .B1(n566), .B2(n362), .ZN(n289) );
  AOI21_X1 U751 ( .B1(n566), .B2(n462), .A(n360), .ZN(n264) );
  OAI22_X1 U752 ( .A1(n480), .A2(n468), .B1(n372), .B2(n462), .ZN(n282) );
  AND2_X1 U753 ( .A1(n1), .A2(n265), .ZN(n297) );
  INV_X1 U754 ( .A(n160), .ZN(n161) );
  NAND2_X1 U755 ( .A1(n288), .A2(n154), .ZN(n27) );
  INV_X1 U756 ( .A(n154), .ZN(n155) );
  INV_X1 U757 ( .A(n264), .ZN(n288) );
  XNOR2_X1 U758 ( .A(a[7]), .B(a[8]), .ZN(n487) );
  OR2_X1 U759 ( .A1(n326), .A2(n316), .ZN(n212) );
  XNOR2_X1 U760 ( .A(n316), .B(n326), .ZN(n213) );
  OAI22_X1 U761 ( .A1(n370), .A2(n462), .B1(n480), .B2(n371), .ZN(n296) );
  INV_X1 U762 ( .A(n605), .ZN(n275) );
  XNOR2_X1 U763 ( .A(n439), .B(n605), .ZN(n400) );
  XNOR2_X1 U764 ( .A(n446), .B(n605), .ZN(n407) );
  XNOR2_X1 U765 ( .A(n441), .B(n604), .ZN(n402) );
  NOR2_X1 U766 ( .A1(n77), .A2(n72), .ZN(n70) );
  INV_X1 U767 ( .A(n77), .ZN(n75) );
  NAND2_X1 U768 ( .A1(n75), .A2(n583), .ZN(n13) );
  OAI21_X1 U769 ( .B1(n582), .B2(n78), .A(n73), .ZN(n71) );
  INV_X1 U770 ( .A(n583), .ZN(n76) );
  NOR2_X1 U771 ( .A1(n205), .A2(n214), .ZN(n77) );
  OAI22_X1 U772 ( .A1(n393), .A2(n458), .B1(n392), .B2(n464), .ZN(n317) );
  OAI22_X1 U773 ( .A1(n392), .A2(n458), .B1(n391), .B2(n464), .ZN(n316) );
  NAND2_X1 U774 ( .A1(n454), .A2(n490), .ZN(n484) );
  XNOR2_X1 U775 ( .A(a[1]), .B(a[2]), .ZN(n490) );
  XNOR2_X1 U776 ( .A(n567), .B(n571), .ZN(n423) );
  XNOR2_X1 U777 ( .A(n448), .B(n561), .ZN(n422) );
  INV_X1 U778 ( .A(n478), .ZN(n278) );
  XNOR2_X1 U779 ( .A(n478), .B(n447), .ZN(n421) );
  XNOR2_X1 U780 ( .A(n561), .B(n590), .ZN(n419) );
  XNOR2_X1 U781 ( .A(n478), .B(n446), .ZN(n420) );
  XNOR2_X1 U782 ( .A(n478), .B(n444), .ZN(n418) );
  XNOR2_X1 U783 ( .A(n478), .B(n443), .ZN(n417) );
  XNOR2_X1 U784 ( .A(n478), .B(n439), .ZN(n413) );
  XNOR2_X1 U785 ( .A(n478), .B(n442), .ZN(n416) );
  XNOR2_X1 U786 ( .A(n552), .B(n478), .ZN(n412) );
  OAI22_X1 U787 ( .A1(n460), .A2(n416), .B1(n466), .B2(n415), .ZN(n339) );
  XOR2_X1 U788 ( .A(a[5]), .B(a[4]), .Z(n453) );
  XNOR2_X1 U789 ( .A(n440), .B(n604), .ZN(n401) );
  XNOR2_X1 U790 ( .A(n448), .B(n605), .ZN(n409) );
  XNOR2_X1 U791 ( .A(n1), .B(n604), .ZN(n410) );
  XNOR2_X1 U792 ( .A(n590), .B(n604), .ZN(n406) );
  XNOR2_X1 U793 ( .A(n444), .B(n605), .ZN(n405) );
  AOI21_X1 U794 ( .B1(n595), .B2(n123), .A(n120), .ZN(n118) );
  XNOR2_X1 U795 ( .A(n478), .B(n441), .ZN(n415) );
  NAND2_X1 U796 ( .A1(n144), .A2(n87), .ZN(n15) );
  INV_X1 U797 ( .A(n86), .ZN(n144) );
  NAND2_X1 U798 ( .A1(n205), .A2(n214), .ZN(n78) );
  NAND2_X1 U799 ( .A1(n225), .A2(n232), .ZN(n87) );
  XNOR2_X1 U800 ( .A(n553), .B(n605), .ZN(n399) );
  XNOR2_X1 U801 ( .A(n576), .B(n605), .ZN(n408) );
  OAI22_X1 U802 ( .A1(n415), .A2(n460), .B1(n414), .B2(n466), .ZN(n338) );
  OAI22_X1 U803 ( .A1(n413), .A2(n466), .B1(n584), .B2(n414), .ZN(n337) );
  XNOR2_X1 U804 ( .A(n478), .B(n440), .ZN(n414) );
  OAI21_X1 U805 ( .B1(n116), .B2(n118), .A(n117), .ZN(n115) );
  OAI21_X1 U806 ( .B1(n36), .B2(n34), .A(n35), .ZN(n33) );
  INV_X1 U807 ( .A(n170), .ZN(n171) );
  OAI22_X1 U808 ( .A1(n566), .A2(n365), .B1(n462), .B2(n364), .ZN(n170) );
  XNOR2_X1 U809 ( .A(a[9]), .B(a[10]), .ZN(n486) );
  INV_X1 U810 ( .A(a[0]), .ZN(n491) );
  XNOR2_X1 U811 ( .A(n590), .B(n479), .ZN(n432) );
  INV_X1 U812 ( .A(n479), .ZN(n473) );
  XNOR2_X1 U813 ( .A(n444), .B(n479), .ZN(n431) );
  XNOR2_X1 U814 ( .A(n479), .B(n448), .ZN(n435) );
  XNOR2_X1 U815 ( .A(n479), .B(n443), .ZN(n430) );
  XNOR2_X1 U816 ( .A(n1), .B(n479), .ZN(n436) );
  XNOR2_X1 U817 ( .A(n439), .B(n479), .ZN(n426) );
  XNOR2_X1 U818 ( .A(n479), .B(n441), .ZN(n428) );
  XNOR2_X1 U819 ( .A(n479), .B(n442), .ZN(n429) );
  XNOR2_X1 U820 ( .A(n479), .B(n440), .ZN(n427) );
  XNOR2_X1 U821 ( .A(n576), .B(n479), .ZN(n434) );
  XNOR2_X1 U822 ( .A(n479), .B(n446), .ZN(n433) );
  XNOR2_X1 U823 ( .A(n438), .B(n479), .ZN(n425) );
  INV_X1 U824 ( .A(n184), .ZN(n185) );
  OAI22_X1 U825 ( .A1(n578), .A2(n389), .B1(n388), .B2(n464), .ZN(n184) );
  XNOR2_X1 U826 ( .A(n439), .B(n564), .ZN(n361) );
  XNOR2_X1 U827 ( .A(n553), .B(n564), .ZN(n360) );
  XNOR2_X1 U828 ( .A(n441), .B(n564), .ZN(n363) );
  XNOR2_X1 U829 ( .A(n564), .B(n440), .ZN(n362) );
  INV_X1 U830 ( .A(n564), .ZN(n468) );
  XNOR2_X1 U831 ( .A(n444), .B(n564), .ZN(n366) );
  XNOR2_X1 U832 ( .A(n590), .B(n564), .ZN(n367) );
  XNOR2_X1 U833 ( .A(n447), .B(n564), .ZN(n369) );
  XNOR2_X1 U834 ( .A(n448), .B(n564), .ZN(n370) );
  XNOR2_X1 U835 ( .A(n1), .B(n564), .ZN(n371) );
  XNOR2_X1 U836 ( .A(n446), .B(n564), .ZN(n368) );
  XNOR2_X1 U837 ( .A(n564), .B(n443), .ZN(n365) );
  XNOR2_X1 U838 ( .A(n442), .B(n564), .ZN(n364) );
  XNOR2_X1 U839 ( .A(a[5]), .B(a[6]), .ZN(n488) );
  AOI21_X1 U840 ( .B1(n107), .B2(n597), .A(n104), .ZN(n102) );
  OAI21_X1 U841 ( .B1(n108), .B2(n110), .A(n109), .ZN(n107) );
  OAI22_X1 U842 ( .A1(n434), .A2(n485), .B1(n433), .B2(n467), .ZN(n357) );
  XNOR2_X1 U843 ( .A(n439), .B(n560), .ZN(n387) );
  XNOR2_X1 U844 ( .A(n438), .B(n560), .ZN(n386) );
  XNOR2_X1 U845 ( .A(n1), .B(n476), .ZN(n397) );
  INV_X1 U846 ( .A(n476), .ZN(n470) );
  XNOR2_X1 U847 ( .A(n448), .B(n476), .ZN(n396) );
  XNOR2_X1 U848 ( .A(n590), .B(n476), .ZN(n393) );
  XNOR2_X1 U849 ( .A(n476), .B(n442), .ZN(n390) );
  XNOR2_X1 U850 ( .A(n576), .B(n476), .ZN(n395) );
  XNOR2_X1 U851 ( .A(n444), .B(n476), .ZN(n392) );
  XNOR2_X1 U852 ( .A(n446), .B(n476), .ZN(n394) );
  XNOR2_X1 U853 ( .A(n476), .B(n443), .ZN(n391) );
  XNOR2_X1 U854 ( .A(n476), .B(n441), .ZN(n389) );
  XNOR2_X1 U855 ( .A(n476), .B(n440), .ZN(n388) );
  NAND2_X1 U856 ( .A1(n452), .A2(n488), .ZN(n482) );
  XOR2_X1 U857 ( .A(a[6]), .B(a[7]), .Z(n452) );
  INV_X1 U858 ( .A(n124), .ZN(n123) );
  AOI21_X1 U859 ( .B1(n596), .B2(n129), .A(n126), .ZN(n124) );
  INV_X1 U860 ( .A(n52), .ZN(n50) );
  OAI21_X1 U861 ( .B1(n57), .B2(n53), .A(n54), .ZN(n52) );
  INV_X1 U862 ( .A(n202), .ZN(n203) );
  OAI22_X1 U863 ( .A1(n483), .A2(n402), .B1(n401), .B2(n465), .ZN(n202) );
  OAI21_X1 U864 ( .B1(n90), .B2(n102), .A(n91), .ZN(n89) );
  OAI21_X1 U865 ( .B1(n589), .B2(n60), .A(n61), .ZN(n59) );
  AOI21_X1 U866 ( .B1(n89), .B2(n81), .A(n82), .ZN(n80) );
  AND2_X1 U867 ( .A1(n567), .A2(a[0]), .ZN(product[0]) );
  XNOR2_X1 U868 ( .A(n23), .B(n129), .ZN(product[2]) );
  NAND2_X1 U869 ( .A1(n596), .A2(n128), .ZN(n23) );
  XOR2_X1 U870 ( .A(n21), .B(n118), .Z(product[4]) );
  NAND2_X1 U871 ( .A1(n150), .A2(n117), .ZN(n21) );
  XNOR2_X1 U872 ( .A(n22), .B(n123), .ZN(product[3]) );
  NAND2_X1 U873 ( .A1(n595), .A2(n122), .ZN(n22) );
  XNOR2_X1 U874 ( .A(n20), .B(n569), .ZN(product[5]) );
  NAND2_X1 U875 ( .A1(n598), .A2(n114), .ZN(n20) );
  XOR2_X1 U876 ( .A(n19), .B(n110), .Z(product[6]) );
  NAND2_X1 U877 ( .A1(n148), .A2(n109), .ZN(n19) );
  XNOR2_X1 U878 ( .A(n562), .B(n18), .ZN(product[7]) );
  NAND2_X1 U879 ( .A1(n597), .A2(n106), .ZN(n18) );
  INV_X1 U880 ( .A(n568), .ZN(n101) );
  XOR2_X1 U881 ( .A(n96), .B(n16), .Z(product[9]) );
  AOI21_X1 U882 ( .B1(n101), .B2(n594), .A(n98), .ZN(n96) );
  XOR2_X1 U883 ( .A(n15), .B(n88), .Z(product[10]) );
  INV_X1 U884 ( .A(n89), .ZN(n88) );
  XNOR2_X1 U885 ( .A(n79), .B(n13), .ZN(product[12]) );
  INV_X1 U886 ( .A(n80), .ZN(n79) );
  AOI21_X1 U887 ( .B1(n588), .B2(n37), .A(n38), .ZN(n36) );
  XOR2_X1 U888 ( .A(n58), .B(n9), .Z(product[16]) );
  INV_X1 U889 ( .A(n59), .ZN(n58) );
  AOI21_X1 U890 ( .B1(n79), .B2(n581), .A(n587), .ZN(n69) );
  XOR2_X1 U891 ( .A(n74), .B(n12), .Z(product[13]) );
  AOI21_X1 U892 ( .B1(n79), .B2(n75), .A(n76), .ZN(n74) );
  XNOR2_X1 U893 ( .A(n48), .B(n7), .ZN(product[18]) );
  OAI21_X1 U894 ( .B1(n58), .B2(n49), .A(n50), .ZN(n48) );
  XNOR2_X1 U895 ( .A(n33), .B(n4), .ZN(product[21]) );
  XNOR2_X1 U896 ( .A(n41), .B(n6), .ZN(product[19]) );
  OAI21_X1 U897 ( .B1(n42), .B2(n58), .A(n43), .ZN(n41) );
  XNOR2_X1 U898 ( .A(n55), .B(n8), .ZN(product[17]) );
  OAI21_X1 U899 ( .B1(n56), .B2(n58), .A(n57), .ZN(n55) );
  XNOR2_X1 U900 ( .A(n66), .B(n10), .ZN(product[15]) );
  OAI21_X1 U901 ( .B1(n69), .B2(n586), .A(n547), .ZN(n66) );
  XOR2_X1 U902 ( .A(n28), .B(n3), .Z(product[22]) );
  AOI21_X1 U903 ( .B1(n33), .B2(n546), .A(n30), .ZN(n28) );
  INV_X1 U904 ( .A(n25), .ZN(product[23]) );
  OAI21_X1 U905 ( .B1(n28), .B2(n26), .A(n27), .ZN(n25) );
endmodule


module datapath_DW_mult_tc_22 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n1, n3, n4, n5, n9, n10, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n25, n26, n27, n28, n29, n30, n31, n32, n34, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n57, n59, n60, n61, n62, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n112, n114,
         n115, n117, n119, n120, n121, n123, n125, n126, n127, n128, n129,
         n131, n133, n134, n135, n136, n137, n138, n139, n140, n141, n143,
         n145, n146, n148, n149, n150, n152, n153, n157, n158, n160, n161,
         n165, n167, n168, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n284, n285, n287, n288, n290, n291,
         n293, n294, n296, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n463, n464, n465, n467, n468, n469, n470, n471, n476, n477,
         n479, n480, n481, n482, n483, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n560, n561, n562, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615;

  FA_X1 U194 ( .A(n306), .B(n177), .CI(n315), .CO(n173), .S(n174) );
  FA_X1 U195 ( .A(n316), .B(n178), .CI(n181), .CO(n175), .S(n176) );
  FA_X1 U197 ( .A(n185), .B(n328), .CI(n182), .CO(n179), .S(n180) );
  FA_X1 U198 ( .A(n307), .B(n187), .CI(n317), .CO(n181), .S(n182) );
  FA_X1 U199 ( .A(n186), .B(n193), .CI(n191), .CO(n183), .S(n184) );
  FA_X1 U200 ( .A(n188), .B(n318), .CI(n329), .CO(n185), .S(n186) );
  FA_X1 U202 ( .A(n197), .B(n194), .CI(n192), .CO(n189), .S(n190) );
  FA_X1 U203 ( .A(n339), .B(n308), .CI(n199), .CO(n191), .S(n192) );
  FA_X1 U204 ( .A(n319), .B(n201), .CI(n330), .CO(n193), .S(n194) );
  FA_X1 U205 ( .A(n205), .B(n200), .CI(n198), .CO(n195), .S(n196) );
  FA_X1 U206 ( .A(n209), .B(n202), .CI(n207), .CO(n197), .S(n198) );
  FA_X1 U207 ( .A(n340), .B(n320), .CI(n309), .CO(n199), .S(n200) );
  FA_X1 U209 ( .A(n213), .B(n208), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U210 ( .A(n215), .B(n217), .CI(n210), .CO(n205), .S(n206) );
  FA_X1 U211 ( .A(n310), .B(n321), .CI(n352), .CO(n207), .S(n208) );
  FA_X1 U212 ( .A(n331), .B(n219), .CI(n341), .CO(n209), .S(n210) );
  FA_X1 U213 ( .A(n223), .B(n216), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U214 ( .A(n218), .B(n227), .CI(n225), .CO(n213), .S(n214) );
  FA_X1 U215 ( .A(n220), .B(n322), .CI(n229), .CO(n215), .S(n216) );
  FA_X1 U216 ( .A(n311), .B(n342), .CI(n353), .CO(n217), .S(n218) );
  FA_X1 U218 ( .A(n233), .B(n226), .CI(n224), .CO(n221), .S(n222) );
  FA_X1 U219 ( .A(n228), .B(n237), .CI(n235), .CO(n223), .S(n224) );
  FA_X1 U220 ( .A(n239), .B(n365), .CI(n230), .CO(n225), .S(n226) );
  FA_X1 U221 ( .A(n354), .B(n312), .CI(n323), .CO(n227), .S(n228) );
  FA_X1 U224 ( .A(n243), .B(n236), .CI(n234), .CO(n231), .S(n232) );
  FA_X1 U225 ( .A(n245), .B(n247), .CI(n238), .CO(n233), .S(n234) );
  FA_X1 U226 ( .A(n333), .B(n324), .CI(n240), .CO(n235), .S(n236) );
  FA_X1 U227 ( .A(n366), .B(n313), .CI(n299), .CO(n237), .S(n238) );
  HA_X1 U228 ( .A(n355), .B(n344), .CO(n239), .S(n240) );
  FA_X1 U230 ( .A(n253), .B(n255), .CI(n248), .CO(n243), .S(n244) );
  FA_X1 U231 ( .A(n367), .B(n334), .CI(n325), .CO(n245), .S(n246) );
  FA_X1 U232 ( .A(n356), .B(n314), .CI(n345), .CO(n247), .S(n248) );
  FA_X1 U234 ( .A(n256), .B(n300), .CI(n261), .CO(n251), .S(n252) );
  FA_X1 U235 ( .A(n346), .B(n335), .CI(n326), .CO(n253), .S(n254) );
  HA_X1 U236 ( .A(n368), .B(n357), .CO(n255), .S(n256) );
  FA_X1 U237 ( .A(n262), .B(n265), .CI(n260), .CO(n257), .S(n258) );
  FA_X1 U238 ( .A(n336), .B(n347), .CI(n267), .CO(n259), .S(n260) );
  FA_X1 U239 ( .A(n369), .B(n327), .CI(n358), .CO(n261), .S(n262) );
  FA_X1 U240 ( .A(n271), .B(n268), .CI(n266), .CO(n263), .S(n264) );
  FA_X1 U241 ( .A(n337), .B(n301), .CI(n359), .CO(n265), .S(n266) );
  HA_X1 U242 ( .A(n348), .B(n370), .CO(n267), .S(n268) );
  FA_X1 U244 ( .A(n371), .B(n338), .CI(n360), .CO(n271), .S(n272) );
  FA_X1 U245 ( .A(n372), .B(n350), .CI(n276), .CO(n273), .S(n274) );
  HA_X1 U246 ( .A(n361), .B(n302), .CO(n275), .S(n276) );
  FA_X1 U247 ( .A(n351), .B(n373), .CI(n362), .CO(n277), .S(n278) );
  HA_X1 U248 ( .A(n374), .B(n303), .CO(n279), .S(n280) );
  CLKBUF_X1 U484 ( .A(b[5]), .Z(n461) );
  BUF_X1 U485 ( .A(b[8]), .Z(n458) );
  INV_X1 U486 ( .A(n562), .ZN(n560) );
  CLKBUF_X3 U487 ( .A(a[11]), .Z(n491) );
  CLKBUF_X2 U488 ( .A(b[7]), .Z(n459) );
  FA_X1 U489 ( .A(n223), .B(n216), .CI(n214), .S(n561) );
  AOI21_X1 U490 ( .B1(n108), .B2(n100), .A(n101), .ZN(n562) );
  BUF_X2 U491 ( .A(b[2]), .Z(n464) );
  CLKBUF_X3 U492 ( .A(a[1]), .Z(n496) );
  CLKBUF_X1 U493 ( .A(n70), .Z(n602) );
  AND2_X1 U494 ( .A1(n608), .A2(n148), .ZN(product[1]) );
  AND3_X1 U495 ( .A1(n583), .A2(n584), .A3(n585), .ZN(product[23]) );
  BUF_X1 U496 ( .A(b[9]), .Z(n457) );
  BUF_X1 U497 ( .A(b[3]), .Z(n463) );
  OAI21_X1 U498 ( .B1(n573), .B2(n97), .A(n92), .ZN(n565) );
  BUF_X2 U499 ( .A(n500), .Z(n566) );
  CLKBUF_X3 U500 ( .A(n506), .Z(n482) );
  BUF_X1 U501 ( .A(b[10]), .Z(n456) );
  XNOR2_X1 U502 ( .A(n252), .B(n567), .ZN(n250) );
  XNOR2_X1 U503 ( .A(n254), .B(n259), .ZN(n567) );
  CLKBUF_X1 U504 ( .A(n601), .Z(n568) );
  CLKBUF_X1 U505 ( .A(n1), .Z(n569) );
  BUF_X1 U506 ( .A(b[0]), .Z(n1) );
  BUF_X2 U507 ( .A(n497), .Z(n570) );
  NAND2_X1 U508 ( .A1(n467), .A2(n503), .ZN(n497) );
  OR2_X2 U509 ( .A1(n571), .A2(a[0]), .ZN(n502) );
  XNOR2_X1 U510 ( .A(a[1]), .B(a[0]), .ZN(n571) );
  CLKBUF_X1 U511 ( .A(n496), .Z(n572) );
  BUF_X2 U512 ( .A(n1), .Z(n612) );
  NAND2_X2 U513 ( .A1(n505), .A2(n469), .ZN(n499) );
  NOR2_X1 U514 ( .A1(n561), .A2(n221), .ZN(n573) );
  BUF_X2 U515 ( .A(n501), .Z(n574) );
  NOR2_X1 U516 ( .A1(n212), .A2(n221), .ZN(n91) );
  NOR2_X2 U517 ( .A1(n278), .A2(n279), .ZN(n135) );
  XOR2_X1 U518 ( .A(n251), .B(n246), .Z(n575) );
  XOR2_X1 U519 ( .A(n244), .B(n575), .Z(n242) );
  NAND2_X1 U520 ( .A1(n244), .A2(n251), .ZN(n576) );
  NAND2_X1 U521 ( .A1(n244), .A2(n246), .ZN(n577) );
  NAND2_X1 U522 ( .A1(n251), .A2(n246), .ZN(n578) );
  NAND3_X1 U523 ( .A1(n576), .A2(n577), .A3(n578), .ZN(n241) );
  CLKBUF_X3 U524 ( .A(a[3]), .Z(n495) );
  OAI21_X1 U525 ( .B1(n135), .B2(n137), .A(n136), .ZN(n579) );
  XNOR2_X1 U526 ( .A(n51), .B(n580), .ZN(product[18]) );
  AND2_X1 U527 ( .A1(n153), .A2(n50), .ZN(n580) );
  AOI21_X1 U528 ( .B1(n610), .B2(n579), .A(n131), .ZN(n581) );
  BUF_X1 U529 ( .A(b[6]), .Z(n460) );
  BUF_X2 U530 ( .A(b[1]), .Z(n465) );
  CLKBUF_X3 U531 ( .A(n503), .Z(n479) );
  XOR2_X1 U532 ( .A(n305), .B(n171), .Z(n582) );
  XOR2_X1 U533 ( .A(n149), .B(n582), .Z(product[22]) );
  NAND2_X1 U534 ( .A1(n149), .A2(n305), .ZN(n583) );
  NAND2_X1 U535 ( .A1(n149), .A2(n171), .ZN(n584) );
  NAND2_X1 U536 ( .A1(n305), .A2(n171), .ZN(n585) );
  CLKBUF_X3 U537 ( .A(a[5]), .Z(n494) );
  OR2_X1 U538 ( .A1(n196), .A2(n203), .ZN(n586) );
  INV_X1 U539 ( .A(n95), .ZN(n587) );
  XNOR2_X1 U540 ( .A(n69), .B(n588), .ZN(product[16]) );
  AND2_X1 U541 ( .A1(n61), .A2(n68), .ZN(n588) );
  XNOR2_X1 U542 ( .A(n60), .B(n589), .ZN(product[17]) );
  AND2_X1 U543 ( .A1(n604), .A2(n59), .ZN(n589) );
  BUF_X2 U544 ( .A(b[11]), .Z(n455) );
  XNOR2_X1 U545 ( .A(n93), .B(n590), .ZN(product[13]) );
  AND2_X1 U546 ( .A1(n158), .A2(n92), .ZN(n590) );
  XOR2_X1 U547 ( .A(n275), .B(n349), .Z(n591) );
  XOR2_X1 U548 ( .A(n272), .B(n591), .Z(n270) );
  NAND2_X1 U549 ( .A1(n272), .A2(n275), .ZN(n592) );
  NAND2_X1 U550 ( .A1(n272), .A2(n349), .ZN(n593) );
  NAND2_X1 U551 ( .A1(n275), .A2(n349), .ZN(n594) );
  NAND3_X1 U552 ( .A1(n592), .A2(n593), .A3(n594), .ZN(n269) );
  BUF_X2 U553 ( .A(n1), .Z(n611) );
  NAND2_X1 U554 ( .A1(n252), .A2(n254), .ZN(n595) );
  NAND2_X1 U555 ( .A1(n252), .A2(n259), .ZN(n596) );
  NAND2_X1 U556 ( .A1(n254), .A2(n259), .ZN(n597) );
  NAND3_X1 U557 ( .A1(n595), .A2(n596), .A3(n597), .ZN(n249) );
  OR2_X1 U558 ( .A1(n502), .A2(n446), .ZN(n598) );
  OR2_X1 U559 ( .A1(n445), .A2(n508), .ZN(n599) );
  NAND2_X1 U560 ( .A1(n598), .A2(n599), .ZN(n369) );
  NOR2_X1 U561 ( .A1(n232), .A2(n241), .ZN(n600) );
  XNOR2_X1 U562 ( .A(n569), .B(n491), .ZN(n388) );
  NAND2_X1 U563 ( .A1(n468), .A2(n504), .ZN(n601) );
  XOR2_X1 U564 ( .A(n107), .B(n14), .Z(product[10]) );
  XOR2_X1 U565 ( .A(n115), .B(n15), .Z(product[9]) );
  XNOR2_X1 U566 ( .A(n104), .B(n13), .ZN(product[11]) );
  OR2_X1 U567 ( .A1(n258), .A2(n263), .ZN(n603) );
  OR2_X1 U568 ( .A1(n189), .A2(n184), .ZN(n604) );
  OR2_X1 U569 ( .A1(n250), .A2(n257), .ZN(n605) );
  OR2_X1 U570 ( .A1(n175), .A2(n174), .ZN(n606) );
  OR2_X1 U571 ( .A1(n375), .A2(n364), .ZN(n607) );
  OR2_X1 U572 ( .A1(n376), .A2(n304), .ZN(n608) );
  OR2_X1 U573 ( .A1(n264), .A2(n269), .ZN(n609) );
  OR2_X1 U574 ( .A1(n274), .A2(n277), .ZN(n610) );
  BUF_X2 U575 ( .A(n504), .Z(n480) );
  BUF_X2 U576 ( .A(n507), .Z(n483) );
  BUF_X1 U577 ( .A(n492), .Z(n613) );
  BUF_X1 U578 ( .A(n492), .Z(n615) );
  BUF_X1 U579 ( .A(n492), .Z(n614) );
  BUF_X2 U580 ( .A(a[7]), .Z(n493) );
  BUF_X1 U581 ( .A(a[9]), .Z(n492) );
  INV_X1 U582 ( .A(n28), .ZN(n150) );
  NAND2_X1 U583 ( .A1(n150), .A2(n29), .ZN(n3) );
  NOR2_X1 U584 ( .A1(n173), .A2(n172), .ZN(n28) );
  NAND2_X1 U585 ( .A1(n173), .A2(n172), .ZN(n29) );
  NOR2_X1 U586 ( .A1(n190), .A2(n195), .ZN(n67) );
  NAND2_X1 U587 ( .A1(n606), .A2(n36), .ZN(n4) );
  INV_X1 U588 ( .A(n36), .ZN(n34) );
  NAND2_X1 U589 ( .A1(n175), .A2(n174), .ZN(n36) );
  INV_X1 U590 ( .A(n68), .ZN(n62) );
  OAI21_X1 U591 ( .B1(n68), .B2(n54), .A(n59), .ZN(n53) );
  INV_X1 U592 ( .A(n67), .ZN(n61) );
  NOR2_X1 U593 ( .A1(n67), .A2(n54), .ZN(n52) );
  NOR2_X1 U594 ( .A1(n176), .A2(n179), .ZN(n46) );
  INV_X1 U595 ( .A(n157), .ZN(n80) );
  AOI21_X1 U596 ( .B1(n120), .B2(n603), .A(n117), .ZN(n115) );
  INV_X1 U597 ( .A(n87), .ZN(n85) );
  NOR2_X1 U598 ( .A1(n87), .A2(n80), .ZN(n78) );
  INV_X1 U599 ( .A(n88), .ZN(n86) );
  XOR2_X1 U600 ( .A(a[9]), .B(a[8]), .Z(n468) );
  NAND2_X1 U601 ( .A1(n278), .A2(n279), .ZN(n136) );
  OAI21_X1 U602 ( .B1(n71), .B2(n99), .A(n72), .ZN(n70) );
  BUF_X2 U603 ( .A(n505), .Z(n481) );
  NAND2_X1 U604 ( .A1(n270), .A2(n273), .ZN(n128) );
  OAI22_X1 U605 ( .A1(n499), .A2(n406), .B1(n405), .B2(n481), .ZN(n201) );
  NAND2_X1 U606 ( .A1(n190), .A2(n195), .ZN(n68) );
  OAI22_X1 U607 ( .A1(n378), .A2(n570), .B1(n377), .B2(n479), .ZN(n171) );
  BUF_X2 U608 ( .A(n500), .Z(n476) );
  NAND2_X1 U609 ( .A1(n603), .A2(n119), .ZN(n16) );
  INV_X1 U610 ( .A(n46), .ZN(n152) );
  NAND2_X1 U611 ( .A1(n152), .A2(n47), .ZN(n5) );
  XNOR2_X1 U612 ( .A(n463), .B(n615), .ZN(n398) );
  OAI22_X1 U613 ( .A1(n566), .A2(n427), .B1(n426), .B2(n482), .ZN(n350) );
  OAI22_X1 U614 ( .A1(n423), .A2(n482), .B1(n566), .B2(n424), .ZN(n347) );
  INV_X1 U615 ( .A(n290), .ZN(n339) );
  INV_X1 U616 ( .A(n604), .ZN(n54) );
  OAI22_X1 U617 ( .A1(n417), .A2(n482), .B1(n566), .B2(n418), .ZN(n341) );
  INV_X1 U618 ( .A(n40), .ZN(n38) );
  NOR2_X1 U619 ( .A1(n67), .A2(n42), .ZN(n40) );
  OAI22_X1 U620 ( .A1(n476), .A2(n419), .B1(n418), .B2(n482), .ZN(n342) );
  NAND2_X1 U621 ( .A1(n586), .A2(n76), .ZN(n9) );
  BUF_X2 U622 ( .A(n501), .Z(n477) );
  NAND2_X1 U623 ( .A1(n280), .A2(n363), .ZN(n140) );
  XOR2_X1 U624 ( .A(a[11]), .B(a[10]), .Z(n467) );
  OAI22_X1 U625 ( .A1(n502), .A2(n453), .B1(n452), .B2(n508), .ZN(n376) );
  OAI22_X1 U626 ( .A1(n449), .A2(n508), .B1(n502), .B2(n450), .ZN(n373) );
  AOI21_X1 U627 ( .B1(n502), .B2(n508), .A(n442), .ZN(n296) );
  OAI22_X1 U628 ( .A1(n451), .A2(n502), .B1(n450), .B2(n508), .ZN(n374) );
  XNOR2_X1 U629 ( .A(b[4]), .B(n613), .ZN(n397) );
  NAND2_X1 U630 ( .A1(n176), .A2(n179), .ZN(n47) );
  NAND2_X1 U631 ( .A1(n183), .A2(n180), .ZN(n50) );
  OAI22_X1 U632 ( .A1(n502), .A2(n445), .B1(n444), .B2(n508), .ZN(n368) );
  OAI22_X1 U633 ( .A1(n477), .A2(n440), .B1(n439), .B2(n483), .ZN(n363) );
  AOI21_X1 U634 ( .B1(n477), .B2(n483), .A(n429), .ZN(n293) );
  OAI22_X1 U635 ( .A1(n436), .A2(n483), .B1(n574), .B2(n437), .ZN(n360) );
  OAI22_X1 U636 ( .A1(n574), .A2(n434), .B1(n433), .B2(n483), .ZN(n357) );
  OAI22_X1 U637 ( .A1(n423), .A2(n566), .B1(n422), .B2(n482), .ZN(n346) );
  OAI22_X1 U638 ( .A1(n422), .A2(n566), .B1(n421), .B2(n482), .ZN(n345) );
  OAI22_X1 U639 ( .A1(n449), .A2(n502), .B1(n448), .B2(n508), .ZN(n372) );
  OAI22_X1 U640 ( .A1(n448), .A2(n502), .B1(n447), .B2(n508), .ZN(n371) );
  XNOR2_X1 U641 ( .A(b[4]), .B(n496), .ZN(n449) );
  XNOR2_X1 U642 ( .A(n496), .B(n460), .ZN(n447) );
  XNOR2_X1 U643 ( .A(n463), .B(n496), .ZN(n450) );
  NOR2_X1 U644 ( .A1(n242), .A2(n249), .ZN(n105) );
  AOI21_X1 U645 ( .B1(n568), .B2(n480), .A(n390), .ZN(n284) );
  INV_X1 U646 ( .A(n125), .ZN(n123) );
  XNOR2_X1 U647 ( .A(a[3]), .B(a[4]), .ZN(n506) );
  INV_X1 U648 ( .A(n482), .ZN(n291) );
  INV_X1 U649 ( .A(n145), .ZN(n143) );
  OAI22_X1 U650 ( .A1(n477), .A2(n433), .B1(n432), .B2(n483), .ZN(n356) );
  NAND2_X1 U651 ( .A1(n258), .A2(n263), .ZN(n119) );
  OAI22_X1 U652 ( .A1(n430), .A2(n483), .B1(n574), .B2(n431), .ZN(n354) );
  OAI22_X1 U653 ( .A1(n399), .A2(n601), .B1(n398), .B2(n480), .ZN(n324) );
  OAI22_X1 U654 ( .A1(n397), .A2(n601), .B1(n396), .B2(n480), .ZN(n322) );
  OAI22_X1 U655 ( .A1(n568), .A2(n394), .B1(n393), .B2(n480), .ZN(n319) );
  OAI22_X1 U656 ( .A1(n568), .A2(n393), .B1(n392), .B2(n480), .ZN(n318) );
  OAI22_X1 U657 ( .A1(n391), .A2(n480), .B1(n568), .B2(n392), .ZN(n317) );
  OAI22_X1 U658 ( .A1(n391), .A2(n568), .B1(n390), .B2(n480), .ZN(n316) );
  OAI22_X1 U659 ( .A1(n601), .A2(n486), .B1(n402), .B2(n480), .ZN(n300) );
  INV_X1 U660 ( .A(n284), .ZN(n315) );
  NAND2_X1 U661 ( .A1(n161), .A2(n106), .ZN(n14) );
  OAI21_X1 U662 ( .B1(n107), .B2(n105), .A(n106), .ZN(n104) );
  NOR2_X1 U663 ( .A1(n204), .A2(n211), .ZN(n82) );
  XNOR2_X1 U664 ( .A(n496), .B(n457), .ZN(n444) );
  XNOR2_X1 U665 ( .A(n613), .B(n457), .ZN(n392) );
  OAI22_X1 U666 ( .A1(n502), .A2(n490), .B1(n454), .B2(n508), .ZN(n304) );
  NAND2_X1 U667 ( .A1(n196), .A2(n203), .ZN(n76) );
  NAND2_X1 U668 ( .A1(n264), .A2(n269), .ZN(n125) );
  INV_X1 U669 ( .A(n82), .ZN(n157) );
  AND2_X1 U670 ( .A1(n612), .A2(n294), .ZN(n364) );
  NOR2_X1 U671 ( .A1(n222), .A2(n231), .ZN(n96) );
  OAI22_X1 U672 ( .A1(n601), .A2(n401), .B1(n400), .B2(n480), .ZN(n326) );
  INV_X1 U673 ( .A(n133), .ZN(n131) );
  XNOR2_X1 U674 ( .A(n496), .B(n458), .ZN(n445) );
  XNOR2_X1 U675 ( .A(n613), .B(n458), .ZN(n393) );
  OAI22_X1 U676 ( .A1(n397), .A2(n480), .B1(n601), .B2(n398), .ZN(n323) );
  INV_X1 U677 ( .A(n600), .ZN(n160) );
  NAND2_X1 U678 ( .A1(n605), .A2(n114), .ZN(n15) );
  NAND2_X1 U679 ( .A1(n242), .A2(n249), .ZN(n106) );
  NOR2_X1 U680 ( .A1(n196), .A2(n203), .ZN(n75) );
  NAND2_X1 U681 ( .A1(n375), .A2(n364), .ZN(n145) );
  OAI22_X1 U682 ( .A1(n502), .A2(n452), .B1(n451), .B2(n508), .ZN(n375) );
  OAI21_X1 U683 ( .B1(n32), .B2(n28), .A(n29), .ZN(n27) );
  AOI21_X1 U684 ( .B1(n41), .B2(n606), .A(n34), .ZN(n32) );
  NAND2_X1 U685 ( .A1(n605), .A2(n603), .ZN(n109) );
  OAI22_X1 U686 ( .A1(n417), .A2(n566), .B1(n416), .B2(n482), .ZN(n340) );
  AOI21_X1 U687 ( .B1(n566), .B2(n482), .A(n416), .ZN(n290) );
  INV_X1 U688 ( .A(n135), .ZN(n167) );
  INV_X1 U689 ( .A(n127), .ZN(n165) );
  NOR2_X1 U690 ( .A1(n270), .A2(n273), .ZN(n127) );
  NOR2_X1 U691 ( .A1(n31), .A2(n28), .ZN(n26) );
  NAND2_X1 U692 ( .A1(n40), .A2(n606), .ZN(n31) );
  NAND2_X1 U693 ( .A1(n274), .A2(n277), .ZN(n133) );
  NAND2_X1 U694 ( .A1(n250), .A2(n257), .ZN(n114) );
  INV_X1 U695 ( .A(n119), .ZN(n117) );
  XNOR2_X1 U696 ( .A(a[7]), .B(a[8]), .ZN(n504) );
  OAI22_X1 U697 ( .A1(n438), .A2(n483), .B1(n439), .B2(n574), .ZN(n362) );
  XNOR2_X1 U698 ( .A(a[1]), .B(a[2]), .ZN(n507) );
  INV_X1 U699 ( .A(n483), .ZN(n294) );
  INV_X1 U700 ( .A(n614), .ZN(n486) );
  OAI22_X1 U701 ( .A1(n438), .A2(n477), .B1(n437), .B2(n483), .ZN(n361) );
  NAND2_X1 U702 ( .A1(n157), .A2(n83), .ZN(n10) );
  OAI21_X1 U703 ( .B1(n88), .B2(n80), .A(n83), .ZN(n79) );
  INV_X1 U704 ( .A(n293), .ZN(n352) );
  OAI22_X1 U705 ( .A1(n396), .A2(n601), .B1(n395), .B2(n480), .ZN(n321) );
  OAI22_X1 U706 ( .A1(n568), .A2(n395), .B1(n394), .B2(n480), .ZN(n320) );
  XNOR2_X1 U707 ( .A(n613), .B(n460), .ZN(n395) );
  INV_X1 U708 ( .A(n573), .ZN(n158) );
  NOR2_X1 U709 ( .A1(n96), .A2(n91), .ZN(n89) );
  OAI21_X1 U710 ( .B1(n91), .B2(n97), .A(n92), .ZN(n90) );
  OAI22_X1 U711 ( .A1(n502), .A2(n447), .B1(n446), .B2(n508), .ZN(n370) );
  INV_X1 U712 ( .A(n41), .ZN(n39) );
  OAI21_X1 U713 ( .B1(n42), .B2(n68), .A(n43), .ZN(n41) );
  NAND2_X1 U714 ( .A1(n561), .A2(n221), .ZN(n92) );
  XNOR2_X1 U715 ( .A(b[4]), .B(n494), .ZN(n423) );
  XNOR2_X1 U716 ( .A(n494), .B(n457), .ZN(n418) );
  XNOR2_X1 U717 ( .A(n494), .B(n458), .ZN(n419) );
  XNOR2_X1 U718 ( .A(n463), .B(n494), .ZN(n424) );
  OAI22_X1 U719 ( .A1(n476), .A2(n420), .B1(n419), .B2(n482), .ZN(n343) );
  INV_X1 U720 ( .A(n296), .ZN(n365) );
  OAI22_X1 U721 ( .A1(n443), .A2(n502), .B1(n442), .B2(n508), .ZN(n366) );
  OAI22_X1 U722 ( .A1(n425), .A2(n482), .B1(n426), .B2(n566), .ZN(n349) );
  OAI22_X1 U723 ( .A1(n425), .A2(n476), .B1(n424), .B2(n482), .ZN(n348) );
  AOI21_X1 U724 ( .B1(n607), .B2(n146), .A(n143), .ZN(n141) );
  AOI21_X1 U725 ( .B1(n605), .B2(n117), .A(n112), .ZN(n110) );
  INV_X1 U726 ( .A(n114), .ZN(n112) );
  OAI22_X1 U727 ( .A1(n436), .A2(n574), .B1(n435), .B2(n483), .ZN(n359) );
  OAI22_X1 U728 ( .A1(n435), .A2(n477), .B1(n434), .B2(n483), .ZN(n358) );
  XNOR2_X1 U729 ( .A(n496), .B(n459), .ZN(n446) );
  XNOR2_X1 U730 ( .A(n494), .B(n459), .ZN(n420) );
  XNOR2_X1 U731 ( .A(n615), .B(n459), .ZN(n394) );
  XNOR2_X1 U732 ( .A(n464), .B(n496), .ZN(n451) );
  XNOR2_X1 U733 ( .A(n464), .B(n494), .ZN(n425) );
  XNOR2_X1 U734 ( .A(n464), .B(n614), .ZN(n399) );
  OAI21_X1 U735 ( .B1(n102), .B2(n106), .A(n103), .ZN(n101) );
  NOR2_X1 U736 ( .A1(n600), .A2(n105), .ZN(n100) );
  NAND2_X1 U737 ( .A1(n160), .A2(n103), .ZN(n13) );
  NOR2_X1 U738 ( .A1(n232), .A2(n241), .ZN(n102) );
  XNOR2_X1 U739 ( .A(n465), .B(n496), .ZN(n452) );
  XNOR2_X1 U740 ( .A(n465), .B(n494), .ZN(n426) );
  XNOR2_X1 U741 ( .A(n465), .B(n614), .ZN(n400) );
  XNOR2_X1 U742 ( .A(n461), .B(n572), .ZN(n448) );
  XNOR2_X1 U743 ( .A(n461), .B(n494), .ZN(n422) );
  XNOR2_X1 U744 ( .A(n461), .B(n615), .ZN(n396) );
  INV_X1 U745 ( .A(n96), .ZN(n94) );
  NAND2_X1 U746 ( .A1(n94), .A2(n587), .ZN(n12) );
  INV_X1 U747 ( .A(n97), .ZN(n95) );
  INV_X1 U748 ( .A(n89), .ZN(n87) );
  INV_X1 U749 ( .A(n565), .ZN(n88) );
  XNOR2_X1 U750 ( .A(n456), .B(n496), .ZN(n443) );
  XNOR2_X1 U751 ( .A(n456), .B(n494), .ZN(n417) );
  XNOR2_X1 U752 ( .A(n456), .B(n615), .ZN(n391) );
  XNOR2_X1 U753 ( .A(n455), .B(n496), .ZN(n442) );
  XNOR2_X1 U754 ( .A(n455), .B(n494), .ZN(n416) );
  XNOR2_X1 U755 ( .A(n455), .B(n613), .ZN(n390) );
  INV_X1 U756 ( .A(n480), .ZN(n285) );
  AND2_X1 U757 ( .A1(n611), .A2(n291), .ZN(n351) );
  XNOR2_X1 U758 ( .A(n611), .B(n494), .ZN(n427) );
  OR2_X1 U759 ( .A1(n611), .A2(n486), .ZN(n402) );
  OR2_X1 U760 ( .A1(n611), .A2(n489), .ZN(n441) );
  XNOR2_X1 U761 ( .A(n612), .B(n572), .ZN(n453) );
  OR2_X1 U762 ( .A1(n611), .A2(n490), .ZN(n454) );
  OR2_X1 U763 ( .A1(n611), .A2(n487), .ZN(n415) );
  AND2_X1 U764 ( .A1(n611), .A2(n285), .ZN(n327) );
  OR2_X1 U765 ( .A1(n611), .A2(n488), .ZN(n428) );
  XNOR2_X1 U766 ( .A(n611), .B(n614), .ZN(n401) );
  OR2_X1 U767 ( .A1(n612), .A2(n485), .ZN(n389) );
  NAND2_X1 U768 ( .A1(n222), .A2(n231), .ZN(n97) );
  INV_X1 U769 ( .A(n49), .ZN(n153) );
  NOR2_X1 U770 ( .A1(n49), .A2(n46), .ZN(n44) );
  NOR2_X1 U771 ( .A1(n183), .A2(n180), .ZN(n49) );
  NAND2_X1 U772 ( .A1(n232), .A2(n241), .ZN(n103) );
  OAI22_X1 U773 ( .A1(n443), .A2(n508), .B1(n502), .B2(n444), .ZN(n367) );
  OAI22_X1 U774 ( .A1(n399), .A2(n480), .B1(n400), .B2(n601), .ZN(n325) );
  INV_X1 U775 ( .A(n59), .ZN(n57) );
  OAI22_X1 U776 ( .A1(n430), .A2(n477), .B1(n429), .B2(n483), .ZN(n353) );
  OAI22_X1 U777 ( .A1(n421), .A2(n476), .B1(n420), .B2(n482), .ZN(n344) );
  XNOR2_X1 U778 ( .A(n494), .B(n460), .ZN(n421) );
  OAI22_X1 U779 ( .A1(n477), .A2(n432), .B1(n431), .B2(n483), .ZN(n355) );
  INV_X1 U780 ( .A(n479), .ZN(n282) );
  OAI22_X1 U781 ( .A1(n387), .A2(n479), .B1(n388), .B2(n497), .ZN(n313) );
  OAI22_X1 U782 ( .A1(n386), .A2(n479), .B1(n387), .B2(n497), .ZN(n312) );
  OAI22_X1 U783 ( .A1(n386), .A2(n497), .B1(n385), .B2(n479), .ZN(n311) );
  OAI22_X1 U784 ( .A1(n384), .A2(n479), .B1(n497), .B2(n385), .ZN(n310) );
  OAI22_X1 U785 ( .A1(n384), .A2(n570), .B1(n383), .B2(n479), .ZN(n309) );
  OAI22_X1 U786 ( .A1(n383), .A2(n570), .B1(n479), .B2(n382), .ZN(n308) );
  OAI22_X1 U787 ( .A1(n570), .A2(n382), .B1(n479), .B2(n381), .ZN(n187) );
  OAI22_X1 U788 ( .A1(n570), .A2(n381), .B1(n479), .B2(n380), .ZN(n307) );
  OAI22_X1 U789 ( .A1(n570), .A2(n380), .B1(n479), .B2(n379), .ZN(n177) );
  OAI22_X1 U790 ( .A1(n378), .A2(n479), .B1(n570), .B2(n379), .ZN(n306) );
  AOI21_X1 U791 ( .B1(n570), .B2(n479), .A(n377), .ZN(n281) );
  OAI22_X1 U792 ( .A1(n389), .A2(n479), .B1(n497), .B2(n485), .ZN(n299) );
  AND2_X1 U793 ( .A1(n612), .A2(n282), .ZN(n314) );
  INV_X1 U794 ( .A(n171), .ZN(n172) );
  INV_X1 U795 ( .A(n281), .ZN(n305) );
  XNOR2_X1 U796 ( .A(n612), .B(n495), .ZN(n440) );
  XNOR2_X1 U797 ( .A(n465), .B(n495), .ZN(n439) );
  XNOR2_X1 U798 ( .A(b[4]), .B(n495), .ZN(n436) );
  XNOR2_X1 U799 ( .A(n464), .B(n495), .ZN(n438) );
  XNOR2_X1 U800 ( .A(n463), .B(n495), .ZN(n437) );
  XNOR2_X1 U801 ( .A(n461), .B(n495), .ZN(n435) );
  XNOR2_X1 U802 ( .A(n495), .B(n460), .ZN(n434) );
  XNOR2_X1 U803 ( .A(n456), .B(n495), .ZN(n430) );
  XNOR2_X1 U804 ( .A(n495), .B(n459), .ZN(n433) );
  XNOR2_X1 U805 ( .A(n455), .B(n495), .ZN(n429) );
  XNOR2_X1 U806 ( .A(n495), .B(n457), .ZN(n431) );
  XNOR2_X1 U807 ( .A(n495), .B(n458), .ZN(n432) );
  NAND2_X1 U808 ( .A1(n470), .A2(n506), .ZN(n500) );
  XOR2_X1 U809 ( .A(a[5]), .B(a[4]), .Z(n470) );
  INV_X1 U810 ( .A(n105), .ZN(n161) );
  NAND2_X1 U811 ( .A1(n471), .A2(n507), .ZN(n501) );
  XOR2_X1 U812 ( .A(a[3]), .B(a[2]), .Z(n471) );
  INV_X1 U813 ( .A(n177), .ZN(n178) );
  OAI22_X1 U814 ( .A1(n574), .A2(n489), .B1(n441), .B2(n483), .ZN(n303) );
  INV_X1 U815 ( .A(n495), .ZN(n489) );
  INV_X1 U816 ( .A(n496), .ZN(n490) );
  INV_X1 U817 ( .A(n139), .ZN(n168) );
  NOR2_X1 U818 ( .A1(n280), .A2(n363), .ZN(n139) );
  OAI22_X1 U819 ( .A1(n476), .A2(n488), .B1(n428), .B2(n482), .ZN(n302) );
  INV_X1 U820 ( .A(n494), .ZN(n488) );
  INV_X1 U821 ( .A(n481), .ZN(n288) );
  AND2_X1 U822 ( .A1(n612), .A2(n288), .ZN(n338) );
  INV_X1 U823 ( .A(n201), .ZN(n202) );
  INV_X1 U824 ( .A(n287), .ZN(n328) );
  OR2_X1 U825 ( .A1(n332), .A2(n343), .ZN(n229) );
  XNOR2_X1 U826 ( .A(n332), .B(n343), .ZN(n230) );
  INV_X1 U827 ( .A(n148), .ZN(n146) );
  NAND2_X1 U828 ( .A1(n376), .A2(n304), .ZN(n148) );
  XNOR2_X1 U829 ( .A(a[5]), .B(a[6]), .ZN(n505) );
  OAI22_X1 U830 ( .A1(n499), .A2(n408), .B1(n407), .B2(n481), .ZN(n219) );
  INV_X1 U831 ( .A(n219), .ZN(n220) );
  OAI21_X1 U832 ( .B1(n139), .B2(n141), .A(n140), .ZN(n138) );
  NAND2_X1 U833 ( .A1(n89), .A2(n73), .ZN(n71) );
  NOR2_X1 U834 ( .A1(n82), .A2(n75), .ZN(n73) );
  OAI22_X1 U835 ( .A1(n412), .A2(n499), .B1(n411), .B2(n481), .ZN(n335) );
  OAI22_X1 U836 ( .A1(n499), .A2(n407), .B1(n406), .B2(n481), .ZN(n331) );
  OAI22_X1 U837 ( .A1(n410), .A2(n499), .B1(n409), .B2(n481), .ZN(n333) );
  OAI22_X1 U838 ( .A1(n404), .A2(n481), .B1(n499), .B2(n405), .ZN(n330) );
  OAI22_X1 U839 ( .A1(n499), .A2(n487), .B1(n415), .B2(n481), .ZN(n301) );
  AOI21_X1 U840 ( .B1(n499), .B2(n481), .A(n403), .ZN(n287) );
  OAI22_X1 U841 ( .A1(n499), .A2(n414), .B1(n413), .B2(n481), .ZN(n337) );
  OAI22_X1 U842 ( .A1(n412), .A2(n481), .B1(n413), .B2(n499), .ZN(n336) );
  OAI22_X1 U843 ( .A1(n404), .A2(n499), .B1(n403), .B2(n481), .ZN(n329) );
  OAI22_X1 U844 ( .A1(n409), .A2(n499), .B1(n408), .B2(n481), .ZN(n332) );
  OAI22_X1 U845 ( .A1(n410), .A2(n481), .B1(n499), .B2(n411), .ZN(n334) );
  INV_X1 U846 ( .A(n493), .ZN(n487) );
  XNOR2_X1 U847 ( .A(n612), .B(n493), .ZN(n414) );
  XNOR2_X1 U848 ( .A(n465), .B(n493), .ZN(n413) );
  XNOR2_X1 U849 ( .A(n456), .B(n493), .ZN(n404) );
  XNOR2_X1 U850 ( .A(n455), .B(n493), .ZN(n403) );
  XNOR2_X1 U851 ( .A(n461), .B(n493), .ZN(n409) );
  XNOR2_X1 U852 ( .A(b[4]), .B(n493), .ZN(n410) );
  XNOR2_X1 U853 ( .A(n464), .B(n493), .ZN(n412) );
  XNOR2_X1 U854 ( .A(n463), .B(n493), .ZN(n411) );
  XNOR2_X1 U855 ( .A(n493), .B(n458), .ZN(n406) );
  XNOR2_X1 U856 ( .A(n493), .B(n457), .ZN(n405) );
  XNOR2_X1 U857 ( .A(n493), .B(n460), .ZN(n408) );
  XNOR2_X1 U858 ( .A(n493), .B(n459), .ZN(n407) );
  OAI21_X1 U859 ( .B1(n135), .B2(n137), .A(n136), .ZN(n134) );
  INV_X1 U860 ( .A(n138), .ZN(n137) );
  INV_X1 U861 ( .A(a[0]), .ZN(n508) );
  INV_X1 U862 ( .A(n187), .ZN(n188) );
  OAI21_X1 U863 ( .B1(n129), .B2(n127), .A(n128), .ZN(n126) );
  XOR2_X1 U864 ( .A(a[7]), .B(a[6]), .Z(n469) );
  AOI21_X1 U865 ( .B1(n126), .B2(n609), .A(n123), .ZN(n121) );
  XNOR2_X1 U866 ( .A(n456), .B(n491), .ZN(n378) );
  XNOR2_X1 U867 ( .A(n455), .B(n491), .ZN(n377) );
  XNOR2_X1 U868 ( .A(b[4]), .B(n491), .ZN(n384) );
  XNOR2_X1 U869 ( .A(n464), .B(n491), .ZN(n386) );
  XNOR2_X1 U870 ( .A(n461), .B(n491), .ZN(n383) );
  XNOR2_X1 U871 ( .A(n463), .B(n491), .ZN(n385) );
  INV_X1 U872 ( .A(n491), .ZN(n485) );
  XNOR2_X1 U873 ( .A(n465), .B(n491), .ZN(n387) );
  XNOR2_X1 U874 ( .A(n458), .B(n491), .ZN(n380) );
  XNOR2_X1 U875 ( .A(n457), .B(n491), .ZN(n379) );
  XNOR2_X1 U876 ( .A(n491), .B(n460), .ZN(n382) );
  XNOR2_X1 U877 ( .A(n459), .B(n491), .ZN(n381) );
  AOI21_X1 U878 ( .B1(n90), .B2(n73), .A(n74), .ZN(n72) );
  OAI21_X1 U879 ( .B1(n83), .B2(n75), .A(n76), .ZN(n74) );
  NAND2_X1 U880 ( .A1(n189), .A2(n184), .ZN(n59) );
  NAND2_X1 U881 ( .A1(n204), .A2(n211), .ZN(n83) );
  AOI21_X1 U882 ( .B1(n44), .B2(n57), .A(n45), .ZN(n43) );
  OAI21_X1 U883 ( .B1(n50), .B2(n46), .A(n47), .ZN(n45) );
  XNOR2_X1 U884 ( .A(a[9]), .B(a[10]), .ZN(n503) );
  AOI21_X1 U885 ( .B1(n108), .B2(n100), .A(n101), .ZN(n99) );
  OAI21_X1 U886 ( .B1(n121), .B2(n109), .A(n110), .ZN(n108) );
  NAND2_X1 U887 ( .A1(n604), .A2(n44), .ZN(n42) );
  AOI21_X1 U888 ( .B1(n602), .B2(n26), .A(n27), .ZN(n25) );
  AND2_X1 U889 ( .A1(n611), .A2(a[0]), .ZN(product[0]) );
  XNOR2_X1 U890 ( .A(n22), .B(n146), .ZN(product[2]) );
  NAND2_X1 U891 ( .A1(n607), .A2(n145), .ZN(n22) );
  XOR2_X1 U892 ( .A(n20), .B(n137), .Z(product[4]) );
  NAND2_X1 U893 ( .A1(n167), .A2(n136), .ZN(n20) );
  XOR2_X1 U894 ( .A(n21), .B(n141), .Z(product[3]) );
  NAND2_X1 U895 ( .A1(n168), .A2(n140), .ZN(n21) );
  XOR2_X1 U896 ( .A(n18), .B(n581), .Z(product[6]) );
  NAND2_X1 U897 ( .A1(n165), .A2(n128), .ZN(n18) );
  AOI21_X1 U898 ( .B1(n610), .B2(n134), .A(n131), .ZN(n129) );
  XNOR2_X1 U899 ( .A(n19), .B(n579), .ZN(product[5]) );
  NAND2_X1 U900 ( .A1(n610), .A2(n133), .ZN(n19) );
  XNOR2_X1 U901 ( .A(n126), .B(n17), .ZN(product[7]) );
  NAND2_X1 U902 ( .A1(n609), .A2(n125), .ZN(n17) );
  XNOR2_X1 U903 ( .A(n120), .B(n16), .ZN(product[8]) );
  INV_X1 U904 ( .A(n121), .ZN(n120) );
  INV_X1 U905 ( .A(n108), .ZN(n107) );
  XNOR2_X1 U906 ( .A(n98), .B(n12), .ZN(product[12]) );
  INV_X1 U907 ( .A(n562), .ZN(n98) );
  AOI21_X1 U908 ( .B1(n602), .B2(n52), .A(n53), .ZN(n51) );
  XNOR2_X1 U909 ( .A(n30), .B(n3), .ZN(product[21]) );
  OAI21_X1 U910 ( .B1(n69), .B2(n31), .A(n32), .ZN(n30) );
  AOI21_X1 U911 ( .B1(n560), .B2(n94), .A(n95), .ZN(n93) );
  XNOR2_X1 U912 ( .A(n48), .B(n5), .ZN(product[19]) );
  OAI21_X1 U913 ( .B1(n49), .B2(n51), .A(n50), .ZN(n48) );
  XOR2_X1 U914 ( .A(n84), .B(n10), .Z(product[14]) );
  AOI21_X1 U915 ( .B1(n98), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U916 ( .B1(n61), .B2(n70), .A(n62), .ZN(n60) );
  XNOR2_X1 U917 ( .A(n37), .B(n4), .ZN(product[20]) );
  OAI21_X1 U918 ( .B1(n69), .B2(n38), .A(n39), .ZN(n37) );
  XOR2_X1 U919 ( .A(n77), .B(n9), .Z(product[15]) );
  AOI21_X1 U920 ( .B1(n78), .B2(n98), .A(n79), .ZN(n77) );
  INV_X1 U921 ( .A(n70), .ZN(n69) );
  INV_X1 U922 ( .A(n25), .ZN(n149) );
endmodule


module datapath_DW_mult_tc_23 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n1, n4, n8, n9, n12, n13, n14, n15, n16, n17, n18, n19, n21, n22, n23,
         n24, n26, n27, n28, n29, n30, n31, n32, n33, n35, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n48, n50, n51, n52, n53, n54, n57, n59,
         n60, n61, n62, n63, n64, n65, n66, n69, n70, n71, n75, n76, n77, n78,
         n80, n81, n82, n83, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n139, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n151, n153, n154, n156, n157,
         n161, n162, n163, n164, n165, n166, n168, n169, n170, n172, n173,
         n175, n176, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n292, n293, n295, n296, n298, n299, n301,
         n302, n305, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n467, n468, n469, n470, n471,
         n472, n473, n475, n476, n477, n478, n479, n482, n484, n485, n487,
         n488, n489, n490, n491, n493, n494, n495, n496, n497, n498, n499,
         n500, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n568, n569, n570, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603;
  assign product[23] = n26;

  FA_X1 U203 ( .A(n314), .B(n185), .CI(n322), .CO(n181), .S(n182) );
  FA_X1 U204 ( .A(n186), .B(n323), .CI(n189), .CO(n183), .S(n184) );
  FA_X1 U206 ( .A(n193), .B(n335), .CI(n190), .CO(n187), .S(n188) );
  FA_X1 U207 ( .A(n315), .B(n195), .CI(n324), .CO(n189), .S(n190) );
  FA_X1 U208 ( .A(n194), .B(n201), .CI(n199), .CO(n191), .S(n192) );
  FA_X1 U209 ( .A(n336), .B(n325), .CI(n196), .CO(n193), .S(n194) );
  FA_X1 U211 ( .A(n205), .B(n202), .CI(n200), .CO(n197), .S(n198) );
  FA_X1 U212 ( .A(n347), .B(n209), .CI(n207), .CO(n199), .S(n200) );
  FA_X1 U213 ( .A(n326), .B(n316), .CI(n337), .CO(n201), .S(n202) );
  FA_X1 U214 ( .A(n213), .B(n208), .CI(n206), .CO(n203), .S(n204) );
  FA_X1 U215 ( .A(n217), .B(n210), .CI(n215), .CO(n205), .S(n206) );
  FA_X1 U216 ( .A(n348), .B(n327), .CI(n317), .CO(n207), .S(n208) );
  FA_X1 U218 ( .A(n221), .B(n216), .CI(n214), .CO(n211), .S(n212) );
  FA_X1 U219 ( .A(n223), .B(n225), .CI(n218), .CO(n213), .S(n214) );
  FA_X1 U220 ( .A(n360), .B(n328), .CI(n318), .CO(n215), .S(n216) );
  FA_X1 U221 ( .A(n338), .B(n576), .CI(n349), .CO(n217), .S(n218) );
  FA_X1 U222 ( .A(n231), .B(n224), .CI(n222), .CO(n219), .S(n220) );
  FA_X1 U223 ( .A(n226), .B(n235), .CI(n233), .CO(n221), .S(n222) );
  FA_X1 U224 ( .A(n329), .B(n228), .CI(n237), .CO(n223), .S(n224) );
  FA_X1 U225 ( .A(n350), .B(n339), .CI(n361), .CO(n225), .S(n226) );
  FA_X1 U227 ( .A(n241), .B(n234), .CI(n232), .CO(n229), .S(n230) );
  FA_X1 U228 ( .A(n236), .B(n245), .CI(n243), .CO(n231), .S(n232) );
  FA_X1 U229 ( .A(n247), .B(n330), .CI(n238), .CO(n233), .S(n234) );
  FA_X1 U230 ( .A(n319), .B(n340), .CI(n572), .CO(n235), .S(n236) );
  FA_X1 U233 ( .A(n251), .B(n244), .CI(n242), .CO(n239), .S(n240) );
  FA_X1 U234 ( .A(n253), .B(n255), .CI(n246), .CO(n241), .S(n242) );
  FA_X1 U235 ( .A(n341), .B(n320), .CI(n248), .CO(n243), .S(n244) );
  FA_X1 U236 ( .A(n352), .B(n331), .CI(n374), .CO(n245), .S(n246) );
  HA_X1 U237 ( .A(n307), .B(n363), .CO(n247), .S(n248) );
  FA_X1 U238 ( .A(n259), .B(n254), .CI(n252), .CO(n249), .S(n250) );
  FA_X1 U239 ( .A(n261), .B(n263), .CI(n256), .CO(n251), .S(n252) );
  FA_X1 U240 ( .A(n332), .B(n353), .CI(n342), .CO(n253), .S(n254) );
  FA_X1 U241 ( .A(n364), .B(n321), .CI(n375), .CO(n255), .S(n256) );
  FA_X1 U242 ( .A(n262), .B(n267), .CI(n260), .CO(n257), .S(n258) );
  FA_X1 U243 ( .A(n264), .B(n354), .CI(n269), .CO(n259), .S(n260) );
  FA_X1 U244 ( .A(n333), .B(n308), .CI(n343), .CO(n261), .S(n262) );
  HA_X1 U245 ( .A(n376), .B(n365), .CO(n263), .S(n264) );
  FA_X1 U246 ( .A(n270), .B(n273), .CI(n268), .CO(n265), .S(n266) );
  FA_X1 U247 ( .A(n275), .B(n355), .CI(n344), .CO(n267), .S(n268) );
  FA_X1 U248 ( .A(n377), .B(n334), .CI(n366), .CO(n269), .S(n270) );
  FA_X1 U249 ( .A(n279), .B(n276), .CI(n274), .CO(n271), .S(n272) );
  FA_X1 U250 ( .A(n356), .B(n345), .CI(n367), .CO(n273), .S(n274) );
  HA_X1 U251 ( .A(n378), .B(n309), .CO(n275), .S(n276) );
  FA_X1 U252 ( .A(n283), .B(n368), .CI(n280), .CO(n277), .S(n278) );
  FA_X1 U253 ( .A(n379), .B(n346), .CI(n357), .CO(n279), .S(n280) );
  FA_X1 U254 ( .A(n380), .B(n358), .CI(n284), .CO(n281), .S(n282) );
  HA_X1 U255 ( .A(n310), .B(n369), .CO(n283), .S(n284) );
  FA_X1 U256 ( .A(n370), .B(n359), .CI(n381), .CO(n285), .S(n286) );
  HA_X1 U257 ( .A(n382), .B(n311), .CO(n287), .S(n288) );
  OAI21_X1 U493 ( .B1(n577), .B2(n111), .A(n106), .ZN(n568) );
  CLKBUF_X1 U494 ( .A(n454), .Z(n569) );
  CLKBUF_X1 U495 ( .A(b[5]), .Z(n469) );
  BUF_X4 U496 ( .A(a[1]), .Z(n504) );
  CLKBUF_X3 U497 ( .A(b[7]), .Z(n467) );
  BUF_X2 U498 ( .A(b[2]), .Z(n472) );
  CLKBUF_X3 U499 ( .A(a[11]), .Z(n499) );
  OR2_X1 U500 ( .A1(n181), .A2(n180), .ZN(n570) );
  AND2_X1 U501 ( .A1(n600), .A2(n156), .ZN(product[1]) );
  OR2_X1 U502 ( .A1(n582), .A2(n450), .ZN(n572) );
  OR2_X1 U503 ( .A1(n581), .A2(n271), .ZN(n573) );
  CLKBUF_X3 U504 ( .A(n515), .Z(n491) );
  CLKBUF_X2 U505 ( .A(b[9]), .Z(n465) );
  BUF_X1 U506 ( .A(b[6]), .Z(n468) );
  BUF_X2 U507 ( .A(b[0]), .Z(n1) );
  INV_X1 U508 ( .A(n584), .ZN(n574) );
  BUF_X2 U509 ( .A(b[3]), .Z(n471) );
  BUF_X2 U510 ( .A(n509), .Z(n575) );
  BUF_X2 U511 ( .A(n509), .Z(n485) );
  OAI22_X1 U512 ( .A1(n394), .A2(n505), .B1(n487), .B2(n393), .ZN(n576) );
  NOR2_X1 U513 ( .A1(n220), .A2(n229), .ZN(n577) );
  CLKBUF_X1 U514 ( .A(n507), .Z(n578) );
  BUF_X4 U515 ( .A(n513), .Z(n489) );
  OR2_X2 U516 ( .A1(n579), .A2(a[0]), .ZN(n510) );
  XNOR2_X1 U517 ( .A(a[1]), .B(a[0]), .ZN(n579) );
  BUF_X1 U518 ( .A(n596), .Z(n593) );
  CLKBUF_X1 U519 ( .A(n125), .Z(n580) );
  BUF_X2 U520 ( .A(b[1]), .Z(n473) );
  BUF_X2 U521 ( .A(n506), .Z(n482) );
  CLKBUF_X1 U522 ( .A(n266), .Z(n581) );
  NAND2_X2 U523 ( .A1(n475), .A2(n511), .ZN(n505) );
  CLKBUF_X1 U524 ( .A(b[4]), .Z(n470) );
  AND2_X1 U525 ( .A1(n510), .A2(n516), .ZN(n582) );
  XNOR2_X1 U526 ( .A(n51), .B(n583), .ZN(product[20]) );
  AND2_X1 U527 ( .A1(n597), .A2(n50), .ZN(n583) );
  CLKBUF_X1 U528 ( .A(n83), .Z(n584) );
  CLKBUF_X1 U529 ( .A(n137), .Z(n585) );
  NOR2_X1 U530 ( .A1(n220), .A2(n229), .ZN(n105) );
  CLKBUF_X3 U531 ( .A(a[3]), .Z(n503) );
  BUF_X1 U532 ( .A(n129), .Z(n586) );
  XNOR2_X1 U533 ( .A(n587), .B(n585), .ZN(product[6]) );
  AND2_X1 U534 ( .A1(n173), .A2(n136), .ZN(n587) );
  XNOR2_X1 U535 ( .A(n83), .B(n588), .ZN(product[16]) );
  AND2_X1 U536 ( .A1(n163), .A2(n82), .ZN(n588) );
  XNOR2_X1 U537 ( .A(n60), .B(n589), .ZN(product[19]) );
  AND2_X1 U538 ( .A1(n598), .A2(n59), .ZN(n589) );
  BUF_X2 U539 ( .A(a[7]), .Z(n603) );
  XNOR2_X1 U540 ( .A(n91), .B(n590), .ZN(product[15]) );
  AND2_X1 U541 ( .A1(n164), .A2(n90), .ZN(n590) );
  XNOR2_X1 U542 ( .A(n38), .B(n591), .ZN(product[21]) );
  AND2_X1 U543 ( .A1(n570), .A2(n37), .ZN(n591) );
  NAND2_X2 U544 ( .A1(n513), .A2(n477), .ZN(n507) );
  NOR2_X1 U545 ( .A1(n240), .A2(n249), .ZN(n592) );
  OAI21_X1 U546 ( .B1(n85), .B2(n113), .A(n86), .ZN(n596) );
  NOR2_X1 U547 ( .A1(n266), .A2(n271), .ZN(n594) );
  NOR2_X1 U548 ( .A1(n266), .A2(n271), .ZN(n595) );
  XOR2_X1 U549 ( .A(n133), .B(n19), .Z(product[7]) );
  NOR2_X1 U550 ( .A1(n191), .A2(n188), .ZN(n69) );
  OR2_X1 U551 ( .A1(n183), .A2(n182), .ZN(n597) );
  OR2_X1 U552 ( .A1(n184), .A2(n187), .ZN(n598) );
  OR2_X1 U553 ( .A1(n383), .A2(n372), .ZN(n599) );
  OR2_X1 U554 ( .A1(n384), .A2(n312), .ZN(n600) );
  OR2_X1 U555 ( .A1(n282), .A2(n285), .ZN(n601) );
  BUF_X2 U556 ( .A(n511), .Z(n487) );
  BUF_X2 U557 ( .A(a[5]), .Z(n502) );
  BUF_X2 U558 ( .A(a[9]), .Z(n500) );
  BUF_X1 U559 ( .A(b[10]), .Z(n464) );
  BUF_X1 U560 ( .A(a[7]), .Z(n602) );
  INV_X1 U561 ( .A(n29), .ZN(n157) );
  NAND2_X1 U562 ( .A1(n157), .A2(n30), .ZN(n4) );
  NOR2_X1 U563 ( .A1(n313), .A2(n179), .ZN(n29) );
  INV_X1 U564 ( .A(n37), .ZN(n35) );
  NAND2_X1 U565 ( .A1(n181), .A2(n180), .ZN(n37) );
  INV_X1 U566 ( .A(n295), .ZN(n335) );
  NAND2_X1 U567 ( .A1(n183), .A2(n182), .ZN(n50) );
  INV_X1 U568 ( .A(n50), .ZN(n48) );
  INV_X1 U569 ( .A(n598), .ZN(n54) );
  NOR2_X1 U570 ( .A1(n69), .A2(n45), .ZN(n43) );
  NOR2_X1 U571 ( .A1(n198), .A2(n203), .ZN(n81) );
  NOR2_X1 U572 ( .A1(n197), .A2(n192), .ZN(n76) );
  AND2_X1 U573 ( .A1(n1), .A2(n302), .ZN(n372) );
  OAI21_X1 U574 ( .B1(n41), .B2(n82), .A(n42), .ZN(n40) );
  NAND2_X1 U575 ( .A1(n198), .A2(n203), .ZN(n82) );
  NAND2_X1 U576 ( .A1(n170), .A2(n124), .ZN(n17) );
  XNOR2_X1 U577 ( .A(n602), .B(n468), .ZN(n416) );
  INV_X1 U578 ( .A(n82), .ZN(n80) );
  NAND2_X1 U579 ( .A1(n258), .A2(n265), .ZN(n124) );
  XNOR2_X1 U580 ( .A(n602), .B(n471), .ZN(n419) );
  XNOR2_X1 U581 ( .A(n603), .B(n467), .ZN(n415) );
  AOI21_X1 U582 ( .B1(n599), .B2(n154), .A(n151), .ZN(n149) );
  BUF_X2 U583 ( .A(n514), .Z(n490) );
  BUF_X2 U584 ( .A(n512), .Z(n488) );
  AOI21_X1 U585 ( .B1(n484), .B2(n490), .A(n424), .ZN(n298) );
  INV_X1 U586 ( .A(n59), .ZN(n57) );
  AOI21_X1 U587 ( .B1(n57), .B2(n597), .A(n48), .ZN(n46) );
  INV_X1 U588 ( .A(n292), .ZN(n322) );
  CLKBUF_X1 U589 ( .A(b[11]), .Z(n463) );
  OAI22_X1 U590 ( .A1(n484), .A2(n426), .B1(n425), .B2(n490), .ZN(n349) );
  INV_X1 U591 ( .A(n298), .ZN(n347) );
  OAI22_X1 U592 ( .A1(n484), .A2(n435), .B1(n434), .B2(n490), .ZN(n358) );
  NAND2_X1 U593 ( .A1(n286), .A2(n287), .ZN(n144) );
  OAI22_X1 U594 ( .A1(n510), .A2(n453), .B1(n452), .B2(n516), .ZN(n376) );
  OAI22_X1 U595 ( .A1(n457), .A2(n516), .B1(n510), .B2(n458), .ZN(n381) );
  OAI22_X1 U596 ( .A1(n482), .A2(n402), .B1(n401), .B2(n488), .ZN(n326) );
  OAI22_X1 U597 ( .A1(n482), .A2(n403), .B1(n402), .B2(n488), .ZN(n327) );
  OAI22_X1 U598 ( .A1(n482), .A2(n404), .B1(n403), .B2(n488), .ZN(n328) );
  OAI22_X1 U599 ( .A1(n482), .A2(n494), .B1(n410), .B2(n488), .ZN(n308) );
  AOI21_X1 U600 ( .B1(n482), .B2(n488), .A(n398), .ZN(n292) );
  OAI22_X1 U601 ( .A1(n482), .A2(n401), .B1(n400), .B2(n488), .ZN(n325) );
  INV_X1 U602 ( .A(n76), .ZN(n162) );
  NAND2_X1 U603 ( .A1(n162), .A2(n77), .ZN(n9) );
  INV_X1 U604 ( .A(n77), .ZN(n75) );
  OAI22_X1 U605 ( .A1(n505), .A2(n390), .B1(n487), .B2(n389), .ZN(n195) );
  OAI22_X1 U606 ( .A1(n484), .A2(n427), .B1(n426), .B2(n490), .ZN(n350) );
  XNOR2_X1 U607 ( .A(a[3]), .B(a[4]), .ZN(n514) );
  OAI22_X1 U608 ( .A1(n484), .A2(n429), .B1(n428), .B2(n490), .ZN(n352) );
  BUF_X2 U609 ( .A(n508), .Z(n484) );
  OAI22_X1 U610 ( .A1(n405), .A2(n482), .B1(n404), .B2(n488), .ZN(n329) );
  XOR2_X1 U611 ( .A(a[9]), .B(a[8]), .Z(n476) );
  NAND2_X1 U612 ( .A1(n197), .A2(n192), .ZN(n77) );
  OAI22_X1 U613 ( .A1(n394), .A2(n505), .B1(n487), .B2(n393), .ZN(n227) );
  OAI22_X1 U614 ( .A1(n510), .A2(n569), .B1(n453), .B2(n516), .ZN(n377) );
  OAI22_X1 U615 ( .A1(n578), .A2(n413), .B1(n412), .B2(n489), .ZN(n337) );
  OAI22_X1 U616 ( .A1(n578), .A2(n414), .B1(n413), .B2(n489), .ZN(n209) );
  AOI21_X1 U617 ( .B1(n578), .B2(n489), .A(n411), .ZN(n295) );
  OAI22_X1 U618 ( .A1(n507), .A2(n415), .B1(n414), .B2(n489), .ZN(n338) );
  OAI22_X1 U619 ( .A1(n507), .A2(n416), .B1(n415), .B2(n489), .ZN(n339) );
  NAND2_X1 U620 ( .A1(n204), .A2(n211), .ZN(n90) );
  NOR2_X1 U621 ( .A1(n272), .A2(n277), .ZN(n131) );
  XOR2_X1 U622 ( .A(a[10]), .B(a[11]), .Z(n475) );
  INV_X1 U623 ( .A(n102), .ZN(n100) );
  INV_X1 U624 ( .A(n165), .ZN(n94) );
  XNOR2_X1 U625 ( .A(n602), .B(n465), .ZN(n413) );
  NOR2_X1 U626 ( .A1(n250), .A2(n257), .ZN(n119) );
  NAND2_X1 U627 ( .A1(n598), .A2(n597), .ZN(n45) );
  NOR2_X1 U628 ( .A1(n204), .A2(n211), .ZN(n89) );
  NOR2_X1 U629 ( .A1(n212), .A2(n219), .ZN(n96) );
  INV_X1 U630 ( .A(n156), .ZN(n154) );
  OAI22_X1 U631 ( .A1(n431), .A2(n484), .B1(n430), .B2(n490), .ZN(n354) );
  INV_X1 U632 ( .A(n153), .ZN(n151) );
  OAI22_X1 U633 ( .A1(n507), .A2(n421), .B1(n420), .B2(n489), .ZN(n344) );
  NAND2_X1 U634 ( .A1(n272), .A2(n277), .ZN(n132) );
  XNOR2_X1 U635 ( .A(n473), .B(n602), .ZN(n421) );
  INV_X1 U636 ( .A(n103), .ZN(n101) );
  NOR2_X1 U637 ( .A1(n110), .A2(n105), .ZN(n103) );
  XOR2_X1 U638 ( .A(a[7]), .B(a[6]), .Z(n477) );
  INV_X1 U639 ( .A(n101), .ZN(n99) );
  INV_X1 U640 ( .A(n147), .ZN(n176) );
  NOR2_X1 U641 ( .A1(n288), .A2(n371), .ZN(n147) );
  OAI22_X1 U642 ( .A1(n507), .A2(n417), .B1(n416), .B2(n489), .ZN(n340) );
  XNOR2_X1 U643 ( .A(n469), .B(n602), .ZN(n417) );
  INV_X1 U644 ( .A(n141), .ZN(n139) );
  NAND2_X1 U645 ( .A1(n266), .A2(n271), .ZN(n129) );
  OAI22_X1 U646 ( .A1(n455), .A2(n510), .B1(n454), .B2(n516), .ZN(n378) );
  INV_X1 U647 ( .A(n135), .ZN(n173) );
  NOR2_X1 U648 ( .A1(n278), .A2(n281), .ZN(n135) );
  INV_X1 U649 ( .A(n592), .ZN(n168) );
  NOR2_X1 U650 ( .A1(n32), .A2(n29), .ZN(n27) );
  NOR2_X1 U651 ( .A1(n101), .A2(n94), .ZN(n92) );
  NAND2_X1 U652 ( .A1(n278), .A2(n281), .ZN(n136) );
  INV_X1 U653 ( .A(n143), .ZN(n175) );
  NOR2_X1 U654 ( .A1(n286), .A2(n287), .ZN(n143) );
  OAI22_X1 U655 ( .A1(n507), .A2(n495), .B1(n423), .B2(n489), .ZN(n309) );
  NOR2_X1 U656 ( .A1(n76), .A2(n69), .ZN(n65) );
  OAI22_X1 U657 ( .A1(n484), .A2(n434), .B1(n433), .B2(n490), .ZN(n357) );
  INV_X1 U658 ( .A(n81), .ZN(n163) );
  OAI22_X1 U659 ( .A1(n457), .A2(n510), .B1(n456), .B2(n516), .ZN(n380) );
  OAI22_X1 U660 ( .A1(n456), .A2(n510), .B1(n455), .B2(n516), .ZN(n379) );
  INV_X1 U661 ( .A(n69), .ZN(n161) );
  NAND2_X1 U662 ( .A1(n161), .A2(n70), .ZN(n8) );
  OAI21_X1 U663 ( .B1(n45), .B2(n70), .A(n46), .ZN(n44) );
  OAI21_X1 U664 ( .B1(n77), .B2(n69), .A(n70), .ZN(n66) );
  AOI21_X1 U665 ( .B1(n43), .B2(n75), .A(n44), .ZN(n42) );
  NAND2_X1 U666 ( .A1(n65), .A2(n163), .ZN(n63) );
  NAND2_X1 U667 ( .A1(n282), .A2(n285), .ZN(n141) );
  OAI22_X1 U668 ( .A1(n484), .A2(n496), .B1(n436), .B2(n490), .ZN(n310) );
  OAI22_X1 U669 ( .A1(n431), .A2(n490), .B1(n484), .B2(n432), .ZN(n355) );
  NAND2_X1 U670 ( .A1(n191), .A2(n188), .ZN(n70) );
  INV_X1 U671 ( .A(n489), .ZN(n296) );
  OAI21_X1 U672 ( .B1(n143), .B2(n145), .A(n144), .ZN(n142) );
  OAI22_X1 U673 ( .A1(n459), .A2(n510), .B1(n458), .B2(n516), .ZN(n382) );
  INV_X1 U674 ( .A(n490), .ZN(n299) );
  OAI22_X1 U675 ( .A1(n484), .A2(n425), .B1(n424), .B2(n490), .ZN(n348) );
  NAND2_X1 U676 ( .A1(n384), .A2(n312), .ZN(n156) );
  OAI22_X1 U677 ( .A1(n510), .A2(n461), .B1(n460), .B2(n516), .ZN(n384) );
  AOI21_X1 U678 ( .B1(n601), .B2(n142), .A(n139), .ZN(n137) );
  NAND2_X1 U679 ( .A1(n383), .A2(n372), .ZN(n153) );
  OAI22_X1 U680 ( .A1(n459), .A2(n516), .B1(n510), .B2(n460), .ZN(n383) );
  NOR2_X1 U681 ( .A1(n63), .A2(n54), .ZN(n52) );
  INV_X1 U682 ( .A(n119), .ZN(n169) );
  NAND2_X1 U683 ( .A1(n169), .A2(n120), .ZN(n16) );
  OAI21_X1 U684 ( .B1(n33), .B2(n29), .A(n30), .ZN(n28) );
  AOI21_X1 U685 ( .B1(n40), .B2(n570), .A(n35), .ZN(n33) );
  NAND2_X1 U686 ( .A1(n39), .A2(n570), .ZN(n32) );
  NOR2_X1 U687 ( .A1(n81), .A2(n41), .ZN(n39) );
  INV_X1 U688 ( .A(n488), .ZN(n293) );
  INV_X1 U689 ( .A(n131), .ZN(n172) );
  OAI22_X1 U690 ( .A1(n507), .A2(n420), .B1(n419), .B2(n489), .ZN(n343) );
  OR2_X1 U691 ( .A1(n1), .A2(n496), .ZN(n436) );
  OR2_X1 U692 ( .A1(n1), .A2(n494), .ZN(n410) );
  OR2_X1 U693 ( .A1(n1), .A2(n497), .ZN(n449) );
  AND2_X1 U694 ( .A1(n1), .A2(n296), .ZN(n346) );
  AND2_X1 U695 ( .A1(n1), .A2(n299), .ZN(n359) );
  AND2_X1 U696 ( .A1(n1), .A2(n293), .ZN(n334) );
  OR2_X1 U697 ( .A1(n493), .A2(n1), .ZN(n397) );
  OR2_X1 U698 ( .A1(n1), .A2(n495), .ZN(n423) );
  OR2_X1 U699 ( .A1(n1), .A2(n498), .ZN(n462) );
  INV_X1 U700 ( .A(n63), .ZN(n61) );
  OAI22_X1 U701 ( .A1(n484), .A2(n433), .B1(n432), .B2(n490), .ZN(n356) );
  INV_X1 U702 ( .A(n96), .ZN(n165) );
  NOR2_X1 U703 ( .A1(n96), .A2(n89), .ZN(n87) );
  NAND2_X1 U704 ( .A1(n165), .A2(n97), .ZN(n12) );
  OAI21_X1 U705 ( .B1(n97), .B2(n89), .A(n90), .ZN(n88) );
  OAI21_X1 U706 ( .B1(n102), .B2(n94), .A(n97), .ZN(n93) );
  INV_X1 U707 ( .A(n89), .ZN(n164) );
  INV_X1 U708 ( .A(n146), .ZN(n145) );
  OAI21_X1 U709 ( .B1(n116), .B2(n120), .A(n117), .ZN(n115) );
  NOR2_X1 U710 ( .A1(n592), .A2(n119), .ZN(n114) );
  NAND2_X1 U711 ( .A1(n168), .A2(n117), .ZN(n15) );
  NOR2_X1 U712 ( .A1(n240), .A2(n249), .ZN(n116) );
  NAND2_X1 U713 ( .A1(n573), .A2(n586), .ZN(n18) );
  NAND2_X1 U714 ( .A1(n212), .A2(n219), .ZN(n97) );
  NAND2_X1 U715 ( .A1(n250), .A2(n257), .ZN(n120) );
  OAI22_X1 U716 ( .A1(n482), .A2(n408), .B1(n407), .B2(n488), .ZN(n332) );
  OAI22_X1 U717 ( .A1(n451), .A2(n516), .B1(n510), .B2(n452), .ZN(n375) );
  OAI22_X1 U718 ( .A1(n451), .A2(n510), .B1(n450), .B2(n516), .ZN(n374) );
  XNOR2_X1 U719 ( .A(n472), .B(n603), .ZN(n420) );
  OAI22_X1 U720 ( .A1(n484), .A2(n430), .B1(n429), .B2(n490), .ZN(n353) );
  INV_X1 U721 ( .A(n105), .ZN(n166) );
  NAND2_X1 U722 ( .A1(n166), .A2(n106), .ZN(n13) );
  NAND2_X1 U723 ( .A1(n103), .A2(n87), .ZN(n85) );
  INV_X1 U724 ( .A(n568), .ZN(n102) );
  OAI22_X1 U725 ( .A1(n507), .A2(n422), .B1(n421), .B2(n489), .ZN(n345) );
  XNOR2_X1 U726 ( .A(n1), .B(n602), .ZN(n422) );
  OAI22_X1 U727 ( .A1(n405), .A2(n488), .B1(n482), .B2(n406), .ZN(n330) );
  OAI22_X1 U728 ( .A1(n418), .A2(n489), .B1(n507), .B2(n419), .ZN(n342) );
  OAI22_X1 U729 ( .A1(n418), .A2(n507), .B1(n417), .B2(n489), .ZN(n341) );
  INV_X1 U730 ( .A(n491), .ZN(n302) );
  OAI22_X1 U731 ( .A1(n447), .A2(n491), .B1(n575), .B2(n448), .ZN(n371) );
  OAI22_X1 U732 ( .A1(n446), .A2(n491), .B1(n447), .B2(n575), .ZN(n370) );
  OAI22_X1 U733 ( .A1(n446), .A2(n485), .B1(n445), .B2(n491), .ZN(n369) );
  OAI22_X1 U734 ( .A1(n444), .A2(n491), .B1(n575), .B2(n445), .ZN(n368) );
  OAI22_X1 U735 ( .A1(n444), .A2(n575), .B1(n443), .B2(n491), .ZN(n367) );
  OAI22_X1 U736 ( .A1(n443), .A2(n575), .B1(n442), .B2(n491), .ZN(n366) );
  OAI22_X1 U737 ( .A1(n575), .A2(n442), .B1(n441), .B2(n491), .ZN(n365) );
  OAI22_X1 U738 ( .A1(n485), .A2(n441), .B1(n440), .B2(n491), .ZN(n364) );
  OAI22_X1 U739 ( .A1(n440), .A2(n485), .B1(n439), .B2(n491), .ZN(n363) );
  AOI21_X1 U740 ( .B1(n575), .B2(n491), .A(n437), .ZN(n301) );
  OAI22_X1 U741 ( .A1(n485), .A2(n497), .B1(n449), .B2(n491), .ZN(n311) );
  NAND2_X1 U742 ( .A1(n288), .A2(n371), .ZN(n148) );
  OR2_X1 U743 ( .A1(n351), .A2(n362), .ZN(n237) );
  OAI22_X1 U744 ( .A1(n484), .A2(n428), .B1(n427), .B2(n490), .ZN(n351) );
  OAI22_X1 U745 ( .A1(n482), .A2(n409), .B1(n408), .B2(n488), .ZN(n333) );
  NAND2_X1 U746 ( .A1(n162), .A2(n43), .ZN(n41) );
  OAI22_X1 U747 ( .A1(n482), .A2(n407), .B1(n406), .B2(n488), .ZN(n331) );
  XNOR2_X1 U748 ( .A(n470), .B(n603), .ZN(n418) );
  NAND2_X1 U749 ( .A1(n184), .A2(n187), .ZN(n59) );
  NAND2_X1 U750 ( .A1(n220), .A2(n229), .ZN(n106) );
  INV_X1 U751 ( .A(n64), .ZN(n62) );
  OAI21_X1 U752 ( .B1(n64), .B2(n54), .A(n59), .ZN(n53) );
  AOI21_X1 U753 ( .B1(n65), .B2(n80), .A(n66), .ZN(n64) );
  OAI22_X1 U754 ( .A1(n482), .A2(n400), .B1(n399), .B2(n488), .ZN(n324) );
  OAI22_X1 U755 ( .A1(n482), .A2(n399), .B1(n398), .B2(n488), .ZN(n323) );
  OAI22_X1 U756 ( .A1(n438), .A2(n491), .B1(n485), .B2(n439), .ZN(n362) );
  OAI22_X1 U757 ( .A1(n438), .A2(n575), .B1(n437), .B2(n491), .ZN(n361) );
  OAI22_X1 U758 ( .A1(n578), .A2(n412), .B1(n411), .B2(n489), .ZN(n336) );
  XNOR2_X1 U759 ( .A(n463), .B(n602), .ZN(n411) );
  XNOR2_X1 U760 ( .A(n464), .B(n602), .ZN(n412) );
  NAND2_X1 U761 ( .A1(n478), .A2(n514), .ZN(n508) );
  XOR2_X1 U762 ( .A(a[5]), .B(a[4]), .Z(n478) );
  INV_X1 U763 ( .A(n123), .ZN(n170) );
  OAI21_X1 U764 ( .B1(n125), .B2(n123), .A(n124), .ZN(n122) );
  NOR2_X1 U765 ( .A1(n258), .A2(n265), .ZN(n123) );
  INV_X1 U766 ( .A(n110), .ZN(n108) );
  NAND2_X1 U767 ( .A1(n108), .A2(n111), .ZN(n14) );
  OAI21_X1 U768 ( .B1(n577), .B2(n111), .A(n106), .ZN(n104) );
  INV_X1 U769 ( .A(n111), .ZN(n109) );
  NOR2_X1 U770 ( .A1(n230), .A2(n239), .ZN(n110) );
  XNOR2_X1 U771 ( .A(a[1]), .B(a[2]), .ZN(n515) );
  NAND2_X1 U772 ( .A1(n476), .A2(n512), .ZN(n506) );
  XNOR2_X1 U773 ( .A(a[7]), .B(a[8]), .ZN(n512) );
  AOI21_X1 U774 ( .B1(n104), .B2(n87), .A(n88), .ZN(n86) );
  NAND2_X1 U775 ( .A1(n479), .A2(n515), .ZN(n509) );
  XOR2_X1 U776 ( .A(a[3]), .B(a[2]), .Z(n479) );
  XNOR2_X1 U777 ( .A(n362), .B(n351), .ZN(n238) );
  INV_X1 U778 ( .A(n301), .ZN(n360) );
  AOI21_X1 U779 ( .B1(n122), .B2(n114), .A(n115), .ZN(n113) );
  NOR2_X1 U780 ( .A1(n595), .A2(n131), .ZN(n126) );
  NAND2_X1 U781 ( .A1(n230), .A2(n239), .ZN(n111) );
  XNOR2_X1 U782 ( .A(n470), .B(n504), .ZN(n457) );
  XNOR2_X1 U783 ( .A(n469), .B(n504), .ZN(n456) );
  XNOR2_X1 U784 ( .A(n464), .B(n504), .ZN(n451) );
  XNOR2_X1 U785 ( .A(n504), .B(n465), .ZN(n452) );
  XNOR2_X1 U786 ( .A(n504), .B(b[8]), .ZN(n453) );
  XNOR2_X1 U787 ( .A(n1), .B(n504), .ZN(n461) );
  XNOR2_X1 U788 ( .A(n504), .B(n467), .ZN(n454) );
  XNOR2_X1 U789 ( .A(n504), .B(n468), .ZN(n455) );
  XNOR2_X1 U790 ( .A(n473), .B(n504), .ZN(n460) );
  XNOR2_X1 U791 ( .A(n472), .B(n504), .ZN(n459) );
  XNOR2_X1 U792 ( .A(n463), .B(n504), .ZN(n450) );
  XNOR2_X1 U793 ( .A(n471), .B(n504), .ZN(n458) );
  INV_X1 U794 ( .A(n500), .ZN(n494) );
  XNOR2_X1 U795 ( .A(n1), .B(n500), .ZN(n409) );
  XNOR2_X1 U796 ( .A(n500), .B(n467), .ZN(n402) );
  XNOR2_X1 U797 ( .A(n463), .B(n500), .ZN(n398) );
  XNOR2_X1 U798 ( .A(n470), .B(n500), .ZN(n405) );
  XNOR2_X1 U799 ( .A(n500), .B(n468), .ZN(n403) );
  XNOR2_X1 U800 ( .A(n473), .B(n500), .ZN(n408) );
  XNOR2_X1 U801 ( .A(n469), .B(n500), .ZN(n404) );
  XNOR2_X1 U802 ( .A(n500), .B(b[8]), .ZN(n401) );
  XNOR2_X1 U803 ( .A(n500), .B(n465), .ZN(n400) );
  XNOR2_X1 U804 ( .A(n472), .B(n500), .ZN(n407) );
  XNOR2_X1 U805 ( .A(n464), .B(n500), .ZN(n399) );
  XNOR2_X1 U806 ( .A(n500), .B(n471), .ZN(n406) );
  XNOR2_X1 U807 ( .A(n603), .B(b[8]), .ZN(n414) );
  INV_X1 U808 ( .A(n603), .ZN(n495) );
  NAND2_X1 U809 ( .A1(n240), .A2(n249), .ZN(n117) );
  INV_X1 U810 ( .A(n209), .ZN(n210) );
  XNOR2_X1 U811 ( .A(a[5]), .B(a[6]), .ZN(n513) );
  INV_X1 U812 ( .A(a[0]), .ZN(n516) );
  INV_X1 U813 ( .A(n487), .ZN(n290) );
  OAI22_X1 U814 ( .A1(n505), .A2(n396), .B1(n395), .B2(n487), .ZN(n320) );
  OAI22_X1 U815 ( .A1(n394), .A2(n487), .B1(n505), .B2(n395), .ZN(n319) );
  OAI22_X1 U816 ( .A1(n392), .A2(n487), .B1(n505), .B2(n393), .ZN(n318) );
  OAI22_X1 U817 ( .A1(n392), .A2(n505), .B1(n391), .B2(n487), .ZN(n317) );
  OAI22_X1 U818 ( .A1(n391), .A2(n505), .B1(n487), .B2(n390), .ZN(n316) );
  OAI22_X1 U819 ( .A1(n505), .A2(n389), .B1(n487), .B2(n388), .ZN(n315) );
  OAI22_X1 U820 ( .A1(n505), .A2(n388), .B1(n487), .B2(n387), .ZN(n185) );
  OAI22_X1 U821 ( .A1(n386), .A2(n487), .B1(n505), .B2(n387), .ZN(n314) );
  OAI22_X1 U822 ( .A1(n386), .A2(n505), .B1(n385), .B2(n487), .ZN(n179) );
  AOI21_X1 U823 ( .B1(n505), .B2(n487), .A(n385), .ZN(n289) );
  OAI22_X1 U824 ( .A1(n505), .A2(n493), .B1(n397), .B2(n487), .ZN(n307) );
  AND2_X1 U825 ( .A1(n1), .A2(n290), .ZN(n321) );
  INV_X1 U826 ( .A(n227), .ZN(n228) );
  INV_X1 U827 ( .A(n195), .ZN(n196) );
  INV_X1 U828 ( .A(n185), .ZN(n186) );
  NAND2_X1 U829 ( .A1(n313), .A2(n179), .ZN(n30) );
  INV_X1 U830 ( .A(n179), .ZN(n180) );
  INV_X1 U831 ( .A(n289), .ZN(n313) );
  AOI21_X1 U832 ( .B1(n134), .B2(n126), .A(n127), .ZN(n125) );
  OAI21_X1 U833 ( .B1(n594), .B2(n132), .A(n129), .ZN(n127) );
  OAI21_X1 U834 ( .B1(n135), .B2(n137), .A(n136), .ZN(n134) );
  OAI21_X1 U835 ( .B1(n147), .B2(n149), .A(n148), .ZN(n146) );
  XNOR2_X1 U836 ( .A(n463), .B(n499), .ZN(n385) );
  XNOR2_X1 U837 ( .A(n464), .B(n499), .ZN(n386) );
  XNOR2_X1 U838 ( .A(n469), .B(n499), .ZN(n391) );
  XNOR2_X1 U839 ( .A(n470), .B(n499), .ZN(n392) );
  XNOR2_X1 U840 ( .A(n1), .B(n499), .ZN(n396) );
  INV_X1 U841 ( .A(n499), .ZN(n493) );
  XNOR2_X1 U842 ( .A(n473), .B(n499), .ZN(n395) );
  XNOR2_X1 U843 ( .A(n499), .B(b[8]), .ZN(n388) );
  XNOR2_X1 U844 ( .A(n499), .B(n465), .ZN(n387) );
  XNOR2_X1 U845 ( .A(n499), .B(n468), .ZN(n390) );
  XNOR2_X1 U846 ( .A(n472), .B(n499), .ZN(n394) );
  XNOR2_X1 U847 ( .A(n467), .B(n499), .ZN(n389) );
  XNOR2_X1 U848 ( .A(n471), .B(n499), .ZN(n393) );
  XNOR2_X1 U849 ( .A(a[9]), .B(a[10]), .ZN(n511) );
  XNOR2_X1 U850 ( .A(n463), .B(n502), .ZN(n424) );
  XNOR2_X1 U851 ( .A(n469), .B(n502), .ZN(n430) );
  XNOR2_X1 U852 ( .A(n464), .B(n502), .ZN(n425) );
  XNOR2_X1 U853 ( .A(n1), .B(n502), .ZN(n435) );
  XNOR2_X1 U854 ( .A(n502), .B(n468), .ZN(n429) );
  XNOR2_X1 U855 ( .A(n472), .B(n502), .ZN(n433) );
  XNOR2_X1 U856 ( .A(n502), .B(n465), .ZN(n426) );
  XNOR2_X1 U857 ( .A(n473), .B(n502), .ZN(n434) );
  XNOR2_X1 U858 ( .A(n470), .B(n502), .ZN(n431) );
  INV_X1 U859 ( .A(n502), .ZN(n496) );
  XNOR2_X1 U860 ( .A(n502), .B(n471), .ZN(n432) );
  XNOR2_X1 U861 ( .A(n502), .B(b[8]), .ZN(n427) );
  XNOR2_X1 U862 ( .A(n502), .B(n467), .ZN(n428) );
  XNOR2_X1 U863 ( .A(n503), .B(n467), .ZN(n441) );
  XNOR2_X1 U864 ( .A(n470), .B(n503), .ZN(n444) );
  XNOR2_X1 U865 ( .A(n1), .B(n503), .ZN(n448) );
  XNOR2_X1 U866 ( .A(n469), .B(n503), .ZN(n443) );
  XNOR2_X1 U867 ( .A(n464), .B(n503), .ZN(n438) );
  XNOR2_X1 U868 ( .A(n473), .B(n503), .ZN(n447) );
  XNOR2_X1 U869 ( .A(n503), .B(n468), .ZN(n442) );
  XNOR2_X1 U870 ( .A(n463), .B(n503), .ZN(n437) );
  INV_X1 U871 ( .A(n503), .ZN(n497) );
  XNOR2_X1 U872 ( .A(n503), .B(n465), .ZN(n439) );
  XNOR2_X1 U873 ( .A(n503), .B(b[8]), .ZN(n440) );
  XNOR2_X1 U874 ( .A(n472), .B(n503), .ZN(n446) );
  XNOR2_X1 U875 ( .A(n471), .B(n503), .ZN(n445) );
  OAI22_X1 U876 ( .A1(n510), .A2(n498), .B1(n462), .B2(n516), .ZN(n312) );
  INV_X1 U877 ( .A(n504), .ZN(n498) );
  AND2_X1 U878 ( .A1(n1), .A2(n305), .ZN(product[0]) );
  INV_X1 U879 ( .A(n516), .ZN(n305) );
  XNOR2_X1 U880 ( .A(n24), .B(n154), .ZN(product[2]) );
  NAND2_X1 U881 ( .A1(n599), .A2(n153), .ZN(n24) );
  XOR2_X1 U882 ( .A(n22), .B(n145), .Z(product[4]) );
  NAND2_X1 U883 ( .A1(n175), .A2(n144), .ZN(n22) );
  XOR2_X1 U884 ( .A(n23), .B(n149), .Z(product[3]) );
  NAND2_X1 U885 ( .A1(n176), .A2(n148), .ZN(n23) );
  XNOR2_X1 U886 ( .A(n21), .B(n142), .ZN(product[5]) );
  NAND2_X1 U887 ( .A1(n601), .A2(n141), .ZN(n21) );
  XOR2_X1 U888 ( .A(n580), .B(n17), .Z(product[9]) );
  NAND2_X1 U889 ( .A1(n172), .A2(n132), .ZN(n19) );
  INV_X1 U890 ( .A(n134), .ZN(n133) );
  XNOR2_X1 U891 ( .A(n130), .B(n18), .ZN(product[8]) );
  OAI21_X1 U892 ( .B1(n133), .B2(n131), .A(n132), .ZN(n130) );
  XOR2_X1 U893 ( .A(n121), .B(n16), .Z(product[10]) );
  INV_X1 U894 ( .A(n122), .ZN(n121) );
  XNOR2_X1 U895 ( .A(n118), .B(n15), .ZN(product[11]) );
  OAI21_X1 U896 ( .B1(n121), .B2(n119), .A(n120), .ZN(n118) );
  XNOR2_X1 U897 ( .A(n112), .B(n14), .ZN(product[12]) );
  INV_X1 U898 ( .A(n113), .ZN(n112) );
  XOR2_X1 U899 ( .A(n98), .B(n12), .Z(product[14]) );
  AOI21_X1 U900 ( .B1(n112), .B2(n99), .A(n100), .ZN(n98) );
  XOR2_X1 U901 ( .A(n107), .B(n13), .Z(product[13]) );
  AOI21_X1 U902 ( .B1(n112), .B2(n108), .A(n109), .ZN(n107) );
  AOI21_X1 U903 ( .B1(n92), .B2(n112), .A(n93), .ZN(n91) );
  INV_X1 U904 ( .A(n596), .ZN(n83) );
  AOI21_X1 U905 ( .B1(n593), .B2(n39), .A(n40), .ZN(n38) );
  AOI21_X1 U906 ( .B1(n574), .B2(n27), .A(n28), .ZN(n26) );
  XNOR2_X1 U907 ( .A(n31), .B(n4), .ZN(product[22]) );
  OAI21_X1 U908 ( .B1(n584), .B2(n32), .A(n33), .ZN(n31) );
  AOI21_X1 U909 ( .B1(n593), .B2(n61), .A(n62), .ZN(n60) );
  AOI21_X1 U910 ( .B1(n593), .B2(n52), .A(n53), .ZN(n51) );
  XOR2_X1 U911 ( .A(n78), .B(n9), .Z(product[17]) );
  AOI21_X1 U912 ( .B1(n596), .B2(n163), .A(n80), .ZN(n78) );
  XNOR2_X1 U913 ( .A(n71), .B(n8), .ZN(product[18]) );
  OAI21_X1 U914 ( .B1(n78), .B2(n76), .A(n77), .ZN(n71) );
endmodule


module datapath_DW01_add_16 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n39, n40, n41, n42, n44, n45, n46, n47, n48,
         n52, n53, n54, n55, n56, n57, n59, n61, n62, n65, n66, n67, n68, n69,
         n70, n72, n73, n74, n75, n76, n80, n81, n82, n85, n87, n88, n89, n90,
         n91, n93, n95, n96, n98, n100, n101, n102, n104, n106, n107, n108,
         n109, n110, n112, n114, n115, n116, n117, n118, n120, n122, n123,
         n124, n125, n126, n128, n130, n131, n132, n133, n134, n136, n138,
         n139, n140, n142, n144, n145, n146, n148, n150, n151, n152, n153,
         n155, n158, n162, n168, n170, n172, n174, n178, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n291, n292;

  NOR2_X1 U207 ( .A1(n260), .A2(n40), .ZN(n258) );
  AND2_X1 U208 ( .A1(B[20]), .A2(A[20]), .ZN(n259) );
  INV_X4 U209 ( .A(n259), .ZN(n52) );
  INV_X1 U210 ( .A(n263), .ZN(n80) );
  NOR2_X1 U211 ( .A1(B[22]), .A2(A[22]), .ZN(n260) );
  AOI21_X1 U212 ( .B1(n277), .B2(n85), .A(n263), .ZN(n261) );
  AOI21_X1 U213 ( .B1(n277), .B2(n85), .A(n263), .ZN(n76) );
  AOI21_X1 U214 ( .B1(n107), .B2(n278), .A(n104), .ZN(n262) );
  AOI21_X1 U215 ( .B1(n107), .B2(n278), .A(n104), .ZN(n102) );
  OR2_X2 U216 ( .A1(B[16]), .A2(A[16]), .ZN(n277) );
  AND2_X1 U217 ( .A1(B[16]), .A2(A[16]), .ZN(n263) );
  OR2_X1 U218 ( .A1(B[22]), .A2(A[22]), .ZN(n264) );
  CLKBUF_X1 U219 ( .A(n107), .Z(n265) );
  CLKBUF_X1 U220 ( .A(n115), .Z(n266) );
  OR2_X1 U221 ( .A1(n67), .A2(n47), .ZN(n267) );
  OAI21_X1 U222 ( .B1(n261), .B2(n72), .A(n73), .ZN(n268) );
  OAI21_X1 U223 ( .B1(n76), .B2(n72), .A(n73), .ZN(n269) );
  AOI21_X1 U224 ( .B1(n288), .B2(n123), .A(n120), .ZN(n270) );
  CLKBUF_X1 U225 ( .A(n110), .Z(n271) );
  OAI21_X1 U226 ( .B1(n90), .B2(n102), .A(n91), .ZN(n272) );
  CLKBUF_X1 U227 ( .A(n123), .Z(n273) );
  CLKBUF_X1 U228 ( .A(n126), .Z(n274) );
  AOI21_X1 U229 ( .B1(n272), .B2(n70), .A(n269), .ZN(n275) );
  AOI21_X1 U230 ( .B1(n70), .B2(n89), .A(n269), .ZN(n276) );
  AOI21_X1 U231 ( .B1(n70), .B2(n272), .A(n268), .ZN(n69) );
  OR2_X1 U232 ( .A1(B[12]), .A2(A[12]), .ZN(n278) );
  OR2_X1 U233 ( .A1(B[15]), .A2(A[15]), .ZN(n279) );
  OR2_X1 U234 ( .A1(B[13]), .A2(A[13]), .ZN(n280) );
  OR2_X1 U235 ( .A1(B[20]), .A2(A[20]), .ZN(n281) );
  OR2_X1 U236 ( .A1(B[19]), .A2(A[19]), .ZN(n282) );
  OR2_X1 U237 ( .A1(B[14]), .A2(A[14]), .ZN(n283) );
  OR2_X1 U238 ( .A1(B[10]), .A2(A[10]), .ZN(n284) );
  OR2_X1 U239 ( .A1(B[6]), .A2(A[6]), .ZN(n285) );
  OR2_X1 U240 ( .A1(B[4]), .A2(A[4]), .ZN(n286) );
  OR2_X1 U241 ( .A1(B[3]), .A2(A[3]), .ZN(n287) );
  OR2_X1 U242 ( .A1(B[8]), .A2(A[8]), .ZN(n288) );
  OR2_X1 U243 ( .A1(B[2]), .A2(A[2]), .ZN(n289) );
  AND2_X1 U244 ( .A1(n292), .A2(n155), .ZN(SUM[0]) );
  OR2_X1 U245 ( .A1(B[23]), .A2(A[23]), .ZN(n291) );
  OR2_X1 U246 ( .A1(B[0]), .A2(A[0]), .ZN(n292) );
  NAND2_X1 U247 ( .A1(B[0]), .A2(A[0]), .ZN(n155) );
  NAND2_X1 U248 ( .A1(B[23]), .A2(A[23]), .ZN(n27) );
  NOR2_X1 U249 ( .A1(B[21]), .A2(A[21]), .ZN(n40) );
  NAND2_X1 U250 ( .A1(n291), .A2(n27), .ZN(n2) );
  NAND2_X1 U251 ( .A1(n158), .A2(n41), .ZN(n4) );
  INV_X1 U252 ( .A(n41), .ZN(n39) );
  NAND2_X1 U253 ( .A1(B[21]), .A2(A[21]), .ZN(n41) );
  NAND2_X1 U254 ( .A1(B[7]), .A2(A[7]), .ZN(n125) );
  NAND2_X1 U255 ( .A1(n162), .A2(n73), .ZN(n8) );
  NAND2_X1 U256 ( .A1(B[17]), .A2(A[17]), .ZN(n73) );
  NAND2_X1 U257 ( .A1(B[5]), .A2(A[5]), .ZN(n133) );
  NAND2_X1 U258 ( .A1(B[1]), .A2(A[1]), .ZN(n153) );
  NAND2_X1 U259 ( .A1(n264), .A2(n34), .ZN(n3) );
  NAND2_X1 U260 ( .A1(B[2]), .A2(A[2]), .ZN(n150) );
  NAND2_X1 U261 ( .A1(n168), .A2(n109), .ZN(n14) );
  NAND2_X1 U262 ( .A1(B[11]), .A2(A[11]), .ZN(n109) );
  NAND2_X1 U263 ( .A1(n283), .A2(n95), .ZN(n11) );
  INV_X1 U264 ( .A(n279), .ZN(n82) );
  AOI21_X1 U265 ( .B1(n286), .B2(n139), .A(n136), .ZN(n134) );
  NAND2_X1 U266 ( .A1(n65), .A2(n68), .ZN(n7) );
  INV_X1 U267 ( .A(n68), .ZN(n66) );
  NAND2_X1 U268 ( .A1(B[18]), .A2(A[18]), .ZN(n68) );
  NAND2_X1 U269 ( .A1(B[22]), .A2(A[22]), .ZN(n34) );
  NAND2_X1 U270 ( .A1(B[9]), .A2(A[9]), .ZN(n117) );
  NAND2_X1 U271 ( .A1(n281), .A2(n52), .ZN(n5) );
  NAND2_X1 U272 ( .A1(n280), .A2(n100), .ZN(n12) );
  INV_X1 U273 ( .A(n57), .ZN(n56) );
  NAND2_X1 U274 ( .A1(n279), .A2(n87), .ZN(n10) );
  NAND2_X1 U275 ( .A1(B[3]), .A2(A[3]), .ZN(n144) );
  INV_X1 U276 ( .A(n124), .ZN(n172) );
  OAI21_X1 U277 ( .B1(n126), .B2(n124), .A(n125), .ZN(n123) );
  NOR2_X1 U278 ( .A1(B[7]), .A2(A[7]), .ZN(n124) );
  NAND2_X1 U279 ( .A1(B[14]), .A2(A[14]), .ZN(n95) );
  NAND2_X1 U280 ( .A1(n277), .A2(n80), .ZN(n9) );
  NAND2_X1 U281 ( .A1(n278), .A2(n106), .ZN(n13) );
  INV_X1 U282 ( .A(n106), .ZN(n104) );
  NAND2_X1 U283 ( .A1(B[12]), .A2(A[12]), .ZN(n106) );
  INV_X1 U284 ( .A(n152), .ZN(n178) );
  NOR2_X1 U285 ( .A1(B[1]), .A2(A[1]), .ZN(n152) );
  INV_X1 U286 ( .A(n150), .ZN(n148) );
  NAND2_X1 U287 ( .A1(B[13]), .A2(A[13]), .ZN(n100) );
  NAND2_X1 U288 ( .A1(B[19]), .A2(A[19]), .ZN(n61) );
  INV_X1 U289 ( .A(n108), .ZN(n168) );
  NOR2_X1 U290 ( .A1(B[11]), .A2(A[11]), .ZN(n108) );
  INV_X1 U291 ( .A(n132), .ZN(n174) );
  NOR2_X1 U292 ( .A1(B[5]), .A2(A[5]), .ZN(n132) );
  NAND2_X1 U293 ( .A1(B[10]), .A2(A[10]), .ZN(n114) );
  NAND2_X1 U294 ( .A1(B[15]), .A2(A[15]), .ZN(n87) );
  NAND2_X1 U295 ( .A1(n282), .A2(n61), .ZN(n6) );
  INV_X1 U296 ( .A(n282), .ZN(n57) );
  INV_X1 U297 ( .A(n95), .ZN(n93) );
  INV_X1 U298 ( .A(n100), .ZN(n98) );
  OAI21_X1 U299 ( .B1(n152), .B2(n155), .A(n153), .ZN(n151) );
  INV_X1 U300 ( .A(n122), .ZN(n120) );
  NAND2_X1 U301 ( .A1(B[8]), .A2(A[8]), .ZN(n122) );
  INV_X1 U302 ( .A(n116), .ZN(n170) );
  NOR2_X1 U303 ( .A1(B[9]), .A2(A[9]), .ZN(n116) );
  INV_X1 U304 ( .A(n138), .ZN(n136) );
  NAND2_X1 U305 ( .A1(B[4]), .A2(A[4]), .ZN(n138) );
  INV_X1 U306 ( .A(n87), .ZN(n85) );
  INV_X1 U307 ( .A(n61), .ZN(n59) );
  INV_X1 U308 ( .A(n144), .ZN(n142) );
  AOI21_X1 U309 ( .B1(n289), .B2(n151), .A(n148), .ZN(n146) );
  INV_X1 U310 ( .A(n72), .ZN(n162) );
  NOR2_X1 U311 ( .A1(B[17]), .A2(A[17]), .ZN(n72) );
  INV_X1 U312 ( .A(n130), .ZN(n128) );
  NAND2_X1 U313 ( .A1(B[6]), .A2(A[6]), .ZN(n130) );
  OAI21_X1 U314 ( .B1(n118), .B2(n116), .A(n117), .ZN(n115) );
  INV_X1 U315 ( .A(n114), .ZN(n112) );
  AOI21_X1 U316 ( .B1(n288), .B2(n123), .A(n120), .ZN(n118) );
  AOI21_X1 U317 ( .B1(n284), .B2(n115), .A(n112), .ZN(n110) );
  OAI21_X1 U318 ( .B1(n110), .B2(n108), .A(n109), .ZN(n107) );
  INV_X1 U319 ( .A(n40), .ZN(n158) );
  OAI21_X1 U320 ( .B1(n47), .B2(n68), .A(n48), .ZN(n46) );
  AOI21_X1 U321 ( .B1(n281), .B2(n59), .A(n259), .ZN(n48) );
  AOI21_X1 U322 ( .B1(n283), .B2(n98), .A(n93), .ZN(n91) );
  NAND2_X1 U323 ( .A1(n277), .A2(n279), .ZN(n75) );
  OAI21_X1 U324 ( .B1(n90), .B2(n262), .A(n91), .ZN(n89) );
  NAND2_X1 U325 ( .A1(n283), .A2(n280), .ZN(n90) );
  INV_X1 U326 ( .A(n67), .ZN(n65) );
  NOR2_X1 U327 ( .A1(B[18]), .A2(A[18]), .ZN(n67) );
  NOR2_X1 U328 ( .A1(n75), .A2(n72), .ZN(n70) );
  NOR2_X1 U329 ( .A1(n67), .A2(n47), .ZN(n45) );
  NAND2_X1 U330 ( .A1(n282), .A2(n281), .ZN(n47) );
  NAND2_X1 U331 ( .A1(n65), .A2(n56), .ZN(n54) );
  AOI21_X1 U332 ( .B1(n66), .B2(n56), .A(n59), .ZN(n55) );
  OAI21_X1 U333 ( .B1(n33), .B2(n41), .A(n34), .ZN(n32) );
  NOR2_X1 U334 ( .A1(n260), .A2(n40), .ZN(n31) );
  NOR2_X1 U335 ( .A1(B[22]), .A2(A[22]), .ZN(n33) );
  INV_X1 U336 ( .A(n146), .ZN(n145) );
  AOI21_X1 U337 ( .B1(n46), .B2(n158), .A(n39), .ZN(n37) );
  INV_X1 U338 ( .A(n46), .ZN(n44) );
  AOI21_X1 U339 ( .B1(n46), .B2(n31), .A(n32), .ZN(n30) );
  AOI21_X1 U340 ( .B1(n285), .B2(n131), .A(n128), .ZN(n126) );
  OAI21_X1 U341 ( .B1(n134), .B2(n132), .A(n133), .ZN(n131) );
  NAND2_X1 U342 ( .A1(n258), .A2(n45), .ZN(n29) );
  NAND2_X1 U343 ( .A1(n45), .A2(n158), .ZN(n36) );
  INV_X1 U344 ( .A(n140), .ZN(n139) );
  AOI21_X1 U345 ( .B1(n287), .B2(n145), .A(n142), .ZN(n140) );
  XOR2_X1 U346 ( .A(n24), .B(n155), .Z(SUM[1]) );
  NAND2_X1 U347 ( .A1(n178), .A2(n153), .ZN(n24) );
  XNOR2_X1 U348 ( .A(n23), .B(n151), .ZN(SUM[2]) );
  NAND2_X1 U349 ( .A1(n289), .A2(n150), .ZN(n23) );
  XNOR2_X1 U350 ( .A(n22), .B(n145), .ZN(SUM[3]) );
  NAND2_X1 U351 ( .A1(n287), .A2(n144), .ZN(n22) );
  XNOR2_X1 U352 ( .A(n21), .B(n139), .ZN(SUM[4]) );
  NAND2_X1 U353 ( .A1(n286), .A2(n138), .ZN(n21) );
  XOR2_X1 U354 ( .A(n20), .B(n134), .Z(SUM[5]) );
  NAND2_X1 U355 ( .A1(n174), .A2(n133), .ZN(n20) );
  XOR2_X1 U356 ( .A(n18), .B(n274), .Z(SUM[7]) );
  NAND2_X1 U357 ( .A1(n172), .A2(n125), .ZN(n18) );
  XNOR2_X1 U358 ( .A(n19), .B(n131), .ZN(SUM[6]) );
  NAND2_X1 U359 ( .A1(n285), .A2(n130), .ZN(n19) );
  XNOR2_X1 U360 ( .A(n17), .B(n273), .ZN(SUM[8]) );
  NAND2_X1 U361 ( .A1(n288), .A2(n122), .ZN(n17) );
  XOR2_X1 U362 ( .A(n16), .B(n270), .Z(SUM[9]) );
  NAND2_X1 U363 ( .A1(n170), .A2(n117), .ZN(n16) );
  NAND2_X1 U364 ( .A1(n284), .A2(n114), .ZN(n15) );
  XNOR2_X1 U365 ( .A(n15), .B(n266), .ZN(SUM[10]) );
  XOR2_X1 U366 ( .A(n14), .B(n271), .Z(SUM[11]) );
  XNOR2_X1 U367 ( .A(n13), .B(n265), .ZN(SUM[12]) );
  XNOR2_X1 U368 ( .A(n12), .B(n101), .ZN(SUM[13]) );
  INV_X1 U369 ( .A(n262), .ZN(n101) );
  XOR2_X1 U370 ( .A(n96), .B(n11), .Z(SUM[14]) );
  AOI21_X1 U371 ( .B1(n101), .B2(n280), .A(n98), .ZN(n96) );
  XOR2_X1 U372 ( .A(n88), .B(n10), .Z(SUM[15]) );
  INV_X1 U373 ( .A(n89), .ZN(n88) );
  XNOR2_X1 U374 ( .A(n74), .B(n8), .ZN(SUM[17]) );
  OAI21_X1 U375 ( .B1(n88), .B2(n75), .A(n261), .ZN(n74) );
  XNOR2_X1 U376 ( .A(n81), .B(n9), .ZN(SUM[16]) );
  OAI21_X1 U377 ( .B1(n88), .B2(n82), .A(n87), .ZN(n81) );
  XOR2_X1 U378 ( .A(n275), .B(n7), .Z(SUM[18]) );
  XNOR2_X1 U379 ( .A(n62), .B(n6), .ZN(SUM[19]) );
  OAI21_X1 U380 ( .B1(n276), .B2(n67), .A(n68), .ZN(n62) );
  XNOR2_X1 U381 ( .A(n42), .B(n4), .ZN(SUM[21]) );
  OAI21_X1 U382 ( .B1(n276), .B2(n267), .A(n44), .ZN(n42) );
  XNOR2_X1 U383 ( .A(n35), .B(n3), .ZN(SUM[22]) );
  OAI21_X1 U384 ( .B1(n69), .B2(n36), .A(n37), .ZN(n35) );
  XNOR2_X1 U385 ( .A(n53), .B(n5), .ZN(SUM[20]) );
  OAI21_X1 U386 ( .B1(n275), .B2(n54), .A(n55), .ZN(n53) );
  XNOR2_X1 U387 ( .A(n28), .B(n2), .ZN(SUM[23]) );
  OAI21_X1 U388 ( .B1(n29), .B2(n69), .A(n30), .ZN(n28) );
endmodule


module datapath_DW01_add_17 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n26, n27, n29, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n44, n45, n46, n47, n48, n49, n51, n53,
         n54, n57, n58, n59, n60, n64, n65, n66, n69, n71, n72, n73, n74, n75,
         n77, n79, n80, n82, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n99, n101, n102, n104, n106, n107, n108, n110,
         n112, n113, n114, n115, n116, n118, n120, n121, n122, n123, n124,
         n126, n128, n129, n130, n131, n132, n134, n136, n137, n138, n139,
         n140, n141, n142, n144, n146, n147, n154, n155, n159, n163, n165,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272;

  FA_X1 U181 ( .A(B[2]), .B(A[2]), .CI(n141), .CO(n140), .S(SUM[2]) );
  FA_X1 U182 ( .A(n142), .B(A[1]), .CI(B[1]), .CO(n141), .S(SUM[1]) );
  OR2_X2 U192 ( .A1(B[20]), .A2(A[20]), .ZN(n266) );
  AND2_X1 U193 ( .A1(B[18]), .A2(A[18]), .ZN(n252) );
  INV_X1 U194 ( .A(n250), .ZN(n44) );
  INV_X1 U195 ( .A(n252), .ZN(n64) );
  OR2_X1 U196 ( .A1(A[19]), .A2(B[19]), .ZN(n245) );
  OR2_X1 U197 ( .A1(B[7]), .A2(A[7]), .ZN(n246) );
  NOR2_X1 U198 ( .A1(B[14]), .A2(A[14]), .ZN(n247) );
  NOR2_X1 U199 ( .A1(B[14]), .A2(A[14]), .ZN(n89) );
  OR2_X1 U200 ( .A1(B[12]), .A2(A[12]), .ZN(n267) );
  CLKBUF_X1 U201 ( .A(n121), .Z(n248) );
  CLKBUF_X1 U202 ( .A(n124), .Z(n249) );
  AND2_X1 U203 ( .A1(B[20]), .A2(A[20]), .ZN(n250) );
  OR2_X2 U204 ( .A1(B[18]), .A2(A[18]), .ZN(n264) );
  AOI21_X1 U205 ( .B1(n113), .B2(n260), .A(n110), .ZN(n251) );
  AOI21_X1 U206 ( .B1(n95), .B2(n87), .A(n88), .ZN(n253) );
  AOI21_X1 U207 ( .B1(n87), .B2(n95), .A(n88), .ZN(n86) );
  OAI21_X2 U208 ( .B1(n116), .B2(n114), .A(n115), .ZN(n113) );
  OAI21_X1 U209 ( .B1(n253), .B2(n74), .A(n75), .ZN(n254) );
  AOI21_X1 U210 ( .B1(n254), .B2(n37), .A(n38), .ZN(n255) );
  AOI21_X1 U211 ( .B1(n73), .B2(n37), .A(n38), .ZN(n256) );
  AOI21_X1 U212 ( .B1(n254), .B2(n37), .A(n38), .ZN(n1) );
  AOI21_X1 U213 ( .B1(n264), .B2(n69), .A(n252), .ZN(n257) );
  OR2_X1 U214 ( .A1(n32), .A2(n35), .ZN(n258) );
  AND2_X1 U215 ( .A1(n272), .A2(n144), .ZN(SUM[0]) );
  NOR2_X1 U216 ( .A1(B[22]), .A2(A[22]), .ZN(n32) );
  OR2_X1 U217 ( .A1(B[10]), .A2(A[10]), .ZN(n260) );
  OR2_X1 U218 ( .A1(B[17]), .A2(A[17]), .ZN(n261) );
  OR2_X1 U219 ( .A1(B[15]), .A2(A[15]), .ZN(n262) );
  OR2_X1 U220 ( .A1(B[11]), .A2(A[11]), .ZN(n263) );
  OR2_X1 U221 ( .A1(B[16]), .A2(A[16]), .ZN(n265) );
  OR2_X1 U222 ( .A1(B[8]), .A2(A[8]), .ZN(n268) );
  OR2_X1 U223 ( .A1(B[6]), .A2(A[6]), .ZN(n269) );
  OR2_X1 U224 ( .A1(B[4]), .A2(A[4]), .ZN(n270) );
  OR2_X1 U225 ( .A1(B[23]), .A2(A[23]), .ZN(n271) );
  OR2_X1 U226 ( .A1(B[0]), .A2(A[0]), .ZN(n272) );
  INV_X1 U227 ( .A(n144), .ZN(n142) );
  NAND2_X1 U228 ( .A1(B[0]), .A2(A[0]), .ZN(n144) );
  NAND2_X1 U229 ( .A1(B[23]), .A2(A[23]), .ZN(n26) );
  NAND2_X1 U230 ( .A1(B[9]), .A2(A[9]), .ZN(n115) );
  NAND2_X1 U231 ( .A1(B[3]), .A2(A[3]), .ZN(n139) );
  NAND2_X1 U232 ( .A1(n147), .A2(n36), .ZN(n5) );
  NAND2_X1 U233 ( .A1(B[21]), .A2(A[21]), .ZN(n36) );
  NAND2_X1 U234 ( .A1(n271), .A2(n26), .ZN(n3) );
  INV_X1 U235 ( .A(n138), .ZN(n165) );
  NOR2_X1 U236 ( .A1(B[3]), .A2(A[3]), .ZN(n138) );
  NAND2_X1 U237 ( .A1(n262), .A2(n84), .ZN(n11) );
  NAND2_X1 U238 ( .A1(n154), .A2(n90), .ZN(n12) );
  NAND2_X1 U239 ( .A1(n146), .A2(n33), .ZN(n4) );
  NAND2_X1 U240 ( .A1(n155), .A2(n93), .ZN(n13) );
  INV_X1 U241 ( .A(n114), .ZN(n159) );
  NOR2_X1 U242 ( .A1(B[9]), .A2(A[9]), .ZN(n114) );
  NAND2_X1 U243 ( .A1(B[15]), .A2(A[15]), .ZN(n84) );
  NAND2_X1 U244 ( .A1(B[5]), .A2(A[5]), .ZN(n131) );
  INV_X1 U245 ( .A(n112), .ZN(n110) );
  NAND2_X1 U246 ( .A1(B[10]), .A2(A[10]), .ZN(n112) );
  NAND2_X1 U247 ( .A1(B[7]), .A2(A[7]), .ZN(n123) );
  NAND2_X1 U248 ( .A1(B[14]), .A2(A[14]), .ZN(n90) );
  AOI21_X1 U249 ( .B1(n270), .B2(n137), .A(n134), .ZN(n132) );
  OAI21_X1 U250 ( .B1(n138), .B2(n2), .A(n139), .ZN(n137) );
  NAND2_X1 U251 ( .A1(n267), .A2(n101), .ZN(n14) );
  INV_X1 U252 ( .A(n31), .ZN(n29) );
  INV_X1 U253 ( .A(n84), .ZN(n82) );
  INV_X1 U254 ( .A(n140), .ZN(n2) );
  NAND2_X1 U255 ( .A1(n265), .A2(n79), .ZN(n10) );
  NAND2_X1 U256 ( .A1(B[13]), .A2(A[13]), .ZN(n93) );
  NAND2_X1 U257 ( .A1(B[6]), .A2(A[6]), .ZN(n128) );
  INV_X1 U258 ( .A(n59), .ZN(n57) );
  INV_X1 U259 ( .A(n245), .ZN(n49) );
  NAND2_X1 U260 ( .A1(n245), .A2(n53), .ZN(n7) );
  NAND2_X1 U261 ( .A1(B[22]), .A2(A[22]), .ZN(n33) );
  NAND2_X1 U262 ( .A1(n263), .A2(n106), .ZN(n15) );
  INV_X1 U263 ( .A(n106), .ZN(n104) );
  NAND2_X1 U264 ( .A1(B[11]), .A2(A[11]), .ZN(n106) );
  AOI21_X1 U265 ( .B1(n264), .B2(n69), .A(n252), .ZN(n60) );
  NAND2_X1 U266 ( .A1(n266), .A2(n44), .ZN(n6) );
  NAND2_X1 U267 ( .A1(B[16]), .A2(A[16]), .ZN(n79) );
  NAND2_X1 U268 ( .A1(B[19]), .A2(A[19]), .ZN(n53) );
  INV_X1 U269 ( .A(n130), .ZN(n163) );
  NOR2_X1 U270 ( .A1(B[5]), .A2(A[5]), .ZN(n130) );
  NAND2_X1 U271 ( .A1(n261), .A2(n71), .ZN(n9) );
  NOR2_X1 U272 ( .A1(B[7]), .A2(A[7]), .ZN(n122) );
  INV_X1 U273 ( .A(n136), .ZN(n134) );
  NAND2_X1 U274 ( .A1(B[4]), .A2(A[4]), .ZN(n136) );
  INV_X1 U275 ( .A(n120), .ZN(n118) );
  NAND2_X1 U276 ( .A1(B[8]), .A2(A[8]), .ZN(n120) );
  NAND2_X1 U277 ( .A1(B[17]), .A2(A[17]), .ZN(n71) );
  NAND2_X1 U278 ( .A1(n264), .A2(n261), .ZN(n59) );
  INV_X1 U279 ( .A(n261), .ZN(n66) );
  INV_X1 U280 ( .A(n79), .ZN(n77) );
  INV_X1 U281 ( .A(n53), .ZN(n51) );
  INV_X1 U282 ( .A(n101), .ZN(n99) );
  NAND2_X1 U283 ( .A1(B[12]), .A2(A[12]), .ZN(n101) );
  INV_X1 U284 ( .A(n247), .ZN(n154) );
  OAI21_X1 U285 ( .B1(n89), .B2(n93), .A(n90), .ZN(n88) );
  OAI21_X1 U286 ( .B1(n130), .B2(n132), .A(n131), .ZN(n129) );
  INV_X1 U287 ( .A(n128), .ZN(n126) );
  NAND2_X1 U288 ( .A1(n264), .A2(n64), .ZN(n8) );
  INV_X1 U289 ( .A(n71), .ZN(n69) );
  INV_X1 U290 ( .A(n92), .ZN(n155) );
  NOR2_X1 U291 ( .A1(B[13]), .A2(A[13]), .ZN(n92) );
  NOR2_X1 U292 ( .A1(n247), .A2(n92), .ZN(n87) );
  INV_X1 U293 ( .A(n257), .ZN(n58) );
  OAI21_X1 U294 ( .B1(n122), .B2(n124), .A(n123), .ZN(n121) );
  AOI21_X1 U295 ( .B1(n269), .B2(n129), .A(n126), .ZN(n124) );
  NAND2_X1 U296 ( .A1(n267), .A2(n263), .ZN(n96) );
  INV_X1 U297 ( .A(n49), .ZN(n48) );
  NAND2_X1 U298 ( .A1(n265), .A2(n262), .ZN(n74) );
  AOI21_X1 U299 ( .B1(n265), .B2(n82), .A(n77), .ZN(n75) );
  NAND2_X1 U300 ( .A1(n57), .A2(n48), .ZN(n46) );
  AOI21_X1 U301 ( .B1(n58), .B2(n48), .A(n51), .ZN(n47) );
  INV_X1 U302 ( .A(n35), .ZN(n147) );
  NOR2_X1 U303 ( .A1(B[21]), .A2(A[21]), .ZN(n35) );
  AOI21_X1 U304 ( .B1(n113), .B2(n260), .A(n110), .ZN(n108) );
  NAND2_X1 U305 ( .A1(n266), .A2(n245), .ZN(n39) );
  AOI21_X1 U306 ( .B1(n266), .B2(n51), .A(n250), .ZN(n40) );
  OAI21_X1 U307 ( .B1(n96), .B2(n108), .A(n97), .ZN(n95) );
  AOI21_X1 U308 ( .B1(n267), .B2(n104), .A(n99), .ZN(n97) );
  NOR2_X1 U309 ( .A1(n39), .A2(n59), .ZN(n37) );
  INV_X1 U310 ( .A(n32), .ZN(n146) );
  OAI21_X1 U311 ( .B1(n32), .B2(n36), .A(n33), .ZN(n31) );
  OAI21_X1 U312 ( .B1(n86), .B2(n74), .A(n75), .ZN(n73) );
  OAI21_X1 U313 ( .B1(n39), .B2(n60), .A(n40), .ZN(n38) );
  XNOR2_X1 U314 ( .A(n23), .B(n140), .ZN(SUM[3]) );
  NAND2_X1 U315 ( .A1(n165), .A2(n139), .ZN(n23) );
  XNOR2_X1 U316 ( .A(n22), .B(n137), .ZN(SUM[4]) );
  NAND2_X1 U317 ( .A1(n270), .A2(n136), .ZN(n22) );
  XOR2_X1 U318 ( .A(n21), .B(n132), .Z(SUM[5]) );
  NAND2_X1 U319 ( .A1(n163), .A2(n131), .ZN(n21) );
  XNOR2_X1 U320 ( .A(n20), .B(n129), .ZN(SUM[6]) );
  NAND2_X1 U321 ( .A1(n269), .A2(n128), .ZN(n20) );
  XOR2_X1 U322 ( .A(n19), .B(n249), .Z(SUM[7]) );
  NAND2_X1 U323 ( .A1(n246), .A2(n123), .ZN(n19) );
  XNOR2_X1 U324 ( .A(n18), .B(n248), .ZN(SUM[8]) );
  NAND2_X1 U325 ( .A1(n268), .A2(n120), .ZN(n18) );
  NAND2_X1 U326 ( .A1(n159), .A2(n115), .ZN(n17) );
  XOR2_X1 U327 ( .A(n116), .B(n17), .Z(SUM[9]) );
  AOI21_X1 U328 ( .B1(n121), .B2(n268), .A(n118), .ZN(n116) );
  NAND2_X1 U329 ( .A1(n260), .A2(n112), .ZN(n16) );
  XNOR2_X1 U330 ( .A(n16), .B(n113), .ZN(SUM[10]) );
  XNOR2_X1 U331 ( .A(n15), .B(n107), .ZN(SUM[11]) );
  INV_X1 U332 ( .A(n251), .ZN(n107) );
  XOR2_X1 U333 ( .A(n14), .B(n102), .Z(SUM[12]) );
  AOI21_X1 U334 ( .B1(n107), .B2(n263), .A(n104), .ZN(n102) );
  XOR2_X1 U335 ( .A(n94), .B(n13), .Z(SUM[13]) );
  INV_X1 U336 ( .A(n95), .ZN(n94) );
  XNOR2_X1 U337 ( .A(n91), .B(n12), .ZN(SUM[14]) );
  OAI21_X1 U338 ( .B1(n94), .B2(n92), .A(n93), .ZN(n91) );
  XNOR2_X1 U339 ( .A(n85), .B(n11), .ZN(SUM[15]) );
  INV_X1 U340 ( .A(n253), .ZN(n85) );
  XOR2_X1 U341 ( .A(n80), .B(n10), .Z(SUM[16]) );
  AOI21_X1 U342 ( .B1(n85), .B2(n262), .A(n82), .ZN(n80) );
  XOR2_X1 U343 ( .A(n72), .B(n9), .Z(SUM[17]) );
  INV_X1 U344 ( .A(n73), .ZN(n72) );
  XOR2_X1 U345 ( .A(n1), .B(n5), .Z(SUM[21]) );
  XNOR2_X1 U346 ( .A(n54), .B(n7), .ZN(SUM[19]) );
  OAI21_X1 U347 ( .B1(n72), .B2(n59), .A(n257), .ZN(n54) );
  XNOR2_X1 U348 ( .A(n65), .B(n8), .ZN(SUM[18]) );
  OAI21_X1 U349 ( .B1(n72), .B2(n66), .A(n71), .ZN(n65) );
  XNOR2_X1 U350 ( .A(n45), .B(n6), .ZN(SUM[20]) );
  OAI21_X1 U351 ( .B1(n72), .B2(n46), .A(n47), .ZN(n45) );
  XNOR2_X1 U352 ( .A(n27), .B(n3), .ZN(SUM[23]) );
  OAI21_X1 U353 ( .B1(n255), .B2(n258), .A(n29), .ZN(n27) );
  XNOR2_X1 U354 ( .A(n34), .B(n4), .ZN(SUM[22]) );
  OAI21_X1 U355 ( .B1(n256), .B2(n35), .A(n36), .ZN(n34) );
endmodule


module datapath_DW01_add_18 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n58, n59, n60, n61, n67, n68,
         n69, n71, n72, n73, n74, n76, n78, n79, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n91, n93, n94, n96, n98, n99, n100, n102, n104, n105,
         n106, n107, n109, n111, n112, n114, n116, n117, n118, n120, n122,
         n123, n124, n125, n126, n128, n130, n131, n132, n134, n136, n137,
         n138, n139, n140, n142, n144, n145, n146, n148, n150, n151, n152,
         n154, n155, n157, n158, n159, n160, n164, n171, n174, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281;

  FA_X1 U192 ( .A(B[2]), .B(A[2]), .CI(n152), .CO(n151), .S(SUM[2]) );
  FA_X1 U193 ( .A(n155), .B(A[1]), .CI(B[1]), .CO(n152), .S(SUM[1]) );
  AOI21_X1 U203 ( .B1(n277), .B2(n145), .A(n142), .ZN(n140) );
  INV_X1 U204 ( .A(n263), .ZN(n67) );
  AND2_X1 U205 ( .A1(n280), .A2(n154), .ZN(SUM[0]) );
  INV_X1 U206 ( .A(n85), .ZN(n257) );
  AND2_X1 U207 ( .A1(B[17]), .A2(A[17]), .ZN(n263) );
  OR2_X1 U208 ( .A1(B[18]), .A2(A[18]), .ZN(n272) );
  AOI21_X1 U209 ( .B1(n268), .B2(n257), .A(n76), .ZN(n258) );
  CLKBUF_X1 U210 ( .A(n123), .Z(n259) );
  AOI21_X1 U211 ( .B1(n259), .B2(n275), .A(n120), .ZN(n260) );
  CLKBUF_X1 U212 ( .A(n126), .Z(n261) );
  OR2_X1 U213 ( .A1(B[16]), .A2(A[16]), .ZN(n268) );
  OR2_X2 U214 ( .A1(B[17]), .A2(A[17]), .ZN(n262) );
  NOR2_X2 U215 ( .A1(B[22]), .A2(A[22]), .ZN(n31) );
  CLKBUF_X1 U216 ( .A(n105), .Z(n264) );
  OAI21_X1 U217 ( .B1(n88), .B2(n100), .A(n89), .ZN(n265) );
  AOI21_X2 U218 ( .B1(n105), .B2(n269), .A(n102), .ZN(n100) );
  AOI21_X1 U219 ( .B1(n265), .B2(n51), .A(n52), .ZN(n266) );
  AOI21_X1 U220 ( .B1(n87), .B2(n51), .A(n52), .ZN(n267) );
  AOI21_X1 U221 ( .B1(n87), .B2(n51), .A(n52), .ZN(n50) );
  OR2_X1 U222 ( .A1(B[12]), .A2(A[12]), .ZN(n269) );
  OR2_X1 U223 ( .A1(B[13]), .A2(A[13]), .ZN(n270) );
  OR2_X1 U224 ( .A1(B[10]), .A2(A[10]), .ZN(n271) );
  OR2_X1 U225 ( .A1(B[14]), .A2(A[14]), .ZN(n273) );
  OR2_X1 U226 ( .A1(B[11]), .A2(A[11]), .ZN(n274) );
  OR2_X1 U227 ( .A1(B[9]), .A2(A[9]), .ZN(n275) );
  OR2_X1 U228 ( .A1(B[6]), .A2(A[6]), .ZN(n276) );
  OR2_X1 U229 ( .A1(B[4]), .A2(A[4]), .ZN(n277) );
  OR2_X1 U230 ( .A1(B[3]), .A2(A[3]), .ZN(n278) );
  OR2_X1 U231 ( .A1(B[7]), .A2(A[7]), .ZN(n279) );
  OR2_X1 U232 ( .A1(B[0]), .A2(A[0]), .ZN(n280) );
  OR2_X1 U233 ( .A1(B[23]), .A2(A[23]), .ZN(n281) );
  INV_X1 U234 ( .A(n154), .ZN(n155) );
  NAND2_X1 U235 ( .A1(B[0]), .A2(A[0]), .ZN(n154) );
  NAND2_X1 U236 ( .A1(B[23]), .A2(A[23]), .ZN(n25) );
  NAND2_X1 U237 ( .A1(n281), .A2(n25), .ZN(n2) );
  NAND2_X1 U238 ( .A1(n159), .A2(n46), .ZN(n5) );
  NAND2_X1 U239 ( .A1(n160), .A2(n49), .ZN(n6) );
  NAND2_X1 U240 ( .A1(B[8]), .A2(A[8]), .ZN(n125) );
  NAND2_X1 U241 ( .A1(B[3]), .A2(A[3]), .ZN(n150) );
  NOR2_X1 U242 ( .A1(B[20]), .A2(A[20]), .ZN(n45) );
  NAND2_X1 U243 ( .A1(B[9]), .A2(A[9]), .ZN(n122) );
  NAND2_X1 U244 ( .A1(n158), .A2(n39), .ZN(n4) );
  NAND2_X1 U245 ( .A1(B[21]), .A2(A[21]), .ZN(n39) );
  NAND2_X1 U246 ( .A1(B[20]), .A2(A[20]), .ZN(n46) );
  NAND2_X1 U247 ( .A1(n157), .A2(n32), .ZN(n3) );
  NAND2_X1 U248 ( .A1(B[19]), .A2(A[19]), .ZN(n49) );
  NAND2_X1 U249 ( .A1(n269), .A2(n104), .ZN(n13) );
  INV_X1 U250 ( .A(n39), .ZN(n37) );
  NAND2_X1 U251 ( .A1(B[5]), .A2(A[5]), .ZN(n139) );
  INV_X1 U252 ( .A(n150), .ZN(n148) );
  NOR2_X1 U253 ( .A1(n31), .A2(n38), .ZN(n29) );
  NAND2_X1 U254 ( .A1(n273), .A2(n93), .ZN(n11) );
  NAND2_X1 U255 ( .A1(n270), .A2(n98), .ZN(n12) );
  INV_X1 U256 ( .A(n83), .ZN(n81) );
  AOI21_X1 U257 ( .B1(n278), .B2(n151), .A(n148), .ZN(n146) );
  NAND2_X1 U258 ( .A1(B[4]), .A2(A[4]), .ZN(n144) );
  NAND2_X1 U259 ( .A1(B[22]), .A2(A[22]), .ZN(n32) );
  NAND2_X1 U260 ( .A1(n164), .A2(n85), .ZN(n10) );
  INV_X1 U261 ( .A(n124), .ZN(n171) );
  NOR2_X1 U262 ( .A1(B[8]), .A2(A[8]), .ZN(n124) );
  NAND2_X1 U263 ( .A1(B[6]), .A2(A[6]), .ZN(n136) );
  NAND2_X1 U264 ( .A1(B[14]), .A2(A[14]), .ZN(n93) );
  INV_X1 U265 ( .A(n122), .ZN(n120) );
  INV_X1 U266 ( .A(n43), .ZN(n41) );
  NAND2_X1 U267 ( .A1(n43), .A2(n158), .ZN(n34) );
  NAND2_X1 U268 ( .A1(n29), .A2(n43), .ZN(n27) );
  NOR2_X1 U269 ( .A1(n45), .A2(n48), .ZN(n43) );
  NAND2_X1 U270 ( .A1(B[13]), .A2(A[13]), .ZN(n98) );
  AOI21_X1 U271 ( .B1(n268), .B2(n83), .A(n76), .ZN(n74) );
  NAND2_X1 U272 ( .A1(n262), .A2(n67), .ZN(n8) );
  INV_X1 U273 ( .A(n146), .ZN(n145) );
  INV_X1 U274 ( .A(n44), .ZN(n42) );
  AOI21_X1 U275 ( .B1(n44), .B2(n158), .A(n37), .ZN(n35) );
  OAI21_X1 U276 ( .B1(n45), .B2(n49), .A(n46), .ZN(n44) );
  INV_X1 U277 ( .A(n138), .ZN(n174) );
  NOR2_X1 U278 ( .A1(B[5]), .A2(A[5]), .ZN(n138) );
  NAND2_X1 U279 ( .A1(n272), .A2(n262), .ZN(n53) );
  INV_X1 U280 ( .A(n73), .ZN(n71) );
  INV_X1 U281 ( .A(n74), .ZN(n72) );
  AOI21_X1 U282 ( .B1(n123), .B2(n275), .A(n120), .ZN(n118) );
  OAI21_X1 U283 ( .B1(n126), .B2(n124), .A(n125), .ZN(n123) );
  NAND2_X1 U284 ( .A1(n271), .A2(n116), .ZN(n15) );
  INV_X1 U285 ( .A(n116), .ZN(n114) );
  NAND2_X1 U286 ( .A1(B[10]), .A2(A[10]), .ZN(n116) );
  INV_X1 U287 ( .A(n93), .ZN(n91) );
  INV_X1 U288 ( .A(n98), .ZN(n96) );
  AOI21_X1 U289 ( .B1(n29), .B2(n44), .A(n30), .ZN(n28) );
  NAND2_X1 U290 ( .A1(B[15]), .A2(A[15]), .ZN(n85) );
  INV_X1 U291 ( .A(n104), .ZN(n102) );
  NAND2_X1 U292 ( .A1(B[12]), .A2(A[12]), .ZN(n104) );
  INV_X1 U293 ( .A(n144), .ZN(n142) );
  NAND2_X1 U294 ( .A1(n268), .A2(n78), .ZN(n9) );
  OAI21_X1 U295 ( .B1(n106), .B2(n118), .A(n107), .ZN(n105) );
  AOI21_X1 U296 ( .B1(n274), .B2(n114), .A(n109), .ZN(n107) );
  NAND2_X1 U297 ( .A1(n274), .A2(n271), .ZN(n106) );
  INV_X1 U298 ( .A(n130), .ZN(n128) );
  NAND2_X1 U299 ( .A1(B[7]), .A2(A[7]), .ZN(n130) );
  NAND2_X1 U300 ( .A1(B[16]), .A2(A[16]), .ZN(n78) );
  OAI21_X1 U301 ( .B1(n138), .B2(n140), .A(n139), .ZN(n137) );
  INV_X1 U302 ( .A(n136), .ZN(n134) );
  INV_X1 U303 ( .A(n84), .ZN(n164) );
  INV_X1 U304 ( .A(n84), .ZN(n82) );
  NOR2_X1 U305 ( .A1(A[15]), .A2(B[15]), .ZN(n84) );
  INV_X1 U306 ( .A(n78), .ZN(n76) );
  INV_X1 U307 ( .A(n85), .ZN(n83) );
  NAND2_X1 U308 ( .A1(n268), .A2(n82), .ZN(n73) );
  AOI21_X1 U309 ( .B1(n272), .B2(n263), .A(n56), .ZN(n54) );
  AOI21_X1 U310 ( .B1(n273), .B2(n96), .A(n91), .ZN(n89) );
  NAND2_X1 U311 ( .A1(n272), .A2(n58), .ZN(n7) );
  INV_X1 U312 ( .A(n58), .ZN(n56) );
  NAND2_X1 U313 ( .A1(B[18]), .A2(A[18]), .ZN(n58) );
  OAI21_X1 U314 ( .B1(n88), .B2(n100), .A(n89), .ZN(n87) );
  NAND2_X1 U315 ( .A1(n273), .A2(n270), .ZN(n88) );
  INV_X1 U316 ( .A(n45), .ZN(n159) );
  NAND2_X1 U317 ( .A1(n71), .A2(n262), .ZN(n60) );
  AOI21_X1 U318 ( .B1(n72), .B2(n262), .A(n263), .ZN(n61) );
  NAND2_X1 U319 ( .A1(n274), .A2(n111), .ZN(n14) );
  INV_X1 U320 ( .A(n111), .ZN(n109) );
  NAND2_X1 U321 ( .A1(B[11]), .A2(A[11]), .ZN(n111) );
  INV_X1 U322 ( .A(n71), .ZN(n69) );
  INV_X1 U323 ( .A(n38), .ZN(n158) );
  NOR2_X1 U324 ( .A1(B[21]), .A2(A[21]), .ZN(n38) );
  INV_X1 U325 ( .A(n48), .ZN(n160) );
  NOR2_X1 U326 ( .A1(B[19]), .A2(A[19]), .ZN(n48) );
  NOR2_X1 U327 ( .A1(n73), .A2(n53), .ZN(n51) );
  INV_X1 U328 ( .A(n31), .ZN(n157) );
  OAI21_X1 U329 ( .B1(n31), .B2(n39), .A(n32), .ZN(n30) );
  OAI21_X1 U330 ( .B1(n258), .B2(n53), .A(n54), .ZN(n52) );
  INV_X1 U331 ( .A(n132), .ZN(n131) );
  AOI21_X1 U332 ( .B1(n137), .B2(n276), .A(n134), .ZN(n132) );
  XNOR2_X1 U333 ( .A(n22), .B(n151), .ZN(SUM[3]) );
  NAND2_X1 U334 ( .A1(n278), .A2(n150), .ZN(n22) );
  XNOR2_X1 U335 ( .A(n21), .B(n145), .ZN(SUM[4]) );
  NAND2_X1 U336 ( .A1(n277), .A2(n144), .ZN(n21) );
  XOR2_X1 U337 ( .A(n20), .B(n140), .Z(SUM[5]) );
  NAND2_X1 U338 ( .A1(n174), .A2(n139), .ZN(n20) );
  XNOR2_X1 U339 ( .A(n19), .B(n137), .ZN(SUM[6]) );
  NAND2_X1 U340 ( .A1(n276), .A2(n136), .ZN(n19) );
  XNOR2_X1 U341 ( .A(n18), .B(n131), .ZN(SUM[7]) );
  NAND2_X1 U342 ( .A1(n279), .A2(n130), .ZN(n18) );
  AOI21_X1 U343 ( .B1(n279), .B2(n131), .A(n128), .ZN(n126) );
  XOR2_X1 U344 ( .A(n17), .B(n261), .Z(SUM[8]) );
  NAND2_X1 U345 ( .A1(n171), .A2(n125), .ZN(n17) );
  NAND2_X1 U346 ( .A1(n275), .A2(n122), .ZN(n16) );
  XNOR2_X1 U347 ( .A(n16), .B(n259), .ZN(SUM[9]) );
  XNOR2_X1 U348 ( .A(n15), .B(n117), .ZN(SUM[10]) );
  INV_X1 U349 ( .A(n260), .ZN(n117) );
  XNOR2_X1 U350 ( .A(n13), .B(n264), .ZN(SUM[12]) );
  XOR2_X1 U351 ( .A(n112), .B(n14), .Z(SUM[11]) );
  AOI21_X1 U352 ( .B1(n271), .B2(n117), .A(n114), .ZN(n112) );
  XNOR2_X1 U353 ( .A(n12), .B(n99), .ZN(SUM[13]) );
  INV_X1 U354 ( .A(n100), .ZN(n99) );
  XOR2_X1 U355 ( .A(n94), .B(n11), .Z(SUM[14]) );
  AOI21_X1 U356 ( .B1(n99), .B2(n270), .A(n96), .ZN(n94) );
  XOR2_X1 U357 ( .A(n86), .B(n10), .Z(SUM[15]) );
  INV_X1 U358 ( .A(n265), .ZN(n86) );
  XNOR2_X1 U359 ( .A(n68), .B(n8), .ZN(SUM[17]) );
  OAI21_X1 U360 ( .B1(n86), .B2(n69), .A(n74), .ZN(n68) );
  XNOR2_X1 U361 ( .A(n79), .B(n9), .ZN(SUM[16]) );
  OAI21_X1 U362 ( .B1(n86), .B2(n84), .A(n81), .ZN(n79) );
  XNOR2_X1 U363 ( .A(n59), .B(n7), .ZN(SUM[18]) );
  OAI21_X1 U364 ( .B1(n60), .B2(n86), .A(n61), .ZN(n59) );
  XOR2_X1 U365 ( .A(n266), .B(n6), .Z(SUM[19]) );
  XNOR2_X1 U366 ( .A(n40), .B(n4), .ZN(SUM[21]) );
  OAI21_X1 U367 ( .B1(n267), .B2(n41), .A(n42), .ZN(n40) );
  XNOR2_X1 U368 ( .A(n33), .B(n3), .ZN(SUM[22]) );
  OAI21_X1 U369 ( .B1(n50), .B2(n34), .A(n35), .ZN(n33) );
  XNOR2_X1 U370 ( .A(n26), .B(n2), .ZN(SUM[23]) );
  OAI21_X1 U371 ( .B1(n267), .B2(n27), .A(n28), .ZN(n26) );
  XNOR2_X1 U372 ( .A(n47), .B(n5), .ZN(SUM[20]) );
  OAI21_X1 U373 ( .B1(n50), .B2(n48), .A(n49), .ZN(n47) );
endmodule


module datapath_DW01_add_19 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n27, n28, n30, n32, n33, n34,
         n35, n36, n37, n41, n42, n43, n44, n46, n48, n49, n50, n51, n52, n54,
         n56, n57, n58, n59, n60, n61, n63, n65, n66, n69, n70, n71, n72, n74,
         n76, n77, n78, n79, n81, n83, n84, n85, n86, n87, n89, n91, n92, n94,
         n96, n97, n98, n100, n102, n103, n104, n105, n107, n109, n110, n112,
         n114, n115, n116, n118, n120, n121, n122, n123, n124, n126, n128,
         n129, n130, n131, n132, n134, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n146, n148, n149, n150, n152, n154, n155, n156,
         n157, n159, n161, n174, n176, n178, n179, n182, n262, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294;

  AND2_X1 U211 ( .A1(B[21]), .A2(A[21]), .ZN(n264) );
  INV_X1 U212 ( .A(n264), .ZN(n41) );
  OR2_X1 U213 ( .A1(B[18]), .A2(A[18]), .ZN(n262) );
  AND2_X1 U214 ( .A1(n293), .A2(n159), .ZN(SUM[0]) );
  OR2_X1 U215 ( .A1(B[19]), .A2(A[19]), .ZN(n280) );
  OAI21_X2 U216 ( .B1(n98), .B2(n86), .A(n87), .ZN(n85) );
  CLKBUF_X1 U217 ( .A(n129), .Z(n265) );
  OAI21_X1 U218 ( .B1(n132), .B2(n130), .A(n131), .ZN(n129) );
  AOI21_X1 U219 ( .B1(n280), .B2(n63), .A(n54), .ZN(n266) );
  AOI21_X1 U220 ( .B1(n81), .B2(n278), .A(n74), .ZN(n267) );
  AOI21_X1 U221 ( .B1(n81), .B2(n278), .A(n74), .ZN(n268) );
  AOI21_X1 U222 ( .B1(n81), .B2(n278), .A(n74), .ZN(n72) );
  AOI21_X1 U223 ( .B1(n283), .B2(n46), .A(n264), .ZN(n269) );
  CLKBUF_X1 U224 ( .A(n116), .Z(n270) );
  OAI21_X1 U225 ( .B1(n267), .B2(n51), .A(n266), .ZN(n271) );
  CLKBUF_X1 U226 ( .A(n103), .Z(n272) );
  CLKBUF_X1 U227 ( .A(n132), .Z(n273) );
  AOI21_X1 U228 ( .B1(n265), .B2(n288), .A(n126), .ZN(n274) );
  AOI21_X1 U229 ( .B1(n272), .B2(n287), .A(n100), .ZN(n275) );
  OR2_X1 U230 ( .A1(B[12]), .A2(A[12]), .ZN(n282) );
  AOI21_X1 U231 ( .B1(n85), .B2(n49), .A(n50), .ZN(n276) );
  AOI21_X1 U232 ( .B1(n85), .B2(n49), .A(n271), .ZN(n1) );
  OR2_X1 U233 ( .A1(n33), .A2(n36), .ZN(n277) );
  OR2_X2 U234 ( .A1(B[17]), .A2(A[17]), .ZN(n278) );
  OR2_X1 U235 ( .A1(B[16]), .A2(A[16]), .ZN(n279) );
  OR2_X1 U236 ( .A1(B[15]), .A2(A[15]), .ZN(n281) );
  OR2_X1 U237 ( .A1(B[21]), .A2(A[21]), .ZN(n283) );
  OR2_X1 U238 ( .A1(B[20]), .A2(A[20]), .ZN(n284) );
  OR2_X1 U239 ( .A1(B[14]), .A2(A[14]), .ZN(n285) );
  OR2_X1 U240 ( .A1(B[11]), .A2(A[11]), .ZN(n286) );
  OR2_X1 U241 ( .A1(B[13]), .A2(A[13]), .ZN(n287) );
  OR2_X1 U242 ( .A1(B[8]), .A2(A[8]), .ZN(n288) );
  OR2_X1 U243 ( .A1(B[10]), .A2(A[10]), .ZN(n289) );
  OR2_X1 U244 ( .A1(B[6]), .A2(A[6]), .ZN(n290) );
  OR2_X1 U245 ( .A1(B[3]), .A2(A[3]), .ZN(n291) );
  OR2_X1 U246 ( .A1(B[2]), .A2(A[2]), .ZN(n292) );
  OR2_X1 U247 ( .A1(B[0]), .A2(A[0]), .ZN(n293) );
  OR2_X1 U248 ( .A1(B[23]), .A2(A[23]), .ZN(n294) );
  NAND2_X1 U249 ( .A1(B[0]), .A2(A[0]), .ZN(n159) );
  NAND2_X1 U250 ( .A1(B[23]), .A2(A[23]), .ZN(n27) );
  NAND2_X1 U251 ( .A1(n294), .A2(n27), .ZN(n2) );
  NAND2_X1 U252 ( .A1(n161), .A2(n34), .ZN(n3) );
  INV_X1 U253 ( .A(n61), .ZN(n60) );
  INV_X1 U254 ( .A(n284), .ZN(n43) );
  NAND2_X1 U255 ( .A1(B[1]), .A2(A[1]), .ZN(n157) );
  NAND2_X1 U256 ( .A1(B[22]), .A2(A[22]), .ZN(n34) );
  NAND2_X1 U257 ( .A1(n174), .A2(n123), .ZN(n16) );
  NAND2_X1 U258 ( .A1(B[9]), .A2(A[9]), .ZN(n123) );
  NAND2_X1 U259 ( .A1(B[2]), .A2(A[2]), .ZN(n154) );
  NAND2_X1 U260 ( .A1(B[5]), .A2(A[5]), .ZN(n139) );
  NAND2_X1 U261 ( .A1(B[4]), .A2(A[4]), .ZN(n143) );
  INV_X1 U262 ( .A(n71), .ZN(n69) );
  NAND2_X1 U263 ( .A1(B[3]), .A2(A[3]), .ZN(n148) );
  INV_X1 U264 ( .A(n262), .ZN(n61) );
  NAND2_X1 U265 ( .A1(n262), .A2(n65), .ZN(n7) );
  INV_X1 U266 ( .A(n279), .ZN(n78) );
  NAND2_X1 U267 ( .A1(n286), .A2(n114), .ZN(n14) );
  NAND2_X1 U268 ( .A1(n280), .A2(n56), .ZN(n6) );
  NAND2_X1 U269 ( .A1(B[7]), .A2(A[7]), .ZN(n131) );
  INV_X1 U270 ( .A(n32), .ZN(n30) );
  INV_X1 U271 ( .A(n81), .ZN(n79) );
  INV_X1 U272 ( .A(n46), .ZN(n44) );
  NAND2_X1 U273 ( .A1(n283), .A2(n41), .ZN(n4) );
  NAND2_X1 U274 ( .A1(B[18]), .A2(A[18]), .ZN(n65) );
  INV_X1 U275 ( .A(n156), .ZN(n182) );
  NOR2_X1 U276 ( .A1(B[1]), .A2(A[1]), .ZN(n156) );
  INV_X1 U277 ( .A(n154), .ZN(n152) );
  NAND2_X1 U278 ( .A1(B[6]), .A2(A[6]), .ZN(n136) );
  NAND2_X1 U279 ( .A1(B[19]), .A2(A[19]), .ZN(n56) );
  NAND2_X1 U280 ( .A1(B[11]), .A2(A[11]), .ZN(n114) );
  INV_X1 U281 ( .A(n122), .ZN(n174) );
  NOR2_X1 U282 ( .A1(B[9]), .A2(A[9]), .ZN(n122) );
  NAND2_X1 U283 ( .A1(n284), .A2(n48), .ZN(n5) );
  AOI21_X1 U284 ( .B1(n281), .B2(n94), .A(n89), .ZN(n87) );
  NAND2_X1 U285 ( .A1(n285), .A2(n281), .ZN(n86) );
  INV_X1 U286 ( .A(n268), .ZN(n70) );
  INV_X1 U287 ( .A(n142), .ZN(n179) );
  NOR2_X1 U288 ( .A1(B[4]), .A2(A[4]), .ZN(n142) );
  INV_X1 U289 ( .A(n138), .ZN(n178) );
  NOR2_X1 U290 ( .A1(B[5]), .A2(A[5]), .ZN(n138) );
  INV_X1 U291 ( .A(n128), .ZN(n126) );
  NAND2_X1 U292 ( .A1(B[8]), .A2(A[8]), .ZN(n128) );
  OAI21_X1 U293 ( .B1(n156), .B2(n159), .A(n157), .ZN(n155) );
  INV_X1 U294 ( .A(n148), .ZN(n146) );
  NAND2_X1 U295 ( .A1(n287), .A2(n102), .ZN(n12) );
  INV_X1 U296 ( .A(n102), .ZN(n100) );
  NAND2_X1 U297 ( .A1(B[13]), .A2(A[13]), .ZN(n102) );
  NAND2_X1 U298 ( .A1(B[20]), .A2(A[20]), .ZN(n48) );
  INV_X1 U299 ( .A(n56), .ZN(n54) );
  INV_X1 U300 ( .A(n65), .ZN(n63) );
  NAND2_X1 U301 ( .A1(n281), .A2(n91), .ZN(n10) );
  INV_X1 U302 ( .A(n91), .ZN(n89) );
  NAND2_X1 U303 ( .A1(B[15]), .A2(A[15]), .ZN(n91) );
  AOI21_X1 U304 ( .B1(n291), .B2(n149), .A(n146), .ZN(n144) );
  INV_X1 U305 ( .A(n136), .ZN(n134) );
  INV_X1 U306 ( .A(n114), .ZN(n112) );
  NAND2_X1 U307 ( .A1(n285), .A2(n96), .ZN(n11) );
  INV_X1 U308 ( .A(n96), .ZN(n94) );
  NAND2_X1 U309 ( .A1(B[14]), .A2(A[14]), .ZN(n96) );
  INV_X1 U310 ( .A(n48), .ZN(n46) );
  NAND2_X1 U311 ( .A1(n289), .A2(n120), .ZN(n15) );
  INV_X1 U312 ( .A(n120), .ZN(n118) );
  NAND2_X1 U313 ( .A1(B[10]), .A2(A[10]), .ZN(n120) );
  AOI21_X1 U314 ( .B1(n129), .B2(n288), .A(n126), .ZN(n124) );
  INV_X1 U315 ( .A(n130), .ZN(n176) );
  NOR2_X1 U316 ( .A1(B[7]), .A2(A[7]), .ZN(n130) );
  NAND2_X1 U317 ( .A1(n279), .A2(n83), .ZN(n9) );
  INV_X1 U318 ( .A(n83), .ZN(n81) );
  NAND2_X1 U319 ( .A1(B[16]), .A2(A[16]), .ZN(n83) );
  NAND2_X1 U320 ( .A1(n278), .A2(n76), .ZN(n8) );
  INV_X1 U321 ( .A(n76), .ZN(n74) );
  NAND2_X1 U322 ( .A1(B[17]), .A2(A[17]), .ZN(n76) );
  AOI21_X1 U323 ( .B1(n290), .B2(n137), .A(n134), .ZN(n132) );
  OAI21_X1 U324 ( .B1(n138), .B2(n140), .A(n139), .ZN(n137) );
  AOI21_X1 U325 ( .B1(n282), .B2(n112), .A(n107), .ZN(n105) );
  NAND2_X1 U326 ( .A1(n282), .A2(n109), .ZN(n13) );
  INV_X1 U327 ( .A(n109), .ZN(n107) );
  NAND2_X1 U328 ( .A1(B[12]), .A2(A[12]), .ZN(n109) );
  OAI21_X1 U329 ( .B1(n122), .B2(n124), .A(n123), .ZN(n121) );
  NAND2_X1 U330 ( .A1(n286), .A2(n282), .ZN(n104) );
  NAND2_X1 U331 ( .A1(n262), .A2(n280), .ZN(n51) );
  AOI21_X1 U332 ( .B1(n280), .B2(n63), .A(n54), .ZN(n52) );
  NAND2_X1 U333 ( .A1(n278), .A2(n279), .ZN(n71) );
  NAND2_X1 U334 ( .A1(n284), .A2(n283), .ZN(n36) );
  AOI21_X1 U335 ( .B1(n289), .B2(n121), .A(n118), .ZN(n116) );
  AOI21_X1 U336 ( .B1(n283), .B2(n46), .A(n264), .ZN(n37) );
  AOI21_X1 U337 ( .B1(n103), .B2(n287), .A(n100), .ZN(n98) );
  OAI21_X1 U338 ( .B1(n116), .B2(n104), .A(n105), .ZN(n103) );
  NAND2_X1 U339 ( .A1(n69), .A2(n60), .ZN(n58) );
  AOI21_X1 U340 ( .B1(n70), .B2(n60), .A(n63), .ZN(n59) );
  OAI21_X1 U341 ( .B1(n72), .B2(n51), .A(n52), .ZN(n50) );
  INV_X1 U342 ( .A(n33), .ZN(n161) );
  OAI21_X1 U343 ( .B1(n33), .B2(n37), .A(n34), .ZN(n32) );
  NOR2_X1 U344 ( .A1(B[22]), .A2(A[22]), .ZN(n33) );
  NOR2_X1 U345 ( .A1(n51), .A2(n71), .ZN(n49) );
  INV_X1 U346 ( .A(n141), .ZN(n140) );
  OAI21_X1 U347 ( .B1(n144), .B2(n142), .A(n143), .ZN(n141) );
  INV_X1 U348 ( .A(n150), .ZN(n149) );
  AOI21_X1 U349 ( .B1(n292), .B2(n155), .A(n152), .ZN(n150) );
  XOR2_X1 U350 ( .A(n24), .B(n159), .Z(SUM[1]) );
  NAND2_X1 U351 ( .A1(n182), .A2(n157), .ZN(n24) );
  XNOR2_X1 U352 ( .A(n23), .B(n155), .ZN(SUM[2]) );
  NAND2_X1 U353 ( .A1(n292), .A2(n154), .ZN(n23) );
  XNOR2_X1 U354 ( .A(n22), .B(n149), .ZN(SUM[3]) );
  NAND2_X1 U355 ( .A1(n291), .A2(n148), .ZN(n22) );
  XOR2_X1 U356 ( .A(n21), .B(n144), .Z(SUM[4]) );
  NAND2_X1 U357 ( .A1(n179), .A2(n143), .ZN(n21) );
  XOR2_X1 U358 ( .A(n20), .B(n140), .Z(SUM[5]) );
  NAND2_X1 U359 ( .A1(n178), .A2(n139), .ZN(n20) );
  XNOR2_X1 U360 ( .A(n19), .B(n137), .ZN(SUM[6]) );
  NAND2_X1 U361 ( .A1(n290), .A2(n136), .ZN(n19) );
  NAND2_X1 U362 ( .A1(n288), .A2(n128), .ZN(n17) );
  XOR2_X1 U363 ( .A(n18), .B(n273), .Z(SUM[7]) );
  NAND2_X1 U364 ( .A1(n176), .A2(n131), .ZN(n18) );
  XNOR2_X1 U365 ( .A(n17), .B(n265), .ZN(SUM[8]) );
  XOR2_X1 U366 ( .A(n16), .B(n274), .Z(SUM[9]) );
  XNOR2_X1 U367 ( .A(n15), .B(n121), .ZN(SUM[10]) );
  XNOR2_X1 U368 ( .A(n14), .B(n115), .ZN(SUM[11]) );
  INV_X1 U369 ( .A(n270), .ZN(n115) );
  XNOR2_X1 U370 ( .A(n12), .B(n272), .ZN(SUM[13]) );
  XOR2_X1 U371 ( .A(n110), .B(n13), .Z(SUM[12]) );
  AOI21_X1 U372 ( .B1(n286), .B2(n115), .A(n112), .ZN(n110) );
  XNOR2_X1 U373 ( .A(n97), .B(n11), .ZN(SUM[14]) );
  INV_X1 U374 ( .A(n275), .ZN(n97) );
  XOR2_X1 U375 ( .A(n92), .B(n10), .Z(SUM[15]) );
  AOI21_X1 U376 ( .B1(n97), .B2(n285), .A(n94), .ZN(n92) );
  XOR2_X1 U377 ( .A(n84), .B(n9), .Z(SUM[16]) );
  INV_X1 U378 ( .A(n85), .ZN(n84) );
  XOR2_X1 U379 ( .A(n276), .B(n5), .Z(SUM[20]) );
  XNOR2_X1 U380 ( .A(n66), .B(n7), .ZN(SUM[18]) );
  OAI21_X1 U381 ( .B1(n84), .B2(n71), .A(n268), .ZN(n66) );
  XNOR2_X1 U382 ( .A(n77), .B(n8), .ZN(SUM[17]) );
  OAI21_X1 U383 ( .B1(n84), .B2(n78), .A(n79), .ZN(n77) );
  XNOR2_X1 U384 ( .A(n57), .B(n6), .ZN(SUM[19]) );
  OAI21_X1 U385 ( .B1(n84), .B2(n58), .A(n59), .ZN(n57) );
  XNOR2_X1 U386 ( .A(n35), .B(n3), .ZN(SUM[22]) );
  OAI21_X1 U387 ( .B1(n1), .B2(n36), .A(n269), .ZN(n35) );
  XNOR2_X1 U388 ( .A(n42), .B(n4), .ZN(SUM[21]) );
  OAI21_X1 U389 ( .B1(n276), .B2(n43), .A(n44), .ZN(n42) );
  XNOR2_X1 U390 ( .A(n28), .B(n2), .ZN(SUM[23]) );
  OAI21_X1 U391 ( .B1(n1), .B2(n277), .A(n30), .ZN(n28) );
endmodule


module datapath_DW01_add_20 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n46, n47,
         n48, n49, n50, n57, n59, n60, n61, n62, n63, n65, n66, n67, n68, n69,
         n70, n71, n73, n74, n75, n77, n79, n80, n81, n82, n83, n84, n86, n87,
         n88, n89, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n104, n106, n107, n108, n109, n110, n112, n114, n115, n116,
         n117, n118, n120, n122, n123, n124, n125, n126, n128, n130, n131,
         n132, n134, n136, n137, n138, n139, n140, n141, n142, n143, n145,
         n147, n148, n149, n150, n152, n153, n154, n155, n156, n157, n158,
         n160, n162, n164, n167, n168, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n267, n268;

  AOI21_X2 U197 ( .B1(n91), .B2(n99), .A(n92), .ZN(n251) );
  NOR2_X2 U198 ( .A1(B[21]), .A2(A[21]), .ZN(n33) );
  CLKBUF_X1 U199 ( .A(n115), .Z(n248) );
  OAI21_X1 U200 ( .B1(n251), .B2(n62), .A(n63), .ZN(n249) );
  CLKBUF_X1 U201 ( .A(n93), .Z(n250) );
  CLKBUF_X1 U202 ( .A(n107), .Z(n252) );
  OR2_X1 U203 ( .A1(n87), .A2(n82), .ZN(n253) );
  NOR2_X1 U204 ( .A1(A[15]), .A2(B[15]), .ZN(n254) );
  INV_X1 U205 ( .A(n46), .ZN(n255) );
  CLKBUF_X1 U206 ( .A(n37), .Z(n256) );
  NOR2_X1 U207 ( .A1(A[20]), .A2(B[20]), .ZN(n257) );
  NOR2_X1 U208 ( .A1(n73), .A2(n66), .ZN(n258) );
  AOI21_X1 U209 ( .B1(n249), .B2(n31), .A(n32), .ZN(n259) );
  OR2_X1 U210 ( .A1(B[18]), .A2(A[18]), .ZN(n260) );
  OR2_X1 U211 ( .A1(B[10]), .A2(A[10]), .ZN(n261) );
  OR2_X1 U212 ( .A1(B[4]), .A2(A[4]), .ZN(n262) );
  OR2_X1 U213 ( .A1(B[6]), .A2(A[6]), .ZN(n263) );
  OR2_X1 U214 ( .A1(B[3]), .A2(A[3]), .ZN(n264) );
  OR2_X1 U215 ( .A1(B[8]), .A2(A[8]), .ZN(n265) );
  AND2_X1 U216 ( .A1(n268), .A2(n145), .ZN(SUM[0]) );
  OR2_X1 U217 ( .A1(B[23]), .A2(A[23]), .ZN(n267) );
  OR2_X1 U218 ( .A1(B[0]), .A2(A[0]), .ZN(n268) );
  NAND2_X1 U219 ( .A1(B[0]), .A2(A[0]), .ZN(n145) );
  NAND2_X1 U220 ( .A1(B[23]), .A2(A[23]), .ZN(n26) );
  NAND2_X1 U221 ( .A1(n158), .A2(n101), .ZN(n13) );
  NAND2_X1 U222 ( .A1(B[11]), .A2(A[11]), .ZN(n101) );
  NAND2_X1 U223 ( .A1(B[2]), .A2(A[2]), .ZN(n139) );
  NAND2_X1 U224 ( .A1(n267), .A2(n26), .ZN(n1) );
  NAND2_X1 U225 ( .A1(B[7]), .A2(A[7]), .ZN(n117) );
  NAND2_X1 U226 ( .A1(B[5]), .A2(A[5]), .ZN(n125) );
  INV_X1 U227 ( .A(n79), .ZN(n77) );
  NOR2_X1 U228 ( .A1(n253), .A2(n71), .ZN(n69) );
  INV_X1 U229 ( .A(n153), .ZN(n71) );
  NAND2_X1 U230 ( .A1(B[1]), .A2(A[1]), .ZN(n143) );
  NAND2_X1 U231 ( .A1(n157), .A2(n97), .ZN(n12) );
  NAND2_X1 U232 ( .A1(B[12]), .A2(A[12]), .ZN(n97) );
  NAND2_X1 U233 ( .A1(B[22]), .A2(A[22]), .ZN(n29) );
  INV_X1 U234 ( .A(n260), .ZN(n50) );
  NAND2_X1 U235 ( .A1(n260), .A2(n150), .ZN(n43) );
  NAND2_X1 U236 ( .A1(n152), .A2(n67), .ZN(n7) );
  NAND2_X1 U237 ( .A1(n148), .A2(n34), .ZN(n3) );
  NAND2_X1 U238 ( .A1(B[21]), .A2(A[21]), .ZN(n34) );
  AOI21_X1 U239 ( .B1(n150), .B2(n57), .A(n46), .ZN(n44) );
  NAND2_X1 U240 ( .A1(n154), .A2(n83), .ZN(n9) );
  NAND2_X1 U241 ( .A1(n156), .A2(n94), .ZN(n11) );
  NAND2_X1 U242 ( .A1(B[9]), .A2(A[9]), .ZN(n109) );
  INV_X1 U243 ( .A(n138), .ZN(n167) );
  NOR2_X1 U244 ( .A1(B[2]), .A2(A[2]), .ZN(n138) );
  NAND2_X1 U245 ( .A1(n149), .A2(n41), .ZN(n4) );
  NAND2_X1 U246 ( .A1(n153), .A2(n74), .ZN(n8) );
  OAI21_X1 U247 ( .B1(n79), .B2(n71), .A(n74), .ZN(n70) );
  INV_X1 U248 ( .A(n100), .ZN(n158) );
  NOR2_X1 U249 ( .A1(B[11]), .A2(A[11]), .ZN(n100) );
  NAND2_X1 U250 ( .A1(B[17]), .A2(A[17]), .ZN(n67) );
  NAND2_X1 U251 ( .A1(n147), .A2(n29), .ZN(n2) );
  INV_X1 U252 ( .A(n116), .ZN(n162) );
  NOR2_X1 U253 ( .A1(B[7]), .A2(A[7]), .ZN(n116) );
  INV_X1 U254 ( .A(n124), .ZN(n164) );
  NOR2_X1 U255 ( .A1(B[5]), .A2(A[5]), .ZN(n124) );
  NAND2_X1 U256 ( .A1(n155), .A2(n88), .ZN(n10) );
  INV_X1 U257 ( .A(n88), .ZN(n86) );
  NAND2_X1 U258 ( .A1(B[3]), .A2(A[3]), .ZN(n136) );
  NAND2_X1 U259 ( .A1(B[15]), .A2(A[15]), .ZN(n83) );
  NAND2_X1 U260 ( .A1(B[13]), .A2(A[13]), .ZN(n94) );
  NAND2_X1 U261 ( .A1(B[20]), .A2(A[20]), .ZN(n41) );
  NAND2_X1 U262 ( .A1(B[16]), .A2(A[16]), .ZN(n74) );
  NAND2_X1 U263 ( .A1(n261), .A2(n106), .ZN(n14) );
  INV_X1 U264 ( .A(n106), .ZN(n104) );
  NAND2_X1 U265 ( .A1(B[10]), .A2(A[10]), .ZN(n106) );
  OAI21_X1 U266 ( .B1(n138), .B2(n140), .A(n139), .ZN(n137) );
  INV_X1 U267 ( .A(n141), .ZN(n140) );
  NAND2_X1 U268 ( .A1(A[14]), .A2(B[14]), .ZN(n88) );
  NOR2_X1 U269 ( .A1(n87), .A2(n82), .ZN(n80) );
  NAND2_X1 U270 ( .A1(n150), .A2(n255), .ZN(n5) );
  INV_X1 U271 ( .A(n48), .ZN(n46) );
  NAND2_X1 U272 ( .A1(B[19]), .A2(A[19]), .ZN(n48) );
  INV_X1 U273 ( .A(n96), .ZN(n157) );
  NOR2_X1 U274 ( .A1(B[12]), .A2(A[12]), .ZN(n96) );
  INV_X1 U275 ( .A(n108), .ZN(n160) );
  NOR2_X1 U276 ( .A1(B[9]), .A2(A[9]), .ZN(n108) );
  INV_X1 U277 ( .A(n130), .ZN(n128) );
  NAND2_X1 U278 ( .A1(B[4]), .A2(A[4]), .ZN(n130) );
  INV_X1 U279 ( .A(n122), .ZN(n120) );
  NAND2_X1 U280 ( .A1(A[6]), .A2(B[6]), .ZN(n122) );
  INV_X1 U281 ( .A(n114), .ZN(n112) );
  NAND2_X1 U282 ( .A1(B[8]), .A2(A[8]), .ZN(n114) );
  INV_X1 U283 ( .A(n81), .ZN(n79) );
  OAI21_X1 U284 ( .B1(n254), .B2(n88), .A(n83), .ZN(n81) );
  INV_X1 U285 ( .A(n136), .ZN(n134) );
  AOI21_X1 U286 ( .B1(n107), .B2(n261), .A(n104), .ZN(n102) );
  NAND2_X1 U287 ( .A1(n260), .A2(n59), .ZN(n6) );
  INV_X1 U288 ( .A(n59), .ZN(n57) );
  NAND2_X1 U289 ( .A1(B[18]), .A2(A[18]), .ZN(n59) );
  INV_X1 U290 ( .A(n87), .ZN(n155) );
  NOR2_X1 U291 ( .A1(B[14]), .A2(A[14]), .ZN(n87) );
  INV_X1 U292 ( .A(n250), .ZN(n156) );
  OAI21_X1 U293 ( .B1(n93), .B2(n97), .A(n94), .ZN(n92) );
  NOR2_X1 U294 ( .A1(n93), .A2(n96), .ZN(n91) );
  NOR2_X1 U295 ( .A1(B[13]), .A2(A[13]), .ZN(n93) );
  AOI21_X1 U296 ( .B1(n264), .B2(n137), .A(n134), .ZN(n132) );
  INV_X1 U297 ( .A(n40), .ZN(n149) );
  OAI21_X1 U298 ( .B1(n257), .B2(n48), .A(n41), .ZN(n39) );
  NOR2_X1 U299 ( .A1(B[20]), .A2(A[20]), .ZN(n40) );
  INV_X1 U300 ( .A(n73), .ZN(n153) );
  NOR2_X1 U301 ( .A1(B[16]), .A2(A[16]), .ZN(n73) );
  INV_X1 U302 ( .A(n47), .ZN(n150) );
  NOR2_X1 U303 ( .A1(B[19]), .A2(A[19]), .ZN(n47) );
  INV_X1 U304 ( .A(n254), .ZN(n154) );
  NOR2_X1 U305 ( .A1(B[15]), .A2(A[15]), .ZN(n82) );
  INV_X1 U306 ( .A(n66), .ZN(n152) );
  OAI21_X1 U307 ( .B1(n66), .B2(n74), .A(n67), .ZN(n65) );
  NOR2_X1 U308 ( .A1(B[17]), .A2(A[17]), .ZN(n66) );
  NOR2_X1 U309 ( .A1(n40), .A2(n47), .ZN(n38) );
  AOI21_X1 U310 ( .B1(n262), .B2(n131), .A(n128), .ZN(n126) );
  INV_X1 U311 ( .A(n132), .ZN(n131) );
  NAND2_X1 U312 ( .A1(n258), .A2(n80), .ZN(n62) );
  AOI21_X1 U313 ( .B1(n81), .B2(n258), .A(n65), .ZN(n63) );
  NAND2_X1 U314 ( .A1(n38), .A2(n260), .ZN(n36) );
  INV_X1 U315 ( .A(n33), .ZN(n148) );
  AOI21_X1 U316 ( .B1(n38), .B2(n57), .A(n39), .ZN(n37) );
  NOR2_X1 U317 ( .A1(n36), .A2(n33), .ZN(n31) );
  OAI21_X1 U318 ( .B1(n251), .B2(n62), .A(n63), .ZN(n61) );
  OAI21_X1 U319 ( .B1(n37), .B2(n33), .A(n34), .ZN(n32) );
  INV_X1 U320 ( .A(n28), .ZN(n147) );
  NOR2_X1 U321 ( .A1(B[22]), .A2(A[22]), .ZN(n28) );
  OAI21_X1 U322 ( .B1(n126), .B2(n124), .A(n125), .ZN(n123) );
  INV_X1 U323 ( .A(n142), .ZN(n168) );
  OAI21_X1 U324 ( .B1(n142), .B2(n145), .A(n143), .ZN(n141) );
  NOR2_X1 U325 ( .A1(B[1]), .A2(A[1]), .ZN(n142) );
  OAI21_X1 U326 ( .B1(n102), .B2(n100), .A(n101), .ZN(n99) );
  XOR2_X1 U327 ( .A(n23), .B(n145), .Z(SUM[1]) );
  NAND2_X1 U328 ( .A1(n168), .A2(n143), .ZN(n23) );
  XOR2_X1 U329 ( .A(n22), .B(n140), .Z(SUM[2]) );
  NAND2_X1 U330 ( .A1(n167), .A2(n139), .ZN(n22) );
  XNOR2_X1 U331 ( .A(n21), .B(n137), .ZN(SUM[3]) );
  NAND2_X1 U332 ( .A1(n264), .A2(n136), .ZN(n21) );
  XNOR2_X1 U333 ( .A(n20), .B(n131), .ZN(SUM[4]) );
  NAND2_X1 U334 ( .A1(n262), .A2(n130), .ZN(n20) );
  XOR2_X1 U335 ( .A(n19), .B(n126), .Z(SUM[5]) );
  NAND2_X1 U336 ( .A1(n164), .A2(n125), .ZN(n19) );
  XNOR2_X1 U337 ( .A(n18), .B(n123), .ZN(SUM[6]) );
  NAND2_X1 U338 ( .A1(n263), .A2(n122), .ZN(n18) );
  AOI21_X1 U339 ( .B1(n263), .B2(n123), .A(n120), .ZN(n118) );
  XOR2_X1 U340 ( .A(n118), .B(n17), .Z(SUM[7]) );
  NAND2_X1 U341 ( .A1(n162), .A2(n117), .ZN(n17) );
  XNOR2_X1 U342 ( .A(n16), .B(n248), .ZN(SUM[8]) );
  NAND2_X1 U343 ( .A1(n265), .A2(n114), .ZN(n16) );
  OAI21_X1 U344 ( .B1(n118), .B2(n116), .A(n117), .ZN(n115) );
  XOR2_X1 U345 ( .A(n15), .B(n110), .Z(SUM[9]) );
  AOI21_X1 U346 ( .B1(n265), .B2(n115), .A(n112), .ZN(n110) );
  NAND2_X1 U347 ( .A1(n160), .A2(n109), .ZN(n15) );
  XNOR2_X1 U348 ( .A(n14), .B(n252), .ZN(SUM[10]) );
  OAI21_X1 U349 ( .B1(n108), .B2(n110), .A(n109), .ZN(n107) );
  XOR2_X1 U350 ( .A(n102), .B(n13), .Z(SUM[11]) );
  XOR2_X1 U351 ( .A(n12), .B(n98), .Z(SUM[12]) );
  INV_X1 U352 ( .A(n99), .ZN(n98) );
  XNOR2_X1 U353 ( .A(n95), .B(n11), .ZN(SUM[13]) );
  OAI21_X1 U354 ( .B1(n98), .B2(n96), .A(n97), .ZN(n95) );
  XNOR2_X1 U355 ( .A(n89), .B(n10), .ZN(SUM[14]) );
  INV_X1 U356 ( .A(n251), .ZN(n89) );
  XOR2_X1 U357 ( .A(n60), .B(n6), .Z(SUM[18]) );
  INV_X1 U358 ( .A(n61), .ZN(n60) );
  XOR2_X1 U359 ( .A(n75), .B(n8), .Z(SUM[16]) );
  AOI21_X1 U360 ( .B1(n89), .B2(n80), .A(n77), .ZN(n75) );
  XOR2_X1 U361 ( .A(n84), .B(n9), .Z(SUM[15]) );
  AOI21_X1 U362 ( .B1(n89), .B2(n155), .A(n86), .ZN(n84) );
  XOR2_X1 U363 ( .A(n68), .B(n7), .Z(SUM[17]) );
  AOI21_X1 U364 ( .B1(n69), .B2(n89), .A(n70), .ZN(n68) );
  XOR2_X1 U365 ( .A(n30), .B(n2), .Z(SUM[22]) );
  AOI21_X1 U366 ( .B1(n249), .B2(n31), .A(n32), .ZN(n30) );
  XNOR2_X1 U367 ( .A(n49), .B(n5), .ZN(SUM[19]) );
  OAI21_X1 U368 ( .B1(n60), .B2(n50), .A(n59), .ZN(n49) );
  XNOR2_X1 U369 ( .A(n42), .B(n4), .ZN(SUM[20]) );
  OAI21_X1 U370 ( .B1(n60), .B2(n43), .A(n44), .ZN(n42) );
  XNOR2_X1 U371 ( .A(n35), .B(n3), .ZN(SUM[21]) );
  OAI21_X1 U372 ( .B1(n60), .B2(n36), .A(n256), .ZN(n35) );
  XNOR2_X1 U373 ( .A(n27), .B(n1), .ZN(SUM[23]) );
  OAI21_X1 U374 ( .B1(n259), .B2(n28), .A(n29), .ZN(n27) );
endmodule


module datapath_DW01_add_21 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n40, n41, n42, n45, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n61, n62, n63, n65, n66, n67, n68, n69,
         n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n91, n93, n94, n96, n98, n99, n100, n102,
         n104, n105, n106, n107, n108, n110, n112, n113, n114, n115, n116,
         n118, n120, n121, n122, n123, n124, n126, n128, n129, n130, n131,
         n132, n133, n134, n136, n138, n139, n142, n143, n144, n145, n146,
         n147, n151, n153, n155, n157, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262;

  FA_X1 U173 ( .A(B[2]), .B(A[2]), .CI(n133), .CO(n132), .S(SUM[2]) );
  FA_X1 U174 ( .A(n134), .B(A[1]), .CI(B[1]), .CO(n133), .S(SUM[1]) );
  INV_X1 U184 ( .A(n245), .ZN(n40) );
  AND2_X1 U185 ( .A1(n261), .A2(n136), .ZN(SUM[0]) );
  AOI21_X1 U186 ( .B1(n259), .B2(n121), .A(n118), .ZN(n238) );
  AOI21_X1 U187 ( .B1(n256), .B2(n45), .A(n245), .ZN(n239) );
  CLKBUF_X1 U188 ( .A(n61), .Z(n240) );
  NOR2_X1 U189 ( .A1(B[21]), .A2(A[21]), .ZN(n241) );
  CLKBUF_X1 U190 ( .A(n105), .Z(n242) );
  CLKBUF_X1 U191 ( .A(n108), .Z(n243) );
  CLKBUF_X1 U192 ( .A(n100), .Z(n244) );
  AND2_X1 U193 ( .A1(B[20]), .A2(A[20]), .ZN(n245) );
  CLKBUF_X1 U194 ( .A(n55), .Z(n246) );
  CLKBUF_X1 U195 ( .A(n62), .Z(n247) );
  CLKBUF_X1 U196 ( .A(n76), .Z(n248) );
  NOR2_X2 U197 ( .A1(B[14]), .A2(A[14]), .ZN(n81) );
  CLKBUF_X1 U198 ( .A(n252), .Z(n249) );
  NOR2_X1 U199 ( .A1(A[16]), .A2(B[16]), .ZN(n250) );
  AOI21_X1 U200 ( .B1(n258), .B2(n129), .A(n126), .ZN(n251) );
  NOR2_X1 U201 ( .A1(B[18]), .A2(A[18]), .ZN(n252) );
  OR2_X1 U202 ( .A1(B[10]), .A2(A[10]), .ZN(n253) );
  OR2_X1 U203 ( .A1(B[19]), .A2(A[19]), .ZN(n254) );
  OR2_X1 U204 ( .A1(B[11]), .A2(A[11]), .ZN(n255) );
  OR2_X1 U205 ( .A1(B[20]), .A2(A[20]), .ZN(n256) );
  OR2_X1 U206 ( .A1(B[12]), .A2(A[12]), .ZN(n257) );
  OR2_X1 U207 ( .A1(B[4]), .A2(A[4]), .ZN(n258) );
  OR2_X1 U208 ( .A1(A[6]), .A2(B[6]), .ZN(n259) );
  OR2_X1 U209 ( .A1(B[8]), .A2(A[8]), .ZN(n260) );
  OR2_X1 U210 ( .A1(B[0]), .A2(A[0]), .ZN(n261) );
  OR2_X1 U211 ( .A1(B[23]), .A2(A[23]), .ZN(n262) );
  INV_X1 U212 ( .A(n136), .ZN(n134) );
  NAND2_X1 U213 ( .A1(B[0]), .A2(A[0]), .ZN(n136) );
  NAND2_X1 U214 ( .A1(B[23]), .A2(A[23]), .ZN(n25) );
  NAND2_X1 U215 ( .A1(B[3]), .A2(A[3]), .ZN(n131) );
  NAND2_X1 U216 ( .A1(B[7]), .A2(A[7]), .ZN(n115) );
  NAND2_X1 U217 ( .A1(n262), .A2(n25), .ZN(n2) );
  NAND2_X1 U218 ( .A1(B[5]), .A2(A[5]), .ZN(n123) );
  NAND2_X1 U219 ( .A1(B[9]), .A2(A[9]), .ZN(n107) );
  INV_X1 U220 ( .A(n130), .ZN(n157) );
  NOR2_X1 U221 ( .A1(B[3]), .A2(A[3]), .ZN(n130) );
  NAND2_X1 U222 ( .A1(B[22]), .A2(A[22]), .ZN(n28) );
  NAND2_X1 U223 ( .A1(n139), .A2(n33), .ZN(n4) );
  NAND2_X1 U224 ( .A1(B[21]), .A2(A[21]), .ZN(n33) );
  INV_X1 U225 ( .A(n114), .ZN(n153) );
  NOR2_X1 U226 ( .A1(B[7]), .A2(A[7]), .ZN(n114) );
  INV_X1 U227 ( .A(n67), .ZN(n65) );
  NAND2_X1 U228 ( .A1(n146), .A2(n82), .ZN(n11) );
  NAND2_X1 U229 ( .A1(n144), .A2(n71), .ZN(n9) );
  NAND2_X1 U230 ( .A1(n147), .A2(n85), .ZN(n12) );
  NAND2_X1 U231 ( .A1(n256), .A2(n40), .ZN(n5) );
  NAND2_X1 U232 ( .A1(n255), .A2(n98), .ZN(n14) );
  OAI21_X1 U233 ( .B1(n130), .B2(n1), .A(n131), .ZN(n129) );
  INV_X1 U234 ( .A(n132), .ZN(n1) );
  NAND2_X1 U235 ( .A1(n138), .A2(n28), .ZN(n3) );
  INV_X1 U236 ( .A(n122), .ZN(n155) );
  NOR2_X1 U237 ( .A1(B[5]), .A2(A[5]), .ZN(n122) );
  NAND2_X1 U238 ( .A1(B[6]), .A2(A[6]), .ZN(n120) );
  NAND2_X1 U239 ( .A1(B[11]), .A2(A[11]), .ZN(n98) );
  NAND2_X1 U240 ( .A1(B[16]), .A2(A[16]), .ZN(n71) );
  NAND2_X1 U241 ( .A1(n142), .A2(n246), .ZN(n7) );
  NAND2_X1 U242 ( .A1(n256), .A2(n254), .ZN(n35) );
  INV_X1 U243 ( .A(n254), .ZN(n42) );
  INV_X1 U244 ( .A(n104), .ZN(n102) );
  NAND2_X1 U245 ( .A1(B[10]), .A2(A[10]), .ZN(n104) );
  NAND2_X1 U246 ( .A1(n143), .A2(n247), .ZN(n8) );
  NAND2_X1 U247 ( .A1(n254), .A2(n47), .ZN(n6) );
  NAND2_X1 U248 ( .A1(B[13]), .A2(A[13]), .ZN(n85) );
  NAND2_X1 U249 ( .A1(B[14]), .A2(A[14]), .ZN(n82) );
  NAND2_X1 U250 ( .A1(n257), .A2(n255), .ZN(n88) );
  INV_X1 U251 ( .A(n106), .ZN(n151) );
  NOR2_X1 U252 ( .A1(B[9]), .A2(A[9]), .ZN(n106) );
  NAND2_X1 U253 ( .A1(n145), .A2(n248), .ZN(n10) );
  INV_X1 U254 ( .A(n248), .ZN(n74) );
  NAND2_X1 U255 ( .A1(B[15]), .A2(A[15]), .ZN(n76) );
  INV_X1 U256 ( .A(n68), .ZN(n66) );
  NOR2_X1 U257 ( .A1(n75), .A2(n250), .ZN(n68) );
  NOR2_X1 U258 ( .A1(B[16]), .A2(A[16]), .ZN(n70) );
  INV_X1 U259 ( .A(n112), .ZN(n110) );
  NAND2_X1 U260 ( .A1(B[8]), .A2(A[8]), .ZN(n112) );
  NAND2_X1 U261 ( .A1(B[18]), .A2(A[18]), .ZN(n55) );
  NAND2_X1 U262 ( .A1(B[17]), .A2(A[17]), .ZN(n62) );
  NAND2_X1 U263 ( .A1(B[19]), .A2(A[19]), .ZN(n47) );
  INV_X1 U264 ( .A(n128), .ZN(n126) );
  NAND2_X1 U265 ( .A1(B[4]), .A2(A[4]), .ZN(n128) );
  AOI21_X1 U266 ( .B1(n257), .B2(n96), .A(n91), .ZN(n89) );
  INV_X1 U267 ( .A(n98), .ZN(n96) );
  INV_X1 U268 ( .A(n120), .ZN(n118) );
  INV_X1 U269 ( .A(n69), .ZN(n67) );
  OAI21_X1 U270 ( .B1(n70), .B2(n76), .A(n71), .ZN(n69) );
  INV_X1 U271 ( .A(n47), .ZN(n45) );
  AOI21_X1 U272 ( .B1(n258), .B2(n129), .A(n126), .ZN(n124) );
  NAND2_X1 U273 ( .A1(n257), .A2(n93), .ZN(n13) );
  INV_X1 U274 ( .A(n93), .ZN(n91) );
  NAND2_X1 U275 ( .A1(B[12]), .A2(A[12]), .ZN(n93) );
  OAI21_X1 U276 ( .B1(n124), .B2(n122), .A(n123), .ZN(n121) );
  AOI21_X1 U277 ( .B1(n256), .B2(n45), .A(n245), .ZN(n36) );
  INV_X1 U278 ( .A(n81), .ZN(n146) );
  OAI21_X1 U279 ( .B1(n81), .B2(n85), .A(n82), .ZN(n80) );
  INV_X1 U280 ( .A(n84), .ZN(n147) );
  NOR2_X1 U281 ( .A1(n81), .A2(n84), .ZN(n79) );
  NOR2_X1 U282 ( .A1(B[13]), .A2(A[13]), .ZN(n84) );
  INV_X1 U283 ( .A(n75), .ZN(n145) );
  NOR2_X1 U284 ( .A1(B[15]), .A2(A[15]), .ZN(n75) );
  INV_X1 U285 ( .A(n70), .ZN(n144) );
  NOR2_X1 U286 ( .A1(n66), .A2(n240), .ZN(n57) );
  OAI21_X1 U287 ( .B1(n67), .B2(n240), .A(n247), .ZN(n58) );
  INV_X1 U288 ( .A(n32), .ZN(n139) );
  NOR2_X1 U289 ( .A1(B[21]), .A2(A[21]), .ZN(n32) );
  OAI21_X1 U290 ( .B1(n116), .B2(n114), .A(n115), .ZN(n113) );
  AOI21_X1 U291 ( .B1(n259), .B2(n121), .A(n118), .ZN(n116) );
  INV_X1 U292 ( .A(n240), .ZN(n143) );
  NOR2_X1 U293 ( .A1(n252), .A2(n61), .ZN(n52) );
  NOR2_X1 U294 ( .A1(B[17]), .A2(A[17]), .ZN(n61) );
  OAI21_X1 U295 ( .B1(n36), .B2(n32), .A(n33), .ZN(n31) );
  NAND2_X1 U296 ( .A1(n52), .A2(n68), .ZN(n50) );
  NOR2_X1 U297 ( .A1(n35), .A2(n241), .ZN(n30) );
  AOI21_X1 U298 ( .B1(n69), .B2(n52), .A(n53), .ZN(n51) );
  INV_X1 U299 ( .A(n249), .ZN(n142) );
  OAI21_X1 U300 ( .B1(n54), .B2(n62), .A(n55), .ZN(n53) );
  NOR2_X1 U301 ( .A1(B[18]), .A2(A[18]), .ZN(n54) );
  OAI21_X1 U302 ( .B1(n50), .B2(n78), .A(n51), .ZN(n49) );
  AOI21_X1 U303 ( .B1(n87), .B2(n79), .A(n80), .ZN(n78) );
  INV_X1 U304 ( .A(n27), .ZN(n138) );
  NOR2_X1 U305 ( .A1(B[22]), .A2(A[22]), .ZN(n27) );
  AOI21_X1 U306 ( .B1(n113), .B2(n260), .A(n110), .ZN(n108) );
  OAI21_X1 U307 ( .B1(n88), .B2(n100), .A(n89), .ZN(n87) );
  AOI21_X1 U308 ( .B1(n253), .B2(n105), .A(n102), .ZN(n100) );
  OAI21_X1 U309 ( .B1(n108), .B2(n106), .A(n107), .ZN(n105) );
  XNOR2_X1 U310 ( .A(n22), .B(n132), .ZN(SUM[3]) );
  NAND2_X1 U311 ( .A1(n157), .A2(n131), .ZN(n22) );
  XNOR2_X1 U312 ( .A(n21), .B(n129), .ZN(SUM[4]) );
  NAND2_X1 U313 ( .A1(n258), .A2(n128), .ZN(n21) );
  XOR2_X1 U314 ( .A(n20), .B(n251), .Z(SUM[5]) );
  NAND2_X1 U315 ( .A1(n155), .A2(n123), .ZN(n20) );
  XOR2_X1 U316 ( .A(n238), .B(n18), .Z(SUM[7]) );
  NAND2_X1 U317 ( .A1(n153), .A2(n115), .ZN(n18) );
  XNOR2_X1 U318 ( .A(n19), .B(n121), .ZN(SUM[6]) );
  NAND2_X1 U319 ( .A1(n259), .A2(n120), .ZN(n19) );
  XNOR2_X1 U320 ( .A(n113), .B(n17), .ZN(SUM[8]) );
  NAND2_X1 U321 ( .A1(n260), .A2(n112), .ZN(n17) );
  XOR2_X1 U322 ( .A(n243), .B(n16), .Z(SUM[9]) );
  NAND2_X1 U323 ( .A1(n151), .A2(n107), .ZN(n16) );
  XNOR2_X1 U324 ( .A(n15), .B(n242), .ZN(SUM[10]) );
  NAND2_X1 U325 ( .A1(n253), .A2(n104), .ZN(n15) );
  XNOR2_X1 U326 ( .A(n99), .B(n14), .ZN(SUM[11]) );
  INV_X1 U327 ( .A(n244), .ZN(n99) );
  XOR2_X1 U328 ( .A(n94), .B(n13), .Z(SUM[12]) );
  AOI21_X1 U329 ( .B1(n99), .B2(n255), .A(n96), .ZN(n94) );
  XOR2_X1 U330 ( .A(n86), .B(n12), .Z(SUM[13]) );
  INV_X1 U331 ( .A(n87), .ZN(n86) );
  XNOR2_X1 U332 ( .A(n83), .B(n11), .ZN(SUM[14]) );
  OAI21_X1 U333 ( .B1(n86), .B2(n84), .A(n85), .ZN(n83) );
  XNOR2_X1 U334 ( .A(n77), .B(n10), .ZN(SUM[15]) );
  INV_X1 U335 ( .A(n78), .ZN(n77) );
  XOR2_X1 U336 ( .A(n63), .B(n8), .Z(SUM[17]) );
  AOI21_X1 U337 ( .B1(n77), .B2(n68), .A(n65), .ZN(n63) );
  XOR2_X1 U338 ( .A(n72), .B(n9), .Z(SUM[16]) );
  AOI21_X1 U339 ( .B1(n77), .B2(n145), .A(n74), .ZN(n72) );
  XOR2_X1 U340 ( .A(n56), .B(n7), .Z(SUM[18]) );
  AOI21_X1 U341 ( .B1(n57), .B2(n77), .A(n58), .ZN(n56) );
  XOR2_X1 U342 ( .A(n48), .B(n6), .Z(SUM[19]) );
  INV_X1 U343 ( .A(n49), .ZN(n48) );
  XOR2_X1 U344 ( .A(n29), .B(n3), .Z(SUM[22]) );
  AOI21_X1 U345 ( .B1(n49), .B2(n30), .A(n31), .ZN(n29) );
  XNOR2_X1 U346 ( .A(n41), .B(n5), .ZN(SUM[20]) );
  OAI21_X1 U347 ( .B1(n48), .B2(n42), .A(n47), .ZN(n41) );
  XNOR2_X1 U348 ( .A(n34), .B(n4), .ZN(SUM[21]) );
  OAI21_X1 U349 ( .B1(n48), .B2(n35), .A(n239), .ZN(n34) );
  XNOR2_X1 U350 ( .A(n26), .B(n2), .ZN(SUM[23]) );
  OAI21_X1 U351 ( .B1(n29), .B2(n27), .A(n28), .ZN(n26) );
endmodule


module datapath_DW01_add_22 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n27, n28, n29, n30, n32, n34,
         n35, n36, n37, n38, n39, n40, n41, n43, n45, n46, n47, n48, n51, n52,
         n53, n54, n55, n57, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n71, n73, n74, n75, n76, n78, n80, n81, n82, n83, n84, n86, n88,
         n89, n91, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n109, n111, n112, n113, n114, n115, n117,
         n119, n120, n121, n122, n123, n125, n127, n128, n129, n130, n131,
         n133, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n148, n152, n153, n154, n160, n161, n163, n165, n167,
         n169, n170, n171, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279;

  AND2_X1 U200 ( .A1(n265), .A2(n266), .ZN(n251) );
  AND2_X1 U201 ( .A1(n265), .A2(n266), .ZN(n62) );
  CLKBUF_X1 U202 ( .A(n120), .Z(n252) );
  CLKBUF_X1 U203 ( .A(n123), .Z(n253) );
  NOR2_X1 U204 ( .A1(A[13]), .A2(B[13]), .ZN(n254) );
  CLKBUF_X1 U205 ( .A(n65), .Z(n255) );
  CLKBUF_X1 U206 ( .A(n104), .Z(n256) );
  CLKBUF_X1 U207 ( .A(n112), .Z(n257) );
  NOR2_X1 U208 ( .A1(B[18]), .A2(A[18]), .ZN(n65) );
  AOI21_X1 U209 ( .B1(n257), .B2(n269), .A(n109), .ZN(n258) );
  OR2_X2 U210 ( .A1(B[22]), .A2(A[22]), .ZN(n273) );
  AOI21_X1 U211 ( .B1(n268), .B2(n78), .A(n71), .ZN(n259) );
  CLKBUF_X1 U212 ( .A(n82), .Z(n260) );
  CLKBUF_X1 U213 ( .A(n95), .Z(n261) );
  CLKBUF_X1 U214 ( .A(B[13]), .Z(n262) );
  OR2_X1 U215 ( .A1(n262), .A2(A[13]), .ZN(n263) );
  AOI21_X1 U216 ( .B1(n279), .B2(n120), .A(n117), .ZN(n264) );
  NAND2_X1 U217 ( .A1(n82), .A2(n63), .ZN(n265) );
  INV_X1 U218 ( .A(n64), .ZN(n266) );
  AND2_X1 U219 ( .A1(n270), .A2(n148), .ZN(SUM[0]) );
  OR2_X1 U220 ( .A1(B[17]), .A2(A[17]), .ZN(n268) );
  OR2_X1 U221 ( .A1(B[10]), .A2(A[10]), .ZN(n269) );
  OR2_X1 U222 ( .A1(B[0]), .A2(A[0]), .ZN(n270) );
  OR2_X1 U223 ( .A1(B[15]), .A2(A[15]), .ZN(n271) );
  OR2_X1 U224 ( .A1(A[16]), .A2(B[16]), .ZN(n272) );
  OR2_X1 U225 ( .A1(B[14]), .A2(A[14]), .ZN(n274) );
  OR2_X1 U226 ( .A1(B[21]), .A2(A[21]), .ZN(n275) );
  OR2_X1 U227 ( .A1(B[23]), .A2(A[23]), .ZN(n276) );
  OR2_X1 U228 ( .A1(B[6]), .A2(A[6]), .ZN(n277) );
  OR2_X1 U229 ( .A1(A[4]), .A2(B[4]), .ZN(n278) );
  OR2_X1 U230 ( .A1(B[8]), .A2(A[8]), .ZN(n279) );
  NOR2_X1 U231 ( .A1(B[13]), .A2(A[13]), .ZN(n98) );
  NAND2_X1 U232 ( .A1(B[0]), .A2(A[0]), .ZN(n148) );
  NAND2_X1 U233 ( .A1(B[23]), .A2(A[23]), .ZN(n27) );
  NAND2_X1 U234 ( .A1(n276), .A2(n27), .ZN(n2) );
  INV_X1 U235 ( .A(n59), .ZN(n57) );
  NAND2_X1 U236 ( .A1(B[7]), .A2(A[7]), .ZN(n122) );
  NAND2_X1 U237 ( .A1(n161), .A2(n106), .ZN(n14) );
  NAND2_X1 U238 ( .A1(B[11]), .A2(A[11]), .ZN(n106) );
  NAND2_X1 U239 ( .A1(n153), .A2(n152), .ZN(n47) );
  NAND2_X1 U240 ( .A1(B[3]), .A2(A[3]), .ZN(n138) );
  NAND2_X1 U241 ( .A1(n273), .A2(n34), .ZN(n3) );
  NAND2_X1 U242 ( .A1(n163), .A2(n114), .ZN(n16) );
  NAND2_X1 U243 ( .A1(B[9]), .A2(A[9]), .ZN(n114) );
  NAND2_X1 U244 ( .A1(B[5]), .A2(A[5]), .ZN(n130) );
  AOI21_X1 U245 ( .B1(n278), .B2(n136), .A(n133), .ZN(n131) );
  NAND2_X1 U246 ( .A1(n154), .A2(n66), .ZN(n7) );
  NAND2_X1 U247 ( .A1(B[18]), .A2(A[18]), .ZN(n66) );
  OAI21_X1 U248 ( .B1(n95), .B2(n83), .A(n84), .ZN(n82) );
  NAND2_X1 U249 ( .A1(B[22]), .A2(A[22]), .ZN(n34) );
  NAND2_X1 U250 ( .A1(n160), .A2(n102), .ZN(n13) );
  NAND2_X1 U251 ( .A1(B[12]), .A2(A[12]), .ZN(n102) );
  NAND2_X1 U252 ( .A1(n263), .A2(n99), .ZN(n12) );
  NAND2_X1 U253 ( .A1(n153), .A2(n61), .ZN(n6) );
  INV_X1 U254 ( .A(n61), .ZN(n59) );
  NAND2_X1 U255 ( .A1(B[19]), .A2(A[19]), .ZN(n61) );
  AOI21_X1 U256 ( .B1(n128), .B2(n277), .A(n125), .ZN(n123) );
  OAI21_X1 U257 ( .B1(n137), .B2(n139), .A(n138), .ZN(n136) );
  INV_X1 U258 ( .A(n140), .ZN(n139) );
  INV_X1 U259 ( .A(n272), .ZN(n75) );
  NAND2_X1 U260 ( .A1(B[2]), .A2(A[2]), .ZN(n142) );
  INV_X1 U261 ( .A(n121), .ZN(n165) );
  NOR2_X1 U262 ( .A1(B[7]), .A2(A[7]), .ZN(n121) );
  INV_X1 U263 ( .A(n105), .ZN(n161) );
  NOR2_X1 U264 ( .A1(B[11]), .A2(A[11]), .ZN(n105) );
  AOI21_X1 U265 ( .B1(n271), .B2(n91), .A(n86), .ZN(n84) );
  NAND2_X1 U266 ( .A1(n274), .A2(n271), .ZN(n83) );
  NAND2_X1 U267 ( .A1(B[13]), .A2(A[13]), .ZN(n99) );
  INV_X1 U268 ( .A(n34), .ZN(n32) );
  INV_X1 U269 ( .A(n113), .ZN(n163) );
  NOR2_X1 U270 ( .A1(B[9]), .A2(A[9]), .ZN(n113) );
  INV_X1 U271 ( .A(n78), .ZN(n76) );
  INV_X1 U272 ( .A(n38), .ZN(n36) );
  INV_X1 U273 ( .A(n101), .ZN(n160) );
  NOR2_X1 U274 ( .A1(B[12]), .A2(A[12]), .ZN(n101) );
  INV_X1 U275 ( .A(n129), .ZN(n167) );
  NOR2_X1 U276 ( .A1(B[5]), .A2(A[5]), .ZN(n129) );
  NAND2_X1 U277 ( .A1(n272), .A2(n80), .ZN(n9) );
  INV_X1 U278 ( .A(n135), .ZN(n133) );
  NAND2_X1 U279 ( .A1(B[4]), .A2(A[4]), .ZN(n135) );
  INV_X1 U280 ( .A(n39), .ZN(n37) );
  AOI21_X1 U281 ( .B1(n39), .B2(n273), .A(n32), .ZN(n30) );
  OAI21_X1 U282 ( .B1(n61), .B2(n40), .A(n41), .ZN(n39) );
  INV_X1 U283 ( .A(n137), .ZN(n169) );
  NOR2_X1 U284 ( .A1(B[3]), .A2(A[3]), .ZN(n137) );
  NAND2_X1 U285 ( .A1(n269), .A2(n111), .ZN(n15) );
  INV_X1 U286 ( .A(n111), .ZN(n109) );
  NAND2_X1 U287 ( .A1(B[10]), .A2(A[10]), .ZN(n111) );
  INV_X1 U288 ( .A(n119), .ZN(n117) );
  NAND2_X1 U289 ( .A1(B[8]), .A2(A[8]), .ZN(n119) );
  AOI21_X1 U290 ( .B1(n275), .B2(n52), .A(n43), .ZN(n41) );
  INV_X1 U291 ( .A(n127), .ZN(n125) );
  NAND2_X1 U292 ( .A1(B[6]), .A2(A[6]), .ZN(n127) );
  NAND2_X1 U293 ( .A1(n271), .A2(n88), .ZN(n10) );
  INV_X1 U294 ( .A(n88), .ZN(n86) );
  NAND2_X1 U295 ( .A1(B[15]), .A2(A[15]), .ZN(n88) );
  NAND2_X1 U296 ( .A1(B[16]), .A2(A[16]), .ZN(n80) );
  NAND2_X1 U297 ( .A1(n274), .A2(n93), .ZN(n11) );
  INV_X1 U298 ( .A(n93), .ZN(n91) );
  NAND2_X1 U299 ( .A1(B[14]), .A2(A[14]), .ZN(n93) );
  NAND2_X1 U300 ( .A1(n38), .A2(n273), .ZN(n29) );
  NOR2_X1 U301 ( .A1(n40), .A2(n60), .ZN(n38) );
  INV_X1 U302 ( .A(n144), .ZN(n143) );
  AOI21_X1 U303 ( .B1(n152), .B2(n59), .A(n52), .ZN(n48) );
  INV_X1 U304 ( .A(n141), .ZN(n170) );
  OAI21_X1 U305 ( .B1(n141), .B2(n143), .A(n142), .ZN(n140) );
  NOR2_X1 U306 ( .A1(B[2]), .A2(A[2]), .ZN(n141) );
  INV_X1 U307 ( .A(n80), .ZN(n78) );
  NAND2_X1 U308 ( .A1(n275), .A2(n51), .ZN(n40) );
  NAND2_X1 U309 ( .A1(n268), .A2(n73), .ZN(n8) );
  INV_X1 U310 ( .A(n73), .ZN(n71) );
  NAND2_X1 U311 ( .A1(B[17]), .A2(A[17]), .ZN(n73) );
  OAI21_X1 U312 ( .B1(n98), .B2(n102), .A(n99), .ZN(n97) );
  NOR2_X1 U313 ( .A1(n101), .A2(n254), .ZN(n96) );
  INV_X1 U314 ( .A(n255), .ZN(n154) );
  NAND2_X1 U315 ( .A1(n272), .A2(n268), .ZN(n68) );
  NAND2_X1 U316 ( .A1(n275), .A2(n45), .ZN(n4) );
  INV_X1 U317 ( .A(n45), .ZN(n43) );
  NAND2_X1 U318 ( .A1(B[21]), .A2(A[21]), .ZN(n45) );
  NAND2_X1 U319 ( .A1(n152), .A2(n54), .ZN(n5) );
  INV_X1 U320 ( .A(n54), .ZN(n52) );
  NAND2_X1 U321 ( .A1(B[20]), .A2(A[20]), .ZN(n54) );
  OAI21_X1 U322 ( .B1(n131), .B2(n129), .A(n130), .ZN(n128) );
  AOI21_X1 U323 ( .B1(n112), .B2(n269), .A(n109), .ZN(n107) );
  AOI21_X1 U324 ( .B1(n268), .B2(n78), .A(n71), .ZN(n69) );
  OAI21_X1 U325 ( .B1(n145), .B2(n148), .A(n146), .ZN(n144) );
  NAND2_X1 U326 ( .A1(B[1]), .A2(A[1]), .ZN(n146) );
  INV_X1 U327 ( .A(n60), .ZN(n153) );
  NOR2_X1 U328 ( .A1(B[19]), .A2(A[19]), .ZN(n60) );
  NOR2_X1 U329 ( .A1(n68), .A2(n65), .ZN(n63) );
  INV_X1 U330 ( .A(n53), .ZN(n152) );
  INV_X1 U331 ( .A(n53), .ZN(n51) );
  NOR2_X1 U332 ( .A1(B[20]), .A2(A[20]), .ZN(n53) );
  OAI21_X1 U333 ( .B1(n65), .B2(n69), .A(n66), .ZN(n64) );
  INV_X1 U334 ( .A(n145), .ZN(n171) );
  NOR2_X1 U335 ( .A1(B[1]), .A2(A[1]), .ZN(n145) );
  AOI21_X1 U336 ( .B1(n104), .B2(n96), .A(n97), .ZN(n95) );
  OAI21_X1 U337 ( .B1(n107), .B2(n105), .A(n106), .ZN(n104) );
  XOR2_X1 U338 ( .A(n24), .B(n148), .Z(SUM[1]) );
  NAND2_X1 U339 ( .A1(n171), .A2(n146), .ZN(n24) );
  XOR2_X1 U340 ( .A(n23), .B(n143), .Z(SUM[2]) );
  NAND2_X1 U341 ( .A1(n170), .A2(n142), .ZN(n23) );
  XOR2_X1 U342 ( .A(n22), .B(n139), .Z(SUM[3]) );
  NAND2_X1 U343 ( .A1(n169), .A2(n138), .ZN(n22) );
  XNOR2_X1 U344 ( .A(n21), .B(n136), .ZN(SUM[4]) );
  NAND2_X1 U345 ( .A1(n278), .A2(n135), .ZN(n21) );
  XOR2_X1 U346 ( .A(n20), .B(n131), .Z(SUM[5]) );
  NAND2_X1 U347 ( .A1(n167), .A2(n130), .ZN(n20) );
  NAND2_X1 U348 ( .A1(n165), .A2(n122), .ZN(n18) );
  XNOR2_X1 U349 ( .A(n19), .B(n128), .ZN(SUM[6]) );
  NAND2_X1 U350 ( .A1(n277), .A2(n127), .ZN(n19) );
  XOR2_X1 U351 ( .A(n18), .B(n253), .Z(SUM[7]) );
  NAND2_X1 U352 ( .A1(n279), .A2(n119), .ZN(n17) );
  XNOR2_X1 U353 ( .A(n17), .B(n252), .ZN(SUM[8]) );
  OAI21_X1 U354 ( .B1(n121), .B2(n123), .A(n122), .ZN(n120) );
  XOR2_X1 U355 ( .A(n16), .B(n264), .Z(SUM[9]) );
  AOI21_X1 U356 ( .B1(n120), .B2(n279), .A(n117), .ZN(n115) );
  XNOR2_X1 U357 ( .A(n15), .B(n257), .ZN(SUM[10]) );
  OAI21_X1 U358 ( .B1(n115), .B2(n113), .A(n114), .ZN(n112) );
  XOR2_X1 U359 ( .A(n258), .B(n14), .Z(SUM[11]) );
  XOR2_X1 U360 ( .A(n13), .B(n103), .Z(SUM[12]) );
  INV_X1 U361 ( .A(n256), .ZN(n103) );
  XNOR2_X1 U362 ( .A(n100), .B(n12), .ZN(SUM[13]) );
  OAI21_X1 U363 ( .B1(n103), .B2(n101), .A(n102), .ZN(n100) );
  XNOR2_X1 U364 ( .A(n94), .B(n11), .ZN(SUM[14]) );
  INV_X1 U365 ( .A(n261), .ZN(n94) );
  XOR2_X1 U366 ( .A(n89), .B(n10), .Z(SUM[15]) );
  AOI21_X1 U367 ( .B1(n94), .B2(n274), .A(n91), .ZN(n89) );
  XOR2_X1 U368 ( .A(n81), .B(n9), .Z(SUM[16]) );
  INV_X1 U369 ( .A(n260), .ZN(n81) );
  XNOR2_X1 U370 ( .A(n74), .B(n8), .ZN(SUM[17]) );
  OAI21_X1 U371 ( .B1(n81), .B2(n75), .A(n76), .ZN(n74) );
  XNOR2_X1 U372 ( .A(n67), .B(n7), .ZN(SUM[18]) );
  OAI21_X1 U373 ( .B1(n81), .B2(n68), .A(n259), .ZN(n67) );
  XOR2_X1 U374 ( .A(n251), .B(n6), .Z(SUM[19]) );
  XNOR2_X1 U375 ( .A(n55), .B(n5), .ZN(SUM[20]) );
  OAI21_X1 U376 ( .B1(n251), .B2(n60), .A(n57), .ZN(n55) );
  XNOR2_X1 U377 ( .A(n35), .B(n3), .ZN(SUM[22]) );
  OAI21_X1 U378 ( .B1(n62), .B2(n36), .A(n37), .ZN(n35) );
  XNOR2_X1 U379 ( .A(n28), .B(n2), .ZN(SUM[23]) );
  OAI21_X1 U380 ( .B1(n62), .B2(n29), .A(n30), .ZN(n28) );
  XNOR2_X1 U381 ( .A(n46), .B(n4), .ZN(SUM[21]) );
  OAI21_X1 U382 ( .B1(n62), .B2(n47), .A(n48), .ZN(n46) );
endmodule


module datapath_DW01_add_23 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n2, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n26, n27, n29, n31, n32, n33, n34, n35, n36, n37,
         n38, n39, n40, n41, n42, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n72, n73, n74, n75, n77, n79, n80, n81, n82, n83, n85, n87, n88,
         n90, n92, n93, n94, n96, n98, n99, n100, n101, n105, n106, n108, n110,
         n111, n112, n114, n116, n117, n118, n119, n120, n122, n124, n125,
         n126, n127, n128, n130, n132, n133, n134, n135, n136, n138, n140,
         n141, n142, n144, n146, n147, n148, n149, n151, n155, n157, n158,
         n167, n169, n171, n174, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n291;

  BUF_X1 U203 ( .A(n32), .Z(n254) );
  AND2_X1 U204 ( .A1(B[16]), .A2(A[16]), .ZN(n267) );
  INV_X1 U205 ( .A(n267), .ZN(n72) );
  OAI21_X1 U206 ( .B1(n120), .B2(n118), .A(n119), .ZN(n117) );
  OR2_X1 U207 ( .A1(B[21]), .A2(A[21]), .ZN(n255) );
  OR2_X1 U208 ( .A1(n264), .A2(A[19]), .ZN(n256) );
  BUF_X1 U209 ( .A(n81), .Z(n260) );
  INV_X1 U210 ( .A(n269), .ZN(n105) );
  INV_X1 U211 ( .A(n79), .ZN(n257) );
  XNOR2_X1 U212 ( .A(n55), .B(n258), .ZN(SUM[19]) );
  AND2_X1 U213 ( .A1(n256), .A2(n54), .ZN(n258) );
  CLKBUF_X1 U214 ( .A(n120), .Z(n259) );
  CLKBUF_X1 U215 ( .A(n60), .Z(n261) );
  NOR2_X1 U216 ( .A1(B[21]), .A2(A[21]), .ZN(n262) );
  NOR2_X1 U217 ( .A1(B[21]), .A2(A[21]), .ZN(n37) );
  NOR2_X1 U218 ( .A1(A[19]), .A2(B[19]), .ZN(n263) );
  CLKBUF_X1 U219 ( .A(B[19]), .Z(n264) );
  NOR2_X1 U220 ( .A1(B[19]), .A2(A[19]), .ZN(n53) );
  AOI21_X1 U221 ( .B1(n283), .B2(n108), .A(n269), .ZN(n265) );
  CLKBUF_X1 U222 ( .A(n276), .Z(n266) );
  OAI21_X1 U223 ( .B1(n100), .B2(n112), .A(n265), .ZN(n268) );
  AND2_X1 U224 ( .A1(B[11]), .A2(A[11]), .ZN(n269) );
  XNOR2_X1 U225 ( .A(n46), .B(n270), .ZN(SUM[20]) );
  AND2_X1 U226 ( .A1(n155), .A2(n45), .ZN(n270) );
  XNOR2_X1 U227 ( .A(n39), .B(n271), .ZN(SUM[21]) );
  AND2_X1 U228 ( .A1(n255), .A2(n38), .ZN(n271) );
  XNOR2_X1 U229 ( .A(n27), .B(n272), .ZN(SUM[23]) );
  AND2_X1 U230 ( .A1(n291), .A2(n26), .ZN(n272) );
  AOI21_X1 U231 ( .B1(n277), .B2(n268), .A(n96), .ZN(n273) );
  OR2_X2 U232 ( .A1(B[11]), .A2(A[11]), .ZN(n283) );
  AOI21_X1 U233 ( .B1(n266), .B2(n77), .A(n267), .ZN(n274) );
  AOI21_X1 U234 ( .B1(n81), .B2(n62), .A(n63), .ZN(n275) );
  OR2_X1 U235 ( .A1(B[16]), .A2(A[16]), .ZN(n276) );
  OR2_X1 U236 ( .A1(B[12]), .A2(A[12]), .ZN(n277) );
  OR2_X1 U237 ( .A1(B[0]), .A2(A[0]), .ZN(n278) );
  OR2_X1 U238 ( .A1(B[15]), .A2(A[15]), .ZN(n279) );
  OR2_X1 U239 ( .A1(B[10]), .A2(A[10]), .ZN(n280) );
  OR2_X1 U240 ( .A1(B[14]), .A2(A[14]), .ZN(n281) );
  OR2_X1 U241 ( .A1(B[13]), .A2(A[13]), .ZN(n282) );
  OR2_X1 U242 ( .A1(B[9]), .A2(A[9]), .ZN(n284) );
  OR2_X1 U243 ( .A1(B[22]), .A2(A[22]), .ZN(n285) );
  OR2_X1 U244 ( .A1(B[5]), .A2(A[5]), .ZN(n286) );
  OR2_X1 U245 ( .A1(B[3]), .A2(A[3]), .ZN(n287) );
  OR2_X1 U246 ( .A1(B[2]), .A2(A[2]), .ZN(n288) );
  OR2_X1 U247 ( .A1(B[7]), .A2(A[7]), .ZN(n289) );
  AND2_X1 U248 ( .A1(n278), .A2(n151), .ZN(SUM[0]) );
  OR2_X1 U249 ( .A1(B[23]), .A2(A[23]), .ZN(n291) );
  NAND2_X1 U250 ( .A1(B[0]), .A2(A[0]), .ZN(n151) );
  NAND2_X1 U251 ( .A1(B[23]), .A2(A[23]), .ZN(n26) );
  NAND2_X1 U252 ( .A1(n285), .A2(n31), .ZN(n2) );
  INV_X1 U253 ( .A(n31), .ZN(n29) );
  NAND2_X1 U254 ( .A1(B[22]), .A2(A[22]), .ZN(n31) );
  NAND2_X1 U255 ( .A1(B[1]), .A2(A[1]), .ZN(n149) );
  NAND2_X1 U256 ( .A1(B[8]), .A2(A[8]), .ZN(n119) );
  NAND2_X1 U257 ( .A1(B[19]), .A2(A[19]), .ZN(n54) );
  INV_X1 U258 ( .A(n155), .ZN(n42) );
  NAND2_X1 U259 ( .A1(B[21]), .A2(A[21]), .ZN(n38) );
  NAND2_X1 U260 ( .A1(B[2]), .A2(A[2]), .ZN(n146) );
  NAND2_X1 U261 ( .A1(B[20]), .A2(A[20]), .ZN(n45) );
  NAND2_X1 U262 ( .A1(B[3]), .A2(A[3]), .ZN(n140) );
  NAND2_X1 U263 ( .A1(n284), .A2(n116), .ZN(n15) );
  INV_X1 U264 ( .A(n116), .ZN(n114) );
  NAND2_X1 U265 ( .A1(B[9]), .A2(A[9]), .ZN(n116) );
  INV_X1 U266 ( .A(n279), .ZN(n74) );
  INV_X1 U267 ( .A(n49), .ZN(n47) );
  NAND2_X1 U268 ( .A1(B[6]), .A2(A[6]), .ZN(n127) );
  INV_X1 U269 ( .A(n148), .ZN(n174) );
  NOR2_X1 U270 ( .A1(B[1]), .A2(A[1]), .ZN(n148) );
  NAND2_X1 U271 ( .A1(B[4]), .A2(A[4]), .ZN(n135) );
  NOR2_X1 U272 ( .A1(B[18]), .A2(A[18]), .ZN(n58) );
  NAND2_X1 U273 ( .A1(n158), .A2(n65), .ZN(n7) );
  NAND2_X1 U274 ( .A1(B[17]), .A2(A[17]), .ZN(n65) );
  NAND2_X1 U275 ( .A1(n279), .A2(n79), .ZN(n9) );
  INV_X1 U276 ( .A(n118), .ZN(n167) );
  NOR2_X1 U277 ( .A1(B[8]), .A2(A[8]), .ZN(n118) );
  NAND2_X1 U278 ( .A1(n157), .A2(n59), .ZN(n6) );
  INV_X1 U279 ( .A(n59), .ZN(n57) );
  NAND2_X1 U280 ( .A1(B[18]), .A2(A[18]), .ZN(n59) );
  NAND2_X1 U281 ( .A1(n283), .A2(n105), .ZN(n13) );
  INV_X1 U282 ( .A(n77), .ZN(n75) );
  INV_X1 U283 ( .A(n134), .ZN(n171) );
  NOR2_X1 U284 ( .A1(B[4]), .A2(A[4]), .ZN(n134) );
  OAI21_X1 U285 ( .B1(n148), .B2(n151), .A(n149), .ZN(n147) );
  INV_X1 U286 ( .A(n146), .ZN(n144) );
  OAI21_X1 U287 ( .B1(n59), .B2(n263), .A(n54), .ZN(n52) );
  INV_X1 U288 ( .A(n132), .ZN(n130) );
  NAND2_X1 U289 ( .A1(B[5]), .A2(A[5]), .ZN(n132) );
  NOR2_X1 U290 ( .A1(n37), .A2(n44), .ZN(n35) );
  NOR2_X1 U291 ( .A1(B[20]), .A2(A[20]), .ZN(n44) );
  NAND2_X1 U292 ( .A1(n277), .A2(n98), .ZN(n12) );
  INV_X1 U293 ( .A(n98), .ZN(n96) );
  NAND2_X1 U294 ( .A1(B[12]), .A2(A[12]), .ZN(n98) );
  INV_X1 U295 ( .A(n51), .ZN(n49) );
  NOR2_X1 U296 ( .A1(n58), .A2(n53), .ZN(n51) );
  INV_X1 U297 ( .A(n50), .ZN(n48) );
  NAND2_X1 U298 ( .A1(n280), .A2(n110), .ZN(n14) );
  INV_X1 U299 ( .A(n110), .ZN(n108) );
  NAND2_X1 U300 ( .A1(B[10]), .A2(A[10]), .ZN(n110) );
  NAND2_X1 U301 ( .A1(n276), .A2(n279), .ZN(n67) );
  INV_X1 U302 ( .A(n124), .ZN(n122) );
  NAND2_X1 U303 ( .A1(B[7]), .A2(A[7]), .ZN(n124) );
  AOI21_X1 U304 ( .B1(n288), .B2(n147), .A(n144), .ZN(n142) );
  INV_X1 U305 ( .A(n140), .ZN(n138) );
  NAND2_X1 U306 ( .A1(B[15]), .A2(A[15]), .ZN(n79) );
  INV_X1 U307 ( .A(n126), .ZN(n169) );
  NOR2_X1 U308 ( .A1(B[6]), .A2(A[6]), .ZN(n126) );
  AOI21_X1 U309 ( .B1(n281), .B2(n90), .A(n85), .ZN(n83) );
  INV_X1 U310 ( .A(n79), .ZN(n77) );
  AOI21_X1 U311 ( .B1(n287), .B2(n141), .A(n138), .ZN(n136) );
  INV_X1 U312 ( .A(n142), .ZN(n141) );
  NAND2_X1 U313 ( .A1(n281), .A2(n87), .ZN(n10) );
  INV_X1 U314 ( .A(n87), .ZN(n85) );
  NAND2_X1 U315 ( .A1(B[14]), .A2(A[14]), .ZN(n87) );
  INV_X1 U316 ( .A(n52), .ZN(n50) );
  AOI21_X1 U317 ( .B1(n52), .B2(n35), .A(n36), .ZN(n34) );
  AOI21_X1 U318 ( .B1(n117), .B2(n284), .A(n114), .ZN(n112) );
  NAND2_X1 U319 ( .A1(n266), .A2(n72), .ZN(n8) );
  INV_X1 U320 ( .A(n64), .ZN(n158) );
  NOR2_X1 U321 ( .A1(n67), .A2(n64), .ZN(n62) );
  NOR2_X1 U322 ( .A1(B[17]), .A2(A[17]), .ZN(n64) );
  OAI21_X1 U323 ( .B1(n262), .B2(n45), .A(n38), .ZN(n36) );
  INV_X1 U324 ( .A(n44), .ZN(n155) );
  OAI21_X1 U325 ( .B1(n61), .B2(n33), .A(n34), .ZN(n32) );
  NAND2_X1 U326 ( .A1(n51), .A2(n35), .ZN(n33) );
  NOR2_X1 U327 ( .A1(n49), .A2(n42), .ZN(n40) );
  OAI21_X1 U328 ( .B1(n50), .B2(n42), .A(n45), .ZN(n41) );
  AOI21_X1 U329 ( .B1(n276), .B2(n257), .A(n267), .ZN(n68) );
  NAND2_X1 U330 ( .A1(n282), .A2(n92), .ZN(n11) );
  INV_X1 U331 ( .A(n92), .ZN(n90) );
  NAND2_X1 U332 ( .A1(B[13]), .A2(A[13]), .ZN(n92) );
  INV_X1 U333 ( .A(n58), .ZN(n157) );
  AOI21_X1 U334 ( .B1(n133), .B2(n286), .A(n130), .ZN(n128) );
  OAI21_X1 U335 ( .B1(n134), .B2(n136), .A(n135), .ZN(n133) );
  NAND2_X1 U336 ( .A1(n283), .A2(n280), .ZN(n100) );
  AOI21_X1 U337 ( .B1(n283), .B2(n108), .A(n269), .ZN(n101) );
  NAND2_X1 U338 ( .A1(n282), .A2(n281), .ZN(n82) );
  AOI21_X1 U339 ( .B1(n277), .B2(n99), .A(n96), .ZN(n94) );
  AOI21_X1 U340 ( .B1(n81), .B2(n62), .A(n63), .ZN(n61) );
  OAI21_X1 U341 ( .B1(n68), .B2(n64), .A(n65), .ZN(n63) );
  OAI21_X1 U342 ( .B1(n82), .B2(n94), .A(n83), .ZN(n81) );
  OAI21_X1 U343 ( .B1(n128), .B2(n126), .A(n127), .ZN(n125) );
  OAI21_X1 U344 ( .B1(n100), .B2(n112), .A(n101), .ZN(n99) );
  XOR2_X1 U345 ( .A(n23), .B(n151), .Z(SUM[1]) );
  NAND2_X1 U346 ( .A1(n174), .A2(n149), .ZN(n23) );
  XNOR2_X1 U347 ( .A(n22), .B(n147), .ZN(SUM[2]) );
  NAND2_X1 U348 ( .A1(n288), .A2(n146), .ZN(n22) );
  XNOR2_X1 U349 ( .A(n21), .B(n141), .ZN(SUM[3]) );
  NAND2_X1 U350 ( .A1(n287), .A2(n140), .ZN(n21) );
  XOR2_X1 U351 ( .A(n20), .B(n136), .Z(SUM[4]) );
  NAND2_X1 U352 ( .A1(n171), .A2(n135), .ZN(n20) );
  XNOR2_X1 U353 ( .A(n19), .B(n133), .ZN(SUM[5]) );
  NAND2_X1 U354 ( .A1(n286), .A2(n132), .ZN(n19) );
  XOR2_X1 U355 ( .A(n18), .B(n128), .Z(SUM[6]) );
  NAND2_X1 U356 ( .A1(n169), .A2(n127), .ZN(n18) );
  XNOR2_X1 U357 ( .A(n17), .B(n125), .ZN(SUM[7]) );
  NAND2_X1 U358 ( .A1(n289), .A2(n124), .ZN(n17) );
  AOI21_X1 U359 ( .B1(n289), .B2(n125), .A(n122), .ZN(n120) );
  XOR2_X1 U360 ( .A(n16), .B(n259), .Z(SUM[8]) );
  NAND2_X1 U361 ( .A1(n167), .A2(n119), .ZN(n16) );
  XNOR2_X1 U362 ( .A(n15), .B(n117), .ZN(SUM[9]) );
  XNOR2_X1 U363 ( .A(n14), .B(n111), .ZN(SUM[10]) );
  INV_X1 U364 ( .A(n112), .ZN(n111) );
  XNOR2_X1 U365 ( .A(n12), .B(n268), .ZN(SUM[12]) );
  XOR2_X1 U366 ( .A(n106), .B(n13), .Z(SUM[11]) );
  AOI21_X1 U367 ( .B1(n111), .B2(n280), .A(n108), .ZN(n106) );
  XNOR2_X1 U368 ( .A(n11), .B(n93), .ZN(SUM[13]) );
  INV_X1 U369 ( .A(n273), .ZN(n93) );
  XOR2_X1 U370 ( .A(n88), .B(n10), .Z(SUM[14]) );
  AOI21_X1 U371 ( .B1(n282), .B2(n93), .A(n90), .ZN(n88) );
  XOR2_X1 U372 ( .A(n80), .B(n9), .Z(SUM[15]) );
  INV_X1 U373 ( .A(n260), .ZN(n80) );
  XNOR2_X1 U374 ( .A(n73), .B(n8), .ZN(SUM[16]) );
  OAI21_X1 U375 ( .B1(n80), .B2(n74), .A(n75), .ZN(n73) );
  XNOR2_X1 U376 ( .A(n66), .B(n7), .ZN(SUM[17]) );
  OAI21_X1 U377 ( .B1(n80), .B2(n67), .A(n274), .ZN(n66) );
  XNOR2_X1 U378 ( .A(n261), .B(n6), .ZN(SUM[18]) );
  INV_X1 U379 ( .A(n275), .ZN(n60) );
  XNOR2_X1 U380 ( .A(n254), .B(n2), .ZN(SUM[22]) );
  AOI21_X1 U381 ( .B1(n60), .B2(n47), .A(n48), .ZN(n46) );
  AOI21_X1 U382 ( .B1(n32), .B2(n285), .A(n29), .ZN(n27) );
  AOI21_X1 U383 ( .B1(n60), .B2(n157), .A(n57), .ZN(n55) );
  AOI21_X1 U384 ( .B1(n60), .B2(n40), .A(n41), .ZN(n39) );
endmodule


module datapath ( clk, data_in, addr_x, wr_en_x, addr_a1, addr_a2, addr_a3, 
        addr_a4, addr_a5, addr_a6, addr_a7, addr_a8, wr_en_a1, wr_en_a2, 
        wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6, wr_en_a7, wr_en_a8, addr_y, 
        wr_en_y, clear_acc, clc, clc1, data_out );
  input [11:0] data_in;
  input [2:0] addr_x;
  input [2:0] addr_a1;
  input [2:0] addr_a2;
  input [2:0] addr_a3;
  input [2:0] addr_a4;
  input [2:0] addr_a5;
  input [2:0] addr_a6;
  input [2:0] addr_a7;
  input [2:0] addr_a8;
  input [2:0] addr_y;
  output [23:0] data_out;
  input clk, wr_en_x, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5,
         wr_en_a6, wr_en_a7, wr_en_a8, wr_en_y, clear_acc, clc, clc1;
  wire   n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n210, n211, n212, n213, n215, n216, n217, n221, n222,
         n223, n224, n227, n228, n231, n232, n235, n236, n239, n240, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n314, n315, n316, n317, n318, n319, n320, n321, n323, n324, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, \mul_out1[9] , \mul_out1[8] ,
         \mul_out1[7] , \mul_out1[6] , \mul_out1[5] , \mul_out1[4] ,
         \mul_out1[3] , \mul_out1[2] , \mul_out1[23] , \mul_out1[22] ,
         \mul_out1[21] , \mul_out1[20] , \mul_out1[1] , \mul_out1[19] ,
         \mul_out1[18] , \mul_out1[17] , \mul_out1[16] , \mul_out1[15] ,
         \mul_out1[14] , \mul_out1[13] , \mul_out1[12] , \mul_out1[11] ,
         \mul_out1[10] , \mul_out1[0] , \mul_out2[9] , \mul_out2[8] ,
         \mul_out2[7] , \mul_out2[6] , \mul_out2[5] , \mul_out2[4] ,
         \mul_out2[3] , \mul_out2[2] , \mul_out2[23] , \mul_out2[22] ,
         \mul_out2[21] , \mul_out2[20] , \mul_out2[1] , \mul_out2[19] ,
         \mul_out2[18] , \mul_out2[17] , \mul_out2[16] , \mul_out2[15] ,
         \mul_out2[14] , \mul_out2[13] , \mul_out2[12] , \mul_out2[11] ,
         \mul_out2[10] , \mul_out2[0] , \mul_out3[9] , \mul_out3[8] ,
         \mul_out3[7] , \mul_out3[6] , \mul_out3[5] , \mul_out3[4] ,
         \mul_out3[3] , \mul_out3[2] , \mul_out3[23] , \mul_out3[22] ,
         \mul_out3[21] , \mul_out3[20] , \mul_out3[1] , \mul_out3[19] ,
         \mul_out3[18] , \mul_out3[17] , \mul_out3[16] , \mul_out3[15] ,
         \mul_out3[14] , \mul_out3[13] , \mul_out3[12] , \mul_out3[11] ,
         \mul_out3[10] , \mul_out3[0] , \mul_out4[9] , \mul_out4[8] ,
         \mul_out4[7] , \mul_out4[6] , \mul_out4[5] , \mul_out4[4] ,
         \mul_out4[3] , \mul_out4[2] , \mul_out4[23] , \mul_out4[22] ,
         \mul_out4[21] , \mul_out4[20] , \mul_out4[1] , \mul_out4[19] ,
         \mul_out4[18] , \mul_out4[17] , \mul_out4[16] , \mul_out4[15] ,
         \mul_out4[14] , \mul_out4[13] , \mul_out4[12] , \mul_out4[11] ,
         \mul_out4[10] , \mul_out4[0] , \mul_out5[9] , \mul_out5[8] ,
         \mul_out5[7] , \mul_out5[6] , \mul_out5[5] , \mul_out5[4] ,
         \mul_out5[3] , \mul_out5[2] , \mul_out5[23] , \mul_out5[22] ,
         \mul_out5[21] , \mul_out5[20] , \mul_out5[1] , \mul_out5[19] ,
         \mul_out5[18] , \mul_out5[17] , \mul_out5[16] , \mul_out5[15] ,
         \mul_out5[14] , \mul_out5[13] , \mul_out5[12] , \mul_out5[11] ,
         \mul_out5[10] , \mul_out5[0] , \mul_out6[9] , \mul_out6[8] ,
         \mul_out6[7] , \mul_out6[6] , \mul_out6[5] , \mul_out6[4] ,
         \mul_out6[3] , \mul_out6[2] , \mul_out6[23] , \mul_out6[22] ,
         \mul_out6[21] , \mul_out6[20] , \mul_out6[1] , \mul_out6[19] ,
         \mul_out6[18] , \mul_out6[17] , \mul_out6[16] , \mul_out6[15] ,
         \mul_out6[14] , \mul_out6[13] , \mul_out6[12] , \mul_out6[11] ,
         \mul_out6[10] , \mul_out6[0] , \mul_out7[9] , \mul_out7[8] ,
         \mul_out7[7] , \mul_out7[6] , \mul_out7[5] , \mul_out7[4] ,
         \mul_out7[3] , \mul_out7[2] , \mul_out7[23] , \mul_out7[22] ,
         \mul_out7[21] , \mul_out7[20] , \mul_out7[1] , \mul_out7[19] ,
         \mul_out7[18] , \mul_out7[17] , \mul_out7[16] , \mul_out7[15] ,
         \mul_out7[14] , \mul_out7[13] , \mul_out7[12] , \mul_out7[11] ,
         \mul_out7[10] , \mul_out7[0] , \mul_out8[9] , \mul_out8[8] ,
         \mul_out8[7] , \mul_out8[6] , \mul_out8[5] , \mul_out8[4] ,
         \mul_out8[3] , \mul_out8[2] , \mul_out8[23] , \mul_out8[22] ,
         \mul_out8[21] , \mul_out8[20] , \mul_out8[1] , \mul_out8[19] ,
         \mul_out8[18] , \mul_out8[17] , \mul_out8[16] , \mul_out8[15] ,
         \mul_out8[14] , \mul_out8[13] , \mul_out8[12] , \mul_out8[11] ,
         \mul_out8[10] , \mul_out8[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n29, n30, n31, n32, n53, n54, n55, n56, n129,
         n130, n131, n132, n133, n134, n153, n154, n155, n156, n157, n158,
         n173, n174, n175, n176, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n214, n218, n219, n220, n225, n226, n229, n230, n233,
         n234, n237, n238, n241, n242, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n322, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822;
  wire   [11:0] data_out_x;
  wire   [11:0] data_out_a1;
  wire   [11:0] data_out_a2;
  wire   [11:0] data_out_a3;
  wire   [11:0] data_out_a4;
  wire   [11:0] data_out_a5;
  wire   [11:0] data_out_a6;
  wire   [11:0] data_out_a7;
  wire   [11:0] data_out_a8;
  wire   [23:0] f;
  wire   [23:0] f1;
  wire   [23:0] f2;
  wire   [23:0] f3;
  wire   [23:0] f4;
  wire   [23:0] f5;
  wire   [23:0] f6;
  wire   [23:0] f7;
  wire   [23:0] f8;
  wire   [23:0] add_r1;
  wire   [23:0] add_r2;
  wire   [23:0] add_r3;
  wire   [23:0] add_r4;
  wire   [23:0] add_r5;
  wire   [23:0] add_r6;
  wire   [23:0] add_r7;
  wire   [23:0] add_r8;

  DFF_X1 \f1_reg[22]  ( .D(n733), .CK(clk), .Q(f1[22]), .QN(n802) );
  DFF_X1 \f1_reg[15]  ( .D(n726), .CK(clk), .Q(f1[15]), .QN(n17) );
  DFF_X1 \f1_reg[14]  ( .D(n725), .CK(clk), .Q(f1[14]), .QN(n18) );
  DFF_X1 \f1_reg[13]  ( .D(n724), .CK(clk), .Q(f1[13]), .QN(n19) );
  DFF_X1 \f2_reg[19]  ( .D(n706), .CK(clk), .Q(n454), .QN(n37) );
  DFF_X1 \f2_reg[18]  ( .D(n705), .CK(clk), .Q(n456), .QN(n38) );
  DFF_X1 \f2_reg[17]  ( .D(n704), .CK(clk), .Q(f2[17]), .QN(n39) );
  DFF_X1 \f2_reg[16]  ( .D(n703), .CK(clk), .Q(f2[16]), .QN(n40) );
  DFF_X1 \f2_reg[15]  ( .D(n702), .CK(clk), .Q(f2[15]), .QN(n41) );
  DFF_X1 \f2_reg[14]  ( .D(n701), .CK(clk), .Q(f2[14]), .QN(n42) );
  DFF_X1 \f2_reg[13]  ( .D(n700), .CK(clk), .Q(f2[13]), .QN(n43) );
  DFF_X1 \f2_reg[12]  ( .D(n699), .CK(clk), .Q(f2[12]), .QN(n44) );
  DFF_X1 \f2_reg[11]  ( .D(n698), .CK(clk), .Q(f2[11]), .QN(n45) );
  DFF_X1 \f3_reg[22]  ( .D(n685), .CK(clk), .Q(n477), .QN(n58) );
  DFF_X1 \f3_reg[19]  ( .D(n682), .CK(clk), .Q(n481), .QN(n61) );
  DFF_X1 \f3_reg[18]  ( .D(n681), .CK(clk), .Q(n483), .QN(n62) );
  DFF_X1 \f3_reg[17]  ( .D(n680), .CK(clk), .Q(f3[17]), .QN(n63) );
  DFF_X1 \f3_reg[16]  ( .D(n679), .CK(clk), .Q(f3[16]), .QN(n64) );
  DFF_X1 \f3_reg[15]  ( .D(n678), .CK(clk), .Q(f3[15]), .QN(n65) );
  DFF_X1 \f3_reg[14]  ( .D(n677), .CK(clk), .Q(f3[14]), .QN(n66) );
  DFF_X1 \f3_reg[13]  ( .D(n676), .CK(clk), .Q(f3[13]), .QN(n67) );
  DFF_X1 \f3_reg[12]  ( .D(n675), .CK(clk), .Q(f3[12]), .QN(n68) );
  DFF_X1 \f4_reg[22]  ( .D(n661), .CK(clk), .Q(f4[22]), .QN(n82) );
  DFF_X1 \f4_reg[18]  ( .D(n657), .CK(clk), .Q(f4[18]), .QN(n86) );
  DFF_X1 \f4_reg[17]  ( .D(n656), .CK(clk), .Q(f4[17]), .QN(n87) );
  DFF_X1 \f4_reg[16]  ( .D(n655), .CK(clk), .Q(f4[16]), .QN(n88) );
  DFF_X1 \f4_reg[15]  ( .D(n654), .CK(clk), .Q(f4[15]), .QN(n89) );
  DFF_X1 \f4_reg[14]  ( .D(n653), .CK(clk), .Q(f4[14]), .QN(n90) );
  DFF_X1 \f4_reg[13]  ( .D(n652), .CK(clk), .Q(f4[13]), .QN(n91) );
  DFF_X1 \f4_reg[12]  ( .D(n651), .CK(clk), .Q(f4[12]), .QN(n92) );
  DFF_X1 \f5_reg[20]  ( .D(n635), .CK(clk), .Q(n513), .QN(n108) );
  DFF_X1 \f5_reg[16]  ( .D(n631), .CK(clk), .Q(f5[16]), .QN(n112) );
  DFF_X1 \f5_reg[15]  ( .D(n630), .CK(clk), .Q(f5[15]), .QN(n113) );
  DFF_X1 \f5_reg[14]  ( .D(n629), .CK(clk), .Q(f5[14]), .QN(n114) );
  DFF_X1 \f5_reg[13]  ( .D(n628), .CK(clk), .Q(f5[13]), .QN(n115) );
  DFF_X1 \f5_reg[12]  ( .D(n627), .CK(clk), .Q(f5[12]), .QN(n116) );
  DFF_X1 \f6_reg[23]  ( .D(n614), .CK(clk), .Q(n814) );
  DFF_X1 \f6_reg[22]  ( .D(n613), .CK(clk), .Q(n805) );
  DFF_X1 \f6_reg[21]  ( .D(n612), .CK(clk), .Q(n800) );
  DFF_X1 \f6_reg[20]  ( .D(n611), .CK(clk), .Q(n795) );
  DFF_X1 \f6_reg[19]  ( .D(n610), .CK(clk), .Q(n791) );
  DFF_X1 \f6_reg[18]  ( .D(n609), .CK(clk), .Q(n787) );
  DFF_X1 \f6_reg[17]  ( .D(n608), .CK(clk), .Q(f6[17]), .QN(n135) );
  DFF_X1 \f6_reg[16]  ( .D(n607), .CK(clk), .Q(f6[16]), .QN(n136) );
  DFF_X1 \f6_reg[15]  ( .D(n606), .CK(clk), .Q(f6[15]), .QN(n137) );
  DFF_X1 \f6_reg[14]  ( .D(n605), .CK(clk), .Q(f6[14]), .QN(n138) );
  DFF_X1 \f6_reg[13]  ( .D(n604), .CK(clk), .Q(f6[13]), .QN(n139) );
  DFF_X1 \f6_reg[11]  ( .D(n602), .CK(clk), .Q(f6[11]), .QN(n141) );
  DFF_X1 \f7_reg[23]  ( .D(n590), .CK(clk), .Q(n812) );
  DFF_X1 \f7_reg[22]  ( .D(n589), .CK(clk), .Q(n804) );
  DFF_X1 \f7_reg[21]  ( .D(n588), .CK(clk), .Q(n799) );
  DFF_X1 \f7_reg[17]  ( .D(n584), .CK(clk), .Q(f7[17]), .QN(n159) );
  DFF_X1 \f7_reg[16]  ( .D(n583), .CK(clk), .Q(f7[16]), .QN(n160) );
  DFF_X1 \f7_reg[15]  ( .D(n582), .CK(clk), .Q(f7[15]), .QN(n161) );
  DFF_X1 \f7_reg[14]  ( .D(n581), .CK(clk), .Q(f7[14]), .QN(n162) );
  DFF_X1 \f7_reg[13]  ( .D(n580), .CK(clk), .Q(f7[13]), .QN(n163) );
  DFF_X1 \f7_reg[12]  ( .D(n579), .CK(clk), .Q(f7[12]), .QN(n164) );
  DFF_X1 \f_reg[23]  ( .D(n519), .CK(clk), .Q(f[23]), .QN(n7) );
  DFF_X1 \f_reg[22]  ( .D(n520), .CK(clk), .Q(f[22]), .QN(n6) );
  DFF_X1 \f_reg[21]  ( .D(n521), .CK(clk), .Q(f[21]), .QN(n5) );
  DFF_X1 \f8_reg[20]  ( .D(n563), .CK(clk), .Q(f8[20]), .QN(n180) );
  DFF_X1 \f_reg[20]  ( .D(n522), .CK(clk), .Q(f[20]), .QN(n4) );
  DFF_X1 \f_reg[19]  ( .D(n523), .CK(clk), .Q(f[19]), .QN(n3) );
  DFF_X1 \f8_reg[18]  ( .D(n561), .CK(clk), .Q(f8[18]), .QN(n182) );
  DFF_X1 \f_reg[18]  ( .D(n524), .CK(clk), .Q(f[18]), .QN(n2) );
  DFF_X1 \f8_reg[17]  ( .D(n560), .CK(clk), .Q(f8[17]), .QN(n183) );
  DFF_X1 \f_reg[17]  ( .D(n525), .CK(clk), .Q(f[17]) );
  DFF_X1 \f_reg[16]  ( .D(n526), .CK(clk), .Q(f[16]) );
  DFF_X1 \f8_reg[15]  ( .D(n558), .CK(clk), .Q(f8[15]), .QN(n185) );
  DFF_X1 \f_reg[15]  ( .D(n527), .CK(clk), .Q(f[15]) );
  DFF_X1 \f8_reg[14]  ( .D(n557), .CK(clk), .Q(f8[14]), .QN(n186) );
  DFF_X1 \f_reg[14]  ( .D(n528), .CK(clk), .Q(f[14]) );
  DFF_X1 \f8_reg[13]  ( .D(n556), .CK(clk), .Q(f8[13]), .QN(n187) );
  DFF_X1 \f_reg[13]  ( .D(n529), .CK(clk), .Q(f[13]) );
  DFF_X1 \f8_reg[12]  ( .D(n555), .CK(clk), .Q(f8[12]), .QN(n188) );
  DFF_X1 \f_reg[12]  ( .D(n530), .CK(clk), .Q(f[12]) );
  DFF_X1 \f_reg[11]  ( .D(n531), .CK(clk), .Q(f[11]) );
  DFF_X1 \f_reg[10]  ( .D(n532), .CK(clk), .Q(f[10]) );
  DFF_X1 \f_reg[9]  ( .D(n533), .CK(clk), .Q(f[9]) );
  DFF_X1 \f_reg[8]  ( .D(n534), .CK(clk), .Q(f[8]) );
  DFF_X1 \f_reg[7]  ( .D(n535), .CK(clk), .Q(f[7]) );
  DFF_X1 \f_reg[6]  ( .D(n536), .CK(clk), .Q(f[6]) );
  DFF_X1 \f_reg[5]  ( .D(n537), .CK(clk), .Q(f[5]) );
  DFF_X1 \f_reg[4]  ( .D(n538), .CK(clk), .Q(f[4]) );
  DFF_X1 \f_reg[3]  ( .D(n539), .CK(clk), .Q(f[3]), .QN(n8) );
  DFF_X1 \f_reg[2]  ( .D(n540), .CK(clk), .Q(f[2]), .QN(n9) );
  DFF_X1 \f_reg[1]  ( .D(n541), .CK(clk), .Q(f[1]), .QN(n10) );
  DFF_X1 \f_reg[0]  ( .D(n542), .CK(clk), .Q(f[0]), .QN(n11) );
  memory_WIDTH12_SIZE8_LOGSIZE3_0 mem_x ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_x), .addr(addr_x), .wr_en(wr_en_x) );
  memory_WIDTH12_SIZE8_LOGSIZE3_8 mem_a1 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a1), .addr(addr_a1), .wr_en(wr_en_a1) );
  memory_WIDTH12_SIZE8_LOGSIZE3_7 mem_a2 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a2), .addr(addr_a2), .wr_en(wr_en_a2) );
  memory_WIDTH12_SIZE8_LOGSIZE3_6 mem_a3 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a3), .addr(addr_a3), .wr_en(wr_en_a3) );
  memory_WIDTH12_SIZE8_LOGSIZE3_5 mem_a4 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a4), .addr(addr_a4), .wr_en(wr_en_a4) );
  memory_WIDTH12_SIZE8_LOGSIZE3_4 mem_a5 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a5), .addr(addr_a5), .wr_en(wr_en_a5) );
  memory_WIDTH12_SIZE8_LOGSIZE3_3 mem_a6 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a6), .addr(addr_a6), .wr_en(wr_en_a6) );
  memory_WIDTH12_SIZE8_LOGSIZE3_2 mem_a7 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a7), .addr(addr_a7), .wr_en(wr_en_a7) );
  memory_WIDTH12_SIZE8_LOGSIZE3_1 mem_a8 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a8), .addr(addr_a8), .wr_en(wr_en_a8) );
  memory_WIDTH24_SIZE8_LOGSIZE3 mem_y ( .clk(clk), .data_in(f), .data_out(
        data_out), .addr(addr_y), .wr_en(wr_en_y) );
  datapath_DW_mult_tc_16 mult_98 ( .a(data_out_a8), .b({data_out_x[11:3], n29, 
        n14, data_out_x[0]}), .product({\mul_out8[23] , \mul_out8[22] , 
        \mul_out8[21] , \mul_out8[20] , \mul_out8[19] , \mul_out8[18] , 
        \mul_out8[17] , \mul_out8[16] , \mul_out8[15] , \mul_out8[14] , 
        \mul_out8[13] , \mul_out8[12] , \mul_out8[11] , \mul_out8[10] , 
        \mul_out8[9] , \mul_out8[8] , \mul_out8[7] , \mul_out8[6] , 
        \mul_out8[5] , \mul_out8[4] , \mul_out8[3] , \mul_out8[2] , 
        \mul_out8[1] , \mul_out8[0] }) );
  datapath_DW_mult_tc_17 mult_96 ( .a(data_out_a7), .b(data_out_x), .product({
        \mul_out7[23] , \mul_out7[22] , \mul_out7[21] , \mul_out7[20] , 
        \mul_out7[19] , \mul_out7[18] , \mul_out7[17] , \mul_out7[16] , 
        \mul_out7[15] , \mul_out7[14] , \mul_out7[13] , \mul_out7[12] , 
        \mul_out7[11] , \mul_out7[10] , \mul_out7[9] , \mul_out7[8] , 
        \mul_out7[7] , \mul_out7[6] , \mul_out7[5] , \mul_out7[4] , 
        \mul_out7[3] , \mul_out7[2] , \mul_out7[1] , \mul_out7[0] }) );
  datapath_DW_mult_tc_18 mult_94 ( .a(data_out_a6), .b(data_out_x), .product({
        \mul_out6[23] , \mul_out6[22] , \mul_out6[21] , \mul_out6[20] , 
        \mul_out6[19] , \mul_out6[18] , \mul_out6[17] , \mul_out6[16] , 
        \mul_out6[15] , \mul_out6[14] , \mul_out6[13] , \mul_out6[12] , 
        \mul_out6[11] , \mul_out6[10] , \mul_out6[9] , \mul_out6[8] , 
        \mul_out6[7] , \mul_out6[6] , \mul_out6[5] , \mul_out6[4] , 
        \mul_out6[3] , \mul_out6[2] , \mul_out6[1] , \mul_out6[0] }) );
  datapath_DW_mult_tc_19 mult_92 ( .a(data_out_a5), .b({data_out_x[11:5], n134, 
        data_out_x[3:0]}), .product({\mul_out5[23] , \mul_out5[22] , 
        \mul_out5[21] , \mul_out5[20] , \mul_out5[19] , \mul_out5[18] , 
        \mul_out5[17] , \mul_out5[16] , \mul_out5[15] , \mul_out5[14] , 
        \mul_out5[13] , \mul_out5[12] , \mul_out5[11] , \mul_out5[10] , 
        \mul_out5[9] , \mul_out5[8] , \mul_out5[7] , \mul_out5[6] , 
        \mul_out5[5] , \mul_out5[4] , \mul_out5[3] , \mul_out5[2] , 
        \mul_out5[1] , \mul_out5[0] }) );
  datapath_DW_mult_tc_20 mult_90 ( .a(data_out_a4), .b({n31, n133, 
        data_out_x[9:6], n129, n134, data_out_x[3:0]}), .product({
        \mul_out4[23] , \mul_out4[22] , \mul_out4[21] , \mul_out4[20] , 
        \mul_out4[19] , \mul_out4[18] , \mul_out4[17] , \mul_out4[16] , 
        \mul_out4[15] , \mul_out4[14] , \mul_out4[13] , \mul_out4[12] , 
        \mul_out4[11] , \mul_out4[10] , \mul_out4[9] , \mul_out4[8] , 
        \mul_out4[7] , \mul_out4[6] , \mul_out4[5] , \mul_out4[4] , 
        \mul_out4[3] , \mul_out4[2] , \mul_out4[1] , \mul_out4[0] }) );
  datapath_DW_mult_tc_21 mult_88 ( .a(data_out_a3), .b(data_out_x), .product({
        \mul_out3[23] , \mul_out3[22] , \mul_out3[21] , \mul_out3[20] , 
        \mul_out3[19] , \mul_out3[18] , \mul_out3[17] , \mul_out3[16] , 
        \mul_out3[15] , \mul_out3[14] , \mul_out3[13] , \mul_out3[12] , 
        \mul_out3[11] , \mul_out3[10] , \mul_out3[9] , \mul_out3[8] , 
        \mul_out3[7] , \mul_out3[6] , \mul_out3[5] , \mul_out3[4] , 
        \mul_out3[3] , \mul_out3[2] , \mul_out3[1] , \mul_out3[0] }) );
  datapath_DW_mult_tc_22 mult_86 ( .a(data_out_a2), .b({data_out_x[11:5], n134, 
        data_out_x[3:0]}), .product({\mul_out2[23] , \mul_out2[22] , 
        \mul_out2[21] , \mul_out2[20] , \mul_out2[19] , \mul_out2[18] , 
        \mul_out2[17] , \mul_out2[16] , \mul_out2[15] , \mul_out2[14] , 
        \mul_out2[13] , \mul_out2[12] , \mul_out2[11] , \mul_out2[10] , 
        \mul_out2[9] , \mul_out2[8] , \mul_out2[7] , \mul_out2[6] , 
        \mul_out2[5] , \mul_out2[4] , \mul_out2[3] , \mul_out2[2] , 
        \mul_out2[1] , \mul_out2[0] }) );
  datapath_DW_mult_tc_23 mult_84 ( .a(data_out_a1), .b({data_out_x[11:9], n132, 
        data_out_x[7:0]}), .product({\mul_out1[23] , \mul_out1[22] , 
        \mul_out1[21] , \mul_out1[20] , \mul_out1[19] , \mul_out1[18] , 
        \mul_out1[17] , \mul_out1[16] , \mul_out1[15] , \mul_out1[14] , 
        \mul_out1[13] , \mul_out1[12] , \mul_out1[11] , \mul_out1[10] , 
        \mul_out1[9] , \mul_out1[8] , \mul_out1[7] , \mul_out1[6] , 
        \mul_out1[5] , \mul_out1[4] , \mul_out1[3] , \mul_out1[2] , 
        \mul_out1[1] , \mul_out1[0] }) );
  datapath_DW01_add_16 add_99 ( .A(f8), .B({\mul_out8[23] , \mul_out8[22] , 
        \mul_out8[21] , \mul_out8[20] , \mul_out8[19] , \mul_out8[18] , 
        \mul_out8[17] , \mul_out8[16] , \mul_out8[15] , \mul_out8[14] , 
        \mul_out8[13] , \mul_out8[12] , \mul_out8[11] , \mul_out8[10] , 
        \mul_out8[9] , \mul_out8[8] , \mul_out8[7] , \mul_out8[6] , 
        \mul_out8[5] , \mul_out8[4] , \mul_out8[3] , \mul_out8[2] , 
        \mul_out8[1] , \mul_out8[0] }), .CI(1'b0), .SUM(add_r8) );
  datapath_DW01_add_17 add_97 ( .A({n812, n804, n799, f7[20:4], n758, n765, 
        n772, n779}), .B({\mul_out7[23] , \mul_out7[22] , \mul_out7[21] , 
        \mul_out7[20] , \mul_out7[19] , \mul_out7[18] , \mul_out7[17] , 
        \mul_out7[16] , \mul_out7[15] , \mul_out7[14] , \mul_out7[13] , 
        \mul_out7[12] , \mul_out7[11] , \mul_out7[10] , \mul_out7[9] , 
        \mul_out7[8] , \mul_out7[7] , \mul_out7[6] , \mul_out7[5] , 
        \mul_out7[4] , \mul_out7[3] , \mul_out7[2] , \mul_out7[1] , 
        \mul_out7[0] }), .CI(1'b0), .SUM(add_r7) );
  datapath_DW01_add_18 add_95 ( .A({n814, n805, n800, n795, n791, n787, 
        f6[17:4], n376, n370, n372, n374}), .B({\mul_out6[23] , \mul_out6[22] , 
        \mul_out6[21] , \mul_out6[20] , \mul_out6[19] , \mul_out6[18] , 
        \mul_out6[17] , \mul_out6[16] , \mul_out6[15] , \mul_out6[14] , 
        \mul_out6[13] , \mul_out6[12] , \mul_out6[11] , \mul_out6[10] , 
        \mul_out6[9] , \mul_out6[8] , \mul_out6[7] , \mul_out6[6] , 
        \mul_out6[5] , \mul_out6[4] , \mul_out6[3] , \mul_out6[2] , 
        \mul_out6[1] , \mul_out6[0] }), .CI(1'b0), .SUM(add_r6) );
  datapath_DW01_add_19 add_93 ( .A({n507, n509, n511, n513, f5[19:4], n753, 
        n747, n749, n751}), .B({\mul_out5[23] , \mul_out5[22] , \mul_out5[21] , 
        \mul_out5[20] , \mul_out5[19] , \mul_out5[18] , \mul_out5[17] , 
        \mul_out5[16] , \mul_out5[15] , \mul_out5[14] , \mul_out5[13] , 
        \mul_out5[12] , \mul_out5[11] , \mul_out5[10] , \mul_out5[9] , 
        \mul_out5[8] , \mul_out5[7] , \mul_out5[6] , \mul_out5[5] , 
        \mul_out5[4] , \mul_out5[3] , \mul_out5[2] , \mul_out5[1] , 
        \mul_out5[0] }), .CI(1'b0), .SUM(add_r5) );
  datapath_DW01_add_20 add_91 ( .A(f4), .B({\mul_out4[23] , \mul_out4[22] , 
        \mul_out4[21] , \mul_out4[20] , \mul_out4[19] , \mul_out4[18] , 
        \mul_out4[17] , \mul_out4[16] , \mul_out4[15] , \mul_out4[14] , 
        \mul_out4[13] , \mul_out4[12] , \mul_out4[11] , \mul_out4[10] , 
        \mul_out4[9] , \mul_out4[8] , \mul_out4[7] , \mul_out4[6] , 
        \mul_out4[5] , \mul_out4[4] , \mul_out4[3] , \mul_out4[2] , 
        \mul_out4[1] , \mul_out4[0] }), .CI(1'b0), .SUM(add_r4) );
  datapath_DW01_add_21 add_89 ( .A({n476, n477, f3[21:20], n481, n483, 
        f3[17:4], n505, n499, n501, n503}), .B({\mul_out3[23] , \mul_out3[22] , 
        \mul_out3[21] , \mul_out3[20] , \mul_out3[19] , \mul_out3[18] , 
        \mul_out3[17] , \mul_out3[16] , \mul_out3[15] , \mul_out3[14] , 
        \mul_out3[13] , \mul_out3[12] , \mul_out3[11] , \mul_out3[10] , 
        \mul_out3[9] , \mul_out3[8] , \mul_out3[7] , \mul_out3[6] , 
        \mul_out3[5] , \mul_out3[4] , \mul_out3[3] , \mul_out3[2] , 
        \mul_out3[1] , \mul_out3[0] }), .CI(1'b0), .SUM(add_r3) );
  datapath_DW01_add_22 add_87 ( .A({f2[23:20], n454, n456, f2[17:4], n760, 
        n767, n774, n782}), .B({\mul_out2[23] , \mul_out2[22] , \mul_out2[21] , 
        \mul_out2[20] , \mul_out2[19] , \mul_out2[18] , \mul_out2[17] , 
        \mul_out2[16] , \mul_out2[15] , \mul_out2[14] , \mul_out2[13] , 
        \mul_out2[12] , \mul_out2[11] , \mul_out2[10] , \mul_out2[9] , 
        \mul_out2[8] , \mul_out2[7] , \mul_out2[6] , \mul_out2[5] , 
        \mul_out2[4] , \mul_out2[3] , \mul_out2[2] , \mul_out2[1] , 
        \mul_out2[0] }), .CI(1'b0), .SUM(add_r2) );
  datapath_DW01_add_23 add_85 ( .A(f1), .B({\mul_out1[23] , \mul_out1[22] , 
        \mul_out1[21] , \mul_out1[20] , \mul_out1[19] , \mul_out1[18] , 
        \mul_out1[17] , \mul_out1[16] , \mul_out1[15] , \mul_out1[14] , 
        \mul_out1[13] , \mul_out1[12] , \mul_out1[11] , \mul_out1[10] , 
        \mul_out1[9] , \mul_out1[8] , \mul_out1[7] , \mul_out1[6] , 
        \mul_out1[5] , \mul_out1[4] , \mul_out1[3] , \mul_out1[2] , 
        \mul_out1[1] , \mul_out1[0] }), .CI(1'b0), .SUM(add_r1) );
  DFF_X1 \f6_reg[2]  ( .D(n593), .CK(clk), .Q(n370), .QN(n150) );
  DFF_X1 \f6_reg[1]  ( .D(n592), .CK(clk), .Q(n372), .QN(n151) );
  DFF_X1 \f6_reg[0]  ( .D(n591), .CK(clk), .Q(n374), .QN(n152) );
  DFF_X1 \f7_reg[2]  ( .D(n569), .CK(clk), .Q(n765) );
  DFF_X1 \f7_reg[1]  ( .D(n568), .CK(clk), .Q(n772) );
  DFF_X1 \f7_reg[0]  ( .D(n567), .CK(clk), .Q(n779) );
  DFF_X1 \f8_reg[1]  ( .D(n544), .CK(clk), .Q(f8[1]), .QN(n199) );
  DFF_X1 \f8_reg[0]  ( .D(n543), .CK(clk), .Q(f8[0]), .QN(n200) );
  DFF_X1 \f4_reg[2]  ( .D(n641), .CK(clk), .Q(f4[2]), .QN(n102) );
  DFF_X1 \f4_reg[1]  ( .D(n640), .CK(clk), .Q(f4[1]), .QN(n103) );
  DFF_X1 \f4_reg[0]  ( .D(n639), .CK(clk), .Q(f4[0]), .QN(n104) );
  DFF_X1 \f8_reg[2]  ( .D(n545), .CK(clk), .Q(f8[2]), .QN(n198) );
  DFF_X1 \f1_reg[2]  ( .D(n713), .CK(clk), .Q(f1[2]), .QN(n763) );
  DFF_X1 \f1_reg[1]  ( .D(n712), .CK(clk), .Q(f1[1]), .QN(n770) );
  DFF_X1 \f1_reg[0]  ( .D(n711), .CK(clk), .Q(f1[0]), .QN(n777) );
  DFF_X1 \f5_reg[2]  ( .D(n617), .CK(clk), .Q(n747), .QN(n126) );
  DFF_X1 \f5_reg[1]  ( .D(n616), .CK(clk), .Q(n749), .QN(n127) );
  DFF_X1 \f5_reg[0]  ( .D(n615), .CK(clk), .Q(n751), .QN(n128) );
  DFF_X1 \f3_reg[2]  ( .D(n665), .CK(clk), .Q(n499), .QN(n78) );
  DFF_X1 \f3_reg[1]  ( .D(n664), .CK(clk), .Q(n501), .QN(n79) );
  DFF_X1 \f3_reg[0]  ( .D(n663), .CK(clk), .Q(n503), .QN(n80) );
  DFF_X1 \f2_reg[2]  ( .D(n689), .CK(clk), .Q(n767) );
  DFF_X1 \f2_reg[1]  ( .D(n688), .CK(clk), .Q(n774) );
  DFF_X1 \f2_reg[0]  ( .D(n687), .CK(clk), .Q(n782) );
  DFF_X1 \f3_reg[3]  ( .D(n666), .CK(clk), .Q(n505), .QN(n77) );
  DFF_X1 \f4_reg[3]  ( .D(n642), .CK(clk), .Q(f4[3]), .QN(n101) );
  DFF_X1 \f8_reg[3]  ( .D(n546), .CK(clk), .Q(f8[3]), .QN(n197) );
  DFF_X1 \f5_reg[3]  ( .D(n618), .CK(clk), .Q(n753), .QN(n125) );
  DFF_X1 \f6_reg[3]  ( .D(n594), .CK(clk), .Q(n376), .QN(n149) );
  DFF_X1 \f1_reg[3]  ( .D(n714), .CK(clk), .Q(f1[3]), .QN(n756) );
  DFF_X1 \f7_reg[3]  ( .D(n570), .CK(clk), .Q(n758) );
  DFF_X1 \f2_reg[3]  ( .D(n690), .CK(clk), .Q(n760) );
  DFF_X1 \f8_reg[4]  ( .D(n547), .CK(clk), .Q(f8[4]), .QN(n196) );
  DFF_X1 \f4_reg[4]  ( .D(n643), .CK(clk), .Q(f4[4]), .QN(n100) );
  DFF_X1 \f7_reg[4]  ( .D(n571), .CK(clk), .Q(f7[4]), .QN(n172) );
  DFF_X1 \f2_reg[4]  ( .D(n691), .CK(clk), .Q(f2[4]), .QN(n52) );
  DFF_X1 \f6_reg[4]  ( .D(n595), .CK(clk), .Q(f6[4]), .QN(n148) );
  DFF_X1 \f3_reg[4]  ( .D(n667), .CK(clk), .Q(f3[4]), .QN(n76) );
  DFF_X1 \f1_reg[4]  ( .D(n715), .CK(clk), .Q(f1[4]), .QN(n28) );
  DFF_X1 \f5_reg[4]  ( .D(n619), .CK(clk), .Q(f5[4]), .QN(n124) );
  DFF_X1 \f1_reg[5]  ( .D(n716), .CK(clk), .Q(f1[5]), .QN(n27) );
  DFF_X1 \f4_reg[5]  ( .D(n644), .CK(clk), .Q(f4[5]), .QN(n99) );
  DFF_X1 \f8_reg[5]  ( .D(n548), .CK(clk), .Q(f8[5]), .QN(n195) );
  DFF_X1 \f3_reg[5]  ( .D(n668), .CK(clk), .Q(f3[5]), .QN(n75) );
  DFF_X1 \f7_reg[5]  ( .D(n572), .CK(clk), .Q(f7[5]), .QN(n171) );
  DFF_X1 \f6_reg[5]  ( .D(n596), .CK(clk), .Q(f6[5]), .QN(n147) );
  DFF_X1 \f5_reg[5]  ( .D(n620), .CK(clk), .Q(f5[5]), .QN(n123) );
  DFF_X1 \f2_reg[5]  ( .D(n692), .CK(clk), .Q(f2[5]), .QN(n51) );
  DFF_X1 \f2_reg[6]  ( .D(n693), .CK(clk), .Q(f2[6]), .QN(n50) );
  DFF_X1 \f4_reg[6]  ( .D(n645), .CK(clk), .Q(f4[6]), .QN(n98) );
  DFF_X1 \f7_reg[6]  ( .D(n573), .CK(clk), .Q(f7[6]), .QN(n170) );
  DFF_X1 \f8_reg[6]  ( .D(n549), .CK(clk), .Q(f8[6]), .QN(n194) );
  DFF_X1 \f5_reg[6]  ( .D(n621), .CK(clk), .Q(f5[6]), .QN(n122) );
  DFF_X1 \f3_reg[6]  ( .D(n669), .CK(clk), .Q(f3[6]), .QN(n74) );
  DFF_X1 \f1_reg[6]  ( .D(n717), .CK(clk), .Q(f1[6]), .QN(n26) );
  DFF_X1 \f4_reg[7]  ( .D(n646), .CK(clk), .Q(f4[7]), .QN(n97) );
  DFF_X1 \f6_reg[6]  ( .D(n597), .CK(clk), .Q(f6[6]), .QN(n146) );
  DFF_X1 \f1_reg[7]  ( .D(n718), .CK(clk), .Q(f1[7]), .QN(n25) );
  DFF_X1 \f6_reg[7]  ( .D(n598), .CK(clk), .Q(f6[7]), .QN(n145) );
  DFF_X1 \f7_reg[7]  ( .D(n574), .CK(clk), .Q(f7[7]), .QN(n169) );
  DFF_X1 \f3_reg[8]  ( .D(n671), .CK(clk), .Q(f3[8]), .QN(n72) );
  DFF_X1 \f3_reg[7]  ( .D(n670), .CK(clk), .Q(f3[7]), .QN(n73) );
  DFF_X1 \f8_reg[7]  ( .D(n550), .CK(clk), .Q(f8[7]), .QN(n193) );
  DFF_X1 \f2_reg[7]  ( .D(n694), .CK(clk), .Q(f2[7]), .QN(n49) );
  DFF_X1 \f5_reg[7]  ( .D(n622), .CK(clk), .Q(f5[7]), .QN(n121) );
  DFF_X1 \f4_reg[8]  ( .D(n647), .CK(clk), .Q(f4[8]), .QN(n96) );
  DFF_X1 \f7_reg[8]  ( .D(n575), .CK(clk), .Q(f7[8]), .QN(n168) );
  DFF_X1 \f2_reg[8]  ( .D(n695), .CK(clk), .Q(f2[8]), .QN(n48) );
  DFF_X1 \f5_reg[8]  ( .D(n623), .CK(clk), .Q(f5[8]), .QN(n120) );
  DFF_X1 \f8_reg[8]  ( .D(n551), .CK(clk), .Q(f8[8]), .QN(n192) );
  DFF_X1 \f1_reg[9]  ( .D(n720), .CK(clk), .Q(f1[9]), .QN(n23) );
  DFF_X1 \f1_reg[8]  ( .D(n719), .CK(clk), .Q(f1[8]), .QN(n24) );
  DFF_X1 \f4_reg[9]  ( .D(n648), .CK(clk), .Q(f4[9]), .QN(n95) );
  DFF_X1 \f7_reg[9]  ( .D(n576), .CK(clk), .Q(f7[9]), .QN(n167) );
  DFF_X1 \f6_reg[8]  ( .D(n599), .CK(clk), .Q(f6[8]), .QN(n144) );
  DFF_X1 \f2_reg[9]  ( .D(n696), .CK(clk), .Q(f2[9]), .QN(n47) );
  DFF_X1 \f8_reg[9]  ( .D(n552), .CK(clk), .Q(f8[9]), .QN(n191) );
  DFF_X1 \f3_reg[9]  ( .D(n672), .CK(clk), .Q(f3[9]), .QN(n71) );
  DFF_X1 \f5_reg[9]  ( .D(n624), .CK(clk), .Q(f5[9]), .QN(n119) );
  DFF_X1 \f7_reg[10]  ( .D(n577), .CK(clk), .Q(f7[10]), .QN(n166) );
  DFF_X1 \f5_reg[10]  ( .D(n625), .CK(clk), .Q(f5[10]), .QN(n118) );
  DFF_X1 \f3_reg[10]  ( .D(n673), .CK(clk), .Q(f3[10]), .QN(n70) );
  DFF_X1 \f8_reg[10]  ( .D(n553), .CK(clk), .Q(f8[10]), .QN(n190) );
  DFF_X1 \f4_reg[10]  ( .D(n649), .CK(clk), .Q(f4[10]), .QN(n94) );
  DFF_X1 \f6_reg[9]  ( .D(n600), .CK(clk), .Q(f6[9]), .QN(n143) );
  DFF_X1 \f1_reg[10]  ( .D(n721), .CK(clk), .Q(f1[10]), .QN(n22) );
  DFF_X1 \f4_reg[11]  ( .D(n650), .CK(clk), .Q(f4[11]), .QN(n93) );
  DFF_X1 \f2_reg[10]  ( .D(n697), .CK(clk), .Q(f2[10]), .QN(n46) );
  DFF_X1 \f1_reg[12]  ( .D(n723), .CK(clk), .Q(f1[12]), .QN(n20) );
  DFF_X1 \f8_reg[11]  ( .D(n554), .CK(clk), .Q(f8[11]), .QN(n189) );
  DFF_X1 \f7_reg[11]  ( .D(n578), .CK(clk), .Q(f7[11]), .QN(n165) );
  DFF_X1 \f3_reg[11]  ( .D(n674), .CK(clk), .Q(f3[11]), .QN(n69) );
  DFF_X1 \f6_reg[10]  ( .D(n601), .CK(clk), .Q(f6[10]), .QN(n142) );
  DFF_X1 \f1_reg[11]  ( .D(n722), .CK(clk), .Q(f1[11]), .QN(n21) );
  DFF_X1 \f5_reg[11]  ( .D(n626), .CK(clk), .Q(f5[11]), .QN(n117) );
  DFF_X1 \f6_reg[12]  ( .D(n603), .CK(clk), .Q(f6[12]), .QN(n140) );
  DFF_X1 \f4_reg[19]  ( .D(n658), .CK(clk), .Q(f4[19]), .QN(n85) );
  DFF_X1 \f1_reg[19]  ( .D(n730), .CK(clk), .Q(f1[19]), .QN(n789) );
  DFF_X1 \f3_reg[20]  ( .D(n683), .CK(clk), .Q(f3[20]), .QN(n60) );
  DFF_X1 \f3_reg[21]  ( .D(n684), .CK(clk), .Q(f3[21]), .QN(n59) );
  DFF_X1 \f4_reg[21]  ( .D(n660), .CK(clk), .Q(f4[21]), .QN(n83) );
  DFF_X1 \f7_reg[19]  ( .D(n586), .CK(clk), .Q(f7[19]) );
  DFF_X1 \f7_reg[18]  ( .D(n585), .CK(clk), .Q(f7[18]) );
  DFF_X1 \f7_reg[20]  ( .D(n587), .CK(clk), .Q(f7[20]) );
  DFF_X1 \f8_reg[16]  ( .D(n559), .CK(clk), .Q(f8[16]), .QN(n184) );
  DFF_X1 \f1_reg[20]  ( .D(n731), .CK(clk), .Q(f1[20]), .QN(n793) );
  DFF_X1 \f1_reg[18]  ( .D(n729), .CK(clk), .Q(f1[18]), .QN(n785) );
  DFF_X1 \f5_reg[22]  ( .D(n637), .CK(clk), .Q(n509), .QN(n106) );
  DFF_X1 \f5_reg[18]  ( .D(n633), .CK(clk), .Q(f5[18]), .QN(n110) );
  DFF_X1 \f5_reg[17]  ( .D(n632), .CK(clk), .Q(f5[17]), .QN(n111) );
  DFF_X1 \f5_reg[19]  ( .D(n634), .CK(clk), .Q(f5[19]), .QN(n109) );
  DFF_X1 \f4_reg[23]  ( .D(n662), .CK(clk), .Q(f4[23]), .QN(n81) );
  DFF_X1 \f1_reg[23]  ( .D(n734), .CK(clk), .Q(f1[23]), .QN(n807) );
  DFF_X1 \f8_reg[19]  ( .D(n562), .CK(clk), .Q(f8[19]), .QN(n181) );
  DFF_X1 \f8_reg[21]  ( .D(n564), .CK(clk), .Q(f8[21]), .QN(n179) );
  DFF_X1 \f1_reg[16]  ( .D(n727), .CK(clk), .Q(f1[16]), .QN(n16) );
  DFF_X1 \f1_reg[17]  ( .D(n728), .CK(clk), .Q(f1[17]), .QN(n15) );
  DFF_X1 \f5_reg[23]  ( .D(n638), .CK(clk), .Q(n507), .QN(n105) );
  DFF_X1 \f8_reg[23]  ( .D(n566), .CK(clk), .Q(f8[23]), .QN(n177) );
  DFF_X1 \f5_reg[21]  ( .D(n636), .CK(clk), .Q(n511), .QN(n107) );
  DFF_X1 \f2_reg[22]  ( .D(n709), .CK(clk), .Q(f2[22]), .QN(n34) );
  DFF_X1 \f2_reg[20]  ( .D(n707), .CK(clk), .Q(f2[20]), .QN(n36) );
  DFF_X1 \f2_reg[21]  ( .D(n708), .CK(clk), .Q(f2[21]), .QN(n35) );
  DFF_X1 \f2_reg[23]  ( .D(n710), .CK(clk), .Q(f2[23]), .QN(n33) );
  DFF_X1 \f1_reg[21]  ( .D(n732), .CK(clk), .Q(f1[21]), .QN(n797) );
  DFF_X1 \f8_reg[22]  ( .D(n565), .CK(clk), .Q(f8[22]), .QN(n178) );
  DFF_X1 \f3_reg[23]  ( .D(n686), .CK(clk), .Q(n476), .QN(n57) );
  DFF_X1 \f4_reg[20]  ( .D(n659), .CK(clk), .Q(f4[20]), .QN(n84) );
  CLKBUF_X2 U3 ( .A(data_out_x[5]), .Z(n129) );
  BUF_X4 U4 ( .A(data_out_x[4]), .Z(n134) );
  BUF_X1 U5 ( .A(data_out_x[8]), .Z(n132) );
  CLKBUF_X2 U6 ( .A(data_out_x[11]), .Z(n31) );
  BUF_X1 U7 ( .A(data_out_x[10]), .Z(n133) );
  BUF_X1 U8 ( .A(data_out_x[2]), .Z(n29) );
  AND2_X1 U9 ( .A1(n299), .A2(n818), .ZN(n1) );
  AOI22_X1 U10 ( .A1(n754), .A2(n476), .B1(add_r3[23]), .B2(n156), .ZN(n12) );
  INV_X1 U11 ( .A(n12), .ZN(n686) );
  OR2_X1 U12 ( .A1(n793), .A2(n300), .ZN(n13) );
  NAND2_X1 U13 ( .A1(n13), .A2(n329), .ZN(n731) );
  BUF_X2 U14 ( .A(data_out_x[1]), .Z(n14) );
  OR2_X1 U15 ( .A1(n807), .A2(n299), .ZN(n30) );
  NAND2_X1 U16 ( .A1(n30), .A2(n326), .ZN(n734) );
  OR2_X1 U17 ( .A1(n178), .A2(n303), .ZN(n32) );
  NAND2_X1 U18 ( .A1(n32), .A2(n403), .ZN(n565) );
  OR2_X1 U19 ( .A1(n177), .A2(n303), .ZN(n53) );
  NAND2_X1 U20 ( .A1(n402), .A2(n53), .ZN(n566) );
  OR2_X1 U21 ( .A1(n84), .A2(n306), .ZN(n54) );
  NAND2_X1 U22 ( .A1(n54), .A2(n429), .ZN(n659) );
  OR2_X1 U23 ( .A1(n83), .A2(n306), .ZN(n55) );
  NAND2_X1 U24 ( .A1(n55), .A2(n428), .ZN(n660) );
  OR2_X1 U25 ( .A1(n85), .A2(n307), .ZN(n56) );
  NAND2_X1 U26 ( .A1(n56), .A2(n430), .ZN(n658) );
  OR2_X1 U27 ( .A1(n789), .A2(n300), .ZN(n130) );
  NAND2_X1 U28 ( .A1(n330), .A2(n130), .ZN(n730) );
  OR2_X1 U29 ( .A1(n81), .A2(n306), .ZN(n131) );
  NAND2_X1 U30 ( .A1(n426), .A2(n131), .ZN(n662) );
  INV_X1 U31 ( .A(n299), .ZN(n226) );
  INV_X1 U32 ( .A(n299), .ZN(n225) );
  INV_X1 U33 ( .A(n242), .ZN(n241) );
  NAND2_X1 U34 ( .A1(n315), .A2(n819), .ZN(n154) );
  NAND2_X1 U35 ( .A1(n315), .A2(n819), .ZN(n215) );
  BUF_X1 U36 ( .A(n155), .Z(n174) );
  BUF_X1 U37 ( .A(n155), .Z(n175) );
  BUF_X1 U38 ( .A(n155), .Z(n173) );
  BUF_X1 U39 ( .A(n155), .Z(n201) );
  BUF_X1 U40 ( .A(n155), .Z(n176) );
  BUF_X1 U41 ( .A(n155), .Z(n158) );
  BUF_X1 U42 ( .A(n157), .Z(n209) );
  BUF_X1 U43 ( .A(n157), .Z(n214) );
  BUF_X1 U44 ( .A(n157), .Z(n218) );
  BUF_X1 U45 ( .A(n156), .Z(n203) );
  BUF_X1 U46 ( .A(n156), .Z(n202) );
  BUF_X1 U47 ( .A(n156), .Z(n204) );
  BUF_X1 U48 ( .A(n156), .Z(n206) );
  BUF_X1 U49 ( .A(n156), .Z(n205) );
  BUF_X1 U50 ( .A(n156), .Z(n207) );
  BUF_X1 U51 ( .A(n157), .Z(n208) );
  BUF_X1 U52 ( .A(n311), .Z(n299) );
  BUF_X1 U53 ( .A(n310), .Z(n242) );
  BUF_X1 U54 ( .A(n310), .Z(n305) );
  BUF_X1 U55 ( .A(n310), .Z(n304) );
  BUF_X1 U56 ( .A(n310), .Z(n308) );
  BUF_X1 U57 ( .A(n311), .Z(n307) );
  BUF_X1 U58 ( .A(n311), .Z(n306) );
  BUF_X1 U59 ( .A(n311), .Z(n302) );
  BUF_X1 U60 ( .A(n310), .Z(n301) );
  BUF_X1 U61 ( .A(n311), .Z(n300) );
  BUF_X1 U62 ( .A(n310), .Z(n309) );
  INV_X1 U63 ( .A(n318), .ZN(n820) );
  NAND2_X1 U64 ( .A1(n323), .A2(n822), .ZN(n222) );
  INV_X1 U65 ( .A(n809), .ZN(n816) );
  NOR3_X1 U66 ( .A1(n314), .A2(n317), .A3(n318), .ZN(n315) );
  NAND2_X1 U67 ( .A1(n320), .A2(n319), .ZN(n221) );
  NAND2_X1 U68 ( .A1(n319), .A2(n821), .ZN(n318) );
  INV_X1 U69 ( .A(n320), .ZN(n821) );
  NAND2_X1 U70 ( .A1(n315), .A2(n316), .ZN(n216) );
  NAND2_X1 U71 ( .A1(n314), .A2(n820), .ZN(n217) );
  BUF_X1 U72 ( .A(n1), .Z(n156) );
  BUF_X1 U73 ( .A(n1), .Z(n155) );
  INV_X1 U74 ( .A(n316), .ZN(n819) );
  AND2_X1 U75 ( .A1(n321), .A2(n822), .ZN(n212) );
  BUF_X1 U76 ( .A(n1), .Z(n157) );
  AND2_X1 U77 ( .A1(n317), .A2(n820), .ZN(n213) );
  INV_X1 U78 ( .A(n219), .ZN(n310) );
  INV_X1 U79 ( .A(n219), .ZN(n311) );
  INV_X1 U80 ( .A(n808), .ZN(n817) );
  NOR3_X1 U81 ( .A1(n321), .A2(n323), .A3(n324), .ZN(n319) );
  NOR3_X1 U82 ( .A1(n312), .A2(addr_y[1]), .A3(n322), .ZN(n323) );
  NOR3_X1 U83 ( .A1(n312), .A2(addr_y[2]), .A3(n313), .ZN(n314) );
  NOR3_X1 U84 ( .A1(n322), .A2(addr_y[0]), .A3(n313), .ZN(n321) );
  NOR2_X1 U85 ( .A1(n322), .A2(addr_y[0]), .ZN(n320) );
  NOR2_X1 U86 ( .A1(n312), .A2(addr_y[1]), .ZN(n316) );
  NOR2_X1 U87 ( .A1(n313), .A2(addr_y[0]), .ZN(n317) );
  BUF_X1 U88 ( .A(n754), .Z(n219) );
  INV_X1 U89 ( .A(n324), .ZN(n822) );
  OAI222_X1 U90 ( .A1(n154), .A2(n41), .B1(n216), .B2(n65), .C1(n217), .C2(
        n113), .ZN(n253) );
  OAI222_X1 U91 ( .A1(n215), .A2(n40), .B1(n216), .B2(n64), .C1(n217), .C2(
        n112), .ZN(n249) );
  OAI222_X1 U92 ( .A1(n215), .A2(n52), .B1(n216), .B2(n76), .C1(n217), .C2(
        n124), .ZN(n297) );
  OAI222_X1 U93 ( .A1(n154), .A2(n51), .B1(n216), .B2(n75), .C1(n217), .C2(
        n123), .ZN(n293) );
  OAI222_X1 U94 ( .A1(n215), .A2(n50), .B1(n216), .B2(n74), .C1(n217), .C2(
        n122), .ZN(n289) );
  OAI222_X1 U95 ( .A1(n154), .A2(n49), .B1(n216), .B2(n73), .C1(n217), .C2(
        n121), .ZN(n285) );
  OAI222_X1 U96 ( .A1(n215), .A2(n48), .B1(n216), .B2(n72), .C1(n217), .C2(
        n120), .ZN(n281) );
  OAI222_X1 U97 ( .A1(n154), .A2(n47), .B1(n216), .B2(n71), .C1(n217), .C2(
        n119), .ZN(n277) );
  OAI222_X1 U98 ( .A1(n215), .A2(n46), .B1(n216), .B2(n70), .C1(n217), .C2(
        n118), .ZN(n273) );
  OAI222_X1 U99 ( .A1(n154), .A2(n45), .B1(n216), .B2(n69), .C1(n217), .C2(
        n117), .ZN(n269) );
  OAI222_X1 U100 ( .A1(n215), .A2(n44), .B1(n216), .B2(n68), .C1(n217), .C2(
        n116), .ZN(n265) );
  OAI222_X1 U101 ( .A1(n154), .A2(n43), .B1(n216), .B2(n67), .C1(n217), .C2(
        n115), .ZN(n261) );
  OAI222_X1 U102 ( .A1(n154), .A2(n42), .B1(n216), .B2(n66), .C1(n217), .C2(
        n114), .ZN(n257) );
  OAI222_X1 U103 ( .A1(n215), .A2(n39), .B1(n216), .B2(n63), .C1(n217), .C2(
        n111), .ZN(n245) );
  NAND3_X1 U104 ( .A1(clc), .A2(n818), .A3(n325), .ZN(n808) );
  NAND2_X1 U105 ( .A1(clc1), .A2(n818), .ZN(n324) );
  NAND2_X1 U106 ( .A1(n239), .A2(n240), .ZN(n524) );
  NAND2_X1 U107 ( .A1(n235), .A2(n236), .ZN(n523) );
  NAND2_X1 U108 ( .A1(n231), .A2(n232), .ZN(n522) );
  NAND2_X1 U109 ( .A1(n227), .A2(n228), .ZN(n521) );
  NAND2_X1 U110 ( .A1(n223), .A2(n224), .ZN(n520) );
  NAND2_X1 U111 ( .A1(n210), .A2(n211), .ZN(n519) );
  NAND2_X1 U112 ( .A1(n295), .A2(n296), .ZN(n538) );
  AOI221_X1 U113 ( .B1(f1[4]), .B2(n817), .C1(f[4]), .C2(n816), .A(n298), .ZN(
        n295) );
  AOI221_X1 U114 ( .B1(f8[4]), .B2(n212), .C1(f4[4]), .C2(n213), .A(n297), 
        .ZN(n296) );
  OAI22_X1 U115 ( .A1(n221), .A2(n148), .B1(n222), .B2(n172), .ZN(n298) );
  NAND2_X1 U116 ( .A1(n291), .A2(n292), .ZN(n537) );
  AOI221_X1 U117 ( .B1(f1[5]), .B2(n817), .C1(f[5]), .C2(n816), .A(n294), .ZN(
        n291) );
  AOI221_X1 U118 ( .B1(f8[5]), .B2(n212), .C1(f4[5]), .C2(n213), .A(n293), 
        .ZN(n292) );
  OAI22_X1 U119 ( .A1(n221), .A2(n147), .B1(n222), .B2(n171), .ZN(n294) );
  NAND2_X1 U120 ( .A1(n287), .A2(n288), .ZN(n536) );
  AOI221_X1 U121 ( .B1(f1[6]), .B2(n817), .C1(f[6]), .C2(n816), .A(n290), .ZN(
        n287) );
  AOI221_X1 U122 ( .B1(f8[6]), .B2(n212), .C1(f4[6]), .C2(n213), .A(n289), 
        .ZN(n288) );
  OAI22_X1 U123 ( .A1(n221), .A2(n146), .B1(n222), .B2(n170), .ZN(n290) );
  NAND2_X1 U124 ( .A1(n283), .A2(n284), .ZN(n535) );
  AOI221_X1 U125 ( .B1(f1[7]), .B2(n817), .C1(f[7]), .C2(n816), .A(n286), .ZN(
        n283) );
  AOI221_X1 U126 ( .B1(f8[7]), .B2(n212), .C1(f4[7]), .C2(n213), .A(n285), 
        .ZN(n284) );
  OAI22_X1 U127 ( .A1(n221), .A2(n145), .B1(n222), .B2(n169), .ZN(n286) );
  NAND2_X1 U128 ( .A1(n279), .A2(n280), .ZN(n534) );
  AOI221_X1 U129 ( .B1(f1[8]), .B2(n817), .C1(f[8]), .C2(n816), .A(n282), .ZN(
        n279) );
  AOI221_X1 U130 ( .B1(f8[8]), .B2(n212), .C1(f4[8]), .C2(n213), .A(n281), 
        .ZN(n280) );
  OAI22_X1 U131 ( .A1(n221), .A2(n144), .B1(n222), .B2(n168), .ZN(n282) );
  NAND2_X1 U132 ( .A1(n275), .A2(n276), .ZN(n533) );
  AOI221_X1 U133 ( .B1(f1[9]), .B2(n817), .C1(f[9]), .C2(n816), .A(n278), .ZN(
        n275) );
  AOI221_X1 U134 ( .B1(f8[9]), .B2(n212), .C1(f4[9]), .C2(n213), .A(n277), 
        .ZN(n276) );
  OAI22_X1 U135 ( .A1(n221), .A2(n143), .B1(n222), .B2(n167), .ZN(n278) );
  NAND2_X1 U136 ( .A1(n271), .A2(n272), .ZN(n532) );
  AOI221_X1 U137 ( .B1(f1[10]), .B2(n817), .C1(f[10]), .C2(n816), .A(n274), 
        .ZN(n271) );
  AOI221_X1 U138 ( .B1(f8[10]), .B2(n212), .C1(f4[10]), .C2(n213), .A(n273), 
        .ZN(n272) );
  OAI22_X1 U139 ( .A1(n221), .A2(n142), .B1(n222), .B2(n166), .ZN(n274) );
  NAND2_X1 U140 ( .A1(n267), .A2(n268), .ZN(n531) );
  AOI221_X1 U141 ( .B1(f1[11]), .B2(n817), .C1(f[11]), .C2(n816), .A(n270), 
        .ZN(n267) );
  AOI221_X1 U142 ( .B1(f8[11]), .B2(n212), .C1(f4[11]), .C2(n213), .A(n269), 
        .ZN(n268) );
  OAI22_X1 U143 ( .A1(n221), .A2(n141), .B1(n222), .B2(n165), .ZN(n270) );
  NAND2_X1 U144 ( .A1(n263), .A2(n264), .ZN(n530) );
  AOI221_X1 U145 ( .B1(f1[12]), .B2(n817), .C1(f[12]), .C2(n816), .A(n266), 
        .ZN(n263) );
  AOI221_X1 U146 ( .B1(f8[12]), .B2(n212), .C1(f4[12]), .C2(n213), .A(n265), 
        .ZN(n264) );
  OAI22_X1 U147 ( .A1(n221), .A2(n140), .B1(n222), .B2(n164), .ZN(n266) );
  NAND2_X1 U148 ( .A1(n259), .A2(n260), .ZN(n529) );
  AOI221_X1 U149 ( .B1(f1[13]), .B2(n817), .C1(f[13]), .C2(n816), .A(n262), 
        .ZN(n259) );
  AOI221_X1 U150 ( .B1(f8[13]), .B2(n212), .C1(f4[13]), .C2(n213), .A(n261), 
        .ZN(n260) );
  OAI22_X1 U151 ( .A1(n221), .A2(n139), .B1(n222), .B2(n163), .ZN(n262) );
  NAND2_X1 U152 ( .A1(n255), .A2(n256), .ZN(n528) );
  AOI221_X1 U153 ( .B1(f1[14]), .B2(n817), .C1(f[14]), .C2(n816), .A(n258), 
        .ZN(n255) );
  AOI221_X1 U154 ( .B1(f8[14]), .B2(n212), .C1(f4[14]), .C2(n213), .A(n257), 
        .ZN(n256) );
  OAI22_X1 U155 ( .A1(n221), .A2(n138), .B1(n222), .B2(n162), .ZN(n258) );
  NAND2_X1 U156 ( .A1(n251), .A2(n252), .ZN(n527) );
  AOI221_X1 U157 ( .B1(f1[15]), .B2(n817), .C1(f[15]), .C2(n816), .A(n254), 
        .ZN(n251) );
  AOI221_X1 U158 ( .B1(f8[15]), .B2(n212), .C1(f4[15]), .C2(n213), .A(n253), 
        .ZN(n252) );
  OAI22_X1 U159 ( .A1(n221), .A2(n137), .B1(n222), .B2(n161), .ZN(n254) );
  NAND2_X1 U160 ( .A1(n247), .A2(n248), .ZN(n526) );
  AOI221_X1 U161 ( .B1(f1[16]), .B2(n817), .C1(f[16]), .C2(n816), .A(n250), 
        .ZN(n247) );
  AOI221_X1 U162 ( .B1(f8[16]), .B2(n212), .C1(f4[16]), .C2(n213), .A(n249), 
        .ZN(n248) );
  OAI22_X1 U163 ( .A1(n221), .A2(n136), .B1(n222), .B2(n160), .ZN(n250) );
  NAND2_X1 U164 ( .A1(n243), .A2(n244), .ZN(n525) );
  AOI221_X1 U165 ( .B1(f1[17]), .B2(n817), .C1(f[17]), .C2(n816), .A(n246), 
        .ZN(n243) );
  AOI221_X1 U166 ( .B1(f8[17]), .B2(n212), .C1(f4[17]), .C2(n213), .A(n245), 
        .ZN(n244) );
  OAI22_X1 U167 ( .A1(n221), .A2(n135), .B1(n222), .B2(n159), .ZN(n246) );
  OR2_X1 U168 ( .A1(n183), .A2(n303), .ZN(n153) );
  NAND2_X1 U169 ( .A1(n153), .A2(n408), .ZN(n560) );
  BUF_X1 U170 ( .A(n311), .Z(n303) );
  INV_X1 U171 ( .A(n299), .ZN(n220) );
  INV_X1 U172 ( .A(n242), .ZN(n229) );
  INV_X1 U173 ( .A(n242), .ZN(n230) );
  INV_X1 U174 ( .A(n242), .ZN(n233) );
  INV_X1 U175 ( .A(n242), .ZN(n234) );
  INV_X1 U176 ( .A(n242), .ZN(n237) );
  INV_X1 U177 ( .A(n242), .ZN(n238) );
  INV_X1 U178 ( .A(addr_y[0]), .ZN(n312) );
  INV_X1 U179 ( .A(addr_y[1]), .ZN(n313) );
  INV_X1 U180 ( .A(addr_y[2]), .ZN(n322) );
  INV_X1 U181 ( .A(clc1), .ZN(n325) );
  INV_X1 U182 ( .A(clear_acc), .ZN(n818) );
  OAI21_X1 U183 ( .B1(clear_acc), .B2(n325), .A(n808), .ZN(n754) );
  NAND2_X1 U184 ( .A1(add_r1[23]), .A2(n158), .ZN(n326) );
  NAND2_X1 U185 ( .A1(add_r1[22]), .A2(n176), .ZN(n327) );
  OAI21_X1 U186 ( .B1(n802), .B2(n299), .A(n327), .ZN(n733) );
  NAND2_X1 U187 ( .A1(add_r1[21]), .A2(n201), .ZN(n328) );
  OAI21_X1 U188 ( .B1(n797), .B2(n299), .A(n328), .ZN(n732) );
  NAND2_X1 U189 ( .A1(add_r1[20]), .A2(n201), .ZN(n329) );
  NAND2_X1 U190 ( .A1(add_r1[19]), .A2(n176), .ZN(n330) );
  NAND2_X1 U191 ( .A1(add_r1[18]), .A2(n176), .ZN(n331) );
  OAI21_X1 U192 ( .B1(n785), .B2(n300), .A(n331), .ZN(n729) );
  NAND2_X1 U193 ( .A1(add_r1[17]), .A2(n176), .ZN(n332) );
  OAI21_X1 U194 ( .B1(n15), .B2(n300), .A(n332), .ZN(n728) );
  NAND2_X1 U195 ( .A1(add_r1[16]), .A2(n201), .ZN(n333) );
  OAI21_X1 U196 ( .B1(n16), .B2(n300), .A(n333), .ZN(n727) );
  NAND2_X1 U197 ( .A1(add_r1[15]), .A2(n176), .ZN(n334) );
  OAI21_X1 U198 ( .B1(n17), .B2(n300), .A(n334), .ZN(n726) );
  NAND2_X1 U199 ( .A1(add_r1[14]), .A2(n201), .ZN(n335) );
  OAI21_X1 U200 ( .B1(n18), .B2(n300), .A(n335), .ZN(n725) );
  NAND2_X1 U201 ( .A1(add_r1[13]), .A2(n201), .ZN(n336) );
  OAI21_X1 U202 ( .B1(n19), .B2(n301), .A(n336), .ZN(n724) );
  NAND2_X1 U203 ( .A1(add_r1[12]), .A2(n176), .ZN(n337) );
  OAI21_X1 U204 ( .B1(n20), .B2(n301), .A(n337), .ZN(n723) );
  NAND2_X1 U205 ( .A1(add_r1[11]), .A2(n201), .ZN(n338) );
  OAI21_X1 U206 ( .B1(n21), .B2(n301), .A(n338), .ZN(n722) );
  NAND2_X1 U207 ( .A1(add_r1[10]), .A2(n201), .ZN(n339) );
  OAI21_X1 U208 ( .B1(n22), .B2(n301), .A(n339), .ZN(n721) );
  NAND2_X1 U209 ( .A1(add_r1[9]), .A2(n176), .ZN(n340) );
  OAI21_X1 U210 ( .B1(n23), .B2(n301), .A(n340), .ZN(n720) );
  NAND2_X1 U211 ( .A1(add_r1[8]), .A2(n201), .ZN(n341) );
  OAI21_X1 U212 ( .B1(n24), .B2(n301), .A(n341), .ZN(n719) );
  NAND2_X1 U213 ( .A1(add_r1[7]), .A2(n201), .ZN(n342) );
  OAI21_X1 U214 ( .B1(n25), .B2(n301), .A(n342), .ZN(n718) );
  NAND2_X1 U215 ( .A1(add_r1[6]), .A2(n176), .ZN(n343) );
  OAI21_X1 U216 ( .B1(n26), .B2(n302), .A(n343), .ZN(n717) );
  NAND2_X1 U217 ( .A1(add_r1[5]), .A2(n176), .ZN(n344) );
  OAI21_X1 U218 ( .B1(n27), .B2(n302), .A(n344), .ZN(n716) );
  NAND2_X1 U219 ( .A1(add_r1[4]), .A2(n201), .ZN(n345) );
  OAI21_X1 U220 ( .B1(n28), .B2(n302), .A(n345), .ZN(n715) );
  NAND2_X1 U221 ( .A1(add_r1[2]), .A2(n176), .ZN(n346) );
  OAI21_X1 U222 ( .B1(n763), .B2(n302), .A(n346), .ZN(n713) );
  NAND2_X1 U223 ( .A1(add_r1[1]), .A2(n201), .ZN(n347) );
  OAI21_X1 U224 ( .B1(n770), .B2(n302), .A(n347), .ZN(n712) );
  NAND2_X1 U225 ( .A1(add_r1[0]), .A2(n176), .ZN(n348) );
  OAI21_X1 U226 ( .B1(n777), .B2(n302), .A(n348), .ZN(n711) );
  NAND2_X1 U227 ( .A1(add_r1[3]), .A2(n201), .ZN(n349) );
  OAI21_X1 U228 ( .B1(n756), .B2(n302), .A(n349), .ZN(n714) );
  AOI22_X1 U229 ( .A1(n220), .A2(n814), .B1(add_r6[23]), .B2(n205), .ZN(n350)
         );
  INV_X1 U230 ( .A(n350), .ZN(n614) );
  AOI22_X1 U231 ( .A1(n220), .A2(n805), .B1(add_r6[22]), .B2(n218), .ZN(n351)
         );
  INV_X1 U232 ( .A(n351), .ZN(n613) );
  AOI22_X1 U233 ( .A1(n220), .A2(n800), .B1(add_r6[21]), .B2(n218), .ZN(n352)
         );
  INV_X1 U234 ( .A(n352), .ZN(n612) );
  AOI22_X1 U235 ( .A1(n220), .A2(n795), .B1(add_r6[20]), .B2(n218), .ZN(n353)
         );
  INV_X1 U236 ( .A(n353), .ZN(n611) );
  AOI22_X1 U237 ( .A1(n220), .A2(n791), .B1(add_r6[19]), .B2(n218), .ZN(n354)
         );
  INV_X1 U238 ( .A(n354), .ZN(n610) );
  AOI22_X1 U239 ( .A1(n220), .A2(n787), .B1(add_r6[18]), .B2(n218), .ZN(n355)
         );
  INV_X1 U240 ( .A(n355), .ZN(n609) );
  AOI22_X1 U241 ( .A1(n220), .A2(f6[17]), .B1(add_r6[17]), .B2(n218), .ZN(n356) );
  INV_X1 U242 ( .A(n356), .ZN(n608) );
  AOI22_X1 U243 ( .A1(n220), .A2(f6[16]), .B1(add_r6[16]), .B2(n218), .ZN(n357) );
  INV_X1 U244 ( .A(n357), .ZN(n607) );
  AOI22_X1 U245 ( .A1(n220), .A2(f6[15]), .B1(add_r6[15]), .B2(n218), .ZN(n358) );
  INV_X1 U246 ( .A(n358), .ZN(n606) );
  AOI22_X1 U247 ( .A1(n220), .A2(f6[14]), .B1(add_r6[14]), .B2(n218), .ZN(n359) );
  INV_X1 U248 ( .A(n359), .ZN(n605) );
  AOI22_X1 U249 ( .A1(n220), .A2(f6[13]), .B1(add_r6[13]), .B2(n218), .ZN(n360) );
  INV_X1 U250 ( .A(n360), .ZN(n604) );
  AOI22_X1 U251 ( .A1(n220), .A2(f6[12]), .B1(add_r6[12]), .B2(n218), .ZN(n361) );
  INV_X1 U252 ( .A(n361), .ZN(n603) );
  AOI22_X1 U253 ( .A1(n225), .A2(f6[11]), .B1(add_r6[11]), .B2(n218), .ZN(n362) );
  INV_X1 U254 ( .A(n362), .ZN(n602) );
  AOI22_X1 U255 ( .A1(n225), .A2(f6[10]), .B1(add_r6[10]), .B2(n214), .ZN(n363) );
  INV_X1 U256 ( .A(n363), .ZN(n601) );
  AOI22_X1 U257 ( .A1(n225), .A2(f6[9]), .B1(add_r6[9]), .B2(n214), .ZN(n364)
         );
  INV_X1 U258 ( .A(n364), .ZN(n600) );
  AOI22_X1 U259 ( .A1(n225), .A2(f6[8]), .B1(add_r6[8]), .B2(n214), .ZN(n365)
         );
  INV_X1 U260 ( .A(n365), .ZN(n599) );
  AOI22_X1 U261 ( .A1(n225), .A2(f6[7]), .B1(add_r6[7]), .B2(n214), .ZN(n366)
         );
  INV_X1 U262 ( .A(n366), .ZN(n598) );
  AOI22_X1 U263 ( .A1(n225), .A2(f6[6]), .B1(add_r6[6]), .B2(n214), .ZN(n367)
         );
  INV_X1 U264 ( .A(n367), .ZN(n597) );
  AOI22_X1 U265 ( .A1(n225), .A2(f6[5]), .B1(add_r6[5]), .B2(n214), .ZN(n368)
         );
  INV_X1 U266 ( .A(n368), .ZN(n596) );
  AOI22_X1 U267 ( .A1(n225), .A2(f6[4]), .B1(add_r6[4]), .B2(n214), .ZN(n369)
         );
  INV_X1 U268 ( .A(n369), .ZN(n595) );
  AOI22_X1 U269 ( .A1(n225), .A2(n370), .B1(add_r6[2]), .B2(n214), .ZN(n371)
         );
  INV_X1 U270 ( .A(n371), .ZN(n593) );
  AOI22_X1 U271 ( .A1(n225), .A2(n372), .B1(add_r6[1]), .B2(n214), .ZN(n373)
         );
  INV_X1 U272 ( .A(n373), .ZN(n592) );
  AOI22_X1 U273 ( .A1(n225), .A2(n374), .B1(add_r6[0]), .B2(n214), .ZN(n375)
         );
  INV_X1 U274 ( .A(n375), .ZN(n591) );
  AOI22_X1 U275 ( .A1(n225), .A2(n376), .B1(add_r6[3]), .B2(n214), .ZN(n377)
         );
  INV_X1 U276 ( .A(n377), .ZN(n594) );
  AOI22_X1 U277 ( .A1(n226), .A2(n812), .B1(add_r7[23]), .B2(n214), .ZN(n378)
         );
  INV_X1 U278 ( .A(n378), .ZN(n590) );
  AOI22_X1 U279 ( .A1(n226), .A2(n804), .B1(add_r7[22]), .B2(n209), .ZN(n379)
         );
  INV_X1 U280 ( .A(n379), .ZN(n589) );
  AOI22_X1 U281 ( .A1(n226), .A2(n799), .B1(add_r7[21]), .B2(n209), .ZN(n380)
         );
  INV_X1 U282 ( .A(n380), .ZN(n588) );
  AOI22_X1 U283 ( .A1(n226), .A2(f7[20]), .B1(add_r7[20]), .B2(n209), .ZN(n381) );
  INV_X1 U284 ( .A(n381), .ZN(n587) );
  AOI22_X1 U285 ( .A1(n226), .A2(f7[19]), .B1(add_r7[19]), .B2(n209), .ZN(n382) );
  INV_X1 U286 ( .A(n382), .ZN(n586) );
  AOI22_X1 U287 ( .A1(n226), .A2(f7[18]), .B1(add_r7[18]), .B2(n209), .ZN(n383) );
  INV_X1 U288 ( .A(n383), .ZN(n585) );
  AOI22_X1 U289 ( .A1(n226), .A2(f7[17]), .B1(add_r7[17]), .B2(n209), .ZN(n384) );
  INV_X1 U290 ( .A(n384), .ZN(n584) );
  AOI22_X1 U291 ( .A1(n226), .A2(f7[16]), .B1(add_r7[16]), .B2(n209), .ZN(n385) );
  INV_X1 U292 ( .A(n385), .ZN(n583) );
  AOI22_X1 U293 ( .A1(n226), .A2(f7[15]), .B1(add_r7[15]), .B2(n209), .ZN(n386) );
  INV_X1 U294 ( .A(n386), .ZN(n582) );
  AOI22_X1 U295 ( .A1(n226), .A2(f7[14]), .B1(add_r7[14]), .B2(n209), .ZN(n387) );
  INV_X1 U296 ( .A(n387), .ZN(n581) );
  AOI22_X1 U297 ( .A1(n226), .A2(f7[13]), .B1(add_r7[13]), .B2(n209), .ZN(n388) );
  INV_X1 U298 ( .A(n388), .ZN(n580) );
  AOI22_X1 U299 ( .A1(n226), .A2(f7[12]), .B1(add_r7[12]), .B2(n209), .ZN(n389) );
  INV_X1 U300 ( .A(n389), .ZN(n579) );
  AOI22_X1 U301 ( .A1(n229), .A2(f7[11]), .B1(add_r7[11]), .B2(n209), .ZN(n390) );
  INV_X1 U302 ( .A(n390), .ZN(n578) );
  AOI22_X1 U303 ( .A1(n229), .A2(f7[10]), .B1(add_r7[10]), .B2(n208), .ZN(n391) );
  INV_X1 U304 ( .A(n391), .ZN(n577) );
  AOI22_X1 U305 ( .A1(n229), .A2(f7[9]), .B1(add_r7[9]), .B2(n208), .ZN(n392)
         );
  INV_X1 U306 ( .A(n392), .ZN(n576) );
  AOI22_X1 U307 ( .A1(n229), .A2(f7[8]), .B1(add_r7[8]), .B2(n208), .ZN(n393)
         );
  INV_X1 U308 ( .A(n393), .ZN(n575) );
  AOI22_X1 U309 ( .A1(n229), .A2(f7[7]), .B1(add_r7[7]), .B2(n208), .ZN(n394)
         );
  INV_X1 U310 ( .A(n394), .ZN(n574) );
  AOI22_X1 U311 ( .A1(n229), .A2(f7[6]), .B1(add_r7[6]), .B2(n208), .ZN(n395)
         );
  INV_X1 U312 ( .A(n395), .ZN(n573) );
  AOI22_X1 U313 ( .A1(n229), .A2(f7[5]), .B1(add_r7[5]), .B2(n208), .ZN(n396)
         );
  INV_X1 U314 ( .A(n396), .ZN(n572) );
  AOI22_X1 U315 ( .A1(n229), .A2(f7[4]), .B1(add_r7[4]), .B2(n208), .ZN(n397)
         );
  INV_X1 U316 ( .A(n397), .ZN(n571) );
  AOI22_X1 U317 ( .A1(n229), .A2(n765), .B1(add_r7[2]), .B2(n208), .ZN(n398)
         );
  INV_X1 U318 ( .A(n398), .ZN(n569) );
  AOI22_X1 U319 ( .A1(n229), .A2(n772), .B1(add_r7[1]), .B2(n208), .ZN(n399)
         );
  INV_X1 U320 ( .A(n399), .ZN(n568) );
  AOI22_X1 U321 ( .A1(n229), .A2(n779), .B1(add_r7[0]), .B2(n208), .ZN(n400)
         );
  INV_X1 U322 ( .A(n400), .ZN(n567) );
  AOI22_X1 U323 ( .A1(n229), .A2(n758), .B1(add_r7[3]), .B2(n208), .ZN(n401)
         );
  INV_X1 U324 ( .A(n401), .ZN(n570) );
  NAND2_X1 U325 ( .A1(add_r8[23]), .A2(n175), .ZN(n402) );
  NAND2_X1 U326 ( .A1(add_r8[22]), .A2(n175), .ZN(n403) );
  NAND2_X1 U327 ( .A1(add_r8[21]), .A2(n175), .ZN(n404) );
  OAI21_X1 U328 ( .B1(n179), .B2(n303), .A(n404), .ZN(n564) );
  NAND2_X1 U329 ( .A1(add_r8[20]), .A2(n175), .ZN(n405) );
  OAI21_X1 U330 ( .B1(n180), .B2(n303), .A(n405), .ZN(n563) );
  NAND2_X1 U331 ( .A1(add_r8[19]), .A2(n175), .ZN(n406) );
  OAI21_X1 U332 ( .B1(n181), .B2(n303), .A(n406), .ZN(n562) );
  NAND2_X1 U333 ( .A1(add_r8[18]), .A2(n175), .ZN(n407) );
  OAI21_X1 U334 ( .B1(n182), .B2(n303), .A(n407), .ZN(n561) );
  NAND2_X1 U335 ( .A1(add_r8[17]), .A2(n175), .ZN(n408) );
  NAND2_X1 U336 ( .A1(add_r8[16]), .A2(n175), .ZN(n409) );
  OAI21_X1 U337 ( .B1(n184), .B2(n304), .A(n409), .ZN(n559) );
  NAND2_X1 U338 ( .A1(add_r8[15]), .A2(n175), .ZN(n410) );
  OAI21_X1 U339 ( .B1(n185), .B2(n304), .A(n410), .ZN(n558) );
  NAND2_X1 U340 ( .A1(add_r8[14]), .A2(n175), .ZN(n411) );
  OAI21_X1 U341 ( .B1(n186), .B2(n304), .A(n411), .ZN(n557) );
  NAND2_X1 U342 ( .A1(add_r8[13]), .A2(n175), .ZN(n412) );
  OAI21_X1 U343 ( .B1(n187), .B2(n304), .A(n412), .ZN(n556) );
  NAND2_X1 U344 ( .A1(add_r8[12]), .A2(n175), .ZN(n413) );
  OAI21_X1 U345 ( .B1(n188), .B2(n304), .A(n413), .ZN(n555) );
  NAND2_X1 U346 ( .A1(add_r8[11]), .A2(n174), .ZN(n414) );
  OAI21_X1 U347 ( .B1(n189), .B2(n304), .A(n414), .ZN(n554) );
  NAND2_X1 U348 ( .A1(add_r8[10]), .A2(n174), .ZN(n415) );
  OAI21_X1 U349 ( .B1(n190), .B2(n304), .A(n415), .ZN(n553) );
  NAND2_X1 U350 ( .A1(add_r8[9]), .A2(n174), .ZN(n416) );
  OAI21_X1 U351 ( .B1(n191), .B2(n305), .A(n416), .ZN(n552) );
  NAND2_X1 U352 ( .A1(add_r8[8]), .A2(n174), .ZN(n417) );
  OAI21_X1 U353 ( .B1(n192), .B2(n305), .A(n417), .ZN(n551) );
  NAND2_X1 U354 ( .A1(add_r8[7]), .A2(n174), .ZN(n418) );
  OAI21_X1 U355 ( .B1(n193), .B2(n305), .A(n418), .ZN(n550) );
  NAND2_X1 U356 ( .A1(add_r8[6]), .A2(n174), .ZN(n419) );
  OAI21_X1 U357 ( .B1(n194), .B2(n305), .A(n419), .ZN(n549) );
  NAND2_X1 U358 ( .A1(add_r8[5]), .A2(n174), .ZN(n420) );
  OAI21_X1 U359 ( .B1(n195), .B2(n305), .A(n420), .ZN(n548) );
  NAND2_X1 U360 ( .A1(add_r8[4]), .A2(n174), .ZN(n421) );
  OAI21_X1 U361 ( .B1(n196), .B2(n305), .A(n421), .ZN(n547) );
  NAND2_X1 U362 ( .A1(add_r8[2]), .A2(n174), .ZN(n422) );
  OAI21_X1 U363 ( .B1(n198), .B2(n305), .A(n422), .ZN(n545) );
  NAND2_X1 U364 ( .A1(add_r8[1]), .A2(n174), .ZN(n423) );
  OAI21_X1 U365 ( .B1(n199), .B2(n306), .A(n423), .ZN(n544) );
  NAND2_X1 U366 ( .A1(add_r8[0]), .A2(n174), .ZN(n424) );
  OAI21_X1 U367 ( .B1(n200), .B2(n306), .A(n424), .ZN(n543) );
  NAND2_X1 U368 ( .A1(add_r8[3]), .A2(n174), .ZN(n425) );
  OAI21_X1 U369 ( .B1(n197), .B2(n306), .A(n425), .ZN(n546) );
  NAND2_X1 U370 ( .A1(add_r4[23]), .A2(n173), .ZN(n426) );
  NAND2_X1 U371 ( .A1(add_r4[22]), .A2(n173), .ZN(n427) );
  OAI21_X1 U372 ( .B1(n82), .B2(n306), .A(n427), .ZN(n661) );
  NAND2_X1 U373 ( .A1(add_r4[21]), .A2(n173), .ZN(n428) );
  NAND2_X1 U374 ( .A1(add_r4[20]), .A2(n176), .ZN(n429) );
  NAND2_X1 U375 ( .A1(add_r4[19]), .A2(n173), .ZN(n430) );
  NAND2_X1 U376 ( .A1(add_r4[18]), .A2(n173), .ZN(n431) );
  OAI21_X1 U377 ( .B1(n86), .B2(n307), .A(n431), .ZN(n657) );
  NAND2_X1 U378 ( .A1(add_r4[17]), .A2(n173), .ZN(n432) );
  OAI21_X1 U379 ( .B1(n87), .B2(n307), .A(n432), .ZN(n656) );
  NAND2_X1 U380 ( .A1(add_r4[16]), .A2(n173), .ZN(n433) );
  OAI21_X1 U381 ( .B1(n88), .B2(n307), .A(n433), .ZN(n655) );
  NAND2_X1 U382 ( .A1(add_r4[15]), .A2(n173), .ZN(n434) );
  OAI21_X1 U383 ( .B1(n89), .B2(n307), .A(n434), .ZN(n654) );
  NAND2_X1 U384 ( .A1(add_r4[14]), .A2(n173), .ZN(n435) );
  OAI21_X1 U385 ( .B1(n90), .B2(n307), .A(n435), .ZN(n653) );
  NAND2_X1 U386 ( .A1(add_r4[13]), .A2(n173), .ZN(n436) );
  OAI21_X1 U387 ( .B1(n91), .B2(n307), .A(n436), .ZN(n652) );
  NAND2_X1 U388 ( .A1(add_r4[12]), .A2(n173), .ZN(n437) );
  OAI21_X1 U389 ( .B1(n92), .B2(n308), .A(n437), .ZN(n651) );
  NAND2_X1 U390 ( .A1(add_r4[11]), .A2(n173), .ZN(n438) );
  OAI21_X1 U391 ( .B1(n93), .B2(n308), .A(n438), .ZN(n650) );
  NAND2_X1 U392 ( .A1(add_r4[10]), .A2(n158), .ZN(n439) );
  OAI21_X1 U393 ( .B1(n94), .B2(n308), .A(n439), .ZN(n649) );
  NAND2_X1 U394 ( .A1(add_r4[9]), .A2(n158), .ZN(n440) );
  OAI21_X1 U395 ( .B1(n95), .B2(n308), .A(n440), .ZN(n648) );
  NAND2_X1 U396 ( .A1(add_r4[8]), .A2(n158), .ZN(n441) );
  OAI21_X1 U397 ( .B1(n96), .B2(n308), .A(n441), .ZN(n647) );
  NAND2_X1 U398 ( .A1(add_r4[7]), .A2(n158), .ZN(n442) );
  OAI21_X1 U399 ( .B1(n97), .B2(n308), .A(n442), .ZN(n646) );
  NAND2_X1 U400 ( .A1(add_r4[6]), .A2(n158), .ZN(n443) );
  OAI21_X1 U401 ( .B1(n98), .B2(n308), .A(n443), .ZN(n645) );
  NAND2_X1 U402 ( .A1(add_r4[5]), .A2(n158), .ZN(n444) );
  OAI21_X1 U403 ( .B1(n99), .B2(n309), .A(n444), .ZN(n644) );
  NAND2_X1 U404 ( .A1(add_r4[4]), .A2(n158), .ZN(n445) );
  OAI21_X1 U405 ( .B1(n100), .B2(n309), .A(n445), .ZN(n643) );
  NAND2_X1 U406 ( .A1(add_r4[2]), .A2(n158), .ZN(n446) );
  OAI21_X1 U407 ( .B1(n102), .B2(n309), .A(n446), .ZN(n641) );
  NAND2_X1 U408 ( .A1(add_r4[1]), .A2(n158), .ZN(n447) );
  OAI21_X1 U409 ( .B1(n103), .B2(n309), .A(n447), .ZN(n640) );
  NAND2_X1 U410 ( .A1(add_r4[0]), .A2(n158), .ZN(n448) );
  OAI21_X1 U411 ( .B1(n104), .B2(n309), .A(n448), .ZN(n639) );
  NAND2_X1 U412 ( .A1(add_r4[3]), .A2(n158), .ZN(n449) );
  OAI21_X1 U413 ( .B1(n101), .B2(n309), .A(n449), .ZN(n642) );
  AOI22_X1 U414 ( .A1(n230), .A2(f2[23]), .B1(add_r2[23]), .B2(n208), .ZN(n450) );
  INV_X1 U415 ( .A(n450), .ZN(n710) );
  AOI22_X1 U416 ( .A1(n230), .A2(f2[22]), .B1(add_r2[22]), .B2(n207), .ZN(n451) );
  INV_X1 U417 ( .A(n451), .ZN(n709) );
  AOI22_X1 U418 ( .A1(n230), .A2(f2[21]), .B1(add_r2[21]), .B2(n207), .ZN(n452) );
  INV_X1 U419 ( .A(n452), .ZN(n708) );
  AOI22_X1 U420 ( .A1(n230), .A2(f2[20]), .B1(add_r2[20]), .B2(n207), .ZN(n453) );
  INV_X1 U421 ( .A(n453), .ZN(n707) );
  AOI22_X1 U422 ( .A1(n230), .A2(n454), .B1(add_r2[19]), .B2(n207), .ZN(n455)
         );
  INV_X1 U423 ( .A(n455), .ZN(n706) );
  AOI22_X1 U424 ( .A1(n230), .A2(n456), .B1(add_r2[18]), .B2(n207), .ZN(n457)
         );
  INV_X1 U425 ( .A(n457), .ZN(n705) );
  AOI22_X1 U426 ( .A1(n230), .A2(f2[17]), .B1(add_r2[17]), .B2(n207), .ZN(n458) );
  INV_X1 U427 ( .A(n458), .ZN(n704) );
  AOI22_X1 U428 ( .A1(n230), .A2(f2[16]), .B1(add_r2[16]), .B2(n207), .ZN(n459) );
  INV_X1 U429 ( .A(n459), .ZN(n703) );
  AOI22_X1 U430 ( .A1(n230), .A2(f2[15]), .B1(add_r2[15]), .B2(n207), .ZN(n460) );
  INV_X1 U431 ( .A(n460), .ZN(n702) );
  AOI22_X1 U432 ( .A1(n230), .A2(f2[14]), .B1(add_r2[14]), .B2(n207), .ZN(n461) );
  INV_X1 U433 ( .A(n461), .ZN(n701) );
  AOI22_X1 U434 ( .A1(n230), .A2(f2[13]), .B1(add_r2[13]), .B2(n207), .ZN(n462) );
  INV_X1 U435 ( .A(n462), .ZN(n700) );
  AOI22_X1 U436 ( .A1(n230), .A2(f2[12]), .B1(add_r2[12]), .B2(n207), .ZN(n463) );
  INV_X1 U437 ( .A(n463), .ZN(n699) );
  AOI22_X1 U438 ( .A1(n233), .A2(f2[11]), .B1(add_r2[11]), .B2(n205), .ZN(n464) );
  INV_X1 U439 ( .A(n464), .ZN(n698) );
  AOI22_X1 U440 ( .A1(n233), .A2(f2[10]), .B1(add_r2[10]), .B2(n206), .ZN(n465) );
  INV_X1 U441 ( .A(n465), .ZN(n697) );
  AOI22_X1 U442 ( .A1(n233), .A2(f2[9]), .B1(add_r2[9]), .B2(n206), .ZN(n466)
         );
  INV_X1 U443 ( .A(n466), .ZN(n696) );
  AOI22_X1 U444 ( .A1(n233), .A2(f2[8]), .B1(add_r2[8]), .B2(n206), .ZN(n467)
         );
  INV_X1 U445 ( .A(n467), .ZN(n695) );
  AOI22_X1 U446 ( .A1(n233), .A2(f2[7]), .B1(add_r2[7]), .B2(n206), .ZN(n468)
         );
  INV_X1 U447 ( .A(n468), .ZN(n694) );
  AOI22_X1 U448 ( .A1(n233), .A2(f2[6]), .B1(add_r2[6]), .B2(n206), .ZN(n469)
         );
  INV_X1 U449 ( .A(n469), .ZN(n693) );
  AOI22_X1 U450 ( .A1(n233), .A2(f2[5]), .B1(add_r2[5]), .B2(n206), .ZN(n470)
         );
  INV_X1 U451 ( .A(n470), .ZN(n692) );
  AOI22_X1 U452 ( .A1(n233), .A2(f2[4]), .B1(add_r2[4]), .B2(n206), .ZN(n471)
         );
  INV_X1 U453 ( .A(n471), .ZN(n691) );
  AOI22_X1 U454 ( .A1(n233), .A2(n767), .B1(add_r2[2]), .B2(n206), .ZN(n472)
         );
  INV_X1 U455 ( .A(n472), .ZN(n689) );
  AOI22_X1 U456 ( .A1(n233), .A2(n774), .B1(add_r2[1]), .B2(n206), .ZN(n473)
         );
  INV_X1 U457 ( .A(n473), .ZN(n688) );
  AOI22_X1 U458 ( .A1(n233), .A2(n782), .B1(add_r2[0]), .B2(n206), .ZN(n474)
         );
  INV_X1 U459 ( .A(n474), .ZN(n687) );
  AOI22_X1 U460 ( .A1(n233), .A2(n760), .B1(add_r2[3]), .B2(n206), .ZN(n475)
         );
  INV_X1 U461 ( .A(n475), .ZN(n690) );
  AOI22_X1 U462 ( .A1(n234), .A2(n477), .B1(add_r3[22]), .B2(n202), .ZN(n478)
         );
  INV_X1 U463 ( .A(n478), .ZN(n685) );
  AOI22_X1 U464 ( .A1(n234), .A2(f3[21]), .B1(add_r3[21]), .B2(n202), .ZN(n479) );
  INV_X1 U465 ( .A(n479), .ZN(n684) );
  AOI22_X1 U466 ( .A1(n234), .A2(f3[20]), .B1(add_r3[20]), .B2(n205), .ZN(n480) );
  INV_X1 U467 ( .A(n480), .ZN(n683) );
  AOI22_X1 U468 ( .A1(n234), .A2(n481), .B1(add_r3[19]), .B2(n205), .ZN(n482)
         );
  INV_X1 U469 ( .A(n482), .ZN(n682) );
  AOI22_X1 U470 ( .A1(n234), .A2(n483), .B1(add_r3[18]), .B2(n202), .ZN(n484)
         );
  INV_X1 U471 ( .A(n484), .ZN(n681) );
  AOI22_X1 U472 ( .A1(n234), .A2(f3[17]), .B1(add_r3[17]), .B2(n204), .ZN(n485) );
  INV_X1 U473 ( .A(n485), .ZN(n680) );
  AOI22_X1 U474 ( .A1(n234), .A2(f3[16]), .B1(add_r3[16]), .B2(n202), .ZN(n486) );
  INV_X1 U475 ( .A(n486), .ZN(n679) );
  AOI22_X1 U476 ( .A1(n234), .A2(f3[15]), .B1(add_r3[15]), .B2(n202), .ZN(n487) );
  INV_X1 U477 ( .A(n487), .ZN(n678) );
  AOI22_X1 U478 ( .A1(n234), .A2(f3[14]), .B1(add_r3[14]), .B2(n204), .ZN(n488) );
  INV_X1 U479 ( .A(n488), .ZN(n677) );
  AOI22_X1 U480 ( .A1(n234), .A2(f3[13]), .B1(add_r3[13]), .B2(n203), .ZN(n489) );
  INV_X1 U481 ( .A(n489), .ZN(n676) );
  AOI22_X1 U482 ( .A1(n234), .A2(f3[12]), .B1(add_r3[12]), .B2(n202), .ZN(n490) );
  INV_X1 U483 ( .A(n490), .ZN(n675) );
  AOI22_X1 U484 ( .A1(n237), .A2(f3[11]), .B1(add_r3[11]), .B2(n203), .ZN(n491) );
  INV_X1 U485 ( .A(n491), .ZN(n674) );
  AOI22_X1 U486 ( .A1(n237), .A2(f3[10]), .B1(add_r3[10]), .B2(n202), .ZN(n492) );
  INV_X1 U487 ( .A(n492), .ZN(n673) );
  AOI22_X1 U488 ( .A1(n237), .A2(f3[9]), .B1(add_r3[9]), .B2(n204), .ZN(n493)
         );
  INV_X1 U489 ( .A(n493), .ZN(n672) );
  AOI22_X1 U490 ( .A1(n237), .A2(f3[8]), .B1(add_r3[8]), .B2(n203), .ZN(n494)
         );
  INV_X1 U491 ( .A(n494), .ZN(n671) );
  AOI22_X1 U492 ( .A1(n237), .A2(f3[7]), .B1(add_r3[7]), .B2(n202), .ZN(n495)
         );
  INV_X1 U493 ( .A(n495), .ZN(n670) );
  AOI22_X1 U494 ( .A1(n237), .A2(f3[6]), .B1(add_r3[6]), .B2(n203), .ZN(n496)
         );
  INV_X1 U495 ( .A(n496), .ZN(n669) );
  AOI22_X1 U496 ( .A1(n237), .A2(f3[5]), .B1(add_r3[5]), .B2(n203), .ZN(n497)
         );
  INV_X1 U497 ( .A(n497), .ZN(n668) );
  AOI22_X1 U498 ( .A1(n237), .A2(f3[4]), .B1(add_r3[4]), .B2(n202), .ZN(n498)
         );
  INV_X1 U499 ( .A(n498), .ZN(n667) );
  AOI22_X1 U500 ( .A1(n237), .A2(n499), .B1(add_r3[2]), .B2(n202), .ZN(n500)
         );
  INV_X1 U501 ( .A(n500), .ZN(n665) );
  AOI22_X1 U502 ( .A1(n237), .A2(n501), .B1(add_r3[1]), .B2(n203), .ZN(n502)
         );
  INV_X1 U503 ( .A(n502), .ZN(n664) );
  AOI22_X1 U504 ( .A1(n237), .A2(n503), .B1(add_r3[0]), .B2(n202), .ZN(n504)
         );
  INV_X1 U505 ( .A(n504), .ZN(n663) );
  AOI22_X1 U506 ( .A1(n237), .A2(n505), .B1(add_r3[3]), .B2(n202), .ZN(n506)
         );
  INV_X1 U507 ( .A(n506), .ZN(n666) );
  AOI22_X1 U508 ( .A1(n238), .A2(n507), .B1(add_r5[23]), .B2(n203), .ZN(n508)
         );
  INV_X1 U509 ( .A(n508), .ZN(n638) );
  AOI22_X1 U510 ( .A1(n238), .A2(n509), .B1(add_r5[22]), .B2(n204), .ZN(n510)
         );
  INV_X1 U511 ( .A(n510), .ZN(n637) );
  AOI22_X1 U512 ( .A1(n238), .A2(n511), .B1(add_r5[21]), .B2(n204), .ZN(n512)
         );
  INV_X1 U513 ( .A(n512), .ZN(n636) );
  AOI22_X1 U514 ( .A1(n238), .A2(n513), .B1(add_r5[20]), .B2(n203), .ZN(n514)
         );
  INV_X1 U515 ( .A(n514), .ZN(n635) );
  AOI22_X1 U516 ( .A1(n238), .A2(f5[19]), .B1(add_r5[19]), .B2(n205), .ZN(n515) );
  INV_X1 U517 ( .A(n515), .ZN(n634) );
  AOI22_X1 U518 ( .A1(n238), .A2(f5[18]), .B1(add_r5[18]), .B2(n203), .ZN(n516) );
  INV_X1 U519 ( .A(n516), .ZN(n633) );
  AOI22_X1 U520 ( .A1(n238), .A2(f5[17]), .B1(add_r5[17]), .B2(n203), .ZN(n517) );
  INV_X1 U521 ( .A(n517), .ZN(n632) );
  AOI22_X1 U522 ( .A1(n238), .A2(f5[16]), .B1(add_r5[16]), .B2(n205), .ZN(n518) );
  INV_X1 U523 ( .A(n518), .ZN(n631) );
  AOI22_X1 U524 ( .A1(n238), .A2(f5[15]), .B1(add_r5[15]), .B2(n203), .ZN(n735) );
  INV_X1 U525 ( .A(n735), .ZN(n630) );
  AOI22_X1 U526 ( .A1(n238), .A2(f5[14]), .B1(add_r5[14]), .B2(n205), .ZN(n736) );
  INV_X1 U527 ( .A(n736), .ZN(n629) );
  AOI22_X1 U528 ( .A1(n238), .A2(f5[13]), .B1(add_r5[13]), .B2(n205), .ZN(n737) );
  INV_X1 U529 ( .A(n737), .ZN(n628) );
  AOI22_X1 U530 ( .A1(n238), .A2(f5[12]), .B1(add_r5[12]), .B2(n203), .ZN(n738) );
  INV_X1 U531 ( .A(n738), .ZN(n627) );
  AOI22_X1 U532 ( .A1(n241), .A2(f5[11]), .B1(add_r5[11]), .B2(n204), .ZN(n739) );
  INV_X1 U533 ( .A(n739), .ZN(n626) );
  AOI22_X1 U534 ( .A1(n241), .A2(f5[10]), .B1(add_r5[10]), .B2(n205), .ZN(n740) );
  INV_X1 U535 ( .A(n740), .ZN(n625) );
  AOI22_X1 U536 ( .A1(n241), .A2(f5[9]), .B1(add_r5[9]), .B2(n204), .ZN(n741)
         );
  INV_X1 U537 ( .A(n741), .ZN(n624) );
  AOI22_X1 U538 ( .A1(n241), .A2(f5[8]), .B1(add_r5[8]), .B2(n204), .ZN(n742)
         );
  INV_X1 U539 ( .A(n742), .ZN(n623) );
  AOI22_X1 U540 ( .A1(n241), .A2(f5[7]), .B1(add_r5[7]), .B2(n205), .ZN(n743)
         );
  INV_X1 U541 ( .A(n743), .ZN(n622) );
  AOI22_X1 U542 ( .A1(n241), .A2(f5[6]), .B1(add_r5[6]), .B2(n204), .ZN(n744)
         );
  INV_X1 U543 ( .A(n744), .ZN(n621) );
  AOI22_X1 U544 ( .A1(n241), .A2(f5[5]), .B1(add_r5[5]), .B2(n204), .ZN(n745)
         );
  INV_X1 U545 ( .A(n745), .ZN(n620) );
  AOI22_X1 U546 ( .A1(n241), .A2(f5[4]), .B1(add_r5[4]), .B2(n205), .ZN(n746)
         );
  INV_X1 U547 ( .A(n746), .ZN(n619) );
  AOI22_X1 U548 ( .A1(n241), .A2(n747), .B1(add_r5[2]), .B2(n204), .ZN(n748)
         );
  INV_X1 U549 ( .A(n748), .ZN(n617) );
  AOI22_X1 U550 ( .A1(n241), .A2(n749), .B1(add_r5[1]), .B2(n206), .ZN(n750)
         );
  INV_X1 U551 ( .A(n750), .ZN(n616) );
  AOI22_X1 U552 ( .A1(n241), .A2(n751), .B1(add_r5[0]), .B2(n205), .ZN(n752)
         );
  INV_X1 U553 ( .A(n752), .ZN(n615) );
  AOI22_X1 U554 ( .A1(n241), .A2(n753), .B1(add_r5[3]), .B2(n207), .ZN(n755)
         );
  INV_X1 U555 ( .A(n755), .ZN(n618) );
  INV_X1 U556 ( .A(n222), .ZN(n811) );
  NAND2_X1 U557 ( .A1(n808), .A2(n324), .ZN(n809) );
  OAI222_X1 U558 ( .A1(n809), .A2(n8), .B1(n808), .B2(n756), .C1(n221), .C2(
        n149), .ZN(n757) );
  AOI221_X1 U559 ( .B1(n758), .B2(n811), .C1(f8[3]), .C2(n212), .A(n757), .ZN(
        n762) );
  INV_X1 U560 ( .A(n215), .ZN(n781) );
  OAI22_X1 U561 ( .A1(n217), .A2(n125), .B1(n216), .B2(n77), .ZN(n759) );
  AOI221_X1 U562 ( .B1(f4[3]), .B2(n213), .C1(n760), .C2(n781), .A(n759), .ZN(
        n761) );
  NAND2_X1 U563 ( .A1(n762), .A2(n761), .ZN(n539) );
  OAI222_X1 U564 ( .A1(n809), .A2(n9), .B1(n808), .B2(n763), .C1(n221), .C2(
        n150), .ZN(n764) );
  AOI221_X1 U565 ( .B1(n765), .B2(n811), .C1(f8[2]), .C2(n212), .A(n764), .ZN(
        n769) );
  OAI22_X1 U566 ( .A1(n217), .A2(n126), .B1(n216), .B2(n78), .ZN(n766) );
  AOI221_X1 U567 ( .B1(f4[2]), .B2(n213), .C1(n767), .C2(n781), .A(n766), .ZN(
        n768) );
  NAND2_X1 U568 ( .A1(n769), .A2(n768), .ZN(n540) );
  OAI222_X1 U569 ( .A1(n809), .A2(n10), .B1(n808), .B2(n770), .C1(n221), .C2(
        n151), .ZN(n771) );
  AOI221_X1 U570 ( .B1(n772), .B2(n811), .C1(f8[1]), .C2(n212), .A(n771), .ZN(
        n776) );
  OAI22_X1 U571 ( .A1(n217), .A2(n127), .B1(n216), .B2(n79), .ZN(n773) );
  AOI221_X1 U572 ( .B1(f4[1]), .B2(n213), .C1(n774), .C2(n781), .A(n773), .ZN(
        n775) );
  NAND2_X1 U573 ( .A1(n776), .A2(n775), .ZN(n541) );
  OAI222_X1 U574 ( .A1(n809), .A2(n11), .B1(n808), .B2(n777), .C1(n221), .C2(
        n152), .ZN(n778) );
  AOI221_X1 U575 ( .B1(n779), .B2(n811), .C1(f8[0]), .C2(n212), .A(n778), .ZN(
        n784) );
  OAI22_X1 U576 ( .A1(n217), .A2(n128), .B1(n216), .B2(n80), .ZN(n780) );
  AOI221_X1 U577 ( .B1(f4[0]), .B2(n213), .C1(n782), .C2(n781), .A(n780), .ZN(
        n783) );
  NAND2_X1 U578 ( .A1(n784), .A2(n783), .ZN(n542) );
  INV_X1 U579 ( .A(n221), .ZN(n813) );
  OAI22_X1 U580 ( .A1(n809), .A2(n2), .B1(n808), .B2(n785), .ZN(n786) );
  AOI221_X1 U581 ( .B1(n787), .B2(n813), .C1(f7[18]), .C2(n811), .A(n786), 
        .ZN(n239) );
  OAI222_X1 U582 ( .A1(n216), .A2(n62), .B1(n154), .B2(n38), .C1(n217), .C2(
        n110), .ZN(n788) );
  AOI221_X1 U583 ( .B1(f4[18]), .B2(n213), .C1(f8[18]), .C2(n212), .A(n788), 
        .ZN(n240) );
  OAI22_X1 U584 ( .A1(n809), .A2(n3), .B1(n808), .B2(n789), .ZN(n790) );
  AOI221_X1 U585 ( .B1(n791), .B2(n813), .C1(f7[19]), .C2(n811), .A(n790), 
        .ZN(n235) );
  OAI222_X1 U586 ( .A1(n216), .A2(n61), .B1(n154), .B2(n37), .C1(n217), .C2(
        n109), .ZN(n792) );
  AOI221_X1 U587 ( .B1(f4[19]), .B2(n213), .C1(f8[19]), .C2(n212), .A(n792), 
        .ZN(n236) );
  OAI22_X1 U588 ( .A1(n809), .A2(n4), .B1(n808), .B2(n793), .ZN(n794) );
  AOI221_X1 U589 ( .B1(n795), .B2(n813), .C1(f7[20]), .C2(n811), .A(n794), 
        .ZN(n231) );
  OAI222_X1 U590 ( .A1(n216), .A2(n60), .B1(n215), .B2(n36), .C1(n217), .C2(
        n108), .ZN(n796) );
  AOI221_X1 U591 ( .B1(f4[20]), .B2(n213), .C1(f8[20]), .C2(n212), .A(n796), 
        .ZN(n232) );
  OAI22_X1 U592 ( .A1(n809), .A2(n5), .B1(n808), .B2(n797), .ZN(n798) );
  AOI221_X1 U593 ( .B1(n800), .B2(n813), .C1(n799), .C2(n811), .A(n798), .ZN(
        n227) );
  OAI222_X1 U594 ( .A1(n216), .A2(n59), .B1(n154), .B2(n35), .C1(n217), .C2(
        n107), .ZN(n801) );
  AOI221_X1 U595 ( .B1(f4[21]), .B2(n213), .C1(f8[21]), .C2(n212), .A(n801), 
        .ZN(n228) );
  OAI22_X1 U596 ( .A1(n809), .A2(n6), .B1(n808), .B2(n802), .ZN(n803) );
  AOI221_X1 U597 ( .B1(n805), .B2(n813), .C1(n804), .C2(n811), .A(n803), .ZN(
        n223) );
  OAI222_X1 U598 ( .A1(n216), .A2(n58), .B1(n215), .B2(n34), .C1(n217), .C2(
        n106), .ZN(n806) );
  AOI221_X1 U599 ( .B1(f4[22]), .B2(n213), .C1(f8[22]), .C2(n212), .A(n806), 
        .ZN(n224) );
  OAI22_X1 U600 ( .A1(n809), .A2(n7), .B1(n808), .B2(n807), .ZN(n810) );
  AOI221_X1 U601 ( .B1(n814), .B2(n813), .C1(n812), .C2(n811), .A(n810), .ZN(
        n210) );
  OAI222_X1 U602 ( .A1(n216), .A2(n57), .B1(n154), .B2(n33), .C1(n217), .C2(
        n105), .ZN(n815) );
  AOI221_X1 U603 ( .B1(f4[23]), .B2(n213), .C1(f8[23]), .C2(n212), .A(n815), 
        .ZN(n211) );
endmodule


module ctrlpath ( clk, reset, start, addr_x, wr_en_x, addr_a1, addr_a2, 
        addr_a3, addr_a4, addr_a5, addr_a6, addr_a7, addr_a8, wr_en_a1, 
        wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6, wr_en_a7, wr_en_a8, 
        clear_acc, clc, clc1, addr_y, wr_en_y, done, loadMatrix, loadVector );
  output [2:0] addr_x;
  output [2:0] addr_a1;
  output [2:0] addr_a2;
  output [2:0] addr_a3;
  output [2:0] addr_a4;
  output [2:0] addr_a5;
  output [2:0] addr_a6;
  output [2:0] addr_a7;
  output [2:0] addr_a8;
  output [2:0] addr_y;
  input clk, reset, start, loadMatrix, loadVector;
  output wr_en_x, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6,
         wr_en_a7, wr_en_a8, clear_acc, clc, clc1, wr_en_y, done;
  wire   N32, N33, N34, N35, N37, N45, N46, N56, N57, N67, N68, N78, N79, N89,
         N90, N100, N101, N111, N112, N122, N123, N131, N132, N133, N141, N142,
         N143, N146, N147, N148, n76, n79, n80, n81, n83, n84, n85, n86, n87,
         n88, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n111, n112, n113, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39;
  wire   [4:0] state;

  DFF_X1 \state_reg[3]  ( .D(N35), .CK(clk), .Q(state[3]) );
  DFF_X1 done_reg ( .D(N37), .CK(clk), .Q(done) );
  DFF_X1 \addr_x_reg[0]  ( .D(N131), .CK(clk), .Q(addr_x[0]) );
  DFF_X1 \addr_x_reg[1]  ( .D(N132), .CK(clk), .Q(addr_x[1]) );
  DFF_X1 clear_acc_reg ( .D(N146), .CK(clk), .Q(clear_acc) );
  DFF_X1 clc_reg ( .D(N147), .CK(clk), .Q(clc) );
  DFF_X1 clc1_reg ( .D(N148), .CK(clk), .Q(clc1) );
  NAND3_X1 U201 ( .A1(n127), .A2(n97), .A3(addr_a5[0]), .ZN(n129) );
  NAND3_X1 U202 ( .A1(n133), .A2(n121), .A3(n134), .ZN(n132) );
  NAND3_X1 U203 ( .A1(n137), .A2(n94), .A3(addr_a4[0]), .ZN(n139) );
  NAND3_X1 U204 ( .A1(n120), .A2(n119), .A3(n142), .ZN(n141) );
  NAND3_X1 U205 ( .A1(n145), .A2(n91), .A3(addr_a3[0]), .ZN(n147) );
  NAND3_X1 U206 ( .A1(n142), .A2(n120), .A3(n27), .ZN(n149) );
  NAND3_X1 U207 ( .A1(n153), .A2(n87), .A3(addr_a2[0]), .ZN(n155) );
  NAND3_X1 U208 ( .A1(n119), .A2(n118), .A3(n142), .ZN(n157) );
  NAND3_X1 U209 ( .A1(n162), .A2(n84), .A3(addr_a1[0]), .ZN(n164) );
  NAND3_X1 U210 ( .A1(n133), .A2(n167), .A3(n134), .ZN(n166) );
  NAND3_X1 U211 ( .A1(n178), .A2(n179), .A3(n31), .ZN(n175) );
  NAND3_X1 U212 ( .A1(addr_a8[1]), .A2(addr_a8[0]), .A3(addr_a8[2]), .ZN(n170)
         );
  NAND3_X1 U213 ( .A1(addr_a7[1]), .A2(addr_a7[0]), .A3(addr_a7[2]), .ZN(n195)
         );
  NAND3_X1 U214 ( .A1(addr_y[0]), .A2(n112), .A3(n216), .ZN(n218) );
  NAND3_X1 U215 ( .A1(n219), .A2(n30), .A3(addr_y[0]), .ZN(n220) );
  NAND3_X1 U216 ( .A1(addr_x[0]), .A2(n224), .A3(addr_x[1]), .ZN(n223) );
  NAND3_X1 U217 ( .A1(n228), .A2(n106), .A3(addr_a8[0]), .ZN(n230) );
  NAND3_X1 U218 ( .A1(n233), .A2(n172), .A3(n134), .ZN(n232) );
  NAND3_X1 U219 ( .A1(n236), .A2(n103), .A3(addr_a7[0]), .ZN(n238) );
  NAND3_X1 U220 ( .A1(n233), .A2(n173), .A3(n134), .ZN(n240) );
  NAND3_X1 U221 ( .A1(n123), .A2(n100), .A3(addr_a6[0]), .ZN(n244) );
  NAND3_X1 U222 ( .A1(n22), .A2(n158), .A3(n28), .ZN(n245) );
  NAND3_X1 U223 ( .A1(n119), .A2(n118), .A3(n120), .ZN(n246) );
  NAND3_X1 U224 ( .A1(addr_x[1]), .A2(addr_x[0]), .A3(addr_x[2]), .ZN(n205) );
  DFF_X1 \state_reg[4]  ( .D(n21), .CK(clk), .Q(state[4]), .QN(n76) );
  DFF_X1 \state_reg[2]  ( .D(N34), .CK(clk), .Q(state[2]), .QN(n79) );
  DFF_X1 \addr_y_reg[0]  ( .D(N141), .CK(clk), .Q(addr_y[0]), .QN(n113) );
  DFF_X1 \addr_y_reg[1]  ( .D(N142), .CK(clk), .Q(addr_y[1]), .QN(n112) );
  DFF_X1 \state_reg[1]  ( .D(N33), .CK(clk), .Q(state[1]), .QN(n80) );
  DFF_X1 \addr_y_reg[2]  ( .D(N143), .CK(clk), .Q(addr_y[2]), .QN(n111) );
  DFF_X1 \state_reg[0]  ( .D(N32), .CK(clk), .Q(state[0]), .QN(n81) );
  DFF_X1 \addr_x_reg[2]  ( .D(N133), .CK(clk), .Q(addr_x[2]), .QN(n108) );
  DFF_X1 \addr_a8_reg[0]  ( .D(n8), .CK(clk), .Q(addr_a8[0]), .QN(n107) );
  DFF_X1 \addr_a7_reg[0]  ( .D(n6), .CK(clk), .Q(addr_a7[0]), .QN(n104) );
  DFF_X1 \addr_a6_reg[0]  ( .D(n5), .CK(clk), .Q(addr_a6[0]), .QN(n101) );
  DFF_X1 \addr_a5_reg[0]  ( .D(n19), .CK(clk), .Q(addr_a5[0]), .QN(n98) );
  DFF_X1 \addr_a4_reg[0]  ( .D(n17), .CK(clk), .Q(addr_a4[0]), .QN(n95) );
  DFF_X1 \addr_a3_reg[0]  ( .D(n15), .CK(clk), .Q(addr_a3[0]), .QN(n92) );
  DFF_X1 \addr_a2_reg[0]  ( .D(n13), .CK(clk), .Q(addr_a2[0]), .QN(n88) );
  DFF_X1 \addr_a1_reg[0]  ( .D(n11), .CK(clk), .Q(addr_a1[0]), .QN(n85) );
  DFF_X1 \addr_a8_reg[1]  ( .D(N122), .CK(clk), .Q(addr_a8[1]), .QN(n106) );
  DFF_X1 \addr_a7_reg[1]  ( .D(N111), .CK(clk), .Q(addr_a7[1]), .QN(n103) );
  DFF_X1 \addr_a6_reg[1]  ( .D(N100), .CK(clk), .Q(addr_a6[1]), .QN(n100) );
  DFF_X1 \addr_a5_reg[1]  ( .D(N89), .CK(clk), .Q(addr_a5[1]), .QN(n97) );
  DFF_X1 \addr_a4_reg[1]  ( .D(N78), .CK(clk), .Q(addr_a4[1]), .QN(n94) );
  DFF_X1 \addr_a3_reg[1]  ( .D(N67), .CK(clk), .Q(addr_a3[1]), .QN(n91) );
  DFF_X1 \addr_a2_reg[1]  ( .D(N56), .CK(clk), .Q(addr_a2[1]), .QN(n87) );
  DFF_X1 \addr_a1_reg[1]  ( .D(N45), .CK(clk), .Q(addr_a1[1]), .QN(n84) );
  DFF_X1 \addr_a8_reg[2]  ( .D(N123), .CK(clk), .Q(addr_a8[2]), .QN(n105) );
  DFF_X1 \addr_a7_reg[2]  ( .D(N112), .CK(clk), .Q(addr_a7[2]), .QN(n102) );
  DFF_X1 \addr_a6_reg[2]  ( .D(N101), .CK(clk), .Q(addr_a6[2]), .QN(n99) );
  DFF_X1 \addr_a5_reg[2]  ( .D(N90), .CK(clk), .Q(addr_a5[2]), .QN(n96) );
  DFF_X1 \addr_a4_reg[2]  ( .D(N79), .CK(clk), .Q(addr_a4[2]), .QN(n93) );
  DFF_X1 \addr_a3_reg[2]  ( .D(N68), .CK(clk), .Q(addr_a3[2]), .QN(n90) );
  DFF_X1 \addr_a2_reg[2]  ( .D(N57), .CK(clk), .Q(addr_a2[2]), .QN(n86) );
  DFF_X1 \addr_a1_reg[2]  ( .D(N46), .CK(clk), .Q(addr_a1[2]), .QN(n83) );
  INV_X1 U3 ( .A(n248), .ZN(n22) );
  INV_X1 U4 ( .A(n224), .ZN(n10) );
  INV_X1 U5 ( .A(n246), .ZN(n28) );
  NAND2_X1 U6 ( .A1(n233), .A2(n133), .ZN(n248) );
  NAND2_X1 U7 ( .A1(n131), .A2(n245), .ZN(n123) );
  NAND2_X1 U8 ( .A1(n131), .A2(n149), .ZN(n145) );
  INV_X1 U9 ( .A(n150), .ZN(n27) );
  NAND2_X1 U10 ( .A1(n131), .A2(n157), .ZN(n153) );
  NAND2_X1 U11 ( .A1(n131), .A2(n141), .ZN(n137) );
  NAND2_X1 U12 ( .A1(n131), .A2(n132), .ZN(n127) );
  NAND2_X1 U13 ( .A1(n131), .A2(n166), .ZN(n162) );
  NOR2_X1 U14 ( .A1(n32), .A2(n23), .ZN(n133) );
  OAI21_X1 U15 ( .B1(n37), .B2(n117), .A(n131), .ZN(n224) );
  NAND2_X1 U16 ( .A1(n202), .A2(n116), .ZN(N148) );
  AND2_X1 U17 ( .A1(n207), .A2(n180), .ZN(n191) );
  NAND2_X1 U18 ( .A1(n117), .A2(n180), .ZN(N146) );
  INV_X1 U19 ( .A(n210), .ZN(n29) );
  AND2_X1 U20 ( .A1(n121), .A2(n167), .ZN(n233) );
  AND4_X1 U21 ( .A1(n247), .A2(n178), .A3(n210), .A4(n26), .ZN(n158) );
  INV_X1 U22 ( .A(N148), .ZN(n26) );
  OR2_X1 U23 ( .A1(n189), .A2(N37), .ZN(n188) );
  OAI211_X2 U24 ( .C1(n205), .C2(n210), .A(n116), .B(n178), .ZN(n124) );
  OAI221_X1 U25 ( .B1(n169), .B2(n167), .C1(n121), .C2(n35), .A(n28), .ZN(n177) );
  INV_X1 U26 ( .A(n184), .ZN(n35) );
  AOI21_X1 U27 ( .B1(n251), .B2(n33), .A(n189), .ZN(n178) );
  OAI22_X1 U28 ( .A1(n117), .A2(n205), .B1(n173), .B2(n170), .ZN(n176) );
  NAND4_X1 U29 ( .A1(n202), .A2(n159), .A3(n247), .A4(n249), .ZN(n131) );
  NOR3_X1 U30 ( .A1(n124), .A2(n248), .A3(n246), .ZN(n249) );
  OAI22_X1 U31 ( .A1(n37), .A2(n117), .B1(n172), .B2(n195), .ZN(n192) );
  OAI22_X1 U32 ( .A1(n190), .A2(n116), .B1(n184), .B2(n121), .ZN(n204) );
  NAND2_X1 U33 ( .A1(n222), .A2(n252), .ZN(n116) );
  NAND2_X1 U34 ( .A1(n254), .A2(n251), .ZN(n117) );
  OAI21_X1 U35 ( .B1(n119), .B2(n36), .A(n118), .ZN(n150) );
  INV_X1 U36 ( .A(n194), .ZN(n36) );
  OAI21_X1 U37 ( .B1(n190), .B2(n208), .A(n209), .ZN(n183) );
  NAND2_X1 U38 ( .A1(n254), .A2(n252), .ZN(n121) );
  NAND2_X1 U39 ( .A1(n131), .A2(n232), .ZN(n228) );
  NAND2_X1 U40 ( .A1(n131), .A2(n240), .ZN(n236) );
  NAND2_X1 U41 ( .A1(n250), .A2(n252), .ZN(n119) );
  NAND2_X1 U42 ( .A1(n255), .A2(n254), .ZN(n210) );
  NAND2_X1 U43 ( .A1(n255), .A2(n250), .ZN(n167) );
  NAND2_X1 U44 ( .A1(n250), .A2(n251), .ZN(n118) );
  INV_X1 U45 ( .A(n205), .ZN(n37) );
  NAND2_X1 U46 ( .A1(n251), .A2(n222), .ZN(n209) );
  NAND2_X1 U47 ( .A1(n221), .A2(n250), .ZN(n120) );
  INV_X1 U48 ( .A(n216), .ZN(n30) );
  NAND2_X1 U49 ( .A1(n33), .A2(n221), .ZN(n202) );
  INV_X1 U50 ( .A(n212), .ZN(n33) );
  NAND2_X1 U51 ( .A1(n33), .A2(n252), .ZN(n180) );
  NAND2_X1 U52 ( .A1(n255), .A2(n222), .ZN(n208) );
  NOR2_X1 U53 ( .A1(n2), .A2(n116), .ZN(N37) );
  INV_X1 U54 ( .A(n190), .ZN(n2) );
  INV_X1 U55 ( .A(n172), .ZN(n32) );
  NAND2_X1 U56 ( .A1(n221), .A2(n254), .ZN(n207) );
  AND3_X1 U57 ( .A1(n158), .A2(n159), .A3(n28), .ZN(n134) );
  INV_X1 U58 ( .A(n222), .ZN(n34) );
  AND3_X1 U59 ( .A1(n158), .A2(n159), .A3(n22), .ZN(n142) );
  INV_X1 U60 ( .A(n193), .ZN(n3) );
  AND2_X1 U61 ( .A1(n221), .A2(n222), .ZN(n189) );
  INV_X1 U62 ( .A(n173), .ZN(n23) );
  INV_X1 U63 ( .A(n168), .ZN(n21) );
  AOI221_X1 U64 ( .B1(n169), .B2(wr_en_a5), .C1(n170), .C2(wr_en_a8), .A(n171), 
        .ZN(n168) );
  OR2_X1 U65 ( .A1(wr_en_a7), .A2(wr_en_a6), .ZN(n171) );
  AND4_X1 U66 ( .A1(n207), .A2(n25), .A3(n209), .A4(n256), .ZN(n247) );
  AND2_X1 U67 ( .A1(n208), .A2(n31), .ZN(n256) );
  INV_X1 U68 ( .A(N146), .ZN(n25) );
  AOI211_X1 U69 ( .C1(n80), .C2(n81), .A(state[4]), .B(n34), .ZN(n216) );
  NOR3_X1 U70 ( .A1(state[0]), .A2(state[4]), .A3(n80), .ZN(n251) );
  NOR2_X1 U71 ( .A1(state[3]), .A2(state[2]), .ZN(n254) );
  NOR3_X1 U72 ( .A1(n97), .A2(n98), .A3(n96), .ZN(n169) );
  NOR3_X1 U73 ( .A1(n112), .A2(n113), .A3(n111), .ZN(n190) );
  NOR3_X1 U74 ( .A1(n81), .A2(state[4]), .A3(n80), .ZN(n255) );
  AOI211_X1 U75 ( .C1(n205), .C2(n29), .A(n183), .B(n206), .ZN(n193) );
  OAI22_X1 U76 ( .A1(n39), .A2(n191), .B1(n167), .B2(n169), .ZN(n206) );
  INV_X1 U77 ( .A(start), .ZN(n39) );
  NOR2_X1 U78 ( .A1(n79), .A2(state[3]), .ZN(n222) );
  NOR2_X1 U79 ( .A1(n211), .A2(state[0]), .ZN(n221) );
  NOR4_X1 U80 ( .A1(n159), .A2(n101), .A3(n100), .A4(n99), .ZN(n200) );
  NOR4_X1 U81 ( .A1(n120), .A2(n88), .A3(n87), .A4(n86), .ZN(n199) );
  NOR2_X1 U82 ( .A1(n81), .A2(n211), .ZN(n252) );
  NOR3_X1 U83 ( .A1(n84), .A2(n85), .A3(n83), .ZN(n184) );
  NOR3_X1 U84 ( .A1(n91), .A2(n92), .A3(n90), .ZN(n194) );
  OAI221_X1 U85 ( .B1(n191), .B2(n38), .C1(n194), .C2(n119), .A(n202), .ZN(
        n198) );
  INV_X1 U86 ( .A(loadMatrix), .ZN(n38) );
  NAND4_X1 U87 ( .A1(state[4]), .A2(n254), .A3(state[0]), .A4(n80), .ZN(n172)
         );
  AOI22_X1 U88 ( .A1(n113), .A2(n216), .B1(n30), .B2(n219), .ZN(n217) );
  AOI21_X1 U89 ( .B1(n101), .B2(n123), .A(n124), .ZN(n243) );
  AOI21_X1 U90 ( .B1(n92), .B2(n145), .A(n124), .ZN(n146) );
  AOI21_X1 U91 ( .B1(n88), .B2(n153), .A(n124), .ZN(n154) );
  AOI21_X1 U92 ( .B1(n95), .B2(n137), .A(n124), .ZN(n138) );
  AOI21_X1 U93 ( .B1(n98), .B2(n127), .A(n124), .ZN(n128) );
  AOI21_X1 U94 ( .B1(n85), .B2(n162), .A(n124), .ZN(n163) );
  AOI21_X1 U95 ( .B1(n107), .B2(n228), .A(n124), .ZN(n229) );
  AOI21_X1 U96 ( .B1(n104), .B2(n236), .A(n124), .ZN(n237) );
  NOR2_X1 U97 ( .A1(n173), .A2(reset), .ZN(wr_en_a8) );
  NOR2_X1 U98 ( .A1(n167), .A2(reset), .ZN(wr_en_a5) );
  NOR2_X1 U99 ( .A1(n172), .A2(reset), .ZN(wr_en_a7) );
  NAND2_X1 U100 ( .A1(n253), .A2(n80), .ZN(n159) );
  NOR2_X1 U101 ( .A1(n159), .A2(reset), .ZN(wr_en_a6) );
  NOR2_X1 U102 ( .A1(reset), .A2(n117), .ZN(wr_en_x) );
  NOR2_X1 U103 ( .A1(reset), .A2(n116), .ZN(wr_en_y) );
  NOR2_X1 U104 ( .A1(reset), .A2(n121), .ZN(wr_en_a1) );
  OAI211_X1 U105 ( .C1(loadVector), .C2(n180), .A(n24), .B(n193), .ZN(n203) );
  INV_X1 U106 ( .A(n176), .ZN(n24) );
  NOR2_X1 U107 ( .A1(reset), .A2(n118), .ZN(wr_en_a4) );
  NOR2_X1 U108 ( .A1(reset), .A2(n120), .ZN(wr_en_a2) );
  NOR2_X1 U109 ( .A1(reset), .A2(n119), .ZN(wr_en_a3) );
  AND2_X1 U110 ( .A1(state[3]), .A2(state[2]), .ZN(n250) );
  NAND2_X1 U111 ( .A1(n76), .A2(n80), .ZN(n211) );
  NAND2_X1 U112 ( .A1(n253), .A2(state[1]), .ZN(n173) );
  AOI21_X1 U113 ( .B1(n181), .B2(n182), .A(reset), .ZN(N34) );
  AOI21_X1 U114 ( .B1(n29), .B2(n37), .A(N148), .ZN(n182) );
  NOR2_X1 U115 ( .A1(n177), .A2(n183), .ZN(n181) );
  AOI21_X1 U116 ( .B1(n185), .B2(n186), .A(reset), .ZN(N33) );
  AOI221_X1 U117 ( .B1(n187), .B2(loadVector), .C1(n23), .C2(n170), .A(n188), 
        .ZN(n186) );
  NOR3_X1 U118 ( .A1(n192), .A2(n150), .A3(n3), .ZN(n185) );
  NOR2_X1 U119 ( .A1(loadMatrix), .A2(n191), .ZN(n187) );
  AOI21_X1 U120 ( .B1(n196), .B2(n197), .A(reset), .ZN(N32) );
  NOR4_X1 U121 ( .A1(n198), .A2(n199), .A3(n200), .A4(n201), .ZN(n197) );
  AOI211_X1 U122 ( .C1(n32), .C2(n195), .A(n203), .B(n204), .ZN(n196) );
  NOR4_X1 U123 ( .A1(n118), .A2(n95), .A3(n94), .A4(n93), .ZN(n201) );
  NAND2_X1 U124 ( .A1(n221), .A2(n79), .ZN(n219) );
  OAI21_X1 U125 ( .B1(n243), .B2(n100), .A(n244), .ZN(N100) );
  OAI21_X1 U126 ( .B1(n237), .B2(n103), .A(n238), .ZN(N111) );
  OAI21_X1 U127 ( .B1(n229), .B2(n106), .A(n230), .ZN(N122) );
  OAI21_X1 U128 ( .B1(n146), .B2(n91), .A(n147), .ZN(N67) );
  OAI21_X1 U129 ( .B1(n154), .B2(n87), .A(n155), .ZN(N56) );
  OAI21_X1 U130 ( .B1(n138), .B2(n94), .A(n139), .ZN(N78) );
  OAI21_X1 U131 ( .B1(n163), .B2(n84), .A(n164), .ZN(N45) );
  OAI21_X1 U132 ( .B1(n128), .B2(n97), .A(n129), .ZN(N89) );
  OAI21_X1 U133 ( .B1(n217), .B2(n112), .A(n218), .ZN(N142) );
  OAI21_X1 U134 ( .B1(n214), .B2(n111), .A(n215), .ZN(N143) );
  NAND4_X1 U135 ( .A1(n216), .A2(addr_y[1]), .A3(addr_y[0]), .A4(n111), .ZN(
        n215) );
  AOI21_X1 U136 ( .B1(n216), .B2(n112), .A(n1), .ZN(n214) );
  INV_X1 U137 ( .A(n217), .ZN(n1) );
  AND3_X1 U138 ( .A1(n254), .A2(n81), .A3(state[4]), .ZN(n253) );
  NAND2_X1 U139 ( .A1(state[3]), .A2(n79), .ZN(n212) );
  OAI21_X1 U140 ( .B1(n241), .B2(n99), .A(n242), .ZN(N101) );
  NAND4_X1 U141 ( .A1(addr_a6[1]), .A2(addr_a6[0]), .A3(n123), .A4(n99), .ZN(
        n242) );
  AOI21_X1 U142 ( .B1(n123), .B2(n100), .A(n4), .ZN(n241) );
  INV_X1 U143 ( .A(n243), .ZN(n4) );
  OAI21_X1 U144 ( .B1(n151), .B2(n86), .A(n152), .ZN(N57) );
  NAND4_X1 U145 ( .A1(addr_a2[1]), .A2(addr_a2[0]), .A3(n153), .A4(n86), .ZN(
        n152) );
  AOI21_X1 U146 ( .B1(n153), .B2(n87), .A(n14), .ZN(n151) );
  INV_X1 U147 ( .A(n154), .ZN(n14) );
  OAI21_X1 U148 ( .B1(n135), .B2(n93), .A(n136), .ZN(N79) );
  NAND4_X1 U149 ( .A1(addr_a4[1]), .A2(addr_a4[0]), .A3(n137), .A4(n93), .ZN(
        n136) );
  AOI21_X1 U150 ( .B1(n137), .B2(n94), .A(n18), .ZN(n135) );
  INV_X1 U151 ( .A(n138), .ZN(n18) );
  OAI21_X1 U152 ( .B1(n143), .B2(n90), .A(n144), .ZN(N68) );
  NAND4_X1 U153 ( .A1(addr_a3[1]), .A2(addr_a3[0]), .A3(n145), .A4(n90), .ZN(
        n144) );
  AOI21_X1 U154 ( .B1(n145), .B2(n91), .A(n16), .ZN(n143) );
  INV_X1 U155 ( .A(n146), .ZN(n16) );
  OAI21_X1 U156 ( .B1(n125), .B2(n96), .A(n126), .ZN(N90) );
  NAND4_X1 U157 ( .A1(addr_a5[1]), .A2(addr_a5[0]), .A3(n127), .A4(n96), .ZN(
        n126) );
  AOI21_X1 U158 ( .B1(n127), .B2(n97), .A(n20), .ZN(n125) );
  INV_X1 U159 ( .A(n128), .ZN(n20) );
  OAI21_X1 U160 ( .B1(n160), .B2(n83), .A(n161), .ZN(N46) );
  NAND4_X1 U161 ( .A1(addr_a1[1]), .A2(addr_a1[0]), .A3(n162), .A4(n83), .ZN(
        n161) );
  AOI21_X1 U162 ( .B1(n162), .B2(n84), .A(n12), .ZN(n160) );
  INV_X1 U163 ( .A(n163), .ZN(n12) );
  OAI21_X1 U164 ( .B1(addr_y[0]), .B2(n30), .A(n220), .ZN(N141) );
  OAI21_X1 U165 ( .B1(n226), .B2(n105), .A(n227), .ZN(N123) );
  NAND4_X1 U166 ( .A1(addr_a8[1]), .A2(addr_a8[0]), .A3(n228), .A4(n105), .ZN(
        n227) );
  AOI21_X1 U167 ( .B1(n228), .B2(n106), .A(n9), .ZN(n226) );
  INV_X1 U168 ( .A(n229), .ZN(n9) );
  OAI21_X1 U169 ( .B1(n234), .B2(n102), .A(n235), .ZN(N112) );
  NAND4_X1 U170 ( .A1(addr_a7[1]), .A2(addr_a7[0]), .A3(n236), .A4(n102), .ZN(
        n235) );
  AOI21_X1 U171 ( .B1(n236), .B2(n103), .A(n7), .ZN(n234) );
  INV_X1 U172 ( .A(n237), .ZN(n7) );
  OAI21_X1 U173 ( .B1(n10), .B2(n108), .A(n223), .ZN(N133) );
  NOR2_X1 U174 ( .A1(addr_x[0]), .A2(n10), .ZN(N131) );
  NOR2_X1 U175 ( .A1(n10), .A2(n225), .ZN(N132) );
  XNOR2_X1 U176 ( .A(addr_x[1]), .B(addr_x[0]), .ZN(n225) );
  NOR2_X1 U177 ( .A1(reset), .A2(n174), .ZN(N35) );
  NOR3_X1 U178 ( .A1(n175), .A2(n176), .A3(n177), .ZN(n174) );
  OR4_X1 U179 ( .A1(n180), .A2(loadMatrix), .A3(loadVector), .A4(start), .ZN(
        n179) );
  INV_X1 U180 ( .A(n257), .ZN(n31) );
  OAI21_X1 U181 ( .B1(n254), .B2(n76), .A(n258), .ZN(n257) );
  OAI211_X1 U182 ( .C1(n33), .C2(state[4]), .A(state[0]), .B(state[1]), .ZN(
        n258) );
  INV_X1 U183 ( .A(n122), .ZN(n5) );
  AOI22_X1 U184 ( .A1(n101), .A2(n123), .B1(n124), .B2(addr_a6[0]), .ZN(n122)
         );
  INV_X1 U185 ( .A(n148), .ZN(n15) );
  AOI22_X1 U186 ( .A1(n92), .A2(n145), .B1(n124), .B2(addr_a3[0]), .ZN(n148)
         );
  INV_X1 U187 ( .A(n156), .ZN(n13) );
  AOI22_X1 U188 ( .A1(n88), .A2(n153), .B1(n124), .B2(addr_a2[0]), .ZN(n156)
         );
  INV_X1 U189 ( .A(n140), .ZN(n17) );
  AOI22_X1 U190 ( .A1(n95), .A2(n137), .B1(n124), .B2(addr_a4[0]), .ZN(n140)
         );
  INV_X1 U191 ( .A(n130), .ZN(n19) );
  AOI22_X1 U192 ( .A1(n98), .A2(n127), .B1(n124), .B2(addr_a5[0]), .ZN(n130)
         );
  INV_X1 U193 ( .A(n165), .ZN(n11) );
  AOI22_X1 U194 ( .A1(n85), .A2(n162), .B1(n124), .B2(addr_a1[0]), .ZN(n165)
         );
  INV_X1 U195 ( .A(n231), .ZN(n8) );
  AOI22_X1 U196 ( .A1(n107), .A2(n228), .B1(n124), .B2(addr_a8[0]), .ZN(n231)
         );
  INV_X1 U197 ( .A(n239), .ZN(n6) );
  AOI22_X1 U198 ( .A1(n104), .A2(n236), .B1(n124), .B2(addr_a7[0]), .ZN(n239)
         );
  OAI22_X1 U199 ( .A1(n211), .A2(n34), .B1(n212), .B2(n213), .ZN(N147) );
  NAND2_X1 U200 ( .A1(n81), .A2(n76), .ZN(n213) );
endmodule


module mvm_8_8_12_1 ( clk, reset, loadMatrix, loadVector, start, done, data_in, 
        data_out );
  input [11:0] data_in;
  output [23:0] data_out;
  input clk, reset, loadMatrix, loadVector, start;
  output done;
  wire   wr_en_x, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6,
         wr_en_a7, wr_en_a8, wr_en_y, clear_acc, clc, clc1;
  wire   [2:0] addr_x;
  wire   [2:0] addr_a1;
  wire   [2:0] addr_a2;
  wire   [2:0] addr_a3;
  wire   [2:0] addr_a4;
  wire   [2:0] addr_a5;
  wire   [2:0] addr_a6;
  wire   [2:0] addr_a7;
  wire   [2:0] addr_a8;
  wire   [2:0] addr_y;

  datapath d ( .clk(clk), .data_in(data_in), .addr_x(addr_x), .wr_en_x(wr_en_x), .addr_a1(addr_a1), .addr_a2(addr_a2), .addr_a3(addr_a3), .addr_a4(addr_a4), 
        .addr_a5(addr_a5), .addr_a6(addr_a6), .addr_a7(addr_a7), .addr_a8(
        addr_a8), .wr_en_a1(wr_en_a1), .wr_en_a2(wr_en_a2), .wr_en_a3(wr_en_a3), .wr_en_a4(wr_en_a4), .wr_en_a5(wr_en_a5), .wr_en_a6(wr_en_a6), .wr_en_a7(
        wr_en_a7), .wr_en_a8(wr_en_a8), .addr_y(addr_y), .wr_en_y(wr_en_y), 
        .clear_acc(clear_acc), .clc(clc), .clc1(clc1), .data_out(data_out) );
  ctrlpath c ( .clk(clk), .reset(reset), .start(start), .addr_x(addr_x), 
        .wr_en_x(wr_en_x), .addr_a1(addr_a1), .addr_a2(addr_a2), .addr_a3(
        addr_a3), .addr_a4(addr_a4), .addr_a5(addr_a5), .addr_a6(addr_a6), 
        .addr_a7(addr_a7), .addr_a8(addr_a8), .wr_en_a1(wr_en_a1), .wr_en_a2(
        wr_en_a2), .wr_en_a3(wr_en_a3), .wr_en_a4(wr_en_a4), .wr_en_a5(
        wr_en_a5), .wr_en_a6(wr_en_a6), .wr_en_a7(wr_en_a7), .wr_en_a8(
        wr_en_a8), .clear_acc(clear_acc), .clc(clc), .clc1(clc1), .addr_y(
        addr_y), .wr_en_y(wr_en_y), .done(done), .loadMatrix(loadMatrix), 
        .loadVector(loadVector) );
endmodule

