
module memory_WIDTH16_SIZE8_LOGSIZE3_0 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] ,
         \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][15] , \mem[6][14] , \mem[6][13] ,
         \mem[6][12] , \mem[6][11] , \mem[6][10] , \mem[6][9] , \mem[6][8] ,
         \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] ,
         \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[5][15] , \mem[5][14] ,
         \mem[5][13] , \mem[5][12] , \mem[5][11] , \mem[5][10] , \mem[5][9] ,
         \mem[5][8] , \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] ,
         \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][15] ,
         \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] , \mem[4][10] ,
         \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \mem_reg[7][15]  ( .D(n285), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n284), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n283), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n282), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n281), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n280), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n279), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n278), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n277), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n276), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n275), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n274), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n273), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n272), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n271), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n270), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n269), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n268), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n267), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n266), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n265), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n264), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n263), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n262), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n261), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n260), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n259), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n258), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n257), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n256), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n255), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n254), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n253), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n252), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n251), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n250), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n249), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n248), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n247), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n246), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n245), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n244), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n243), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n242), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n241), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n240), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n239), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n238), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n237), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n236), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n235), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n234), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n233), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n232), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n231), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n230), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n229), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n228), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n227), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n226), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n225), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n224), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n223), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n222), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n221), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n220), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n219), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n218), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n217), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n216), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n215), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n214), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n213), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n212), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n211), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n210), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n209), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n208), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n207), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n206), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n205), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n204), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n203), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n202), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n201), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n200), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n199), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n198), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n197), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n196), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n195), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n194), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n193), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n192), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n191), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n190), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n189), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n188), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n187), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n186), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n185), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n184), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n183), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n182), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n181), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n180), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n179), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n178), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n177), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n176), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n175), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n174), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n173), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n172), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n171), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n170), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n169), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n168), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n167), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n166), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n165), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n164), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n163), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n162), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n161), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n160), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n159), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n158), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U280 ( .A1(n376), .A2(n377), .A3(n37), .ZN(n20) );
  NAND3_X1 U281 ( .A1(n37), .A2(n377), .A3(N10), .ZN(n38) );
  NAND3_X1 U282 ( .A1(n37), .A2(n376), .A3(N11), .ZN(n55) );
  NAND3_X1 U283 ( .A1(N10), .A2(n37), .A3(N11), .ZN(n72) );
  NAND3_X1 U284 ( .A1(n376), .A2(n377), .A3(n106), .ZN(n89) );
  NAND3_X1 U285 ( .A1(N10), .A2(n377), .A3(n106), .ZN(n107) );
  NAND3_X1 U286 ( .A1(N11), .A2(n376), .A3(n106), .ZN(n124) );
  NAND3_X1 U287 ( .A1(N11), .A2(N10), .A3(n106), .ZN(n141) );
  SDFF_X1 \data_out_reg[2]  ( .D(n19), .SI(n16), .SE(N12), .CK(clk), .Q(
        data_out[2]) );
  SDFF_X1 \data_out_reg[4]  ( .D(n297), .SI(n294), .SE(N12), .CK(clk), .Q(
        data_out[4]) );
  SDFF_X1 \data_out_reg[14]  ( .D(n357), .SI(n354), .SE(N12), .CK(clk), .Q(
        data_out[14]) );
  SDFF_X1 \data_out_reg[12]  ( .D(n345), .SI(n342), .SE(N12), .CK(clk), .Q(
        data_out[12]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n327), .SI(n324), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[10]  ( .D(n333), .SI(n330), .SE(N12), .CK(clk), .Q(
        data_out[10]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n315), .SI(n312), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n339), .SI(n336), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[0]  ( .D(n7), .SI(n4), .SE(N12), .CK(clk), .Q(
        data_out[0]) );
  SDFF_X1 \data_out_reg[6]  ( .D(n309), .SI(n306), .SE(N12), .CK(clk), .Q(
        data_out[6]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n291), .SI(n288), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n351), .SI(n348), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n303), .SI(n300), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n363), .SI(n360), .SE(N12), .CK(clk), .Q(
        data_out[15]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n13), .SI(n10), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[8]  ( .D(n321), .SI(n318), .SE(N12), .CK(clk), .Q(
        data_out[8]) );
  BUF_X1 U3 ( .A(N10), .Z(n366) );
  BUF_X1 U4 ( .A(N10), .Z(n367) );
  BUF_X1 U5 ( .A(n20), .Z(n375) );
  BUF_X1 U6 ( .A(n38), .Z(n374) );
  BUF_X1 U7 ( .A(n72), .Z(n372) );
  BUF_X1 U8 ( .A(n89), .Z(n371) );
  BUF_X1 U9 ( .A(n107), .Z(n370) );
  BUF_X1 U10 ( .A(n124), .Z(n369) );
  BUF_X1 U11 ( .A(n141), .Z(n368) );
  BUF_X1 U12 ( .A(n55), .Z(n373) );
  BUF_X1 U13 ( .A(N10), .Z(n365) );
  BUF_X1 U14 ( .A(N11), .Z(n364) );
  NOR2_X1 U15 ( .A1(n378), .A2(N12), .ZN(n37) );
  INV_X1 U16 ( .A(wr_en), .ZN(n378) );
  AND2_X1 U17 ( .A1(N12), .A2(wr_en), .ZN(n106) );
  INV_X1 U18 ( .A(N10), .ZN(n376) );
  OAI21_X1 U19 ( .B1(n387), .B2(n72), .A(n80), .ZN(n213) );
  NAND2_X1 U20 ( .A1(\mem[3][7] ), .A2(n372), .ZN(n80) );
  OAI21_X1 U21 ( .B1(n386), .B2(n372), .A(n81), .ZN(n214) );
  NAND2_X1 U22 ( .A1(\mem[3][8] ), .A2(n372), .ZN(n81) );
  OAI21_X1 U23 ( .B1(n385), .B2(n72), .A(n82), .ZN(n215) );
  NAND2_X1 U24 ( .A1(\mem[3][9] ), .A2(n372), .ZN(n82) );
  OAI21_X1 U25 ( .B1(n384), .B2(n72), .A(n83), .ZN(n216) );
  NAND2_X1 U26 ( .A1(\mem[3][10] ), .A2(n372), .ZN(n83) );
  OAI21_X1 U27 ( .B1(n383), .B2(n72), .A(n84), .ZN(n217) );
  NAND2_X1 U28 ( .A1(\mem[3][11] ), .A2(n372), .ZN(n84) );
  OAI21_X1 U29 ( .B1(n382), .B2(n72), .A(n85), .ZN(n218) );
  NAND2_X1 U30 ( .A1(\mem[3][12] ), .A2(n372), .ZN(n85) );
  OAI21_X1 U31 ( .B1(n381), .B2(n72), .A(n86), .ZN(n219) );
  NAND2_X1 U32 ( .A1(\mem[3][13] ), .A2(n372), .ZN(n86) );
  OAI21_X1 U33 ( .B1(n380), .B2(n72), .A(n87), .ZN(n220) );
  NAND2_X1 U34 ( .A1(\mem[3][14] ), .A2(n372), .ZN(n87) );
  OAI21_X1 U35 ( .B1(n387), .B2(n107), .A(n115), .ZN(n245) );
  NAND2_X1 U36 ( .A1(\mem[5][7] ), .A2(n370), .ZN(n115) );
  OAI21_X1 U37 ( .B1(n386), .B2(n370), .A(n116), .ZN(n246) );
  NAND2_X1 U38 ( .A1(\mem[5][8] ), .A2(n370), .ZN(n116) );
  OAI21_X1 U39 ( .B1(n385), .B2(n107), .A(n117), .ZN(n247) );
  NAND2_X1 U40 ( .A1(\mem[5][9] ), .A2(n370), .ZN(n117) );
  OAI21_X1 U41 ( .B1(n384), .B2(n107), .A(n118), .ZN(n248) );
  NAND2_X1 U42 ( .A1(\mem[5][10] ), .A2(n370), .ZN(n118) );
  OAI21_X1 U43 ( .B1(n383), .B2(n107), .A(n119), .ZN(n249) );
  NAND2_X1 U44 ( .A1(\mem[5][11] ), .A2(n370), .ZN(n119) );
  OAI21_X1 U45 ( .B1(n382), .B2(n107), .A(n120), .ZN(n250) );
  NAND2_X1 U46 ( .A1(\mem[5][12] ), .A2(n370), .ZN(n120) );
  OAI21_X1 U47 ( .B1(n381), .B2(n107), .A(n121), .ZN(n251) );
  NAND2_X1 U48 ( .A1(\mem[5][13] ), .A2(n370), .ZN(n121) );
  OAI21_X1 U49 ( .B1(n380), .B2(n107), .A(n122), .ZN(n252) );
  NAND2_X1 U50 ( .A1(\mem[5][14] ), .A2(n370), .ZN(n122) );
  OAI21_X1 U51 ( .B1(n387), .B2(n141), .A(n149), .ZN(n277) );
  NAND2_X1 U52 ( .A1(\mem[7][7] ), .A2(n368), .ZN(n149) );
  OAI21_X1 U53 ( .B1(n386), .B2(n368), .A(n150), .ZN(n278) );
  NAND2_X1 U54 ( .A1(\mem[7][8] ), .A2(n368), .ZN(n150) );
  OAI21_X1 U55 ( .B1(n385), .B2(n141), .A(n151), .ZN(n279) );
  NAND2_X1 U56 ( .A1(\mem[7][9] ), .A2(n368), .ZN(n151) );
  OAI21_X1 U57 ( .B1(n384), .B2(n141), .A(n152), .ZN(n280) );
  NAND2_X1 U58 ( .A1(\mem[7][10] ), .A2(n368), .ZN(n152) );
  OAI21_X1 U59 ( .B1(n383), .B2(n141), .A(n153), .ZN(n281) );
  NAND2_X1 U60 ( .A1(\mem[7][11] ), .A2(n368), .ZN(n153) );
  OAI21_X1 U61 ( .B1(n382), .B2(n141), .A(n154), .ZN(n282) );
  NAND2_X1 U62 ( .A1(\mem[7][12] ), .A2(n368), .ZN(n154) );
  OAI21_X1 U63 ( .B1(n381), .B2(n141), .A(n155), .ZN(n283) );
  NAND2_X1 U64 ( .A1(\mem[7][13] ), .A2(n368), .ZN(n155) );
  OAI21_X1 U65 ( .B1(n380), .B2(n141), .A(n156), .ZN(n284) );
  NAND2_X1 U66 ( .A1(\mem[7][14] ), .A2(n368), .ZN(n156) );
  OAI21_X1 U67 ( .B1(n387), .B2(n124), .A(n132), .ZN(n261) );
  NAND2_X1 U68 ( .A1(\mem[6][7] ), .A2(n369), .ZN(n132) );
  OAI21_X1 U69 ( .B1(n386), .B2(n369), .A(n133), .ZN(n262) );
  NAND2_X1 U70 ( .A1(\mem[6][8] ), .A2(n369), .ZN(n133) );
  OAI21_X1 U71 ( .B1(n385), .B2(n124), .A(n134), .ZN(n263) );
  NAND2_X1 U72 ( .A1(\mem[6][9] ), .A2(n369), .ZN(n134) );
  OAI21_X1 U73 ( .B1(n384), .B2(n124), .A(n135), .ZN(n264) );
  NAND2_X1 U74 ( .A1(\mem[6][10] ), .A2(n369), .ZN(n135) );
  OAI21_X1 U75 ( .B1(n383), .B2(n124), .A(n136), .ZN(n265) );
  NAND2_X1 U76 ( .A1(\mem[6][11] ), .A2(n369), .ZN(n136) );
  OAI21_X1 U77 ( .B1(n382), .B2(n124), .A(n137), .ZN(n266) );
  NAND2_X1 U78 ( .A1(\mem[6][12] ), .A2(n369), .ZN(n137) );
  OAI21_X1 U79 ( .B1(n381), .B2(n124), .A(n138), .ZN(n267) );
  NAND2_X1 U80 ( .A1(\mem[6][13] ), .A2(n369), .ZN(n138) );
  OAI21_X1 U81 ( .B1(n380), .B2(n124), .A(n139), .ZN(n268) );
  NAND2_X1 U82 ( .A1(\mem[6][14] ), .A2(n369), .ZN(n139) );
  OAI21_X1 U83 ( .B1(n387), .B2(n38), .A(n46), .ZN(n181) );
  NAND2_X1 U84 ( .A1(\mem[1][7] ), .A2(n374), .ZN(n46) );
  OAI21_X1 U85 ( .B1(n386), .B2(n374), .A(n47), .ZN(n182) );
  NAND2_X1 U86 ( .A1(\mem[1][8] ), .A2(n374), .ZN(n47) );
  OAI21_X1 U87 ( .B1(n385), .B2(n38), .A(n48), .ZN(n183) );
  NAND2_X1 U88 ( .A1(\mem[1][9] ), .A2(n374), .ZN(n48) );
  OAI21_X1 U89 ( .B1(n384), .B2(n38), .A(n49), .ZN(n184) );
  NAND2_X1 U90 ( .A1(\mem[1][10] ), .A2(n374), .ZN(n49) );
  OAI21_X1 U91 ( .B1(n383), .B2(n38), .A(n50), .ZN(n185) );
  NAND2_X1 U92 ( .A1(\mem[1][11] ), .A2(n374), .ZN(n50) );
  OAI21_X1 U93 ( .B1(n382), .B2(n38), .A(n51), .ZN(n186) );
  NAND2_X1 U94 ( .A1(\mem[1][12] ), .A2(n374), .ZN(n51) );
  OAI21_X1 U95 ( .B1(n381), .B2(n38), .A(n52), .ZN(n187) );
  NAND2_X1 U96 ( .A1(\mem[1][13] ), .A2(n374), .ZN(n52) );
  OAI21_X1 U97 ( .B1(n380), .B2(n38), .A(n53), .ZN(n188) );
  NAND2_X1 U98 ( .A1(\mem[1][14] ), .A2(n374), .ZN(n53) );
  OAI21_X1 U99 ( .B1(n387), .B2(n55), .A(n63), .ZN(n197) );
  NAND2_X1 U100 ( .A1(\mem[2][7] ), .A2(n373), .ZN(n63) );
  OAI21_X1 U101 ( .B1(n386), .B2(n55), .A(n64), .ZN(n198) );
  NAND2_X1 U102 ( .A1(\mem[2][8] ), .A2(n55), .ZN(n64) );
  OAI21_X1 U103 ( .B1(n385), .B2(n55), .A(n65), .ZN(n199) );
  NAND2_X1 U104 ( .A1(\mem[2][9] ), .A2(n55), .ZN(n65) );
  OAI21_X1 U105 ( .B1(n384), .B2(n55), .A(n66), .ZN(n200) );
  NAND2_X1 U106 ( .A1(\mem[2][10] ), .A2(n55), .ZN(n66) );
  OAI21_X1 U107 ( .B1(n383), .B2(n55), .A(n67), .ZN(n201) );
  NAND2_X1 U108 ( .A1(\mem[2][11] ), .A2(n55), .ZN(n67) );
  OAI21_X1 U109 ( .B1(n382), .B2(n55), .A(n68), .ZN(n202) );
  NAND2_X1 U110 ( .A1(\mem[2][12] ), .A2(n55), .ZN(n68) );
  OAI21_X1 U111 ( .B1(n381), .B2(n55), .A(n69), .ZN(n203) );
  NAND2_X1 U112 ( .A1(\mem[2][13] ), .A2(n55), .ZN(n69) );
  OAI21_X1 U113 ( .B1(n380), .B2(n55), .A(n70), .ZN(n204) );
  NAND2_X1 U114 ( .A1(\mem[2][14] ), .A2(n55), .ZN(n70) );
  OAI21_X1 U115 ( .B1(n387), .B2(n89), .A(n97), .ZN(n229) );
  NAND2_X1 U116 ( .A1(\mem[4][7] ), .A2(n371), .ZN(n97) );
  OAI21_X1 U117 ( .B1(n386), .B2(n371), .A(n98), .ZN(n230) );
  NAND2_X1 U118 ( .A1(\mem[4][8] ), .A2(n371), .ZN(n98) );
  OAI21_X1 U119 ( .B1(n385), .B2(n89), .A(n99), .ZN(n231) );
  NAND2_X1 U120 ( .A1(\mem[4][9] ), .A2(n371), .ZN(n99) );
  OAI21_X1 U121 ( .B1(n384), .B2(n89), .A(n100), .ZN(n232) );
  NAND2_X1 U122 ( .A1(\mem[4][10] ), .A2(n371), .ZN(n100) );
  OAI21_X1 U123 ( .B1(n383), .B2(n89), .A(n101), .ZN(n233) );
  NAND2_X1 U124 ( .A1(\mem[4][11] ), .A2(n371), .ZN(n101) );
  OAI21_X1 U125 ( .B1(n382), .B2(n89), .A(n102), .ZN(n234) );
  NAND2_X1 U126 ( .A1(\mem[4][12] ), .A2(n371), .ZN(n102) );
  OAI21_X1 U127 ( .B1(n381), .B2(n89), .A(n103), .ZN(n235) );
  NAND2_X1 U128 ( .A1(\mem[4][13] ), .A2(n371), .ZN(n103) );
  OAI21_X1 U129 ( .B1(n380), .B2(n89), .A(n104), .ZN(n236) );
  NAND2_X1 U130 ( .A1(\mem[4][14] ), .A2(n371), .ZN(n104) );
  OAI21_X1 U131 ( .B1(n20), .B2(n386), .A(n29), .ZN(n166) );
  NAND2_X1 U132 ( .A1(\mem[0][8] ), .A2(n375), .ZN(n29) );
  OAI21_X1 U133 ( .B1(n20), .B2(n385), .A(n30), .ZN(n167) );
  NAND2_X1 U134 ( .A1(\mem[0][9] ), .A2(n20), .ZN(n30) );
  OAI21_X1 U135 ( .B1(n375), .B2(n384), .A(n31), .ZN(n168) );
  NAND2_X1 U136 ( .A1(\mem[0][10] ), .A2(n20), .ZN(n31) );
  OAI21_X1 U137 ( .B1(n20), .B2(n383), .A(n32), .ZN(n169) );
  NAND2_X1 U138 ( .A1(\mem[0][11] ), .A2(n20), .ZN(n32) );
  OAI21_X1 U139 ( .B1(n20), .B2(n382), .A(n33), .ZN(n170) );
  NAND2_X1 U140 ( .A1(\mem[0][12] ), .A2(n20), .ZN(n33) );
  OAI21_X1 U141 ( .B1(n20), .B2(n381), .A(n34), .ZN(n171) );
  NAND2_X1 U142 ( .A1(\mem[0][13] ), .A2(n20), .ZN(n34) );
  OAI21_X1 U143 ( .B1(n20), .B2(n380), .A(n35), .ZN(n172) );
  NAND2_X1 U144 ( .A1(\mem[0][14] ), .A2(n20), .ZN(n35) );
  OAI21_X1 U145 ( .B1(n394), .B2(n38), .A(n39), .ZN(n174) );
  NAND2_X1 U146 ( .A1(\mem[1][0] ), .A2(n374), .ZN(n39) );
  OAI21_X1 U147 ( .B1(n393), .B2(n38), .A(n40), .ZN(n175) );
  NAND2_X1 U148 ( .A1(\mem[1][1] ), .A2(n374), .ZN(n40) );
  OAI21_X1 U149 ( .B1(n392), .B2(n38), .A(n41), .ZN(n176) );
  NAND2_X1 U150 ( .A1(\mem[1][2] ), .A2(n374), .ZN(n41) );
  OAI21_X1 U151 ( .B1(n391), .B2(n38), .A(n42), .ZN(n177) );
  NAND2_X1 U152 ( .A1(\mem[1][3] ), .A2(n374), .ZN(n42) );
  OAI21_X1 U153 ( .B1(n390), .B2(n38), .A(n43), .ZN(n178) );
  NAND2_X1 U154 ( .A1(\mem[1][4] ), .A2(n38), .ZN(n43) );
  OAI21_X1 U155 ( .B1(n389), .B2(n38), .A(n44), .ZN(n179) );
  NAND2_X1 U156 ( .A1(\mem[1][5] ), .A2(n38), .ZN(n44) );
  OAI21_X1 U157 ( .B1(n388), .B2(n38), .A(n45), .ZN(n180) );
  NAND2_X1 U158 ( .A1(\mem[1][6] ), .A2(n38), .ZN(n45) );
  OAI21_X1 U159 ( .B1(n379), .B2(n38), .A(n54), .ZN(n189) );
  NAND2_X1 U160 ( .A1(\mem[1][15] ), .A2(n374), .ZN(n54) );
  OAI21_X1 U161 ( .B1(n394), .B2(n373), .A(n56), .ZN(n190) );
  NAND2_X1 U162 ( .A1(\mem[2][0] ), .A2(n373), .ZN(n56) );
  OAI21_X1 U163 ( .B1(n393), .B2(n373), .A(n57), .ZN(n191) );
  NAND2_X1 U164 ( .A1(\mem[2][1] ), .A2(n55), .ZN(n57) );
  OAI21_X1 U165 ( .B1(n392), .B2(n373), .A(n58), .ZN(n192) );
  NAND2_X1 U166 ( .A1(\mem[2][2] ), .A2(n55), .ZN(n58) );
  OAI21_X1 U167 ( .B1(n391), .B2(n373), .A(n59), .ZN(n193) );
  NAND2_X1 U168 ( .A1(\mem[2][3] ), .A2(n55), .ZN(n59) );
  OAI21_X1 U169 ( .B1(n390), .B2(n373), .A(n60), .ZN(n194) );
  NAND2_X1 U170 ( .A1(\mem[2][4] ), .A2(n373), .ZN(n60) );
  OAI21_X1 U171 ( .B1(n389), .B2(n373), .A(n61), .ZN(n195) );
  NAND2_X1 U172 ( .A1(\mem[2][5] ), .A2(n373), .ZN(n61) );
  OAI21_X1 U173 ( .B1(n388), .B2(n373), .A(n62), .ZN(n196) );
  NAND2_X1 U174 ( .A1(\mem[2][6] ), .A2(n373), .ZN(n62) );
  OAI21_X1 U175 ( .B1(n379), .B2(n373), .A(n71), .ZN(n205) );
  NAND2_X1 U176 ( .A1(\mem[2][15] ), .A2(n373), .ZN(n71) );
  OAI21_X1 U177 ( .B1(n394), .B2(n72), .A(n73), .ZN(n206) );
  NAND2_X1 U178 ( .A1(\mem[3][0] ), .A2(n372), .ZN(n73) );
  OAI21_X1 U179 ( .B1(n393), .B2(n72), .A(n74), .ZN(n207) );
  NAND2_X1 U180 ( .A1(\mem[3][1] ), .A2(n372), .ZN(n74) );
  OAI21_X1 U181 ( .B1(n392), .B2(n72), .A(n75), .ZN(n208) );
  NAND2_X1 U182 ( .A1(\mem[3][2] ), .A2(n372), .ZN(n75) );
  OAI21_X1 U183 ( .B1(n391), .B2(n72), .A(n76), .ZN(n209) );
  NAND2_X1 U184 ( .A1(\mem[3][3] ), .A2(n372), .ZN(n76) );
  OAI21_X1 U185 ( .B1(n390), .B2(n72), .A(n77), .ZN(n210) );
  NAND2_X1 U186 ( .A1(\mem[3][4] ), .A2(n72), .ZN(n77) );
  OAI21_X1 U187 ( .B1(n389), .B2(n72), .A(n78), .ZN(n211) );
  NAND2_X1 U188 ( .A1(\mem[3][5] ), .A2(n72), .ZN(n78) );
  OAI21_X1 U189 ( .B1(n388), .B2(n72), .A(n79), .ZN(n212) );
  NAND2_X1 U190 ( .A1(\mem[3][6] ), .A2(n72), .ZN(n79) );
  OAI21_X1 U191 ( .B1(n379), .B2(n72), .A(n88), .ZN(n221) );
  NAND2_X1 U192 ( .A1(\mem[3][15] ), .A2(n372), .ZN(n88) );
  OAI21_X1 U193 ( .B1(n394), .B2(n89), .A(n90), .ZN(n222) );
  NAND2_X1 U194 ( .A1(\mem[4][0] ), .A2(n371), .ZN(n90) );
  OAI21_X1 U195 ( .B1(n393), .B2(n89), .A(n91), .ZN(n223) );
  NAND2_X1 U196 ( .A1(\mem[4][1] ), .A2(n371), .ZN(n91) );
  OAI21_X1 U197 ( .B1(n392), .B2(n89), .A(n92), .ZN(n224) );
  NAND2_X1 U198 ( .A1(\mem[4][2] ), .A2(n371), .ZN(n92) );
  OAI21_X1 U199 ( .B1(n391), .B2(n89), .A(n93), .ZN(n225) );
  NAND2_X1 U200 ( .A1(\mem[4][3] ), .A2(n371), .ZN(n93) );
  OAI21_X1 U201 ( .B1(n390), .B2(n89), .A(n94), .ZN(n226) );
  NAND2_X1 U202 ( .A1(\mem[4][4] ), .A2(n89), .ZN(n94) );
  OAI21_X1 U203 ( .B1(n389), .B2(n89), .A(n95), .ZN(n227) );
  NAND2_X1 U204 ( .A1(\mem[4][5] ), .A2(n89), .ZN(n95) );
  OAI21_X1 U205 ( .B1(n388), .B2(n89), .A(n96), .ZN(n228) );
  NAND2_X1 U206 ( .A1(\mem[4][6] ), .A2(n89), .ZN(n96) );
  OAI21_X1 U207 ( .B1(n379), .B2(n89), .A(n105), .ZN(n237) );
  NAND2_X1 U208 ( .A1(\mem[4][15] ), .A2(n371), .ZN(n105) );
  OAI21_X1 U209 ( .B1(n394), .B2(n107), .A(n108), .ZN(n238) );
  NAND2_X1 U210 ( .A1(\mem[5][0] ), .A2(n370), .ZN(n108) );
  OAI21_X1 U211 ( .B1(n393), .B2(n107), .A(n109), .ZN(n239) );
  NAND2_X1 U212 ( .A1(\mem[5][1] ), .A2(n370), .ZN(n109) );
  OAI21_X1 U213 ( .B1(n392), .B2(n107), .A(n110), .ZN(n240) );
  NAND2_X1 U214 ( .A1(\mem[5][2] ), .A2(n370), .ZN(n110) );
  OAI21_X1 U215 ( .B1(n391), .B2(n107), .A(n111), .ZN(n241) );
  NAND2_X1 U216 ( .A1(\mem[5][3] ), .A2(n370), .ZN(n111) );
  OAI21_X1 U217 ( .B1(n390), .B2(n107), .A(n112), .ZN(n242) );
  NAND2_X1 U218 ( .A1(\mem[5][4] ), .A2(n107), .ZN(n112) );
  OAI21_X1 U219 ( .B1(n389), .B2(n107), .A(n113), .ZN(n243) );
  NAND2_X1 U220 ( .A1(\mem[5][5] ), .A2(n107), .ZN(n113) );
  OAI21_X1 U221 ( .B1(n388), .B2(n107), .A(n114), .ZN(n244) );
  NAND2_X1 U222 ( .A1(\mem[5][6] ), .A2(n107), .ZN(n114) );
  OAI21_X1 U223 ( .B1(n379), .B2(n107), .A(n123), .ZN(n253) );
  NAND2_X1 U224 ( .A1(\mem[5][15] ), .A2(n370), .ZN(n123) );
  OAI21_X1 U225 ( .B1(n394), .B2(n124), .A(n125), .ZN(n254) );
  NAND2_X1 U226 ( .A1(\mem[6][0] ), .A2(n369), .ZN(n125) );
  OAI21_X1 U227 ( .B1(n393), .B2(n124), .A(n126), .ZN(n255) );
  NAND2_X1 U228 ( .A1(\mem[6][1] ), .A2(n369), .ZN(n126) );
  OAI21_X1 U229 ( .B1(n392), .B2(n124), .A(n127), .ZN(n256) );
  NAND2_X1 U230 ( .A1(\mem[6][2] ), .A2(n369), .ZN(n127) );
  OAI21_X1 U231 ( .B1(n391), .B2(n124), .A(n128), .ZN(n257) );
  NAND2_X1 U232 ( .A1(\mem[6][3] ), .A2(n369), .ZN(n128) );
  OAI21_X1 U233 ( .B1(n390), .B2(n124), .A(n129), .ZN(n258) );
  NAND2_X1 U234 ( .A1(\mem[6][4] ), .A2(n124), .ZN(n129) );
  OAI21_X1 U235 ( .B1(n389), .B2(n124), .A(n130), .ZN(n259) );
  NAND2_X1 U236 ( .A1(\mem[6][5] ), .A2(n124), .ZN(n130) );
  OAI21_X1 U237 ( .B1(n388), .B2(n124), .A(n131), .ZN(n260) );
  NAND2_X1 U238 ( .A1(\mem[6][6] ), .A2(n124), .ZN(n131) );
  OAI21_X1 U239 ( .B1(n379), .B2(n124), .A(n140), .ZN(n269) );
  NAND2_X1 U240 ( .A1(\mem[6][15] ), .A2(n369), .ZN(n140) );
  OAI21_X1 U241 ( .B1(n394), .B2(n141), .A(n142), .ZN(n270) );
  NAND2_X1 U242 ( .A1(\mem[7][0] ), .A2(n368), .ZN(n142) );
  OAI21_X1 U243 ( .B1(n393), .B2(n141), .A(n143), .ZN(n271) );
  NAND2_X1 U244 ( .A1(\mem[7][1] ), .A2(n368), .ZN(n143) );
  OAI21_X1 U245 ( .B1(n392), .B2(n141), .A(n144), .ZN(n272) );
  NAND2_X1 U246 ( .A1(\mem[7][2] ), .A2(n368), .ZN(n144) );
  OAI21_X1 U247 ( .B1(n391), .B2(n141), .A(n145), .ZN(n273) );
  NAND2_X1 U248 ( .A1(\mem[7][3] ), .A2(n368), .ZN(n145) );
  OAI21_X1 U249 ( .B1(n390), .B2(n141), .A(n146), .ZN(n274) );
  NAND2_X1 U250 ( .A1(\mem[7][4] ), .A2(n141), .ZN(n146) );
  OAI21_X1 U251 ( .B1(n389), .B2(n141), .A(n147), .ZN(n275) );
  NAND2_X1 U252 ( .A1(\mem[7][5] ), .A2(n141), .ZN(n147) );
  OAI21_X1 U253 ( .B1(n388), .B2(n141), .A(n148), .ZN(n276) );
  NAND2_X1 U254 ( .A1(\mem[7][6] ), .A2(n141), .ZN(n148) );
  OAI21_X1 U255 ( .B1(n379), .B2(n141), .A(n157), .ZN(n285) );
  NAND2_X1 U256 ( .A1(\mem[7][15] ), .A2(n368), .ZN(n157) );
  OAI21_X1 U257 ( .B1(n375), .B2(n394), .A(n21), .ZN(n158) );
  NAND2_X1 U258 ( .A1(\mem[0][0] ), .A2(n20), .ZN(n21) );
  OAI21_X1 U259 ( .B1(n375), .B2(n393), .A(n22), .ZN(n159) );
  NAND2_X1 U260 ( .A1(\mem[0][1] ), .A2(n20), .ZN(n22) );
  OAI21_X1 U261 ( .B1(n375), .B2(n392), .A(n23), .ZN(n160) );
  NAND2_X1 U262 ( .A1(\mem[0][2] ), .A2(n20), .ZN(n23) );
  OAI21_X1 U263 ( .B1(n375), .B2(n391), .A(n24), .ZN(n161) );
  NAND2_X1 U264 ( .A1(\mem[0][3] ), .A2(n20), .ZN(n24) );
  OAI21_X1 U265 ( .B1(n375), .B2(n390), .A(n25), .ZN(n162) );
  NAND2_X1 U266 ( .A1(\mem[0][4] ), .A2(n375), .ZN(n25) );
  OAI21_X1 U267 ( .B1(n375), .B2(n389), .A(n26), .ZN(n163) );
  NAND2_X1 U268 ( .A1(\mem[0][5] ), .A2(n375), .ZN(n26) );
  OAI21_X1 U269 ( .B1(n375), .B2(n388), .A(n27), .ZN(n164) );
  NAND2_X1 U270 ( .A1(\mem[0][6] ), .A2(n375), .ZN(n27) );
  OAI21_X1 U271 ( .B1(n375), .B2(n387), .A(n28), .ZN(n165) );
  NAND2_X1 U272 ( .A1(\mem[0][7] ), .A2(n375), .ZN(n28) );
  OAI21_X1 U273 ( .B1(n375), .B2(n379), .A(n36), .ZN(n173) );
  NAND2_X1 U274 ( .A1(\mem[0][15] ), .A2(n20), .ZN(n36) );
  INV_X1 U275 ( .A(N11), .ZN(n377) );
  INV_X1 U276 ( .A(data_in[0]), .ZN(n394) );
  INV_X1 U277 ( .A(data_in[1]), .ZN(n393) );
  INV_X1 U278 ( .A(data_in[2]), .ZN(n392) );
  INV_X1 U279 ( .A(data_in[3]), .ZN(n391) );
  INV_X1 U288 ( .A(data_in[4]), .ZN(n390) );
  INV_X1 U289 ( .A(data_in[5]), .ZN(n389) );
  INV_X1 U290 ( .A(data_in[6]), .ZN(n388) );
  INV_X1 U291 ( .A(data_in[7]), .ZN(n387) );
  INV_X1 U292 ( .A(data_in[8]), .ZN(n386) );
  INV_X1 U293 ( .A(data_in[9]), .ZN(n385) );
  INV_X1 U294 ( .A(data_in[10]), .ZN(n384) );
  INV_X1 U295 ( .A(data_in[11]), .ZN(n383) );
  INV_X1 U296 ( .A(data_in[12]), .ZN(n382) );
  INV_X1 U297 ( .A(data_in[13]), .ZN(n381) );
  INV_X1 U298 ( .A(data_in[14]), .ZN(n380) );
  INV_X1 U299 ( .A(data_in[15]), .ZN(n379) );
  MUX2_X1 U300 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n366), .Z(n2) );
  MUX2_X1 U301 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n367), .Z(n3) );
  MUX2_X1 U302 ( .A(n3), .B(n2), .S(n364), .Z(n4) );
  MUX2_X1 U303 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n365), .Z(n5) );
  MUX2_X1 U304 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n366), .Z(n6) );
  MUX2_X1 U305 ( .A(n6), .B(n5), .S(n364), .Z(n7) );
  MUX2_X1 U306 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n365), .Z(n8) );
  MUX2_X1 U307 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n365), .Z(n9) );
  MUX2_X1 U308 ( .A(n9), .B(n8), .S(n364), .Z(n10) );
  MUX2_X1 U309 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n365), .Z(n11) );
  MUX2_X1 U310 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n365), .Z(n12) );
  MUX2_X1 U311 ( .A(n12), .B(n11), .S(N11), .Z(n13) );
  MUX2_X1 U312 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n365), .Z(n14) );
  MUX2_X1 U313 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n365), .Z(n15) );
  MUX2_X1 U314 ( .A(n15), .B(n14), .S(n364), .Z(n16) );
  MUX2_X1 U315 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n365), .Z(n17) );
  MUX2_X1 U316 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n365), .Z(n18) );
  MUX2_X1 U317 ( .A(n18), .B(n17), .S(n364), .Z(n19) );
  MUX2_X1 U318 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n365), .Z(n286) );
  MUX2_X1 U319 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n365), .Z(n287) );
  MUX2_X1 U320 ( .A(n287), .B(n286), .S(N11), .Z(n288) );
  MUX2_X1 U321 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n365), .Z(n289) );
  MUX2_X1 U322 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n365), .Z(n290) );
  MUX2_X1 U323 ( .A(n290), .B(n289), .S(N11), .Z(n291) );
  MUX2_X1 U324 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n366), .Z(n292) );
  MUX2_X1 U325 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n366), .Z(n293) );
  MUX2_X1 U326 ( .A(n293), .B(n292), .S(n364), .Z(n294) );
  MUX2_X1 U327 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n367), .Z(n295) );
  MUX2_X1 U328 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n365), .Z(n296) );
  MUX2_X1 U329 ( .A(n296), .B(n295), .S(n364), .Z(n297) );
  MUX2_X1 U330 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n367), .Z(n298) );
  MUX2_X1 U331 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n367), .Z(n299) );
  MUX2_X1 U332 ( .A(n299), .B(n298), .S(n364), .Z(n300) );
  MUX2_X1 U333 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n365), .Z(n301) );
  MUX2_X1 U334 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n366), .Z(n302) );
  MUX2_X1 U335 ( .A(n302), .B(n301), .S(n364), .Z(n303) );
  MUX2_X1 U336 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n365), .Z(n304) );
  MUX2_X1 U337 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n365), .Z(n305) );
  MUX2_X1 U338 ( .A(n305), .B(n304), .S(n364), .Z(n306) );
  MUX2_X1 U339 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n366), .Z(n307) );
  MUX2_X1 U340 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n367), .Z(n308) );
  MUX2_X1 U341 ( .A(n308), .B(n307), .S(n364), .Z(n309) );
  MUX2_X1 U342 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n366), .Z(n310) );
  MUX2_X1 U343 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n366), .Z(n311) );
  MUX2_X1 U344 ( .A(n311), .B(n310), .S(n364), .Z(n312) );
  MUX2_X1 U345 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n365), .Z(n313) );
  MUX2_X1 U346 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n367), .Z(n314) );
  MUX2_X1 U347 ( .A(n314), .B(n313), .S(n364), .Z(n315) );
  MUX2_X1 U348 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n367), .Z(n316) );
  MUX2_X1 U349 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n366), .Z(n317) );
  MUX2_X1 U350 ( .A(n317), .B(n316), .S(n364), .Z(n318) );
  MUX2_X1 U351 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n367), .Z(n319) );
  MUX2_X1 U352 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n365), .Z(n320) );
  MUX2_X1 U353 ( .A(n320), .B(n319), .S(n364), .Z(n321) );
  MUX2_X1 U354 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n365), .Z(n322) );
  MUX2_X1 U355 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n367), .Z(n323) );
  MUX2_X1 U356 ( .A(n323), .B(n322), .S(n364), .Z(n324) );
  MUX2_X1 U357 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n366), .Z(n325) );
  MUX2_X1 U358 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n365), .Z(n326) );
  MUX2_X1 U359 ( .A(n326), .B(n325), .S(n364), .Z(n327) );
  MUX2_X1 U360 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n366), .Z(n328) );
  MUX2_X1 U361 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n366), .Z(n329) );
  MUX2_X1 U362 ( .A(n329), .B(n328), .S(n364), .Z(n330) );
  MUX2_X1 U363 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n366), .Z(n331) );
  MUX2_X1 U364 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n366), .Z(n332) );
  MUX2_X1 U365 ( .A(n332), .B(n331), .S(N11), .Z(n333) );
  MUX2_X1 U366 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n366), .Z(n334) );
  MUX2_X1 U367 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n366), .Z(n335) );
  MUX2_X1 U368 ( .A(n335), .B(n334), .S(n364), .Z(n336) );
  MUX2_X1 U369 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n366), .Z(n337) );
  MUX2_X1 U370 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n366), .Z(n338) );
  MUX2_X1 U371 ( .A(n338), .B(n337), .S(N11), .Z(n339) );
  MUX2_X1 U372 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n366), .Z(n340) );
  MUX2_X1 U373 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n366), .Z(n341) );
  MUX2_X1 U374 ( .A(n341), .B(n340), .S(n364), .Z(n342) );
  MUX2_X1 U375 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n366), .Z(n343) );
  MUX2_X1 U376 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n366), .Z(n344) );
  MUX2_X1 U377 ( .A(n344), .B(n343), .S(N11), .Z(n345) );
  MUX2_X1 U378 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n367), .Z(n346) );
  MUX2_X1 U379 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n367), .Z(n347) );
  MUX2_X1 U380 ( .A(n347), .B(n346), .S(n364), .Z(n348) );
  MUX2_X1 U381 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n367), .Z(n349) );
  MUX2_X1 U382 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n367), .Z(n350) );
  MUX2_X1 U383 ( .A(n350), .B(n349), .S(N11), .Z(n351) );
  MUX2_X1 U384 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n367), .Z(n352) );
  MUX2_X1 U385 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n367), .Z(n353) );
  MUX2_X1 U386 ( .A(n353), .B(n352), .S(n364), .Z(n354) );
  MUX2_X1 U387 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n367), .Z(n355) );
  MUX2_X1 U388 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n367), .Z(n356) );
  MUX2_X1 U389 ( .A(n356), .B(n355), .S(N11), .Z(n357) );
  MUX2_X1 U390 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n367), .Z(n358) );
  MUX2_X1 U391 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n367), .Z(n359) );
  MUX2_X1 U392 ( .A(n359), .B(n358), .S(n364), .Z(n360) );
  MUX2_X1 U393 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n367), .Z(n361) );
  MUX2_X1 U394 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n367), .Z(n362) );
  MUX2_X1 U395 ( .A(n362), .B(n361), .S(N11), .Z(n363) );
endmodule


module memory_WIDTH16_SIZE8_LOGSIZE3_8 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] ,
         \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][15] , \mem[6][14] , \mem[6][13] ,
         \mem[6][12] , \mem[6][11] , \mem[6][10] , \mem[6][9] , \mem[6][8] ,
         \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] ,
         \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[5][15] , \mem[5][14] ,
         \mem[5][13] , \mem[5][12] , \mem[5][11] , \mem[5][10] , \mem[5][9] ,
         \mem[5][8] , \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] ,
         \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][15] ,
         \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] , \mem[4][10] ,
         \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N13, N14, N16,
         N18, N20, N22, N24, N25, N26, N27, N28, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[15]  ( .D(N13), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N14), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N16), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N18), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[8]  ( .D(N20), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N22), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N24), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N25), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N26), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N28), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][15]  ( .D(n394), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n395), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n396), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n397), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n398), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n399), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n400), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n401), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n402), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n403), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n404), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n405), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n406), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n407), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n408), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n409), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n410), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n411), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n412), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n413), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n414), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n415), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n416), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n417), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n418), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n419), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n420), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n421), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n422), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n423), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n424), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n425), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n426), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n427), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n428), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n429), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n430), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n431), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n432), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n433), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n434), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n435), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n436), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n437), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n438), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n439), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n440), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n441), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n442), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n443), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n444), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n445), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n446), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n447), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n448), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n449), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n450), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n451), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n452), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n453), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n454), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n455), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n456), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n457), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n458), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n459), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n460), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n461), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n462), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n463), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n464), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n465), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n466), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n467), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n468), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n469), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n470), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n471), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n472), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n473), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n474), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n475), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n476), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n477), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n478), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n479), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n480), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n481), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n482), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n483), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n484), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n485), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n486), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n487), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n488), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n489), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n490), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n491), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n492), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n493), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n494), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n495), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n496), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n497), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n498), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n499), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n500), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n501), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n502), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n503), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n504), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n505), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n506), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n507), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n508), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n509), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n510), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n511), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n512), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n513), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n514), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n515), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n516), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n517), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n518), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n519), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n520), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n521), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U280 ( .A1(n375), .A2(n376), .A3(n642), .ZN(n659) );
  NAND3_X1 U281 ( .A1(n642), .A2(n376), .A3(N10), .ZN(n641) );
  NAND3_X1 U282 ( .A1(n642), .A2(n375), .A3(N11), .ZN(n624) );
  NAND3_X1 U283 ( .A1(N10), .A2(n642), .A3(N11), .ZN(n607) );
  NAND3_X1 U284 ( .A1(n375), .A2(n376), .A3(n573), .ZN(n590) );
  NAND3_X1 U285 ( .A1(N10), .A2(n376), .A3(n573), .ZN(n572) );
  NAND3_X1 U286 ( .A1(N11), .A2(n375), .A3(n573), .ZN(n555) );
  NAND3_X1 U287 ( .A1(N11), .A2(N10), .A3(n573), .ZN(n538) );
  DFF_X1 \data_out_reg[1]  ( .D(N27), .CK(clk), .Q(data_out[1]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n350), .SI(n347), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n302), .SI(n299), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n338), .SI(n335), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n326), .SI(n323), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n314), .SI(n311), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  BUF_X1 U3 ( .A(N10), .Z(n365) );
  BUF_X1 U4 ( .A(N10), .Z(n366) );
  BUF_X1 U5 ( .A(n659), .Z(n374) );
  BUF_X1 U6 ( .A(n624), .Z(n372) );
  BUF_X1 U7 ( .A(n607), .Z(n371) );
  BUF_X1 U8 ( .A(n590), .Z(n370) );
  BUF_X1 U9 ( .A(n555), .Z(n368) );
  BUF_X1 U10 ( .A(n538), .Z(n367) );
  BUF_X1 U11 ( .A(n572), .Z(n369) );
  BUF_X1 U12 ( .A(n641), .Z(n373) );
  BUF_X1 U13 ( .A(N10), .Z(n364) );
  BUF_X1 U14 ( .A(N11), .Z(n363) );
  NOR2_X1 U15 ( .A1(n377), .A2(N12), .ZN(n642) );
  INV_X1 U16 ( .A(wr_en), .ZN(n377) );
  AND2_X1 U17 ( .A1(N12), .A2(wr_en), .ZN(n573) );
  OAI21_X1 U18 ( .B1(n386), .B2(n607), .A(n599), .ZN(n466) );
  NAND2_X1 U19 ( .A1(\mem[3][7] ), .A2(n371), .ZN(n599) );
  OAI21_X1 U20 ( .B1(n385), .B2(n371), .A(n598), .ZN(n465) );
  NAND2_X1 U21 ( .A1(\mem[3][8] ), .A2(n371), .ZN(n598) );
  OAI21_X1 U22 ( .B1(n384), .B2(n607), .A(n597), .ZN(n464) );
  NAND2_X1 U23 ( .A1(\mem[3][9] ), .A2(n371), .ZN(n597) );
  OAI21_X1 U24 ( .B1(n383), .B2(n607), .A(n596), .ZN(n463) );
  NAND2_X1 U25 ( .A1(\mem[3][10] ), .A2(n371), .ZN(n596) );
  OAI21_X1 U26 ( .B1(n382), .B2(n607), .A(n595), .ZN(n462) );
  NAND2_X1 U27 ( .A1(\mem[3][11] ), .A2(n371), .ZN(n595) );
  OAI21_X1 U28 ( .B1(n381), .B2(n607), .A(n594), .ZN(n461) );
  NAND2_X1 U29 ( .A1(\mem[3][12] ), .A2(n371), .ZN(n594) );
  OAI21_X1 U30 ( .B1(n380), .B2(n607), .A(n593), .ZN(n460) );
  NAND2_X1 U31 ( .A1(\mem[3][13] ), .A2(n371), .ZN(n593) );
  OAI21_X1 U32 ( .B1(n379), .B2(n607), .A(n592), .ZN(n459) );
  NAND2_X1 U33 ( .A1(\mem[3][14] ), .A2(n371), .ZN(n592) );
  OAI21_X1 U34 ( .B1(n386), .B2(n572), .A(n564), .ZN(n434) );
  NAND2_X1 U35 ( .A1(\mem[5][7] ), .A2(n369), .ZN(n564) );
  OAI21_X1 U36 ( .B1(n385), .B2(n572), .A(n563), .ZN(n433) );
  NAND2_X1 U37 ( .A1(\mem[5][8] ), .A2(n572), .ZN(n563) );
  OAI21_X1 U38 ( .B1(n384), .B2(n572), .A(n562), .ZN(n432) );
  NAND2_X1 U39 ( .A1(\mem[5][9] ), .A2(n572), .ZN(n562) );
  OAI21_X1 U40 ( .B1(n383), .B2(n572), .A(n561), .ZN(n431) );
  NAND2_X1 U41 ( .A1(\mem[5][10] ), .A2(n572), .ZN(n561) );
  OAI21_X1 U42 ( .B1(n382), .B2(n572), .A(n560), .ZN(n430) );
  NAND2_X1 U43 ( .A1(\mem[5][11] ), .A2(n572), .ZN(n560) );
  OAI21_X1 U44 ( .B1(n381), .B2(n572), .A(n559), .ZN(n429) );
  NAND2_X1 U45 ( .A1(\mem[5][12] ), .A2(n572), .ZN(n559) );
  OAI21_X1 U46 ( .B1(n380), .B2(n572), .A(n558), .ZN(n428) );
  NAND2_X1 U47 ( .A1(\mem[5][13] ), .A2(n572), .ZN(n558) );
  OAI21_X1 U48 ( .B1(n379), .B2(n572), .A(n557), .ZN(n427) );
  NAND2_X1 U49 ( .A1(\mem[5][14] ), .A2(n572), .ZN(n557) );
  OAI21_X1 U50 ( .B1(n386), .B2(n538), .A(n530), .ZN(n402) );
  NAND2_X1 U51 ( .A1(\mem[7][7] ), .A2(n367), .ZN(n530) );
  OAI21_X1 U52 ( .B1(n385), .B2(n367), .A(n529), .ZN(n401) );
  NAND2_X1 U53 ( .A1(\mem[7][8] ), .A2(n367), .ZN(n529) );
  OAI21_X1 U54 ( .B1(n384), .B2(n538), .A(n528), .ZN(n400) );
  NAND2_X1 U55 ( .A1(\mem[7][9] ), .A2(n367), .ZN(n528) );
  OAI21_X1 U56 ( .B1(n383), .B2(n538), .A(n527), .ZN(n399) );
  NAND2_X1 U57 ( .A1(\mem[7][10] ), .A2(n367), .ZN(n527) );
  OAI21_X1 U58 ( .B1(n382), .B2(n538), .A(n526), .ZN(n398) );
  NAND2_X1 U59 ( .A1(\mem[7][11] ), .A2(n367), .ZN(n526) );
  OAI21_X1 U60 ( .B1(n381), .B2(n538), .A(n525), .ZN(n397) );
  NAND2_X1 U61 ( .A1(\mem[7][12] ), .A2(n367), .ZN(n525) );
  OAI21_X1 U62 ( .B1(n380), .B2(n538), .A(n524), .ZN(n396) );
  NAND2_X1 U63 ( .A1(\mem[7][13] ), .A2(n367), .ZN(n524) );
  OAI21_X1 U64 ( .B1(n379), .B2(n538), .A(n523), .ZN(n395) );
  NAND2_X1 U65 ( .A1(\mem[7][14] ), .A2(n367), .ZN(n523) );
  OAI21_X1 U66 ( .B1(n386), .B2(n373), .A(n633), .ZN(n498) );
  NAND2_X1 U67 ( .A1(\mem[1][7] ), .A2(n373), .ZN(n633) );
  OAI21_X1 U68 ( .B1(n385), .B2(n373), .A(n632), .ZN(n497) );
  NAND2_X1 U69 ( .A1(\mem[1][8] ), .A2(n641), .ZN(n632) );
  OAI21_X1 U70 ( .B1(n384), .B2(n373), .A(n631), .ZN(n496) );
  NAND2_X1 U71 ( .A1(\mem[1][9] ), .A2(n641), .ZN(n631) );
  OAI21_X1 U72 ( .B1(n383), .B2(n373), .A(n630), .ZN(n495) );
  NAND2_X1 U73 ( .A1(\mem[1][10] ), .A2(n641), .ZN(n630) );
  OAI21_X1 U74 ( .B1(n382), .B2(n373), .A(n629), .ZN(n494) );
  NAND2_X1 U75 ( .A1(\mem[1][11] ), .A2(n641), .ZN(n629) );
  OAI21_X1 U76 ( .B1(n381), .B2(n373), .A(n628), .ZN(n493) );
  NAND2_X1 U77 ( .A1(\mem[1][12] ), .A2(n641), .ZN(n628) );
  OAI21_X1 U78 ( .B1(n380), .B2(n373), .A(n627), .ZN(n492) );
  NAND2_X1 U79 ( .A1(\mem[1][13] ), .A2(n641), .ZN(n627) );
  OAI21_X1 U80 ( .B1(n379), .B2(n373), .A(n626), .ZN(n491) );
  NAND2_X1 U81 ( .A1(\mem[1][14] ), .A2(n641), .ZN(n626) );
  OAI21_X1 U82 ( .B1(n386), .B2(n555), .A(n547), .ZN(n418) );
  NAND2_X1 U83 ( .A1(\mem[6][7] ), .A2(n368), .ZN(n547) );
  OAI21_X1 U84 ( .B1(n385), .B2(n368), .A(n546), .ZN(n417) );
  NAND2_X1 U85 ( .A1(\mem[6][8] ), .A2(n368), .ZN(n546) );
  OAI21_X1 U86 ( .B1(n384), .B2(n555), .A(n545), .ZN(n416) );
  NAND2_X1 U87 ( .A1(\mem[6][9] ), .A2(n368), .ZN(n545) );
  OAI21_X1 U88 ( .B1(n383), .B2(n555), .A(n544), .ZN(n415) );
  NAND2_X1 U89 ( .A1(\mem[6][10] ), .A2(n368), .ZN(n544) );
  OAI21_X1 U90 ( .B1(n382), .B2(n555), .A(n543), .ZN(n414) );
  NAND2_X1 U91 ( .A1(\mem[6][11] ), .A2(n368), .ZN(n543) );
  OAI21_X1 U92 ( .B1(n381), .B2(n555), .A(n542), .ZN(n413) );
  NAND2_X1 U93 ( .A1(\mem[6][12] ), .A2(n368), .ZN(n542) );
  OAI21_X1 U94 ( .B1(n380), .B2(n555), .A(n541), .ZN(n412) );
  NAND2_X1 U95 ( .A1(\mem[6][13] ), .A2(n368), .ZN(n541) );
  OAI21_X1 U96 ( .B1(n379), .B2(n555), .A(n540), .ZN(n411) );
  NAND2_X1 U97 ( .A1(\mem[6][14] ), .A2(n368), .ZN(n540) );
  OAI21_X1 U98 ( .B1(n386), .B2(n624), .A(n616), .ZN(n482) );
  NAND2_X1 U99 ( .A1(\mem[2][7] ), .A2(n372), .ZN(n616) );
  OAI21_X1 U100 ( .B1(n385), .B2(n372), .A(n615), .ZN(n481) );
  NAND2_X1 U101 ( .A1(\mem[2][8] ), .A2(n372), .ZN(n615) );
  OAI21_X1 U102 ( .B1(n384), .B2(n624), .A(n614), .ZN(n480) );
  NAND2_X1 U103 ( .A1(\mem[2][9] ), .A2(n372), .ZN(n614) );
  OAI21_X1 U104 ( .B1(n383), .B2(n624), .A(n613), .ZN(n479) );
  NAND2_X1 U105 ( .A1(\mem[2][10] ), .A2(n372), .ZN(n613) );
  OAI21_X1 U106 ( .B1(n382), .B2(n624), .A(n612), .ZN(n478) );
  NAND2_X1 U107 ( .A1(\mem[2][11] ), .A2(n372), .ZN(n612) );
  OAI21_X1 U108 ( .B1(n381), .B2(n624), .A(n611), .ZN(n477) );
  NAND2_X1 U109 ( .A1(\mem[2][12] ), .A2(n372), .ZN(n611) );
  OAI21_X1 U110 ( .B1(n380), .B2(n624), .A(n610), .ZN(n476) );
  NAND2_X1 U111 ( .A1(\mem[2][13] ), .A2(n372), .ZN(n610) );
  OAI21_X1 U112 ( .B1(n379), .B2(n624), .A(n609), .ZN(n475) );
  NAND2_X1 U113 ( .A1(\mem[2][14] ), .A2(n372), .ZN(n609) );
  OAI21_X1 U114 ( .B1(n386), .B2(n590), .A(n582), .ZN(n450) );
  NAND2_X1 U115 ( .A1(\mem[4][7] ), .A2(n370), .ZN(n582) );
  OAI21_X1 U116 ( .B1(n385), .B2(n370), .A(n581), .ZN(n449) );
  NAND2_X1 U117 ( .A1(\mem[4][8] ), .A2(n370), .ZN(n581) );
  OAI21_X1 U118 ( .B1(n384), .B2(n590), .A(n580), .ZN(n448) );
  NAND2_X1 U119 ( .A1(\mem[4][9] ), .A2(n370), .ZN(n580) );
  OAI21_X1 U120 ( .B1(n383), .B2(n590), .A(n579), .ZN(n447) );
  NAND2_X1 U121 ( .A1(\mem[4][10] ), .A2(n370), .ZN(n579) );
  OAI21_X1 U122 ( .B1(n382), .B2(n590), .A(n578), .ZN(n446) );
  NAND2_X1 U123 ( .A1(\mem[4][11] ), .A2(n370), .ZN(n578) );
  OAI21_X1 U124 ( .B1(n381), .B2(n590), .A(n577), .ZN(n445) );
  NAND2_X1 U125 ( .A1(\mem[4][12] ), .A2(n370), .ZN(n577) );
  OAI21_X1 U126 ( .B1(n380), .B2(n590), .A(n576), .ZN(n444) );
  NAND2_X1 U127 ( .A1(\mem[4][13] ), .A2(n370), .ZN(n576) );
  OAI21_X1 U128 ( .B1(n379), .B2(n590), .A(n575), .ZN(n443) );
  NAND2_X1 U129 ( .A1(\mem[4][14] ), .A2(n370), .ZN(n575) );
  OAI21_X1 U130 ( .B1(n659), .B2(n385), .A(n650), .ZN(n513) );
  NAND2_X1 U131 ( .A1(\mem[0][8] ), .A2(n374), .ZN(n650) );
  OAI21_X1 U132 ( .B1(n659), .B2(n384), .A(n649), .ZN(n512) );
  NAND2_X1 U133 ( .A1(\mem[0][9] ), .A2(n659), .ZN(n649) );
  OAI21_X1 U134 ( .B1(n374), .B2(n383), .A(n648), .ZN(n511) );
  NAND2_X1 U135 ( .A1(\mem[0][10] ), .A2(n659), .ZN(n648) );
  OAI21_X1 U136 ( .B1(n659), .B2(n382), .A(n647), .ZN(n510) );
  NAND2_X1 U137 ( .A1(\mem[0][11] ), .A2(n659), .ZN(n647) );
  OAI21_X1 U138 ( .B1(n659), .B2(n381), .A(n646), .ZN(n509) );
  NAND2_X1 U139 ( .A1(\mem[0][12] ), .A2(n659), .ZN(n646) );
  OAI21_X1 U140 ( .B1(n659), .B2(n380), .A(n645), .ZN(n508) );
  NAND2_X1 U141 ( .A1(\mem[0][13] ), .A2(n659), .ZN(n645) );
  OAI21_X1 U142 ( .B1(n659), .B2(n379), .A(n644), .ZN(n507) );
  NAND2_X1 U143 ( .A1(\mem[0][14] ), .A2(n659), .ZN(n644) );
  INV_X1 U144 ( .A(N10), .ZN(n375) );
  OAI21_X1 U145 ( .B1(n393), .B2(n373), .A(n640), .ZN(n505) );
  NAND2_X1 U146 ( .A1(\mem[1][0] ), .A2(n373), .ZN(n640) );
  OAI21_X1 U147 ( .B1(n392), .B2(n641), .A(n639), .ZN(n504) );
  NAND2_X1 U148 ( .A1(\mem[1][1] ), .A2(n641), .ZN(n639) );
  OAI21_X1 U149 ( .B1(n391), .B2(n373), .A(n638), .ZN(n503) );
  NAND2_X1 U150 ( .A1(\mem[1][2] ), .A2(n641), .ZN(n638) );
  OAI21_X1 U151 ( .B1(n390), .B2(n641), .A(n637), .ZN(n502) );
  NAND2_X1 U152 ( .A1(\mem[1][3] ), .A2(n641), .ZN(n637) );
  OAI21_X1 U153 ( .B1(n389), .B2(n641), .A(n636), .ZN(n501) );
  NAND2_X1 U154 ( .A1(\mem[1][4] ), .A2(n373), .ZN(n636) );
  OAI21_X1 U155 ( .B1(n388), .B2(n641), .A(n635), .ZN(n500) );
  NAND2_X1 U156 ( .A1(\mem[1][5] ), .A2(n373), .ZN(n635) );
  OAI21_X1 U157 ( .B1(n387), .B2(n641), .A(n634), .ZN(n499) );
  NAND2_X1 U158 ( .A1(\mem[1][6] ), .A2(n373), .ZN(n634) );
  OAI21_X1 U159 ( .B1(n378), .B2(n641), .A(n625), .ZN(n490) );
  NAND2_X1 U160 ( .A1(\mem[1][15] ), .A2(n641), .ZN(n625) );
  OAI21_X1 U161 ( .B1(n393), .B2(n624), .A(n623), .ZN(n489) );
  NAND2_X1 U162 ( .A1(\mem[2][0] ), .A2(n372), .ZN(n623) );
  OAI21_X1 U163 ( .B1(n392), .B2(n624), .A(n622), .ZN(n488) );
  NAND2_X1 U164 ( .A1(\mem[2][1] ), .A2(n372), .ZN(n622) );
  OAI21_X1 U165 ( .B1(n391), .B2(n624), .A(n621), .ZN(n487) );
  NAND2_X1 U166 ( .A1(\mem[2][2] ), .A2(n372), .ZN(n621) );
  OAI21_X1 U167 ( .B1(n390), .B2(n624), .A(n620), .ZN(n486) );
  NAND2_X1 U168 ( .A1(\mem[2][3] ), .A2(n372), .ZN(n620) );
  OAI21_X1 U169 ( .B1(n389), .B2(n624), .A(n619), .ZN(n485) );
  NAND2_X1 U170 ( .A1(\mem[2][4] ), .A2(n624), .ZN(n619) );
  OAI21_X1 U171 ( .B1(n388), .B2(n624), .A(n618), .ZN(n484) );
  NAND2_X1 U172 ( .A1(\mem[2][5] ), .A2(n624), .ZN(n618) );
  OAI21_X1 U173 ( .B1(n387), .B2(n624), .A(n617), .ZN(n483) );
  NAND2_X1 U174 ( .A1(\mem[2][6] ), .A2(n624), .ZN(n617) );
  OAI21_X1 U175 ( .B1(n378), .B2(n624), .A(n608), .ZN(n474) );
  NAND2_X1 U176 ( .A1(\mem[2][15] ), .A2(n372), .ZN(n608) );
  OAI21_X1 U177 ( .B1(n393), .B2(n607), .A(n606), .ZN(n473) );
  NAND2_X1 U178 ( .A1(\mem[3][0] ), .A2(n371), .ZN(n606) );
  OAI21_X1 U179 ( .B1(n392), .B2(n607), .A(n605), .ZN(n472) );
  NAND2_X1 U180 ( .A1(\mem[3][1] ), .A2(n371), .ZN(n605) );
  OAI21_X1 U181 ( .B1(n391), .B2(n607), .A(n604), .ZN(n471) );
  NAND2_X1 U182 ( .A1(\mem[3][2] ), .A2(n371), .ZN(n604) );
  OAI21_X1 U183 ( .B1(n390), .B2(n607), .A(n603), .ZN(n470) );
  NAND2_X1 U184 ( .A1(\mem[3][3] ), .A2(n371), .ZN(n603) );
  OAI21_X1 U185 ( .B1(n389), .B2(n607), .A(n602), .ZN(n469) );
  NAND2_X1 U186 ( .A1(\mem[3][4] ), .A2(n607), .ZN(n602) );
  OAI21_X1 U187 ( .B1(n388), .B2(n607), .A(n601), .ZN(n468) );
  NAND2_X1 U188 ( .A1(\mem[3][5] ), .A2(n607), .ZN(n601) );
  OAI21_X1 U189 ( .B1(n387), .B2(n607), .A(n600), .ZN(n467) );
  NAND2_X1 U190 ( .A1(\mem[3][6] ), .A2(n607), .ZN(n600) );
  OAI21_X1 U191 ( .B1(n378), .B2(n607), .A(n591), .ZN(n458) );
  NAND2_X1 U192 ( .A1(\mem[3][15] ), .A2(n371), .ZN(n591) );
  OAI21_X1 U193 ( .B1(n393), .B2(n590), .A(n589), .ZN(n457) );
  NAND2_X1 U194 ( .A1(\mem[4][0] ), .A2(n370), .ZN(n589) );
  OAI21_X1 U195 ( .B1(n392), .B2(n590), .A(n588), .ZN(n456) );
  NAND2_X1 U196 ( .A1(\mem[4][1] ), .A2(n370), .ZN(n588) );
  OAI21_X1 U197 ( .B1(n391), .B2(n590), .A(n587), .ZN(n455) );
  NAND2_X1 U198 ( .A1(\mem[4][2] ), .A2(n370), .ZN(n587) );
  OAI21_X1 U199 ( .B1(n390), .B2(n590), .A(n586), .ZN(n454) );
  NAND2_X1 U200 ( .A1(\mem[4][3] ), .A2(n370), .ZN(n586) );
  OAI21_X1 U201 ( .B1(n389), .B2(n590), .A(n585), .ZN(n453) );
  NAND2_X1 U202 ( .A1(\mem[4][4] ), .A2(n590), .ZN(n585) );
  OAI21_X1 U203 ( .B1(n388), .B2(n590), .A(n584), .ZN(n452) );
  NAND2_X1 U204 ( .A1(\mem[4][5] ), .A2(n590), .ZN(n584) );
  OAI21_X1 U205 ( .B1(n387), .B2(n590), .A(n583), .ZN(n451) );
  NAND2_X1 U206 ( .A1(\mem[4][6] ), .A2(n590), .ZN(n583) );
  OAI21_X1 U207 ( .B1(n378), .B2(n590), .A(n574), .ZN(n442) );
  NAND2_X1 U208 ( .A1(\mem[4][15] ), .A2(n370), .ZN(n574) );
  OAI21_X1 U209 ( .B1(n393), .B2(n369), .A(n571), .ZN(n441) );
  NAND2_X1 U210 ( .A1(\mem[5][0] ), .A2(n369), .ZN(n571) );
  OAI21_X1 U211 ( .B1(n392), .B2(n369), .A(n570), .ZN(n440) );
  NAND2_X1 U212 ( .A1(\mem[5][1] ), .A2(n572), .ZN(n570) );
  OAI21_X1 U213 ( .B1(n391), .B2(n369), .A(n569), .ZN(n439) );
  NAND2_X1 U214 ( .A1(\mem[5][2] ), .A2(n572), .ZN(n569) );
  OAI21_X1 U215 ( .B1(n390), .B2(n369), .A(n568), .ZN(n438) );
  NAND2_X1 U216 ( .A1(\mem[5][3] ), .A2(n572), .ZN(n568) );
  OAI21_X1 U217 ( .B1(n389), .B2(n369), .A(n567), .ZN(n437) );
  NAND2_X1 U218 ( .A1(\mem[5][4] ), .A2(n369), .ZN(n567) );
  OAI21_X1 U219 ( .B1(n388), .B2(n369), .A(n566), .ZN(n436) );
  NAND2_X1 U220 ( .A1(\mem[5][5] ), .A2(n369), .ZN(n566) );
  OAI21_X1 U221 ( .B1(n387), .B2(n369), .A(n565), .ZN(n435) );
  NAND2_X1 U222 ( .A1(\mem[5][6] ), .A2(n369), .ZN(n565) );
  OAI21_X1 U223 ( .B1(n378), .B2(n369), .A(n556), .ZN(n426) );
  NAND2_X1 U224 ( .A1(\mem[5][15] ), .A2(n369), .ZN(n556) );
  OAI21_X1 U225 ( .B1(n393), .B2(n555), .A(n554), .ZN(n425) );
  NAND2_X1 U226 ( .A1(\mem[6][0] ), .A2(n368), .ZN(n554) );
  OAI21_X1 U227 ( .B1(n392), .B2(n555), .A(n553), .ZN(n424) );
  NAND2_X1 U228 ( .A1(\mem[6][1] ), .A2(n368), .ZN(n553) );
  OAI21_X1 U229 ( .B1(n391), .B2(n555), .A(n552), .ZN(n423) );
  NAND2_X1 U230 ( .A1(\mem[6][2] ), .A2(n368), .ZN(n552) );
  OAI21_X1 U231 ( .B1(n390), .B2(n555), .A(n551), .ZN(n422) );
  NAND2_X1 U232 ( .A1(\mem[6][3] ), .A2(n368), .ZN(n551) );
  OAI21_X1 U233 ( .B1(n389), .B2(n555), .A(n550), .ZN(n421) );
  NAND2_X1 U234 ( .A1(\mem[6][4] ), .A2(n555), .ZN(n550) );
  OAI21_X1 U235 ( .B1(n388), .B2(n555), .A(n549), .ZN(n420) );
  NAND2_X1 U236 ( .A1(\mem[6][5] ), .A2(n555), .ZN(n549) );
  OAI21_X1 U237 ( .B1(n387), .B2(n555), .A(n548), .ZN(n419) );
  NAND2_X1 U238 ( .A1(\mem[6][6] ), .A2(n555), .ZN(n548) );
  OAI21_X1 U239 ( .B1(n378), .B2(n555), .A(n539), .ZN(n410) );
  NAND2_X1 U240 ( .A1(\mem[6][15] ), .A2(n368), .ZN(n539) );
  OAI21_X1 U241 ( .B1(n393), .B2(n538), .A(n537), .ZN(n409) );
  NAND2_X1 U242 ( .A1(\mem[7][0] ), .A2(n367), .ZN(n537) );
  OAI21_X1 U243 ( .B1(n392), .B2(n538), .A(n536), .ZN(n408) );
  NAND2_X1 U244 ( .A1(\mem[7][1] ), .A2(n367), .ZN(n536) );
  OAI21_X1 U245 ( .B1(n391), .B2(n538), .A(n535), .ZN(n407) );
  NAND2_X1 U246 ( .A1(\mem[7][2] ), .A2(n367), .ZN(n535) );
  OAI21_X1 U247 ( .B1(n390), .B2(n538), .A(n534), .ZN(n406) );
  NAND2_X1 U248 ( .A1(\mem[7][3] ), .A2(n367), .ZN(n534) );
  OAI21_X1 U249 ( .B1(n389), .B2(n538), .A(n533), .ZN(n405) );
  NAND2_X1 U250 ( .A1(\mem[7][4] ), .A2(n538), .ZN(n533) );
  OAI21_X1 U251 ( .B1(n388), .B2(n538), .A(n532), .ZN(n404) );
  NAND2_X1 U252 ( .A1(\mem[7][5] ), .A2(n538), .ZN(n532) );
  OAI21_X1 U253 ( .B1(n387), .B2(n538), .A(n531), .ZN(n403) );
  NAND2_X1 U254 ( .A1(\mem[7][6] ), .A2(n538), .ZN(n531) );
  OAI21_X1 U255 ( .B1(n378), .B2(n538), .A(n522), .ZN(n394) );
  NAND2_X1 U256 ( .A1(\mem[7][15] ), .A2(n367), .ZN(n522) );
  OAI21_X1 U257 ( .B1(n374), .B2(n393), .A(n658), .ZN(n521) );
  NAND2_X1 U258 ( .A1(\mem[0][0] ), .A2(n659), .ZN(n658) );
  OAI21_X1 U259 ( .B1(n374), .B2(n392), .A(n657), .ZN(n520) );
  NAND2_X1 U260 ( .A1(\mem[0][1] ), .A2(n659), .ZN(n657) );
  OAI21_X1 U261 ( .B1(n374), .B2(n391), .A(n656), .ZN(n519) );
  NAND2_X1 U262 ( .A1(\mem[0][2] ), .A2(n659), .ZN(n656) );
  OAI21_X1 U263 ( .B1(n374), .B2(n390), .A(n655), .ZN(n518) );
  NAND2_X1 U264 ( .A1(\mem[0][3] ), .A2(n659), .ZN(n655) );
  OAI21_X1 U265 ( .B1(n374), .B2(n389), .A(n654), .ZN(n517) );
  NAND2_X1 U266 ( .A1(\mem[0][4] ), .A2(n374), .ZN(n654) );
  OAI21_X1 U267 ( .B1(n374), .B2(n388), .A(n653), .ZN(n516) );
  NAND2_X1 U268 ( .A1(\mem[0][5] ), .A2(n374), .ZN(n653) );
  OAI21_X1 U269 ( .B1(n374), .B2(n387), .A(n652), .ZN(n515) );
  NAND2_X1 U270 ( .A1(\mem[0][6] ), .A2(n374), .ZN(n652) );
  OAI21_X1 U271 ( .B1(n374), .B2(n386), .A(n651), .ZN(n514) );
  NAND2_X1 U272 ( .A1(\mem[0][7] ), .A2(n374), .ZN(n651) );
  OAI21_X1 U273 ( .B1(n374), .B2(n378), .A(n643), .ZN(n506) );
  NAND2_X1 U274 ( .A1(\mem[0][15] ), .A2(n659), .ZN(n643) );
  INV_X1 U275 ( .A(N11), .ZN(n376) );
  INV_X1 U276 ( .A(data_in[0]), .ZN(n393) );
  INV_X1 U277 ( .A(data_in[1]), .ZN(n392) );
  INV_X1 U278 ( .A(data_in[2]), .ZN(n391) );
  INV_X1 U279 ( .A(data_in[3]), .ZN(n390) );
  INV_X1 U288 ( .A(data_in[4]), .ZN(n389) );
  INV_X1 U289 ( .A(data_in[5]), .ZN(n388) );
  INV_X1 U290 ( .A(data_in[6]), .ZN(n387) );
  INV_X1 U291 ( .A(data_in[7]), .ZN(n386) );
  INV_X1 U292 ( .A(data_in[8]), .ZN(n385) );
  INV_X1 U293 ( .A(data_in[9]), .ZN(n384) );
  INV_X1 U294 ( .A(data_in[10]), .ZN(n383) );
  INV_X1 U295 ( .A(data_in[11]), .ZN(n382) );
  INV_X1 U296 ( .A(data_in[12]), .ZN(n381) );
  INV_X1 U297 ( .A(data_in[13]), .ZN(n380) );
  INV_X1 U298 ( .A(data_in[14]), .ZN(n379) );
  INV_X1 U299 ( .A(data_in[15]), .ZN(n378) );
  MUX2_X1 U300 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n365), .Z(n1) );
  MUX2_X1 U301 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n364), .Z(n2) );
  MUX2_X1 U302 ( .A(n2), .B(n1), .S(n363), .Z(n3) );
  MUX2_X1 U303 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n366), .Z(n4) );
  MUX2_X1 U304 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n365), .Z(n5) );
  MUX2_X1 U305 ( .A(n5), .B(n4), .S(n363), .Z(n6) );
  MUX2_X1 U306 ( .A(n6), .B(n3), .S(N12), .Z(N28) );
  MUX2_X1 U307 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n364), .Z(n7) );
  MUX2_X1 U308 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n364), .Z(n8) );
  MUX2_X1 U309 ( .A(n8), .B(n7), .S(n363), .Z(n9) );
  MUX2_X1 U310 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n364), .Z(n10) );
  MUX2_X1 U311 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n364), .Z(n11) );
  MUX2_X1 U312 ( .A(n11), .B(n10), .S(N11), .Z(n12) );
  MUX2_X1 U313 ( .A(n12), .B(n9), .S(N12), .Z(N27) );
  MUX2_X1 U314 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n364), .Z(n13) );
  MUX2_X1 U315 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n364), .Z(n14) );
  MUX2_X1 U316 ( .A(n14), .B(n13), .S(n363), .Z(n15) );
  MUX2_X1 U317 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n364), .Z(n16) );
  MUX2_X1 U318 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n364), .Z(n17) );
  MUX2_X1 U319 ( .A(n17), .B(n16), .S(n363), .Z(n18) );
  MUX2_X1 U320 ( .A(n18), .B(n15), .S(N12), .Z(N26) );
  MUX2_X1 U321 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n364), .Z(n19) );
  MUX2_X1 U322 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n364), .Z(n286) );
  MUX2_X1 U323 ( .A(n286), .B(n19), .S(n363), .Z(n287) );
  MUX2_X1 U324 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n364), .Z(n288) );
  MUX2_X1 U325 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n364), .Z(n289) );
  MUX2_X1 U326 ( .A(n289), .B(n288), .S(N11), .Z(n290) );
  MUX2_X1 U327 ( .A(n290), .B(n287), .S(N12), .Z(N25) );
  MUX2_X1 U328 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n365), .Z(n291) );
  MUX2_X1 U329 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n366), .Z(n292) );
  MUX2_X1 U330 ( .A(n292), .B(n291), .S(n363), .Z(n293) );
  MUX2_X1 U331 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n364), .Z(n294) );
  MUX2_X1 U332 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n365), .Z(n295) );
  MUX2_X1 U333 ( .A(n295), .B(n294), .S(n363), .Z(n296) );
  MUX2_X1 U334 ( .A(n296), .B(n293), .S(N12), .Z(N24) );
  MUX2_X1 U335 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n366), .Z(n297) );
  MUX2_X1 U336 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n364), .Z(n298) );
  MUX2_X1 U337 ( .A(n298), .B(n297), .S(n363), .Z(n299) );
  MUX2_X1 U338 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n366), .Z(n300) );
  MUX2_X1 U339 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n364), .Z(n301) );
  MUX2_X1 U340 ( .A(n301), .B(n300), .S(n363), .Z(n302) );
  MUX2_X1 U341 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n366), .Z(n303) );
  MUX2_X1 U342 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n364), .Z(n304) );
  MUX2_X1 U343 ( .A(n304), .B(n303), .S(n363), .Z(n305) );
  MUX2_X1 U344 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n365), .Z(n306) );
  MUX2_X1 U345 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n366), .Z(n307) );
  MUX2_X1 U346 ( .A(n307), .B(n306), .S(n363), .Z(n308) );
  MUX2_X1 U347 ( .A(n308), .B(n305), .S(N12), .Z(N22) );
  MUX2_X1 U348 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n365), .Z(n309) );
  MUX2_X1 U349 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n364), .Z(n310) );
  MUX2_X1 U350 ( .A(n310), .B(n309), .S(n363), .Z(n311) );
  MUX2_X1 U351 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n365), .Z(n312) );
  MUX2_X1 U352 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n364), .Z(n313) );
  MUX2_X1 U353 ( .A(n313), .B(n312), .S(n363), .Z(n314) );
  MUX2_X1 U354 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n365), .Z(n315) );
  MUX2_X1 U355 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n364), .Z(n316) );
  MUX2_X1 U356 ( .A(n316), .B(n315), .S(n363), .Z(n317) );
  MUX2_X1 U357 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n366), .Z(n318) );
  MUX2_X1 U358 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n364), .Z(n319) );
  MUX2_X1 U359 ( .A(n319), .B(n318), .S(n363), .Z(n320) );
  MUX2_X1 U360 ( .A(n320), .B(n317), .S(N12), .Z(N20) );
  MUX2_X1 U361 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n366), .Z(n321) );
  MUX2_X1 U362 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n365), .Z(n322) );
  MUX2_X1 U363 ( .A(n322), .B(n321), .S(n363), .Z(n323) );
  MUX2_X1 U364 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n366), .Z(n324) );
  MUX2_X1 U365 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(N10), .Z(n325) );
  MUX2_X1 U366 ( .A(n325), .B(n324), .S(n363), .Z(n326) );
  MUX2_X1 U367 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n365), .Z(n327) );
  MUX2_X1 U368 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n365), .Z(n328) );
  MUX2_X1 U369 ( .A(n328), .B(n327), .S(n363), .Z(n329) );
  MUX2_X1 U370 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n365), .Z(n330) );
  MUX2_X1 U371 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n365), .Z(n331) );
  MUX2_X1 U372 ( .A(n331), .B(n330), .S(n363), .Z(n332) );
  MUX2_X1 U373 ( .A(n332), .B(n329), .S(N12), .Z(N18) );
  MUX2_X1 U374 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n365), .Z(n333) );
  MUX2_X1 U375 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n365), .Z(n334) );
  MUX2_X1 U376 ( .A(n334), .B(n333), .S(N11), .Z(n335) );
  MUX2_X1 U377 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n365), .Z(n336) );
  MUX2_X1 U378 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n365), .Z(n337) );
  MUX2_X1 U379 ( .A(n337), .B(n336), .S(N11), .Z(n338) );
  MUX2_X1 U380 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n365), .Z(n339) );
  MUX2_X1 U381 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n365), .Z(n340) );
  MUX2_X1 U382 ( .A(n340), .B(n339), .S(n363), .Z(n341) );
  MUX2_X1 U383 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n365), .Z(n342) );
  MUX2_X1 U384 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n365), .Z(n343) );
  MUX2_X1 U385 ( .A(n343), .B(n342), .S(N11), .Z(n344) );
  MUX2_X1 U386 ( .A(n344), .B(n341), .S(N12), .Z(N16) );
  MUX2_X1 U387 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n366), .Z(n345) );
  MUX2_X1 U388 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n366), .Z(n346) );
  MUX2_X1 U389 ( .A(n346), .B(n345), .S(N11), .Z(n347) );
  MUX2_X1 U390 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n366), .Z(n348) );
  MUX2_X1 U391 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n366), .Z(n349) );
  MUX2_X1 U392 ( .A(n349), .B(n348), .S(N11), .Z(n350) );
  MUX2_X1 U393 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n366), .Z(n351) );
  MUX2_X1 U394 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n366), .Z(n352) );
  MUX2_X1 U395 ( .A(n352), .B(n351), .S(n363), .Z(n353) );
  MUX2_X1 U396 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n366), .Z(n354) );
  MUX2_X1 U397 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n366), .Z(n355) );
  MUX2_X1 U398 ( .A(n355), .B(n354), .S(N11), .Z(n356) );
  MUX2_X1 U399 ( .A(n356), .B(n353), .S(N12), .Z(N14) );
  MUX2_X1 U400 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n366), .Z(n357) );
  MUX2_X1 U401 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n366), .Z(n358) );
  MUX2_X1 U402 ( .A(n358), .B(n357), .S(n363), .Z(n359) );
  MUX2_X1 U403 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n366), .Z(n360) );
  MUX2_X1 U404 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n366), .Z(n361) );
  MUX2_X1 U405 ( .A(n361), .B(n360), .S(N11), .Z(n362) );
  MUX2_X1 U406 ( .A(n362), .B(n359), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH16_SIZE8_LOGSIZE3_7 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] ,
         \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][15] , \mem[6][14] , \mem[6][13] ,
         \mem[6][12] , \mem[6][11] , \mem[6][10] , \mem[6][9] , \mem[6][8] ,
         \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] ,
         \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[5][15] , \mem[5][14] ,
         \mem[5][13] , \mem[5][12] , \mem[5][11] , \mem[5][10] , \mem[5][9] ,
         \mem[5][8] , \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] ,
         \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][15] ,
         \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] , \mem[4][10] ,
         \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N13, N14, N16,
         N18, N20, N21, N22, N24, N26, N28, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[15]  ( .D(N13), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N14), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N16), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N18), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[8]  ( .D(N20), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N22), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N24), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N26), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N28), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][15]  ( .D(n394), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n395), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n396), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n397), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n398), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n399), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n400), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n401), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n402), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n403), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n404), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n405), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n406), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n407), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n408), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n409), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n410), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n411), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n412), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n413), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n414), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n415), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n416), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n417), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n418), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n419), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n420), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n421), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n422), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n423), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n424), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n425), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n426), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n427), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n428), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n429), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n430), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n431), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n432), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n433), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n434), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n435), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n436), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n437), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n438), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n439), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n440), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n441), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n442), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n443), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n444), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n445), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n446), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n447), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n448), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n449), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n450), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n451), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n452), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n453), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n454), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n455), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n456), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n457), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n458), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n459), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n460), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n461), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n462), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n463), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n464), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n465), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n466), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n467), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n468), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n469), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n470), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n471), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n472), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n473), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n474), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n475), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n476), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n477), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n478), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n479), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n480), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n481), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n482), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n483), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n484), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n485), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n486), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n487), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n488), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n489), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n490), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n491), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n492), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n493), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n494), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n495), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n496), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n497), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n498), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n499), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n500), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n501), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n502), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n503), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n504), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n505), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n506), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n507), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n508), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n509), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n510), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n511), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n512), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n513), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n514), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n515), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n516), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n517), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n518), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n519), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n520), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n521), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U280 ( .A1(n375), .A2(n376), .A3(n642), .ZN(n659) );
  NAND3_X1 U281 ( .A1(n642), .A2(n376), .A3(N10), .ZN(n641) );
  NAND3_X1 U282 ( .A1(n642), .A2(n375), .A3(N11), .ZN(n624) );
  NAND3_X1 U283 ( .A1(N10), .A2(n642), .A3(N11), .ZN(n607) );
  NAND3_X1 U284 ( .A1(n375), .A2(n376), .A3(n573), .ZN(n590) );
  NAND3_X1 U285 ( .A1(N10), .A2(n376), .A3(n573), .ZN(n572) );
  NAND3_X1 U286 ( .A1(N11), .A2(n375), .A3(n573), .ZN(n555) );
  NAND3_X1 U287 ( .A1(N11), .A2(N10), .A3(n573), .ZN(n538) );
  DFF_X1 \data_out_reg[7]  ( .D(N21), .CK(clk), .Q(data_out[7]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n12), .SI(n9), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n326), .SI(n323), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n302), .SI(n299), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n338), .SI(n335), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n290), .SI(n287), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n350), .SI(n347), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  BUF_X1 U3 ( .A(n624), .Z(n372) );
  BUF_X1 U4 ( .A(n607), .Z(n371) );
  BUF_X1 U5 ( .A(n590), .Z(n370) );
  BUF_X1 U6 ( .A(n572), .Z(n369) );
  BUF_X1 U7 ( .A(n538), .Z(n367) );
  BUF_X1 U8 ( .A(n555), .Z(n368) );
  BUF_X1 U9 ( .A(n641), .Z(n373) );
  BUF_X1 U10 ( .A(N10), .Z(n364) );
  BUF_X1 U11 ( .A(N10), .Z(n365) );
  BUF_X1 U12 ( .A(N10), .Z(n366) );
  BUF_X1 U13 ( .A(n659), .Z(n374) );
  BUF_X1 U14 ( .A(N11), .Z(n363) );
  AND2_X1 U15 ( .A1(N12), .A2(wr_en), .ZN(n573) );
  OAI21_X1 U16 ( .B1(n386), .B2(n607), .A(n599), .ZN(n466) );
  NAND2_X1 U17 ( .A1(\mem[3][7] ), .A2(n371), .ZN(n599) );
  OAI21_X1 U18 ( .B1(n385), .B2(n371), .A(n598), .ZN(n465) );
  NAND2_X1 U19 ( .A1(\mem[3][8] ), .A2(n371), .ZN(n598) );
  OAI21_X1 U20 ( .B1(n384), .B2(n607), .A(n597), .ZN(n464) );
  NAND2_X1 U21 ( .A1(\mem[3][9] ), .A2(n371), .ZN(n597) );
  OAI21_X1 U22 ( .B1(n383), .B2(n607), .A(n596), .ZN(n463) );
  NAND2_X1 U23 ( .A1(\mem[3][10] ), .A2(n371), .ZN(n596) );
  OAI21_X1 U24 ( .B1(n382), .B2(n607), .A(n595), .ZN(n462) );
  NAND2_X1 U25 ( .A1(\mem[3][11] ), .A2(n371), .ZN(n595) );
  OAI21_X1 U26 ( .B1(n381), .B2(n607), .A(n594), .ZN(n461) );
  NAND2_X1 U27 ( .A1(\mem[3][12] ), .A2(n371), .ZN(n594) );
  OAI21_X1 U28 ( .B1(n380), .B2(n607), .A(n593), .ZN(n460) );
  NAND2_X1 U29 ( .A1(\mem[3][13] ), .A2(n371), .ZN(n593) );
  OAI21_X1 U30 ( .B1(n379), .B2(n607), .A(n592), .ZN(n459) );
  NAND2_X1 U31 ( .A1(\mem[3][14] ), .A2(n371), .ZN(n592) );
  OAI21_X1 U32 ( .B1(n386), .B2(n572), .A(n564), .ZN(n434) );
  NAND2_X1 U33 ( .A1(\mem[5][7] ), .A2(n369), .ZN(n564) );
  OAI21_X1 U34 ( .B1(n385), .B2(n369), .A(n563), .ZN(n433) );
  NAND2_X1 U35 ( .A1(\mem[5][8] ), .A2(n369), .ZN(n563) );
  OAI21_X1 U36 ( .B1(n384), .B2(n572), .A(n562), .ZN(n432) );
  NAND2_X1 U37 ( .A1(\mem[5][9] ), .A2(n369), .ZN(n562) );
  OAI21_X1 U38 ( .B1(n383), .B2(n572), .A(n561), .ZN(n431) );
  NAND2_X1 U39 ( .A1(\mem[5][10] ), .A2(n369), .ZN(n561) );
  OAI21_X1 U40 ( .B1(n382), .B2(n572), .A(n560), .ZN(n430) );
  NAND2_X1 U41 ( .A1(\mem[5][11] ), .A2(n369), .ZN(n560) );
  OAI21_X1 U42 ( .B1(n381), .B2(n572), .A(n559), .ZN(n429) );
  NAND2_X1 U43 ( .A1(\mem[5][12] ), .A2(n369), .ZN(n559) );
  OAI21_X1 U44 ( .B1(n380), .B2(n572), .A(n558), .ZN(n428) );
  NAND2_X1 U45 ( .A1(\mem[5][13] ), .A2(n369), .ZN(n558) );
  OAI21_X1 U46 ( .B1(n379), .B2(n572), .A(n557), .ZN(n427) );
  NAND2_X1 U47 ( .A1(\mem[5][14] ), .A2(n369), .ZN(n557) );
  OAI21_X1 U48 ( .B1(n386), .B2(n538), .A(n530), .ZN(n402) );
  NAND2_X1 U49 ( .A1(\mem[7][7] ), .A2(n367), .ZN(n530) );
  OAI21_X1 U50 ( .B1(n385), .B2(n367), .A(n529), .ZN(n401) );
  NAND2_X1 U51 ( .A1(\mem[7][8] ), .A2(n367), .ZN(n529) );
  OAI21_X1 U52 ( .B1(n384), .B2(n538), .A(n528), .ZN(n400) );
  NAND2_X1 U53 ( .A1(\mem[7][9] ), .A2(n367), .ZN(n528) );
  OAI21_X1 U54 ( .B1(n383), .B2(n538), .A(n527), .ZN(n399) );
  NAND2_X1 U55 ( .A1(\mem[7][10] ), .A2(n367), .ZN(n527) );
  OAI21_X1 U56 ( .B1(n382), .B2(n538), .A(n526), .ZN(n398) );
  NAND2_X1 U57 ( .A1(\mem[7][11] ), .A2(n367), .ZN(n526) );
  OAI21_X1 U58 ( .B1(n381), .B2(n538), .A(n525), .ZN(n397) );
  NAND2_X1 U59 ( .A1(\mem[7][12] ), .A2(n367), .ZN(n525) );
  OAI21_X1 U60 ( .B1(n380), .B2(n538), .A(n524), .ZN(n396) );
  NAND2_X1 U61 ( .A1(\mem[7][13] ), .A2(n367), .ZN(n524) );
  OAI21_X1 U62 ( .B1(n379), .B2(n538), .A(n523), .ZN(n395) );
  NAND2_X1 U63 ( .A1(\mem[7][14] ), .A2(n367), .ZN(n523) );
  OAI21_X1 U64 ( .B1(n386), .B2(n373), .A(n633), .ZN(n498) );
  NAND2_X1 U65 ( .A1(\mem[1][7] ), .A2(n373), .ZN(n633) );
  OAI21_X1 U66 ( .B1(n385), .B2(n373), .A(n632), .ZN(n497) );
  NAND2_X1 U67 ( .A1(\mem[1][8] ), .A2(n641), .ZN(n632) );
  OAI21_X1 U68 ( .B1(n384), .B2(n373), .A(n631), .ZN(n496) );
  NAND2_X1 U69 ( .A1(\mem[1][9] ), .A2(n641), .ZN(n631) );
  OAI21_X1 U70 ( .B1(n383), .B2(n373), .A(n630), .ZN(n495) );
  NAND2_X1 U71 ( .A1(\mem[1][10] ), .A2(n641), .ZN(n630) );
  OAI21_X1 U72 ( .B1(n382), .B2(n373), .A(n629), .ZN(n494) );
  NAND2_X1 U73 ( .A1(\mem[1][11] ), .A2(n641), .ZN(n629) );
  OAI21_X1 U74 ( .B1(n381), .B2(n373), .A(n628), .ZN(n493) );
  NAND2_X1 U75 ( .A1(\mem[1][12] ), .A2(n641), .ZN(n628) );
  OAI21_X1 U76 ( .B1(n380), .B2(n373), .A(n627), .ZN(n492) );
  NAND2_X1 U77 ( .A1(\mem[1][13] ), .A2(n641), .ZN(n627) );
  OAI21_X1 U78 ( .B1(n379), .B2(n373), .A(n626), .ZN(n491) );
  NAND2_X1 U79 ( .A1(\mem[1][14] ), .A2(n641), .ZN(n626) );
  OAI21_X1 U80 ( .B1(n386), .B2(n555), .A(n547), .ZN(n418) );
  NAND2_X1 U81 ( .A1(\mem[6][7] ), .A2(n368), .ZN(n547) );
  OAI21_X1 U82 ( .B1(n385), .B2(n555), .A(n546), .ZN(n417) );
  NAND2_X1 U83 ( .A1(\mem[6][8] ), .A2(n555), .ZN(n546) );
  OAI21_X1 U84 ( .B1(n384), .B2(n555), .A(n545), .ZN(n416) );
  NAND2_X1 U85 ( .A1(\mem[6][9] ), .A2(n555), .ZN(n545) );
  OAI21_X1 U86 ( .B1(n383), .B2(n555), .A(n544), .ZN(n415) );
  NAND2_X1 U87 ( .A1(\mem[6][10] ), .A2(n555), .ZN(n544) );
  OAI21_X1 U88 ( .B1(n382), .B2(n555), .A(n543), .ZN(n414) );
  NAND2_X1 U89 ( .A1(\mem[6][11] ), .A2(n555), .ZN(n543) );
  OAI21_X1 U90 ( .B1(n381), .B2(n555), .A(n542), .ZN(n413) );
  NAND2_X1 U91 ( .A1(\mem[6][12] ), .A2(n555), .ZN(n542) );
  OAI21_X1 U92 ( .B1(n380), .B2(n555), .A(n541), .ZN(n412) );
  NAND2_X1 U93 ( .A1(\mem[6][13] ), .A2(n555), .ZN(n541) );
  OAI21_X1 U94 ( .B1(n379), .B2(n555), .A(n540), .ZN(n411) );
  NAND2_X1 U95 ( .A1(\mem[6][14] ), .A2(n555), .ZN(n540) );
  OAI21_X1 U96 ( .B1(n386), .B2(n624), .A(n616), .ZN(n482) );
  NAND2_X1 U97 ( .A1(\mem[2][7] ), .A2(n372), .ZN(n616) );
  OAI21_X1 U98 ( .B1(n385), .B2(n372), .A(n615), .ZN(n481) );
  NAND2_X1 U99 ( .A1(\mem[2][8] ), .A2(n372), .ZN(n615) );
  OAI21_X1 U100 ( .B1(n384), .B2(n624), .A(n614), .ZN(n480) );
  NAND2_X1 U101 ( .A1(\mem[2][9] ), .A2(n372), .ZN(n614) );
  OAI21_X1 U102 ( .B1(n383), .B2(n624), .A(n613), .ZN(n479) );
  NAND2_X1 U103 ( .A1(\mem[2][10] ), .A2(n372), .ZN(n613) );
  OAI21_X1 U104 ( .B1(n382), .B2(n624), .A(n612), .ZN(n478) );
  NAND2_X1 U105 ( .A1(\mem[2][11] ), .A2(n372), .ZN(n612) );
  OAI21_X1 U106 ( .B1(n381), .B2(n624), .A(n611), .ZN(n477) );
  NAND2_X1 U107 ( .A1(\mem[2][12] ), .A2(n372), .ZN(n611) );
  OAI21_X1 U108 ( .B1(n380), .B2(n624), .A(n610), .ZN(n476) );
  NAND2_X1 U109 ( .A1(\mem[2][13] ), .A2(n372), .ZN(n610) );
  OAI21_X1 U110 ( .B1(n379), .B2(n624), .A(n609), .ZN(n475) );
  NAND2_X1 U111 ( .A1(\mem[2][14] ), .A2(n372), .ZN(n609) );
  OAI21_X1 U112 ( .B1(n386), .B2(n590), .A(n582), .ZN(n450) );
  NAND2_X1 U113 ( .A1(\mem[4][7] ), .A2(n370), .ZN(n582) );
  OAI21_X1 U114 ( .B1(n385), .B2(n370), .A(n581), .ZN(n449) );
  NAND2_X1 U115 ( .A1(\mem[4][8] ), .A2(n370), .ZN(n581) );
  OAI21_X1 U116 ( .B1(n384), .B2(n590), .A(n580), .ZN(n448) );
  NAND2_X1 U117 ( .A1(\mem[4][9] ), .A2(n370), .ZN(n580) );
  OAI21_X1 U118 ( .B1(n383), .B2(n590), .A(n579), .ZN(n447) );
  NAND2_X1 U119 ( .A1(\mem[4][10] ), .A2(n370), .ZN(n579) );
  OAI21_X1 U120 ( .B1(n382), .B2(n590), .A(n578), .ZN(n446) );
  NAND2_X1 U121 ( .A1(\mem[4][11] ), .A2(n370), .ZN(n578) );
  OAI21_X1 U122 ( .B1(n381), .B2(n590), .A(n577), .ZN(n445) );
  NAND2_X1 U123 ( .A1(\mem[4][12] ), .A2(n370), .ZN(n577) );
  OAI21_X1 U124 ( .B1(n380), .B2(n590), .A(n576), .ZN(n444) );
  NAND2_X1 U125 ( .A1(\mem[4][13] ), .A2(n370), .ZN(n576) );
  OAI21_X1 U126 ( .B1(n379), .B2(n590), .A(n575), .ZN(n443) );
  NAND2_X1 U127 ( .A1(\mem[4][14] ), .A2(n370), .ZN(n575) );
  OAI21_X1 U128 ( .B1(n374), .B2(n385), .A(n650), .ZN(n513) );
  NAND2_X1 U129 ( .A1(\mem[0][8] ), .A2(n374), .ZN(n650) );
  OAI21_X1 U130 ( .B1(n374), .B2(n384), .A(n649), .ZN(n512) );
  NAND2_X1 U131 ( .A1(\mem[0][9] ), .A2(n374), .ZN(n649) );
  OAI21_X1 U132 ( .B1(n374), .B2(n383), .A(n648), .ZN(n511) );
  NAND2_X1 U133 ( .A1(\mem[0][10] ), .A2(n659), .ZN(n648) );
  OAI21_X1 U134 ( .B1(n374), .B2(n382), .A(n647), .ZN(n510) );
  NAND2_X1 U135 ( .A1(\mem[0][11] ), .A2(n374), .ZN(n647) );
  OAI21_X1 U136 ( .B1(n374), .B2(n381), .A(n646), .ZN(n509) );
  NAND2_X1 U137 ( .A1(\mem[0][12] ), .A2(n659), .ZN(n646) );
  OAI21_X1 U138 ( .B1(n374), .B2(n380), .A(n645), .ZN(n508) );
  NAND2_X1 U139 ( .A1(\mem[0][13] ), .A2(n659), .ZN(n645) );
  OAI21_X1 U140 ( .B1(n374), .B2(n379), .A(n644), .ZN(n507) );
  NAND2_X1 U141 ( .A1(\mem[0][14] ), .A2(n659), .ZN(n644) );
  INV_X1 U142 ( .A(N10), .ZN(n375) );
  OAI21_X1 U143 ( .B1(n393), .B2(n373), .A(n640), .ZN(n505) );
  NAND2_X1 U144 ( .A1(\mem[1][0] ), .A2(n373), .ZN(n640) );
  OAI21_X1 U145 ( .B1(n392), .B2(n641), .A(n639), .ZN(n504) );
  NAND2_X1 U146 ( .A1(\mem[1][1] ), .A2(n641), .ZN(n639) );
  OAI21_X1 U147 ( .B1(n391), .B2(n373), .A(n638), .ZN(n503) );
  NAND2_X1 U148 ( .A1(\mem[1][2] ), .A2(n641), .ZN(n638) );
  OAI21_X1 U149 ( .B1(n390), .B2(n641), .A(n637), .ZN(n502) );
  NAND2_X1 U150 ( .A1(\mem[1][3] ), .A2(n641), .ZN(n637) );
  OAI21_X1 U151 ( .B1(n389), .B2(n641), .A(n636), .ZN(n501) );
  NAND2_X1 U152 ( .A1(\mem[1][4] ), .A2(n373), .ZN(n636) );
  OAI21_X1 U153 ( .B1(n388), .B2(n641), .A(n635), .ZN(n500) );
  NAND2_X1 U154 ( .A1(\mem[1][5] ), .A2(n373), .ZN(n635) );
  OAI21_X1 U155 ( .B1(n387), .B2(n641), .A(n634), .ZN(n499) );
  NAND2_X1 U156 ( .A1(\mem[1][6] ), .A2(n373), .ZN(n634) );
  OAI21_X1 U157 ( .B1(n378), .B2(n641), .A(n625), .ZN(n490) );
  NAND2_X1 U158 ( .A1(\mem[1][15] ), .A2(n641), .ZN(n625) );
  OAI21_X1 U159 ( .B1(n393), .B2(n624), .A(n623), .ZN(n489) );
  NAND2_X1 U160 ( .A1(\mem[2][0] ), .A2(n372), .ZN(n623) );
  OAI21_X1 U161 ( .B1(n392), .B2(n624), .A(n622), .ZN(n488) );
  NAND2_X1 U162 ( .A1(\mem[2][1] ), .A2(n372), .ZN(n622) );
  OAI21_X1 U163 ( .B1(n391), .B2(n624), .A(n621), .ZN(n487) );
  NAND2_X1 U164 ( .A1(\mem[2][2] ), .A2(n372), .ZN(n621) );
  OAI21_X1 U165 ( .B1(n390), .B2(n624), .A(n620), .ZN(n486) );
  NAND2_X1 U166 ( .A1(\mem[2][3] ), .A2(n372), .ZN(n620) );
  OAI21_X1 U167 ( .B1(n389), .B2(n624), .A(n619), .ZN(n485) );
  NAND2_X1 U168 ( .A1(\mem[2][4] ), .A2(n624), .ZN(n619) );
  OAI21_X1 U169 ( .B1(n388), .B2(n624), .A(n618), .ZN(n484) );
  NAND2_X1 U170 ( .A1(\mem[2][5] ), .A2(n624), .ZN(n618) );
  OAI21_X1 U171 ( .B1(n387), .B2(n624), .A(n617), .ZN(n483) );
  NAND2_X1 U172 ( .A1(\mem[2][6] ), .A2(n624), .ZN(n617) );
  OAI21_X1 U173 ( .B1(n378), .B2(n624), .A(n608), .ZN(n474) );
  NAND2_X1 U174 ( .A1(\mem[2][15] ), .A2(n372), .ZN(n608) );
  OAI21_X1 U175 ( .B1(n393), .B2(n607), .A(n606), .ZN(n473) );
  NAND2_X1 U176 ( .A1(\mem[3][0] ), .A2(n371), .ZN(n606) );
  OAI21_X1 U177 ( .B1(n392), .B2(n607), .A(n605), .ZN(n472) );
  NAND2_X1 U178 ( .A1(\mem[3][1] ), .A2(n371), .ZN(n605) );
  OAI21_X1 U179 ( .B1(n391), .B2(n607), .A(n604), .ZN(n471) );
  NAND2_X1 U180 ( .A1(\mem[3][2] ), .A2(n371), .ZN(n604) );
  OAI21_X1 U181 ( .B1(n390), .B2(n607), .A(n603), .ZN(n470) );
  NAND2_X1 U182 ( .A1(\mem[3][3] ), .A2(n371), .ZN(n603) );
  OAI21_X1 U183 ( .B1(n389), .B2(n607), .A(n602), .ZN(n469) );
  NAND2_X1 U184 ( .A1(\mem[3][4] ), .A2(n607), .ZN(n602) );
  OAI21_X1 U185 ( .B1(n388), .B2(n607), .A(n601), .ZN(n468) );
  NAND2_X1 U186 ( .A1(\mem[3][5] ), .A2(n607), .ZN(n601) );
  OAI21_X1 U187 ( .B1(n387), .B2(n607), .A(n600), .ZN(n467) );
  NAND2_X1 U188 ( .A1(\mem[3][6] ), .A2(n607), .ZN(n600) );
  OAI21_X1 U189 ( .B1(n378), .B2(n607), .A(n591), .ZN(n458) );
  NAND2_X1 U190 ( .A1(\mem[3][15] ), .A2(n371), .ZN(n591) );
  OAI21_X1 U191 ( .B1(n393), .B2(n590), .A(n589), .ZN(n457) );
  NAND2_X1 U192 ( .A1(\mem[4][0] ), .A2(n370), .ZN(n589) );
  OAI21_X1 U193 ( .B1(n392), .B2(n590), .A(n588), .ZN(n456) );
  NAND2_X1 U194 ( .A1(\mem[4][1] ), .A2(n370), .ZN(n588) );
  OAI21_X1 U195 ( .B1(n391), .B2(n590), .A(n587), .ZN(n455) );
  NAND2_X1 U196 ( .A1(\mem[4][2] ), .A2(n370), .ZN(n587) );
  OAI21_X1 U197 ( .B1(n390), .B2(n590), .A(n586), .ZN(n454) );
  NAND2_X1 U198 ( .A1(\mem[4][3] ), .A2(n370), .ZN(n586) );
  OAI21_X1 U199 ( .B1(n389), .B2(n590), .A(n585), .ZN(n453) );
  NAND2_X1 U200 ( .A1(\mem[4][4] ), .A2(n590), .ZN(n585) );
  OAI21_X1 U201 ( .B1(n388), .B2(n590), .A(n584), .ZN(n452) );
  NAND2_X1 U202 ( .A1(\mem[4][5] ), .A2(n590), .ZN(n584) );
  OAI21_X1 U203 ( .B1(n387), .B2(n590), .A(n583), .ZN(n451) );
  NAND2_X1 U204 ( .A1(\mem[4][6] ), .A2(n590), .ZN(n583) );
  OAI21_X1 U205 ( .B1(n378), .B2(n590), .A(n574), .ZN(n442) );
  NAND2_X1 U206 ( .A1(\mem[4][15] ), .A2(n370), .ZN(n574) );
  OAI21_X1 U207 ( .B1(n393), .B2(n572), .A(n571), .ZN(n441) );
  NAND2_X1 U208 ( .A1(\mem[5][0] ), .A2(n369), .ZN(n571) );
  OAI21_X1 U209 ( .B1(n392), .B2(n572), .A(n570), .ZN(n440) );
  NAND2_X1 U210 ( .A1(\mem[5][1] ), .A2(n369), .ZN(n570) );
  OAI21_X1 U211 ( .B1(n391), .B2(n572), .A(n569), .ZN(n439) );
  NAND2_X1 U212 ( .A1(\mem[5][2] ), .A2(n369), .ZN(n569) );
  OAI21_X1 U213 ( .B1(n390), .B2(n572), .A(n568), .ZN(n438) );
  NAND2_X1 U214 ( .A1(\mem[5][3] ), .A2(n369), .ZN(n568) );
  OAI21_X1 U215 ( .B1(n389), .B2(n572), .A(n567), .ZN(n437) );
  NAND2_X1 U216 ( .A1(\mem[5][4] ), .A2(n572), .ZN(n567) );
  OAI21_X1 U217 ( .B1(n388), .B2(n572), .A(n566), .ZN(n436) );
  NAND2_X1 U218 ( .A1(\mem[5][5] ), .A2(n572), .ZN(n566) );
  OAI21_X1 U219 ( .B1(n387), .B2(n572), .A(n565), .ZN(n435) );
  NAND2_X1 U220 ( .A1(\mem[5][6] ), .A2(n572), .ZN(n565) );
  OAI21_X1 U221 ( .B1(n378), .B2(n572), .A(n556), .ZN(n426) );
  NAND2_X1 U222 ( .A1(\mem[5][15] ), .A2(n369), .ZN(n556) );
  OAI21_X1 U223 ( .B1(n393), .B2(n368), .A(n554), .ZN(n425) );
  NAND2_X1 U224 ( .A1(\mem[6][0] ), .A2(n368), .ZN(n554) );
  OAI21_X1 U225 ( .B1(n392), .B2(n368), .A(n553), .ZN(n424) );
  NAND2_X1 U226 ( .A1(\mem[6][1] ), .A2(n555), .ZN(n553) );
  OAI21_X1 U227 ( .B1(n391), .B2(n368), .A(n552), .ZN(n423) );
  NAND2_X1 U228 ( .A1(\mem[6][2] ), .A2(n555), .ZN(n552) );
  OAI21_X1 U229 ( .B1(n390), .B2(n368), .A(n551), .ZN(n422) );
  NAND2_X1 U230 ( .A1(\mem[6][3] ), .A2(n555), .ZN(n551) );
  OAI21_X1 U231 ( .B1(n389), .B2(n368), .A(n550), .ZN(n421) );
  NAND2_X1 U232 ( .A1(\mem[6][4] ), .A2(n368), .ZN(n550) );
  OAI21_X1 U233 ( .B1(n388), .B2(n368), .A(n549), .ZN(n420) );
  NAND2_X1 U234 ( .A1(\mem[6][5] ), .A2(n368), .ZN(n549) );
  OAI21_X1 U235 ( .B1(n387), .B2(n368), .A(n548), .ZN(n419) );
  NAND2_X1 U236 ( .A1(\mem[6][6] ), .A2(n368), .ZN(n548) );
  OAI21_X1 U237 ( .B1(n378), .B2(n368), .A(n539), .ZN(n410) );
  NAND2_X1 U238 ( .A1(\mem[6][15] ), .A2(n368), .ZN(n539) );
  OAI21_X1 U239 ( .B1(n393), .B2(n538), .A(n537), .ZN(n409) );
  NAND2_X1 U240 ( .A1(\mem[7][0] ), .A2(n367), .ZN(n537) );
  OAI21_X1 U241 ( .B1(n392), .B2(n538), .A(n536), .ZN(n408) );
  NAND2_X1 U242 ( .A1(\mem[7][1] ), .A2(n367), .ZN(n536) );
  OAI21_X1 U243 ( .B1(n391), .B2(n538), .A(n535), .ZN(n407) );
  NAND2_X1 U244 ( .A1(\mem[7][2] ), .A2(n367), .ZN(n535) );
  OAI21_X1 U245 ( .B1(n390), .B2(n538), .A(n534), .ZN(n406) );
  NAND2_X1 U246 ( .A1(\mem[7][3] ), .A2(n367), .ZN(n534) );
  OAI21_X1 U247 ( .B1(n389), .B2(n538), .A(n533), .ZN(n405) );
  NAND2_X1 U248 ( .A1(\mem[7][4] ), .A2(n538), .ZN(n533) );
  OAI21_X1 U249 ( .B1(n388), .B2(n538), .A(n532), .ZN(n404) );
  NAND2_X1 U250 ( .A1(\mem[7][5] ), .A2(n538), .ZN(n532) );
  OAI21_X1 U251 ( .B1(n387), .B2(n538), .A(n531), .ZN(n403) );
  NAND2_X1 U252 ( .A1(\mem[7][6] ), .A2(n538), .ZN(n531) );
  OAI21_X1 U253 ( .B1(n378), .B2(n538), .A(n522), .ZN(n394) );
  NAND2_X1 U254 ( .A1(\mem[7][15] ), .A2(n367), .ZN(n522) );
  OAI21_X1 U255 ( .B1(n659), .B2(n393), .A(n658), .ZN(n521) );
  NAND2_X1 U256 ( .A1(\mem[0][0] ), .A2(n374), .ZN(n658) );
  OAI21_X1 U257 ( .B1(n659), .B2(n392), .A(n657), .ZN(n520) );
  NAND2_X1 U258 ( .A1(\mem[0][1] ), .A2(n374), .ZN(n657) );
  OAI21_X1 U259 ( .B1(n659), .B2(n391), .A(n656), .ZN(n519) );
  NAND2_X1 U260 ( .A1(\mem[0][2] ), .A2(n374), .ZN(n656) );
  OAI21_X1 U261 ( .B1(n659), .B2(n390), .A(n655), .ZN(n518) );
  NAND2_X1 U262 ( .A1(\mem[0][3] ), .A2(n374), .ZN(n655) );
  OAI21_X1 U263 ( .B1(n659), .B2(n389), .A(n654), .ZN(n517) );
  NAND2_X1 U264 ( .A1(\mem[0][4] ), .A2(n374), .ZN(n654) );
  OAI21_X1 U265 ( .B1(n659), .B2(n388), .A(n653), .ZN(n516) );
  NAND2_X1 U266 ( .A1(\mem[0][5] ), .A2(n659), .ZN(n653) );
  OAI21_X1 U267 ( .B1(n659), .B2(n387), .A(n652), .ZN(n515) );
  NAND2_X1 U268 ( .A1(\mem[0][6] ), .A2(n659), .ZN(n652) );
  OAI21_X1 U269 ( .B1(n659), .B2(n386), .A(n651), .ZN(n514) );
  NAND2_X1 U270 ( .A1(\mem[0][7] ), .A2(n659), .ZN(n651) );
  OAI21_X1 U271 ( .B1(n659), .B2(n378), .A(n643), .ZN(n506) );
  NAND2_X1 U272 ( .A1(\mem[0][15] ), .A2(n374), .ZN(n643) );
  NOR2_X1 U273 ( .A1(n377), .A2(N12), .ZN(n642) );
  INV_X1 U274 ( .A(wr_en), .ZN(n377) );
  INV_X1 U275 ( .A(N11), .ZN(n376) );
  INV_X1 U276 ( .A(data_in[0]), .ZN(n393) );
  INV_X1 U277 ( .A(data_in[1]), .ZN(n392) );
  INV_X1 U278 ( .A(data_in[2]), .ZN(n391) );
  INV_X1 U279 ( .A(data_in[3]), .ZN(n390) );
  INV_X1 U288 ( .A(data_in[4]), .ZN(n389) );
  INV_X1 U289 ( .A(data_in[5]), .ZN(n388) );
  INV_X1 U290 ( .A(data_in[6]), .ZN(n387) );
  INV_X1 U291 ( .A(data_in[7]), .ZN(n386) );
  INV_X1 U292 ( .A(data_in[8]), .ZN(n385) );
  INV_X1 U293 ( .A(data_in[9]), .ZN(n384) );
  INV_X1 U294 ( .A(data_in[10]), .ZN(n383) );
  INV_X1 U295 ( .A(data_in[11]), .ZN(n382) );
  INV_X1 U296 ( .A(data_in[12]), .ZN(n381) );
  INV_X1 U297 ( .A(data_in[13]), .ZN(n380) );
  INV_X1 U298 ( .A(data_in[14]), .ZN(n379) );
  INV_X1 U299 ( .A(data_in[15]), .ZN(n378) );
  MUX2_X1 U300 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n366), .Z(n1) );
  MUX2_X1 U301 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n365), .Z(n2) );
  MUX2_X1 U302 ( .A(n2), .B(n1), .S(n363), .Z(n3) );
  MUX2_X1 U303 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n365), .Z(n4) );
  MUX2_X1 U304 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n364), .Z(n5) );
  MUX2_X1 U305 ( .A(n5), .B(n4), .S(n363), .Z(n6) );
  MUX2_X1 U306 ( .A(n6), .B(n3), .S(N12), .Z(N28) );
  MUX2_X1 U307 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n364), .Z(n7) );
  MUX2_X1 U308 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n364), .Z(n8) );
  MUX2_X1 U309 ( .A(n8), .B(n7), .S(n363), .Z(n9) );
  MUX2_X1 U310 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n364), .Z(n10) );
  MUX2_X1 U311 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n364), .Z(n11) );
  MUX2_X1 U312 ( .A(n11), .B(n10), .S(n363), .Z(n12) );
  MUX2_X1 U313 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n364), .Z(n13) );
  MUX2_X1 U314 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n364), .Z(n14) );
  MUX2_X1 U315 ( .A(n14), .B(n13), .S(n363), .Z(n15) );
  MUX2_X1 U316 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n364), .Z(n16) );
  MUX2_X1 U317 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n364), .Z(n17) );
  MUX2_X1 U318 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U319 ( .A(n18), .B(n15), .S(N12), .Z(N26) );
  MUX2_X1 U320 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n364), .Z(n19) );
  MUX2_X1 U321 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n364), .Z(n286) );
  MUX2_X1 U322 ( .A(n286), .B(n19), .S(N11), .Z(n287) );
  MUX2_X1 U323 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n364), .Z(n288) );
  MUX2_X1 U324 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n364), .Z(n289) );
  MUX2_X1 U325 ( .A(n289), .B(n288), .S(N11), .Z(n290) );
  MUX2_X1 U326 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n365), .Z(n291) );
  MUX2_X1 U327 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n365), .Z(n292) );
  MUX2_X1 U328 ( .A(n292), .B(n291), .S(n363), .Z(n293) );
  MUX2_X1 U329 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n365), .Z(n294) );
  MUX2_X1 U330 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n365), .Z(n295) );
  MUX2_X1 U331 ( .A(n295), .B(n294), .S(n363), .Z(n296) );
  MUX2_X1 U332 ( .A(n296), .B(n293), .S(N12), .Z(N24) );
  MUX2_X1 U333 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n365), .Z(n297) );
  MUX2_X1 U334 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n365), .Z(n298) );
  MUX2_X1 U335 ( .A(n298), .B(n297), .S(n363), .Z(n299) );
  MUX2_X1 U336 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n365), .Z(n300) );
  MUX2_X1 U337 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n365), .Z(n301) );
  MUX2_X1 U338 ( .A(n301), .B(n300), .S(n363), .Z(n302) );
  MUX2_X1 U339 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n365), .Z(n303) );
  MUX2_X1 U340 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n365), .Z(n304) );
  MUX2_X1 U341 ( .A(n304), .B(n303), .S(n363), .Z(n305) );
  MUX2_X1 U342 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n365), .Z(n306) );
  MUX2_X1 U343 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n365), .Z(n307) );
  MUX2_X1 U344 ( .A(n307), .B(n306), .S(n363), .Z(n308) );
  MUX2_X1 U345 ( .A(n308), .B(n305), .S(N12), .Z(N22) );
  MUX2_X1 U346 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n366), .Z(n309) );
  MUX2_X1 U347 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n366), .Z(n310) );
  MUX2_X1 U348 ( .A(n310), .B(n309), .S(n363), .Z(n311) );
  MUX2_X1 U349 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n366), .Z(n312) );
  MUX2_X1 U350 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n366), .Z(n313) );
  MUX2_X1 U351 ( .A(n313), .B(n312), .S(n363), .Z(n314) );
  MUX2_X1 U352 ( .A(n314), .B(n311), .S(N12), .Z(N21) );
  MUX2_X1 U353 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n366), .Z(n315) );
  MUX2_X1 U354 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n366), .Z(n316) );
  MUX2_X1 U355 ( .A(n316), .B(n315), .S(n363), .Z(n317) );
  MUX2_X1 U356 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n366), .Z(n318) );
  MUX2_X1 U357 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n366), .Z(n319) );
  MUX2_X1 U358 ( .A(n319), .B(n318), .S(n363), .Z(n320) );
  MUX2_X1 U359 ( .A(n320), .B(n317), .S(N12), .Z(N20) );
  MUX2_X1 U360 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n366), .Z(n321) );
  MUX2_X1 U361 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n366), .Z(n322) );
  MUX2_X1 U362 ( .A(n322), .B(n321), .S(n363), .Z(n323) );
  MUX2_X1 U363 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n366), .Z(n324) );
  MUX2_X1 U364 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n366), .Z(n325) );
  MUX2_X1 U365 ( .A(n325), .B(n324), .S(n363), .Z(n326) );
  MUX2_X1 U366 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n364), .Z(n327) );
  MUX2_X1 U367 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n366), .Z(n328) );
  MUX2_X1 U368 ( .A(n328), .B(n327), .S(n363), .Z(n329) );
  MUX2_X1 U369 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n366), .Z(n330) );
  MUX2_X1 U370 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n365), .Z(n331) );
  MUX2_X1 U371 ( .A(n331), .B(n330), .S(n363), .Z(n332) );
  MUX2_X1 U372 ( .A(n332), .B(n329), .S(N12), .Z(N18) );
  MUX2_X1 U373 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n366), .Z(n333) );
  MUX2_X1 U374 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n364), .Z(n334) );
  MUX2_X1 U375 ( .A(n334), .B(n333), .S(N11), .Z(n335) );
  MUX2_X1 U376 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n365), .Z(n336) );
  MUX2_X1 U377 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n366), .Z(n337) );
  MUX2_X1 U378 ( .A(n337), .B(n336), .S(N11), .Z(n338) );
  MUX2_X1 U379 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n365), .Z(n339) );
  MUX2_X1 U380 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n364), .Z(n340) );
  MUX2_X1 U381 ( .A(n340), .B(n339), .S(n363), .Z(n341) );
  MUX2_X1 U382 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n364), .Z(n342) );
  MUX2_X1 U383 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n366), .Z(n343) );
  MUX2_X1 U384 ( .A(n343), .B(n342), .S(n363), .Z(n344) );
  MUX2_X1 U385 ( .A(n344), .B(n341), .S(N12), .Z(N16) );
  MUX2_X1 U386 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n365), .Z(n345) );
  MUX2_X1 U387 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n366), .Z(n346) );
  MUX2_X1 U388 ( .A(n346), .B(n345), .S(N11), .Z(n347) );
  MUX2_X1 U389 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n365), .Z(n348) );
  MUX2_X1 U390 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(N10), .Z(n349) );
  MUX2_X1 U391 ( .A(n349), .B(n348), .S(N11), .Z(n350) );
  MUX2_X1 U392 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n364), .Z(n351) );
  MUX2_X1 U393 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n366), .Z(n352) );
  MUX2_X1 U394 ( .A(n352), .B(n351), .S(n363), .Z(n353) );
  MUX2_X1 U395 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n365), .Z(n354) );
  MUX2_X1 U396 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n364), .Z(n355) );
  MUX2_X1 U397 ( .A(n355), .B(n354), .S(N11), .Z(n356) );
  MUX2_X1 U398 ( .A(n356), .B(n353), .S(N12), .Z(N14) );
  MUX2_X1 U399 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n365), .Z(n357) );
  MUX2_X1 U400 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n364), .Z(n358) );
  MUX2_X1 U401 ( .A(n358), .B(n357), .S(n363), .Z(n359) );
  MUX2_X1 U402 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n366), .Z(n360) );
  MUX2_X1 U403 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n364), .Z(n361) );
  MUX2_X1 U404 ( .A(n361), .B(n360), .S(N11), .Z(n362) );
  MUX2_X1 U405 ( .A(n362), .B(n359), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH16_SIZE8_LOGSIZE3_6 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] ,
         \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][15] , \mem[6][14] , \mem[6][13] ,
         \mem[6][12] , \mem[6][11] , \mem[6][10] , \mem[6][9] , \mem[6][8] ,
         \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] ,
         \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[5][15] , \mem[5][14] ,
         \mem[5][13] , \mem[5][12] , \mem[5][11] , \mem[5][10] , \mem[5][9] ,
         \mem[5][8] , \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] ,
         \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][15] ,
         \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] , \mem[4][10] ,
         \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14, N16, N18,
         N20, N22, N25, N26, N28, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[14]  ( .D(N14), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N16), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N18), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[8]  ( .D(N20), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N22), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[3]  ( .D(N25), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N26), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N28), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][15]  ( .D(n394), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n395), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n396), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n397), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n398), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n399), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n400), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n401), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n402), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n403), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n404), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n405), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n406), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n407), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n408), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n409), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n410), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n411), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n412), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n413), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n414), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n415), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n416), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n417), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n418), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n419), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n420), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n421), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n422), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n423), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n424), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n425), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n426), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n427), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n428), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n429), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n430), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n431), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n432), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n433), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n434), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n435), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n436), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n437), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n438), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n439), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n440), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n441), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n442), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n443), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n444), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n445), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n446), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n447), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n448), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n449), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n450), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n451), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n452), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n453), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n454), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n455), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n456), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n457), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n458), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n459), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n460), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n461), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n462), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n463), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n464), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n465), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n466), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n467), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n468), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n469), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n470), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n471), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n472), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n473), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n474), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n475), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n476), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n477), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n478), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n479), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n480), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n481), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n482), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n483), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n484), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n485), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n486), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n487), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n488), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n489), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n490), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n491), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n492), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n493), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n494), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n495), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n496), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n497), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n498), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n499), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n500), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n501), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n502), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n503), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n504), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n505), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n506), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n507), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n508), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n509), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n510), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n511), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n512), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n513), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n514), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n515), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n516), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n517), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n518), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n519), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n520), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n521), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U280 ( .A1(n375), .A2(n376), .A3(n642), .ZN(n659) );
  NAND3_X1 U281 ( .A1(n642), .A2(n376), .A3(N10), .ZN(n641) );
  NAND3_X1 U282 ( .A1(n642), .A2(n375), .A3(N11), .ZN(n624) );
  NAND3_X1 U283 ( .A1(N10), .A2(n642), .A3(N11), .ZN(n607) );
  NAND3_X1 U284 ( .A1(n375), .A2(n376), .A3(n573), .ZN(n590) );
  NAND3_X1 U285 ( .A1(N10), .A2(n376), .A3(n573), .ZN(n572) );
  NAND3_X1 U286 ( .A1(N11), .A2(n375), .A3(n573), .ZN(n555) );
  NAND3_X1 U287 ( .A1(N11), .A2(N10), .A3(n573), .ZN(n538) );
  SDFF_X1 \data_out_reg[5]  ( .D(n302), .SI(n299), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n338), .SI(n335), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n314), .SI(n311), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n350), .SI(n347), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n362), .SI(n359), .SE(N12), .CK(clk), .Q(
        data_out[15]) );
  SDFF_X1 \data_out_reg[4]  ( .D(n296), .SI(n293), .SE(N12), .CK(clk), .Q(
        data_out[4]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n12), .SI(n9), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n326), .SI(n323), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  BUF_X1 U3 ( .A(N10), .Z(n365) );
  BUF_X1 U4 ( .A(N10), .Z(n366) );
  BUF_X1 U5 ( .A(n659), .Z(n374) );
  BUF_X1 U6 ( .A(n641), .Z(n373) );
  BUF_X1 U7 ( .A(n607), .Z(n371) );
  BUF_X1 U8 ( .A(n590), .Z(n370) );
  BUF_X1 U9 ( .A(n555), .Z(n368) );
  BUF_X1 U10 ( .A(n572), .Z(n369) );
  BUF_X1 U11 ( .A(n538), .Z(n367) );
  BUF_X1 U12 ( .A(n624), .Z(n372) );
  BUF_X1 U13 ( .A(N10), .Z(n364) );
  BUF_X1 U14 ( .A(N11), .Z(n363) );
  NOR2_X1 U15 ( .A1(n377), .A2(N12), .ZN(n642) );
  INV_X1 U16 ( .A(wr_en), .ZN(n377) );
  AND2_X1 U17 ( .A1(N12), .A2(wr_en), .ZN(n573) );
  OAI21_X1 U18 ( .B1(n386), .B2(n607), .A(n599), .ZN(n466) );
  NAND2_X1 U19 ( .A1(\mem[3][7] ), .A2(n371), .ZN(n599) );
  OAI21_X1 U20 ( .B1(n385), .B2(n371), .A(n598), .ZN(n465) );
  NAND2_X1 U21 ( .A1(\mem[3][8] ), .A2(n371), .ZN(n598) );
  OAI21_X1 U22 ( .B1(n384), .B2(n607), .A(n597), .ZN(n464) );
  NAND2_X1 U23 ( .A1(\mem[3][9] ), .A2(n371), .ZN(n597) );
  OAI21_X1 U24 ( .B1(n383), .B2(n607), .A(n596), .ZN(n463) );
  NAND2_X1 U25 ( .A1(\mem[3][10] ), .A2(n371), .ZN(n596) );
  OAI21_X1 U26 ( .B1(n382), .B2(n607), .A(n595), .ZN(n462) );
  NAND2_X1 U27 ( .A1(\mem[3][11] ), .A2(n371), .ZN(n595) );
  OAI21_X1 U28 ( .B1(n381), .B2(n607), .A(n594), .ZN(n461) );
  NAND2_X1 U29 ( .A1(\mem[3][12] ), .A2(n371), .ZN(n594) );
  OAI21_X1 U30 ( .B1(n380), .B2(n607), .A(n593), .ZN(n460) );
  NAND2_X1 U31 ( .A1(\mem[3][13] ), .A2(n371), .ZN(n593) );
  OAI21_X1 U32 ( .B1(n379), .B2(n607), .A(n592), .ZN(n459) );
  NAND2_X1 U33 ( .A1(\mem[3][14] ), .A2(n371), .ZN(n592) );
  OAI21_X1 U34 ( .B1(n386), .B2(n572), .A(n564), .ZN(n434) );
  NAND2_X1 U35 ( .A1(\mem[5][7] ), .A2(n369), .ZN(n564) );
  OAI21_X1 U36 ( .B1(n385), .B2(n572), .A(n563), .ZN(n433) );
  NAND2_X1 U37 ( .A1(\mem[5][8] ), .A2(n572), .ZN(n563) );
  OAI21_X1 U38 ( .B1(n384), .B2(n572), .A(n562), .ZN(n432) );
  NAND2_X1 U39 ( .A1(\mem[5][9] ), .A2(n572), .ZN(n562) );
  OAI21_X1 U40 ( .B1(n383), .B2(n572), .A(n561), .ZN(n431) );
  NAND2_X1 U41 ( .A1(\mem[5][10] ), .A2(n572), .ZN(n561) );
  OAI21_X1 U42 ( .B1(n382), .B2(n572), .A(n560), .ZN(n430) );
  NAND2_X1 U43 ( .A1(\mem[5][11] ), .A2(n572), .ZN(n560) );
  OAI21_X1 U44 ( .B1(n381), .B2(n572), .A(n559), .ZN(n429) );
  NAND2_X1 U45 ( .A1(\mem[5][12] ), .A2(n572), .ZN(n559) );
  OAI21_X1 U46 ( .B1(n380), .B2(n572), .A(n558), .ZN(n428) );
  NAND2_X1 U47 ( .A1(\mem[5][13] ), .A2(n572), .ZN(n558) );
  OAI21_X1 U48 ( .B1(n379), .B2(n572), .A(n557), .ZN(n427) );
  NAND2_X1 U49 ( .A1(\mem[5][14] ), .A2(n572), .ZN(n557) );
  OAI21_X1 U50 ( .B1(n386), .B2(n538), .A(n530), .ZN(n402) );
  NAND2_X1 U51 ( .A1(\mem[7][7] ), .A2(n367), .ZN(n530) );
  OAI21_X1 U52 ( .B1(n385), .B2(n538), .A(n529), .ZN(n401) );
  NAND2_X1 U53 ( .A1(\mem[7][8] ), .A2(n538), .ZN(n529) );
  OAI21_X1 U54 ( .B1(n384), .B2(n538), .A(n528), .ZN(n400) );
  NAND2_X1 U55 ( .A1(\mem[7][9] ), .A2(n538), .ZN(n528) );
  OAI21_X1 U56 ( .B1(n383), .B2(n538), .A(n527), .ZN(n399) );
  NAND2_X1 U57 ( .A1(\mem[7][10] ), .A2(n538), .ZN(n527) );
  OAI21_X1 U58 ( .B1(n382), .B2(n538), .A(n526), .ZN(n398) );
  NAND2_X1 U59 ( .A1(\mem[7][11] ), .A2(n538), .ZN(n526) );
  OAI21_X1 U60 ( .B1(n381), .B2(n538), .A(n525), .ZN(n397) );
  NAND2_X1 U61 ( .A1(\mem[7][12] ), .A2(n538), .ZN(n525) );
  OAI21_X1 U62 ( .B1(n380), .B2(n538), .A(n524), .ZN(n396) );
  NAND2_X1 U63 ( .A1(\mem[7][13] ), .A2(n538), .ZN(n524) );
  OAI21_X1 U64 ( .B1(n379), .B2(n538), .A(n523), .ZN(n395) );
  NAND2_X1 U65 ( .A1(\mem[7][14] ), .A2(n538), .ZN(n523) );
  OAI21_X1 U66 ( .B1(n386), .B2(n641), .A(n633), .ZN(n498) );
  NAND2_X1 U67 ( .A1(\mem[1][7] ), .A2(n373), .ZN(n633) );
  OAI21_X1 U68 ( .B1(n385), .B2(n373), .A(n632), .ZN(n497) );
  NAND2_X1 U69 ( .A1(\mem[1][8] ), .A2(n373), .ZN(n632) );
  OAI21_X1 U70 ( .B1(n384), .B2(n641), .A(n631), .ZN(n496) );
  NAND2_X1 U71 ( .A1(\mem[1][9] ), .A2(n373), .ZN(n631) );
  OAI21_X1 U72 ( .B1(n383), .B2(n641), .A(n630), .ZN(n495) );
  NAND2_X1 U73 ( .A1(\mem[1][10] ), .A2(n373), .ZN(n630) );
  OAI21_X1 U74 ( .B1(n382), .B2(n641), .A(n629), .ZN(n494) );
  NAND2_X1 U75 ( .A1(\mem[1][11] ), .A2(n373), .ZN(n629) );
  OAI21_X1 U76 ( .B1(n381), .B2(n641), .A(n628), .ZN(n493) );
  NAND2_X1 U77 ( .A1(\mem[1][12] ), .A2(n373), .ZN(n628) );
  OAI21_X1 U78 ( .B1(n380), .B2(n641), .A(n627), .ZN(n492) );
  NAND2_X1 U79 ( .A1(\mem[1][13] ), .A2(n373), .ZN(n627) );
  OAI21_X1 U80 ( .B1(n379), .B2(n641), .A(n626), .ZN(n491) );
  NAND2_X1 U81 ( .A1(\mem[1][14] ), .A2(n373), .ZN(n626) );
  OAI21_X1 U82 ( .B1(n386), .B2(n555), .A(n547), .ZN(n418) );
  NAND2_X1 U83 ( .A1(\mem[6][7] ), .A2(n368), .ZN(n547) );
  OAI21_X1 U84 ( .B1(n385), .B2(n368), .A(n546), .ZN(n417) );
  NAND2_X1 U85 ( .A1(\mem[6][8] ), .A2(n368), .ZN(n546) );
  OAI21_X1 U86 ( .B1(n384), .B2(n555), .A(n545), .ZN(n416) );
  NAND2_X1 U87 ( .A1(\mem[6][9] ), .A2(n368), .ZN(n545) );
  OAI21_X1 U88 ( .B1(n383), .B2(n555), .A(n544), .ZN(n415) );
  NAND2_X1 U89 ( .A1(\mem[6][10] ), .A2(n368), .ZN(n544) );
  OAI21_X1 U90 ( .B1(n382), .B2(n555), .A(n543), .ZN(n414) );
  NAND2_X1 U91 ( .A1(\mem[6][11] ), .A2(n368), .ZN(n543) );
  OAI21_X1 U92 ( .B1(n381), .B2(n555), .A(n542), .ZN(n413) );
  NAND2_X1 U93 ( .A1(\mem[6][12] ), .A2(n368), .ZN(n542) );
  OAI21_X1 U94 ( .B1(n380), .B2(n555), .A(n541), .ZN(n412) );
  NAND2_X1 U95 ( .A1(\mem[6][13] ), .A2(n368), .ZN(n541) );
  OAI21_X1 U96 ( .B1(n379), .B2(n555), .A(n540), .ZN(n411) );
  NAND2_X1 U97 ( .A1(\mem[6][14] ), .A2(n368), .ZN(n540) );
  OAI21_X1 U98 ( .B1(n380), .B2(n372), .A(n610), .ZN(n476) );
  NAND2_X1 U99 ( .A1(\mem[2][13] ), .A2(n624), .ZN(n610) );
  OAI21_X1 U100 ( .B1(n386), .B2(n372), .A(n616), .ZN(n482) );
  NAND2_X1 U101 ( .A1(\mem[2][7] ), .A2(n372), .ZN(n616) );
  OAI21_X1 U102 ( .B1(n385), .B2(n372), .A(n615), .ZN(n481) );
  NAND2_X1 U103 ( .A1(\mem[2][8] ), .A2(n624), .ZN(n615) );
  OAI21_X1 U104 ( .B1(n384), .B2(n372), .A(n614), .ZN(n480) );
  NAND2_X1 U105 ( .A1(\mem[2][9] ), .A2(n624), .ZN(n614) );
  OAI21_X1 U106 ( .B1(n383), .B2(n372), .A(n613), .ZN(n479) );
  NAND2_X1 U107 ( .A1(\mem[2][10] ), .A2(n624), .ZN(n613) );
  OAI21_X1 U108 ( .B1(n382), .B2(n372), .A(n612), .ZN(n478) );
  NAND2_X1 U109 ( .A1(\mem[2][11] ), .A2(n624), .ZN(n612) );
  OAI21_X1 U110 ( .B1(n381), .B2(n372), .A(n611), .ZN(n477) );
  NAND2_X1 U111 ( .A1(\mem[2][12] ), .A2(n624), .ZN(n611) );
  OAI21_X1 U112 ( .B1(n379), .B2(n372), .A(n609), .ZN(n475) );
  NAND2_X1 U113 ( .A1(\mem[2][14] ), .A2(n624), .ZN(n609) );
  OAI21_X1 U114 ( .B1(n386), .B2(n590), .A(n582), .ZN(n450) );
  NAND2_X1 U115 ( .A1(\mem[4][7] ), .A2(n370), .ZN(n582) );
  OAI21_X1 U116 ( .B1(n385), .B2(n370), .A(n581), .ZN(n449) );
  NAND2_X1 U117 ( .A1(\mem[4][8] ), .A2(n370), .ZN(n581) );
  OAI21_X1 U118 ( .B1(n384), .B2(n590), .A(n580), .ZN(n448) );
  NAND2_X1 U119 ( .A1(\mem[4][9] ), .A2(n370), .ZN(n580) );
  OAI21_X1 U120 ( .B1(n383), .B2(n590), .A(n579), .ZN(n447) );
  NAND2_X1 U121 ( .A1(\mem[4][10] ), .A2(n370), .ZN(n579) );
  OAI21_X1 U122 ( .B1(n382), .B2(n590), .A(n578), .ZN(n446) );
  NAND2_X1 U123 ( .A1(\mem[4][11] ), .A2(n370), .ZN(n578) );
  OAI21_X1 U124 ( .B1(n381), .B2(n590), .A(n577), .ZN(n445) );
  NAND2_X1 U125 ( .A1(\mem[4][12] ), .A2(n370), .ZN(n577) );
  OAI21_X1 U126 ( .B1(n380), .B2(n590), .A(n576), .ZN(n444) );
  NAND2_X1 U127 ( .A1(\mem[4][13] ), .A2(n370), .ZN(n576) );
  OAI21_X1 U128 ( .B1(n379), .B2(n590), .A(n575), .ZN(n443) );
  NAND2_X1 U129 ( .A1(\mem[4][14] ), .A2(n370), .ZN(n575) );
  OAI21_X1 U130 ( .B1(n659), .B2(n385), .A(n650), .ZN(n513) );
  NAND2_X1 U131 ( .A1(\mem[0][8] ), .A2(n374), .ZN(n650) );
  OAI21_X1 U132 ( .B1(n659), .B2(n384), .A(n649), .ZN(n512) );
  NAND2_X1 U133 ( .A1(\mem[0][9] ), .A2(n659), .ZN(n649) );
  OAI21_X1 U134 ( .B1(n374), .B2(n383), .A(n648), .ZN(n511) );
  NAND2_X1 U135 ( .A1(\mem[0][10] ), .A2(n659), .ZN(n648) );
  OAI21_X1 U136 ( .B1(n659), .B2(n382), .A(n647), .ZN(n510) );
  NAND2_X1 U137 ( .A1(\mem[0][11] ), .A2(n659), .ZN(n647) );
  OAI21_X1 U138 ( .B1(n659), .B2(n381), .A(n646), .ZN(n509) );
  NAND2_X1 U139 ( .A1(\mem[0][12] ), .A2(n659), .ZN(n646) );
  OAI21_X1 U140 ( .B1(n659), .B2(n380), .A(n645), .ZN(n508) );
  NAND2_X1 U141 ( .A1(\mem[0][13] ), .A2(n659), .ZN(n645) );
  OAI21_X1 U142 ( .B1(n659), .B2(n379), .A(n644), .ZN(n507) );
  NAND2_X1 U143 ( .A1(\mem[0][14] ), .A2(n659), .ZN(n644) );
  INV_X1 U144 ( .A(N10), .ZN(n375) );
  OAI21_X1 U145 ( .B1(n393), .B2(n641), .A(n640), .ZN(n505) );
  NAND2_X1 U146 ( .A1(\mem[1][0] ), .A2(n373), .ZN(n640) );
  OAI21_X1 U147 ( .B1(n392), .B2(n641), .A(n639), .ZN(n504) );
  NAND2_X1 U148 ( .A1(\mem[1][1] ), .A2(n373), .ZN(n639) );
  OAI21_X1 U149 ( .B1(n391), .B2(n641), .A(n638), .ZN(n503) );
  NAND2_X1 U150 ( .A1(\mem[1][2] ), .A2(n373), .ZN(n638) );
  OAI21_X1 U151 ( .B1(n390), .B2(n641), .A(n637), .ZN(n502) );
  NAND2_X1 U152 ( .A1(\mem[1][3] ), .A2(n373), .ZN(n637) );
  OAI21_X1 U153 ( .B1(n389), .B2(n641), .A(n636), .ZN(n501) );
  NAND2_X1 U154 ( .A1(\mem[1][4] ), .A2(n641), .ZN(n636) );
  OAI21_X1 U155 ( .B1(n388), .B2(n641), .A(n635), .ZN(n500) );
  NAND2_X1 U156 ( .A1(\mem[1][5] ), .A2(n641), .ZN(n635) );
  OAI21_X1 U157 ( .B1(n387), .B2(n641), .A(n634), .ZN(n499) );
  NAND2_X1 U158 ( .A1(\mem[1][6] ), .A2(n641), .ZN(n634) );
  OAI21_X1 U159 ( .B1(n378), .B2(n641), .A(n625), .ZN(n490) );
  NAND2_X1 U160 ( .A1(\mem[1][15] ), .A2(n373), .ZN(n625) );
  OAI21_X1 U161 ( .B1(n393), .B2(n372), .A(n623), .ZN(n489) );
  NAND2_X1 U162 ( .A1(\mem[2][0] ), .A2(n372), .ZN(n623) );
  OAI21_X1 U163 ( .B1(n392), .B2(n624), .A(n622), .ZN(n488) );
  NAND2_X1 U164 ( .A1(\mem[2][1] ), .A2(n624), .ZN(n622) );
  OAI21_X1 U165 ( .B1(n391), .B2(n372), .A(n621), .ZN(n487) );
  NAND2_X1 U166 ( .A1(\mem[2][2] ), .A2(n624), .ZN(n621) );
  OAI21_X1 U167 ( .B1(n390), .B2(n624), .A(n620), .ZN(n486) );
  NAND2_X1 U168 ( .A1(\mem[2][3] ), .A2(n624), .ZN(n620) );
  OAI21_X1 U169 ( .B1(n389), .B2(n624), .A(n619), .ZN(n485) );
  NAND2_X1 U170 ( .A1(\mem[2][4] ), .A2(n372), .ZN(n619) );
  OAI21_X1 U171 ( .B1(n388), .B2(n624), .A(n618), .ZN(n484) );
  NAND2_X1 U172 ( .A1(\mem[2][5] ), .A2(n372), .ZN(n618) );
  OAI21_X1 U173 ( .B1(n387), .B2(n624), .A(n617), .ZN(n483) );
  NAND2_X1 U174 ( .A1(\mem[2][6] ), .A2(n372), .ZN(n617) );
  OAI21_X1 U175 ( .B1(n378), .B2(n624), .A(n608), .ZN(n474) );
  NAND2_X1 U176 ( .A1(\mem[2][15] ), .A2(n624), .ZN(n608) );
  OAI21_X1 U177 ( .B1(n393), .B2(n607), .A(n606), .ZN(n473) );
  NAND2_X1 U178 ( .A1(\mem[3][0] ), .A2(n371), .ZN(n606) );
  OAI21_X1 U179 ( .B1(n392), .B2(n607), .A(n605), .ZN(n472) );
  NAND2_X1 U180 ( .A1(\mem[3][1] ), .A2(n371), .ZN(n605) );
  OAI21_X1 U181 ( .B1(n391), .B2(n607), .A(n604), .ZN(n471) );
  NAND2_X1 U182 ( .A1(\mem[3][2] ), .A2(n371), .ZN(n604) );
  OAI21_X1 U183 ( .B1(n390), .B2(n607), .A(n603), .ZN(n470) );
  NAND2_X1 U184 ( .A1(\mem[3][3] ), .A2(n371), .ZN(n603) );
  OAI21_X1 U185 ( .B1(n389), .B2(n607), .A(n602), .ZN(n469) );
  NAND2_X1 U186 ( .A1(\mem[3][4] ), .A2(n607), .ZN(n602) );
  OAI21_X1 U187 ( .B1(n388), .B2(n607), .A(n601), .ZN(n468) );
  NAND2_X1 U188 ( .A1(\mem[3][5] ), .A2(n607), .ZN(n601) );
  OAI21_X1 U189 ( .B1(n387), .B2(n607), .A(n600), .ZN(n467) );
  NAND2_X1 U190 ( .A1(\mem[3][6] ), .A2(n607), .ZN(n600) );
  OAI21_X1 U191 ( .B1(n378), .B2(n607), .A(n591), .ZN(n458) );
  NAND2_X1 U192 ( .A1(\mem[3][15] ), .A2(n371), .ZN(n591) );
  OAI21_X1 U193 ( .B1(n393), .B2(n590), .A(n589), .ZN(n457) );
  NAND2_X1 U194 ( .A1(\mem[4][0] ), .A2(n370), .ZN(n589) );
  OAI21_X1 U195 ( .B1(n392), .B2(n590), .A(n588), .ZN(n456) );
  NAND2_X1 U196 ( .A1(\mem[4][1] ), .A2(n370), .ZN(n588) );
  OAI21_X1 U197 ( .B1(n391), .B2(n590), .A(n587), .ZN(n455) );
  NAND2_X1 U198 ( .A1(\mem[4][2] ), .A2(n370), .ZN(n587) );
  OAI21_X1 U199 ( .B1(n390), .B2(n590), .A(n586), .ZN(n454) );
  NAND2_X1 U200 ( .A1(\mem[4][3] ), .A2(n370), .ZN(n586) );
  OAI21_X1 U201 ( .B1(n389), .B2(n590), .A(n585), .ZN(n453) );
  NAND2_X1 U202 ( .A1(\mem[4][4] ), .A2(n590), .ZN(n585) );
  OAI21_X1 U203 ( .B1(n388), .B2(n590), .A(n584), .ZN(n452) );
  NAND2_X1 U204 ( .A1(\mem[4][5] ), .A2(n590), .ZN(n584) );
  OAI21_X1 U205 ( .B1(n387), .B2(n590), .A(n583), .ZN(n451) );
  NAND2_X1 U206 ( .A1(\mem[4][6] ), .A2(n590), .ZN(n583) );
  OAI21_X1 U207 ( .B1(n378), .B2(n590), .A(n574), .ZN(n442) );
  NAND2_X1 U208 ( .A1(\mem[4][15] ), .A2(n370), .ZN(n574) );
  OAI21_X1 U209 ( .B1(n393), .B2(n369), .A(n571), .ZN(n441) );
  NAND2_X1 U210 ( .A1(\mem[5][0] ), .A2(n369), .ZN(n571) );
  OAI21_X1 U211 ( .B1(n392), .B2(n369), .A(n570), .ZN(n440) );
  NAND2_X1 U212 ( .A1(\mem[5][1] ), .A2(n572), .ZN(n570) );
  OAI21_X1 U213 ( .B1(n391), .B2(n369), .A(n569), .ZN(n439) );
  NAND2_X1 U214 ( .A1(\mem[5][2] ), .A2(n572), .ZN(n569) );
  OAI21_X1 U215 ( .B1(n390), .B2(n369), .A(n568), .ZN(n438) );
  NAND2_X1 U216 ( .A1(\mem[5][3] ), .A2(n572), .ZN(n568) );
  OAI21_X1 U217 ( .B1(n389), .B2(n369), .A(n567), .ZN(n437) );
  NAND2_X1 U218 ( .A1(\mem[5][4] ), .A2(n369), .ZN(n567) );
  OAI21_X1 U219 ( .B1(n388), .B2(n369), .A(n566), .ZN(n436) );
  NAND2_X1 U220 ( .A1(\mem[5][5] ), .A2(n369), .ZN(n566) );
  OAI21_X1 U221 ( .B1(n387), .B2(n369), .A(n565), .ZN(n435) );
  NAND2_X1 U222 ( .A1(\mem[5][6] ), .A2(n369), .ZN(n565) );
  OAI21_X1 U223 ( .B1(n378), .B2(n369), .A(n556), .ZN(n426) );
  NAND2_X1 U224 ( .A1(\mem[5][15] ), .A2(n369), .ZN(n556) );
  OAI21_X1 U225 ( .B1(n393), .B2(n555), .A(n554), .ZN(n425) );
  NAND2_X1 U226 ( .A1(\mem[6][0] ), .A2(n368), .ZN(n554) );
  OAI21_X1 U227 ( .B1(n392), .B2(n555), .A(n553), .ZN(n424) );
  NAND2_X1 U228 ( .A1(\mem[6][1] ), .A2(n368), .ZN(n553) );
  OAI21_X1 U229 ( .B1(n391), .B2(n555), .A(n552), .ZN(n423) );
  NAND2_X1 U230 ( .A1(\mem[6][2] ), .A2(n368), .ZN(n552) );
  OAI21_X1 U231 ( .B1(n390), .B2(n555), .A(n551), .ZN(n422) );
  NAND2_X1 U232 ( .A1(\mem[6][3] ), .A2(n368), .ZN(n551) );
  OAI21_X1 U233 ( .B1(n389), .B2(n555), .A(n550), .ZN(n421) );
  NAND2_X1 U234 ( .A1(\mem[6][4] ), .A2(n555), .ZN(n550) );
  OAI21_X1 U235 ( .B1(n388), .B2(n555), .A(n549), .ZN(n420) );
  NAND2_X1 U236 ( .A1(\mem[6][5] ), .A2(n555), .ZN(n549) );
  OAI21_X1 U237 ( .B1(n387), .B2(n555), .A(n548), .ZN(n419) );
  NAND2_X1 U238 ( .A1(\mem[6][6] ), .A2(n555), .ZN(n548) );
  OAI21_X1 U239 ( .B1(n378), .B2(n555), .A(n539), .ZN(n410) );
  NAND2_X1 U240 ( .A1(\mem[6][15] ), .A2(n368), .ZN(n539) );
  OAI21_X1 U241 ( .B1(n393), .B2(n367), .A(n537), .ZN(n409) );
  NAND2_X1 U242 ( .A1(\mem[7][0] ), .A2(n367), .ZN(n537) );
  OAI21_X1 U243 ( .B1(n392), .B2(n367), .A(n536), .ZN(n408) );
  NAND2_X1 U244 ( .A1(\mem[7][1] ), .A2(n538), .ZN(n536) );
  OAI21_X1 U245 ( .B1(n391), .B2(n367), .A(n535), .ZN(n407) );
  NAND2_X1 U246 ( .A1(\mem[7][2] ), .A2(n538), .ZN(n535) );
  OAI21_X1 U247 ( .B1(n390), .B2(n367), .A(n534), .ZN(n406) );
  NAND2_X1 U248 ( .A1(\mem[7][3] ), .A2(n538), .ZN(n534) );
  OAI21_X1 U249 ( .B1(n389), .B2(n367), .A(n533), .ZN(n405) );
  NAND2_X1 U250 ( .A1(\mem[7][4] ), .A2(n367), .ZN(n533) );
  OAI21_X1 U251 ( .B1(n388), .B2(n367), .A(n532), .ZN(n404) );
  NAND2_X1 U252 ( .A1(\mem[7][5] ), .A2(n367), .ZN(n532) );
  OAI21_X1 U253 ( .B1(n387), .B2(n367), .A(n531), .ZN(n403) );
  NAND2_X1 U254 ( .A1(\mem[7][6] ), .A2(n367), .ZN(n531) );
  OAI21_X1 U255 ( .B1(n378), .B2(n367), .A(n522), .ZN(n394) );
  NAND2_X1 U256 ( .A1(\mem[7][15] ), .A2(n367), .ZN(n522) );
  OAI21_X1 U257 ( .B1(n374), .B2(n393), .A(n658), .ZN(n521) );
  NAND2_X1 U258 ( .A1(\mem[0][0] ), .A2(n659), .ZN(n658) );
  OAI21_X1 U259 ( .B1(n374), .B2(n392), .A(n657), .ZN(n520) );
  NAND2_X1 U260 ( .A1(\mem[0][1] ), .A2(n659), .ZN(n657) );
  OAI21_X1 U261 ( .B1(n374), .B2(n391), .A(n656), .ZN(n519) );
  NAND2_X1 U262 ( .A1(\mem[0][2] ), .A2(n659), .ZN(n656) );
  OAI21_X1 U263 ( .B1(n374), .B2(n390), .A(n655), .ZN(n518) );
  NAND2_X1 U264 ( .A1(\mem[0][3] ), .A2(n659), .ZN(n655) );
  OAI21_X1 U265 ( .B1(n374), .B2(n389), .A(n654), .ZN(n517) );
  NAND2_X1 U266 ( .A1(\mem[0][4] ), .A2(n374), .ZN(n654) );
  OAI21_X1 U267 ( .B1(n374), .B2(n388), .A(n653), .ZN(n516) );
  NAND2_X1 U268 ( .A1(\mem[0][5] ), .A2(n374), .ZN(n653) );
  OAI21_X1 U269 ( .B1(n374), .B2(n387), .A(n652), .ZN(n515) );
  NAND2_X1 U270 ( .A1(\mem[0][6] ), .A2(n374), .ZN(n652) );
  OAI21_X1 U271 ( .B1(n374), .B2(n386), .A(n651), .ZN(n514) );
  NAND2_X1 U272 ( .A1(\mem[0][7] ), .A2(n374), .ZN(n651) );
  OAI21_X1 U273 ( .B1(n374), .B2(n378), .A(n643), .ZN(n506) );
  NAND2_X1 U274 ( .A1(\mem[0][15] ), .A2(n659), .ZN(n643) );
  INV_X1 U275 ( .A(N11), .ZN(n376) );
  INV_X1 U276 ( .A(data_in[0]), .ZN(n393) );
  INV_X1 U277 ( .A(data_in[1]), .ZN(n392) );
  INV_X1 U278 ( .A(data_in[2]), .ZN(n391) );
  INV_X1 U279 ( .A(data_in[3]), .ZN(n390) );
  INV_X1 U288 ( .A(data_in[4]), .ZN(n389) );
  INV_X1 U289 ( .A(data_in[5]), .ZN(n388) );
  INV_X1 U290 ( .A(data_in[6]), .ZN(n387) );
  INV_X1 U291 ( .A(data_in[7]), .ZN(n386) );
  INV_X1 U292 ( .A(data_in[8]), .ZN(n385) );
  INV_X1 U293 ( .A(data_in[9]), .ZN(n384) );
  INV_X1 U294 ( .A(data_in[10]), .ZN(n383) );
  INV_X1 U295 ( .A(data_in[11]), .ZN(n382) );
  INV_X1 U296 ( .A(data_in[12]), .ZN(n381) );
  INV_X1 U297 ( .A(data_in[13]), .ZN(n380) );
  INV_X1 U298 ( .A(data_in[14]), .ZN(n379) );
  INV_X1 U299 ( .A(data_in[15]), .ZN(n378) );
  MUX2_X1 U300 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n364), .Z(n1) );
  MUX2_X1 U301 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n366), .Z(n2) );
  MUX2_X1 U302 ( .A(n2), .B(n1), .S(n363), .Z(n3) );
  MUX2_X1 U303 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n365), .Z(n4) );
  MUX2_X1 U304 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n365), .Z(n5) );
  MUX2_X1 U305 ( .A(n5), .B(n4), .S(N11), .Z(n6) );
  MUX2_X1 U306 ( .A(n6), .B(n3), .S(N12), .Z(N28) );
  MUX2_X1 U307 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n364), .Z(n7) );
  MUX2_X1 U308 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n364), .Z(n8) );
  MUX2_X1 U309 ( .A(n8), .B(n7), .S(N11), .Z(n9) );
  MUX2_X1 U310 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n364), .Z(n10) );
  MUX2_X1 U311 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n364), .Z(n11) );
  MUX2_X1 U312 ( .A(n11), .B(n10), .S(N11), .Z(n12) );
  MUX2_X1 U313 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n364), .Z(n13) );
  MUX2_X1 U314 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n364), .Z(n14) );
  MUX2_X1 U315 ( .A(n14), .B(n13), .S(N11), .Z(n15) );
  MUX2_X1 U316 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n364), .Z(n16) );
  MUX2_X1 U317 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n364), .Z(n17) );
  MUX2_X1 U318 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U319 ( .A(n18), .B(n15), .S(N12), .Z(N26) );
  MUX2_X1 U320 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n364), .Z(n19) );
  MUX2_X1 U321 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n364), .Z(n286) );
  MUX2_X1 U322 ( .A(n286), .B(n19), .S(N11), .Z(n287) );
  MUX2_X1 U323 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n364), .Z(n288) );
  MUX2_X1 U324 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n364), .Z(n289) );
  MUX2_X1 U325 ( .A(n289), .B(n288), .S(N11), .Z(n290) );
  MUX2_X1 U326 ( .A(n290), .B(n287), .S(N12), .Z(N25) );
  MUX2_X1 U327 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n365), .Z(n291) );
  MUX2_X1 U328 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n364), .Z(n292) );
  MUX2_X1 U329 ( .A(n292), .B(n291), .S(n363), .Z(n293) );
  MUX2_X1 U330 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n364), .Z(n294) );
  MUX2_X1 U331 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n366), .Z(n295) );
  MUX2_X1 U332 ( .A(n295), .B(n294), .S(n363), .Z(n296) );
  MUX2_X1 U333 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n366), .Z(n297) );
  MUX2_X1 U334 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n365), .Z(n298) );
  MUX2_X1 U335 ( .A(n298), .B(n297), .S(n363), .Z(n299) );
  MUX2_X1 U336 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n365), .Z(n300) );
  MUX2_X1 U337 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n364), .Z(n301) );
  MUX2_X1 U338 ( .A(n301), .B(n300), .S(n363), .Z(n302) );
  MUX2_X1 U339 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n366), .Z(n303) );
  MUX2_X1 U340 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n365), .Z(n304) );
  MUX2_X1 U341 ( .A(n304), .B(n303), .S(n363), .Z(n305) );
  MUX2_X1 U342 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n364), .Z(n306) );
  MUX2_X1 U343 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n364), .Z(n307) );
  MUX2_X1 U344 ( .A(n307), .B(n306), .S(n363), .Z(n308) );
  MUX2_X1 U345 ( .A(n308), .B(n305), .S(N12), .Z(N22) );
  MUX2_X1 U346 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n364), .Z(n309) );
  MUX2_X1 U347 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n366), .Z(n310) );
  MUX2_X1 U348 ( .A(n310), .B(n309), .S(n363), .Z(n311) );
  MUX2_X1 U349 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n364), .Z(n312) );
  MUX2_X1 U350 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n365), .Z(n313) );
  MUX2_X1 U351 ( .A(n313), .B(n312), .S(n363), .Z(n314) );
  MUX2_X1 U352 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n364), .Z(n315) );
  MUX2_X1 U353 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n366), .Z(n316) );
  MUX2_X1 U354 ( .A(n316), .B(n315), .S(n363), .Z(n317) );
  MUX2_X1 U355 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n365), .Z(n318) );
  MUX2_X1 U356 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n366), .Z(n319) );
  MUX2_X1 U357 ( .A(n319), .B(n318), .S(n363), .Z(n320) );
  MUX2_X1 U358 ( .A(n320), .B(n317), .S(N12), .Z(N20) );
  MUX2_X1 U359 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n365), .Z(n321) );
  MUX2_X1 U360 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n366), .Z(n322) );
  MUX2_X1 U361 ( .A(n322), .B(n321), .S(n363), .Z(n323) );
  MUX2_X1 U362 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n365), .Z(n324) );
  MUX2_X1 U363 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n366), .Z(n325) );
  MUX2_X1 U364 ( .A(n325), .B(n324), .S(n363), .Z(n326) );
  MUX2_X1 U365 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n365), .Z(n327) );
  MUX2_X1 U366 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n365), .Z(n328) );
  MUX2_X1 U367 ( .A(n328), .B(n327), .S(n363), .Z(n329) );
  MUX2_X1 U368 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n365), .Z(n330) );
  MUX2_X1 U369 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n365), .Z(n331) );
  MUX2_X1 U370 ( .A(n331), .B(n330), .S(N11), .Z(n332) );
  MUX2_X1 U371 ( .A(n332), .B(n329), .S(N12), .Z(N18) );
  MUX2_X1 U372 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n365), .Z(n333) );
  MUX2_X1 U373 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n365), .Z(n334) );
  MUX2_X1 U374 ( .A(n334), .B(n333), .S(N11), .Z(n335) );
  MUX2_X1 U375 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n365), .Z(n336) );
  MUX2_X1 U376 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n365), .Z(n337) );
  MUX2_X1 U377 ( .A(n337), .B(n336), .S(N11), .Z(n338) );
  MUX2_X1 U378 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n365), .Z(n339) );
  MUX2_X1 U379 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n365), .Z(n340) );
  MUX2_X1 U380 ( .A(n340), .B(n339), .S(n363), .Z(n341) );
  MUX2_X1 U381 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n365), .Z(n342) );
  MUX2_X1 U382 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n365), .Z(n343) );
  MUX2_X1 U383 ( .A(n343), .B(n342), .S(N11), .Z(n344) );
  MUX2_X1 U384 ( .A(n344), .B(n341), .S(N12), .Z(N16) );
  MUX2_X1 U385 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n366), .Z(n345) );
  MUX2_X1 U386 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n366), .Z(n346) );
  MUX2_X1 U387 ( .A(n346), .B(n345), .S(N11), .Z(n347) );
  MUX2_X1 U388 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n366), .Z(n348) );
  MUX2_X1 U389 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n366), .Z(n349) );
  MUX2_X1 U390 ( .A(n349), .B(n348), .S(N11), .Z(n350) );
  MUX2_X1 U391 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n366), .Z(n351) );
  MUX2_X1 U392 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n366), .Z(n352) );
  MUX2_X1 U393 ( .A(n352), .B(n351), .S(N11), .Z(n353) );
  MUX2_X1 U394 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n366), .Z(n354) );
  MUX2_X1 U395 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n366), .Z(n355) );
  MUX2_X1 U396 ( .A(n355), .B(n354), .S(N11), .Z(n356) );
  MUX2_X1 U397 ( .A(n356), .B(n353), .S(N12), .Z(N14) );
  MUX2_X1 U398 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n366), .Z(n357) );
  MUX2_X1 U399 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n366), .Z(n358) );
  MUX2_X1 U400 ( .A(n358), .B(n357), .S(N11), .Z(n359) );
  MUX2_X1 U401 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n366), .Z(n360) );
  MUX2_X1 U402 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n366), .Z(n361) );
  MUX2_X1 U403 ( .A(n361), .B(n360), .S(N11), .Z(n362) );
endmodule


module memory_WIDTH16_SIZE8_LOGSIZE3_5 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] ,
         \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][15] , \mem[6][14] , \mem[6][13] ,
         \mem[6][12] , \mem[6][11] , \mem[6][10] , \mem[6][9] , \mem[6][8] ,
         \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] ,
         \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[5][15] , \mem[5][14] ,
         \mem[5][13] , \mem[5][12] , \mem[5][11] , \mem[5][10] , \mem[5][9] ,
         \mem[5][8] , \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] ,
         \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][15] ,
         \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] , \mem[4][10] ,
         \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N13, N14, N15,
         N16, N17, N18, N19, N20, N21, N22, N23, N26, N28, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[15]  ( .D(N13), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N14), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(N15), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(N16), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N18), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N19), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N20), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N21), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N22), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N23), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[2]  ( .D(N26), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N28), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][15]  ( .D(n394), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n395), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n396), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n397), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n398), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n399), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n400), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n401), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n402), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n403), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n404), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n405), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n406), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n407), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n408), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n409), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n410), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n411), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n412), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n413), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n414), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n415), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n416), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n417), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n418), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n419), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n420), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n421), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n422), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n423), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n424), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n425), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n426), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n427), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n428), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n429), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n430), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n431), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n432), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n433), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n434), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n435), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n436), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n437), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n438), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n439), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n440), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n441), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n442), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n443), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n444), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n445), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n446), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n447), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n448), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n449), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n450), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n451), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n452), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n453), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n454), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n455), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n456), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n457), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n458), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n459), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n460), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n461), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n462), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n463), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n464), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n465), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n466), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n467), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n468), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n469), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n470), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n471), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n472), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n473), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n474), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n475), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n476), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n477), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n478), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n479), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n480), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n481), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n482), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n483), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n484), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n485), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n486), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n487), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n488), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n489), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n490), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n491), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n492), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n493), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n494), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n495), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n496), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n497), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n498), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n499), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n500), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n501), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n502), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n503), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n504), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n505), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n506), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n507), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n508), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n509), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n510), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n511), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n512), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n513), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n514), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n515), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n516), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n517), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n518), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n519), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n520), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n521), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U280 ( .A1(n375), .A2(n376), .A3(n642), .ZN(n659) );
  NAND3_X1 U281 ( .A1(n642), .A2(n376), .A3(N10), .ZN(n641) );
  NAND3_X1 U282 ( .A1(n642), .A2(n375), .A3(N11), .ZN(n624) );
  NAND3_X1 U283 ( .A1(N10), .A2(n642), .A3(N11), .ZN(n607) );
  NAND3_X1 U284 ( .A1(n375), .A2(n376), .A3(n573), .ZN(n590) );
  NAND3_X1 U285 ( .A1(N10), .A2(n376), .A3(n573), .ZN(n572) );
  NAND3_X1 U286 ( .A1(N11), .A2(n375), .A3(n573), .ZN(n555) );
  NAND3_X1 U287 ( .A1(N11), .A2(N10), .A3(n573), .ZN(n538) );
  DFF_X1 \data_out_reg[11]  ( .D(N17), .CK(clk), .Q(data_out[11]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n12), .SI(n9), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[4]  ( .D(n296), .SI(n293), .SE(N12), .CK(clk), .Q(
        data_out[4]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n290), .SI(n287), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  BUF_X1 U3 ( .A(n659), .Z(n374) );
  BUF_X1 U4 ( .A(n641), .Z(n373) );
  BUF_X1 U5 ( .A(n607), .Z(n371) );
  BUF_X1 U6 ( .A(n590), .Z(n370) );
  BUF_X1 U7 ( .A(n572), .Z(n369) );
  BUF_X1 U8 ( .A(n555), .Z(n368) );
  BUF_X1 U9 ( .A(n538), .Z(n367) );
  BUF_X1 U10 ( .A(n624), .Z(n372) );
  BUF_X1 U11 ( .A(N10), .Z(n365) );
  BUF_X1 U12 ( .A(N10), .Z(n366) );
  BUF_X1 U13 ( .A(N11), .Z(n363) );
  NOR2_X1 U14 ( .A1(n377), .A2(N12), .ZN(n642) );
  INV_X1 U15 ( .A(wr_en), .ZN(n377) );
  AND2_X1 U16 ( .A1(N12), .A2(wr_en), .ZN(n573) );
  OAI21_X1 U17 ( .B1(n386), .B2(n607), .A(n599), .ZN(n466) );
  NAND2_X1 U18 ( .A1(\mem[3][7] ), .A2(n371), .ZN(n599) );
  OAI21_X1 U19 ( .B1(n385), .B2(n371), .A(n598), .ZN(n465) );
  NAND2_X1 U20 ( .A1(\mem[3][8] ), .A2(n371), .ZN(n598) );
  OAI21_X1 U21 ( .B1(n384), .B2(n607), .A(n597), .ZN(n464) );
  NAND2_X1 U22 ( .A1(\mem[3][9] ), .A2(n371), .ZN(n597) );
  OAI21_X1 U23 ( .B1(n383), .B2(n607), .A(n596), .ZN(n463) );
  NAND2_X1 U24 ( .A1(\mem[3][10] ), .A2(n371), .ZN(n596) );
  OAI21_X1 U25 ( .B1(n382), .B2(n607), .A(n595), .ZN(n462) );
  NAND2_X1 U26 ( .A1(\mem[3][11] ), .A2(n371), .ZN(n595) );
  OAI21_X1 U27 ( .B1(n381), .B2(n607), .A(n594), .ZN(n461) );
  NAND2_X1 U28 ( .A1(\mem[3][12] ), .A2(n371), .ZN(n594) );
  OAI21_X1 U29 ( .B1(n380), .B2(n607), .A(n593), .ZN(n460) );
  NAND2_X1 U30 ( .A1(\mem[3][13] ), .A2(n371), .ZN(n593) );
  OAI21_X1 U31 ( .B1(n379), .B2(n607), .A(n592), .ZN(n459) );
  NAND2_X1 U32 ( .A1(\mem[3][14] ), .A2(n371), .ZN(n592) );
  OAI21_X1 U33 ( .B1(n386), .B2(n572), .A(n564), .ZN(n434) );
  NAND2_X1 U34 ( .A1(\mem[5][7] ), .A2(n369), .ZN(n564) );
  OAI21_X1 U35 ( .B1(n385), .B2(n369), .A(n563), .ZN(n433) );
  NAND2_X1 U36 ( .A1(\mem[5][8] ), .A2(n369), .ZN(n563) );
  OAI21_X1 U37 ( .B1(n384), .B2(n572), .A(n562), .ZN(n432) );
  NAND2_X1 U38 ( .A1(\mem[5][9] ), .A2(n369), .ZN(n562) );
  OAI21_X1 U39 ( .B1(n383), .B2(n572), .A(n561), .ZN(n431) );
  NAND2_X1 U40 ( .A1(\mem[5][10] ), .A2(n369), .ZN(n561) );
  OAI21_X1 U41 ( .B1(n382), .B2(n572), .A(n560), .ZN(n430) );
  NAND2_X1 U42 ( .A1(\mem[5][11] ), .A2(n369), .ZN(n560) );
  OAI21_X1 U43 ( .B1(n381), .B2(n572), .A(n559), .ZN(n429) );
  NAND2_X1 U44 ( .A1(\mem[5][12] ), .A2(n369), .ZN(n559) );
  OAI21_X1 U45 ( .B1(n380), .B2(n572), .A(n558), .ZN(n428) );
  NAND2_X1 U46 ( .A1(\mem[5][13] ), .A2(n369), .ZN(n558) );
  OAI21_X1 U47 ( .B1(n379), .B2(n572), .A(n557), .ZN(n427) );
  NAND2_X1 U48 ( .A1(\mem[5][14] ), .A2(n369), .ZN(n557) );
  OAI21_X1 U49 ( .B1(n386), .B2(n538), .A(n530), .ZN(n402) );
  NAND2_X1 U50 ( .A1(\mem[7][7] ), .A2(n367), .ZN(n530) );
  OAI21_X1 U51 ( .B1(n385), .B2(n538), .A(n529), .ZN(n401) );
  NAND2_X1 U52 ( .A1(\mem[7][8] ), .A2(n538), .ZN(n529) );
  OAI21_X1 U53 ( .B1(n384), .B2(n538), .A(n528), .ZN(n400) );
  NAND2_X1 U54 ( .A1(\mem[7][9] ), .A2(n538), .ZN(n528) );
  OAI21_X1 U55 ( .B1(n383), .B2(n538), .A(n527), .ZN(n399) );
  NAND2_X1 U56 ( .A1(\mem[7][10] ), .A2(n538), .ZN(n527) );
  OAI21_X1 U57 ( .B1(n382), .B2(n538), .A(n526), .ZN(n398) );
  NAND2_X1 U58 ( .A1(\mem[7][11] ), .A2(n538), .ZN(n526) );
  OAI21_X1 U59 ( .B1(n381), .B2(n538), .A(n525), .ZN(n397) );
  NAND2_X1 U60 ( .A1(\mem[7][12] ), .A2(n538), .ZN(n525) );
  OAI21_X1 U61 ( .B1(n380), .B2(n538), .A(n524), .ZN(n396) );
  NAND2_X1 U62 ( .A1(\mem[7][13] ), .A2(n538), .ZN(n524) );
  OAI21_X1 U63 ( .B1(n379), .B2(n538), .A(n523), .ZN(n395) );
  NAND2_X1 U64 ( .A1(\mem[7][14] ), .A2(n538), .ZN(n523) );
  OAI21_X1 U65 ( .B1(n386), .B2(n641), .A(n633), .ZN(n498) );
  NAND2_X1 U66 ( .A1(\mem[1][7] ), .A2(n373), .ZN(n633) );
  OAI21_X1 U67 ( .B1(n385), .B2(n373), .A(n632), .ZN(n497) );
  NAND2_X1 U68 ( .A1(\mem[1][8] ), .A2(n373), .ZN(n632) );
  OAI21_X1 U69 ( .B1(n384), .B2(n641), .A(n631), .ZN(n496) );
  NAND2_X1 U70 ( .A1(\mem[1][9] ), .A2(n373), .ZN(n631) );
  OAI21_X1 U71 ( .B1(n383), .B2(n641), .A(n630), .ZN(n495) );
  NAND2_X1 U72 ( .A1(\mem[1][10] ), .A2(n373), .ZN(n630) );
  OAI21_X1 U73 ( .B1(n382), .B2(n641), .A(n629), .ZN(n494) );
  NAND2_X1 U74 ( .A1(\mem[1][11] ), .A2(n373), .ZN(n629) );
  OAI21_X1 U75 ( .B1(n381), .B2(n641), .A(n628), .ZN(n493) );
  NAND2_X1 U76 ( .A1(\mem[1][12] ), .A2(n373), .ZN(n628) );
  OAI21_X1 U77 ( .B1(n380), .B2(n641), .A(n627), .ZN(n492) );
  NAND2_X1 U78 ( .A1(\mem[1][13] ), .A2(n373), .ZN(n627) );
  OAI21_X1 U79 ( .B1(n379), .B2(n641), .A(n626), .ZN(n491) );
  NAND2_X1 U80 ( .A1(\mem[1][14] ), .A2(n373), .ZN(n626) );
  OAI21_X1 U81 ( .B1(n386), .B2(n555), .A(n547), .ZN(n418) );
  NAND2_X1 U82 ( .A1(\mem[6][7] ), .A2(n368), .ZN(n547) );
  OAI21_X1 U83 ( .B1(n385), .B2(n368), .A(n546), .ZN(n417) );
  NAND2_X1 U84 ( .A1(\mem[6][8] ), .A2(n368), .ZN(n546) );
  OAI21_X1 U85 ( .B1(n384), .B2(n555), .A(n545), .ZN(n416) );
  NAND2_X1 U86 ( .A1(\mem[6][9] ), .A2(n368), .ZN(n545) );
  OAI21_X1 U87 ( .B1(n383), .B2(n555), .A(n544), .ZN(n415) );
  NAND2_X1 U88 ( .A1(\mem[6][10] ), .A2(n368), .ZN(n544) );
  OAI21_X1 U89 ( .B1(n382), .B2(n555), .A(n543), .ZN(n414) );
  NAND2_X1 U90 ( .A1(\mem[6][11] ), .A2(n368), .ZN(n543) );
  OAI21_X1 U91 ( .B1(n381), .B2(n555), .A(n542), .ZN(n413) );
  NAND2_X1 U92 ( .A1(\mem[6][12] ), .A2(n368), .ZN(n542) );
  OAI21_X1 U93 ( .B1(n380), .B2(n555), .A(n541), .ZN(n412) );
  NAND2_X1 U94 ( .A1(\mem[6][13] ), .A2(n368), .ZN(n541) );
  OAI21_X1 U95 ( .B1(n379), .B2(n555), .A(n540), .ZN(n411) );
  NAND2_X1 U96 ( .A1(\mem[6][14] ), .A2(n368), .ZN(n540) );
  OAI21_X1 U97 ( .B1(n386), .B2(n372), .A(n616), .ZN(n482) );
  NAND2_X1 U98 ( .A1(\mem[2][7] ), .A2(n372), .ZN(n616) );
  OAI21_X1 U99 ( .B1(n385), .B2(n372), .A(n615), .ZN(n481) );
  NAND2_X1 U100 ( .A1(\mem[2][8] ), .A2(n624), .ZN(n615) );
  OAI21_X1 U101 ( .B1(n384), .B2(n372), .A(n614), .ZN(n480) );
  NAND2_X1 U102 ( .A1(\mem[2][9] ), .A2(n624), .ZN(n614) );
  OAI21_X1 U103 ( .B1(n383), .B2(n372), .A(n613), .ZN(n479) );
  NAND2_X1 U104 ( .A1(\mem[2][10] ), .A2(n624), .ZN(n613) );
  OAI21_X1 U105 ( .B1(n382), .B2(n372), .A(n612), .ZN(n478) );
  NAND2_X1 U106 ( .A1(\mem[2][11] ), .A2(n624), .ZN(n612) );
  OAI21_X1 U107 ( .B1(n381), .B2(n372), .A(n611), .ZN(n477) );
  NAND2_X1 U108 ( .A1(\mem[2][12] ), .A2(n624), .ZN(n611) );
  OAI21_X1 U109 ( .B1(n380), .B2(n372), .A(n610), .ZN(n476) );
  NAND2_X1 U110 ( .A1(\mem[2][13] ), .A2(n624), .ZN(n610) );
  OAI21_X1 U111 ( .B1(n379), .B2(n372), .A(n609), .ZN(n475) );
  NAND2_X1 U112 ( .A1(\mem[2][14] ), .A2(n624), .ZN(n609) );
  OAI21_X1 U113 ( .B1(n386), .B2(n590), .A(n582), .ZN(n450) );
  NAND2_X1 U114 ( .A1(\mem[4][7] ), .A2(n370), .ZN(n582) );
  OAI21_X1 U115 ( .B1(n385), .B2(n370), .A(n581), .ZN(n449) );
  NAND2_X1 U116 ( .A1(\mem[4][8] ), .A2(n370), .ZN(n581) );
  OAI21_X1 U117 ( .B1(n384), .B2(n590), .A(n580), .ZN(n448) );
  NAND2_X1 U118 ( .A1(\mem[4][9] ), .A2(n370), .ZN(n580) );
  OAI21_X1 U119 ( .B1(n383), .B2(n590), .A(n579), .ZN(n447) );
  NAND2_X1 U120 ( .A1(\mem[4][10] ), .A2(n370), .ZN(n579) );
  OAI21_X1 U121 ( .B1(n382), .B2(n590), .A(n578), .ZN(n446) );
  NAND2_X1 U122 ( .A1(\mem[4][11] ), .A2(n370), .ZN(n578) );
  OAI21_X1 U123 ( .B1(n381), .B2(n590), .A(n577), .ZN(n445) );
  NAND2_X1 U124 ( .A1(\mem[4][12] ), .A2(n370), .ZN(n577) );
  OAI21_X1 U125 ( .B1(n380), .B2(n590), .A(n576), .ZN(n444) );
  NAND2_X1 U126 ( .A1(\mem[4][13] ), .A2(n370), .ZN(n576) );
  OAI21_X1 U127 ( .B1(n379), .B2(n590), .A(n575), .ZN(n443) );
  NAND2_X1 U128 ( .A1(\mem[4][14] ), .A2(n370), .ZN(n575) );
  OAI21_X1 U129 ( .B1(n659), .B2(n385), .A(n650), .ZN(n513) );
  NAND2_X1 U130 ( .A1(\mem[0][8] ), .A2(n374), .ZN(n650) );
  OAI21_X1 U131 ( .B1(n659), .B2(n384), .A(n649), .ZN(n512) );
  NAND2_X1 U132 ( .A1(\mem[0][9] ), .A2(n374), .ZN(n649) );
  OAI21_X1 U133 ( .B1(n659), .B2(n383), .A(n648), .ZN(n511) );
  NAND2_X1 U134 ( .A1(\mem[0][10] ), .A2(n374), .ZN(n648) );
  OAI21_X1 U135 ( .B1(n659), .B2(n382), .A(n647), .ZN(n510) );
  NAND2_X1 U136 ( .A1(\mem[0][11] ), .A2(n374), .ZN(n647) );
  OAI21_X1 U137 ( .B1(n659), .B2(n381), .A(n646), .ZN(n509) );
  NAND2_X1 U138 ( .A1(\mem[0][12] ), .A2(n374), .ZN(n646) );
  OAI21_X1 U139 ( .B1(n659), .B2(n380), .A(n645), .ZN(n508) );
  NAND2_X1 U140 ( .A1(\mem[0][13] ), .A2(n374), .ZN(n645) );
  OAI21_X1 U141 ( .B1(n659), .B2(n379), .A(n644), .ZN(n507) );
  NAND2_X1 U142 ( .A1(\mem[0][14] ), .A2(n374), .ZN(n644) );
  INV_X1 U143 ( .A(N10), .ZN(n375) );
  OAI21_X1 U144 ( .B1(n393), .B2(n641), .A(n640), .ZN(n505) );
  NAND2_X1 U145 ( .A1(\mem[1][0] ), .A2(n373), .ZN(n640) );
  OAI21_X1 U146 ( .B1(n392), .B2(n641), .A(n639), .ZN(n504) );
  NAND2_X1 U147 ( .A1(\mem[1][1] ), .A2(n373), .ZN(n639) );
  OAI21_X1 U148 ( .B1(n391), .B2(n641), .A(n638), .ZN(n503) );
  NAND2_X1 U149 ( .A1(\mem[1][2] ), .A2(n373), .ZN(n638) );
  OAI21_X1 U150 ( .B1(n390), .B2(n641), .A(n637), .ZN(n502) );
  NAND2_X1 U151 ( .A1(\mem[1][3] ), .A2(n373), .ZN(n637) );
  OAI21_X1 U152 ( .B1(n389), .B2(n641), .A(n636), .ZN(n501) );
  NAND2_X1 U153 ( .A1(\mem[1][4] ), .A2(n641), .ZN(n636) );
  OAI21_X1 U154 ( .B1(n388), .B2(n641), .A(n635), .ZN(n500) );
  NAND2_X1 U155 ( .A1(\mem[1][5] ), .A2(n641), .ZN(n635) );
  OAI21_X1 U156 ( .B1(n387), .B2(n641), .A(n634), .ZN(n499) );
  NAND2_X1 U157 ( .A1(\mem[1][6] ), .A2(n641), .ZN(n634) );
  OAI21_X1 U158 ( .B1(n378), .B2(n641), .A(n625), .ZN(n490) );
  NAND2_X1 U159 ( .A1(\mem[1][15] ), .A2(n373), .ZN(n625) );
  OAI21_X1 U160 ( .B1(n393), .B2(n372), .A(n623), .ZN(n489) );
  NAND2_X1 U161 ( .A1(\mem[2][0] ), .A2(n372), .ZN(n623) );
  OAI21_X1 U162 ( .B1(n392), .B2(n624), .A(n622), .ZN(n488) );
  NAND2_X1 U163 ( .A1(\mem[2][1] ), .A2(n624), .ZN(n622) );
  OAI21_X1 U164 ( .B1(n391), .B2(n372), .A(n621), .ZN(n487) );
  NAND2_X1 U165 ( .A1(\mem[2][2] ), .A2(n624), .ZN(n621) );
  OAI21_X1 U166 ( .B1(n390), .B2(n624), .A(n620), .ZN(n486) );
  NAND2_X1 U167 ( .A1(\mem[2][3] ), .A2(n624), .ZN(n620) );
  OAI21_X1 U168 ( .B1(n389), .B2(n624), .A(n619), .ZN(n485) );
  NAND2_X1 U169 ( .A1(\mem[2][4] ), .A2(n372), .ZN(n619) );
  OAI21_X1 U170 ( .B1(n388), .B2(n624), .A(n618), .ZN(n484) );
  NAND2_X1 U171 ( .A1(\mem[2][5] ), .A2(n372), .ZN(n618) );
  OAI21_X1 U172 ( .B1(n387), .B2(n624), .A(n617), .ZN(n483) );
  NAND2_X1 U173 ( .A1(\mem[2][6] ), .A2(n372), .ZN(n617) );
  OAI21_X1 U174 ( .B1(n378), .B2(n624), .A(n608), .ZN(n474) );
  NAND2_X1 U175 ( .A1(\mem[2][15] ), .A2(n624), .ZN(n608) );
  OAI21_X1 U176 ( .B1(n393), .B2(n607), .A(n606), .ZN(n473) );
  NAND2_X1 U177 ( .A1(\mem[3][0] ), .A2(n371), .ZN(n606) );
  OAI21_X1 U178 ( .B1(n392), .B2(n607), .A(n605), .ZN(n472) );
  NAND2_X1 U179 ( .A1(\mem[3][1] ), .A2(n371), .ZN(n605) );
  OAI21_X1 U180 ( .B1(n391), .B2(n607), .A(n604), .ZN(n471) );
  NAND2_X1 U181 ( .A1(\mem[3][2] ), .A2(n371), .ZN(n604) );
  OAI21_X1 U182 ( .B1(n390), .B2(n607), .A(n603), .ZN(n470) );
  NAND2_X1 U183 ( .A1(\mem[3][3] ), .A2(n371), .ZN(n603) );
  OAI21_X1 U184 ( .B1(n389), .B2(n607), .A(n602), .ZN(n469) );
  NAND2_X1 U185 ( .A1(\mem[3][4] ), .A2(n607), .ZN(n602) );
  OAI21_X1 U186 ( .B1(n388), .B2(n607), .A(n601), .ZN(n468) );
  NAND2_X1 U187 ( .A1(\mem[3][5] ), .A2(n607), .ZN(n601) );
  OAI21_X1 U188 ( .B1(n387), .B2(n607), .A(n600), .ZN(n467) );
  NAND2_X1 U189 ( .A1(\mem[3][6] ), .A2(n607), .ZN(n600) );
  OAI21_X1 U190 ( .B1(n378), .B2(n607), .A(n591), .ZN(n458) );
  NAND2_X1 U191 ( .A1(\mem[3][15] ), .A2(n371), .ZN(n591) );
  OAI21_X1 U192 ( .B1(n393), .B2(n590), .A(n589), .ZN(n457) );
  NAND2_X1 U193 ( .A1(\mem[4][0] ), .A2(n370), .ZN(n589) );
  OAI21_X1 U194 ( .B1(n392), .B2(n590), .A(n588), .ZN(n456) );
  NAND2_X1 U195 ( .A1(\mem[4][1] ), .A2(n370), .ZN(n588) );
  OAI21_X1 U196 ( .B1(n391), .B2(n590), .A(n587), .ZN(n455) );
  NAND2_X1 U197 ( .A1(\mem[4][2] ), .A2(n370), .ZN(n587) );
  OAI21_X1 U198 ( .B1(n390), .B2(n590), .A(n586), .ZN(n454) );
  NAND2_X1 U199 ( .A1(\mem[4][3] ), .A2(n370), .ZN(n586) );
  OAI21_X1 U200 ( .B1(n389), .B2(n590), .A(n585), .ZN(n453) );
  NAND2_X1 U201 ( .A1(\mem[4][4] ), .A2(n590), .ZN(n585) );
  OAI21_X1 U202 ( .B1(n388), .B2(n590), .A(n584), .ZN(n452) );
  NAND2_X1 U203 ( .A1(\mem[4][5] ), .A2(n590), .ZN(n584) );
  OAI21_X1 U204 ( .B1(n387), .B2(n590), .A(n583), .ZN(n451) );
  NAND2_X1 U205 ( .A1(\mem[4][6] ), .A2(n590), .ZN(n583) );
  OAI21_X1 U206 ( .B1(n378), .B2(n590), .A(n574), .ZN(n442) );
  NAND2_X1 U207 ( .A1(\mem[4][15] ), .A2(n370), .ZN(n574) );
  OAI21_X1 U208 ( .B1(n393), .B2(n572), .A(n571), .ZN(n441) );
  NAND2_X1 U209 ( .A1(\mem[5][0] ), .A2(n369), .ZN(n571) );
  OAI21_X1 U210 ( .B1(n392), .B2(n572), .A(n570), .ZN(n440) );
  NAND2_X1 U211 ( .A1(\mem[5][1] ), .A2(n369), .ZN(n570) );
  OAI21_X1 U212 ( .B1(n391), .B2(n572), .A(n569), .ZN(n439) );
  NAND2_X1 U213 ( .A1(\mem[5][2] ), .A2(n369), .ZN(n569) );
  OAI21_X1 U214 ( .B1(n390), .B2(n572), .A(n568), .ZN(n438) );
  NAND2_X1 U215 ( .A1(\mem[5][3] ), .A2(n369), .ZN(n568) );
  OAI21_X1 U216 ( .B1(n389), .B2(n572), .A(n567), .ZN(n437) );
  NAND2_X1 U217 ( .A1(\mem[5][4] ), .A2(n572), .ZN(n567) );
  OAI21_X1 U218 ( .B1(n388), .B2(n572), .A(n566), .ZN(n436) );
  NAND2_X1 U219 ( .A1(\mem[5][5] ), .A2(n572), .ZN(n566) );
  OAI21_X1 U220 ( .B1(n387), .B2(n572), .A(n565), .ZN(n435) );
  NAND2_X1 U221 ( .A1(\mem[5][6] ), .A2(n572), .ZN(n565) );
  OAI21_X1 U222 ( .B1(n378), .B2(n572), .A(n556), .ZN(n426) );
  NAND2_X1 U223 ( .A1(\mem[5][15] ), .A2(n369), .ZN(n556) );
  OAI21_X1 U224 ( .B1(n393), .B2(n555), .A(n554), .ZN(n425) );
  NAND2_X1 U225 ( .A1(\mem[6][0] ), .A2(n368), .ZN(n554) );
  OAI21_X1 U226 ( .B1(n392), .B2(n555), .A(n553), .ZN(n424) );
  NAND2_X1 U227 ( .A1(\mem[6][1] ), .A2(n368), .ZN(n553) );
  OAI21_X1 U228 ( .B1(n391), .B2(n555), .A(n552), .ZN(n423) );
  NAND2_X1 U229 ( .A1(\mem[6][2] ), .A2(n368), .ZN(n552) );
  OAI21_X1 U230 ( .B1(n390), .B2(n555), .A(n551), .ZN(n422) );
  NAND2_X1 U231 ( .A1(\mem[6][3] ), .A2(n368), .ZN(n551) );
  OAI21_X1 U232 ( .B1(n389), .B2(n555), .A(n550), .ZN(n421) );
  NAND2_X1 U233 ( .A1(\mem[6][4] ), .A2(n555), .ZN(n550) );
  OAI21_X1 U234 ( .B1(n388), .B2(n555), .A(n549), .ZN(n420) );
  NAND2_X1 U235 ( .A1(\mem[6][5] ), .A2(n555), .ZN(n549) );
  OAI21_X1 U236 ( .B1(n387), .B2(n555), .A(n548), .ZN(n419) );
  NAND2_X1 U237 ( .A1(\mem[6][6] ), .A2(n555), .ZN(n548) );
  OAI21_X1 U238 ( .B1(n378), .B2(n555), .A(n539), .ZN(n410) );
  NAND2_X1 U239 ( .A1(\mem[6][15] ), .A2(n368), .ZN(n539) );
  OAI21_X1 U240 ( .B1(n393), .B2(n367), .A(n537), .ZN(n409) );
  NAND2_X1 U241 ( .A1(\mem[7][0] ), .A2(n367), .ZN(n537) );
  OAI21_X1 U242 ( .B1(n392), .B2(n367), .A(n536), .ZN(n408) );
  NAND2_X1 U243 ( .A1(\mem[7][1] ), .A2(n538), .ZN(n536) );
  OAI21_X1 U244 ( .B1(n391), .B2(n367), .A(n535), .ZN(n407) );
  NAND2_X1 U245 ( .A1(\mem[7][2] ), .A2(n538), .ZN(n535) );
  OAI21_X1 U246 ( .B1(n390), .B2(n367), .A(n534), .ZN(n406) );
  NAND2_X1 U247 ( .A1(\mem[7][3] ), .A2(n538), .ZN(n534) );
  OAI21_X1 U248 ( .B1(n389), .B2(n367), .A(n533), .ZN(n405) );
  NAND2_X1 U249 ( .A1(\mem[7][4] ), .A2(n367), .ZN(n533) );
  OAI21_X1 U250 ( .B1(n388), .B2(n367), .A(n532), .ZN(n404) );
  NAND2_X1 U251 ( .A1(\mem[7][5] ), .A2(n367), .ZN(n532) );
  OAI21_X1 U252 ( .B1(n387), .B2(n367), .A(n531), .ZN(n403) );
  NAND2_X1 U253 ( .A1(\mem[7][6] ), .A2(n367), .ZN(n531) );
  OAI21_X1 U254 ( .B1(n378), .B2(n367), .A(n522), .ZN(n394) );
  NAND2_X1 U255 ( .A1(\mem[7][15] ), .A2(n367), .ZN(n522) );
  OAI21_X1 U256 ( .B1(n659), .B2(n393), .A(n658), .ZN(n521) );
  NAND2_X1 U257 ( .A1(\mem[0][0] ), .A2(n374), .ZN(n658) );
  OAI21_X1 U258 ( .B1(n374), .B2(n392), .A(n657), .ZN(n520) );
  NAND2_X1 U259 ( .A1(\mem[0][1] ), .A2(n374), .ZN(n657) );
  OAI21_X1 U260 ( .B1(n659), .B2(n391), .A(n656), .ZN(n519) );
  NAND2_X1 U261 ( .A1(\mem[0][2] ), .A2(n374), .ZN(n656) );
  OAI21_X1 U262 ( .B1(n659), .B2(n390), .A(n655), .ZN(n518) );
  NAND2_X1 U263 ( .A1(\mem[0][3] ), .A2(n374), .ZN(n655) );
  OAI21_X1 U264 ( .B1(n659), .B2(n389), .A(n654), .ZN(n517) );
  NAND2_X1 U265 ( .A1(\mem[0][4] ), .A2(n374), .ZN(n654) );
  OAI21_X1 U266 ( .B1(n659), .B2(n388), .A(n653), .ZN(n516) );
  NAND2_X1 U267 ( .A1(\mem[0][5] ), .A2(n659), .ZN(n653) );
  OAI21_X1 U268 ( .B1(n659), .B2(n387), .A(n652), .ZN(n515) );
  NAND2_X1 U269 ( .A1(\mem[0][6] ), .A2(n659), .ZN(n652) );
  OAI21_X1 U270 ( .B1(n659), .B2(n386), .A(n651), .ZN(n514) );
  NAND2_X1 U271 ( .A1(\mem[0][7] ), .A2(n659), .ZN(n651) );
  OAI21_X1 U272 ( .B1(n659), .B2(n378), .A(n643), .ZN(n506) );
  NAND2_X1 U273 ( .A1(\mem[0][15] ), .A2(n374), .ZN(n643) );
  INV_X1 U274 ( .A(N11), .ZN(n376) );
  INV_X1 U275 ( .A(data_in[0]), .ZN(n393) );
  INV_X1 U276 ( .A(data_in[1]), .ZN(n392) );
  INV_X1 U277 ( .A(data_in[2]), .ZN(n391) );
  INV_X1 U278 ( .A(data_in[3]), .ZN(n390) );
  INV_X1 U279 ( .A(data_in[4]), .ZN(n389) );
  INV_X1 U288 ( .A(data_in[5]), .ZN(n388) );
  INV_X1 U289 ( .A(data_in[6]), .ZN(n387) );
  INV_X1 U290 ( .A(data_in[7]), .ZN(n386) );
  INV_X1 U291 ( .A(data_in[8]), .ZN(n385) );
  INV_X1 U292 ( .A(data_in[9]), .ZN(n384) );
  INV_X1 U293 ( .A(data_in[10]), .ZN(n383) );
  INV_X1 U294 ( .A(data_in[11]), .ZN(n382) );
  INV_X1 U295 ( .A(data_in[12]), .ZN(n381) );
  INV_X1 U296 ( .A(data_in[13]), .ZN(n380) );
  INV_X1 U297 ( .A(data_in[14]), .ZN(n379) );
  INV_X1 U298 ( .A(data_in[15]), .ZN(n378) );
  MUX2_X1 U299 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n364), .Z(n1) );
  MUX2_X1 U300 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n364), .Z(n2) );
  MUX2_X1 U301 ( .A(n2), .B(n1), .S(n363), .Z(n3) );
  MUX2_X1 U302 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n364), .Z(n4) );
  MUX2_X1 U303 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n364), .Z(n5) );
  MUX2_X1 U304 ( .A(n5), .B(n4), .S(N11), .Z(n6) );
  MUX2_X1 U305 ( .A(n6), .B(n3), .S(N12), .Z(N28) );
  MUX2_X1 U306 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n364), .Z(n7) );
  MUX2_X1 U307 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n364), .Z(n8) );
  MUX2_X1 U308 ( .A(n8), .B(n7), .S(N11), .Z(n9) );
  MUX2_X1 U309 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n366), .Z(n10) );
  MUX2_X1 U310 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(N10), .Z(n11) );
  MUX2_X1 U311 ( .A(n11), .B(n10), .S(N11), .Z(n12) );
  MUX2_X1 U312 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n364), .Z(n13) );
  MUX2_X1 U313 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n364), .Z(n14) );
  MUX2_X1 U314 ( .A(n14), .B(n13), .S(N11), .Z(n15) );
  MUX2_X1 U315 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n364), .Z(n16) );
  MUX2_X1 U316 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n364), .Z(n17) );
  MUX2_X1 U317 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U318 ( .A(n18), .B(n15), .S(N12), .Z(N26) );
  MUX2_X1 U319 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n364), .Z(n19) );
  MUX2_X1 U320 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n365), .Z(n286) );
  MUX2_X1 U321 ( .A(n286), .B(n19), .S(N11), .Z(n287) );
  MUX2_X1 U322 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n288) );
  MUX2_X1 U323 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n364), .Z(n289) );
  MUX2_X1 U324 ( .A(n289), .B(n288), .S(N11), .Z(n290) );
  MUX2_X1 U325 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n365), .Z(n291) );
  MUX2_X1 U326 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n365), .Z(n292) );
  MUX2_X1 U327 ( .A(n292), .B(n291), .S(n363), .Z(n293) );
  MUX2_X1 U328 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n365), .Z(n294) );
  MUX2_X1 U329 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n365), .Z(n295) );
  MUX2_X1 U330 ( .A(n295), .B(n294), .S(n363), .Z(n296) );
  MUX2_X1 U331 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n365), .Z(n297) );
  MUX2_X1 U332 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n365), .Z(n298) );
  MUX2_X1 U333 ( .A(n298), .B(n297), .S(n363), .Z(n299) );
  MUX2_X1 U334 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n365), .Z(n300) );
  MUX2_X1 U335 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n365), .Z(n301) );
  MUX2_X1 U336 ( .A(n301), .B(n300), .S(n363), .Z(n302) );
  MUX2_X1 U337 ( .A(n302), .B(n299), .S(N12), .Z(N23) );
  MUX2_X1 U338 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n365), .Z(n303) );
  MUX2_X1 U339 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n365), .Z(n304) );
  MUX2_X1 U340 ( .A(n304), .B(n303), .S(n363), .Z(n305) );
  MUX2_X1 U341 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n365), .Z(n306) );
  MUX2_X1 U342 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n365), .Z(n307) );
  MUX2_X1 U343 ( .A(n307), .B(n306), .S(n363), .Z(n308) );
  MUX2_X1 U344 ( .A(n308), .B(n305), .S(N12), .Z(N22) );
  MUX2_X1 U345 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n366), .Z(n309) );
  MUX2_X1 U346 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n366), .Z(n310) );
  MUX2_X1 U347 ( .A(n310), .B(n309), .S(n363), .Z(n311) );
  MUX2_X1 U348 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n366), .Z(n312) );
  MUX2_X1 U349 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n366), .Z(n313) );
  MUX2_X1 U350 ( .A(n313), .B(n312), .S(n363), .Z(n314) );
  MUX2_X1 U351 ( .A(n314), .B(n311), .S(N12), .Z(N21) );
  MUX2_X1 U352 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n366), .Z(n315) );
  MUX2_X1 U353 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n366), .Z(n316) );
  MUX2_X1 U354 ( .A(n316), .B(n315), .S(n363), .Z(n317) );
  MUX2_X1 U355 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n366), .Z(n318) );
  MUX2_X1 U356 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n366), .Z(n319) );
  MUX2_X1 U357 ( .A(n319), .B(n318), .S(n363), .Z(n320) );
  MUX2_X1 U358 ( .A(n320), .B(n317), .S(N12), .Z(N20) );
  MUX2_X1 U359 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n366), .Z(n321) );
  MUX2_X1 U360 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n366), .Z(n322) );
  MUX2_X1 U361 ( .A(n322), .B(n321), .S(n363), .Z(n323) );
  MUX2_X1 U362 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n366), .Z(n324) );
  MUX2_X1 U363 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n366), .Z(n325) );
  MUX2_X1 U364 ( .A(n325), .B(n324), .S(n363), .Z(n326) );
  MUX2_X1 U365 ( .A(n326), .B(n323), .S(N12), .Z(N19) );
  MUX2_X1 U366 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n364), .Z(n327) );
  MUX2_X1 U367 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n366), .Z(n328) );
  MUX2_X1 U368 ( .A(n328), .B(n327), .S(n363), .Z(n329) );
  MUX2_X1 U369 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n364), .Z(n330) );
  MUX2_X1 U370 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n366), .Z(n331) );
  MUX2_X1 U371 ( .A(n331), .B(n330), .S(N11), .Z(n332) );
  MUX2_X1 U372 ( .A(n332), .B(n329), .S(N12), .Z(N18) );
  MUX2_X1 U373 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n365), .Z(n333) );
  MUX2_X1 U374 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n364), .Z(n334) );
  MUX2_X1 U375 ( .A(n334), .B(n333), .S(n363), .Z(n335) );
  MUX2_X1 U376 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n365), .Z(n336) );
  MUX2_X1 U377 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n364), .Z(n337) );
  MUX2_X1 U378 ( .A(n337), .B(n336), .S(N11), .Z(n338) );
  MUX2_X1 U379 ( .A(n338), .B(n335), .S(N12), .Z(N17) );
  MUX2_X1 U380 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n365), .Z(n339) );
  MUX2_X1 U381 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n365), .Z(n340) );
  MUX2_X1 U382 ( .A(n340), .B(n339), .S(N11), .Z(n341) );
  MUX2_X1 U383 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n366), .Z(n342) );
  MUX2_X1 U384 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n365), .Z(n343) );
  MUX2_X1 U385 ( .A(n343), .B(n342), .S(N11), .Z(n344) );
  MUX2_X1 U386 ( .A(n344), .B(n341), .S(N12), .Z(N16) );
  MUX2_X1 U387 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n366), .Z(n345) );
  MUX2_X1 U388 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n366), .Z(n346) );
  MUX2_X1 U389 ( .A(n346), .B(n345), .S(N11), .Z(n347) );
  MUX2_X1 U390 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n364), .Z(n348) );
  MUX2_X1 U391 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n365), .Z(n349) );
  MUX2_X1 U392 ( .A(n349), .B(n348), .S(N11), .Z(n350) );
  MUX2_X1 U393 ( .A(n350), .B(n347), .S(N12), .Z(N15) );
  MUX2_X1 U394 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n365), .Z(n351) );
  MUX2_X1 U395 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n364), .Z(n352) );
  MUX2_X1 U396 ( .A(n352), .B(n351), .S(N11), .Z(n353) );
  MUX2_X1 U397 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n364), .Z(n354) );
  MUX2_X1 U398 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n366), .Z(n355) );
  MUX2_X1 U399 ( .A(n355), .B(n354), .S(N11), .Z(n356) );
  MUX2_X1 U400 ( .A(n356), .B(n353), .S(N12), .Z(N14) );
  MUX2_X1 U401 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n366), .Z(n357) );
  MUX2_X1 U402 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n366), .Z(n358) );
  MUX2_X1 U403 ( .A(n358), .B(n357), .S(N11), .Z(n359) );
  MUX2_X1 U404 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n365), .Z(n360) );
  MUX2_X1 U405 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n364), .Z(n361) );
  MUX2_X1 U406 ( .A(n361), .B(n360), .S(N11), .Z(n362) );
  MUX2_X1 U407 ( .A(n362), .B(n359), .S(N12), .Z(N13) );
  CLKBUF_X1 U408 ( .A(N10), .Z(n364) );
endmodule


module memory_WIDTH16_SIZE8_LOGSIZE3_4 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] ,
         \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][15] , \mem[6][14] , \mem[6][13] ,
         \mem[6][12] , \mem[6][11] , \mem[6][10] , \mem[6][9] , \mem[6][8] ,
         \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] ,
         \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[5][15] , \mem[5][14] ,
         \mem[5][13] , \mem[5][12] , \mem[5][11] , \mem[5][10] , \mem[5][9] ,
         \mem[5][8] , \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] ,
         \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][15] ,
         \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] , \mem[4][10] ,
         \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14, N16, N18,
         N19, N20, N22, N24, N26, N27, N28, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[14]  ( .D(N14), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N16), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N18), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N19), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N20), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N22), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N24), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N26), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N27), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N28), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][15]  ( .D(n394), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n395), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n396), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n397), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n398), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n399), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n400), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n401), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n402), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n403), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n404), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n405), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n406), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n407), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n408), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n409), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n410), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n411), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n412), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n413), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n414), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n415), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n416), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n417), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n418), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n419), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n420), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n421), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n422), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n423), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n424), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n425), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n426), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n427), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n428), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n429), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n430), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n431), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n432), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n433), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n434), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n435), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n436), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n437), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n438), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n439), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n440), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n441), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n442), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n443), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n444), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n445), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n446), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n447), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n448), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n449), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n450), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n451), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n452), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n453), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n454), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n455), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n456), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n457), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n458), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n459), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n460), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n461), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n462), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n463), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n464), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n465), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n466), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n467), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n468), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n469), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n470), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n471), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n472), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n473), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n474), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n475), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n476), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n477), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n478), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n479), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n480), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n481), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n482), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n483), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n484), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n485), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n486), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n487), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n488), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n489), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n490), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n491), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n492), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n493), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n494), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n495), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n496), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n497), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n498), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n499), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n500), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n501), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n502), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n503), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n504), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n505), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n506), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n507), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n508), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n509), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n510), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n511), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n512), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n513), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n514), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n515), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n516), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n517), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n518), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n519), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n520), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n521), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U280 ( .A1(n375), .A2(n376), .A3(n642), .ZN(n659) );
  NAND3_X1 U281 ( .A1(n642), .A2(n376), .A3(N10), .ZN(n641) );
  NAND3_X1 U282 ( .A1(n642), .A2(n375), .A3(N11), .ZN(n624) );
  NAND3_X1 U283 ( .A1(N10), .A2(n642), .A3(N11), .ZN(n607) );
  NAND3_X1 U284 ( .A1(n375), .A2(n376), .A3(n573), .ZN(n590) );
  NAND3_X1 U285 ( .A1(N10), .A2(n376), .A3(n573), .ZN(n572) );
  NAND3_X1 U286 ( .A1(N11), .A2(n375), .A3(n573), .ZN(n555) );
  NAND3_X1 U287 ( .A1(N11), .A2(N10), .A3(n573), .ZN(n538) );
  SDFF_X1 \data_out_reg[11]  ( .D(n338), .SI(n335), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n302), .SI(n299), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n314), .SI(n311), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n290), .SI(n287), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n362), .SI(n359), .SE(N12), .CK(clk), .Q(
        data_out[15]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n350), .SI(n347), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  BUF_X1 U3 ( .A(N10), .Z(n365) );
  BUF_X1 U4 ( .A(N10), .Z(n366) );
  BUF_X1 U5 ( .A(n659), .Z(n374) );
  BUF_X1 U6 ( .A(n641), .Z(n373) );
  BUF_X1 U7 ( .A(n624), .Z(n372) );
  BUF_X1 U8 ( .A(n590), .Z(n370) );
  BUF_X1 U9 ( .A(n572), .Z(n369) );
  BUF_X1 U10 ( .A(n555), .Z(n368) );
  BUF_X1 U11 ( .A(n538), .Z(n367) );
  BUF_X1 U12 ( .A(n607), .Z(n371) );
  BUF_X1 U13 ( .A(N10), .Z(n364) );
  BUF_X1 U14 ( .A(N11), .Z(n363) );
  NOR2_X1 U15 ( .A1(n377), .A2(N12), .ZN(n642) );
  INV_X1 U16 ( .A(wr_en), .ZN(n377) );
  AND2_X1 U17 ( .A1(N12), .A2(wr_en), .ZN(n573) );
  OAI21_X1 U18 ( .B1(n386), .B2(n607), .A(n599), .ZN(n466) );
  NAND2_X1 U19 ( .A1(\mem[3][7] ), .A2(n371), .ZN(n599) );
  OAI21_X1 U20 ( .B1(n385), .B2(n607), .A(n598), .ZN(n465) );
  NAND2_X1 U21 ( .A1(\mem[3][8] ), .A2(n607), .ZN(n598) );
  OAI21_X1 U22 ( .B1(n384), .B2(n607), .A(n597), .ZN(n464) );
  NAND2_X1 U23 ( .A1(\mem[3][9] ), .A2(n607), .ZN(n597) );
  OAI21_X1 U24 ( .B1(n383), .B2(n607), .A(n596), .ZN(n463) );
  NAND2_X1 U25 ( .A1(\mem[3][10] ), .A2(n607), .ZN(n596) );
  OAI21_X1 U26 ( .B1(n382), .B2(n607), .A(n595), .ZN(n462) );
  NAND2_X1 U27 ( .A1(\mem[3][11] ), .A2(n607), .ZN(n595) );
  OAI21_X1 U28 ( .B1(n381), .B2(n607), .A(n594), .ZN(n461) );
  NAND2_X1 U29 ( .A1(\mem[3][12] ), .A2(n607), .ZN(n594) );
  OAI21_X1 U30 ( .B1(n380), .B2(n607), .A(n593), .ZN(n460) );
  NAND2_X1 U31 ( .A1(\mem[3][13] ), .A2(n607), .ZN(n593) );
  OAI21_X1 U32 ( .B1(n379), .B2(n607), .A(n592), .ZN(n459) );
  NAND2_X1 U33 ( .A1(\mem[3][14] ), .A2(n607), .ZN(n592) );
  OAI21_X1 U34 ( .B1(n386), .B2(n572), .A(n564), .ZN(n434) );
  NAND2_X1 U35 ( .A1(\mem[5][7] ), .A2(n369), .ZN(n564) );
  OAI21_X1 U36 ( .B1(n385), .B2(n369), .A(n563), .ZN(n433) );
  NAND2_X1 U37 ( .A1(\mem[5][8] ), .A2(n369), .ZN(n563) );
  OAI21_X1 U38 ( .B1(n384), .B2(n572), .A(n562), .ZN(n432) );
  NAND2_X1 U39 ( .A1(\mem[5][9] ), .A2(n369), .ZN(n562) );
  OAI21_X1 U40 ( .B1(n383), .B2(n572), .A(n561), .ZN(n431) );
  NAND2_X1 U41 ( .A1(\mem[5][10] ), .A2(n369), .ZN(n561) );
  OAI21_X1 U42 ( .B1(n382), .B2(n572), .A(n560), .ZN(n430) );
  NAND2_X1 U43 ( .A1(\mem[5][11] ), .A2(n369), .ZN(n560) );
  OAI21_X1 U44 ( .B1(n381), .B2(n572), .A(n559), .ZN(n429) );
  NAND2_X1 U45 ( .A1(\mem[5][12] ), .A2(n369), .ZN(n559) );
  OAI21_X1 U46 ( .B1(n380), .B2(n572), .A(n558), .ZN(n428) );
  NAND2_X1 U47 ( .A1(\mem[5][13] ), .A2(n369), .ZN(n558) );
  OAI21_X1 U48 ( .B1(n379), .B2(n572), .A(n557), .ZN(n427) );
  NAND2_X1 U49 ( .A1(\mem[5][14] ), .A2(n369), .ZN(n557) );
  OAI21_X1 U50 ( .B1(n386), .B2(n538), .A(n530), .ZN(n402) );
  NAND2_X1 U51 ( .A1(\mem[7][7] ), .A2(n367), .ZN(n530) );
  OAI21_X1 U52 ( .B1(n385), .B2(n367), .A(n529), .ZN(n401) );
  NAND2_X1 U53 ( .A1(\mem[7][8] ), .A2(n367), .ZN(n529) );
  OAI21_X1 U54 ( .B1(n384), .B2(n538), .A(n528), .ZN(n400) );
  NAND2_X1 U55 ( .A1(\mem[7][9] ), .A2(n367), .ZN(n528) );
  OAI21_X1 U56 ( .B1(n383), .B2(n538), .A(n527), .ZN(n399) );
  NAND2_X1 U57 ( .A1(\mem[7][10] ), .A2(n367), .ZN(n527) );
  OAI21_X1 U58 ( .B1(n382), .B2(n538), .A(n526), .ZN(n398) );
  NAND2_X1 U59 ( .A1(\mem[7][11] ), .A2(n367), .ZN(n526) );
  OAI21_X1 U60 ( .B1(n381), .B2(n538), .A(n525), .ZN(n397) );
  NAND2_X1 U61 ( .A1(\mem[7][12] ), .A2(n367), .ZN(n525) );
  OAI21_X1 U62 ( .B1(n380), .B2(n538), .A(n524), .ZN(n396) );
  NAND2_X1 U63 ( .A1(\mem[7][13] ), .A2(n367), .ZN(n524) );
  OAI21_X1 U64 ( .B1(n379), .B2(n538), .A(n523), .ZN(n395) );
  NAND2_X1 U65 ( .A1(\mem[7][14] ), .A2(n367), .ZN(n523) );
  OAI21_X1 U66 ( .B1(n386), .B2(n641), .A(n633), .ZN(n498) );
  NAND2_X1 U67 ( .A1(\mem[1][7] ), .A2(n373), .ZN(n633) );
  OAI21_X1 U68 ( .B1(n385), .B2(n373), .A(n632), .ZN(n497) );
  NAND2_X1 U69 ( .A1(\mem[1][8] ), .A2(n373), .ZN(n632) );
  OAI21_X1 U70 ( .B1(n384), .B2(n641), .A(n631), .ZN(n496) );
  NAND2_X1 U71 ( .A1(\mem[1][9] ), .A2(n373), .ZN(n631) );
  OAI21_X1 U72 ( .B1(n383), .B2(n641), .A(n630), .ZN(n495) );
  NAND2_X1 U73 ( .A1(\mem[1][10] ), .A2(n373), .ZN(n630) );
  OAI21_X1 U74 ( .B1(n382), .B2(n641), .A(n629), .ZN(n494) );
  NAND2_X1 U75 ( .A1(\mem[1][11] ), .A2(n373), .ZN(n629) );
  OAI21_X1 U76 ( .B1(n381), .B2(n641), .A(n628), .ZN(n493) );
  NAND2_X1 U77 ( .A1(\mem[1][12] ), .A2(n373), .ZN(n628) );
  OAI21_X1 U78 ( .B1(n380), .B2(n641), .A(n627), .ZN(n492) );
  NAND2_X1 U79 ( .A1(\mem[1][13] ), .A2(n373), .ZN(n627) );
  OAI21_X1 U80 ( .B1(n379), .B2(n641), .A(n626), .ZN(n491) );
  NAND2_X1 U81 ( .A1(\mem[1][14] ), .A2(n373), .ZN(n626) );
  OAI21_X1 U82 ( .B1(n386), .B2(n555), .A(n547), .ZN(n418) );
  NAND2_X1 U83 ( .A1(\mem[6][7] ), .A2(n368), .ZN(n547) );
  OAI21_X1 U84 ( .B1(n385), .B2(n368), .A(n546), .ZN(n417) );
  NAND2_X1 U85 ( .A1(\mem[6][8] ), .A2(n368), .ZN(n546) );
  OAI21_X1 U86 ( .B1(n384), .B2(n555), .A(n545), .ZN(n416) );
  NAND2_X1 U87 ( .A1(\mem[6][9] ), .A2(n368), .ZN(n545) );
  OAI21_X1 U88 ( .B1(n383), .B2(n555), .A(n544), .ZN(n415) );
  NAND2_X1 U89 ( .A1(\mem[6][10] ), .A2(n368), .ZN(n544) );
  OAI21_X1 U90 ( .B1(n382), .B2(n555), .A(n543), .ZN(n414) );
  NAND2_X1 U91 ( .A1(\mem[6][11] ), .A2(n368), .ZN(n543) );
  OAI21_X1 U92 ( .B1(n381), .B2(n555), .A(n542), .ZN(n413) );
  NAND2_X1 U93 ( .A1(\mem[6][12] ), .A2(n368), .ZN(n542) );
  OAI21_X1 U94 ( .B1(n380), .B2(n555), .A(n541), .ZN(n412) );
  NAND2_X1 U95 ( .A1(\mem[6][13] ), .A2(n368), .ZN(n541) );
  OAI21_X1 U96 ( .B1(n379), .B2(n555), .A(n540), .ZN(n411) );
  NAND2_X1 U97 ( .A1(\mem[6][14] ), .A2(n368), .ZN(n540) );
  OAI21_X1 U98 ( .B1(n386), .B2(n624), .A(n616), .ZN(n482) );
  NAND2_X1 U99 ( .A1(\mem[2][7] ), .A2(n372), .ZN(n616) );
  OAI21_X1 U100 ( .B1(n385), .B2(n372), .A(n615), .ZN(n481) );
  NAND2_X1 U101 ( .A1(\mem[2][8] ), .A2(n372), .ZN(n615) );
  OAI21_X1 U102 ( .B1(n384), .B2(n624), .A(n614), .ZN(n480) );
  NAND2_X1 U103 ( .A1(\mem[2][9] ), .A2(n372), .ZN(n614) );
  OAI21_X1 U104 ( .B1(n383), .B2(n624), .A(n613), .ZN(n479) );
  NAND2_X1 U105 ( .A1(\mem[2][10] ), .A2(n372), .ZN(n613) );
  OAI21_X1 U106 ( .B1(n382), .B2(n624), .A(n612), .ZN(n478) );
  NAND2_X1 U107 ( .A1(\mem[2][11] ), .A2(n372), .ZN(n612) );
  OAI21_X1 U108 ( .B1(n381), .B2(n624), .A(n611), .ZN(n477) );
  NAND2_X1 U109 ( .A1(\mem[2][12] ), .A2(n372), .ZN(n611) );
  OAI21_X1 U110 ( .B1(n380), .B2(n624), .A(n610), .ZN(n476) );
  NAND2_X1 U111 ( .A1(\mem[2][13] ), .A2(n372), .ZN(n610) );
  OAI21_X1 U112 ( .B1(n379), .B2(n624), .A(n609), .ZN(n475) );
  NAND2_X1 U113 ( .A1(\mem[2][14] ), .A2(n372), .ZN(n609) );
  OAI21_X1 U114 ( .B1(n386), .B2(n590), .A(n582), .ZN(n450) );
  NAND2_X1 U115 ( .A1(\mem[4][7] ), .A2(n370), .ZN(n582) );
  OAI21_X1 U116 ( .B1(n385), .B2(n370), .A(n581), .ZN(n449) );
  NAND2_X1 U117 ( .A1(\mem[4][8] ), .A2(n370), .ZN(n581) );
  OAI21_X1 U118 ( .B1(n384), .B2(n590), .A(n580), .ZN(n448) );
  NAND2_X1 U119 ( .A1(\mem[4][9] ), .A2(n370), .ZN(n580) );
  OAI21_X1 U120 ( .B1(n383), .B2(n590), .A(n579), .ZN(n447) );
  NAND2_X1 U121 ( .A1(\mem[4][10] ), .A2(n370), .ZN(n579) );
  OAI21_X1 U122 ( .B1(n382), .B2(n590), .A(n578), .ZN(n446) );
  NAND2_X1 U123 ( .A1(\mem[4][11] ), .A2(n370), .ZN(n578) );
  OAI21_X1 U124 ( .B1(n381), .B2(n590), .A(n577), .ZN(n445) );
  NAND2_X1 U125 ( .A1(\mem[4][12] ), .A2(n370), .ZN(n577) );
  OAI21_X1 U126 ( .B1(n380), .B2(n590), .A(n576), .ZN(n444) );
  NAND2_X1 U127 ( .A1(\mem[4][13] ), .A2(n370), .ZN(n576) );
  OAI21_X1 U128 ( .B1(n379), .B2(n590), .A(n575), .ZN(n443) );
  NAND2_X1 U129 ( .A1(\mem[4][14] ), .A2(n370), .ZN(n575) );
  OAI21_X1 U130 ( .B1(n659), .B2(n385), .A(n650), .ZN(n513) );
  NAND2_X1 U131 ( .A1(\mem[0][8] ), .A2(n374), .ZN(n650) );
  OAI21_X1 U132 ( .B1(n659), .B2(n384), .A(n649), .ZN(n512) );
  NAND2_X1 U133 ( .A1(\mem[0][9] ), .A2(n659), .ZN(n649) );
  OAI21_X1 U134 ( .B1(n374), .B2(n383), .A(n648), .ZN(n511) );
  NAND2_X1 U135 ( .A1(\mem[0][10] ), .A2(n659), .ZN(n648) );
  OAI21_X1 U136 ( .B1(n659), .B2(n382), .A(n647), .ZN(n510) );
  NAND2_X1 U137 ( .A1(\mem[0][11] ), .A2(n659), .ZN(n647) );
  OAI21_X1 U138 ( .B1(n659), .B2(n381), .A(n646), .ZN(n509) );
  NAND2_X1 U139 ( .A1(\mem[0][12] ), .A2(n659), .ZN(n646) );
  OAI21_X1 U140 ( .B1(n659), .B2(n380), .A(n645), .ZN(n508) );
  NAND2_X1 U141 ( .A1(\mem[0][13] ), .A2(n659), .ZN(n645) );
  OAI21_X1 U142 ( .B1(n659), .B2(n379), .A(n644), .ZN(n507) );
  NAND2_X1 U143 ( .A1(\mem[0][14] ), .A2(n659), .ZN(n644) );
  INV_X1 U144 ( .A(N10), .ZN(n375) );
  OAI21_X1 U145 ( .B1(n393), .B2(n641), .A(n640), .ZN(n505) );
  NAND2_X1 U146 ( .A1(\mem[1][0] ), .A2(n373), .ZN(n640) );
  OAI21_X1 U147 ( .B1(n392), .B2(n641), .A(n639), .ZN(n504) );
  NAND2_X1 U148 ( .A1(\mem[1][1] ), .A2(n373), .ZN(n639) );
  OAI21_X1 U149 ( .B1(n391), .B2(n641), .A(n638), .ZN(n503) );
  NAND2_X1 U150 ( .A1(\mem[1][2] ), .A2(n373), .ZN(n638) );
  OAI21_X1 U151 ( .B1(n390), .B2(n641), .A(n637), .ZN(n502) );
  NAND2_X1 U152 ( .A1(\mem[1][3] ), .A2(n373), .ZN(n637) );
  OAI21_X1 U153 ( .B1(n389), .B2(n641), .A(n636), .ZN(n501) );
  NAND2_X1 U154 ( .A1(\mem[1][4] ), .A2(n641), .ZN(n636) );
  OAI21_X1 U155 ( .B1(n388), .B2(n641), .A(n635), .ZN(n500) );
  NAND2_X1 U156 ( .A1(\mem[1][5] ), .A2(n641), .ZN(n635) );
  OAI21_X1 U157 ( .B1(n387), .B2(n641), .A(n634), .ZN(n499) );
  NAND2_X1 U158 ( .A1(\mem[1][6] ), .A2(n641), .ZN(n634) );
  OAI21_X1 U159 ( .B1(n378), .B2(n641), .A(n625), .ZN(n490) );
  NAND2_X1 U160 ( .A1(\mem[1][15] ), .A2(n373), .ZN(n625) );
  OAI21_X1 U161 ( .B1(n393), .B2(n624), .A(n623), .ZN(n489) );
  NAND2_X1 U162 ( .A1(\mem[2][0] ), .A2(n372), .ZN(n623) );
  OAI21_X1 U163 ( .B1(n392), .B2(n624), .A(n622), .ZN(n488) );
  NAND2_X1 U164 ( .A1(\mem[2][1] ), .A2(n372), .ZN(n622) );
  OAI21_X1 U165 ( .B1(n391), .B2(n624), .A(n621), .ZN(n487) );
  NAND2_X1 U166 ( .A1(\mem[2][2] ), .A2(n372), .ZN(n621) );
  OAI21_X1 U167 ( .B1(n390), .B2(n624), .A(n620), .ZN(n486) );
  NAND2_X1 U168 ( .A1(\mem[2][3] ), .A2(n372), .ZN(n620) );
  OAI21_X1 U169 ( .B1(n389), .B2(n624), .A(n619), .ZN(n485) );
  NAND2_X1 U170 ( .A1(\mem[2][4] ), .A2(n624), .ZN(n619) );
  OAI21_X1 U171 ( .B1(n388), .B2(n624), .A(n618), .ZN(n484) );
  NAND2_X1 U172 ( .A1(\mem[2][5] ), .A2(n624), .ZN(n618) );
  OAI21_X1 U173 ( .B1(n387), .B2(n624), .A(n617), .ZN(n483) );
  NAND2_X1 U174 ( .A1(\mem[2][6] ), .A2(n624), .ZN(n617) );
  OAI21_X1 U175 ( .B1(n378), .B2(n624), .A(n608), .ZN(n474) );
  NAND2_X1 U176 ( .A1(\mem[2][15] ), .A2(n372), .ZN(n608) );
  OAI21_X1 U177 ( .B1(n393), .B2(n371), .A(n606), .ZN(n473) );
  NAND2_X1 U178 ( .A1(\mem[3][0] ), .A2(n371), .ZN(n606) );
  OAI21_X1 U179 ( .B1(n392), .B2(n371), .A(n605), .ZN(n472) );
  NAND2_X1 U180 ( .A1(\mem[3][1] ), .A2(n607), .ZN(n605) );
  OAI21_X1 U181 ( .B1(n391), .B2(n371), .A(n604), .ZN(n471) );
  NAND2_X1 U182 ( .A1(\mem[3][2] ), .A2(n607), .ZN(n604) );
  OAI21_X1 U183 ( .B1(n390), .B2(n371), .A(n603), .ZN(n470) );
  NAND2_X1 U184 ( .A1(\mem[3][3] ), .A2(n607), .ZN(n603) );
  OAI21_X1 U185 ( .B1(n389), .B2(n371), .A(n602), .ZN(n469) );
  NAND2_X1 U186 ( .A1(\mem[3][4] ), .A2(n371), .ZN(n602) );
  OAI21_X1 U187 ( .B1(n388), .B2(n371), .A(n601), .ZN(n468) );
  NAND2_X1 U188 ( .A1(\mem[3][5] ), .A2(n371), .ZN(n601) );
  OAI21_X1 U189 ( .B1(n387), .B2(n371), .A(n600), .ZN(n467) );
  NAND2_X1 U190 ( .A1(\mem[3][6] ), .A2(n371), .ZN(n600) );
  OAI21_X1 U191 ( .B1(n378), .B2(n371), .A(n591), .ZN(n458) );
  NAND2_X1 U192 ( .A1(\mem[3][15] ), .A2(n371), .ZN(n591) );
  OAI21_X1 U193 ( .B1(n393), .B2(n590), .A(n589), .ZN(n457) );
  NAND2_X1 U194 ( .A1(\mem[4][0] ), .A2(n370), .ZN(n589) );
  OAI21_X1 U195 ( .B1(n392), .B2(n590), .A(n588), .ZN(n456) );
  NAND2_X1 U196 ( .A1(\mem[4][1] ), .A2(n370), .ZN(n588) );
  OAI21_X1 U197 ( .B1(n391), .B2(n590), .A(n587), .ZN(n455) );
  NAND2_X1 U198 ( .A1(\mem[4][2] ), .A2(n370), .ZN(n587) );
  OAI21_X1 U199 ( .B1(n390), .B2(n590), .A(n586), .ZN(n454) );
  NAND2_X1 U200 ( .A1(\mem[4][3] ), .A2(n370), .ZN(n586) );
  OAI21_X1 U201 ( .B1(n389), .B2(n590), .A(n585), .ZN(n453) );
  NAND2_X1 U202 ( .A1(\mem[4][4] ), .A2(n590), .ZN(n585) );
  OAI21_X1 U203 ( .B1(n388), .B2(n590), .A(n584), .ZN(n452) );
  NAND2_X1 U204 ( .A1(\mem[4][5] ), .A2(n590), .ZN(n584) );
  OAI21_X1 U205 ( .B1(n387), .B2(n590), .A(n583), .ZN(n451) );
  NAND2_X1 U206 ( .A1(\mem[4][6] ), .A2(n590), .ZN(n583) );
  OAI21_X1 U207 ( .B1(n378), .B2(n590), .A(n574), .ZN(n442) );
  NAND2_X1 U208 ( .A1(\mem[4][15] ), .A2(n370), .ZN(n574) );
  OAI21_X1 U209 ( .B1(n393), .B2(n572), .A(n571), .ZN(n441) );
  NAND2_X1 U210 ( .A1(\mem[5][0] ), .A2(n369), .ZN(n571) );
  OAI21_X1 U211 ( .B1(n392), .B2(n572), .A(n570), .ZN(n440) );
  NAND2_X1 U212 ( .A1(\mem[5][1] ), .A2(n369), .ZN(n570) );
  OAI21_X1 U213 ( .B1(n391), .B2(n572), .A(n569), .ZN(n439) );
  NAND2_X1 U214 ( .A1(\mem[5][2] ), .A2(n369), .ZN(n569) );
  OAI21_X1 U215 ( .B1(n390), .B2(n572), .A(n568), .ZN(n438) );
  NAND2_X1 U216 ( .A1(\mem[5][3] ), .A2(n369), .ZN(n568) );
  OAI21_X1 U217 ( .B1(n389), .B2(n572), .A(n567), .ZN(n437) );
  NAND2_X1 U218 ( .A1(\mem[5][4] ), .A2(n572), .ZN(n567) );
  OAI21_X1 U219 ( .B1(n388), .B2(n572), .A(n566), .ZN(n436) );
  NAND2_X1 U220 ( .A1(\mem[5][5] ), .A2(n572), .ZN(n566) );
  OAI21_X1 U221 ( .B1(n387), .B2(n572), .A(n565), .ZN(n435) );
  NAND2_X1 U222 ( .A1(\mem[5][6] ), .A2(n572), .ZN(n565) );
  OAI21_X1 U223 ( .B1(n378), .B2(n572), .A(n556), .ZN(n426) );
  NAND2_X1 U224 ( .A1(\mem[5][15] ), .A2(n369), .ZN(n556) );
  OAI21_X1 U225 ( .B1(n393), .B2(n555), .A(n554), .ZN(n425) );
  NAND2_X1 U226 ( .A1(\mem[6][0] ), .A2(n368), .ZN(n554) );
  OAI21_X1 U227 ( .B1(n392), .B2(n555), .A(n553), .ZN(n424) );
  NAND2_X1 U228 ( .A1(\mem[6][1] ), .A2(n368), .ZN(n553) );
  OAI21_X1 U229 ( .B1(n391), .B2(n555), .A(n552), .ZN(n423) );
  NAND2_X1 U230 ( .A1(\mem[6][2] ), .A2(n368), .ZN(n552) );
  OAI21_X1 U231 ( .B1(n390), .B2(n555), .A(n551), .ZN(n422) );
  NAND2_X1 U232 ( .A1(\mem[6][3] ), .A2(n368), .ZN(n551) );
  OAI21_X1 U233 ( .B1(n389), .B2(n555), .A(n550), .ZN(n421) );
  NAND2_X1 U234 ( .A1(\mem[6][4] ), .A2(n555), .ZN(n550) );
  OAI21_X1 U235 ( .B1(n388), .B2(n555), .A(n549), .ZN(n420) );
  NAND2_X1 U236 ( .A1(\mem[6][5] ), .A2(n555), .ZN(n549) );
  OAI21_X1 U237 ( .B1(n387), .B2(n555), .A(n548), .ZN(n419) );
  NAND2_X1 U238 ( .A1(\mem[6][6] ), .A2(n555), .ZN(n548) );
  OAI21_X1 U239 ( .B1(n378), .B2(n555), .A(n539), .ZN(n410) );
  NAND2_X1 U240 ( .A1(\mem[6][15] ), .A2(n368), .ZN(n539) );
  OAI21_X1 U241 ( .B1(n393), .B2(n538), .A(n537), .ZN(n409) );
  NAND2_X1 U242 ( .A1(\mem[7][0] ), .A2(n367), .ZN(n537) );
  OAI21_X1 U243 ( .B1(n392), .B2(n538), .A(n536), .ZN(n408) );
  NAND2_X1 U244 ( .A1(\mem[7][1] ), .A2(n367), .ZN(n536) );
  OAI21_X1 U245 ( .B1(n391), .B2(n538), .A(n535), .ZN(n407) );
  NAND2_X1 U246 ( .A1(\mem[7][2] ), .A2(n367), .ZN(n535) );
  OAI21_X1 U247 ( .B1(n390), .B2(n538), .A(n534), .ZN(n406) );
  NAND2_X1 U248 ( .A1(\mem[7][3] ), .A2(n367), .ZN(n534) );
  OAI21_X1 U249 ( .B1(n389), .B2(n538), .A(n533), .ZN(n405) );
  NAND2_X1 U250 ( .A1(\mem[7][4] ), .A2(n538), .ZN(n533) );
  OAI21_X1 U251 ( .B1(n388), .B2(n538), .A(n532), .ZN(n404) );
  NAND2_X1 U252 ( .A1(\mem[7][5] ), .A2(n538), .ZN(n532) );
  OAI21_X1 U253 ( .B1(n387), .B2(n538), .A(n531), .ZN(n403) );
  NAND2_X1 U254 ( .A1(\mem[7][6] ), .A2(n538), .ZN(n531) );
  OAI21_X1 U255 ( .B1(n378), .B2(n538), .A(n522), .ZN(n394) );
  NAND2_X1 U256 ( .A1(\mem[7][15] ), .A2(n367), .ZN(n522) );
  OAI21_X1 U257 ( .B1(n374), .B2(n393), .A(n658), .ZN(n521) );
  NAND2_X1 U258 ( .A1(\mem[0][0] ), .A2(n659), .ZN(n658) );
  OAI21_X1 U259 ( .B1(n374), .B2(n392), .A(n657), .ZN(n520) );
  NAND2_X1 U260 ( .A1(\mem[0][1] ), .A2(n659), .ZN(n657) );
  OAI21_X1 U261 ( .B1(n374), .B2(n391), .A(n656), .ZN(n519) );
  NAND2_X1 U262 ( .A1(\mem[0][2] ), .A2(n659), .ZN(n656) );
  OAI21_X1 U263 ( .B1(n374), .B2(n390), .A(n655), .ZN(n518) );
  NAND2_X1 U264 ( .A1(\mem[0][3] ), .A2(n659), .ZN(n655) );
  OAI21_X1 U265 ( .B1(n374), .B2(n389), .A(n654), .ZN(n517) );
  NAND2_X1 U266 ( .A1(\mem[0][4] ), .A2(n374), .ZN(n654) );
  OAI21_X1 U267 ( .B1(n374), .B2(n388), .A(n653), .ZN(n516) );
  NAND2_X1 U268 ( .A1(\mem[0][5] ), .A2(n374), .ZN(n653) );
  OAI21_X1 U269 ( .B1(n374), .B2(n387), .A(n652), .ZN(n515) );
  NAND2_X1 U270 ( .A1(\mem[0][6] ), .A2(n374), .ZN(n652) );
  OAI21_X1 U271 ( .B1(n374), .B2(n386), .A(n651), .ZN(n514) );
  NAND2_X1 U272 ( .A1(\mem[0][7] ), .A2(n374), .ZN(n651) );
  OAI21_X1 U273 ( .B1(n374), .B2(n378), .A(n643), .ZN(n506) );
  NAND2_X1 U274 ( .A1(\mem[0][15] ), .A2(n659), .ZN(n643) );
  INV_X1 U275 ( .A(N11), .ZN(n376) );
  INV_X1 U276 ( .A(data_in[0]), .ZN(n393) );
  INV_X1 U277 ( .A(data_in[1]), .ZN(n392) );
  INV_X1 U278 ( .A(data_in[2]), .ZN(n391) );
  INV_X1 U279 ( .A(data_in[3]), .ZN(n390) );
  INV_X1 U288 ( .A(data_in[4]), .ZN(n389) );
  INV_X1 U289 ( .A(data_in[5]), .ZN(n388) );
  INV_X1 U290 ( .A(data_in[6]), .ZN(n387) );
  INV_X1 U291 ( .A(data_in[7]), .ZN(n386) );
  INV_X1 U292 ( .A(data_in[8]), .ZN(n385) );
  INV_X1 U293 ( .A(data_in[9]), .ZN(n384) );
  INV_X1 U294 ( .A(data_in[10]), .ZN(n383) );
  INV_X1 U295 ( .A(data_in[11]), .ZN(n382) );
  INV_X1 U296 ( .A(data_in[12]), .ZN(n381) );
  INV_X1 U297 ( .A(data_in[13]), .ZN(n380) );
  INV_X1 U298 ( .A(data_in[14]), .ZN(n379) );
  INV_X1 U299 ( .A(data_in[15]), .ZN(n378) );
  MUX2_X1 U300 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n365), .Z(n1) );
  MUX2_X1 U301 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n366), .Z(n2) );
  MUX2_X1 U302 ( .A(n2), .B(n1), .S(n363), .Z(n3) );
  MUX2_X1 U303 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n364), .Z(n4) );
  MUX2_X1 U304 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n366), .Z(n5) );
  MUX2_X1 U305 ( .A(n5), .B(n4), .S(N11), .Z(n6) );
  MUX2_X1 U306 ( .A(n6), .B(n3), .S(N12), .Z(N28) );
  MUX2_X1 U307 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n364), .Z(n7) );
  MUX2_X1 U308 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n364), .Z(n8) );
  MUX2_X1 U309 ( .A(n8), .B(n7), .S(n363), .Z(n9) );
  MUX2_X1 U310 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n364), .Z(n10) );
  MUX2_X1 U311 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n364), .Z(n11) );
  MUX2_X1 U312 ( .A(n11), .B(n10), .S(n363), .Z(n12) );
  MUX2_X1 U313 ( .A(n12), .B(n9), .S(N12), .Z(N27) );
  MUX2_X1 U314 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n364), .Z(n13) );
  MUX2_X1 U315 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n364), .Z(n14) );
  MUX2_X1 U316 ( .A(n14), .B(n13), .S(n363), .Z(n15) );
  MUX2_X1 U317 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n364), .Z(n16) );
  MUX2_X1 U318 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n364), .Z(n17) );
  MUX2_X1 U319 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U320 ( .A(n18), .B(n15), .S(N12), .Z(N26) );
  MUX2_X1 U321 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n364), .Z(n19) );
  MUX2_X1 U322 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n364), .Z(n286) );
  MUX2_X1 U323 ( .A(n286), .B(n19), .S(n363), .Z(n287) );
  MUX2_X1 U324 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n364), .Z(n288) );
  MUX2_X1 U325 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n364), .Z(n289) );
  MUX2_X1 U326 ( .A(n289), .B(n288), .S(N11), .Z(n290) );
  MUX2_X1 U327 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n365), .Z(n291) );
  MUX2_X1 U328 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n364), .Z(n292) );
  MUX2_X1 U329 ( .A(n292), .B(n291), .S(n363), .Z(n293) );
  MUX2_X1 U330 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n364), .Z(n294) );
  MUX2_X1 U331 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n366), .Z(n295) );
  MUX2_X1 U332 ( .A(n295), .B(n294), .S(n363), .Z(n296) );
  MUX2_X1 U333 ( .A(n296), .B(n293), .S(N12), .Z(N24) );
  MUX2_X1 U334 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n364), .Z(n297) );
  MUX2_X1 U335 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n365), .Z(n298) );
  MUX2_X1 U336 ( .A(n298), .B(n297), .S(n363), .Z(n299) );
  MUX2_X1 U337 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n366), .Z(n300) );
  MUX2_X1 U338 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n364), .Z(n301) );
  MUX2_X1 U339 ( .A(n301), .B(n300), .S(n363), .Z(n302) );
  MUX2_X1 U340 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n366), .Z(n303) );
  MUX2_X1 U341 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n365), .Z(n304) );
  MUX2_X1 U342 ( .A(n304), .B(n303), .S(n363), .Z(n305) );
  MUX2_X1 U343 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n365), .Z(n306) );
  MUX2_X1 U344 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n364), .Z(n307) );
  MUX2_X1 U345 ( .A(n307), .B(n306), .S(n363), .Z(n308) );
  MUX2_X1 U346 ( .A(n308), .B(n305), .S(N12), .Z(N22) );
  MUX2_X1 U347 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n365), .Z(n309) );
  MUX2_X1 U348 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n366), .Z(n310) );
  MUX2_X1 U349 ( .A(n310), .B(n309), .S(n363), .Z(n311) );
  MUX2_X1 U350 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n364), .Z(n312) );
  MUX2_X1 U351 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n313) );
  MUX2_X1 U352 ( .A(n313), .B(n312), .S(n363), .Z(n314) );
  MUX2_X1 U353 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n365), .Z(n315) );
  MUX2_X1 U354 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n365), .Z(n316) );
  MUX2_X1 U355 ( .A(n316), .B(n315), .S(n363), .Z(n317) );
  MUX2_X1 U356 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n364), .Z(n318) );
  MUX2_X1 U357 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n364), .Z(n319) );
  MUX2_X1 U358 ( .A(n319), .B(n318), .S(n363), .Z(n320) );
  MUX2_X1 U359 ( .A(n320), .B(n317), .S(N12), .Z(N20) );
  MUX2_X1 U360 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n366), .Z(n321) );
  MUX2_X1 U361 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n366), .Z(n322) );
  MUX2_X1 U362 ( .A(n322), .B(n321), .S(n363), .Z(n323) );
  MUX2_X1 U363 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n366), .Z(n324) );
  MUX2_X1 U364 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n365), .Z(n325) );
  MUX2_X1 U365 ( .A(n325), .B(n324), .S(n363), .Z(n326) );
  MUX2_X1 U366 ( .A(n326), .B(n323), .S(N12), .Z(N19) );
  MUX2_X1 U367 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n365), .Z(n327) );
  MUX2_X1 U368 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n365), .Z(n328) );
  MUX2_X1 U369 ( .A(n328), .B(n327), .S(n363), .Z(n329) );
  MUX2_X1 U370 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n365), .Z(n330) );
  MUX2_X1 U371 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n365), .Z(n331) );
  MUX2_X1 U372 ( .A(n331), .B(n330), .S(n363), .Z(n332) );
  MUX2_X1 U373 ( .A(n332), .B(n329), .S(N12), .Z(N18) );
  MUX2_X1 U374 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n365), .Z(n333) );
  MUX2_X1 U375 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n365), .Z(n334) );
  MUX2_X1 U376 ( .A(n334), .B(n333), .S(N11), .Z(n335) );
  MUX2_X1 U377 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n365), .Z(n336) );
  MUX2_X1 U378 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n365), .Z(n337) );
  MUX2_X1 U379 ( .A(n337), .B(n336), .S(N11), .Z(n338) );
  MUX2_X1 U380 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n365), .Z(n339) );
  MUX2_X1 U381 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n365), .Z(n340) );
  MUX2_X1 U382 ( .A(n340), .B(n339), .S(n363), .Z(n341) );
  MUX2_X1 U383 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n365), .Z(n342) );
  MUX2_X1 U384 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n365), .Z(n343) );
  MUX2_X1 U385 ( .A(n343), .B(n342), .S(n363), .Z(n344) );
  MUX2_X1 U386 ( .A(n344), .B(n341), .S(N12), .Z(N16) );
  MUX2_X1 U387 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n366), .Z(n345) );
  MUX2_X1 U388 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n366), .Z(n346) );
  MUX2_X1 U389 ( .A(n346), .B(n345), .S(N11), .Z(n347) );
  MUX2_X1 U390 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n366), .Z(n348) );
  MUX2_X1 U391 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n366), .Z(n349) );
  MUX2_X1 U392 ( .A(n349), .B(n348), .S(N11), .Z(n350) );
  MUX2_X1 U393 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n366), .Z(n351) );
  MUX2_X1 U394 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n366), .Z(n352) );
  MUX2_X1 U395 ( .A(n352), .B(n351), .S(n363), .Z(n353) );
  MUX2_X1 U396 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n366), .Z(n354) );
  MUX2_X1 U397 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n366), .Z(n355) );
  MUX2_X1 U398 ( .A(n355), .B(n354), .S(n363), .Z(n356) );
  MUX2_X1 U399 ( .A(n356), .B(n353), .S(N12), .Z(N14) );
  MUX2_X1 U400 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n366), .Z(n357) );
  MUX2_X1 U401 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n366), .Z(n358) );
  MUX2_X1 U402 ( .A(n358), .B(n357), .S(N11), .Z(n359) );
  MUX2_X1 U403 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n366), .Z(n360) );
  MUX2_X1 U404 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n366), .Z(n361) );
  MUX2_X1 U405 ( .A(n361), .B(n360), .S(N11), .Z(n362) );
endmodule


module memory_WIDTH16_SIZE8_LOGSIZE3_3 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] ,
         \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][15] , \mem[6][14] , \mem[6][13] ,
         \mem[6][12] , \mem[6][11] , \mem[6][10] , \mem[6][9] , \mem[6][8] ,
         \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] ,
         \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[5][15] , \mem[5][14] ,
         \mem[5][13] , \mem[5][12] , \mem[5][11] , \mem[5][10] , \mem[5][9] ,
         \mem[5][8] , \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] ,
         \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][15] ,
         \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] , \mem[4][10] ,
         \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N14, N16, N18,
         N20, N22, N24, N26, N27, N28, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[14]  ( .D(N14), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N16), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N18), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[8]  ( .D(N20), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N22), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N24), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N26), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N28), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][15]  ( .D(n394), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n395), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n396), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n397), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n398), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n399), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n400), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n401), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n402), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n403), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n404), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n405), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n406), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n407), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n408), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n409), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n410), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n411), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n412), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n413), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n414), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n415), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n416), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n417), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n418), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n419), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n420), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n421), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n422), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n423), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n424), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n425), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n426), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n427), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n428), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n429), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n430), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n431), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n432), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n433), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n434), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n435), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n436), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n437), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n438), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n439), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n440), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n441), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n442), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n443), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n444), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n445), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n446), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n447), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n448), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n449), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n450), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n451), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n452), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n453), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n454), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n455), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n456), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n457), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n458), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n459), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n460), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n461), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n462), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n463), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n464), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n465), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n466), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n467), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n468), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n469), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n470), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n471), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n472), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n473), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n474), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n475), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n476), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n477), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n478), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n479), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n480), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n481), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n482), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n483), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n484), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n485), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n486), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n487), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n488), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n489), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n490), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n491), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n492), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n493), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n494), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n495), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n496), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n497), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n498), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n499), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n500), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n501), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n502), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n503), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n504), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n505), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n506), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n507), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n508), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n509), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n510), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n511), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n512), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n513), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n514), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n515), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n516), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n517), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n518), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n519), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n520), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n521), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U280 ( .A1(n375), .A2(n376), .A3(n642), .ZN(n659) );
  NAND3_X1 U281 ( .A1(n642), .A2(n376), .A3(N10), .ZN(n641) );
  NAND3_X1 U282 ( .A1(n642), .A2(n375), .A3(N11), .ZN(n624) );
  NAND3_X1 U283 ( .A1(N10), .A2(n642), .A3(N11), .ZN(n607) );
  NAND3_X1 U284 ( .A1(n375), .A2(n376), .A3(n573), .ZN(n590) );
  NAND3_X1 U285 ( .A1(N10), .A2(n376), .A3(n573), .ZN(n572) );
  NAND3_X1 U286 ( .A1(N11), .A2(n375), .A3(n573), .ZN(n555) );
  NAND3_X1 U287 ( .A1(N11), .A2(N10), .A3(n573), .ZN(n538) );
  DFF_X1 \data_out_reg[1]  ( .D(N27), .CK(clk), .Q(data_out[1]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n350), .SI(n347), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n326), .SI(n323), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n302), .SI(n299), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n290), .SI(n287), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[15]  ( .D(n362), .SI(n359), .SE(N12), .CK(clk), .Q(
        data_out[15]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n338), .SI(n335), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n314), .SI(n311), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  BUF_X1 U3 ( .A(N10), .Z(n366) );
  BUF_X1 U4 ( .A(n641), .Z(n373) );
  BUF_X1 U5 ( .A(n624), .Z(n372) );
  BUF_X1 U6 ( .A(n607), .Z(n371) );
  BUF_X1 U7 ( .A(n590), .Z(n370) );
  BUF_X1 U8 ( .A(n572), .Z(n369) );
  BUF_X1 U9 ( .A(n555), .Z(n368) );
  BUF_X1 U10 ( .A(n538), .Z(n367) );
  BUF_X1 U11 ( .A(N10), .Z(n364) );
  BUF_X1 U12 ( .A(N10), .Z(n365) );
  BUF_X1 U13 ( .A(n659), .Z(n374) );
  BUF_X1 U14 ( .A(N11), .Z(n363) );
  NOR2_X1 U15 ( .A1(n377), .A2(N12), .ZN(n642) );
  INV_X1 U16 ( .A(wr_en), .ZN(n377) );
  AND2_X1 U17 ( .A1(N12), .A2(wr_en), .ZN(n573) );
  OAI21_X1 U18 ( .B1(n386), .B2(n607), .A(n599), .ZN(n466) );
  NAND2_X1 U19 ( .A1(\mem[3][7] ), .A2(n371), .ZN(n599) );
  OAI21_X1 U20 ( .B1(n385), .B2(n371), .A(n598), .ZN(n465) );
  NAND2_X1 U21 ( .A1(\mem[3][8] ), .A2(n371), .ZN(n598) );
  OAI21_X1 U22 ( .B1(n384), .B2(n607), .A(n597), .ZN(n464) );
  NAND2_X1 U23 ( .A1(\mem[3][9] ), .A2(n371), .ZN(n597) );
  OAI21_X1 U24 ( .B1(n383), .B2(n607), .A(n596), .ZN(n463) );
  NAND2_X1 U25 ( .A1(\mem[3][10] ), .A2(n371), .ZN(n596) );
  OAI21_X1 U26 ( .B1(n382), .B2(n607), .A(n595), .ZN(n462) );
  NAND2_X1 U27 ( .A1(\mem[3][11] ), .A2(n371), .ZN(n595) );
  OAI21_X1 U28 ( .B1(n381), .B2(n607), .A(n594), .ZN(n461) );
  NAND2_X1 U29 ( .A1(\mem[3][12] ), .A2(n371), .ZN(n594) );
  OAI21_X1 U30 ( .B1(n380), .B2(n607), .A(n593), .ZN(n460) );
  NAND2_X1 U31 ( .A1(\mem[3][13] ), .A2(n371), .ZN(n593) );
  OAI21_X1 U32 ( .B1(n379), .B2(n607), .A(n592), .ZN(n459) );
  NAND2_X1 U33 ( .A1(\mem[3][14] ), .A2(n371), .ZN(n592) );
  OAI21_X1 U34 ( .B1(n386), .B2(n572), .A(n564), .ZN(n434) );
  NAND2_X1 U35 ( .A1(\mem[5][7] ), .A2(n369), .ZN(n564) );
  OAI21_X1 U36 ( .B1(n385), .B2(n369), .A(n563), .ZN(n433) );
  NAND2_X1 U37 ( .A1(\mem[5][8] ), .A2(n369), .ZN(n563) );
  OAI21_X1 U38 ( .B1(n384), .B2(n572), .A(n562), .ZN(n432) );
  NAND2_X1 U39 ( .A1(\mem[5][9] ), .A2(n369), .ZN(n562) );
  OAI21_X1 U40 ( .B1(n383), .B2(n572), .A(n561), .ZN(n431) );
  NAND2_X1 U41 ( .A1(\mem[5][10] ), .A2(n369), .ZN(n561) );
  OAI21_X1 U42 ( .B1(n382), .B2(n572), .A(n560), .ZN(n430) );
  NAND2_X1 U43 ( .A1(\mem[5][11] ), .A2(n369), .ZN(n560) );
  OAI21_X1 U44 ( .B1(n381), .B2(n572), .A(n559), .ZN(n429) );
  NAND2_X1 U45 ( .A1(\mem[5][12] ), .A2(n369), .ZN(n559) );
  OAI21_X1 U46 ( .B1(n380), .B2(n572), .A(n558), .ZN(n428) );
  NAND2_X1 U47 ( .A1(\mem[5][13] ), .A2(n369), .ZN(n558) );
  OAI21_X1 U48 ( .B1(n379), .B2(n572), .A(n557), .ZN(n427) );
  NAND2_X1 U49 ( .A1(\mem[5][14] ), .A2(n369), .ZN(n557) );
  OAI21_X1 U50 ( .B1(n386), .B2(n538), .A(n530), .ZN(n402) );
  NAND2_X1 U51 ( .A1(\mem[7][7] ), .A2(n367), .ZN(n530) );
  OAI21_X1 U52 ( .B1(n385), .B2(n367), .A(n529), .ZN(n401) );
  NAND2_X1 U53 ( .A1(\mem[7][8] ), .A2(n367), .ZN(n529) );
  OAI21_X1 U54 ( .B1(n384), .B2(n538), .A(n528), .ZN(n400) );
  NAND2_X1 U55 ( .A1(\mem[7][9] ), .A2(n367), .ZN(n528) );
  OAI21_X1 U56 ( .B1(n383), .B2(n538), .A(n527), .ZN(n399) );
  NAND2_X1 U57 ( .A1(\mem[7][10] ), .A2(n367), .ZN(n527) );
  OAI21_X1 U58 ( .B1(n382), .B2(n538), .A(n526), .ZN(n398) );
  NAND2_X1 U59 ( .A1(\mem[7][11] ), .A2(n367), .ZN(n526) );
  OAI21_X1 U60 ( .B1(n381), .B2(n538), .A(n525), .ZN(n397) );
  NAND2_X1 U61 ( .A1(\mem[7][12] ), .A2(n367), .ZN(n525) );
  OAI21_X1 U62 ( .B1(n380), .B2(n538), .A(n524), .ZN(n396) );
  NAND2_X1 U63 ( .A1(\mem[7][13] ), .A2(n367), .ZN(n524) );
  OAI21_X1 U64 ( .B1(n379), .B2(n538), .A(n523), .ZN(n395) );
  NAND2_X1 U65 ( .A1(\mem[7][14] ), .A2(n367), .ZN(n523) );
  OAI21_X1 U66 ( .B1(n382), .B2(n641), .A(n629), .ZN(n494) );
  NAND2_X1 U67 ( .A1(\mem[1][11] ), .A2(n373), .ZN(n629) );
  OAI21_X1 U68 ( .B1(n386), .B2(n555), .A(n547), .ZN(n418) );
  NAND2_X1 U69 ( .A1(\mem[6][7] ), .A2(n368), .ZN(n547) );
  OAI21_X1 U70 ( .B1(n385), .B2(n368), .A(n546), .ZN(n417) );
  NAND2_X1 U71 ( .A1(\mem[6][8] ), .A2(n368), .ZN(n546) );
  OAI21_X1 U72 ( .B1(n384), .B2(n555), .A(n545), .ZN(n416) );
  NAND2_X1 U73 ( .A1(\mem[6][9] ), .A2(n368), .ZN(n545) );
  OAI21_X1 U74 ( .B1(n383), .B2(n555), .A(n544), .ZN(n415) );
  NAND2_X1 U75 ( .A1(\mem[6][10] ), .A2(n368), .ZN(n544) );
  OAI21_X1 U76 ( .B1(n382), .B2(n555), .A(n543), .ZN(n414) );
  NAND2_X1 U77 ( .A1(\mem[6][11] ), .A2(n368), .ZN(n543) );
  OAI21_X1 U78 ( .B1(n381), .B2(n555), .A(n542), .ZN(n413) );
  NAND2_X1 U79 ( .A1(\mem[6][12] ), .A2(n368), .ZN(n542) );
  OAI21_X1 U80 ( .B1(n380), .B2(n555), .A(n541), .ZN(n412) );
  NAND2_X1 U81 ( .A1(\mem[6][13] ), .A2(n368), .ZN(n541) );
  OAI21_X1 U82 ( .B1(n379), .B2(n555), .A(n540), .ZN(n411) );
  NAND2_X1 U83 ( .A1(\mem[6][14] ), .A2(n368), .ZN(n540) );
  OAI21_X1 U84 ( .B1(n386), .B2(n373), .A(n633), .ZN(n498) );
  NAND2_X1 U85 ( .A1(\mem[1][7] ), .A2(n641), .ZN(n633) );
  OAI21_X1 U86 ( .B1(n385), .B2(n641), .A(n632), .ZN(n497) );
  NAND2_X1 U87 ( .A1(\mem[1][8] ), .A2(n373), .ZN(n632) );
  OAI21_X1 U88 ( .B1(n384), .B2(n641), .A(n631), .ZN(n496) );
  NAND2_X1 U89 ( .A1(\mem[1][9] ), .A2(n373), .ZN(n631) );
  OAI21_X1 U90 ( .B1(n383), .B2(n641), .A(n630), .ZN(n495) );
  NAND2_X1 U91 ( .A1(\mem[1][10] ), .A2(n373), .ZN(n630) );
  OAI21_X1 U92 ( .B1(n381), .B2(n641), .A(n628), .ZN(n493) );
  NAND2_X1 U93 ( .A1(\mem[1][12] ), .A2(n373), .ZN(n628) );
  OAI21_X1 U94 ( .B1(n380), .B2(n641), .A(n627), .ZN(n492) );
  NAND2_X1 U95 ( .A1(\mem[1][13] ), .A2(n373), .ZN(n627) );
  OAI21_X1 U96 ( .B1(n379), .B2(n641), .A(n626), .ZN(n491) );
  NAND2_X1 U97 ( .A1(\mem[1][14] ), .A2(n373), .ZN(n626) );
  OAI21_X1 U98 ( .B1(n386), .B2(n624), .A(n616), .ZN(n482) );
  NAND2_X1 U99 ( .A1(\mem[2][7] ), .A2(n372), .ZN(n616) );
  OAI21_X1 U100 ( .B1(n385), .B2(n372), .A(n615), .ZN(n481) );
  NAND2_X1 U101 ( .A1(\mem[2][8] ), .A2(n372), .ZN(n615) );
  OAI21_X1 U102 ( .B1(n384), .B2(n624), .A(n614), .ZN(n480) );
  NAND2_X1 U103 ( .A1(\mem[2][9] ), .A2(n372), .ZN(n614) );
  OAI21_X1 U104 ( .B1(n383), .B2(n624), .A(n613), .ZN(n479) );
  NAND2_X1 U105 ( .A1(\mem[2][10] ), .A2(n372), .ZN(n613) );
  OAI21_X1 U106 ( .B1(n382), .B2(n624), .A(n612), .ZN(n478) );
  NAND2_X1 U107 ( .A1(\mem[2][11] ), .A2(n372), .ZN(n612) );
  OAI21_X1 U108 ( .B1(n381), .B2(n624), .A(n611), .ZN(n477) );
  NAND2_X1 U109 ( .A1(\mem[2][12] ), .A2(n372), .ZN(n611) );
  OAI21_X1 U110 ( .B1(n380), .B2(n624), .A(n610), .ZN(n476) );
  NAND2_X1 U111 ( .A1(\mem[2][13] ), .A2(n372), .ZN(n610) );
  OAI21_X1 U112 ( .B1(n379), .B2(n624), .A(n609), .ZN(n475) );
  NAND2_X1 U113 ( .A1(\mem[2][14] ), .A2(n372), .ZN(n609) );
  OAI21_X1 U114 ( .B1(n386), .B2(n590), .A(n582), .ZN(n450) );
  NAND2_X1 U115 ( .A1(\mem[4][7] ), .A2(n370), .ZN(n582) );
  OAI21_X1 U116 ( .B1(n385), .B2(n370), .A(n581), .ZN(n449) );
  NAND2_X1 U117 ( .A1(\mem[4][8] ), .A2(n370), .ZN(n581) );
  OAI21_X1 U118 ( .B1(n384), .B2(n590), .A(n580), .ZN(n448) );
  NAND2_X1 U119 ( .A1(\mem[4][9] ), .A2(n370), .ZN(n580) );
  OAI21_X1 U120 ( .B1(n383), .B2(n590), .A(n579), .ZN(n447) );
  NAND2_X1 U121 ( .A1(\mem[4][10] ), .A2(n370), .ZN(n579) );
  OAI21_X1 U122 ( .B1(n382), .B2(n590), .A(n578), .ZN(n446) );
  NAND2_X1 U123 ( .A1(\mem[4][11] ), .A2(n370), .ZN(n578) );
  OAI21_X1 U124 ( .B1(n381), .B2(n590), .A(n577), .ZN(n445) );
  NAND2_X1 U125 ( .A1(\mem[4][12] ), .A2(n370), .ZN(n577) );
  OAI21_X1 U126 ( .B1(n380), .B2(n590), .A(n576), .ZN(n444) );
  NAND2_X1 U127 ( .A1(\mem[4][13] ), .A2(n370), .ZN(n576) );
  OAI21_X1 U128 ( .B1(n379), .B2(n590), .A(n575), .ZN(n443) );
  NAND2_X1 U129 ( .A1(\mem[4][14] ), .A2(n370), .ZN(n575) );
  OAI21_X1 U130 ( .B1(n374), .B2(n385), .A(n650), .ZN(n513) );
  NAND2_X1 U131 ( .A1(\mem[0][8] ), .A2(n374), .ZN(n650) );
  OAI21_X1 U132 ( .B1(n374), .B2(n384), .A(n649), .ZN(n512) );
  NAND2_X1 U133 ( .A1(\mem[0][9] ), .A2(n374), .ZN(n649) );
  OAI21_X1 U134 ( .B1(n374), .B2(n383), .A(n648), .ZN(n511) );
  NAND2_X1 U135 ( .A1(\mem[0][10] ), .A2(n659), .ZN(n648) );
  OAI21_X1 U136 ( .B1(n374), .B2(n382), .A(n647), .ZN(n510) );
  NAND2_X1 U137 ( .A1(\mem[0][11] ), .A2(n374), .ZN(n647) );
  OAI21_X1 U138 ( .B1(n374), .B2(n381), .A(n646), .ZN(n509) );
  NAND2_X1 U139 ( .A1(\mem[0][12] ), .A2(n659), .ZN(n646) );
  OAI21_X1 U140 ( .B1(n374), .B2(n380), .A(n645), .ZN(n508) );
  NAND2_X1 U141 ( .A1(\mem[0][13] ), .A2(n659), .ZN(n645) );
  OAI21_X1 U142 ( .B1(n374), .B2(n379), .A(n644), .ZN(n507) );
  NAND2_X1 U143 ( .A1(\mem[0][14] ), .A2(n659), .ZN(n644) );
  INV_X1 U144 ( .A(N10), .ZN(n375) );
  OAI21_X1 U145 ( .B1(n393), .B2(n641), .A(n640), .ZN(n505) );
  NAND2_X1 U146 ( .A1(\mem[1][0] ), .A2(n373), .ZN(n640) );
  OAI21_X1 U147 ( .B1(n392), .B2(n641), .A(n639), .ZN(n504) );
  NAND2_X1 U148 ( .A1(\mem[1][1] ), .A2(n373), .ZN(n639) );
  OAI21_X1 U149 ( .B1(n391), .B2(n641), .A(n638), .ZN(n503) );
  NAND2_X1 U150 ( .A1(\mem[1][2] ), .A2(n373), .ZN(n638) );
  OAI21_X1 U151 ( .B1(n390), .B2(n641), .A(n637), .ZN(n502) );
  NAND2_X1 U152 ( .A1(\mem[1][3] ), .A2(n373), .ZN(n637) );
  OAI21_X1 U153 ( .B1(n389), .B2(n641), .A(n636), .ZN(n501) );
  NAND2_X1 U154 ( .A1(\mem[1][4] ), .A2(n373), .ZN(n636) );
  OAI21_X1 U155 ( .B1(n388), .B2(n641), .A(n635), .ZN(n500) );
  NAND2_X1 U156 ( .A1(\mem[1][5] ), .A2(n641), .ZN(n635) );
  OAI21_X1 U157 ( .B1(n387), .B2(n641), .A(n634), .ZN(n499) );
  NAND2_X1 U158 ( .A1(\mem[1][6] ), .A2(n641), .ZN(n634) );
  OAI21_X1 U159 ( .B1(n378), .B2(n641), .A(n625), .ZN(n490) );
  NAND2_X1 U160 ( .A1(\mem[1][15] ), .A2(n373), .ZN(n625) );
  OAI21_X1 U161 ( .B1(n393), .B2(n624), .A(n623), .ZN(n489) );
  NAND2_X1 U162 ( .A1(\mem[2][0] ), .A2(n372), .ZN(n623) );
  OAI21_X1 U163 ( .B1(n392), .B2(n624), .A(n622), .ZN(n488) );
  NAND2_X1 U164 ( .A1(\mem[2][1] ), .A2(n372), .ZN(n622) );
  OAI21_X1 U165 ( .B1(n391), .B2(n624), .A(n621), .ZN(n487) );
  NAND2_X1 U166 ( .A1(\mem[2][2] ), .A2(n372), .ZN(n621) );
  OAI21_X1 U167 ( .B1(n390), .B2(n624), .A(n620), .ZN(n486) );
  NAND2_X1 U168 ( .A1(\mem[2][3] ), .A2(n372), .ZN(n620) );
  OAI21_X1 U169 ( .B1(n389), .B2(n624), .A(n619), .ZN(n485) );
  NAND2_X1 U170 ( .A1(\mem[2][4] ), .A2(n624), .ZN(n619) );
  OAI21_X1 U171 ( .B1(n388), .B2(n624), .A(n618), .ZN(n484) );
  NAND2_X1 U172 ( .A1(\mem[2][5] ), .A2(n624), .ZN(n618) );
  OAI21_X1 U173 ( .B1(n387), .B2(n624), .A(n617), .ZN(n483) );
  NAND2_X1 U174 ( .A1(\mem[2][6] ), .A2(n624), .ZN(n617) );
  OAI21_X1 U175 ( .B1(n378), .B2(n624), .A(n608), .ZN(n474) );
  NAND2_X1 U176 ( .A1(\mem[2][15] ), .A2(n372), .ZN(n608) );
  OAI21_X1 U177 ( .B1(n393), .B2(n607), .A(n606), .ZN(n473) );
  NAND2_X1 U178 ( .A1(\mem[3][0] ), .A2(n371), .ZN(n606) );
  OAI21_X1 U179 ( .B1(n392), .B2(n607), .A(n605), .ZN(n472) );
  NAND2_X1 U180 ( .A1(\mem[3][1] ), .A2(n371), .ZN(n605) );
  OAI21_X1 U181 ( .B1(n391), .B2(n607), .A(n604), .ZN(n471) );
  NAND2_X1 U182 ( .A1(\mem[3][2] ), .A2(n371), .ZN(n604) );
  OAI21_X1 U183 ( .B1(n390), .B2(n607), .A(n603), .ZN(n470) );
  NAND2_X1 U184 ( .A1(\mem[3][3] ), .A2(n371), .ZN(n603) );
  OAI21_X1 U185 ( .B1(n389), .B2(n607), .A(n602), .ZN(n469) );
  NAND2_X1 U186 ( .A1(\mem[3][4] ), .A2(n607), .ZN(n602) );
  OAI21_X1 U187 ( .B1(n388), .B2(n607), .A(n601), .ZN(n468) );
  NAND2_X1 U188 ( .A1(\mem[3][5] ), .A2(n607), .ZN(n601) );
  OAI21_X1 U189 ( .B1(n387), .B2(n607), .A(n600), .ZN(n467) );
  NAND2_X1 U190 ( .A1(\mem[3][6] ), .A2(n607), .ZN(n600) );
  OAI21_X1 U191 ( .B1(n378), .B2(n607), .A(n591), .ZN(n458) );
  NAND2_X1 U192 ( .A1(\mem[3][15] ), .A2(n371), .ZN(n591) );
  OAI21_X1 U193 ( .B1(n393), .B2(n590), .A(n589), .ZN(n457) );
  NAND2_X1 U194 ( .A1(\mem[4][0] ), .A2(n370), .ZN(n589) );
  OAI21_X1 U195 ( .B1(n392), .B2(n590), .A(n588), .ZN(n456) );
  NAND2_X1 U196 ( .A1(\mem[4][1] ), .A2(n370), .ZN(n588) );
  OAI21_X1 U197 ( .B1(n391), .B2(n590), .A(n587), .ZN(n455) );
  NAND2_X1 U198 ( .A1(\mem[4][2] ), .A2(n370), .ZN(n587) );
  OAI21_X1 U199 ( .B1(n390), .B2(n590), .A(n586), .ZN(n454) );
  NAND2_X1 U200 ( .A1(\mem[4][3] ), .A2(n370), .ZN(n586) );
  OAI21_X1 U201 ( .B1(n389), .B2(n590), .A(n585), .ZN(n453) );
  NAND2_X1 U202 ( .A1(\mem[4][4] ), .A2(n590), .ZN(n585) );
  OAI21_X1 U203 ( .B1(n388), .B2(n590), .A(n584), .ZN(n452) );
  NAND2_X1 U204 ( .A1(\mem[4][5] ), .A2(n590), .ZN(n584) );
  OAI21_X1 U205 ( .B1(n387), .B2(n590), .A(n583), .ZN(n451) );
  NAND2_X1 U206 ( .A1(\mem[4][6] ), .A2(n590), .ZN(n583) );
  OAI21_X1 U207 ( .B1(n378), .B2(n590), .A(n574), .ZN(n442) );
  NAND2_X1 U208 ( .A1(\mem[4][15] ), .A2(n370), .ZN(n574) );
  OAI21_X1 U209 ( .B1(n393), .B2(n572), .A(n571), .ZN(n441) );
  NAND2_X1 U210 ( .A1(\mem[5][0] ), .A2(n369), .ZN(n571) );
  OAI21_X1 U211 ( .B1(n392), .B2(n572), .A(n570), .ZN(n440) );
  NAND2_X1 U212 ( .A1(\mem[5][1] ), .A2(n369), .ZN(n570) );
  OAI21_X1 U213 ( .B1(n391), .B2(n572), .A(n569), .ZN(n439) );
  NAND2_X1 U214 ( .A1(\mem[5][2] ), .A2(n369), .ZN(n569) );
  OAI21_X1 U215 ( .B1(n390), .B2(n572), .A(n568), .ZN(n438) );
  NAND2_X1 U216 ( .A1(\mem[5][3] ), .A2(n369), .ZN(n568) );
  OAI21_X1 U217 ( .B1(n389), .B2(n572), .A(n567), .ZN(n437) );
  NAND2_X1 U218 ( .A1(\mem[5][4] ), .A2(n572), .ZN(n567) );
  OAI21_X1 U219 ( .B1(n388), .B2(n572), .A(n566), .ZN(n436) );
  NAND2_X1 U220 ( .A1(\mem[5][5] ), .A2(n572), .ZN(n566) );
  OAI21_X1 U221 ( .B1(n387), .B2(n572), .A(n565), .ZN(n435) );
  NAND2_X1 U222 ( .A1(\mem[5][6] ), .A2(n572), .ZN(n565) );
  OAI21_X1 U223 ( .B1(n378), .B2(n572), .A(n556), .ZN(n426) );
  NAND2_X1 U224 ( .A1(\mem[5][15] ), .A2(n369), .ZN(n556) );
  OAI21_X1 U225 ( .B1(n393), .B2(n555), .A(n554), .ZN(n425) );
  NAND2_X1 U226 ( .A1(\mem[6][0] ), .A2(n368), .ZN(n554) );
  OAI21_X1 U227 ( .B1(n392), .B2(n555), .A(n553), .ZN(n424) );
  NAND2_X1 U228 ( .A1(\mem[6][1] ), .A2(n368), .ZN(n553) );
  OAI21_X1 U229 ( .B1(n391), .B2(n555), .A(n552), .ZN(n423) );
  NAND2_X1 U230 ( .A1(\mem[6][2] ), .A2(n368), .ZN(n552) );
  OAI21_X1 U231 ( .B1(n390), .B2(n555), .A(n551), .ZN(n422) );
  NAND2_X1 U232 ( .A1(\mem[6][3] ), .A2(n368), .ZN(n551) );
  OAI21_X1 U233 ( .B1(n389), .B2(n555), .A(n550), .ZN(n421) );
  NAND2_X1 U234 ( .A1(\mem[6][4] ), .A2(n555), .ZN(n550) );
  OAI21_X1 U235 ( .B1(n388), .B2(n555), .A(n549), .ZN(n420) );
  NAND2_X1 U236 ( .A1(\mem[6][5] ), .A2(n555), .ZN(n549) );
  OAI21_X1 U237 ( .B1(n387), .B2(n555), .A(n548), .ZN(n419) );
  NAND2_X1 U238 ( .A1(\mem[6][6] ), .A2(n555), .ZN(n548) );
  OAI21_X1 U239 ( .B1(n378), .B2(n555), .A(n539), .ZN(n410) );
  NAND2_X1 U240 ( .A1(\mem[6][15] ), .A2(n368), .ZN(n539) );
  OAI21_X1 U241 ( .B1(n393), .B2(n538), .A(n537), .ZN(n409) );
  NAND2_X1 U242 ( .A1(\mem[7][0] ), .A2(n367), .ZN(n537) );
  OAI21_X1 U243 ( .B1(n392), .B2(n538), .A(n536), .ZN(n408) );
  NAND2_X1 U244 ( .A1(\mem[7][1] ), .A2(n367), .ZN(n536) );
  OAI21_X1 U245 ( .B1(n391), .B2(n538), .A(n535), .ZN(n407) );
  NAND2_X1 U246 ( .A1(\mem[7][2] ), .A2(n367), .ZN(n535) );
  OAI21_X1 U247 ( .B1(n390), .B2(n538), .A(n534), .ZN(n406) );
  NAND2_X1 U248 ( .A1(\mem[7][3] ), .A2(n367), .ZN(n534) );
  OAI21_X1 U249 ( .B1(n389), .B2(n538), .A(n533), .ZN(n405) );
  NAND2_X1 U250 ( .A1(\mem[7][4] ), .A2(n538), .ZN(n533) );
  OAI21_X1 U251 ( .B1(n388), .B2(n538), .A(n532), .ZN(n404) );
  NAND2_X1 U252 ( .A1(\mem[7][5] ), .A2(n538), .ZN(n532) );
  OAI21_X1 U253 ( .B1(n387), .B2(n538), .A(n531), .ZN(n403) );
  NAND2_X1 U254 ( .A1(\mem[7][6] ), .A2(n538), .ZN(n531) );
  OAI21_X1 U255 ( .B1(n378), .B2(n538), .A(n522), .ZN(n394) );
  NAND2_X1 U256 ( .A1(\mem[7][15] ), .A2(n367), .ZN(n522) );
  OAI21_X1 U257 ( .B1(n659), .B2(n393), .A(n658), .ZN(n521) );
  NAND2_X1 U258 ( .A1(\mem[0][0] ), .A2(n374), .ZN(n658) );
  OAI21_X1 U259 ( .B1(n659), .B2(n392), .A(n657), .ZN(n520) );
  NAND2_X1 U260 ( .A1(\mem[0][1] ), .A2(n374), .ZN(n657) );
  OAI21_X1 U261 ( .B1(n659), .B2(n391), .A(n656), .ZN(n519) );
  NAND2_X1 U262 ( .A1(\mem[0][2] ), .A2(n374), .ZN(n656) );
  OAI21_X1 U263 ( .B1(n659), .B2(n390), .A(n655), .ZN(n518) );
  NAND2_X1 U264 ( .A1(\mem[0][3] ), .A2(n374), .ZN(n655) );
  OAI21_X1 U265 ( .B1(n659), .B2(n389), .A(n654), .ZN(n517) );
  NAND2_X1 U266 ( .A1(\mem[0][4] ), .A2(n374), .ZN(n654) );
  OAI21_X1 U267 ( .B1(n659), .B2(n388), .A(n653), .ZN(n516) );
  NAND2_X1 U268 ( .A1(\mem[0][5] ), .A2(n659), .ZN(n653) );
  OAI21_X1 U269 ( .B1(n659), .B2(n387), .A(n652), .ZN(n515) );
  NAND2_X1 U270 ( .A1(\mem[0][6] ), .A2(n659), .ZN(n652) );
  OAI21_X1 U271 ( .B1(n659), .B2(n386), .A(n651), .ZN(n514) );
  NAND2_X1 U272 ( .A1(\mem[0][7] ), .A2(n659), .ZN(n651) );
  OAI21_X1 U273 ( .B1(n659), .B2(n378), .A(n643), .ZN(n506) );
  NAND2_X1 U274 ( .A1(\mem[0][15] ), .A2(n374), .ZN(n643) );
  INV_X1 U275 ( .A(N11), .ZN(n376) );
  INV_X1 U276 ( .A(data_in[0]), .ZN(n393) );
  INV_X1 U277 ( .A(data_in[1]), .ZN(n392) );
  INV_X1 U278 ( .A(data_in[2]), .ZN(n391) );
  INV_X1 U279 ( .A(data_in[3]), .ZN(n390) );
  INV_X1 U288 ( .A(data_in[4]), .ZN(n389) );
  INV_X1 U289 ( .A(data_in[5]), .ZN(n388) );
  INV_X1 U290 ( .A(data_in[6]), .ZN(n387) );
  INV_X1 U291 ( .A(data_in[7]), .ZN(n386) );
  INV_X1 U292 ( .A(data_in[8]), .ZN(n385) );
  INV_X1 U293 ( .A(data_in[9]), .ZN(n384) );
  INV_X1 U294 ( .A(data_in[10]), .ZN(n383) );
  INV_X1 U295 ( .A(data_in[11]), .ZN(n382) );
  INV_X1 U296 ( .A(data_in[12]), .ZN(n381) );
  INV_X1 U297 ( .A(data_in[13]), .ZN(n380) );
  INV_X1 U298 ( .A(data_in[14]), .ZN(n379) );
  INV_X1 U299 ( .A(data_in[15]), .ZN(n378) );
  MUX2_X1 U300 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n366), .Z(n1) );
  MUX2_X1 U301 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n364), .Z(n2) );
  MUX2_X1 U302 ( .A(n2), .B(n1), .S(n363), .Z(n3) );
  MUX2_X1 U303 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n365), .Z(n4) );
  MUX2_X1 U304 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n365), .Z(n5) );
  MUX2_X1 U305 ( .A(n5), .B(n4), .S(n363), .Z(n6) );
  MUX2_X1 U306 ( .A(n6), .B(n3), .S(N12), .Z(N28) );
  MUX2_X1 U307 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n364), .Z(n7) );
  MUX2_X1 U308 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n364), .Z(n8) );
  MUX2_X1 U309 ( .A(n8), .B(n7), .S(n363), .Z(n9) );
  MUX2_X1 U310 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n364), .Z(n10) );
  MUX2_X1 U311 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n364), .Z(n11) );
  MUX2_X1 U312 ( .A(n11), .B(n10), .S(n363), .Z(n12) );
  MUX2_X1 U313 ( .A(n12), .B(n9), .S(N12), .Z(N27) );
  MUX2_X1 U314 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n364), .Z(n13) );
  MUX2_X1 U315 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n364), .Z(n14) );
  MUX2_X1 U316 ( .A(n14), .B(n13), .S(n363), .Z(n15) );
  MUX2_X1 U317 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n364), .Z(n16) );
  MUX2_X1 U318 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n364), .Z(n17) );
  MUX2_X1 U319 ( .A(n17), .B(n16), .S(n363), .Z(n18) );
  MUX2_X1 U320 ( .A(n18), .B(n15), .S(N12), .Z(N26) );
  MUX2_X1 U321 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n364), .Z(n19) );
  MUX2_X1 U322 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n364), .Z(n286) );
  MUX2_X1 U323 ( .A(n286), .B(n19), .S(n363), .Z(n287) );
  MUX2_X1 U324 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n364), .Z(n288) );
  MUX2_X1 U325 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n364), .Z(n289) );
  MUX2_X1 U326 ( .A(n289), .B(n288), .S(n363), .Z(n290) );
  MUX2_X1 U327 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n365), .Z(n291) );
  MUX2_X1 U328 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n365), .Z(n292) );
  MUX2_X1 U329 ( .A(n292), .B(n291), .S(n363), .Z(n293) );
  MUX2_X1 U330 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n365), .Z(n294) );
  MUX2_X1 U331 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n365), .Z(n295) );
  MUX2_X1 U332 ( .A(n295), .B(n294), .S(N11), .Z(n296) );
  MUX2_X1 U333 ( .A(n296), .B(n293), .S(N12), .Z(N24) );
  MUX2_X1 U334 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n365), .Z(n297) );
  MUX2_X1 U335 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n365), .Z(n298) );
  MUX2_X1 U336 ( .A(n298), .B(n297), .S(N11), .Z(n299) );
  MUX2_X1 U337 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n365), .Z(n300) );
  MUX2_X1 U338 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n365), .Z(n301) );
  MUX2_X1 U339 ( .A(n301), .B(n300), .S(N11), .Z(n302) );
  MUX2_X1 U340 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n365), .Z(n303) );
  MUX2_X1 U341 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n365), .Z(n304) );
  MUX2_X1 U342 ( .A(n304), .B(n303), .S(N11), .Z(n305) );
  MUX2_X1 U343 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n365), .Z(n306) );
  MUX2_X1 U344 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n365), .Z(n307) );
  MUX2_X1 U345 ( .A(n307), .B(n306), .S(N11), .Z(n308) );
  MUX2_X1 U346 ( .A(n308), .B(n305), .S(N12), .Z(N22) );
  MUX2_X1 U347 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n364), .Z(n309) );
  MUX2_X1 U348 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n366), .Z(n310) );
  MUX2_X1 U349 ( .A(n310), .B(n309), .S(N11), .Z(n311) );
  MUX2_X1 U350 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n366), .Z(n312) );
  MUX2_X1 U351 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n365), .Z(n313) );
  MUX2_X1 U352 ( .A(n313), .B(n312), .S(n363), .Z(n314) );
  MUX2_X1 U353 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n364), .Z(n315) );
  MUX2_X1 U354 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n364), .Z(n316) );
  MUX2_X1 U355 ( .A(n316), .B(n315), .S(N11), .Z(n317) );
  MUX2_X1 U356 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n366), .Z(n318) );
  MUX2_X1 U357 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n366), .Z(n319) );
  MUX2_X1 U358 ( .A(n319), .B(n318), .S(N11), .Z(n320) );
  MUX2_X1 U359 ( .A(n320), .B(n317), .S(N12), .Z(N20) );
  MUX2_X1 U360 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n365), .Z(n321) );
  MUX2_X1 U361 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n364), .Z(n322) );
  MUX2_X1 U362 ( .A(n322), .B(n321), .S(N11), .Z(n323) );
  MUX2_X1 U363 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n364), .Z(n324) );
  MUX2_X1 U364 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n366), .Z(n325) );
  MUX2_X1 U365 ( .A(n325), .B(n324), .S(n363), .Z(n326) );
  MUX2_X1 U366 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n366), .Z(n327) );
  MUX2_X1 U367 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n365), .Z(n328) );
  MUX2_X1 U368 ( .A(n328), .B(n327), .S(n363), .Z(n329) );
  MUX2_X1 U369 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n364), .Z(n330) );
  MUX2_X1 U370 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n364), .Z(n331) );
  MUX2_X1 U371 ( .A(n331), .B(n330), .S(n363), .Z(n332) );
  MUX2_X1 U372 ( .A(n332), .B(n329), .S(N12), .Z(N18) );
  MUX2_X1 U373 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n366), .Z(n333) );
  MUX2_X1 U374 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n365), .Z(n334) );
  MUX2_X1 U375 ( .A(n334), .B(n333), .S(N11), .Z(n335) );
  MUX2_X1 U376 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n365), .Z(n336) );
  MUX2_X1 U377 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n365), .Z(n337) );
  MUX2_X1 U378 ( .A(n337), .B(n336), .S(N11), .Z(n338) );
  MUX2_X1 U379 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n364), .Z(n339) );
  MUX2_X1 U380 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n366), .Z(n340) );
  MUX2_X1 U381 ( .A(n340), .B(n339), .S(n363), .Z(n341) );
  MUX2_X1 U382 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n365), .Z(n342) );
  MUX2_X1 U383 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n366), .Z(n343) );
  MUX2_X1 U384 ( .A(n343), .B(n342), .S(N11), .Z(n344) );
  MUX2_X1 U385 ( .A(n344), .B(n341), .S(N12), .Z(N16) );
  MUX2_X1 U386 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n366), .Z(n345) );
  MUX2_X1 U387 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n366), .Z(n346) );
  MUX2_X1 U388 ( .A(n346), .B(n345), .S(N11), .Z(n347) );
  MUX2_X1 U389 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n366), .Z(n348) );
  MUX2_X1 U390 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n366), .Z(n349) );
  MUX2_X1 U391 ( .A(n349), .B(n348), .S(N11), .Z(n350) );
  MUX2_X1 U392 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n366), .Z(n351) );
  MUX2_X1 U393 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n366), .Z(n352) );
  MUX2_X1 U394 ( .A(n352), .B(n351), .S(n363), .Z(n353) );
  MUX2_X1 U395 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n366), .Z(n354) );
  MUX2_X1 U396 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n366), .Z(n355) );
  MUX2_X1 U397 ( .A(n355), .B(n354), .S(N11), .Z(n356) );
  MUX2_X1 U398 ( .A(n356), .B(n353), .S(N12), .Z(N14) );
  MUX2_X1 U399 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n366), .Z(n357) );
  MUX2_X1 U400 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n366), .Z(n358) );
  MUX2_X1 U401 ( .A(n358), .B(n357), .S(N11), .Z(n359) );
  MUX2_X1 U402 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n366), .Z(n360) );
  MUX2_X1 U403 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n366), .Z(n361) );
  MUX2_X1 U404 ( .A(n361), .B(n360), .S(N11), .Z(n362) );
endmodule


module memory_WIDTH16_SIZE8_LOGSIZE3_2 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] ,
         \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][15] , \mem[6][14] , \mem[6][13] ,
         \mem[6][12] , \mem[6][11] , \mem[6][10] , \mem[6][9] , \mem[6][8] ,
         \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] ,
         \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[5][15] , \mem[5][14] ,
         \mem[5][13] , \mem[5][12] , \mem[5][11] , \mem[5][10] , \mem[5][9] ,
         \mem[5][8] , \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] ,
         \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][15] ,
         \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] , \mem[4][10] ,
         \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N13, N14, N16,
         N18, N21, N22, N24, N26, N28, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[14]  ( .D(N14), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N16), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N18), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[7]  ( .D(N21), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N22), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N24), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N26), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N28), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][15]  ( .D(n394), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n395), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n396), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n397), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n398), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n399), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n400), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n401), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n402), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n403), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n404), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n405), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n406), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n407), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n408), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n409), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n410), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n411), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n412), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n413), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n414), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n415), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n416), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n417), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n418), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n419), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n420), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n421), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n422), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n423), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n424), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n425), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n426), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n427), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n428), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n429), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n430), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n431), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n432), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n433), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n434), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n435), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n436), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n437), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n438), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n439), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n440), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n441), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n442), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n443), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n444), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n445), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n446), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n447), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n448), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n449), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n450), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n451), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n452), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n453), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n454), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n455), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n456), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n457), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n458), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n459), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n460), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n461), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n462), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n463), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n464), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n465), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n466), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n467), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n468), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n469), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n470), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n471), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n472), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n473), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n474), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n475), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n476), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n477), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n478), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n479), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n480), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n481), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n482), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n483), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n484), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n485), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n486), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n487), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n488), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n489), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n490), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n491), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n492), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n493), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n494), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n495), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n496), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n497), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n498), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n499), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n500), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n501), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n502), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n503), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n504), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n505), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n506), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n507), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n508), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n509), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n510), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n511), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n512), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n513), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n514), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n515), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n516), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n517), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n518), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n519), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n520), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n521), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U280 ( .A1(n375), .A2(n376), .A3(n642), .ZN(n659) );
  NAND3_X1 U281 ( .A1(n642), .A2(n376), .A3(N10), .ZN(n641) );
  NAND3_X1 U282 ( .A1(n642), .A2(n375), .A3(N11), .ZN(n624) );
  NAND3_X1 U283 ( .A1(N10), .A2(n642), .A3(N11), .ZN(n607) );
  NAND3_X1 U284 ( .A1(n375), .A2(n376), .A3(n573), .ZN(n590) );
  NAND3_X1 U285 ( .A1(N10), .A2(n376), .A3(n573), .ZN(n572) );
  NAND3_X1 U286 ( .A1(N11), .A2(n375), .A3(n573), .ZN(n555) );
  NAND3_X1 U287 ( .A1(N11), .A2(N10), .A3(n573), .ZN(n538) );
  DFF_X1 \data_out_reg[15]  ( .D(N13), .CK(clk), .Q(data_out[15]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n302), .SI(n299), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n338), .SI(n335), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[8]  ( .D(n320), .SI(n317), .SE(N12), .CK(clk), .Q(
        data_out[8]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n290), .SI(n287), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[1]  ( .D(n12), .SI(n9), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n326), .SI(n323), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n350), .SI(n347), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  BUF_X1 U3 ( .A(N10), .Z(n365) );
  BUF_X1 U4 ( .A(N10), .Z(n366) );
  BUF_X1 U5 ( .A(n659), .Z(n374) );
  BUF_X1 U6 ( .A(n641), .Z(n373) );
  BUF_X1 U7 ( .A(n624), .Z(n372) );
  BUF_X1 U8 ( .A(n572), .Z(n369) );
  BUF_X1 U9 ( .A(n555), .Z(n368) );
  BUF_X1 U10 ( .A(n538), .Z(n367) );
  BUF_X1 U11 ( .A(n607), .Z(n371) );
  BUF_X1 U12 ( .A(n590), .Z(n370) );
  BUF_X1 U13 ( .A(N11), .Z(n363) );
  AND2_X1 U14 ( .A1(N12), .A2(wr_en), .ZN(n573) );
  OAI21_X1 U15 ( .B1(n386), .B2(n607), .A(n599), .ZN(n466) );
  NAND2_X1 U16 ( .A1(\mem[3][7] ), .A2(n371), .ZN(n599) );
  OAI21_X1 U17 ( .B1(n385), .B2(n607), .A(n598), .ZN(n465) );
  NAND2_X1 U18 ( .A1(\mem[3][8] ), .A2(n607), .ZN(n598) );
  OAI21_X1 U19 ( .B1(n384), .B2(n607), .A(n597), .ZN(n464) );
  NAND2_X1 U20 ( .A1(\mem[3][9] ), .A2(n607), .ZN(n597) );
  OAI21_X1 U21 ( .B1(n383), .B2(n607), .A(n596), .ZN(n463) );
  NAND2_X1 U22 ( .A1(\mem[3][10] ), .A2(n607), .ZN(n596) );
  OAI21_X1 U23 ( .B1(n382), .B2(n607), .A(n595), .ZN(n462) );
  NAND2_X1 U24 ( .A1(\mem[3][11] ), .A2(n607), .ZN(n595) );
  OAI21_X1 U25 ( .B1(n381), .B2(n607), .A(n594), .ZN(n461) );
  NAND2_X1 U26 ( .A1(\mem[3][12] ), .A2(n607), .ZN(n594) );
  OAI21_X1 U27 ( .B1(n380), .B2(n607), .A(n593), .ZN(n460) );
  NAND2_X1 U28 ( .A1(\mem[3][13] ), .A2(n607), .ZN(n593) );
  OAI21_X1 U29 ( .B1(n379), .B2(n607), .A(n592), .ZN(n459) );
  NAND2_X1 U30 ( .A1(\mem[3][14] ), .A2(n607), .ZN(n592) );
  OAI21_X1 U31 ( .B1(n386), .B2(n572), .A(n564), .ZN(n434) );
  NAND2_X1 U32 ( .A1(\mem[5][7] ), .A2(n369), .ZN(n564) );
  OAI21_X1 U33 ( .B1(n385), .B2(n369), .A(n563), .ZN(n433) );
  NAND2_X1 U34 ( .A1(\mem[5][8] ), .A2(n369), .ZN(n563) );
  OAI21_X1 U35 ( .B1(n384), .B2(n572), .A(n562), .ZN(n432) );
  NAND2_X1 U36 ( .A1(\mem[5][9] ), .A2(n369), .ZN(n562) );
  OAI21_X1 U37 ( .B1(n383), .B2(n572), .A(n561), .ZN(n431) );
  NAND2_X1 U38 ( .A1(\mem[5][10] ), .A2(n369), .ZN(n561) );
  OAI21_X1 U39 ( .B1(n382), .B2(n572), .A(n560), .ZN(n430) );
  NAND2_X1 U40 ( .A1(\mem[5][11] ), .A2(n369), .ZN(n560) );
  OAI21_X1 U41 ( .B1(n381), .B2(n572), .A(n559), .ZN(n429) );
  NAND2_X1 U42 ( .A1(\mem[5][12] ), .A2(n369), .ZN(n559) );
  OAI21_X1 U43 ( .B1(n380), .B2(n572), .A(n558), .ZN(n428) );
  NAND2_X1 U44 ( .A1(\mem[5][13] ), .A2(n369), .ZN(n558) );
  OAI21_X1 U45 ( .B1(n379), .B2(n572), .A(n557), .ZN(n427) );
  NAND2_X1 U46 ( .A1(\mem[5][14] ), .A2(n369), .ZN(n557) );
  OAI21_X1 U47 ( .B1(n386), .B2(n538), .A(n530), .ZN(n402) );
  NAND2_X1 U48 ( .A1(\mem[7][7] ), .A2(n367), .ZN(n530) );
  OAI21_X1 U49 ( .B1(n385), .B2(n367), .A(n529), .ZN(n401) );
  NAND2_X1 U50 ( .A1(\mem[7][8] ), .A2(n367), .ZN(n529) );
  OAI21_X1 U51 ( .B1(n384), .B2(n538), .A(n528), .ZN(n400) );
  NAND2_X1 U52 ( .A1(\mem[7][9] ), .A2(n367), .ZN(n528) );
  OAI21_X1 U53 ( .B1(n383), .B2(n538), .A(n527), .ZN(n399) );
  NAND2_X1 U54 ( .A1(\mem[7][10] ), .A2(n367), .ZN(n527) );
  OAI21_X1 U55 ( .B1(n382), .B2(n538), .A(n526), .ZN(n398) );
  NAND2_X1 U56 ( .A1(\mem[7][11] ), .A2(n367), .ZN(n526) );
  OAI21_X1 U57 ( .B1(n381), .B2(n538), .A(n525), .ZN(n397) );
  NAND2_X1 U58 ( .A1(\mem[7][12] ), .A2(n367), .ZN(n525) );
  OAI21_X1 U59 ( .B1(n380), .B2(n538), .A(n524), .ZN(n396) );
  NAND2_X1 U60 ( .A1(\mem[7][13] ), .A2(n367), .ZN(n524) );
  OAI21_X1 U61 ( .B1(n379), .B2(n538), .A(n523), .ZN(n395) );
  NAND2_X1 U62 ( .A1(\mem[7][14] ), .A2(n367), .ZN(n523) );
  OAI21_X1 U63 ( .B1(n384), .B2(n641), .A(n631), .ZN(n496) );
  NAND2_X1 U64 ( .A1(\mem[1][9] ), .A2(n373), .ZN(n631) );
  OAI21_X1 U65 ( .B1(n383), .B2(n373), .A(n630), .ZN(n495) );
  NAND2_X1 U66 ( .A1(\mem[1][10] ), .A2(n373), .ZN(n630) );
  OAI21_X1 U67 ( .B1(n382), .B2(n641), .A(n629), .ZN(n494) );
  NAND2_X1 U68 ( .A1(\mem[1][11] ), .A2(n373), .ZN(n629) );
  OAI21_X1 U69 ( .B1(n380), .B2(n641), .A(n627), .ZN(n492) );
  NAND2_X1 U70 ( .A1(\mem[1][13] ), .A2(n373), .ZN(n627) );
  OAI21_X1 U71 ( .B1(n379), .B2(n641), .A(n626), .ZN(n491) );
  NAND2_X1 U72 ( .A1(\mem[1][14] ), .A2(n373), .ZN(n626) );
  OAI21_X1 U73 ( .B1(n386), .B2(n555), .A(n547), .ZN(n418) );
  NAND2_X1 U74 ( .A1(\mem[6][7] ), .A2(n368), .ZN(n547) );
  OAI21_X1 U75 ( .B1(n385), .B2(n368), .A(n546), .ZN(n417) );
  NAND2_X1 U76 ( .A1(\mem[6][8] ), .A2(n368), .ZN(n546) );
  OAI21_X1 U77 ( .B1(n384), .B2(n555), .A(n545), .ZN(n416) );
  NAND2_X1 U78 ( .A1(\mem[6][9] ), .A2(n368), .ZN(n545) );
  OAI21_X1 U79 ( .B1(n383), .B2(n555), .A(n544), .ZN(n415) );
  NAND2_X1 U80 ( .A1(\mem[6][10] ), .A2(n368), .ZN(n544) );
  OAI21_X1 U81 ( .B1(n382), .B2(n555), .A(n543), .ZN(n414) );
  NAND2_X1 U82 ( .A1(\mem[6][11] ), .A2(n368), .ZN(n543) );
  OAI21_X1 U83 ( .B1(n381), .B2(n555), .A(n542), .ZN(n413) );
  NAND2_X1 U84 ( .A1(\mem[6][12] ), .A2(n368), .ZN(n542) );
  OAI21_X1 U85 ( .B1(n380), .B2(n555), .A(n541), .ZN(n412) );
  NAND2_X1 U86 ( .A1(\mem[6][13] ), .A2(n368), .ZN(n541) );
  OAI21_X1 U87 ( .B1(n379), .B2(n555), .A(n540), .ZN(n411) );
  NAND2_X1 U88 ( .A1(\mem[6][14] ), .A2(n368), .ZN(n540) );
  OAI21_X1 U89 ( .B1(n386), .B2(n641), .A(n633), .ZN(n498) );
  NAND2_X1 U90 ( .A1(\mem[1][7] ), .A2(n641), .ZN(n633) );
  OAI21_X1 U91 ( .B1(n385), .B2(n641), .A(n632), .ZN(n497) );
  NAND2_X1 U92 ( .A1(\mem[1][8] ), .A2(n373), .ZN(n632) );
  OAI21_X1 U93 ( .B1(n381), .B2(n641), .A(n628), .ZN(n493) );
  NAND2_X1 U94 ( .A1(\mem[1][12] ), .A2(n373), .ZN(n628) );
  OAI21_X1 U95 ( .B1(n386), .B2(n624), .A(n616), .ZN(n482) );
  NAND2_X1 U96 ( .A1(\mem[2][7] ), .A2(n372), .ZN(n616) );
  OAI21_X1 U97 ( .B1(n385), .B2(n372), .A(n615), .ZN(n481) );
  NAND2_X1 U98 ( .A1(\mem[2][8] ), .A2(n372), .ZN(n615) );
  OAI21_X1 U99 ( .B1(n384), .B2(n624), .A(n614), .ZN(n480) );
  NAND2_X1 U100 ( .A1(\mem[2][9] ), .A2(n372), .ZN(n614) );
  OAI21_X1 U101 ( .B1(n383), .B2(n624), .A(n613), .ZN(n479) );
  NAND2_X1 U102 ( .A1(\mem[2][10] ), .A2(n372), .ZN(n613) );
  OAI21_X1 U103 ( .B1(n382), .B2(n624), .A(n612), .ZN(n478) );
  NAND2_X1 U104 ( .A1(\mem[2][11] ), .A2(n372), .ZN(n612) );
  OAI21_X1 U105 ( .B1(n381), .B2(n624), .A(n611), .ZN(n477) );
  NAND2_X1 U106 ( .A1(\mem[2][12] ), .A2(n372), .ZN(n611) );
  OAI21_X1 U107 ( .B1(n380), .B2(n624), .A(n610), .ZN(n476) );
  NAND2_X1 U108 ( .A1(\mem[2][13] ), .A2(n372), .ZN(n610) );
  OAI21_X1 U109 ( .B1(n379), .B2(n624), .A(n609), .ZN(n475) );
  NAND2_X1 U110 ( .A1(\mem[2][14] ), .A2(n372), .ZN(n609) );
  OAI21_X1 U111 ( .B1(n386), .B2(n370), .A(n582), .ZN(n450) );
  NAND2_X1 U112 ( .A1(\mem[4][7] ), .A2(n370), .ZN(n582) );
  OAI21_X1 U113 ( .B1(n385), .B2(n370), .A(n581), .ZN(n449) );
  NAND2_X1 U114 ( .A1(\mem[4][8] ), .A2(n590), .ZN(n581) );
  OAI21_X1 U115 ( .B1(n384), .B2(n370), .A(n580), .ZN(n448) );
  NAND2_X1 U116 ( .A1(\mem[4][9] ), .A2(n590), .ZN(n580) );
  OAI21_X1 U117 ( .B1(n383), .B2(n370), .A(n579), .ZN(n447) );
  NAND2_X1 U118 ( .A1(\mem[4][10] ), .A2(n590), .ZN(n579) );
  OAI21_X1 U119 ( .B1(n382), .B2(n370), .A(n578), .ZN(n446) );
  NAND2_X1 U120 ( .A1(\mem[4][11] ), .A2(n590), .ZN(n578) );
  OAI21_X1 U121 ( .B1(n381), .B2(n370), .A(n577), .ZN(n445) );
  NAND2_X1 U122 ( .A1(\mem[4][12] ), .A2(n590), .ZN(n577) );
  OAI21_X1 U123 ( .B1(n380), .B2(n370), .A(n576), .ZN(n444) );
  NAND2_X1 U124 ( .A1(\mem[4][13] ), .A2(n590), .ZN(n576) );
  OAI21_X1 U125 ( .B1(n379), .B2(n370), .A(n575), .ZN(n443) );
  NAND2_X1 U126 ( .A1(\mem[4][14] ), .A2(n590), .ZN(n575) );
  INV_X1 U127 ( .A(N10), .ZN(n375) );
  OAI21_X1 U128 ( .B1(n659), .B2(n385), .A(n650), .ZN(n513) );
  NAND2_X1 U129 ( .A1(\mem[0][8] ), .A2(n374), .ZN(n650) );
  OAI21_X1 U130 ( .B1(n659), .B2(n384), .A(n649), .ZN(n512) );
  NAND2_X1 U131 ( .A1(\mem[0][9] ), .A2(n659), .ZN(n649) );
  OAI21_X1 U132 ( .B1(n374), .B2(n383), .A(n648), .ZN(n511) );
  NAND2_X1 U133 ( .A1(\mem[0][10] ), .A2(n659), .ZN(n648) );
  OAI21_X1 U134 ( .B1(n659), .B2(n382), .A(n647), .ZN(n510) );
  NAND2_X1 U135 ( .A1(\mem[0][11] ), .A2(n659), .ZN(n647) );
  OAI21_X1 U136 ( .B1(n659), .B2(n381), .A(n646), .ZN(n509) );
  NAND2_X1 U137 ( .A1(\mem[0][12] ), .A2(n659), .ZN(n646) );
  OAI21_X1 U138 ( .B1(n659), .B2(n380), .A(n645), .ZN(n508) );
  NAND2_X1 U139 ( .A1(\mem[0][13] ), .A2(n659), .ZN(n645) );
  OAI21_X1 U140 ( .B1(n659), .B2(n379), .A(n644), .ZN(n507) );
  NAND2_X1 U141 ( .A1(\mem[0][14] ), .A2(n659), .ZN(n644) );
  OAI21_X1 U142 ( .B1(n393), .B2(n641), .A(n640), .ZN(n505) );
  NAND2_X1 U143 ( .A1(\mem[1][0] ), .A2(n373), .ZN(n640) );
  OAI21_X1 U144 ( .B1(n392), .B2(n641), .A(n639), .ZN(n504) );
  NAND2_X1 U145 ( .A1(\mem[1][1] ), .A2(n373), .ZN(n639) );
  OAI21_X1 U146 ( .B1(n391), .B2(n641), .A(n638), .ZN(n503) );
  NAND2_X1 U147 ( .A1(\mem[1][2] ), .A2(n373), .ZN(n638) );
  OAI21_X1 U148 ( .B1(n390), .B2(n641), .A(n637), .ZN(n502) );
  NAND2_X1 U149 ( .A1(\mem[1][3] ), .A2(n373), .ZN(n637) );
  OAI21_X1 U150 ( .B1(n389), .B2(n641), .A(n636), .ZN(n501) );
  NAND2_X1 U151 ( .A1(\mem[1][4] ), .A2(n373), .ZN(n636) );
  OAI21_X1 U152 ( .B1(n388), .B2(n641), .A(n635), .ZN(n500) );
  NAND2_X1 U153 ( .A1(\mem[1][5] ), .A2(n641), .ZN(n635) );
  OAI21_X1 U154 ( .B1(n387), .B2(n641), .A(n634), .ZN(n499) );
  NAND2_X1 U155 ( .A1(\mem[1][6] ), .A2(n641), .ZN(n634) );
  OAI21_X1 U156 ( .B1(n378), .B2(n641), .A(n625), .ZN(n490) );
  NAND2_X1 U157 ( .A1(\mem[1][15] ), .A2(n373), .ZN(n625) );
  OAI21_X1 U158 ( .B1(n393), .B2(n624), .A(n623), .ZN(n489) );
  NAND2_X1 U159 ( .A1(\mem[2][0] ), .A2(n372), .ZN(n623) );
  OAI21_X1 U160 ( .B1(n392), .B2(n624), .A(n622), .ZN(n488) );
  NAND2_X1 U161 ( .A1(\mem[2][1] ), .A2(n372), .ZN(n622) );
  OAI21_X1 U162 ( .B1(n391), .B2(n624), .A(n621), .ZN(n487) );
  NAND2_X1 U163 ( .A1(\mem[2][2] ), .A2(n372), .ZN(n621) );
  OAI21_X1 U164 ( .B1(n390), .B2(n624), .A(n620), .ZN(n486) );
  NAND2_X1 U165 ( .A1(\mem[2][3] ), .A2(n372), .ZN(n620) );
  OAI21_X1 U166 ( .B1(n389), .B2(n624), .A(n619), .ZN(n485) );
  NAND2_X1 U167 ( .A1(\mem[2][4] ), .A2(n624), .ZN(n619) );
  OAI21_X1 U168 ( .B1(n388), .B2(n624), .A(n618), .ZN(n484) );
  NAND2_X1 U169 ( .A1(\mem[2][5] ), .A2(n624), .ZN(n618) );
  OAI21_X1 U170 ( .B1(n387), .B2(n624), .A(n617), .ZN(n483) );
  NAND2_X1 U171 ( .A1(\mem[2][6] ), .A2(n624), .ZN(n617) );
  OAI21_X1 U172 ( .B1(n378), .B2(n624), .A(n608), .ZN(n474) );
  NAND2_X1 U173 ( .A1(\mem[2][15] ), .A2(n372), .ZN(n608) );
  OAI21_X1 U174 ( .B1(n393), .B2(n371), .A(n606), .ZN(n473) );
  NAND2_X1 U175 ( .A1(\mem[3][0] ), .A2(n371), .ZN(n606) );
  OAI21_X1 U176 ( .B1(n392), .B2(n371), .A(n605), .ZN(n472) );
  NAND2_X1 U177 ( .A1(\mem[3][1] ), .A2(n607), .ZN(n605) );
  OAI21_X1 U178 ( .B1(n391), .B2(n371), .A(n604), .ZN(n471) );
  NAND2_X1 U179 ( .A1(\mem[3][2] ), .A2(n607), .ZN(n604) );
  OAI21_X1 U180 ( .B1(n390), .B2(n371), .A(n603), .ZN(n470) );
  NAND2_X1 U181 ( .A1(\mem[3][3] ), .A2(n607), .ZN(n603) );
  OAI21_X1 U182 ( .B1(n389), .B2(n371), .A(n602), .ZN(n469) );
  NAND2_X1 U183 ( .A1(\mem[3][4] ), .A2(n371), .ZN(n602) );
  OAI21_X1 U184 ( .B1(n388), .B2(n371), .A(n601), .ZN(n468) );
  NAND2_X1 U185 ( .A1(\mem[3][5] ), .A2(n371), .ZN(n601) );
  OAI21_X1 U186 ( .B1(n387), .B2(n371), .A(n600), .ZN(n467) );
  NAND2_X1 U187 ( .A1(\mem[3][6] ), .A2(n371), .ZN(n600) );
  OAI21_X1 U188 ( .B1(n378), .B2(n371), .A(n591), .ZN(n458) );
  NAND2_X1 U189 ( .A1(\mem[3][15] ), .A2(n371), .ZN(n591) );
  OAI21_X1 U190 ( .B1(n393), .B2(n370), .A(n589), .ZN(n457) );
  NAND2_X1 U191 ( .A1(\mem[4][0] ), .A2(n590), .ZN(n589) );
  OAI21_X1 U192 ( .B1(n392), .B2(n590), .A(n588), .ZN(n456) );
  NAND2_X1 U193 ( .A1(\mem[4][1] ), .A2(n370), .ZN(n588) );
  OAI21_X1 U194 ( .B1(n391), .B2(n590), .A(n587), .ZN(n455) );
  NAND2_X1 U195 ( .A1(\mem[4][2] ), .A2(n590), .ZN(n587) );
  OAI21_X1 U196 ( .B1(n390), .B2(n590), .A(n586), .ZN(n454) );
  NAND2_X1 U197 ( .A1(\mem[4][3] ), .A2(n590), .ZN(n586) );
  OAI21_X1 U198 ( .B1(n389), .B2(n590), .A(n585), .ZN(n453) );
  NAND2_X1 U199 ( .A1(\mem[4][4] ), .A2(n370), .ZN(n585) );
  OAI21_X1 U200 ( .B1(n388), .B2(n590), .A(n584), .ZN(n452) );
  NAND2_X1 U201 ( .A1(\mem[4][5] ), .A2(n370), .ZN(n584) );
  OAI21_X1 U202 ( .B1(n387), .B2(n590), .A(n583), .ZN(n451) );
  NAND2_X1 U203 ( .A1(\mem[4][6] ), .A2(n370), .ZN(n583) );
  OAI21_X1 U204 ( .B1(n378), .B2(n590), .A(n574), .ZN(n442) );
  NAND2_X1 U205 ( .A1(\mem[4][15] ), .A2(n590), .ZN(n574) );
  OAI21_X1 U206 ( .B1(n393), .B2(n572), .A(n571), .ZN(n441) );
  NAND2_X1 U207 ( .A1(\mem[5][0] ), .A2(n369), .ZN(n571) );
  OAI21_X1 U208 ( .B1(n392), .B2(n572), .A(n570), .ZN(n440) );
  NAND2_X1 U209 ( .A1(\mem[5][1] ), .A2(n369), .ZN(n570) );
  OAI21_X1 U210 ( .B1(n391), .B2(n572), .A(n569), .ZN(n439) );
  NAND2_X1 U211 ( .A1(\mem[5][2] ), .A2(n369), .ZN(n569) );
  OAI21_X1 U212 ( .B1(n390), .B2(n572), .A(n568), .ZN(n438) );
  NAND2_X1 U213 ( .A1(\mem[5][3] ), .A2(n369), .ZN(n568) );
  OAI21_X1 U214 ( .B1(n389), .B2(n572), .A(n567), .ZN(n437) );
  NAND2_X1 U215 ( .A1(\mem[5][4] ), .A2(n572), .ZN(n567) );
  OAI21_X1 U216 ( .B1(n388), .B2(n572), .A(n566), .ZN(n436) );
  NAND2_X1 U217 ( .A1(\mem[5][5] ), .A2(n572), .ZN(n566) );
  OAI21_X1 U218 ( .B1(n387), .B2(n572), .A(n565), .ZN(n435) );
  NAND2_X1 U219 ( .A1(\mem[5][6] ), .A2(n572), .ZN(n565) );
  OAI21_X1 U220 ( .B1(n378), .B2(n572), .A(n556), .ZN(n426) );
  NAND2_X1 U221 ( .A1(\mem[5][15] ), .A2(n369), .ZN(n556) );
  OAI21_X1 U222 ( .B1(n393), .B2(n555), .A(n554), .ZN(n425) );
  NAND2_X1 U223 ( .A1(\mem[6][0] ), .A2(n368), .ZN(n554) );
  OAI21_X1 U224 ( .B1(n392), .B2(n555), .A(n553), .ZN(n424) );
  NAND2_X1 U225 ( .A1(\mem[6][1] ), .A2(n368), .ZN(n553) );
  OAI21_X1 U226 ( .B1(n391), .B2(n555), .A(n552), .ZN(n423) );
  NAND2_X1 U227 ( .A1(\mem[6][2] ), .A2(n368), .ZN(n552) );
  OAI21_X1 U228 ( .B1(n390), .B2(n555), .A(n551), .ZN(n422) );
  NAND2_X1 U229 ( .A1(\mem[6][3] ), .A2(n368), .ZN(n551) );
  OAI21_X1 U230 ( .B1(n389), .B2(n555), .A(n550), .ZN(n421) );
  NAND2_X1 U231 ( .A1(\mem[6][4] ), .A2(n555), .ZN(n550) );
  OAI21_X1 U232 ( .B1(n388), .B2(n555), .A(n549), .ZN(n420) );
  NAND2_X1 U233 ( .A1(\mem[6][5] ), .A2(n555), .ZN(n549) );
  OAI21_X1 U234 ( .B1(n387), .B2(n555), .A(n548), .ZN(n419) );
  NAND2_X1 U235 ( .A1(\mem[6][6] ), .A2(n555), .ZN(n548) );
  OAI21_X1 U236 ( .B1(n378), .B2(n555), .A(n539), .ZN(n410) );
  NAND2_X1 U237 ( .A1(\mem[6][15] ), .A2(n368), .ZN(n539) );
  OAI21_X1 U238 ( .B1(n393), .B2(n538), .A(n537), .ZN(n409) );
  NAND2_X1 U239 ( .A1(\mem[7][0] ), .A2(n367), .ZN(n537) );
  OAI21_X1 U240 ( .B1(n392), .B2(n538), .A(n536), .ZN(n408) );
  NAND2_X1 U241 ( .A1(\mem[7][1] ), .A2(n367), .ZN(n536) );
  OAI21_X1 U242 ( .B1(n391), .B2(n538), .A(n535), .ZN(n407) );
  NAND2_X1 U243 ( .A1(\mem[7][2] ), .A2(n367), .ZN(n535) );
  OAI21_X1 U244 ( .B1(n390), .B2(n538), .A(n534), .ZN(n406) );
  NAND2_X1 U245 ( .A1(\mem[7][3] ), .A2(n367), .ZN(n534) );
  OAI21_X1 U246 ( .B1(n389), .B2(n538), .A(n533), .ZN(n405) );
  NAND2_X1 U247 ( .A1(\mem[7][4] ), .A2(n538), .ZN(n533) );
  OAI21_X1 U248 ( .B1(n388), .B2(n538), .A(n532), .ZN(n404) );
  NAND2_X1 U249 ( .A1(\mem[7][5] ), .A2(n538), .ZN(n532) );
  OAI21_X1 U250 ( .B1(n387), .B2(n538), .A(n531), .ZN(n403) );
  NAND2_X1 U251 ( .A1(\mem[7][6] ), .A2(n538), .ZN(n531) );
  OAI21_X1 U252 ( .B1(n378), .B2(n538), .A(n522), .ZN(n394) );
  NAND2_X1 U253 ( .A1(\mem[7][15] ), .A2(n367), .ZN(n522) );
  OAI21_X1 U254 ( .B1(n374), .B2(n393), .A(n658), .ZN(n521) );
  NAND2_X1 U255 ( .A1(\mem[0][0] ), .A2(n659), .ZN(n658) );
  OAI21_X1 U256 ( .B1(n374), .B2(n392), .A(n657), .ZN(n520) );
  NAND2_X1 U257 ( .A1(\mem[0][1] ), .A2(n659), .ZN(n657) );
  OAI21_X1 U258 ( .B1(n374), .B2(n391), .A(n656), .ZN(n519) );
  NAND2_X1 U259 ( .A1(\mem[0][2] ), .A2(n659), .ZN(n656) );
  OAI21_X1 U260 ( .B1(n374), .B2(n390), .A(n655), .ZN(n518) );
  NAND2_X1 U261 ( .A1(\mem[0][3] ), .A2(n659), .ZN(n655) );
  OAI21_X1 U262 ( .B1(n374), .B2(n389), .A(n654), .ZN(n517) );
  NAND2_X1 U263 ( .A1(\mem[0][4] ), .A2(n374), .ZN(n654) );
  OAI21_X1 U264 ( .B1(n374), .B2(n388), .A(n653), .ZN(n516) );
  NAND2_X1 U265 ( .A1(\mem[0][5] ), .A2(n374), .ZN(n653) );
  OAI21_X1 U266 ( .B1(n374), .B2(n387), .A(n652), .ZN(n515) );
  NAND2_X1 U267 ( .A1(\mem[0][6] ), .A2(n374), .ZN(n652) );
  OAI21_X1 U268 ( .B1(n374), .B2(n386), .A(n651), .ZN(n514) );
  NAND2_X1 U269 ( .A1(\mem[0][7] ), .A2(n374), .ZN(n651) );
  OAI21_X1 U270 ( .B1(n374), .B2(n378), .A(n643), .ZN(n506) );
  NAND2_X1 U271 ( .A1(\mem[0][15] ), .A2(n659), .ZN(n643) );
  NOR2_X1 U272 ( .A1(n377), .A2(N12), .ZN(n642) );
  INV_X1 U273 ( .A(wr_en), .ZN(n377) );
  INV_X1 U274 ( .A(N11), .ZN(n376) );
  INV_X1 U275 ( .A(data_in[0]), .ZN(n393) );
  INV_X1 U276 ( .A(data_in[1]), .ZN(n392) );
  INV_X1 U277 ( .A(data_in[2]), .ZN(n391) );
  INV_X1 U278 ( .A(data_in[3]), .ZN(n390) );
  INV_X1 U279 ( .A(data_in[4]), .ZN(n389) );
  INV_X1 U288 ( .A(data_in[5]), .ZN(n388) );
  INV_X1 U289 ( .A(data_in[6]), .ZN(n387) );
  INV_X1 U290 ( .A(data_in[7]), .ZN(n386) );
  INV_X1 U291 ( .A(data_in[8]), .ZN(n385) );
  INV_X1 U292 ( .A(data_in[9]), .ZN(n384) );
  INV_X1 U293 ( .A(data_in[10]), .ZN(n383) );
  INV_X1 U294 ( .A(data_in[11]), .ZN(n382) );
  INV_X1 U295 ( .A(data_in[12]), .ZN(n381) );
  INV_X1 U296 ( .A(data_in[13]), .ZN(n380) );
  INV_X1 U297 ( .A(data_in[14]), .ZN(n379) );
  INV_X1 U298 ( .A(data_in[15]), .ZN(n378) );
  MUX2_X1 U299 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n364), .Z(n1) );
  MUX2_X1 U300 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n364), .Z(n2) );
  MUX2_X1 U301 ( .A(n2), .B(n1), .S(n363), .Z(n3) );
  MUX2_X1 U302 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n364), .Z(n4) );
  MUX2_X1 U303 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n364), .Z(n5) );
  MUX2_X1 U304 ( .A(n5), .B(n4), .S(n363), .Z(n6) );
  MUX2_X1 U305 ( .A(n6), .B(n3), .S(N12), .Z(N28) );
  MUX2_X1 U306 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n365), .Z(n7) );
  MUX2_X1 U307 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n366), .Z(n8) );
  MUX2_X1 U308 ( .A(n8), .B(n7), .S(n363), .Z(n9) );
  MUX2_X1 U309 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n364), .Z(n10) );
  MUX2_X1 U310 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(N10), .Z(n11) );
  MUX2_X1 U311 ( .A(n11), .B(n10), .S(n363), .Z(n12) );
  MUX2_X1 U312 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n366), .Z(n13) );
  MUX2_X1 U313 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n366), .Z(n14) );
  MUX2_X1 U314 ( .A(n14), .B(n13), .S(n363), .Z(n15) );
  MUX2_X1 U315 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n364), .Z(n16) );
  MUX2_X1 U316 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n366), .Z(n17) );
  MUX2_X1 U317 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U318 ( .A(n18), .B(n15), .S(N12), .Z(N26) );
  MUX2_X1 U319 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n364), .Z(n19) );
  MUX2_X1 U320 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n365), .Z(n286) );
  MUX2_X1 U321 ( .A(n286), .B(n19), .S(N11), .Z(n287) );
  MUX2_X1 U322 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n366), .Z(n288) );
  MUX2_X1 U323 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n289) );
  MUX2_X1 U324 ( .A(n289), .B(n288), .S(N11), .Z(n290) );
  MUX2_X1 U325 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n365), .Z(n291) );
  MUX2_X1 U326 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n365), .Z(n292) );
  MUX2_X1 U327 ( .A(n292), .B(n291), .S(n363), .Z(n293) );
  MUX2_X1 U328 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n364), .Z(n294) );
  MUX2_X1 U329 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n365), .Z(n295) );
  MUX2_X1 U330 ( .A(n295), .B(n294), .S(n363), .Z(n296) );
  MUX2_X1 U331 ( .A(n296), .B(n293), .S(N12), .Z(N24) );
  MUX2_X1 U332 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n365), .Z(n297) );
  MUX2_X1 U333 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n366), .Z(n298) );
  MUX2_X1 U334 ( .A(n298), .B(n297), .S(n363), .Z(n299) );
  MUX2_X1 U335 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n365), .Z(n300) );
  MUX2_X1 U336 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n364), .Z(n301) );
  MUX2_X1 U337 ( .A(n301), .B(n300), .S(n363), .Z(n302) );
  MUX2_X1 U338 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n366), .Z(n303) );
  MUX2_X1 U339 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n366), .Z(n304) );
  MUX2_X1 U340 ( .A(n304), .B(n303), .S(n363), .Z(n305) );
  MUX2_X1 U341 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n364), .Z(n306) );
  MUX2_X1 U342 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n364), .Z(n307) );
  MUX2_X1 U343 ( .A(n307), .B(n306), .S(n363), .Z(n308) );
  MUX2_X1 U344 ( .A(n308), .B(n305), .S(N12), .Z(N22) );
  MUX2_X1 U345 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n364), .Z(n309) );
  MUX2_X1 U346 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n364), .Z(n310) );
  MUX2_X1 U347 ( .A(n310), .B(n309), .S(n363), .Z(n311) );
  MUX2_X1 U348 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n364), .Z(n312) );
  MUX2_X1 U349 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n364), .Z(n313) );
  MUX2_X1 U350 ( .A(n313), .B(n312), .S(n363), .Z(n314) );
  MUX2_X1 U351 ( .A(n314), .B(n311), .S(N12), .Z(N21) );
  MUX2_X1 U352 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n364), .Z(n315) );
  MUX2_X1 U353 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n364), .Z(n316) );
  MUX2_X1 U354 ( .A(n316), .B(n315), .S(n363), .Z(n317) );
  MUX2_X1 U355 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n366), .Z(n318) );
  MUX2_X1 U356 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n365), .Z(n319) );
  MUX2_X1 U357 ( .A(n319), .B(n318), .S(n363), .Z(n320) );
  MUX2_X1 U358 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n364), .Z(n321) );
  MUX2_X1 U359 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n365), .Z(n322) );
  MUX2_X1 U360 ( .A(n322), .B(n321), .S(n363), .Z(n323) );
  MUX2_X1 U361 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(N10), .Z(n324) );
  MUX2_X1 U362 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n364), .Z(n325) );
  MUX2_X1 U363 ( .A(n325), .B(n324), .S(n363), .Z(n326) );
  MUX2_X1 U364 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n365), .Z(n327) );
  MUX2_X1 U365 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n365), .Z(n328) );
  MUX2_X1 U366 ( .A(n328), .B(n327), .S(n363), .Z(n329) );
  MUX2_X1 U367 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n365), .Z(n330) );
  MUX2_X1 U368 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n365), .Z(n331) );
  MUX2_X1 U369 ( .A(n331), .B(n330), .S(n363), .Z(n332) );
  MUX2_X1 U370 ( .A(n332), .B(n329), .S(N12), .Z(N18) );
  MUX2_X1 U371 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n365), .Z(n333) );
  MUX2_X1 U372 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n365), .Z(n334) );
  MUX2_X1 U373 ( .A(n334), .B(n333), .S(N11), .Z(n335) );
  MUX2_X1 U374 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n365), .Z(n336) );
  MUX2_X1 U375 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n365), .Z(n337) );
  MUX2_X1 U376 ( .A(n337), .B(n336), .S(N11), .Z(n338) );
  MUX2_X1 U377 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n365), .Z(n339) );
  MUX2_X1 U378 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n365), .Z(n340) );
  MUX2_X1 U379 ( .A(n340), .B(n339), .S(n363), .Z(n341) );
  MUX2_X1 U380 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n365), .Z(n342) );
  MUX2_X1 U381 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n365), .Z(n343) );
  MUX2_X1 U382 ( .A(n343), .B(n342), .S(n363), .Z(n344) );
  MUX2_X1 U383 ( .A(n344), .B(n341), .S(N12), .Z(N16) );
  MUX2_X1 U384 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n366), .Z(n345) );
  MUX2_X1 U385 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n366), .Z(n346) );
  MUX2_X1 U386 ( .A(n346), .B(n345), .S(N11), .Z(n347) );
  MUX2_X1 U387 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n366), .Z(n348) );
  MUX2_X1 U388 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n366), .Z(n349) );
  MUX2_X1 U389 ( .A(n349), .B(n348), .S(N11), .Z(n350) );
  MUX2_X1 U390 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n366), .Z(n351) );
  MUX2_X1 U391 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n366), .Z(n352) );
  MUX2_X1 U392 ( .A(n352), .B(n351), .S(n363), .Z(n353) );
  MUX2_X1 U393 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n366), .Z(n354) );
  MUX2_X1 U394 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n366), .Z(n355) );
  MUX2_X1 U395 ( .A(n355), .B(n354), .S(N11), .Z(n356) );
  MUX2_X1 U396 ( .A(n356), .B(n353), .S(N12), .Z(N14) );
  MUX2_X1 U397 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n366), .Z(n357) );
  MUX2_X1 U398 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n366), .Z(n358) );
  MUX2_X1 U399 ( .A(n358), .B(n357), .S(n363), .Z(n359) );
  MUX2_X1 U400 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n366), .Z(n360) );
  MUX2_X1 U401 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n366), .Z(n361) );
  MUX2_X1 U402 ( .A(n361), .B(n360), .S(N11), .Z(n362) );
  MUX2_X1 U403 ( .A(n362), .B(n359), .S(N12), .Z(N13) );
  CLKBUF_X1 U404 ( .A(N10), .Z(n364) );
endmodule


module memory_WIDTH16_SIZE8_LOGSIZE3_1 ( clk, data_in, data_out, addr, wr_en
 );
  input [15:0] data_in;
  output [15:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][15] , \mem[7][14] , \mem[7][13] , \mem[7][12] ,
         \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][15] , \mem[6][14] , \mem[6][13] ,
         \mem[6][12] , \mem[6][11] , \mem[6][10] , \mem[6][9] , \mem[6][8] ,
         \mem[6][7] , \mem[6][6] , \mem[6][5] , \mem[6][4] , \mem[6][3] ,
         \mem[6][2] , \mem[6][1] , \mem[6][0] , \mem[5][15] , \mem[5][14] ,
         \mem[5][13] , \mem[5][12] , \mem[5][11] , \mem[5][10] , \mem[5][9] ,
         \mem[5][8] , \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] ,
         \mem[5][3] , \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][15] ,
         \mem[4][14] , \mem[4][13] , \mem[4][12] , \mem[4][11] , \mem[4][10] ,
         \mem[4][9] , \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] ,
         \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][15] , \mem[2][14] , \mem[2][13] , \mem[2][12] ,
         \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][15] , \mem[1][14] , \mem[1][13] ,
         \mem[1][12] , \mem[1][11] , \mem[1][10] , \mem[1][9] , \mem[1][8] ,
         \mem[1][7] , \mem[1][6] , \mem[1][5] , \mem[1][4] , \mem[1][3] ,
         \mem[1][2] , \mem[1][1] , \mem[1][0] , \mem[0][15] , \mem[0][14] ,
         \mem[0][13] , \mem[0][12] , \mem[0][11] , \mem[0][10] , \mem[0][9] ,
         \mem[0][8] , \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] ,
         \mem[0][3] , \mem[0][2] , \mem[0][1] , \mem[0][0] , N13, N14, N16,
         N18, N20, N22, N24, N28, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[15]  ( .D(N13), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N14), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[12]  ( .D(N16), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[10]  ( .D(N18), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[8]  ( .D(N20), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[6]  ( .D(N22), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N24), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[0]  ( .D(N28), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][15]  ( .D(n394), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n395), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n396), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n397), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n398), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n399), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n400), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n401), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n402), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n403), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n404), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n405), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n406), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n407), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n408), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n409), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n410), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n411), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n412), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n413), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n414), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n415), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n416), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n417), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n418), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n419), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n420), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n421), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n422), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n423), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n424), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n425), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n426), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n427), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n428), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n429), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n430), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n431), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n432), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n433), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n434), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n435), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n436), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n437), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n438), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n439), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n440), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n441), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n442), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n443), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n444), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n445), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n446), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n447), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n448), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n449), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n450), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n451), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n452), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n453), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n454), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n455), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n456), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n457), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n458), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n459), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n460), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n461), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n462), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n463), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n464), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n465), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n466), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n467), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n468), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n469), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n470), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n471), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n472), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n473), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n474), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n475), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n476), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n477), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n478), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n479), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n480), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n481), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n482), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n483), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n484), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n485), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n486), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n487), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n488), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n489), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n490), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n491), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n492), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n493), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n494), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n495), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n496), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n497), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n498), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n499), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n500), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n501), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n502), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n503), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n504), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n505), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n506), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n507), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n508), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n509), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n510), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n511), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n512), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n513), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n514), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n515), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n516), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n517), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n518), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n519), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n520), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n521), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U280 ( .A1(n375), .A2(n376), .A3(n642), .ZN(n659) );
  NAND3_X1 U281 ( .A1(n642), .A2(n376), .A3(N10), .ZN(n641) );
  NAND3_X1 U282 ( .A1(n642), .A2(n375), .A3(N11), .ZN(n624) );
  NAND3_X1 U283 ( .A1(N10), .A2(n642), .A3(N11), .ZN(n607) );
  NAND3_X1 U284 ( .A1(n375), .A2(n376), .A3(n573), .ZN(n590) );
  NAND3_X1 U285 ( .A1(N10), .A2(n376), .A3(n573), .ZN(n572) );
  NAND3_X1 U286 ( .A1(N11), .A2(n375), .A3(n573), .ZN(n555) );
  NAND3_X1 U287 ( .A1(N11), .A2(N10), .A3(n573), .ZN(n538) );
  SDFF_X1 \data_out_reg[1]  ( .D(n12), .SI(n9), .SE(N12), .CK(clk), .Q(
        data_out[1]) );
  SDFF_X1 \data_out_reg[5]  ( .D(n302), .SI(n299), .SE(N12), .CK(clk), .Q(
        data_out[5]) );
  SDFF_X1 \data_out_reg[3]  ( .D(n290), .SI(n287), .SE(N12), .CK(clk), .Q(
        data_out[3]) );
  SDFF_X1 \data_out_reg[9]  ( .D(n326), .SI(n323), .SE(N12), .CK(clk), .Q(
        data_out[9]) );
  SDFF_X1 \data_out_reg[7]  ( .D(n314), .SI(n311), .SE(N12), .CK(clk), .Q(
        data_out[7]) );
  SDFF_X1 \data_out_reg[2]  ( .D(n18), .SI(n15), .SE(N12), .CK(clk), .Q(
        data_out[2]) );
  SDFF_X1 \data_out_reg[11]  ( .D(n338), .SI(n335), .SE(N12), .CK(clk), .Q(
        data_out[11]) );
  SDFF_X1 \data_out_reg[13]  ( .D(n350), .SI(n347), .SE(N12), .CK(clk), .Q(
        data_out[13]) );
  BUF_X1 U3 ( .A(n659), .Z(n374) );
  BUF_X1 U4 ( .A(n641), .Z(n373) );
  BUF_X1 U5 ( .A(n624), .Z(n372) );
  BUF_X1 U6 ( .A(n607), .Z(n371) );
  BUF_X1 U7 ( .A(n590), .Z(n370) );
  BUF_X1 U8 ( .A(n572), .Z(n369) );
  BUF_X1 U9 ( .A(n555), .Z(n368) );
  BUF_X1 U10 ( .A(n538), .Z(n367) );
  BUF_X1 U11 ( .A(N10), .Z(n364) );
  BUF_X1 U12 ( .A(N10), .Z(n365) );
  BUF_X1 U13 ( .A(N10), .Z(n366) );
  BUF_X1 U14 ( .A(N11), .Z(n363) );
  NOR2_X1 U15 ( .A1(n377), .A2(N12), .ZN(n642) );
  INV_X1 U16 ( .A(wr_en), .ZN(n377) );
  AND2_X1 U17 ( .A1(N12), .A2(wr_en), .ZN(n573) );
  OAI21_X1 U18 ( .B1(n386), .B2(n607), .A(n599), .ZN(n466) );
  NAND2_X1 U19 ( .A1(\mem[3][7] ), .A2(n371), .ZN(n599) );
  OAI21_X1 U20 ( .B1(n385), .B2(n371), .A(n598), .ZN(n465) );
  NAND2_X1 U21 ( .A1(\mem[3][8] ), .A2(n371), .ZN(n598) );
  OAI21_X1 U22 ( .B1(n384), .B2(n607), .A(n597), .ZN(n464) );
  NAND2_X1 U23 ( .A1(\mem[3][9] ), .A2(n371), .ZN(n597) );
  OAI21_X1 U24 ( .B1(n383), .B2(n607), .A(n596), .ZN(n463) );
  NAND2_X1 U25 ( .A1(\mem[3][10] ), .A2(n371), .ZN(n596) );
  OAI21_X1 U26 ( .B1(n382), .B2(n607), .A(n595), .ZN(n462) );
  NAND2_X1 U27 ( .A1(\mem[3][11] ), .A2(n371), .ZN(n595) );
  OAI21_X1 U28 ( .B1(n381), .B2(n607), .A(n594), .ZN(n461) );
  NAND2_X1 U29 ( .A1(\mem[3][12] ), .A2(n371), .ZN(n594) );
  OAI21_X1 U30 ( .B1(n380), .B2(n607), .A(n593), .ZN(n460) );
  NAND2_X1 U31 ( .A1(\mem[3][13] ), .A2(n371), .ZN(n593) );
  OAI21_X1 U32 ( .B1(n379), .B2(n607), .A(n592), .ZN(n459) );
  NAND2_X1 U33 ( .A1(\mem[3][14] ), .A2(n371), .ZN(n592) );
  OAI21_X1 U34 ( .B1(n386), .B2(n572), .A(n564), .ZN(n434) );
  NAND2_X1 U35 ( .A1(\mem[5][7] ), .A2(n369), .ZN(n564) );
  OAI21_X1 U36 ( .B1(n385), .B2(n369), .A(n563), .ZN(n433) );
  NAND2_X1 U37 ( .A1(\mem[5][8] ), .A2(n369), .ZN(n563) );
  OAI21_X1 U38 ( .B1(n384), .B2(n572), .A(n562), .ZN(n432) );
  NAND2_X1 U39 ( .A1(\mem[5][9] ), .A2(n369), .ZN(n562) );
  OAI21_X1 U40 ( .B1(n383), .B2(n572), .A(n561), .ZN(n431) );
  NAND2_X1 U41 ( .A1(\mem[5][10] ), .A2(n369), .ZN(n561) );
  OAI21_X1 U42 ( .B1(n382), .B2(n572), .A(n560), .ZN(n430) );
  NAND2_X1 U43 ( .A1(\mem[5][11] ), .A2(n369), .ZN(n560) );
  OAI21_X1 U44 ( .B1(n381), .B2(n572), .A(n559), .ZN(n429) );
  NAND2_X1 U45 ( .A1(\mem[5][12] ), .A2(n369), .ZN(n559) );
  OAI21_X1 U46 ( .B1(n380), .B2(n572), .A(n558), .ZN(n428) );
  NAND2_X1 U47 ( .A1(\mem[5][13] ), .A2(n369), .ZN(n558) );
  OAI21_X1 U48 ( .B1(n379), .B2(n572), .A(n557), .ZN(n427) );
  NAND2_X1 U49 ( .A1(\mem[5][14] ), .A2(n369), .ZN(n557) );
  OAI21_X1 U50 ( .B1(n386), .B2(n538), .A(n530), .ZN(n402) );
  NAND2_X1 U51 ( .A1(\mem[7][7] ), .A2(n367), .ZN(n530) );
  OAI21_X1 U52 ( .B1(n385), .B2(n367), .A(n529), .ZN(n401) );
  NAND2_X1 U53 ( .A1(\mem[7][8] ), .A2(n367), .ZN(n529) );
  OAI21_X1 U54 ( .B1(n384), .B2(n538), .A(n528), .ZN(n400) );
  NAND2_X1 U55 ( .A1(\mem[7][9] ), .A2(n367), .ZN(n528) );
  OAI21_X1 U56 ( .B1(n383), .B2(n538), .A(n527), .ZN(n399) );
  NAND2_X1 U57 ( .A1(\mem[7][10] ), .A2(n367), .ZN(n527) );
  OAI21_X1 U58 ( .B1(n382), .B2(n538), .A(n526), .ZN(n398) );
  NAND2_X1 U59 ( .A1(\mem[7][11] ), .A2(n367), .ZN(n526) );
  OAI21_X1 U60 ( .B1(n381), .B2(n538), .A(n525), .ZN(n397) );
  NAND2_X1 U61 ( .A1(\mem[7][12] ), .A2(n367), .ZN(n525) );
  OAI21_X1 U62 ( .B1(n380), .B2(n538), .A(n524), .ZN(n396) );
  NAND2_X1 U63 ( .A1(\mem[7][13] ), .A2(n367), .ZN(n524) );
  OAI21_X1 U64 ( .B1(n379), .B2(n538), .A(n523), .ZN(n395) );
  NAND2_X1 U65 ( .A1(\mem[7][14] ), .A2(n367), .ZN(n523) );
  OAI21_X1 U66 ( .B1(n386), .B2(n555), .A(n547), .ZN(n418) );
  NAND2_X1 U67 ( .A1(\mem[6][7] ), .A2(n368), .ZN(n547) );
  OAI21_X1 U68 ( .B1(n385), .B2(n368), .A(n546), .ZN(n417) );
  NAND2_X1 U69 ( .A1(\mem[6][8] ), .A2(n368), .ZN(n546) );
  OAI21_X1 U70 ( .B1(n384), .B2(n555), .A(n545), .ZN(n416) );
  NAND2_X1 U71 ( .A1(\mem[6][9] ), .A2(n368), .ZN(n545) );
  OAI21_X1 U72 ( .B1(n383), .B2(n555), .A(n544), .ZN(n415) );
  NAND2_X1 U73 ( .A1(\mem[6][10] ), .A2(n368), .ZN(n544) );
  OAI21_X1 U74 ( .B1(n382), .B2(n555), .A(n543), .ZN(n414) );
  NAND2_X1 U75 ( .A1(\mem[6][11] ), .A2(n368), .ZN(n543) );
  OAI21_X1 U76 ( .B1(n381), .B2(n555), .A(n542), .ZN(n413) );
  NAND2_X1 U77 ( .A1(\mem[6][12] ), .A2(n368), .ZN(n542) );
  OAI21_X1 U78 ( .B1(n380), .B2(n555), .A(n541), .ZN(n412) );
  NAND2_X1 U79 ( .A1(\mem[6][13] ), .A2(n368), .ZN(n541) );
  OAI21_X1 U80 ( .B1(n379), .B2(n555), .A(n540), .ZN(n411) );
  NAND2_X1 U81 ( .A1(\mem[6][14] ), .A2(n368), .ZN(n540) );
  OAI21_X1 U82 ( .B1(n386), .B2(n641), .A(n633), .ZN(n498) );
  NAND2_X1 U83 ( .A1(\mem[1][7] ), .A2(n373), .ZN(n633) );
  OAI21_X1 U84 ( .B1(n385), .B2(n373), .A(n632), .ZN(n497) );
  NAND2_X1 U85 ( .A1(\mem[1][8] ), .A2(n373), .ZN(n632) );
  OAI21_X1 U86 ( .B1(n384), .B2(n641), .A(n631), .ZN(n496) );
  NAND2_X1 U87 ( .A1(\mem[1][9] ), .A2(n373), .ZN(n631) );
  OAI21_X1 U88 ( .B1(n383), .B2(n641), .A(n630), .ZN(n495) );
  NAND2_X1 U89 ( .A1(\mem[1][10] ), .A2(n373), .ZN(n630) );
  OAI21_X1 U90 ( .B1(n382), .B2(n641), .A(n629), .ZN(n494) );
  NAND2_X1 U91 ( .A1(\mem[1][11] ), .A2(n373), .ZN(n629) );
  OAI21_X1 U92 ( .B1(n381), .B2(n641), .A(n628), .ZN(n493) );
  NAND2_X1 U93 ( .A1(\mem[1][12] ), .A2(n373), .ZN(n628) );
  OAI21_X1 U94 ( .B1(n380), .B2(n641), .A(n627), .ZN(n492) );
  NAND2_X1 U95 ( .A1(\mem[1][13] ), .A2(n373), .ZN(n627) );
  OAI21_X1 U96 ( .B1(n379), .B2(n641), .A(n626), .ZN(n491) );
  NAND2_X1 U97 ( .A1(\mem[1][14] ), .A2(n373), .ZN(n626) );
  OAI21_X1 U98 ( .B1(n386), .B2(n624), .A(n616), .ZN(n482) );
  NAND2_X1 U99 ( .A1(\mem[2][7] ), .A2(n372), .ZN(n616) );
  OAI21_X1 U100 ( .B1(n385), .B2(n372), .A(n615), .ZN(n481) );
  NAND2_X1 U101 ( .A1(\mem[2][8] ), .A2(n372), .ZN(n615) );
  OAI21_X1 U102 ( .B1(n384), .B2(n624), .A(n614), .ZN(n480) );
  NAND2_X1 U103 ( .A1(\mem[2][9] ), .A2(n372), .ZN(n614) );
  OAI21_X1 U104 ( .B1(n383), .B2(n624), .A(n613), .ZN(n479) );
  NAND2_X1 U105 ( .A1(\mem[2][10] ), .A2(n372), .ZN(n613) );
  OAI21_X1 U106 ( .B1(n382), .B2(n624), .A(n612), .ZN(n478) );
  NAND2_X1 U107 ( .A1(\mem[2][11] ), .A2(n372), .ZN(n612) );
  OAI21_X1 U108 ( .B1(n381), .B2(n624), .A(n611), .ZN(n477) );
  NAND2_X1 U109 ( .A1(\mem[2][12] ), .A2(n372), .ZN(n611) );
  OAI21_X1 U110 ( .B1(n380), .B2(n624), .A(n610), .ZN(n476) );
  NAND2_X1 U111 ( .A1(\mem[2][13] ), .A2(n372), .ZN(n610) );
  OAI21_X1 U112 ( .B1(n379), .B2(n624), .A(n609), .ZN(n475) );
  NAND2_X1 U113 ( .A1(\mem[2][14] ), .A2(n372), .ZN(n609) );
  OAI21_X1 U114 ( .B1(n386), .B2(n590), .A(n582), .ZN(n450) );
  NAND2_X1 U115 ( .A1(\mem[4][7] ), .A2(n370), .ZN(n582) );
  OAI21_X1 U116 ( .B1(n385), .B2(n370), .A(n581), .ZN(n449) );
  NAND2_X1 U117 ( .A1(\mem[4][8] ), .A2(n370), .ZN(n581) );
  OAI21_X1 U118 ( .B1(n384), .B2(n590), .A(n580), .ZN(n448) );
  NAND2_X1 U119 ( .A1(\mem[4][9] ), .A2(n370), .ZN(n580) );
  OAI21_X1 U120 ( .B1(n383), .B2(n590), .A(n579), .ZN(n447) );
  NAND2_X1 U121 ( .A1(\mem[4][10] ), .A2(n370), .ZN(n579) );
  OAI21_X1 U122 ( .B1(n382), .B2(n590), .A(n578), .ZN(n446) );
  NAND2_X1 U123 ( .A1(\mem[4][11] ), .A2(n370), .ZN(n578) );
  OAI21_X1 U124 ( .B1(n381), .B2(n590), .A(n577), .ZN(n445) );
  NAND2_X1 U125 ( .A1(\mem[4][12] ), .A2(n370), .ZN(n577) );
  OAI21_X1 U126 ( .B1(n380), .B2(n590), .A(n576), .ZN(n444) );
  NAND2_X1 U127 ( .A1(\mem[4][13] ), .A2(n370), .ZN(n576) );
  OAI21_X1 U128 ( .B1(n379), .B2(n590), .A(n575), .ZN(n443) );
  NAND2_X1 U129 ( .A1(\mem[4][14] ), .A2(n370), .ZN(n575) );
  INV_X1 U130 ( .A(N10), .ZN(n375) );
  OAI21_X1 U131 ( .B1(n659), .B2(n385), .A(n650), .ZN(n513) );
  NAND2_X1 U132 ( .A1(\mem[0][8] ), .A2(n374), .ZN(n650) );
  OAI21_X1 U133 ( .B1(n659), .B2(n384), .A(n649), .ZN(n512) );
  NAND2_X1 U134 ( .A1(\mem[0][9] ), .A2(n659), .ZN(n649) );
  OAI21_X1 U135 ( .B1(n374), .B2(n383), .A(n648), .ZN(n511) );
  NAND2_X1 U136 ( .A1(\mem[0][10] ), .A2(n659), .ZN(n648) );
  OAI21_X1 U137 ( .B1(n659), .B2(n382), .A(n647), .ZN(n510) );
  NAND2_X1 U138 ( .A1(\mem[0][11] ), .A2(n659), .ZN(n647) );
  OAI21_X1 U139 ( .B1(n659), .B2(n381), .A(n646), .ZN(n509) );
  NAND2_X1 U140 ( .A1(\mem[0][12] ), .A2(n659), .ZN(n646) );
  OAI21_X1 U141 ( .B1(n659), .B2(n380), .A(n645), .ZN(n508) );
  NAND2_X1 U142 ( .A1(\mem[0][13] ), .A2(n659), .ZN(n645) );
  OAI21_X1 U143 ( .B1(n659), .B2(n379), .A(n644), .ZN(n507) );
  NAND2_X1 U144 ( .A1(\mem[0][14] ), .A2(n659), .ZN(n644) );
  OAI21_X1 U145 ( .B1(n393), .B2(n641), .A(n640), .ZN(n505) );
  NAND2_X1 U146 ( .A1(\mem[1][0] ), .A2(n373), .ZN(n640) );
  OAI21_X1 U147 ( .B1(n392), .B2(n641), .A(n639), .ZN(n504) );
  NAND2_X1 U148 ( .A1(\mem[1][1] ), .A2(n373), .ZN(n639) );
  OAI21_X1 U149 ( .B1(n391), .B2(n641), .A(n638), .ZN(n503) );
  NAND2_X1 U150 ( .A1(\mem[1][2] ), .A2(n373), .ZN(n638) );
  OAI21_X1 U151 ( .B1(n390), .B2(n641), .A(n637), .ZN(n502) );
  NAND2_X1 U152 ( .A1(\mem[1][3] ), .A2(n373), .ZN(n637) );
  OAI21_X1 U153 ( .B1(n389), .B2(n641), .A(n636), .ZN(n501) );
  NAND2_X1 U154 ( .A1(\mem[1][4] ), .A2(n641), .ZN(n636) );
  OAI21_X1 U155 ( .B1(n388), .B2(n641), .A(n635), .ZN(n500) );
  NAND2_X1 U156 ( .A1(\mem[1][5] ), .A2(n641), .ZN(n635) );
  OAI21_X1 U157 ( .B1(n387), .B2(n641), .A(n634), .ZN(n499) );
  NAND2_X1 U158 ( .A1(\mem[1][6] ), .A2(n641), .ZN(n634) );
  OAI21_X1 U159 ( .B1(n378), .B2(n641), .A(n625), .ZN(n490) );
  NAND2_X1 U160 ( .A1(\mem[1][15] ), .A2(n373), .ZN(n625) );
  OAI21_X1 U161 ( .B1(n393), .B2(n624), .A(n623), .ZN(n489) );
  NAND2_X1 U162 ( .A1(\mem[2][0] ), .A2(n372), .ZN(n623) );
  OAI21_X1 U163 ( .B1(n392), .B2(n624), .A(n622), .ZN(n488) );
  NAND2_X1 U164 ( .A1(\mem[2][1] ), .A2(n372), .ZN(n622) );
  OAI21_X1 U165 ( .B1(n391), .B2(n624), .A(n621), .ZN(n487) );
  NAND2_X1 U166 ( .A1(\mem[2][2] ), .A2(n372), .ZN(n621) );
  OAI21_X1 U167 ( .B1(n390), .B2(n624), .A(n620), .ZN(n486) );
  NAND2_X1 U168 ( .A1(\mem[2][3] ), .A2(n372), .ZN(n620) );
  OAI21_X1 U169 ( .B1(n389), .B2(n624), .A(n619), .ZN(n485) );
  NAND2_X1 U170 ( .A1(\mem[2][4] ), .A2(n624), .ZN(n619) );
  OAI21_X1 U171 ( .B1(n388), .B2(n624), .A(n618), .ZN(n484) );
  NAND2_X1 U172 ( .A1(\mem[2][5] ), .A2(n624), .ZN(n618) );
  OAI21_X1 U173 ( .B1(n387), .B2(n624), .A(n617), .ZN(n483) );
  NAND2_X1 U174 ( .A1(\mem[2][6] ), .A2(n624), .ZN(n617) );
  OAI21_X1 U175 ( .B1(n378), .B2(n624), .A(n608), .ZN(n474) );
  NAND2_X1 U176 ( .A1(\mem[2][15] ), .A2(n372), .ZN(n608) );
  OAI21_X1 U177 ( .B1(n393), .B2(n607), .A(n606), .ZN(n473) );
  NAND2_X1 U178 ( .A1(\mem[3][0] ), .A2(n371), .ZN(n606) );
  OAI21_X1 U179 ( .B1(n392), .B2(n607), .A(n605), .ZN(n472) );
  NAND2_X1 U180 ( .A1(\mem[3][1] ), .A2(n371), .ZN(n605) );
  OAI21_X1 U181 ( .B1(n391), .B2(n607), .A(n604), .ZN(n471) );
  NAND2_X1 U182 ( .A1(\mem[3][2] ), .A2(n371), .ZN(n604) );
  OAI21_X1 U183 ( .B1(n390), .B2(n607), .A(n603), .ZN(n470) );
  NAND2_X1 U184 ( .A1(\mem[3][3] ), .A2(n371), .ZN(n603) );
  OAI21_X1 U185 ( .B1(n389), .B2(n607), .A(n602), .ZN(n469) );
  NAND2_X1 U186 ( .A1(\mem[3][4] ), .A2(n607), .ZN(n602) );
  OAI21_X1 U187 ( .B1(n388), .B2(n607), .A(n601), .ZN(n468) );
  NAND2_X1 U188 ( .A1(\mem[3][5] ), .A2(n607), .ZN(n601) );
  OAI21_X1 U189 ( .B1(n387), .B2(n607), .A(n600), .ZN(n467) );
  NAND2_X1 U190 ( .A1(\mem[3][6] ), .A2(n607), .ZN(n600) );
  OAI21_X1 U191 ( .B1(n378), .B2(n607), .A(n591), .ZN(n458) );
  NAND2_X1 U192 ( .A1(\mem[3][15] ), .A2(n371), .ZN(n591) );
  OAI21_X1 U193 ( .B1(n393), .B2(n590), .A(n589), .ZN(n457) );
  NAND2_X1 U194 ( .A1(\mem[4][0] ), .A2(n370), .ZN(n589) );
  OAI21_X1 U195 ( .B1(n392), .B2(n590), .A(n588), .ZN(n456) );
  NAND2_X1 U196 ( .A1(\mem[4][1] ), .A2(n370), .ZN(n588) );
  OAI21_X1 U197 ( .B1(n391), .B2(n590), .A(n587), .ZN(n455) );
  NAND2_X1 U198 ( .A1(\mem[4][2] ), .A2(n370), .ZN(n587) );
  OAI21_X1 U199 ( .B1(n390), .B2(n590), .A(n586), .ZN(n454) );
  NAND2_X1 U200 ( .A1(\mem[4][3] ), .A2(n370), .ZN(n586) );
  OAI21_X1 U201 ( .B1(n389), .B2(n590), .A(n585), .ZN(n453) );
  NAND2_X1 U202 ( .A1(\mem[4][4] ), .A2(n590), .ZN(n585) );
  OAI21_X1 U203 ( .B1(n388), .B2(n590), .A(n584), .ZN(n452) );
  NAND2_X1 U204 ( .A1(\mem[4][5] ), .A2(n590), .ZN(n584) );
  OAI21_X1 U205 ( .B1(n387), .B2(n590), .A(n583), .ZN(n451) );
  NAND2_X1 U206 ( .A1(\mem[4][6] ), .A2(n590), .ZN(n583) );
  OAI21_X1 U207 ( .B1(n378), .B2(n590), .A(n574), .ZN(n442) );
  NAND2_X1 U208 ( .A1(\mem[4][15] ), .A2(n370), .ZN(n574) );
  OAI21_X1 U209 ( .B1(n393), .B2(n572), .A(n571), .ZN(n441) );
  NAND2_X1 U210 ( .A1(\mem[5][0] ), .A2(n369), .ZN(n571) );
  OAI21_X1 U211 ( .B1(n392), .B2(n572), .A(n570), .ZN(n440) );
  NAND2_X1 U212 ( .A1(\mem[5][1] ), .A2(n369), .ZN(n570) );
  OAI21_X1 U213 ( .B1(n391), .B2(n572), .A(n569), .ZN(n439) );
  NAND2_X1 U214 ( .A1(\mem[5][2] ), .A2(n369), .ZN(n569) );
  OAI21_X1 U215 ( .B1(n390), .B2(n572), .A(n568), .ZN(n438) );
  NAND2_X1 U216 ( .A1(\mem[5][3] ), .A2(n369), .ZN(n568) );
  OAI21_X1 U217 ( .B1(n389), .B2(n572), .A(n567), .ZN(n437) );
  NAND2_X1 U218 ( .A1(\mem[5][4] ), .A2(n572), .ZN(n567) );
  OAI21_X1 U219 ( .B1(n388), .B2(n572), .A(n566), .ZN(n436) );
  NAND2_X1 U220 ( .A1(\mem[5][5] ), .A2(n572), .ZN(n566) );
  OAI21_X1 U221 ( .B1(n387), .B2(n572), .A(n565), .ZN(n435) );
  NAND2_X1 U222 ( .A1(\mem[5][6] ), .A2(n572), .ZN(n565) );
  OAI21_X1 U223 ( .B1(n378), .B2(n572), .A(n556), .ZN(n426) );
  NAND2_X1 U224 ( .A1(\mem[5][15] ), .A2(n369), .ZN(n556) );
  OAI21_X1 U225 ( .B1(n393), .B2(n555), .A(n554), .ZN(n425) );
  NAND2_X1 U226 ( .A1(\mem[6][0] ), .A2(n368), .ZN(n554) );
  OAI21_X1 U227 ( .B1(n392), .B2(n555), .A(n553), .ZN(n424) );
  NAND2_X1 U228 ( .A1(\mem[6][1] ), .A2(n368), .ZN(n553) );
  OAI21_X1 U229 ( .B1(n391), .B2(n555), .A(n552), .ZN(n423) );
  NAND2_X1 U230 ( .A1(\mem[6][2] ), .A2(n368), .ZN(n552) );
  OAI21_X1 U231 ( .B1(n390), .B2(n555), .A(n551), .ZN(n422) );
  NAND2_X1 U232 ( .A1(\mem[6][3] ), .A2(n368), .ZN(n551) );
  OAI21_X1 U233 ( .B1(n389), .B2(n555), .A(n550), .ZN(n421) );
  NAND2_X1 U234 ( .A1(\mem[6][4] ), .A2(n555), .ZN(n550) );
  OAI21_X1 U235 ( .B1(n388), .B2(n555), .A(n549), .ZN(n420) );
  NAND2_X1 U236 ( .A1(\mem[6][5] ), .A2(n555), .ZN(n549) );
  OAI21_X1 U237 ( .B1(n387), .B2(n555), .A(n548), .ZN(n419) );
  NAND2_X1 U238 ( .A1(\mem[6][6] ), .A2(n555), .ZN(n548) );
  OAI21_X1 U239 ( .B1(n378), .B2(n555), .A(n539), .ZN(n410) );
  NAND2_X1 U240 ( .A1(\mem[6][15] ), .A2(n368), .ZN(n539) );
  OAI21_X1 U241 ( .B1(n393), .B2(n538), .A(n537), .ZN(n409) );
  NAND2_X1 U242 ( .A1(\mem[7][0] ), .A2(n367), .ZN(n537) );
  OAI21_X1 U243 ( .B1(n392), .B2(n538), .A(n536), .ZN(n408) );
  NAND2_X1 U244 ( .A1(\mem[7][1] ), .A2(n367), .ZN(n536) );
  OAI21_X1 U245 ( .B1(n391), .B2(n538), .A(n535), .ZN(n407) );
  NAND2_X1 U246 ( .A1(\mem[7][2] ), .A2(n367), .ZN(n535) );
  OAI21_X1 U247 ( .B1(n390), .B2(n538), .A(n534), .ZN(n406) );
  NAND2_X1 U248 ( .A1(\mem[7][3] ), .A2(n367), .ZN(n534) );
  OAI21_X1 U249 ( .B1(n389), .B2(n538), .A(n533), .ZN(n405) );
  NAND2_X1 U250 ( .A1(\mem[7][4] ), .A2(n538), .ZN(n533) );
  OAI21_X1 U251 ( .B1(n388), .B2(n538), .A(n532), .ZN(n404) );
  NAND2_X1 U252 ( .A1(\mem[7][5] ), .A2(n538), .ZN(n532) );
  OAI21_X1 U253 ( .B1(n387), .B2(n538), .A(n531), .ZN(n403) );
  NAND2_X1 U254 ( .A1(\mem[7][6] ), .A2(n538), .ZN(n531) );
  OAI21_X1 U255 ( .B1(n378), .B2(n538), .A(n522), .ZN(n394) );
  NAND2_X1 U256 ( .A1(\mem[7][15] ), .A2(n367), .ZN(n522) );
  OAI21_X1 U257 ( .B1(n374), .B2(n393), .A(n658), .ZN(n521) );
  NAND2_X1 U258 ( .A1(\mem[0][0] ), .A2(n659), .ZN(n658) );
  OAI21_X1 U259 ( .B1(n374), .B2(n392), .A(n657), .ZN(n520) );
  NAND2_X1 U260 ( .A1(\mem[0][1] ), .A2(n659), .ZN(n657) );
  OAI21_X1 U261 ( .B1(n374), .B2(n391), .A(n656), .ZN(n519) );
  NAND2_X1 U262 ( .A1(\mem[0][2] ), .A2(n659), .ZN(n656) );
  OAI21_X1 U263 ( .B1(n374), .B2(n390), .A(n655), .ZN(n518) );
  NAND2_X1 U264 ( .A1(\mem[0][3] ), .A2(n659), .ZN(n655) );
  OAI21_X1 U265 ( .B1(n374), .B2(n389), .A(n654), .ZN(n517) );
  NAND2_X1 U266 ( .A1(\mem[0][4] ), .A2(n374), .ZN(n654) );
  OAI21_X1 U267 ( .B1(n374), .B2(n388), .A(n653), .ZN(n516) );
  NAND2_X1 U268 ( .A1(\mem[0][5] ), .A2(n374), .ZN(n653) );
  OAI21_X1 U269 ( .B1(n374), .B2(n387), .A(n652), .ZN(n515) );
  NAND2_X1 U270 ( .A1(\mem[0][6] ), .A2(n374), .ZN(n652) );
  OAI21_X1 U271 ( .B1(n374), .B2(n386), .A(n651), .ZN(n514) );
  NAND2_X1 U272 ( .A1(\mem[0][7] ), .A2(n374), .ZN(n651) );
  OAI21_X1 U273 ( .B1(n374), .B2(n378), .A(n643), .ZN(n506) );
  NAND2_X1 U274 ( .A1(\mem[0][15] ), .A2(n659), .ZN(n643) );
  INV_X1 U275 ( .A(N11), .ZN(n376) );
  INV_X1 U276 ( .A(data_in[0]), .ZN(n393) );
  INV_X1 U277 ( .A(data_in[1]), .ZN(n392) );
  INV_X1 U278 ( .A(data_in[2]), .ZN(n391) );
  INV_X1 U279 ( .A(data_in[3]), .ZN(n390) );
  INV_X1 U288 ( .A(data_in[4]), .ZN(n389) );
  INV_X1 U289 ( .A(data_in[5]), .ZN(n388) );
  INV_X1 U290 ( .A(data_in[6]), .ZN(n387) );
  INV_X1 U291 ( .A(data_in[7]), .ZN(n386) );
  INV_X1 U292 ( .A(data_in[8]), .ZN(n385) );
  INV_X1 U293 ( .A(data_in[9]), .ZN(n384) );
  INV_X1 U294 ( .A(data_in[10]), .ZN(n383) );
  INV_X1 U295 ( .A(data_in[11]), .ZN(n382) );
  INV_X1 U296 ( .A(data_in[12]), .ZN(n381) );
  INV_X1 U297 ( .A(data_in[13]), .ZN(n380) );
  INV_X1 U298 ( .A(data_in[14]), .ZN(n379) );
  INV_X1 U299 ( .A(data_in[15]), .ZN(n378) );
  MUX2_X1 U300 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n366), .Z(n1) );
  MUX2_X1 U301 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n365), .Z(n2) );
  MUX2_X1 U302 ( .A(n2), .B(n1), .S(n363), .Z(n3) );
  MUX2_X1 U303 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n366), .Z(n4) );
  MUX2_X1 U304 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n364), .Z(n5) );
  MUX2_X1 U305 ( .A(n5), .B(n4), .S(N11), .Z(n6) );
  MUX2_X1 U306 ( .A(n6), .B(n3), .S(N12), .Z(N28) );
  MUX2_X1 U307 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n364), .Z(n7) );
  MUX2_X1 U308 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n364), .Z(n8) );
  MUX2_X1 U309 ( .A(n8), .B(n7), .S(n363), .Z(n9) );
  MUX2_X1 U310 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n364), .Z(n10) );
  MUX2_X1 U311 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n364), .Z(n11) );
  MUX2_X1 U312 ( .A(n11), .B(n10), .S(N11), .Z(n12) );
  MUX2_X1 U313 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n364), .Z(n13) );
  MUX2_X1 U314 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n364), .Z(n14) );
  MUX2_X1 U315 ( .A(n14), .B(n13), .S(N11), .Z(n15) );
  MUX2_X1 U316 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n364), .Z(n16) );
  MUX2_X1 U317 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n364), .Z(n17) );
  MUX2_X1 U318 ( .A(n17), .B(n16), .S(n363), .Z(n18) );
  MUX2_X1 U319 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n364), .Z(n19) );
  MUX2_X1 U320 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n364), .Z(n286) );
  MUX2_X1 U321 ( .A(n286), .B(n19), .S(n363), .Z(n287) );
  MUX2_X1 U322 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n364), .Z(n288) );
  MUX2_X1 U323 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n364), .Z(n289) );
  MUX2_X1 U324 ( .A(n289), .B(n288), .S(N11), .Z(n290) );
  MUX2_X1 U325 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n365), .Z(n291) );
  MUX2_X1 U326 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n365), .Z(n292) );
  MUX2_X1 U327 ( .A(n292), .B(n291), .S(n363), .Z(n293) );
  MUX2_X1 U328 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n365), .Z(n294) );
  MUX2_X1 U329 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n365), .Z(n295) );
  MUX2_X1 U330 ( .A(n295), .B(n294), .S(n363), .Z(n296) );
  MUX2_X1 U331 ( .A(n296), .B(n293), .S(N12), .Z(N24) );
  MUX2_X1 U332 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n365), .Z(n297) );
  MUX2_X1 U333 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n365), .Z(n298) );
  MUX2_X1 U334 ( .A(n298), .B(n297), .S(n363), .Z(n299) );
  MUX2_X1 U335 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n365), .Z(n300) );
  MUX2_X1 U336 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n365), .Z(n301) );
  MUX2_X1 U337 ( .A(n301), .B(n300), .S(n363), .Z(n302) );
  MUX2_X1 U338 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n365), .Z(n303) );
  MUX2_X1 U339 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n365), .Z(n304) );
  MUX2_X1 U340 ( .A(n304), .B(n303), .S(n363), .Z(n305) );
  MUX2_X1 U341 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n365), .Z(n306) );
  MUX2_X1 U342 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n365), .Z(n307) );
  MUX2_X1 U343 ( .A(n307), .B(n306), .S(n363), .Z(n308) );
  MUX2_X1 U344 ( .A(n308), .B(n305), .S(N12), .Z(N22) );
  MUX2_X1 U345 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n366), .Z(n309) );
  MUX2_X1 U346 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n366), .Z(n310) );
  MUX2_X1 U347 ( .A(n310), .B(n309), .S(n363), .Z(n311) );
  MUX2_X1 U348 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n366), .Z(n312) );
  MUX2_X1 U349 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n366), .Z(n313) );
  MUX2_X1 U350 ( .A(n313), .B(n312), .S(n363), .Z(n314) );
  MUX2_X1 U351 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n366), .Z(n315) );
  MUX2_X1 U352 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n366), .Z(n316) );
  MUX2_X1 U353 ( .A(n316), .B(n315), .S(n363), .Z(n317) );
  MUX2_X1 U354 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n366), .Z(n318) );
  MUX2_X1 U355 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n366), .Z(n319) );
  MUX2_X1 U356 ( .A(n319), .B(n318), .S(n363), .Z(n320) );
  MUX2_X1 U357 ( .A(n320), .B(n317), .S(N12), .Z(N20) );
  MUX2_X1 U358 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n366), .Z(n321) );
  MUX2_X1 U359 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n366), .Z(n322) );
  MUX2_X1 U360 ( .A(n322), .B(n321), .S(n363), .Z(n323) );
  MUX2_X1 U361 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n366), .Z(n324) );
  MUX2_X1 U362 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n366), .Z(n325) );
  MUX2_X1 U363 ( .A(n325), .B(n324), .S(n363), .Z(n326) );
  MUX2_X1 U364 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n364), .Z(n327) );
  MUX2_X1 U365 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n366), .Z(n328) );
  MUX2_X1 U366 ( .A(n328), .B(n327), .S(n363), .Z(n329) );
  MUX2_X1 U367 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n366), .Z(n330) );
  MUX2_X1 U368 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n365), .Z(n331) );
  MUX2_X1 U369 ( .A(n331), .B(n330), .S(n363), .Z(n332) );
  MUX2_X1 U370 ( .A(n332), .B(n329), .S(N12), .Z(N18) );
  MUX2_X1 U371 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n366), .Z(n333) );
  MUX2_X1 U372 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n364), .Z(n334) );
  MUX2_X1 U373 ( .A(n334), .B(n333), .S(N11), .Z(n335) );
  MUX2_X1 U374 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n365), .Z(n336) );
  MUX2_X1 U375 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n366), .Z(n337) );
  MUX2_X1 U376 ( .A(n337), .B(n336), .S(N11), .Z(n338) );
  MUX2_X1 U377 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n365), .Z(n339) );
  MUX2_X1 U378 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n364), .Z(n340) );
  MUX2_X1 U379 ( .A(n340), .B(n339), .S(n363), .Z(n341) );
  MUX2_X1 U380 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n364), .Z(n342) );
  MUX2_X1 U381 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n366), .Z(n343) );
  MUX2_X1 U382 ( .A(n343), .B(n342), .S(n363), .Z(n344) );
  MUX2_X1 U383 ( .A(n344), .B(n341), .S(N12), .Z(N16) );
  MUX2_X1 U384 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n365), .Z(n345) );
  MUX2_X1 U385 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n366), .Z(n346) );
  MUX2_X1 U386 ( .A(n346), .B(n345), .S(N11), .Z(n347) );
  MUX2_X1 U387 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n365), .Z(n348) );
  MUX2_X1 U388 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(N10), .Z(n349) );
  MUX2_X1 U389 ( .A(n349), .B(n348), .S(N11), .Z(n350) );
  MUX2_X1 U390 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n364), .Z(n351) );
  MUX2_X1 U391 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n366), .Z(n352) );
  MUX2_X1 U392 ( .A(n352), .B(n351), .S(n363), .Z(n353) );
  MUX2_X1 U393 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n365), .Z(n354) );
  MUX2_X1 U394 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n364), .Z(n355) );
  MUX2_X1 U395 ( .A(n355), .B(n354), .S(n363), .Z(n356) );
  MUX2_X1 U396 ( .A(n356), .B(n353), .S(N12), .Z(N14) );
  MUX2_X1 U397 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n365), .Z(n357) );
  MUX2_X1 U398 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n364), .Z(n358) );
  MUX2_X1 U399 ( .A(n358), .B(n357), .S(n363), .Z(n359) );
  MUX2_X1 U400 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n365), .Z(n360) );
  MUX2_X1 U401 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n364), .Z(n361) );
  MUX2_X1 U402 ( .A(n361), .B(n360), .S(N11), .Z(n362) );
  MUX2_X1 U403 ( .A(n362), .B(n359), .S(N12), .Z(N13) );
endmodule


module memory_WIDTH32_SIZE8_LOGSIZE3 ( clk, data_in, data_out, addr, wr_en );
  input [31:0] data_in;
  output [31:0] data_out;
  input [2:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, \mem[7][31] , \mem[7][30] , \mem[7][29] , \mem[7][28] ,
         \mem[7][27] , \mem[7][26] , \mem[7][25] , \mem[7][24] , \mem[7][23] ,
         \mem[7][22] , \mem[7][21] , \mem[7][20] , \mem[7][19] , \mem[7][18] ,
         \mem[7][17] , \mem[7][16] , \mem[7][15] , \mem[7][14] , \mem[7][13] ,
         \mem[7][12] , \mem[7][11] , \mem[7][10] , \mem[7][9] , \mem[7][8] ,
         \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] ,
         \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][31] , \mem[6][30] ,
         \mem[6][29] , \mem[6][28] , \mem[6][27] , \mem[6][26] , \mem[6][25] ,
         \mem[6][24] , \mem[6][23] , \mem[6][22] , \mem[6][21] , \mem[6][20] ,
         \mem[6][19] , \mem[6][18] , \mem[6][17] , \mem[6][16] , \mem[6][15] ,
         \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][31] , \mem[5][30] , \mem[5][29] , \mem[5][28] , \mem[5][27] ,
         \mem[5][26] , \mem[5][25] , \mem[5][24] , \mem[5][23] , \mem[5][22] ,
         \mem[5][21] , \mem[5][20] , \mem[5][19] , \mem[5][18] , \mem[5][17] ,
         \mem[5][16] , \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] ,
         \mem[5][11] , \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] ,
         \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] ,
         \mem[5][1] , \mem[5][0] , \mem[4][31] , \mem[4][30] , \mem[4][29] ,
         \mem[4][28] , \mem[4][27] , \mem[4][26] , \mem[4][25] , \mem[4][24] ,
         \mem[4][23] , \mem[4][22] , \mem[4][21] , \mem[4][20] , \mem[4][19] ,
         \mem[4][18] , \mem[4][17] , \mem[4][16] , \mem[4][15] , \mem[4][14] ,
         \mem[4][13] , \mem[4][12] , \mem[4][11] , \mem[4][10] , \mem[4][9] ,
         \mem[4][8] , \mem[4][7] , \mem[4][6] , \mem[4][5] , \mem[4][4] ,
         \mem[4][3] , \mem[4][2] , \mem[4][1] , \mem[4][0] , \mem[3][31] ,
         \mem[3][30] , \mem[3][29] , \mem[3][28] , \mem[3][27] , \mem[3][26] ,
         \mem[3][25] , \mem[3][24] , \mem[3][23] , \mem[3][22] , \mem[3][21] ,
         \mem[3][20] , \mem[3][19] , \mem[3][18] , \mem[3][17] , \mem[3][16] ,
         \mem[3][15] , \mem[3][14] , \mem[3][13] , \mem[3][12] , \mem[3][11] ,
         \mem[3][10] , \mem[3][9] , \mem[3][8] , \mem[3][7] , \mem[3][6] ,
         \mem[3][5] , \mem[3][4] , \mem[3][3] , \mem[3][2] , \mem[3][1] ,
         \mem[3][0] , \mem[2][31] , \mem[2][30] , \mem[2][29] , \mem[2][28] ,
         \mem[2][27] , \mem[2][26] , \mem[2][25] , \mem[2][24] , \mem[2][23] ,
         \mem[2][22] , \mem[2][21] , \mem[2][20] , \mem[2][19] , \mem[2][18] ,
         \mem[2][17] , \mem[2][16] , \mem[2][15] , \mem[2][14] , \mem[2][13] ,
         \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] , \mem[2][8] ,
         \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] ,
         \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][31] , \mem[1][30] ,
         \mem[1][29] , \mem[1][28] , \mem[1][27] , \mem[1][26] , \mem[1][25] ,
         \mem[1][24] , \mem[1][23] , \mem[1][22] , \mem[1][21] , \mem[1][20] ,
         \mem[1][19] , \mem[1][18] , \mem[1][17] , \mem[1][16] , \mem[1][15] ,
         \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][31] , \mem[0][30] , \mem[0][29] , \mem[0][28] , \mem[0][27] ,
         \mem[0][26] , \mem[0][25] , \mem[0][24] , \mem[0][23] , \mem[0][22] ,
         \mem[0][21] , \mem[0][20] , \mem[0][19] , \mem[0][18] , \mem[0][17] ,
         \mem[0][16] , \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] ,
         \mem[0][11] , \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] ,
         \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] ,
         \mem[0][1] , \mem[0][0] , N13, N14, N15, N16, N17, N18, N19, N20, N21,
         N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35,
         N36, N37, N38, N39, N40, N41, N42, N43, N44, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];

  DFF_X1 \data_out_reg[31]  ( .D(N13), .CK(clk), .Q(data_out[31]) );
  DFF_X1 \data_out_reg[30]  ( .D(N14), .CK(clk), .Q(data_out[30]) );
  DFF_X1 \data_out_reg[29]  ( .D(N15), .CK(clk), .Q(data_out[29]) );
  DFF_X1 \data_out_reg[28]  ( .D(N16), .CK(clk), .Q(data_out[28]) );
  DFF_X1 \data_out_reg[27]  ( .D(N17), .CK(clk), .Q(data_out[27]) );
  DFF_X1 \data_out_reg[26]  ( .D(N18), .CK(clk), .Q(data_out[26]) );
  DFF_X1 \data_out_reg[25]  ( .D(N19), .CK(clk), .Q(data_out[25]) );
  DFF_X1 \data_out_reg[24]  ( .D(N20), .CK(clk), .Q(data_out[24]) );
  DFF_X1 \data_out_reg[23]  ( .D(N21), .CK(clk), .Q(data_out[23]) );
  DFF_X1 \data_out_reg[22]  ( .D(N22), .CK(clk), .Q(data_out[22]) );
  DFF_X1 \data_out_reg[21]  ( .D(N23), .CK(clk), .Q(data_out[21]) );
  DFF_X1 \data_out_reg[20]  ( .D(N24), .CK(clk), .Q(data_out[20]) );
  DFF_X1 \data_out_reg[19]  ( .D(N25), .CK(clk), .Q(data_out[19]) );
  DFF_X1 \data_out_reg[18]  ( .D(N26), .CK(clk), .Q(data_out[18]) );
  DFF_X1 \data_out_reg[17]  ( .D(N27), .CK(clk), .Q(data_out[17]) );
  DFF_X1 \data_out_reg[16]  ( .D(N28), .CK(clk), .Q(data_out[16]) );
  DFF_X1 \data_out_reg[15]  ( .D(N29), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N30), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(N31), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(N32), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(N33), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N34), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N35), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N36), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N37), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N38), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N39), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N40), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N41), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N42), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N43), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N44), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[7][31]  ( .D(n557), .CK(clk), .Q(\mem[7][31] ) );
  DFF_X1 \mem_reg[7][30]  ( .D(n556), .CK(clk), .Q(\mem[7][30] ) );
  DFF_X1 \mem_reg[7][29]  ( .D(n555), .CK(clk), .Q(\mem[7][29] ) );
  DFF_X1 \mem_reg[7][28]  ( .D(n554), .CK(clk), .Q(\mem[7][28] ) );
  DFF_X1 \mem_reg[7][27]  ( .D(n553), .CK(clk), .Q(\mem[7][27] ) );
  DFF_X1 \mem_reg[7][26]  ( .D(n552), .CK(clk), .Q(\mem[7][26] ) );
  DFF_X1 \mem_reg[7][25]  ( .D(n551), .CK(clk), .Q(\mem[7][25] ) );
  DFF_X1 \mem_reg[7][24]  ( .D(n550), .CK(clk), .Q(\mem[7][24] ) );
  DFF_X1 \mem_reg[7][23]  ( .D(n549), .CK(clk), .Q(\mem[7][23] ) );
  DFF_X1 \mem_reg[7][22]  ( .D(n548), .CK(clk), .Q(\mem[7][22] ) );
  DFF_X1 \mem_reg[7][21]  ( .D(n547), .CK(clk), .Q(\mem[7][21] ) );
  DFF_X1 \mem_reg[7][20]  ( .D(n546), .CK(clk), .Q(\mem[7][20] ) );
  DFF_X1 \mem_reg[7][19]  ( .D(n545), .CK(clk), .Q(\mem[7][19] ) );
  DFF_X1 \mem_reg[7][18]  ( .D(n544), .CK(clk), .Q(\mem[7][18] ) );
  DFF_X1 \mem_reg[7][17]  ( .D(n543), .CK(clk), .Q(\mem[7][17] ) );
  DFF_X1 \mem_reg[7][16]  ( .D(n542), .CK(clk), .Q(\mem[7][16] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n541), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n540), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n539), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n538), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n537), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n536), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n535), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n534), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n533), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n532), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n531), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n530), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n529), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n528), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n527), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n526), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][31]  ( .D(n525), .CK(clk), .Q(\mem[6][31] ) );
  DFF_X1 \mem_reg[6][30]  ( .D(n524), .CK(clk), .Q(\mem[6][30] ) );
  DFF_X1 \mem_reg[6][29]  ( .D(n523), .CK(clk), .Q(\mem[6][29] ) );
  DFF_X1 \mem_reg[6][28]  ( .D(n522), .CK(clk), .Q(\mem[6][28] ) );
  DFF_X1 \mem_reg[6][27]  ( .D(n521), .CK(clk), .Q(\mem[6][27] ) );
  DFF_X1 \mem_reg[6][26]  ( .D(n520), .CK(clk), .Q(\mem[6][26] ) );
  DFF_X1 \mem_reg[6][25]  ( .D(n519), .CK(clk), .Q(\mem[6][25] ) );
  DFF_X1 \mem_reg[6][24]  ( .D(n518), .CK(clk), .Q(\mem[6][24] ) );
  DFF_X1 \mem_reg[6][23]  ( .D(n517), .CK(clk), .Q(\mem[6][23] ) );
  DFF_X1 \mem_reg[6][22]  ( .D(n516), .CK(clk), .Q(\mem[6][22] ) );
  DFF_X1 \mem_reg[6][21]  ( .D(n515), .CK(clk), .Q(\mem[6][21] ) );
  DFF_X1 \mem_reg[6][20]  ( .D(n514), .CK(clk), .Q(\mem[6][20] ) );
  DFF_X1 \mem_reg[6][19]  ( .D(n513), .CK(clk), .Q(\mem[6][19] ) );
  DFF_X1 \mem_reg[6][18]  ( .D(n512), .CK(clk), .Q(\mem[6][18] ) );
  DFF_X1 \mem_reg[6][17]  ( .D(n511), .CK(clk), .Q(\mem[6][17] ) );
  DFF_X1 \mem_reg[6][16]  ( .D(n510), .CK(clk), .Q(\mem[6][16] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n509), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n508), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n507), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n506), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n505), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n504), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n503), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n502), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n501), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n500), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n499), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n498), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n497), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n496), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n495), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n494), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][31]  ( .D(n493), .CK(clk), .Q(\mem[5][31] ) );
  DFF_X1 \mem_reg[5][30]  ( .D(n492), .CK(clk), .Q(\mem[5][30] ) );
  DFF_X1 \mem_reg[5][29]  ( .D(n491), .CK(clk), .Q(\mem[5][29] ) );
  DFF_X1 \mem_reg[5][28]  ( .D(n490), .CK(clk), .Q(\mem[5][28] ) );
  DFF_X1 \mem_reg[5][27]  ( .D(n489), .CK(clk), .Q(\mem[5][27] ) );
  DFF_X1 \mem_reg[5][26]  ( .D(n488), .CK(clk), .Q(\mem[5][26] ) );
  DFF_X1 \mem_reg[5][25]  ( .D(n487), .CK(clk), .Q(\mem[5][25] ) );
  DFF_X1 \mem_reg[5][24]  ( .D(n486), .CK(clk), .Q(\mem[5][24] ) );
  DFF_X1 \mem_reg[5][23]  ( .D(n485), .CK(clk), .Q(\mem[5][23] ) );
  DFF_X1 \mem_reg[5][22]  ( .D(n484), .CK(clk), .Q(\mem[5][22] ) );
  DFF_X1 \mem_reg[5][21]  ( .D(n483), .CK(clk), .Q(\mem[5][21] ) );
  DFF_X1 \mem_reg[5][20]  ( .D(n482), .CK(clk), .Q(\mem[5][20] ) );
  DFF_X1 \mem_reg[5][19]  ( .D(n481), .CK(clk), .Q(\mem[5][19] ) );
  DFF_X1 \mem_reg[5][18]  ( .D(n480), .CK(clk), .Q(\mem[5][18] ) );
  DFF_X1 \mem_reg[5][17]  ( .D(n479), .CK(clk), .Q(\mem[5][17] ) );
  DFF_X1 \mem_reg[5][16]  ( .D(n478), .CK(clk), .Q(\mem[5][16] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n477), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n476), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n475), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n474), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n473), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n472), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n471), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n470), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n469), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n468), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n467), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n466), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n465), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n464), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n463), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n462), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][31]  ( .D(n461), .CK(clk), .Q(\mem[4][31] ) );
  DFF_X1 \mem_reg[4][30]  ( .D(n460), .CK(clk), .Q(\mem[4][30] ) );
  DFF_X1 \mem_reg[4][29]  ( .D(n459), .CK(clk), .Q(\mem[4][29] ) );
  DFF_X1 \mem_reg[4][28]  ( .D(n458), .CK(clk), .Q(\mem[4][28] ) );
  DFF_X1 \mem_reg[4][27]  ( .D(n457), .CK(clk), .Q(\mem[4][27] ) );
  DFF_X1 \mem_reg[4][26]  ( .D(n456), .CK(clk), .Q(\mem[4][26] ) );
  DFF_X1 \mem_reg[4][25]  ( .D(n455), .CK(clk), .Q(\mem[4][25] ) );
  DFF_X1 \mem_reg[4][24]  ( .D(n454), .CK(clk), .Q(\mem[4][24] ) );
  DFF_X1 \mem_reg[4][23]  ( .D(n453), .CK(clk), .Q(\mem[4][23] ) );
  DFF_X1 \mem_reg[4][22]  ( .D(n452), .CK(clk), .Q(\mem[4][22] ) );
  DFF_X1 \mem_reg[4][21]  ( .D(n451), .CK(clk), .Q(\mem[4][21] ) );
  DFF_X1 \mem_reg[4][20]  ( .D(n450), .CK(clk), .Q(\mem[4][20] ) );
  DFF_X1 \mem_reg[4][19]  ( .D(n449), .CK(clk), .Q(\mem[4][19] ) );
  DFF_X1 \mem_reg[4][18]  ( .D(n448), .CK(clk), .Q(\mem[4][18] ) );
  DFF_X1 \mem_reg[4][17]  ( .D(n447), .CK(clk), .Q(\mem[4][17] ) );
  DFF_X1 \mem_reg[4][16]  ( .D(n446), .CK(clk), .Q(\mem[4][16] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n445), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n444), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n443), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n442), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n441), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n440), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n439), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n438), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n437), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n436), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n435), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n434), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n433), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n432), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n431), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n430), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][31]  ( .D(n429), .CK(clk), .Q(\mem[3][31] ) );
  DFF_X1 \mem_reg[3][30]  ( .D(n428), .CK(clk), .Q(\mem[3][30] ) );
  DFF_X1 \mem_reg[3][29]  ( .D(n427), .CK(clk), .Q(\mem[3][29] ) );
  DFF_X1 \mem_reg[3][28]  ( .D(n426), .CK(clk), .Q(\mem[3][28] ) );
  DFF_X1 \mem_reg[3][27]  ( .D(n425), .CK(clk), .Q(\mem[3][27] ) );
  DFF_X1 \mem_reg[3][26]  ( .D(n424), .CK(clk), .Q(\mem[3][26] ) );
  DFF_X1 \mem_reg[3][25]  ( .D(n423), .CK(clk), .Q(\mem[3][25] ) );
  DFF_X1 \mem_reg[3][24]  ( .D(n422), .CK(clk), .Q(\mem[3][24] ) );
  DFF_X1 \mem_reg[3][23]  ( .D(n421), .CK(clk), .Q(\mem[3][23] ) );
  DFF_X1 \mem_reg[3][22]  ( .D(n420), .CK(clk), .Q(\mem[3][22] ) );
  DFF_X1 \mem_reg[3][21]  ( .D(n419), .CK(clk), .Q(\mem[3][21] ) );
  DFF_X1 \mem_reg[3][20]  ( .D(n418), .CK(clk), .Q(\mem[3][20] ) );
  DFF_X1 \mem_reg[3][19]  ( .D(n417), .CK(clk), .Q(\mem[3][19] ) );
  DFF_X1 \mem_reg[3][18]  ( .D(n416), .CK(clk), .Q(\mem[3][18] ) );
  DFF_X1 \mem_reg[3][17]  ( .D(n415), .CK(clk), .Q(\mem[3][17] ) );
  DFF_X1 \mem_reg[3][16]  ( .D(n414), .CK(clk), .Q(\mem[3][16] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n413), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n412), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n411), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n410), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n409), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n408), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n407), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n406), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n405), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n404), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n403), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n402), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n401), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n400), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n399), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n398), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][31]  ( .D(n397), .CK(clk), .Q(\mem[2][31] ) );
  DFF_X1 \mem_reg[2][30]  ( .D(n396), .CK(clk), .Q(\mem[2][30] ) );
  DFF_X1 \mem_reg[2][29]  ( .D(n395), .CK(clk), .Q(\mem[2][29] ) );
  DFF_X1 \mem_reg[2][28]  ( .D(n394), .CK(clk), .Q(\mem[2][28] ) );
  DFF_X1 \mem_reg[2][27]  ( .D(n393), .CK(clk), .Q(\mem[2][27] ) );
  DFF_X1 \mem_reg[2][26]  ( .D(n392), .CK(clk), .Q(\mem[2][26] ) );
  DFF_X1 \mem_reg[2][25]  ( .D(n391), .CK(clk), .Q(\mem[2][25] ) );
  DFF_X1 \mem_reg[2][24]  ( .D(n390), .CK(clk), .Q(\mem[2][24] ) );
  DFF_X1 \mem_reg[2][23]  ( .D(n389), .CK(clk), .Q(\mem[2][23] ) );
  DFF_X1 \mem_reg[2][22]  ( .D(n388), .CK(clk), .Q(\mem[2][22] ) );
  DFF_X1 \mem_reg[2][21]  ( .D(n387), .CK(clk), .Q(\mem[2][21] ) );
  DFF_X1 \mem_reg[2][20]  ( .D(n386), .CK(clk), .Q(\mem[2][20] ) );
  DFF_X1 \mem_reg[2][19]  ( .D(n385), .CK(clk), .Q(\mem[2][19] ) );
  DFF_X1 \mem_reg[2][18]  ( .D(n384), .CK(clk), .Q(\mem[2][18] ) );
  DFF_X1 \mem_reg[2][17]  ( .D(n383), .CK(clk), .Q(\mem[2][17] ) );
  DFF_X1 \mem_reg[2][16]  ( .D(n382), .CK(clk), .Q(\mem[2][16] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n381), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n380), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n379), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n378), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n377), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n376), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n375), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n374), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n373), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n372), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n371), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n370), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n369), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n368), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n367), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n366), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][31]  ( .D(n365), .CK(clk), .Q(\mem[1][31] ) );
  DFF_X1 \mem_reg[1][30]  ( .D(n364), .CK(clk), .Q(\mem[1][30] ) );
  DFF_X1 \mem_reg[1][29]  ( .D(n363), .CK(clk), .Q(\mem[1][29] ) );
  DFF_X1 \mem_reg[1][28]  ( .D(n362), .CK(clk), .Q(\mem[1][28] ) );
  DFF_X1 \mem_reg[1][27]  ( .D(n361), .CK(clk), .Q(\mem[1][27] ) );
  DFF_X1 \mem_reg[1][26]  ( .D(n360), .CK(clk), .Q(\mem[1][26] ) );
  DFF_X1 \mem_reg[1][25]  ( .D(n359), .CK(clk), .Q(\mem[1][25] ) );
  DFF_X1 \mem_reg[1][24]  ( .D(n358), .CK(clk), .Q(\mem[1][24] ) );
  DFF_X1 \mem_reg[1][23]  ( .D(n357), .CK(clk), .Q(\mem[1][23] ) );
  DFF_X1 \mem_reg[1][22]  ( .D(n356), .CK(clk), .Q(\mem[1][22] ) );
  DFF_X1 \mem_reg[1][21]  ( .D(n355), .CK(clk), .Q(\mem[1][21] ) );
  DFF_X1 \mem_reg[1][20]  ( .D(n354), .CK(clk), .Q(\mem[1][20] ) );
  DFF_X1 \mem_reg[1][19]  ( .D(n353), .CK(clk), .Q(\mem[1][19] ) );
  DFF_X1 \mem_reg[1][18]  ( .D(n352), .CK(clk), .Q(\mem[1][18] ) );
  DFF_X1 \mem_reg[1][17]  ( .D(n351), .CK(clk), .Q(\mem[1][17] ) );
  DFF_X1 \mem_reg[1][16]  ( .D(n350), .CK(clk), .Q(\mem[1][16] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n349), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n348), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n347), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n346), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n345), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n344), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n343), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n342), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n341), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n340), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n339), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n338), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n337), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n336), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n335), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n334), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][31]  ( .D(n333), .CK(clk), .Q(\mem[0][31] ) );
  DFF_X1 \mem_reg[0][30]  ( .D(n332), .CK(clk), .Q(\mem[0][30] ) );
  DFF_X1 \mem_reg[0][29]  ( .D(n331), .CK(clk), .Q(\mem[0][29] ) );
  DFF_X1 \mem_reg[0][28]  ( .D(n330), .CK(clk), .Q(\mem[0][28] ) );
  DFF_X1 \mem_reg[0][27]  ( .D(n329), .CK(clk), .Q(\mem[0][27] ) );
  DFF_X1 \mem_reg[0][26]  ( .D(n328), .CK(clk), .Q(\mem[0][26] ) );
  DFF_X1 \mem_reg[0][25]  ( .D(n327), .CK(clk), .Q(\mem[0][25] ) );
  DFF_X1 \mem_reg[0][24]  ( .D(n326), .CK(clk), .Q(\mem[0][24] ) );
  DFF_X1 \mem_reg[0][23]  ( .D(n325), .CK(clk), .Q(\mem[0][23] ) );
  DFF_X1 \mem_reg[0][22]  ( .D(n324), .CK(clk), .Q(\mem[0][22] ) );
  DFF_X1 \mem_reg[0][21]  ( .D(n323), .CK(clk), .Q(\mem[0][21] ) );
  DFF_X1 \mem_reg[0][20]  ( .D(n322), .CK(clk), .Q(\mem[0][20] ) );
  DFF_X1 \mem_reg[0][19]  ( .D(n321), .CK(clk), .Q(\mem[0][19] ) );
  DFF_X1 \mem_reg[0][18]  ( .D(n320), .CK(clk), .Q(\mem[0][18] ) );
  DFF_X1 \mem_reg[0][17]  ( .D(n319), .CK(clk), .Q(\mem[0][17] ) );
  DFF_X1 \mem_reg[0][16]  ( .D(n318), .CK(clk), .Q(\mem[0][16] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n317), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n316), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n315), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n314), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n313), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n312), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n311), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n310), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n309), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n308), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n307), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n306), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n305), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n304), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n303), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n302), .CK(clk), .Q(\mem[0][0] ) );
  NAND3_X1 U552 ( .A1(n741), .A2(n742), .A3(n69), .ZN(n36) );
  NAND3_X1 U553 ( .A1(n69), .A2(n742), .A3(N10), .ZN(n70) );
  NAND3_X1 U554 ( .A1(n69), .A2(n741), .A3(N11), .ZN(n103) );
  NAND3_X1 U555 ( .A1(N10), .A2(n69), .A3(N11), .ZN(n136) );
  NAND3_X1 U556 ( .A1(n741), .A2(n742), .A3(n202), .ZN(n169) );
  NAND3_X1 U557 ( .A1(N10), .A2(n742), .A3(n202), .ZN(n203) );
  NAND3_X1 U558 ( .A1(N11), .A2(n741), .A3(n202), .ZN(n236) );
  NAND3_X1 U559 ( .A1(N11), .A2(N10), .A3(n202), .ZN(n269) );
  BUF_X1 U3 ( .A(n724), .Z(n720) );
  BUF_X1 U4 ( .A(n724), .Z(n721) );
  BUF_X1 U5 ( .A(n724), .Z(n722) );
  BUF_X1 U6 ( .A(n724), .Z(n723) );
  BUF_X1 U7 ( .A(N11), .Z(n716) );
  BUF_X1 U8 ( .A(N11), .Z(n717) );
  BUF_X1 U9 ( .A(N11), .Z(n718) );
  BUF_X1 U10 ( .A(N10), .Z(n724) );
  BUF_X1 U11 ( .A(n103), .Z(n736) );
  BUF_X1 U12 ( .A(n103), .Z(n735) );
  BUF_X1 U13 ( .A(n169), .Z(n732) );
  BUF_X1 U14 ( .A(n169), .Z(n731) );
  BUF_X1 U15 ( .A(n203), .Z(n730) );
  BUF_X1 U16 ( .A(n203), .Z(n729) );
  BUF_X1 U17 ( .A(n236), .Z(n728) );
  BUF_X1 U18 ( .A(n236), .Z(n727) );
  BUF_X1 U19 ( .A(n269), .Z(n726) );
  BUF_X1 U20 ( .A(n269), .Z(n725) );
  BUF_X1 U21 ( .A(n70), .Z(n737) );
  BUF_X1 U22 ( .A(n36), .Z(n739) );
  BUF_X1 U23 ( .A(n70), .Z(n738) );
  BUF_X1 U24 ( .A(n136), .Z(n733) );
  INV_X1 U25 ( .A(N10), .ZN(n741) );
  INV_X1 U26 ( .A(N11), .ZN(n742) );
  BUF_X1 U27 ( .A(N12), .Z(n715) );
  NOR2_X1 U28 ( .A1(n743), .A2(N12), .ZN(n69) );
  INV_X1 U29 ( .A(wr_en), .ZN(n743) );
  AND2_X1 U30 ( .A1(N12), .A2(wr_en), .ZN(n202) );
  OAI21_X1 U31 ( .B1(n748), .B2(n236), .A(n264), .ZN(n521) );
  NAND2_X1 U32 ( .A1(\mem[6][27] ), .A2(n727), .ZN(n264) );
  OAI21_X1 U33 ( .B1(n747), .B2(n236), .A(n265), .ZN(n522) );
  NAND2_X1 U34 ( .A1(\mem[6][28] ), .A2(n727), .ZN(n265) );
  OAI21_X1 U35 ( .B1(n746), .B2(n236), .A(n266), .ZN(n523) );
  NAND2_X1 U36 ( .A1(\mem[6][29] ), .A2(n727), .ZN(n266) );
  OAI21_X1 U37 ( .B1(n745), .B2(n236), .A(n267), .ZN(n524) );
  NAND2_X1 U38 ( .A1(\mem[6][30] ), .A2(n727), .ZN(n267) );
  OAI21_X1 U39 ( .B1(n748), .B2(n269), .A(n297), .ZN(n553) );
  NAND2_X1 U40 ( .A1(\mem[7][27] ), .A2(n725), .ZN(n297) );
  OAI21_X1 U41 ( .B1(n747), .B2(n269), .A(n298), .ZN(n554) );
  NAND2_X1 U42 ( .A1(\mem[7][28] ), .A2(n725), .ZN(n298) );
  OAI21_X1 U43 ( .B1(n746), .B2(n269), .A(n299), .ZN(n555) );
  NAND2_X1 U44 ( .A1(\mem[7][29] ), .A2(n725), .ZN(n299) );
  OAI21_X1 U45 ( .B1(n745), .B2(n269), .A(n300), .ZN(n556) );
  NAND2_X1 U46 ( .A1(\mem[7][30] ), .A2(n725), .ZN(n300) );
  OAI21_X1 U47 ( .B1(n748), .B2(n70), .A(n98), .ZN(n361) );
  NAND2_X1 U48 ( .A1(\mem[1][27] ), .A2(n70), .ZN(n98) );
  OAI21_X1 U49 ( .B1(n747), .B2(n737), .A(n99), .ZN(n362) );
  NAND2_X1 U50 ( .A1(\mem[1][28] ), .A2(n70), .ZN(n99) );
  OAI21_X1 U51 ( .B1(n746), .B2(n738), .A(n100), .ZN(n363) );
  NAND2_X1 U52 ( .A1(\mem[1][29] ), .A2(n70), .ZN(n100) );
  OAI21_X1 U53 ( .B1(n745), .B2(n737), .A(n101), .ZN(n364) );
  NAND2_X1 U54 ( .A1(\mem[1][30] ), .A2(n70), .ZN(n101) );
  OAI21_X1 U55 ( .B1(n748), .B2(n735), .A(n131), .ZN(n393) );
  NAND2_X1 U56 ( .A1(\mem[2][27] ), .A2(n735), .ZN(n131) );
  OAI21_X1 U57 ( .B1(n747), .B2(n735), .A(n132), .ZN(n394) );
  NAND2_X1 U58 ( .A1(\mem[2][28] ), .A2(n735), .ZN(n132) );
  OAI21_X1 U59 ( .B1(n746), .B2(n736), .A(n133), .ZN(n395) );
  NAND2_X1 U60 ( .A1(\mem[2][29] ), .A2(n735), .ZN(n133) );
  OAI21_X1 U61 ( .B1(n745), .B2(n103), .A(n134), .ZN(n396) );
  NAND2_X1 U62 ( .A1(\mem[2][30] ), .A2(n735), .ZN(n134) );
  OAI21_X1 U63 ( .B1(n748), .B2(n734), .A(n164), .ZN(n425) );
  NAND2_X1 U64 ( .A1(\mem[3][27] ), .A2(n136), .ZN(n164) );
  OAI21_X1 U65 ( .B1(n747), .B2(n734), .A(n165), .ZN(n426) );
  NAND2_X1 U66 ( .A1(\mem[3][28] ), .A2(n136), .ZN(n165) );
  OAI21_X1 U67 ( .B1(n746), .B2(n734), .A(n166), .ZN(n427) );
  NAND2_X1 U68 ( .A1(\mem[3][29] ), .A2(n136), .ZN(n166) );
  OAI21_X1 U69 ( .B1(n745), .B2(n734), .A(n167), .ZN(n428) );
  NAND2_X1 U70 ( .A1(\mem[3][30] ), .A2(n136), .ZN(n167) );
  OAI21_X1 U71 ( .B1(n748), .B2(n731), .A(n197), .ZN(n457) );
  NAND2_X1 U72 ( .A1(\mem[4][27] ), .A2(n731), .ZN(n197) );
  OAI21_X1 U73 ( .B1(n747), .B2(n731), .A(n198), .ZN(n458) );
  NAND2_X1 U74 ( .A1(\mem[4][28] ), .A2(n731), .ZN(n198) );
  OAI21_X1 U75 ( .B1(n746), .B2(n732), .A(n199), .ZN(n459) );
  NAND2_X1 U76 ( .A1(\mem[4][29] ), .A2(n731), .ZN(n199) );
  OAI21_X1 U77 ( .B1(n745), .B2(n169), .A(n200), .ZN(n460) );
  NAND2_X1 U78 ( .A1(\mem[4][30] ), .A2(n731), .ZN(n200) );
  OAI21_X1 U79 ( .B1(n748), .B2(n203), .A(n231), .ZN(n489) );
  NAND2_X1 U80 ( .A1(\mem[5][27] ), .A2(n729), .ZN(n231) );
  OAI21_X1 U81 ( .B1(n747), .B2(n203), .A(n232), .ZN(n490) );
  NAND2_X1 U82 ( .A1(\mem[5][28] ), .A2(n729), .ZN(n232) );
  OAI21_X1 U83 ( .B1(n746), .B2(n203), .A(n233), .ZN(n491) );
  NAND2_X1 U84 ( .A1(\mem[5][29] ), .A2(n729), .ZN(n233) );
  OAI21_X1 U85 ( .B1(n745), .B2(n203), .A(n234), .ZN(n492) );
  NAND2_X1 U86 ( .A1(\mem[5][30] ), .A2(n729), .ZN(n234) );
  OAI21_X1 U87 ( .B1(n774), .B2(n738), .A(n72), .ZN(n335) );
  NAND2_X1 U88 ( .A1(\mem[1][1] ), .A2(n738), .ZN(n72) );
  OAI21_X1 U89 ( .B1(n772), .B2(n70), .A(n74), .ZN(n337) );
  NAND2_X1 U90 ( .A1(\mem[1][3] ), .A2(n70), .ZN(n74) );
  OAI21_X1 U91 ( .B1(n771), .B2(n70), .A(n75), .ZN(n338) );
  NAND2_X1 U92 ( .A1(\mem[1][4] ), .A2(n738), .ZN(n75) );
  OAI21_X1 U93 ( .B1(n744), .B2(n70), .A(n102), .ZN(n365) );
  NAND2_X1 U94 ( .A1(\mem[1][31] ), .A2(n70), .ZN(n102) );
  OAI21_X1 U95 ( .B1(n774), .B2(n735), .A(n105), .ZN(n367) );
  NAND2_X1 U96 ( .A1(\mem[2][1] ), .A2(n735), .ZN(n105) );
  OAI21_X1 U97 ( .B1(n772), .B2(n736), .A(n107), .ZN(n369) );
  NAND2_X1 U98 ( .A1(\mem[2][3] ), .A2(n735), .ZN(n107) );
  OAI21_X1 U99 ( .B1(n771), .B2(n735), .A(n108), .ZN(n370) );
  NAND2_X1 U100 ( .A1(\mem[2][4] ), .A2(n736), .ZN(n108) );
  OAI21_X1 U101 ( .B1(n744), .B2(n736), .A(n135), .ZN(n397) );
  NAND2_X1 U102 ( .A1(\mem[2][31] ), .A2(n735), .ZN(n135) );
  OAI21_X1 U103 ( .B1(n774), .B2(n136), .A(n138), .ZN(n399) );
  NAND2_X1 U104 ( .A1(\mem[3][1] ), .A2(n136), .ZN(n138) );
  OAI21_X1 U105 ( .B1(n772), .B2(n733), .A(n140), .ZN(n401) );
  NAND2_X1 U106 ( .A1(\mem[3][3] ), .A2(n136), .ZN(n140) );
  OAI21_X1 U107 ( .B1(n771), .B2(n136), .A(n141), .ZN(n402) );
  NAND2_X1 U108 ( .A1(\mem[3][4] ), .A2(n136), .ZN(n141) );
  OAI21_X1 U109 ( .B1(n744), .B2(n136), .A(n168), .ZN(n429) );
  NAND2_X1 U110 ( .A1(\mem[3][31] ), .A2(n136), .ZN(n168) );
  OAI21_X1 U111 ( .B1(n774), .B2(n731), .A(n171), .ZN(n431) );
  NAND2_X1 U112 ( .A1(\mem[4][1] ), .A2(n731), .ZN(n171) );
  OAI21_X1 U113 ( .B1(n772), .B2(n732), .A(n173), .ZN(n433) );
  NAND2_X1 U114 ( .A1(\mem[4][3] ), .A2(n731), .ZN(n173) );
  OAI21_X1 U115 ( .B1(n771), .B2(n731), .A(n174), .ZN(n434) );
  NAND2_X1 U116 ( .A1(\mem[4][4] ), .A2(n732), .ZN(n174) );
  OAI21_X1 U117 ( .B1(n744), .B2(n732), .A(n201), .ZN(n461) );
  NAND2_X1 U118 ( .A1(\mem[4][31] ), .A2(n731), .ZN(n201) );
  OAI21_X1 U119 ( .B1(n774), .B2(n730), .A(n205), .ZN(n463) );
  NAND2_X1 U120 ( .A1(\mem[5][1] ), .A2(n729), .ZN(n205) );
  OAI21_X1 U121 ( .B1(n772), .B2(n729), .A(n207), .ZN(n465) );
  NAND2_X1 U122 ( .A1(\mem[5][3] ), .A2(n729), .ZN(n207) );
  OAI21_X1 U123 ( .B1(n771), .B2(n730), .A(n208), .ZN(n466) );
  NAND2_X1 U124 ( .A1(\mem[5][4] ), .A2(n730), .ZN(n208) );
  OAI21_X1 U125 ( .B1(n744), .B2(n729), .A(n235), .ZN(n493) );
  NAND2_X1 U126 ( .A1(\mem[5][31] ), .A2(n729), .ZN(n235) );
  OAI21_X1 U127 ( .B1(n774), .B2(n728), .A(n238), .ZN(n495) );
  NAND2_X1 U128 ( .A1(\mem[6][1] ), .A2(n727), .ZN(n238) );
  OAI21_X1 U129 ( .B1(n772), .B2(n727), .A(n240), .ZN(n497) );
  NAND2_X1 U130 ( .A1(\mem[6][3] ), .A2(n727), .ZN(n240) );
  OAI21_X1 U131 ( .B1(n771), .B2(n728), .A(n241), .ZN(n498) );
  NAND2_X1 U132 ( .A1(\mem[6][4] ), .A2(n728), .ZN(n241) );
  OAI21_X1 U133 ( .B1(n744), .B2(n727), .A(n268), .ZN(n525) );
  NAND2_X1 U134 ( .A1(\mem[6][31] ), .A2(n727), .ZN(n268) );
  OAI21_X1 U135 ( .B1(n774), .B2(n726), .A(n271), .ZN(n527) );
  NAND2_X1 U136 ( .A1(\mem[7][1] ), .A2(n725), .ZN(n271) );
  OAI21_X1 U137 ( .B1(n772), .B2(n725), .A(n273), .ZN(n529) );
  NAND2_X1 U138 ( .A1(\mem[7][3] ), .A2(n725), .ZN(n273) );
  OAI21_X1 U139 ( .B1(n771), .B2(n726), .A(n274), .ZN(n530) );
  NAND2_X1 U140 ( .A1(\mem[7][4] ), .A2(n726), .ZN(n274) );
  OAI21_X1 U141 ( .B1(n744), .B2(n725), .A(n301), .ZN(n557) );
  NAND2_X1 U142 ( .A1(\mem[7][31] ), .A2(n725), .ZN(n301) );
  OAI21_X1 U143 ( .B1(n775), .B2(n737), .A(n71), .ZN(n334) );
  NAND2_X1 U144 ( .A1(\mem[1][0] ), .A2(n738), .ZN(n71) );
  OAI21_X1 U145 ( .B1(n773), .B2(n737), .A(n73), .ZN(n336) );
  NAND2_X1 U146 ( .A1(\mem[1][2] ), .A2(n737), .ZN(n73) );
  OAI21_X1 U147 ( .B1(n770), .B2(n737), .A(n76), .ZN(n339) );
  NAND2_X1 U148 ( .A1(\mem[1][5] ), .A2(n737), .ZN(n76) );
  OAI21_X1 U149 ( .B1(n769), .B2(n737), .A(n77), .ZN(n340) );
  NAND2_X1 U150 ( .A1(\mem[1][6] ), .A2(n738), .ZN(n77) );
  OAI21_X1 U151 ( .B1(n768), .B2(n737), .A(n78), .ZN(n341) );
  NAND2_X1 U152 ( .A1(\mem[1][7] ), .A2(n70), .ZN(n78) );
  OAI21_X1 U153 ( .B1(n767), .B2(n737), .A(n79), .ZN(n342) );
  NAND2_X1 U154 ( .A1(\mem[1][8] ), .A2(n70), .ZN(n79) );
  OAI21_X1 U155 ( .B1(n766), .B2(n737), .A(n80), .ZN(n343) );
  NAND2_X1 U156 ( .A1(\mem[1][9] ), .A2(n70), .ZN(n80) );
  OAI21_X1 U157 ( .B1(n765), .B2(n737), .A(n81), .ZN(n344) );
  NAND2_X1 U158 ( .A1(\mem[1][10] ), .A2(n737), .ZN(n81) );
  OAI21_X1 U159 ( .B1(n764), .B2(n737), .A(n82), .ZN(n345) );
  NAND2_X1 U160 ( .A1(\mem[1][11] ), .A2(n738), .ZN(n82) );
  OAI21_X1 U161 ( .B1(n763), .B2(n737), .A(n83), .ZN(n346) );
  NAND2_X1 U162 ( .A1(\mem[1][12] ), .A2(n737), .ZN(n83) );
  OAI21_X1 U163 ( .B1(n762), .B2(n737), .A(n84), .ZN(n347) );
  NAND2_X1 U164 ( .A1(\mem[1][13] ), .A2(n737), .ZN(n84) );
  OAI21_X1 U165 ( .B1(n761), .B2(n737), .A(n85), .ZN(n348) );
  NAND2_X1 U166 ( .A1(\mem[1][14] ), .A2(n70), .ZN(n85) );
  OAI21_X1 U167 ( .B1(n775), .B2(n103), .A(n104), .ZN(n366) );
  NAND2_X1 U168 ( .A1(\mem[2][0] ), .A2(n735), .ZN(n104) );
  OAI21_X1 U169 ( .B1(n773), .B2(n103), .A(n106), .ZN(n368) );
  NAND2_X1 U170 ( .A1(\mem[2][2] ), .A2(n735), .ZN(n106) );
  OAI21_X1 U171 ( .B1(n770), .B2(n103), .A(n109), .ZN(n371) );
  NAND2_X1 U172 ( .A1(\mem[2][5] ), .A2(n736), .ZN(n109) );
  OAI21_X1 U173 ( .B1(n769), .B2(n103), .A(n110), .ZN(n372) );
  NAND2_X1 U174 ( .A1(\mem[2][6] ), .A2(n736), .ZN(n110) );
  OAI21_X1 U175 ( .B1(n768), .B2(n103), .A(n111), .ZN(n373) );
  NAND2_X1 U176 ( .A1(\mem[2][7] ), .A2(n735), .ZN(n111) );
  OAI21_X1 U177 ( .B1(n767), .B2(n103), .A(n112), .ZN(n374) );
  NAND2_X1 U178 ( .A1(\mem[2][8] ), .A2(n736), .ZN(n112) );
  OAI21_X1 U179 ( .B1(n766), .B2(n103), .A(n113), .ZN(n375) );
  NAND2_X1 U180 ( .A1(\mem[2][9] ), .A2(n103), .ZN(n113) );
  OAI21_X1 U181 ( .B1(n765), .B2(n103), .A(n114), .ZN(n376) );
  NAND2_X1 U182 ( .A1(\mem[2][10] ), .A2(n103), .ZN(n114) );
  OAI21_X1 U183 ( .B1(n764), .B2(n103), .A(n115), .ZN(n377) );
  NAND2_X1 U184 ( .A1(\mem[2][11] ), .A2(n735), .ZN(n115) );
  OAI21_X1 U185 ( .B1(n763), .B2(n103), .A(n116), .ZN(n378) );
  NAND2_X1 U186 ( .A1(\mem[2][12] ), .A2(n736), .ZN(n116) );
  OAI21_X1 U187 ( .B1(n762), .B2(n103), .A(n117), .ZN(n379) );
  NAND2_X1 U188 ( .A1(\mem[2][13] ), .A2(n736), .ZN(n117) );
  OAI21_X1 U189 ( .B1(n761), .B2(n103), .A(n118), .ZN(n380) );
  NAND2_X1 U190 ( .A1(\mem[2][14] ), .A2(n735), .ZN(n118) );
  OAI21_X1 U191 ( .B1(n775), .B2(n734), .A(n137), .ZN(n398) );
  NAND2_X1 U192 ( .A1(\mem[3][0] ), .A2(n136), .ZN(n137) );
  OAI21_X1 U193 ( .B1(n773), .B2(n734), .A(n139), .ZN(n400) );
  NAND2_X1 U194 ( .A1(\mem[3][2] ), .A2(n136), .ZN(n139) );
  OAI21_X1 U195 ( .B1(n770), .B2(n734), .A(n142), .ZN(n403) );
  NAND2_X1 U196 ( .A1(\mem[3][5] ), .A2(n733), .ZN(n142) );
  OAI21_X1 U197 ( .B1(n769), .B2(n733), .A(n143), .ZN(n404) );
  NAND2_X1 U198 ( .A1(\mem[3][6] ), .A2(n136), .ZN(n143) );
  OAI21_X1 U199 ( .B1(n768), .B2(n733), .A(n144), .ZN(n405) );
  NAND2_X1 U200 ( .A1(\mem[3][7] ), .A2(n734), .ZN(n144) );
  OAI21_X1 U201 ( .B1(n767), .B2(n734), .A(n145), .ZN(n406) );
  NAND2_X1 U202 ( .A1(\mem[3][8] ), .A2(n136), .ZN(n145) );
  OAI21_X1 U203 ( .B1(n766), .B2(n733), .A(n146), .ZN(n407) );
  NAND2_X1 U204 ( .A1(\mem[3][9] ), .A2(n733), .ZN(n146) );
  OAI21_X1 U205 ( .B1(n765), .B2(n734), .A(n147), .ZN(n408) );
  NAND2_X1 U206 ( .A1(\mem[3][10] ), .A2(n136), .ZN(n147) );
  OAI21_X1 U207 ( .B1(n764), .B2(n733), .A(n148), .ZN(n409) );
  NAND2_X1 U208 ( .A1(\mem[3][11] ), .A2(n136), .ZN(n148) );
  OAI21_X1 U209 ( .B1(n763), .B2(n734), .A(n149), .ZN(n410) );
  NAND2_X1 U210 ( .A1(\mem[3][12] ), .A2(n136), .ZN(n149) );
  OAI21_X1 U211 ( .B1(n762), .B2(n733), .A(n150), .ZN(n411) );
  NAND2_X1 U212 ( .A1(\mem[3][13] ), .A2(n734), .ZN(n150) );
  OAI21_X1 U213 ( .B1(n761), .B2(n734), .A(n151), .ZN(n412) );
  NAND2_X1 U214 ( .A1(\mem[3][14] ), .A2(n136), .ZN(n151) );
  OAI21_X1 U215 ( .B1(n775), .B2(n169), .A(n170), .ZN(n430) );
  NAND2_X1 U216 ( .A1(\mem[4][0] ), .A2(n731), .ZN(n170) );
  OAI21_X1 U217 ( .B1(n773), .B2(n169), .A(n172), .ZN(n432) );
  NAND2_X1 U218 ( .A1(\mem[4][2] ), .A2(n731), .ZN(n172) );
  OAI21_X1 U219 ( .B1(n770), .B2(n169), .A(n175), .ZN(n435) );
  NAND2_X1 U220 ( .A1(\mem[4][5] ), .A2(n732), .ZN(n175) );
  OAI21_X1 U221 ( .B1(n769), .B2(n169), .A(n176), .ZN(n436) );
  NAND2_X1 U222 ( .A1(\mem[4][6] ), .A2(n732), .ZN(n176) );
  OAI21_X1 U223 ( .B1(n768), .B2(n169), .A(n177), .ZN(n437) );
  NAND2_X1 U224 ( .A1(\mem[4][7] ), .A2(n731), .ZN(n177) );
  OAI21_X1 U225 ( .B1(n767), .B2(n169), .A(n178), .ZN(n438) );
  NAND2_X1 U226 ( .A1(\mem[4][8] ), .A2(n732), .ZN(n178) );
  OAI21_X1 U227 ( .B1(n766), .B2(n169), .A(n179), .ZN(n439) );
  NAND2_X1 U228 ( .A1(\mem[4][9] ), .A2(n169), .ZN(n179) );
  OAI21_X1 U229 ( .B1(n765), .B2(n169), .A(n180), .ZN(n440) );
  NAND2_X1 U230 ( .A1(\mem[4][10] ), .A2(n169), .ZN(n180) );
  OAI21_X1 U231 ( .B1(n764), .B2(n169), .A(n181), .ZN(n441) );
  NAND2_X1 U232 ( .A1(\mem[4][11] ), .A2(n731), .ZN(n181) );
  OAI21_X1 U233 ( .B1(n763), .B2(n169), .A(n182), .ZN(n442) );
  NAND2_X1 U234 ( .A1(\mem[4][12] ), .A2(n732), .ZN(n182) );
  OAI21_X1 U235 ( .B1(n762), .B2(n169), .A(n183), .ZN(n443) );
  NAND2_X1 U236 ( .A1(\mem[4][13] ), .A2(n732), .ZN(n183) );
  OAI21_X1 U237 ( .B1(n761), .B2(n169), .A(n184), .ZN(n444) );
  NAND2_X1 U238 ( .A1(\mem[4][14] ), .A2(n731), .ZN(n184) );
  OAI21_X1 U239 ( .B1(n775), .B2(n730), .A(n204), .ZN(n462) );
  NAND2_X1 U240 ( .A1(\mem[5][0] ), .A2(n729), .ZN(n204) );
  OAI21_X1 U241 ( .B1(n773), .B2(n729), .A(n206), .ZN(n464) );
  NAND2_X1 U242 ( .A1(\mem[5][2] ), .A2(n729), .ZN(n206) );
  OAI21_X1 U243 ( .B1(n770), .B2(n730), .A(n209), .ZN(n467) );
  NAND2_X1 U244 ( .A1(\mem[5][5] ), .A2(n730), .ZN(n209) );
  OAI21_X1 U245 ( .B1(n769), .B2(n203), .A(n210), .ZN(n468) );
  NAND2_X1 U246 ( .A1(\mem[5][6] ), .A2(n730), .ZN(n210) );
  OAI21_X1 U247 ( .B1(n768), .B2(n203), .A(n211), .ZN(n469) );
  NAND2_X1 U248 ( .A1(\mem[5][7] ), .A2(n730), .ZN(n211) );
  OAI21_X1 U249 ( .B1(n767), .B2(n203), .A(n212), .ZN(n470) );
  NAND2_X1 U250 ( .A1(\mem[5][8] ), .A2(n729), .ZN(n212) );
  OAI21_X1 U251 ( .B1(n766), .B2(n203), .A(n213), .ZN(n471) );
  NAND2_X1 U252 ( .A1(\mem[5][9] ), .A2(n203), .ZN(n213) );
  OAI21_X1 U253 ( .B1(n765), .B2(n203), .A(n214), .ZN(n472) );
  NAND2_X1 U254 ( .A1(\mem[5][10] ), .A2(n203), .ZN(n214) );
  OAI21_X1 U255 ( .B1(n764), .B2(n203), .A(n215), .ZN(n473) );
  NAND2_X1 U256 ( .A1(\mem[5][11] ), .A2(n730), .ZN(n215) );
  OAI21_X1 U257 ( .B1(n763), .B2(n203), .A(n216), .ZN(n474) );
  NAND2_X1 U258 ( .A1(\mem[5][12] ), .A2(n729), .ZN(n216) );
  OAI21_X1 U259 ( .B1(n762), .B2(n203), .A(n217), .ZN(n475) );
  NAND2_X1 U260 ( .A1(\mem[5][13] ), .A2(n730), .ZN(n217) );
  OAI21_X1 U261 ( .B1(n761), .B2(n203), .A(n218), .ZN(n476) );
  NAND2_X1 U262 ( .A1(\mem[5][14] ), .A2(n730), .ZN(n218) );
  OAI21_X1 U263 ( .B1(n775), .B2(n728), .A(n237), .ZN(n494) );
  NAND2_X1 U264 ( .A1(\mem[6][0] ), .A2(n727), .ZN(n237) );
  OAI21_X1 U265 ( .B1(n773), .B2(n727), .A(n239), .ZN(n496) );
  NAND2_X1 U266 ( .A1(\mem[6][2] ), .A2(n727), .ZN(n239) );
  OAI21_X1 U267 ( .B1(n770), .B2(n728), .A(n242), .ZN(n499) );
  NAND2_X1 U268 ( .A1(\mem[6][5] ), .A2(n728), .ZN(n242) );
  OAI21_X1 U269 ( .B1(n769), .B2(n236), .A(n243), .ZN(n500) );
  NAND2_X1 U270 ( .A1(\mem[6][6] ), .A2(n728), .ZN(n243) );
  OAI21_X1 U271 ( .B1(n768), .B2(n236), .A(n244), .ZN(n501) );
  NAND2_X1 U272 ( .A1(\mem[6][7] ), .A2(n728), .ZN(n244) );
  OAI21_X1 U273 ( .B1(n767), .B2(n236), .A(n245), .ZN(n502) );
  NAND2_X1 U274 ( .A1(\mem[6][8] ), .A2(n727), .ZN(n245) );
  OAI21_X1 U275 ( .B1(n766), .B2(n236), .A(n246), .ZN(n503) );
  NAND2_X1 U276 ( .A1(\mem[6][9] ), .A2(n236), .ZN(n246) );
  OAI21_X1 U277 ( .B1(n765), .B2(n236), .A(n247), .ZN(n504) );
  NAND2_X1 U278 ( .A1(\mem[6][10] ), .A2(n236), .ZN(n247) );
  OAI21_X1 U279 ( .B1(n764), .B2(n236), .A(n248), .ZN(n505) );
  NAND2_X1 U280 ( .A1(\mem[6][11] ), .A2(n728), .ZN(n248) );
  OAI21_X1 U281 ( .B1(n763), .B2(n236), .A(n249), .ZN(n506) );
  NAND2_X1 U282 ( .A1(\mem[6][12] ), .A2(n727), .ZN(n249) );
  OAI21_X1 U283 ( .B1(n762), .B2(n236), .A(n250), .ZN(n507) );
  NAND2_X1 U284 ( .A1(\mem[6][13] ), .A2(n728), .ZN(n250) );
  OAI21_X1 U285 ( .B1(n761), .B2(n236), .A(n251), .ZN(n508) );
  NAND2_X1 U286 ( .A1(\mem[6][14] ), .A2(n728), .ZN(n251) );
  OAI21_X1 U287 ( .B1(n775), .B2(n726), .A(n270), .ZN(n526) );
  NAND2_X1 U288 ( .A1(\mem[7][0] ), .A2(n725), .ZN(n270) );
  OAI21_X1 U289 ( .B1(n773), .B2(n725), .A(n272), .ZN(n528) );
  NAND2_X1 U290 ( .A1(\mem[7][2] ), .A2(n725), .ZN(n272) );
  OAI21_X1 U291 ( .B1(n770), .B2(n726), .A(n275), .ZN(n531) );
  NAND2_X1 U292 ( .A1(\mem[7][5] ), .A2(n726), .ZN(n275) );
  OAI21_X1 U293 ( .B1(n769), .B2(n269), .A(n276), .ZN(n532) );
  NAND2_X1 U294 ( .A1(\mem[7][6] ), .A2(n726), .ZN(n276) );
  OAI21_X1 U295 ( .B1(n768), .B2(n269), .A(n277), .ZN(n533) );
  NAND2_X1 U296 ( .A1(\mem[7][7] ), .A2(n726), .ZN(n277) );
  OAI21_X1 U297 ( .B1(n767), .B2(n269), .A(n278), .ZN(n534) );
  NAND2_X1 U298 ( .A1(\mem[7][8] ), .A2(n725), .ZN(n278) );
  OAI21_X1 U299 ( .B1(n766), .B2(n269), .A(n279), .ZN(n535) );
  NAND2_X1 U300 ( .A1(\mem[7][9] ), .A2(n269), .ZN(n279) );
  OAI21_X1 U301 ( .B1(n765), .B2(n269), .A(n280), .ZN(n536) );
  NAND2_X1 U302 ( .A1(\mem[7][10] ), .A2(n269), .ZN(n280) );
  OAI21_X1 U303 ( .B1(n764), .B2(n269), .A(n281), .ZN(n537) );
  NAND2_X1 U304 ( .A1(\mem[7][11] ), .A2(n726), .ZN(n281) );
  OAI21_X1 U305 ( .B1(n763), .B2(n269), .A(n282), .ZN(n538) );
  NAND2_X1 U306 ( .A1(\mem[7][12] ), .A2(n725), .ZN(n282) );
  OAI21_X1 U307 ( .B1(n762), .B2(n269), .A(n283), .ZN(n539) );
  NAND2_X1 U308 ( .A1(\mem[7][13] ), .A2(n726), .ZN(n283) );
  OAI21_X1 U309 ( .B1(n761), .B2(n269), .A(n284), .ZN(n540) );
  NAND2_X1 U310 ( .A1(\mem[7][14] ), .A2(n726), .ZN(n284) );
  OAI21_X1 U311 ( .B1(n36), .B2(n774), .A(n38), .ZN(n303) );
  NAND2_X1 U312 ( .A1(\mem[0][1] ), .A2(n36), .ZN(n38) );
  OAI21_X1 U313 ( .B1(n36), .B2(n772), .A(n40), .ZN(n305) );
  NAND2_X1 U314 ( .A1(\mem[0][3] ), .A2(n36), .ZN(n40) );
  OAI21_X1 U315 ( .B1(n36), .B2(n771), .A(n41), .ZN(n306) );
  NAND2_X1 U316 ( .A1(\mem[0][4] ), .A2(n36), .ZN(n41) );
  OAI21_X1 U317 ( .B1(n36), .B2(n744), .A(n68), .ZN(n333) );
  NAND2_X1 U318 ( .A1(\mem[0][31] ), .A2(n36), .ZN(n68) );
  OAI21_X1 U319 ( .B1(n740), .B2(n746), .A(n66), .ZN(n331) );
  NAND2_X1 U320 ( .A1(\mem[0][29] ), .A2(n36), .ZN(n66) );
  OAI21_X1 U321 ( .B1(n740), .B2(n745), .A(n67), .ZN(n332) );
  NAND2_X1 U322 ( .A1(\mem[0][30] ), .A2(n36), .ZN(n67) );
  OAI21_X1 U323 ( .B1(n760), .B2(n738), .A(n86), .ZN(n349) );
  NAND2_X1 U324 ( .A1(\mem[1][15] ), .A2(n737), .ZN(n86) );
  OAI21_X1 U325 ( .B1(n759), .B2(n738), .A(n87), .ZN(n350) );
  NAND2_X1 U326 ( .A1(\mem[1][16] ), .A2(n737), .ZN(n87) );
  OAI21_X1 U327 ( .B1(n758), .B2(n738), .A(n88), .ZN(n351) );
  NAND2_X1 U328 ( .A1(\mem[1][17] ), .A2(n70), .ZN(n88) );
  OAI21_X1 U329 ( .B1(n757), .B2(n738), .A(n89), .ZN(n352) );
  NAND2_X1 U330 ( .A1(\mem[1][18] ), .A2(n70), .ZN(n89) );
  OAI21_X1 U331 ( .B1(n756), .B2(n738), .A(n90), .ZN(n353) );
  NAND2_X1 U332 ( .A1(\mem[1][19] ), .A2(n70), .ZN(n90) );
  OAI21_X1 U333 ( .B1(n760), .B2(n103), .A(n119), .ZN(n381) );
  NAND2_X1 U334 ( .A1(\mem[2][15] ), .A2(n736), .ZN(n119) );
  OAI21_X1 U335 ( .B1(n759), .B2(n103), .A(n120), .ZN(n382) );
  NAND2_X1 U336 ( .A1(\mem[2][16] ), .A2(n736), .ZN(n120) );
  OAI21_X1 U337 ( .B1(n758), .B2(n103), .A(n121), .ZN(n383) );
  NAND2_X1 U338 ( .A1(\mem[2][17] ), .A2(n736), .ZN(n121) );
  OAI21_X1 U339 ( .B1(n757), .B2(n103), .A(n122), .ZN(n384) );
  NAND2_X1 U340 ( .A1(\mem[2][18] ), .A2(n736), .ZN(n122) );
  OAI21_X1 U341 ( .B1(n756), .B2(n736), .A(n123), .ZN(n385) );
  NAND2_X1 U342 ( .A1(\mem[2][19] ), .A2(n736), .ZN(n123) );
  OAI21_X1 U343 ( .B1(n760), .B2(n733), .A(n152), .ZN(n413) );
  NAND2_X1 U344 ( .A1(\mem[3][15] ), .A2(n136), .ZN(n152) );
  OAI21_X1 U345 ( .B1(n759), .B2(n733), .A(n153), .ZN(n414) );
  NAND2_X1 U346 ( .A1(\mem[3][16] ), .A2(n734), .ZN(n153) );
  OAI21_X1 U347 ( .B1(n758), .B2(n733), .A(n154), .ZN(n415) );
  NAND2_X1 U348 ( .A1(\mem[3][17] ), .A2(n733), .ZN(n154) );
  OAI21_X1 U349 ( .B1(n757), .B2(n733), .A(n155), .ZN(n416) );
  NAND2_X1 U350 ( .A1(\mem[3][18] ), .A2(n733), .ZN(n155) );
  OAI21_X1 U351 ( .B1(n756), .B2(n733), .A(n156), .ZN(n417) );
  NAND2_X1 U352 ( .A1(\mem[3][19] ), .A2(n734), .ZN(n156) );
  OAI21_X1 U353 ( .B1(n760), .B2(n169), .A(n185), .ZN(n445) );
  NAND2_X1 U354 ( .A1(\mem[4][15] ), .A2(n732), .ZN(n185) );
  OAI21_X1 U355 ( .B1(n759), .B2(n169), .A(n186), .ZN(n446) );
  NAND2_X1 U356 ( .A1(\mem[4][16] ), .A2(n732), .ZN(n186) );
  OAI21_X1 U357 ( .B1(n758), .B2(n169), .A(n187), .ZN(n447) );
  NAND2_X1 U358 ( .A1(\mem[4][17] ), .A2(n732), .ZN(n187) );
  OAI21_X1 U359 ( .B1(n757), .B2(n169), .A(n188), .ZN(n448) );
  NAND2_X1 U360 ( .A1(\mem[4][18] ), .A2(n732), .ZN(n188) );
  OAI21_X1 U361 ( .B1(n756), .B2(n732), .A(n189), .ZN(n449) );
  NAND2_X1 U362 ( .A1(\mem[4][19] ), .A2(n732), .ZN(n189) );
  OAI21_X1 U363 ( .B1(n760), .B2(n203), .A(n219), .ZN(n477) );
  NAND2_X1 U364 ( .A1(\mem[5][15] ), .A2(n729), .ZN(n219) );
  OAI21_X1 U365 ( .B1(n759), .B2(n203), .A(n220), .ZN(n478) );
  NAND2_X1 U366 ( .A1(\mem[5][16] ), .A2(n730), .ZN(n220) );
  OAI21_X1 U367 ( .B1(n758), .B2(n203), .A(n221), .ZN(n479) );
  NAND2_X1 U368 ( .A1(\mem[5][17] ), .A2(n730), .ZN(n221) );
  OAI21_X1 U369 ( .B1(n757), .B2(n203), .A(n222), .ZN(n480) );
  NAND2_X1 U370 ( .A1(\mem[5][18] ), .A2(n730), .ZN(n222) );
  OAI21_X1 U371 ( .B1(n756), .B2(n203), .A(n223), .ZN(n481) );
  NAND2_X1 U372 ( .A1(\mem[5][19] ), .A2(n730), .ZN(n223) );
  OAI21_X1 U373 ( .B1(n760), .B2(n236), .A(n252), .ZN(n509) );
  NAND2_X1 U374 ( .A1(\mem[6][15] ), .A2(n727), .ZN(n252) );
  OAI21_X1 U375 ( .B1(n759), .B2(n236), .A(n253), .ZN(n510) );
  NAND2_X1 U376 ( .A1(\mem[6][16] ), .A2(n728), .ZN(n253) );
  OAI21_X1 U377 ( .B1(n758), .B2(n236), .A(n254), .ZN(n511) );
  NAND2_X1 U378 ( .A1(\mem[6][17] ), .A2(n728), .ZN(n254) );
  OAI21_X1 U379 ( .B1(n757), .B2(n236), .A(n255), .ZN(n512) );
  NAND2_X1 U380 ( .A1(\mem[6][18] ), .A2(n728), .ZN(n255) );
  OAI21_X1 U381 ( .B1(n756), .B2(n236), .A(n256), .ZN(n513) );
  NAND2_X1 U382 ( .A1(\mem[6][19] ), .A2(n728), .ZN(n256) );
  OAI21_X1 U383 ( .B1(n760), .B2(n269), .A(n285), .ZN(n541) );
  NAND2_X1 U384 ( .A1(\mem[7][15] ), .A2(n725), .ZN(n285) );
  OAI21_X1 U385 ( .B1(n759), .B2(n269), .A(n286), .ZN(n542) );
  NAND2_X1 U386 ( .A1(\mem[7][16] ), .A2(n726), .ZN(n286) );
  OAI21_X1 U387 ( .B1(n758), .B2(n269), .A(n287), .ZN(n543) );
  NAND2_X1 U388 ( .A1(\mem[7][17] ), .A2(n726), .ZN(n287) );
  OAI21_X1 U389 ( .B1(n757), .B2(n269), .A(n288), .ZN(n544) );
  NAND2_X1 U390 ( .A1(\mem[7][18] ), .A2(n726), .ZN(n288) );
  OAI21_X1 U391 ( .B1(n756), .B2(n269), .A(n289), .ZN(n545) );
  NAND2_X1 U392 ( .A1(\mem[7][19] ), .A2(n726), .ZN(n289) );
  OAI21_X1 U393 ( .B1(n755), .B2(n738), .A(n91), .ZN(n354) );
  NAND2_X1 U394 ( .A1(\mem[1][20] ), .A2(n70), .ZN(n91) );
  OAI21_X1 U395 ( .B1(n754), .B2(n738), .A(n92), .ZN(n355) );
  NAND2_X1 U396 ( .A1(\mem[1][21] ), .A2(n70), .ZN(n92) );
  OAI21_X1 U397 ( .B1(n753), .B2(n738), .A(n93), .ZN(n356) );
  NAND2_X1 U398 ( .A1(\mem[1][22] ), .A2(n70), .ZN(n93) );
  OAI21_X1 U399 ( .B1(n752), .B2(n738), .A(n94), .ZN(n357) );
  NAND2_X1 U400 ( .A1(\mem[1][23] ), .A2(n70), .ZN(n94) );
  OAI21_X1 U401 ( .B1(n751), .B2(n738), .A(n95), .ZN(n358) );
  NAND2_X1 U402 ( .A1(\mem[1][24] ), .A2(n70), .ZN(n95) );
  OAI21_X1 U403 ( .B1(n750), .B2(n738), .A(n96), .ZN(n359) );
  NAND2_X1 U404 ( .A1(\mem[1][25] ), .A2(n738), .ZN(n96) );
  OAI21_X1 U405 ( .B1(n749), .B2(n738), .A(n97), .ZN(n360) );
  NAND2_X1 U406 ( .A1(\mem[1][26] ), .A2(n70), .ZN(n97) );
  OAI21_X1 U407 ( .B1(n755), .B2(n735), .A(n124), .ZN(n386) );
  NAND2_X1 U408 ( .A1(\mem[2][20] ), .A2(n736), .ZN(n124) );
  OAI21_X1 U409 ( .B1(n754), .B2(n736), .A(n125), .ZN(n387) );
  NAND2_X1 U410 ( .A1(\mem[2][21] ), .A2(n736), .ZN(n125) );
  OAI21_X1 U411 ( .B1(n753), .B2(n103), .A(n126), .ZN(n388) );
  NAND2_X1 U412 ( .A1(\mem[2][22] ), .A2(n736), .ZN(n126) );
  OAI21_X1 U413 ( .B1(n752), .B2(n103), .A(n127), .ZN(n389) );
  NAND2_X1 U414 ( .A1(\mem[2][23] ), .A2(n736), .ZN(n127) );
  OAI21_X1 U415 ( .B1(n751), .B2(n103), .A(n128), .ZN(n390) );
  NAND2_X1 U416 ( .A1(\mem[2][24] ), .A2(n735), .ZN(n128) );
  OAI21_X1 U417 ( .B1(n750), .B2(n103), .A(n129), .ZN(n391) );
  NAND2_X1 U418 ( .A1(\mem[2][25] ), .A2(n735), .ZN(n129) );
  OAI21_X1 U419 ( .B1(n749), .B2(n103), .A(n130), .ZN(n392) );
  NAND2_X1 U420 ( .A1(\mem[2][26] ), .A2(n735), .ZN(n130) );
  OAI21_X1 U421 ( .B1(n755), .B2(n733), .A(n157), .ZN(n418) );
  NAND2_X1 U422 ( .A1(\mem[3][20] ), .A2(n733), .ZN(n157) );
  OAI21_X1 U423 ( .B1(n754), .B2(n733), .A(n158), .ZN(n419) );
  NAND2_X1 U424 ( .A1(\mem[3][21] ), .A2(n733), .ZN(n158) );
  OAI21_X1 U425 ( .B1(n753), .B2(n733), .A(n159), .ZN(n420) );
  NAND2_X1 U426 ( .A1(\mem[3][22] ), .A2(n734), .ZN(n159) );
  OAI21_X1 U427 ( .B1(n752), .B2(n733), .A(n160), .ZN(n421) );
  NAND2_X1 U428 ( .A1(\mem[3][23] ), .A2(n733), .ZN(n160) );
  OAI21_X1 U429 ( .B1(n751), .B2(n733), .A(n161), .ZN(n422) );
  NAND2_X1 U430 ( .A1(\mem[3][24] ), .A2(n136), .ZN(n161) );
  OAI21_X1 U431 ( .B1(n750), .B2(n733), .A(n162), .ZN(n423) );
  NAND2_X1 U432 ( .A1(\mem[3][25] ), .A2(n136), .ZN(n162) );
  OAI21_X1 U433 ( .B1(n749), .B2(n733), .A(n163), .ZN(n424) );
  NAND2_X1 U434 ( .A1(\mem[3][26] ), .A2(n136), .ZN(n163) );
  OAI21_X1 U435 ( .B1(n755), .B2(n731), .A(n190), .ZN(n450) );
  NAND2_X1 U436 ( .A1(\mem[4][20] ), .A2(n732), .ZN(n190) );
  OAI21_X1 U437 ( .B1(n754), .B2(n732), .A(n191), .ZN(n451) );
  NAND2_X1 U438 ( .A1(\mem[4][21] ), .A2(n732), .ZN(n191) );
  OAI21_X1 U439 ( .B1(n753), .B2(n169), .A(n192), .ZN(n452) );
  NAND2_X1 U440 ( .A1(\mem[4][22] ), .A2(n732), .ZN(n192) );
  OAI21_X1 U441 ( .B1(n752), .B2(n169), .A(n193), .ZN(n453) );
  NAND2_X1 U442 ( .A1(\mem[4][23] ), .A2(n732), .ZN(n193) );
  OAI21_X1 U443 ( .B1(n751), .B2(n169), .A(n194), .ZN(n454) );
  NAND2_X1 U444 ( .A1(\mem[4][24] ), .A2(n731), .ZN(n194) );
  OAI21_X1 U445 ( .B1(n750), .B2(n169), .A(n195), .ZN(n455) );
  NAND2_X1 U446 ( .A1(\mem[4][25] ), .A2(n731), .ZN(n195) );
  OAI21_X1 U447 ( .B1(n749), .B2(n169), .A(n196), .ZN(n456) );
  NAND2_X1 U448 ( .A1(\mem[4][26] ), .A2(n731), .ZN(n196) );
  OAI21_X1 U449 ( .B1(n755), .B2(n203), .A(n224), .ZN(n482) );
  NAND2_X1 U450 ( .A1(\mem[5][20] ), .A2(n730), .ZN(n224) );
  OAI21_X1 U451 ( .B1(n754), .B2(n729), .A(n225), .ZN(n483) );
  NAND2_X1 U452 ( .A1(\mem[5][21] ), .A2(n730), .ZN(n225) );
  OAI21_X1 U453 ( .B1(n753), .B2(n730), .A(n226), .ZN(n484) );
  NAND2_X1 U454 ( .A1(\mem[5][22] ), .A2(n730), .ZN(n226) );
  OAI21_X1 U455 ( .B1(n752), .B2(n729), .A(n227), .ZN(n485) );
  NAND2_X1 U456 ( .A1(\mem[5][23] ), .A2(n730), .ZN(n227) );
  OAI21_X1 U457 ( .B1(n751), .B2(n203), .A(n228), .ZN(n486) );
  NAND2_X1 U458 ( .A1(\mem[5][24] ), .A2(n729), .ZN(n228) );
  OAI21_X1 U459 ( .B1(n750), .B2(n203), .A(n229), .ZN(n487) );
  NAND2_X1 U460 ( .A1(\mem[5][25] ), .A2(n729), .ZN(n229) );
  OAI21_X1 U461 ( .B1(n749), .B2(n203), .A(n230), .ZN(n488) );
  NAND2_X1 U462 ( .A1(\mem[5][26] ), .A2(n729), .ZN(n230) );
  OAI21_X1 U463 ( .B1(n755), .B2(n236), .A(n257), .ZN(n514) );
  NAND2_X1 U464 ( .A1(\mem[6][20] ), .A2(n728), .ZN(n257) );
  OAI21_X1 U465 ( .B1(n754), .B2(n727), .A(n258), .ZN(n515) );
  NAND2_X1 U466 ( .A1(\mem[6][21] ), .A2(n728), .ZN(n258) );
  OAI21_X1 U467 ( .B1(n753), .B2(n728), .A(n259), .ZN(n516) );
  NAND2_X1 U468 ( .A1(\mem[6][22] ), .A2(n728), .ZN(n259) );
  OAI21_X1 U469 ( .B1(n752), .B2(n727), .A(n260), .ZN(n517) );
  NAND2_X1 U470 ( .A1(\mem[6][23] ), .A2(n728), .ZN(n260) );
  OAI21_X1 U471 ( .B1(n751), .B2(n236), .A(n261), .ZN(n518) );
  NAND2_X1 U472 ( .A1(\mem[6][24] ), .A2(n727), .ZN(n261) );
  OAI21_X1 U473 ( .B1(n750), .B2(n236), .A(n262), .ZN(n519) );
  NAND2_X1 U474 ( .A1(\mem[6][25] ), .A2(n727), .ZN(n262) );
  OAI21_X1 U475 ( .B1(n749), .B2(n236), .A(n263), .ZN(n520) );
  NAND2_X1 U476 ( .A1(\mem[6][26] ), .A2(n727), .ZN(n263) );
  OAI21_X1 U477 ( .B1(n755), .B2(n269), .A(n290), .ZN(n546) );
  NAND2_X1 U478 ( .A1(\mem[7][20] ), .A2(n726), .ZN(n290) );
  OAI21_X1 U479 ( .B1(n754), .B2(n725), .A(n291), .ZN(n547) );
  NAND2_X1 U480 ( .A1(\mem[7][21] ), .A2(n726), .ZN(n291) );
  OAI21_X1 U481 ( .B1(n753), .B2(n726), .A(n292), .ZN(n548) );
  NAND2_X1 U482 ( .A1(\mem[7][22] ), .A2(n726), .ZN(n292) );
  OAI21_X1 U483 ( .B1(n752), .B2(n725), .A(n293), .ZN(n549) );
  NAND2_X1 U484 ( .A1(\mem[7][23] ), .A2(n726), .ZN(n293) );
  OAI21_X1 U485 ( .B1(n751), .B2(n269), .A(n294), .ZN(n550) );
  NAND2_X1 U486 ( .A1(\mem[7][24] ), .A2(n725), .ZN(n294) );
  OAI21_X1 U487 ( .B1(n750), .B2(n269), .A(n295), .ZN(n551) );
  NAND2_X1 U488 ( .A1(\mem[7][25] ), .A2(n725), .ZN(n295) );
  OAI21_X1 U489 ( .B1(n749), .B2(n269), .A(n296), .ZN(n552) );
  NAND2_X1 U490 ( .A1(\mem[7][26] ), .A2(n725), .ZN(n296) );
  OAI21_X1 U491 ( .B1(n740), .B2(n775), .A(n37), .ZN(n302) );
  NAND2_X1 U492 ( .A1(\mem[0][0] ), .A2(n36), .ZN(n37) );
  OAI21_X1 U493 ( .B1(n740), .B2(n773), .A(n39), .ZN(n304) );
  NAND2_X1 U494 ( .A1(\mem[0][2] ), .A2(n36), .ZN(n39) );
  OAI21_X1 U495 ( .B1(n740), .B2(n770), .A(n42), .ZN(n307) );
  NAND2_X1 U496 ( .A1(\mem[0][5] ), .A2(n740), .ZN(n42) );
  OAI21_X1 U497 ( .B1(n740), .B2(n769), .A(n43), .ZN(n308) );
  NAND2_X1 U498 ( .A1(\mem[0][6] ), .A2(n739), .ZN(n43) );
  OAI21_X1 U499 ( .B1(n740), .B2(n768), .A(n44), .ZN(n309) );
  NAND2_X1 U500 ( .A1(\mem[0][7] ), .A2(n36), .ZN(n44) );
  OAI21_X1 U501 ( .B1(n739), .B2(n767), .A(n45), .ZN(n310) );
  NAND2_X1 U502 ( .A1(\mem[0][8] ), .A2(n740), .ZN(n45) );
  OAI21_X1 U503 ( .B1(n740), .B2(n766), .A(n46), .ZN(n311) );
  NAND2_X1 U504 ( .A1(\mem[0][9] ), .A2(n36), .ZN(n46) );
  OAI21_X1 U505 ( .B1(n739), .B2(n765), .A(n47), .ZN(n312) );
  NAND2_X1 U506 ( .A1(\mem[0][10] ), .A2(n739), .ZN(n47) );
  OAI21_X1 U507 ( .B1(n740), .B2(n764), .A(n48), .ZN(n313) );
  NAND2_X1 U508 ( .A1(\mem[0][11] ), .A2(n36), .ZN(n48) );
  OAI21_X1 U509 ( .B1(n739), .B2(n763), .A(n49), .ZN(n314) );
  NAND2_X1 U510 ( .A1(\mem[0][12] ), .A2(n36), .ZN(n49) );
  OAI21_X1 U511 ( .B1(n740), .B2(n762), .A(n50), .ZN(n315) );
  NAND2_X1 U512 ( .A1(\mem[0][13] ), .A2(n739), .ZN(n50) );
  OAI21_X1 U513 ( .B1(n739), .B2(n761), .A(n51), .ZN(n316) );
  NAND2_X1 U514 ( .A1(\mem[0][14] ), .A2(n36), .ZN(n51) );
  OAI21_X1 U515 ( .B1(n740), .B2(n760), .A(n52), .ZN(n317) );
  NAND2_X1 U516 ( .A1(\mem[0][15] ), .A2(n36), .ZN(n52) );
  OAI21_X1 U517 ( .B1(n739), .B2(n759), .A(n53), .ZN(n318) );
  NAND2_X1 U518 ( .A1(\mem[0][16] ), .A2(n740), .ZN(n53) );
  OAI21_X1 U519 ( .B1(n739), .B2(n758), .A(n54), .ZN(n319) );
  NAND2_X1 U520 ( .A1(\mem[0][17] ), .A2(n739), .ZN(n54) );
  OAI21_X1 U521 ( .B1(n739), .B2(n757), .A(n55), .ZN(n320) );
  NAND2_X1 U522 ( .A1(\mem[0][18] ), .A2(n739), .ZN(n55) );
  OAI21_X1 U523 ( .B1(n739), .B2(n756), .A(n56), .ZN(n321) );
  NAND2_X1 U524 ( .A1(\mem[0][19] ), .A2(n740), .ZN(n56) );
  OAI21_X1 U525 ( .B1(n739), .B2(n755), .A(n57), .ZN(n322) );
  NAND2_X1 U526 ( .A1(\mem[0][20] ), .A2(n739), .ZN(n57) );
  OAI21_X1 U527 ( .B1(n739), .B2(n754), .A(n58), .ZN(n323) );
  NAND2_X1 U528 ( .A1(\mem[0][21] ), .A2(n739), .ZN(n58) );
  OAI21_X1 U529 ( .B1(n739), .B2(n753), .A(n59), .ZN(n324) );
  NAND2_X1 U530 ( .A1(\mem[0][22] ), .A2(n739), .ZN(n59) );
  OAI21_X1 U531 ( .B1(n739), .B2(n752), .A(n60), .ZN(n325) );
  NAND2_X1 U532 ( .A1(\mem[0][23] ), .A2(n740), .ZN(n60) );
  OAI21_X1 U533 ( .B1(n739), .B2(n751), .A(n61), .ZN(n326) );
  NAND2_X1 U534 ( .A1(\mem[0][24] ), .A2(n36), .ZN(n61) );
  OAI21_X1 U535 ( .B1(n739), .B2(n750), .A(n62), .ZN(n327) );
  NAND2_X1 U536 ( .A1(\mem[0][25] ), .A2(n36), .ZN(n62) );
  OAI21_X1 U537 ( .B1(n739), .B2(n749), .A(n63), .ZN(n328) );
  NAND2_X1 U538 ( .A1(\mem[0][26] ), .A2(n36), .ZN(n63) );
  OAI21_X1 U539 ( .B1(n739), .B2(n748), .A(n64), .ZN(n329) );
  NAND2_X1 U540 ( .A1(\mem[0][27] ), .A2(n36), .ZN(n64) );
  OAI21_X1 U541 ( .B1(n739), .B2(n747), .A(n65), .ZN(n330) );
  NAND2_X1 U542 ( .A1(\mem[0][28] ), .A2(n36), .ZN(n65) );
  INV_X1 U543 ( .A(data_in[0]), .ZN(n775) );
  INV_X1 U544 ( .A(data_in[1]), .ZN(n774) );
  INV_X1 U545 ( .A(data_in[2]), .ZN(n773) );
  INV_X1 U546 ( .A(data_in[3]), .ZN(n772) );
  INV_X1 U547 ( .A(data_in[4]), .ZN(n771) );
  INV_X1 U548 ( .A(data_in[5]), .ZN(n770) );
  INV_X1 U549 ( .A(data_in[6]), .ZN(n769) );
  INV_X1 U550 ( .A(data_in[7]), .ZN(n768) );
  INV_X1 U551 ( .A(data_in[8]), .ZN(n767) );
  INV_X1 U560 ( .A(data_in[9]), .ZN(n766) );
  INV_X1 U561 ( .A(data_in[10]), .ZN(n765) );
  INV_X1 U562 ( .A(data_in[11]), .ZN(n764) );
  INV_X1 U563 ( .A(data_in[12]), .ZN(n763) );
  INV_X1 U564 ( .A(data_in[13]), .ZN(n762) );
  INV_X1 U565 ( .A(data_in[14]), .ZN(n761) );
  INV_X1 U566 ( .A(data_in[15]), .ZN(n760) );
  INV_X1 U567 ( .A(data_in[16]), .ZN(n759) );
  INV_X1 U568 ( .A(data_in[17]), .ZN(n758) );
  INV_X1 U569 ( .A(data_in[18]), .ZN(n757) );
  INV_X1 U570 ( .A(data_in[19]), .ZN(n756) );
  INV_X1 U571 ( .A(data_in[20]), .ZN(n755) );
  INV_X1 U572 ( .A(data_in[21]), .ZN(n754) );
  INV_X1 U573 ( .A(data_in[22]), .ZN(n753) );
  INV_X1 U574 ( .A(data_in[23]), .ZN(n752) );
  INV_X1 U575 ( .A(data_in[24]), .ZN(n751) );
  INV_X1 U576 ( .A(data_in[25]), .ZN(n750) );
  INV_X1 U577 ( .A(data_in[26]), .ZN(n749) );
  INV_X1 U578 ( .A(data_in[27]), .ZN(n748) );
  INV_X1 U579 ( .A(data_in[28]), .ZN(n747) );
  INV_X1 U580 ( .A(data_in[29]), .ZN(n746) );
  INV_X1 U581 ( .A(data_in[30]), .ZN(n745) );
  INV_X1 U582 ( .A(data_in[31]), .ZN(n744) );
  MUX2_X1 U583 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n719), .Z(n1) );
  MUX2_X1 U584 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n719), .Z(n2) );
  MUX2_X1 U585 ( .A(n2), .B(n1), .S(n716), .Z(n3) );
  MUX2_X1 U586 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n719), .Z(n4) );
  MUX2_X1 U587 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n719), .Z(n5) );
  MUX2_X1 U588 ( .A(n5), .B(n4), .S(n717), .Z(n6) );
  MUX2_X1 U589 ( .A(n6), .B(n3), .S(N12), .Z(N44) );
  MUX2_X1 U590 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n719), .Z(n7) );
  MUX2_X1 U591 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n719), .Z(n8) );
  MUX2_X1 U592 ( .A(n8), .B(n7), .S(n717), .Z(n9) );
  MUX2_X1 U593 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n719), .Z(n10) );
  MUX2_X1 U594 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n719), .Z(n11) );
  MUX2_X1 U595 ( .A(n11), .B(n10), .S(n718), .Z(n12) );
  MUX2_X1 U596 ( .A(n12), .B(n9), .S(N12), .Z(N43) );
  MUX2_X1 U597 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n720), .Z(n13) );
  MUX2_X1 U598 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n720), .Z(n14) );
  MUX2_X1 U599 ( .A(n14), .B(n13), .S(n716), .Z(n15) );
  MUX2_X1 U600 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n720), .Z(n16) );
  MUX2_X1 U601 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n720), .Z(n17) );
  MUX2_X1 U602 ( .A(n17), .B(n16), .S(n716), .Z(n18) );
  MUX2_X1 U603 ( .A(n18), .B(n15), .S(N12), .Z(N42) );
  MUX2_X1 U604 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n720), .Z(n19) );
  MUX2_X1 U605 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n720), .Z(n20) );
  MUX2_X1 U606 ( .A(n20), .B(n19), .S(n716), .Z(n21) );
  MUX2_X1 U607 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n720), .Z(n22) );
  MUX2_X1 U608 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n720), .Z(n23) );
  MUX2_X1 U609 ( .A(n23), .B(n22), .S(n716), .Z(n24) );
  MUX2_X1 U610 ( .A(n24), .B(n21), .S(N12), .Z(N41) );
  MUX2_X1 U611 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n720), .Z(n25) );
  MUX2_X1 U612 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n720), .Z(n26) );
  MUX2_X1 U613 ( .A(n26), .B(n25), .S(n716), .Z(n27) );
  MUX2_X1 U614 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n720), .Z(n28) );
  MUX2_X1 U615 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n720), .Z(n29) );
  MUX2_X1 U616 ( .A(n29), .B(n28), .S(n716), .Z(n30) );
  MUX2_X1 U617 ( .A(n30), .B(n27), .S(N12), .Z(N40) );
  MUX2_X1 U618 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n721), .Z(n31) );
  MUX2_X1 U619 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n721), .Z(n32) );
  MUX2_X1 U620 ( .A(n32), .B(n31), .S(n716), .Z(n33) );
  MUX2_X1 U621 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n721), .Z(n34) );
  MUX2_X1 U622 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n721), .Z(n35) );
  MUX2_X1 U623 ( .A(n35), .B(n34), .S(n716), .Z(n558) );
  MUX2_X1 U624 ( .A(n558), .B(n33), .S(N12), .Z(N39) );
  MUX2_X1 U625 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n721), .Z(n559) );
  MUX2_X1 U626 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n721), .Z(n560) );
  MUX2_X1 U627 ( .A(n560), .B(n559), .S(n716), .Z(n561) );
  MUX2_X1 U628 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n721), .Z(n562) );
  MUX2_X1 U629 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n721), .Z(n563) );
  MUX2_X1 U630 ( .A(n563), .B(n562), .S(n716), .Z(n564) );
  MUX2_X1 U631 ( .A(n564), .B(n561), .S(N12), .Z(N38) );
  MUX2_X1 U632 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n721), .Z(n565) );
  MUX2_X1 U633 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n721), .Z(n566) );
  MUX2_X1 U634 ( .A(n566), .B(n565), .S(n716), .Z(n567) );
  MUX2_X1 U635 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n721), .Z(n568) );
  MUX2_X1 U636 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n721), .Z(n569) );
  MUX2_X1 U637 ( .A(n569), .B(n568), .S(n716), .Z(n570) );
  MUX2_X1 U638 ( .A(n570), .B(n567), .S(N12), .Z(N37) );
  MUX2_X1 U639 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n722), .Z(n571) );
  MUX2_X1 U640 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n722), .Z(n572) );
  MUX2_X1 U641 ( .A(n572), .B(n571), .S(n717), .Z(n573) );
  MUX2_X1 U642 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n722), .Z(n574) );
  MUX2_X1 U643 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n722), .Z(n575) );
  MUX2_X1 U644 ( .A(n575), .B(n574), .S(n717), .Z(n576) );
  MUX2_X1 U645 ( .A(n576), .B(n573), .S(n715), .Z(N36) );
  MUX2_X1 U646 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n722), .Z(n577) );
  MUX2_X1 U647 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n722), .Z(n578) );
  MUX2_X1 U648 ( .A(n578), .B(n577), .S(n717), .Z(n579) );
  MUX2_X1 U649 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n722), .Z(n580) );
  MUX2_X1 U650 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n722), .Z(n581) );
  MUX2_X1 U651 ( .A(n581), .B(n580), .S(n717), .Z(n582) );
  MUX2_X1 U652 ( .A(n582), .B(n579), .S(n715), .Z(N35) );
  MUX2_X1 U653 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n722), .Z(n583) );
  MUX2_X1 U654 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n722), .Z(n584) );
  MUX2_X1 U655 ( .A(n584), .B(n583), .S(n717), .Z(n585) );
  MUX2_X1 U656 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n722), .Z(n586) );
  MUX2_X1 U657 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n722), .Z(n587) );
  MUX2_X1 U658 ( .A(n587), .B(n586), .S(n717), .Z(n588) );
  MUX2_X1 U659 ( .A(n588), .B(n585), .S(n715), .Z(N34) );
  MUX2_X1 U660 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n723), .Z(n589) );
  MUX2_X1 U661 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n723), .Z(n590) );
  MUX2_X1 U662 ( .A(n590), .B(n589), .S(n717), .Z(n591) );
  MUX2_X1 U663 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n723), .Z(n592) );
  MUX2_X1 U664 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n723), .Z(n593) );
  MUX2_X1 U665 ( .A(n593), .B(n592), .S(n717), .Z(n594) );
  MUX2_X1 U666 ( .A(n594), .B(n591), .S(n715), .Z(N33) );
  MUX2_X1 U667 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n723), .Z(n595) );
  MUX2_X1 U668 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n723), .Z(n596) );
  MUX2_X1 U669 ( .A(n596), .B(n595), .S(n717), .Z(n597) );
  MUX2_X1 U670 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n723), .Z(n598) );
  MUX2_X1 U671 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n723), .Z(n599) );
  MUX2_X1 U672 ( .A(n599), .B(n598), .S(n717), .Z(n600) );
  MUX2_X1 U673 ( .A(n600), .B(n597), .S(n715), .Z(N32) );
  MUX2_X1 U674 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n723), .Z(n601) );
  MUX2_X1 U675 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n723), .Z(n602) );
  MUX2_X1 U676 ( .A(n602), .B(n601), .S(n717), .Z(n603) );
  MUX2_X1 U677 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n723), .Z(n604) );
  MUX2_X1 U678 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n723), .Z(n605) );
  MUX2_X1 U679 ( .A(n605), .B(n604), .S(n717), .Z(n606) );
  MUX2_X1 U680 ( .A(n606), .B(n603), .S(n715), .Z(N31) );
  MUX2_X1 U681 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n724), .Z(n607) );
  MUX2_X1 U682 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(N10), .Z(n608) );
  MUX2_X1 U683 ( .A(n608), .B(n607), .S(n718), .Z(n609) );
  MUX2_X1 U684 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(N10), .Z(n610) );
  MUX2_X1 U685 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(N10), .Z(n611) );
  MUX2_X1 U686 ( .A(n611), .B(n610), .S(n718), .Z(n612) );
  MUX2_X1 U687 ( .A(n612), .B(n609), .S(n715), .Z(N30) );
  MUX2_X1 U688 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(N10), .Z(n613) );
  MUX2_X1 U689 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(N10), .Z(n614) );
  MUX2_X1 U690 ( .A(n614), .B(n613), .S(n718), .Z(n615) );
  MUX2_X1 U691 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(N10), .Z(n616) );
  MUX2_X1 U692 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n724), .Z(n617) );
  MUX2_X1 U693 ( .A(n617), .B(n616), .S(n718), .Z(n618) );
  MUX2_X1 U694 ( .A(n618), .B(n615), .S(n715), .Z(N29) );
  MUX2_X1 U695 ( .A(\mem[6][16] ), .B(\mem[7][16] ), .S(N10), .Z(n619) );
  MUX2_X1 U696 ( .A(\mem[4][16] ), .B(\mem[5][16] ), .S(N10), .Z(n620) );
  MUX2_X1 U697 ( .A(n620), .B(n619), .S(n718), .Z(n621) );
  MUX2_X1 U698 ( .A(\mem[2][16] ), .B(\mem[3][16] ), .S(N10), .Z(n622) );
  MUX2_X1 U699 ( .A(\mem[0][16] ), .B(\mem[1][16] ), .S(n724), .Z(n623) );
  MUX2_X1 U700 ( .A(n623), .B(n622), .S(n718), .Z(n624) );
  MUX2_X1 U701 ( .A(n624), .B(n621), .S(n715), .Z(N28) );
  MUX2_X1 U702 ( .A(\mem[6][17] ), .B(\mem[7][17] ), .S(n724), .Z(n625) );
  MUX2_X1 U703 ( .A(\mem[4][17] ), .B(\mem[5][17] ), .S(n723), .Z(n626) );
  MUX2_X1 U704 ( .A(n626), .B(n625), .S(n718), .Z(n627) );
  MUX2_X1 U705 ( .A(\mem[2][17] ), .B(\mem[3][17] ), .S(n720), .Z(n628) );
  MUX2_X1 U706 ( .A(\mem[0][17] ), .B(\mem[1][17] ), .S(n724), .Z(n629) );
  MUX2_X1 U707 ( .A(n629), .B(n628), .S(n718), .Z(n630) );
  MUX2_X1 U708 ( .A(n630), .B(n627), .S(n715), .Z(N27) );
  MUX2_X1 U709 ( .A(\mem[6][18] ), .B(\mem[7][18] ), .S(n721), .Z(n631) );
  MUX2_X1 U710 ( .A(\mem[4][18] ), .B(\mem[5][18] ), .S(n723), .Z(n632) );
  MUX2_X1 U711 ( .A(n632), .B(n631), .S(n718), .Z(n633) );
  MUX2_X1 U712 ( .A(\mem[2][18] ), .B(\mem[3][18] ), .S(n721), .Z(n634) );
  MUX2_X1 U713 ( .A(\mem[0][18] ), .B(\mem[1][18] ), .S(n724), .Z(n635) );
  MUX2_X1 U714 ( .A(n635), .B(n634), .S(n718), .Z(n636) );
  MUX2_X1 U715 ( .A(n636), .B(n633), .S(n715), .Z(N26) );
  MUX2_X1 U716 ( .A(\mem[6][19] ), .B(\mem[7][19] ), .S(N10), .Z(n637) );
  MUX2_X1 U717 ( .A(\mem[4][19] ), .B(\mem[5][19] ), .S(n724), .Z(n638) );
  MUX2_X1 U718 ( .A(n638), .B(n637), .S(n718), .Z(n639) );
  MUX2_X1 U719 ( .A(\mem[2][19] ), .B(\mem[3][19] ), .S(n722), .Z(n640) );
  MUX2_X1 U720 ( .A(\mem[0][19] ), .B(\mem[1][19] ), .S(N10), .Z(n641) );
  MUX2_X1 U721 ( .A(n641), .B(n640), .S(n718), .Z(n642) );
  MUX2_X1 U722 ( .A(n642), .B(n639), .S(N12), .Z(N25) );
  MUX2_X1 U723 ( .A(\mem[6][20] ), .B(\mem[7][20] ), .S(n719), .Z(n643) );
  MUX2_X1 U724 ( .A(\mem[4][20] ), .B(\mem[5][20] ), .S(n724), .Z(n644) );
  MUX2_X1 U725 ( .A(n644), .B(n643), .S(n716), .Z(n645) );
  MUX2_X1 U726 ( .A(\mem[2][20] ), .B(\mem[3][20] ), .S(n724), .Z(n646) );
  MUX2_X1 U727 ( .A(\mem[0][20] ), .B(\mem[1][20] ), .S(n724), .Z(n647) );
  MUX2_X1 U728 ( .A(n647), .B(n646), .S(N11), .Z(n648) );
  MUX2_X1 U729 ( .A(n648), .B(n645), .S(n715), .Z(N24) );
  MUX2_X1 U730 ( .A(\mem[6][21] ), .B(\mem[7][21] ), .S(n719), .Z(n649) );
  MUX2_X1 U731 ( .A(\mem[4][21] ), .B(\mem[5][21] ), .S(n724), .Z(n650) );
  MUX2_X1 U732 ( .A(n650), .B(n649), .S(n717), .Z(n651) );
  MUX2_X1 U733 ( .A(\mem[2][21] ), .B(\mem[3][21] ), .S(n724), .Z(n652) );
  MUX2_X1 U734 ( .A(\mem[0][21] ), .B(\mem[1][21] ), .S(n724), .Z(n653) );
  MUX2_X1 U735 ( .A(n653), .B(n652), .S(N11), .Z(n654) );
  MUX2_X1 U736 ( .A(n654), .B(n651), .S(n715), .Z(N23) );
  MUX2_X1 U737 ( .A(\mem[6][22] ), .B(\mem[7][22] ), .S(n719), .Z(n655) );
  MUX2_X1 U738 ( .A(\mem[4][22] ), .B(\mem[5][22] ), .S(n724), .Z(n656) );
  MUX2_X1 U739 ( .A(n656), .B(n655), .S(n718), .Z(n657) );
  MUX2_X1 U740 ( .A(\mem[2][22] ), .B(\mem[3][22] ), .S(n724), .Z(n658) );
  MUX2_X1 U741 ( .A(\mem[0][22] ), .B(\mem[1][22] ), .S(n724), .Z(n659) );
  MUX2_X1 U742 ( .A(n659), .B(n658), .S(N11), .Z(n660) );
  MUX2_X1 U743 ( .A(n660), .B(n657), .S(n715), .Z(N22) );
  MUX2_X1 U744 ( .A(\mem[6][23] ), .B(\mem[7][23] ), .S(n719), .Z(n661) );
  MUX2_X1 U745 ( .A(\mem[4][23] ), .B(\mem[5][23] ), .S(n723), .Z(n662) );
  MUX2_X1 U746 ( .A(n662), .B(n661), .S(N11), .Z(n663) );
  MUX2_X1 U747 ( .A(\mem[2][23] ), .B(\mem[3][23] ), .S(n723), .Z(n664) );
  MUX2_X1 U748 ( .A(\mem[0][23] ), .B(\mem[1][23] ), .S(n722), .Z(n665) );
  MUX2_X1 U749 ( .A(n665), .B(n664), .S(N11), .Z(n666) );
  MUX2_X1 U750 ( .A(n666), .B(n663), .S(n715), .Z(N21) );
  MUX2_X1 U751 ( .A(\mem[6][24] ), .B(\mem[7][24] ), .S(n724), .Z(n667) );
  MUX2_X1 U752 ( .A(\mem[4][24] ), .B(\mem[5][24] ), .S(n722), .Z(n668) );
  MUX2_X1 U753 ( .A(n668), .B(n667), .S(N11), .Z(n669) );
  MUX2_X1 U754 ( .A(\mem[2][24] ), .B(\mem[3][24] ), .S(n721), .Z(n670) );
  MUX2_X1 U755 ( .A(\mem[0][24] ), .B(\mem[1][24] ), .S(n721), .Z(n671) );
  MUX2_X1 U756 ( .A(n671), .B(n670), .S(N11), .Z(n672) );
  MUX2_X1 U757 ( .A(n672), .B(n669), .S(n715), .Z(N20) );
  MUX2_X1 U758 ( .A(\mem[6][25] ), .B(\mem[7][25] ), .S(n720), .Z(n673) );
  MUX2_X1 U759 ( .A(\mem[4][25] ), .B(\mem[5][25] ), .S(n721), .Z(n674) );
  MUX2_X1 U760 ( .A(n674), .B(n673), .S(N11), .Z(n675) );
  MUX2_X1 U761 ( .A(\mem[2][25] ), .B(\mem[3][25] ), .S(n719), .Z(n676) );
  MUX2_X1 U762 ( .A(\mem[0][25] ), .B(\mem[1][25] ), .S(n720), .Z(n677) );
  MUX2_X1 U763 ( .A(n677), .B(n676), .S(N11), .Z(n678) );
  MUX2_X1 U764 ( .A(n678), .B(n675), .S(n715), .Z(N19) );
  MUX2_X1 U765 ( .A(\mem[6][26] ), .B(\mem[7][26] ), .S(n720), .Z(n679) );
  MUX2_X1 U766 ( .A(\mem[4][26] ), .B(\mem[5][26] ), .S(n720), .Z(n680) );
  MUX2_X1 U767 ( .A(n680), .B(n679), .S(n716), .Z(n681) );
  MUX2_X1 U768 ( .A(\mem[2][26] ), .B(\mem[3][26] ), .S(n723), .Z(n682) );
  MUX2_X1 U769 ( .A(\mem[0][26] ), .B(\mem[1][26] ), .S(n722), .Z(n683) );
  MUX2_X1 U770 ( .A(n683), .B(n682), .S(n718), .Z(n684) );
  MUX2_X1 U771 ( .A(n684), .B(n681), .S(n715), .Z(N18) );
  MUX2_X1 U772 ( .A(\mem[6][27] ), .B(\mem[7][27] ), .S(n722), .Z(n685) );
  MUX2_X1 U773 ( .A(\mem[4][27] ), .B(\mem[5][27] ), .S(n719), .Z(n686) );
  MUX2_X1 U774 ( .A(n686), .B(n685), .S(n717), .Z(n687) );
  MUX2_X1 U775 ( .A(\mem[2][27] ), .B(\mem[3][27] ), .S(n722), .Z(n688) );
  MUX2_X1 U776 ( .A(\mem[0][27] ), .B(\mem[1][27] ), .S(n721), .Z(n689) );
  MUX2_X1 U777 ( .A(n689), .B(n688), .S(n716), .Z(n690) );
  MUX2_X1 U778 ( .A(n690), .B(n687), .S(n715), .Z(N17) );
  MUX2_X1 U779 ( .A(\mem[6][28] ), .B(\mem[7][28] ), .S(n719), .Z(n691) );
  MUX2_X1 U780 ( .A(\mem[4][28] ), .B(\mem[5][28] ), .S(n723), .Z(n692) );
  MUX2_X1 U781 ( .A(n692), .B(n691), .S(n718), .Z(n693) );
  MUX2_X1 U782 ( .A(\mem[2][28] ), .B(\mem[3][28] ), .S(n720), .Z(n694) );
  MUX2_X1 U783 ( .A(\mem[0][28] ), .B(\mem[1][28] ), .S(n720), .Z(n695) );
  MUX2_X1 U784 ( .A(n695), .B(n694), .S(n717), .Z(n696) );
  MUX2_X1 U785 ( .A(n696), .B(n693), .S(n715), .Z(N16) );
  MUX2_X1 U786 ( .A(\mem[6][29] ), .B(\mem[7][29] ), .S(n724), .Z(n697) );
  MUX2_X1 U787 ( .A(\mem[4][29] ), .B(\mem[5][29] ), .S(n723), .Z(n698) );
  MUX2_X1 U788 ( .A(n698), .B(n697), .S(n716), .Z(n699) );
  MUX2_X1 U789 ( .A(\mem[2][29] ), .B(\mem[3][29] ), .S(n721), .Z(n700) );
  MUX2_X1 U790 ( .A(\mem[0][29] ), .B(\mem[1][29] ), .S(n721), .Z(n701) );
  MUX2_X1 U791 ( .A(n701), .B(n700), .S(n718), .Z(n702) );
  MUX2_X1 U792 ( .A(n702), .B(n699), .S(n715), .Z(N15) );
  MUX2_X1 U793 ( .A(\mem[6][30] ), .B(\mem[7][30] ), .S(n724), .Z(n703) );
  MUX2_X1 U794 ( .A(\mem[4][30] ), .B(\mem[5][30] ), .S(n719), .Z(n704) );
  MUX2_X1 U795 ( .A(n704), .B(n703), .S(n717), .Z(n705) );
  MUX2_X1 U796 ( .A(\mem[2][30] ), .B(\mem[3][30] ), .S(n720), .Z(n706) );
  MUX2_X1 U797 ( .A(\mem[0][30] ), .B(\mem[1][30] ), .S(n723), .Z(n707) );
  MUX2_X1 U798 ( .A(n707), .B(n706), .S(N11), .Z(n708) );
  MUX2_X1 U799 ( .A(n708), .B(n705), .S(n715), .Z(N14) );
  MUX2_X1 U800 ( .A(\mem[6][31] ), .B(\mem[7][31] ), .S(n724), .Z(n709) );
  MUX2_X1 U801 ( .A(\mem[4][31] ), .B(\mem[5][31] ), .S(n719), .Z(n710) );
  MUX2_X1 U802 ( .A(n710), .B(n709), .S(n718), .Z(n711) );
  MUX2_X1 U803 ( .A(\mem[2][31] ), .B(\mem[3][31] ), .S(n722), .Z(n712) );
  MUX2_X1 U804 ( .A(\mem[0][31] ), .B(\mem[1][31] ), .S(n722), .Z(n713) );
  MUX2_X1 U805 ( .A(n713), .B(n712), .S(n716), .Z(n714) );
  MUX2_X1 U806 ( .A(n714), .B(n711), .S(n715), .Z(N13) );
  CLKBUF_X1 U807 ( .A(n724), .Z(n719) );
  CLKBUF_X1 U808 ( .A(n136), .Z(n734) );
  CLKBUF_X1 U809 ( .A(n36), .Z(n740) );
endmodule


module datapath_DW_mult_tc_8 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n4, n5, n6, n7, n10, n11, n12, n13, n15, n16, n17, n18, n19, n21,
         n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34, n35, n36, n37,
         n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n51, n54, n56, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n84, n85, n86, n87, n88, n90, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n103, n105, n106, n107, n108, n109, n110,
         n114, n116, n117, n118, n119, n122, n123, n124, n125, n127, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n143, n144, n145, n146, n147, n148, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n180, n182, n183, n184, n185, n188, n189, n190,
         n191, n192, n193, n195, n196, n197, n198, n199, n200, n201, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n218, n219, n220, n221, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n244, n246, n247, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n259, n261, n262, n264, n266, n267, n268,
         n270, n272, n273, n274, n275, n276, n278, n280, n281, n282, n283,
         n284, n286, n288, n289, n290, n291, n292, n294, n296, n297, n298,
         n299, n301, n306, n308, n312, n313, n314, n315, n316, n324, n326,
         n328, n330, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n545, n546, n548, n549, n551, n552,
         n554, n555, n557, n558, n560, n561, n563, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033;
  assign product[31] = n84;

  FA_X1 U364 ( .A(n575), .B(n338), .CI(n590), .CO(n334), .S(n335) );
  FA_X1 U365 ( .A(n339), .B(n576), .CI(n342), .CO(n336), .S(n337) );
  FA_X1 U367 ( .A(n346), .B(n577), .CI(n343), .CO(n340), .S(n341) );
  FA_X1 U368 ( .A(n591), .B(n348), .CI(n606), .CO(n342), .S(n343) );
  FA_X1 U369 ( .A(n347), .B(n354), .CI(n352), .CO(n344), .S(n345) );
  FA_X1 U370 ( .A(n578), .B(n592), .CI(n349), .CO(n346), .S(n347) );
  FA_X1 U372 ( .A(n358), .B(n355), .CI(n353), .CO(n350), .S(n351) );
  FA_X1 U373 ( .A(n362), .B(n607), .CI(n360), .CO(n352), .S(n353) );
  FA_X1 U374 ( .A(n593), .B(n579), .CI(n622), .CO(n354), .S(n355) );
  FA_X1 U375 ( .A(n359), .B(n361), .CI(n366), .CO(n356), .S(n357) );
  FA_X1 U376 ( .A(n370), .B(n363), .CI(n368), .CO(n358), .S(n359) );
  FA_X1 U377 ( .A(n580), .B(n594), .CI(n608), .CO(n360), .S(n361) );
  FA_X1 U379 ( .A(n374), .B(n376), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U380 ( .A(n369), .B(n378), .CI(n371), .CO(n366), .S(n367) );
  FA_X1 U381 ( .A(n595), .B(n380), .CI(n609), .CO(n368), .S(n369) );
  FA_X1 U382 ( .A(n623), .B(n581), .CI(n638), .CO(n370), .S(n371) );
  FA_X1 U383 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  FA_X1 U384 ( .A(n379), .B(n388), .CI(n386), .CO(n374), .S(n375) );
  FA_X1 U385 ( .A(n381), .B(n610), .CI(n390), .CO(n376), .S(n377) );
  FA_X1 U386 ( .A(n624), .B(n596), .CI(n582), .CO(n378), .S(n379) );
  FA_X1 U388 ( .A(n394), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U389 ( .A(n391), .B(n389), .CI(n396), .CO(n384), .S(n385) );
  FA_X1 U390 ( .A(n400), .B(n625), .CI(n398), .CO(n386), .S(n387) );
  FA_X1 U391 ( .A(n597), .B(n639), .CI(n611), .CO(n388), .S(n389) );
  FA_X1 U392 ( .A(n654), .B(n583), .CI(n999), .CO(n390), .S(n391) );
  FA_X1 U393 ( .A(n406), .B(n397), .CI(n395), .CO(n392), .S(n393) );
  FA_X1 U394 ( .A(n410), .B(n399), .CI(n408), .CO(n394), .S(n395) );
  FA_X1 U395 ( .A(n412), .B(n414), .CI(n401), .CO(n396), .S(n397) );
  FA_X1 U396 ( .A(n584), .B(n598), .CI(n403), .CO(n398), .S(n399) );
  FA_X1 U397 ( .A(n626), .B(n612), .CI(n640), .CO(n400), .S(n401) );
  FA_X1 U399 ( .A(n418), .B(n409), .CI(n407), .CO(n404), .S(n405) );
  FA_X1 U400 ( .A(n411), .B(n422), .CI(n420), .CO(n406), .S(n407) );
  FA_X1 U401 ( .A(n413), .B(n424), .CI(n415), .CO(n408), .S(n409) );
  FA_X1 U402 ( .A(n613), .B(n627), .CI(n426), .CO(n410), .S(n411) );
  FA_X1 U403 ( .A(n599), .B(n655), .CI(n641), .CO(n412), .S(n413) );
  FA_X1 U404 ( .A(n428), .B(n585), .CI(n670), .CO(n414), .S(n415) );
  FA_X1 U405 ( .A(n432), .B(n421), .CI(n419), .CO(n416), .S(n417) );
  FA_X1 U406 ( .A(n423), .B(n436), .CI(n434), .CO(n418), .S(n419) );
  FA_X1 U409 ( .A(n642), .B(n628), .CI(n600), .CO(n424), .S(n425) );
  FA_X1 U410 ( .A(n614), .B(n586), .CI(n656), .CO(n426), .S(n427) );
  FA_X1 U414 ( .A(n439), .B(n452), .CI(n441), .CO(n434), .S(n435) );
  FA_X1 U415 ( .A(n443), .B(n456), .CI(n454), .CO(n436), .S(n437) );
  FA_X1 U416 ( .A(n671), .B(n615), .CI(n657), .CO(n438), .S(n439) );
  FA_X1 U417 ( .A(n587), .B(n629), .CI(n686), .CO(n440), .S(n441) );
  FA_X1 U420 ( .A(n449), .B(n460), .CI(n447), .CO(n444), .S(n445) );
  FA_X1 U421 ( .A(n462), .B(n455), .CI(n451), .CO(n446), .S(n447) );
  FA_X1 U422 ( .A(n464), .B(n466), .CI(n453), .CO(n448), .S(n449) );
  FA_X1 U423 ( .A(n457), .B(n672), .CI(n468), .CO(n450), .S(n451) );
  FA_X1 U424 ( .A(n687), .B(n630), .CI(n658), .CO(n452), .S(n453) );
  FA_X1 U425 ( .A(n602), .B(n644), .CI(n616), .CO(n454), .S(n455) );
  HA_X1 U426 ( .A(n566), .B(n588), .CO(n456), .S(n457) );
  FA_X1 U427 ( .A(n463), .B(n472), .CI(n461), .CO(n458), .S(n459) );
  FA_X1 U428 ( .A(n465), .B(n467), .CI(n474), .CO(n460), .S(n461) );
  FA_X1 U429 ( .A(n476), .B(n478), .CI(n469), .CO(n462), .S(n463) );
  FA_X1 U430 ( .A(n645), .B(n659), .CI(n480), .CO(n464), .S(n465) );
  FA_X1 U431 ( .A(n603), .B(n673), .CI(n631), .CO(n466), .S(n467) );
  FA_X1 U432 ( .A(n617), .B(n589), .CI(n688), .CO(n468), .S(n469) );
  FA_X1 U435 ( .A(n490), .B(n481), .CI(n488), .CO(n474), .S(n475) );
  FA_X1 U436 ( .A(n618), .B(n660), .CI(n632), .CO(n476), .S(n477) );
  FA_X1 U437 ( .A(n674), .B(n646), .CI(n689), .CO(n478), .S(n479) );
  HA_X1 U438 ( .A(n604), .B(n567), .CO(n480), .S(n481) );
  FA_X1 U439 ( .A(n487), .B(n494), .CI(n485), .CO(n482), .S(n483) );
  FA_X1 U440 ( .A(n489), .B(n491), .CI(n496), .CO(n484), .S(n485) );
  FA_X1 U441 ( .A(n500), .B(n661), .CI(n498), .CO(n486), .S(n487) );
  FA_X1 U442 ( .A(n647), .B(n619), .CI(n675), .CO(n488), .S(n489) );
  FA_X1 U443 ( .A(n633), .B(n605), .CI(n690), .CO(n490), .S(n491) );
  FA_X1 U444 ( .A(n504), .B(n497), .CI(n495), .CO(n492), .S(n493) );
  FA_X1 U445 ( .A(n506), .B(n508), .CI(n499), .CO(n494), .S(n495) );
  FA_X1 U446 ( .A(n648), .B(n676), .CI(n501), .CO(n496), .S(n497) );
  FA_X1 U447 ( .A(n634), .B(n662), .CI(n691), .CO(n498), .S(n499) );
  HA_X1 U448 ( .A(n620), .B(n568), .CO(n500), .S(n501) );
  FA_X1 U449 ( .A(n512), .B(n507), .CI(n505), .CO(n502), .S(n503) );
  FA_X1 U450 ( .A(n514), .B(n516), .CI(n509), .CO(n504), .S(n505) );
  FA_X1 U451 ( .A(n635), .B(n677), .CI(n663), .CO(n506), .S(n507) );
  FA_X1 U452 ( .A(n649), .B(n621), .CI(n692), .CO(n508), .S(n509) );
  FA_X1 U453 ( .A(n515), .B(n520), .CI(n513), .CO(n510), .S(n511) );
  FA_X1 U454 ( .A(n517), .B(n693), .CI(n522), .CO(n512), .S(n513) );
  FA_X1 U455 ( .A(n650), .B(n664), .CI(n678), .CO(n514), .S(n515) );
  HA_X1 U456 ( .A(n569), .B(n636), .CO(n516), .S(n517) );
  FA_X1 U457 ( .A(n523), .B(n526), .CI(n521), .CO(n518), .S(n519) );
  FA_X1 U458 ( .A(n651), .B(n679), .CI(n528), .CO(n520), .S(n521) );
  FA_X1 U459 ( .A(n665), .B(n637), .CI(n694), .CO(n522), .S(n523) );
  FA_X1 U460 ( .A(n532), .B(n529), .CI(n527), .CO(n524), .S(n525) );
  FA_X1 U461 ( .A(n666), .B(n695), .CI(n680), .CO(n526), .S(n527) );
  HA_X1 U462 ( .A(n570), .B(n652), .CO(n528), .S(n529) );
  FA_X1 U463 ( .A(n536), .B(n667), .CI(n533), .CO(n530), .S(n531) );
  FA_X1 U464 ( .A(n696), .B(n653), .CI(n681), .CO(n532), .S(n533) );
  FA_X1 U465 ( .A(n682), .B(n697), .CI(n537), .CO(n534), .S(n535) );
  HA_X1 U466 ( .A(n668), .B(n571), .CO(n536), .S(n537) );
  FA_X1 U467 ( .A(n698), .B(n669), .CI(n683), .CO(n538), .S(n539) );
  HA_X1 U468 ( .A(n684), .B(n699), .CO(n540), .S(n541) );
  CLKBUF_X2 U822 ( .A(b[13]), .Z(n840) );
  CLKBUF_X1 U823 ( .A(n276), .Z(n953) );
  BUF_X2 U824 ( .A(n874), .Z(n21) );
  BUF_X2 U825 ( .A(n870), .Z(n45) );
  XNOR2_X1 U826 ( .A(n954), .B(n486), .ZN(n473) );
  XNOR2_X1 U827 ( .A(n479), .B(n477), .ZN(n954) );
  NOR2_X2 U828 ( .A1(n431), .A2(n444), .ZN(n227) );
  BUF_X2 U829 ( .A(n864), .Z(n36) );
  BUF_X2 U830 ( .A(n872), .Z(n34) );
  XNOR2_X2 U831 ( .A(n448), .B(n955), .ZN(n433) );
  XNOR2_X1 U832 ( .A(n437), .B(n450), .ZN(n955) );
  CLKBUF_X1 U833 ( .A(b[0]), .Z(n49) );
  BUF_X2 U834 ( .A(n49), .Z(n956) );
  CLKBUF_X3 U835 ( .A(b[2]), .Z(n851) );
  CLKBUF_X3 U836 ( .A(b[15]), .Z(n838) );
  CLKBUF_X3 U837 ( .A(n875), .Z(n16) );
  CLKBUF_X3 U838 ( .A(n866), .Z(n23) );
  XOR2_X1 U839 ( .A(n442), .B(n429), .Z(n957) );
  XOR2_X1 U840 ( .A(n440), .B(n957), .Z(n423) );
  NAND2_X1 U841 ( .A1(n440), .A2(n442), .ZN(n958) );
  NAND2_X1 U842 ( .A1(n440), .A2(n429), .ZN(n959) );
  NAND2_X1 U843 ( .A1(n442), .A2(n429), .ZN(n960) );
  NAND3_X1 U844 ( .A1(n958), .A2(n959), .A3(n960), .ZN(n422) );
  XOR2_X1 U845 ( .A(n427), .B(n438), .Z(n961) );
  XOR2_X1 U846 ( .A(n425), .B(n961), .Z(n421) );
  NAND2_X1 U847 ( .A1(n425), .A2(n427), .ZN(n962) );
  NAND2_X1 U848 ( .A1(n425), .A2(n438), .ZN(n963) );
  NAND2_X1 U849 ( .A1(n427), .A2(n438), .ZN(n964) );
  NAND3_X1 U850 ( .A1(n962), .A2(n963), .A3(n964), .ZN(n420) );
  NAND2_X1 U851 ( .A1(n448), .A2(n437), .ZN(n965) );
  NAND2_X1 U852 ( .A1(n448), .A2(n450), .ZN(n966) );
  NAND2_X1 U853 ( .A1(n437), .A2(n450), .ZN(n967) );
  NAND3_X1 U854 ( .A1(n965), .A2(n966), .A3(n967), .ZN(n432) );
  BUF_X4 U855 ( .A(a[3]), .Z(n7) );
  BUF_X2 U856 ( .A(a[9]), .Z(n25) );
  BUF_X2 U857 ( .A(n865), .Z(n29) );
  BUF_X2 U858 ( .A(n206), .Z(n1026) );
  OR2_X1 U859 ( .A1(n503), .A2(n510), .ZN(n968) );
  XNOR2_X1 U860 ( .A(n106), .B(n969), .ZN(product[29]) );
  AND2_X1 U861 ( .A1(n971), .A2(n105), .ZN(n969) );
  OAI21_X1 U862 ( .B1(n199), .B2(n205), .A(n200), .ZN(n970) );
  NOR2_X2 U863 ( .A1(n383), .A2(n392), .ZN(n199) );
  BUF_X1 U864 ( .A(n841), .Z(n1030) );
  BUF_X2 U865 ( .A(b[10]), .Z(n843) );
  BUF_X2 U866 ( .A(b[6]), .Z(n847) );
  BUF_X2 U867 ( .A(n863), .Z(n41) );
  OAI21_X1 U868 ( .B1(n199), .B2(n205), .A(n200), .ZN(n198) );
  OAI22_X1 U869 ( .A1(n48), .A2(n703), .B1(n46), .B2(n702), .ZN(n332) );
  OR2_X1 U870 ( .A1(n334), .A2(n333), .ZN(n971) );
  OR2_X1 U871 ( .A1(n337), .A2(n340), .ZN(n972) );
  OR2_X1 U872 ( .A1(n574), .A2(n332), .ZN(n973) );
  OR2_X1 U873 ( .A1(n541), .A2(n572), .ZN(n974) );
  AND2_X1 U874 ( .A1(n980), .A2(n301), .ZN(product[1]) );
  OR2_X1 U875 ( .A1(n336), .A2(n335), .ZN(n976) );
  OR2_X1 U876 ( .A1(n535), .A2(n538), .ZN(n977) );
  OR2_X1 U877 ( .A1(n511), .A2(n518), .ZN(n978) );
  OR2_X1 U878 ( .A1(n525), .A2(n530), .ZN(n979) );
  OR2_X1 U879 ( .A1(n701), .A2(n573), .ZN(n980) );
  BUF_X2 U880 ( .A(n841), .Z(n1029) );
  CLKBUF_X3 U881 ( .A(b[1]), .Z(n852) );
  BUF_X1 U882 ( .A(n875), .Z(n15) );
  CLKBUF_X1 U883 ( .A(n991), .Z(n981) );
  OR2_X2 U884 ( .A1(n493), .A2(n502), .ZN(n982) );
  BUF_X2 U885 ( .A(n49), .Z(n1033) );
  AOI21_X1 U886 ( .B1(n970), .B2(n151), .A(n152), .ZN(n983) );
  AOI21_X1 U887 ( .B1(n198), .B2(n151), .A(n152), .ZN(n984) );
  CLKBUF_X1 U888 ( .A(n219), .Z(n985) );
  BUF_X2 U889 ( .A(b[8]), .Z(n845) );
  CLKBUF_X3 U890 ( .A(n876), .Z(n10) );
  CLKBUF_X1 U891 ( .A(n281), .Z(n986) );
  BUF_X2 U892 ( .A(n869), .Z(n5) );
  BUF_X4 U893 ( .A(a[7]), .Z(n19) );
  BUF_X2 U894 ( .A(n868), .Z(n12) );
  BUF_X1 U895 ( .A(n873), .Z(n28) );
  BUF_X2 U896 ( .A(n865), .Z(n30) );
  BUF_X2 U897 ( .A(n869), .Z(n6) );
  CLKBUF_X2 U898 ( .A(n863), .Z(n42) );
  CLKBUF_X3 U899 ( .A(n862), .Z(n47) );
  BUF_X4 U900 ( .A(a[15]), .Z(n43) );
  XNOR2_X1 U901 ( .A(n1), .B(n1029), .ZN(n987) );
  CLKBUF_X1 U902 ( .A(n232), .Z(n988) );
  BUF_X2 U903 ( .A(a[13]), .Z(n989) );
  OAI21_X1 U904 ( .B1(n227), .B2(n233), .A(n228), .ZN(n990) );
  NOR2_X1 U905 ( .A1(n405), .A2(n416), .ZN(n991) );
  NOR2_X1 U906 ( .A1(n405), .A2(n416), .ZN(n211) );
  OR2_X1 U907 ( .A1(n365), .A2(n372), .ZN(n992) );
  XNOR2_X1 U908 ( .A(n31), .B(n847), .ZN(n993) );
  AOI21_X1 U909 ( .B1(n1027), .B2(n251), .A(n244), .ZN(n994) );
  CLKBUF_X1 U910 ( .A(n839), .Z(n995) );
  XNOR2_X1 U911 ( .A(n146), .B(n996), .ZN(product[25]) );
  AND2_X1 U912 ( .A1(n143), .A2(n145), .ZN(n996) );
  BUF_X2 U913 ( .A(n866), .Z(n24) );
  AOI21_X1 U914 ( .B1(n255), .B2(n236), .A(n237), .ZN(n997) );
  OR2_X1 U915 ( .A1(n459), .A2(n470), .ZN(n998) );
  OAI22_X1 U916 ( .A1(n18), .A2(n788), .B1(n16), .B2(n787), .ZN(n999) );
  CLKBUF_X2 U917 ( .A(b[3]), .Z(n850) );
  CLKBUF_X1 U918 ( .A(n218), .Z(n1000) );
  BUF_X2 U919 ( .A(a[11]), .Z(n1001) );
  XNOR2_X1 U920 ( .A(n192), .B(n1002), .ZN(product[21]) );
  AND2_X1 U921 ( .A1(n188), .A2(n191), .ZN(n1002) );
  XNOR2_X1 U922 ( .A(n201), .B(n1003), .ZN(product[20]) );
  AND2_X1 U923 ( .A1(n312), .A2(n200), .ZN(n1003) );
  CLKBUF_X1 U924 ( .A(n284), .Z(n1004) );
  BUF_X2 U925 ( .A(b[9]), .Z(n1005) );
  XNOR2_X1 U926 ( .A(n159), .B(n1006), .ZN(product[24]) );
  AND2_X1 U927 ( .A1(n308), .A2(n158), .ZN(n1006) );
  CLKBUF_X1 U928 ( .A(b[11]), .Z(n842) );
  CLKBUF_X1 U929 ( .A(b[11]), .Z(n1008) );
  CLKBUF_X1 U930 ( .A(b[11]), .Z(n1009) );
  XNOR2_X1 U931 ( .A(n433), .B(n1007), .ZN(n431) );
  XNOR2_X1 U932 ( .A(n446), .B(n435), .ZN(n1007) );
  XNOR2_X1 U933 ( .A(n139), .B(n1010), .ZN(product[26]) );
  AND2_X1 U934 ( .A1(n306), .A2(n138), .ZN(n1010) );
  XOR2_X1 U935 ( .A(n484), .B(n475), .Z(n1011) );
  XOR2_X1 U936 ( .A(n1011), .B(n473), .Z(n471) );
  NAND2_X1 U937 ( .A1(n479), .A2(n477), .ZN(n1012) );
  NAND2_X1 U938 ( .A1(n479), .A2(n486), .ZN(n1013) );
  NAND2_X1 U939 ( .A1(n477), .A2(n486), .ZN(n1014) );
  NAND3_X1 U940 ( .A1(n1012), .A2(n1013), .A3(n1014), .ZN(n472) );
  NAND2_X1 U941 ( .A1(n484), .A2(n475), .ZN(n1015) );
  NAND2_X1 U942 ( .A1(n484), .A2(n473), .ZN(n1016) );
  NAND2_X1 U943 ( .A1(n475), .A2(n473), .ZN(n1017) );
  NAND3_X1 U944 ( .A1(n1015), .A2(n1016), .A3(n1017), .ZN(n470) );
  OR2_X1 U945 ( .A1(n17), .A2(n796), .ZN(n1018) );
  OR2_X1 U946 ( .A1(n15), .A2(n795), .ZN(n1019) );
  NAND2_X1 U947 ( .A1(n1018), .A2(n1019), .ZN(n662) );
  BUF_X2 U948 ( .A(b[5]), .Z(n848) );
  NAND2_X1 U949 ( .A1(n433), .A2(n446), .ZN(n1020) );
  NAND2_X1 U950 ( .A1(n433), .A2(n435), .ZN(n1021) );
  NAND2_X1 U951 ( .A1(n446), .A2(n435), .ZN(n1022) );
  NAND3_X1 U952 ( .A1(n1020), .A2(n1021), .A3(n1022), .ZN(n430) );
  BUF_X2 U953 ( .A(n864), .Z(n35) );
  BUF_X1 U954 ( .A(b[12]), .Z(n841) );
  CLKBUF_X2 U955 ( .A(b[7]), .Z(n846) );
  XNOR2_X1 U956 ( .A(n183), .B(n1023), .ZN(product[22]) );
  AND2_X1 U957 ( .A1(n175), .A2(n182), .ZN(n1023) );
  XNOR2_X1 U958 ( .A(n130), .B(n1024), .ZN(product[27]) );
  AND2_X1 U959 ( .A1(n972), .A2(n129), .ZN(n1024) );
  XNOR2_X1 U960 ( .A(n170), .B(n1025), .ZN(product[23]) );
  AND2_X1 U961 ( .A1(n167), .A2(n169), .ZN(n1025) );
  BUF_X2 U962 ( .A(n867), .Z(n18) );
  BUF_X2 U963 ( .A(b[14]), .Z(n839) );
  BUF_X2 U964 ( .A(b[9]), .Z(n844) );
  OR2_X2 U965 ( .A1(n471), .A2(n482), .ZN(n1027) );
  BUF_X1 U966 ( .A(n841), .Z(n1028) );
  BUF_X4 U967 ( .A(a[5]), .Z(n13) );
  BUF_X2 U968 ( .A(b[4]), .Z(n849) );
  BUF_X4 U969 ( .A(a[1]), .Z(n1) );
  BUF_X2 U970 ( .A(n867), .Z(n17) );
  BUF_X2 U971 ( .A(n49), .Z(n1032) );
  NAND2_X1 U972 ( .A1(n197), .A2(n151), .ZN(n1031) );
  NOR2_X1 U973 ( .A1(n345), .A2(n350), .ZN(n144) );
  NOR2_X1 U974 ( .A1(n373), .A2(n382), .ZN(n190) );
  NOR2_X1 U975 ( .A1(n700), .A2(n685), .ZN(n298) );
  NOR2_X1 U976 ( .A1(n539), .A2(n540), .ZN(n290) );
  BUF_X1 U977 ( .A(n873), .Z(n27) );
  BUF_X1 U978 ( .A(n874), .Z(n22) );
  BUF_X2 U979 ( .A(a[13]), .Z(n37) );
  INV_X1 U980 ( .A(n223), .ZN(n221) );
  BUF_X2 U981 ( .A(n206), .Z(n51) );
  INV_X1 U982 ( .A(n225), .ZN(n223) );
  NOR2_X1 U983 ( .A1(n195), .A2(n190), .ZN(n184) );
  NOR2_X1 U984 ( .A1(n195), .A2(n162), .ZN(n160) );
  NOR2_X1 U985 ( .A1(n195), .A2(n173), .ZN(n171) );
  NOR2_X1 U986 ( .A1(n223), .A2(n1000), .ZN(n214) );
  INV_X1 U987 ( .A(n177), .ZN(n175) );
  INV_X1 U988 ( .A(n195), .ZN(n193) );
  INV_X1 U989 ( .A(n98), .ZN(n96) );
  INV_X1 U990 ( .A(n1031), .ZN(n147) );
  NAND2_X1 U991 ( .A1(n230), .A2(n233), .ZN(n69) );
  NAND2_X1 U992 ( .A1(n313), .A2(n205), .ZN(n65) );
  INV_X1 U993 ( .A(n204), .ZN(n313) );
  XOR2_X1 U994 ( .A(n213), .B(n66), .Z(product[18]) );
  NAND2_X1 U995 ( .A1(n314), .A2(n212), .ZN(n66) );
  INV_X1 U996 ( .A(n981), .ZN(n314) );
  XNOR2_X1 U997 ( .A(n240), .B(n70), .ZN(product[14]) );
  NAND2_X1 U998 ( .A1(n998), .A2(n239), .ZN(n70) );
  XOR2_X1 U999 ( .A(n229), .B(n68), .Z(product[16]) );
  NAND2_X1 U1000 ( .A1(n316), .A2(n228), .ZN(n68) );
  INV_X1 U1001 ( .A(n227), .ZN(n316) );
  INV_X1 U1002 ( .A(n197), .ZN(n195) );
  XOR2_X1 U1003 ( .A(n220), .B(n67), .Z(product[17]) );
  NAND2_X1 U1004 ( .A1(n315), .A2(n985), .ZN(n67) );
  NOR2_X1 U1005 ( .A1(n124), .A2(n100), .ZN(n98) );
  NOR2_X1 U1006 ( .A1(n177), .A2(n166), .ZN(n164) );
  INV_X1 U1007 ( .A(n255), .ZN(n254) );
  INV_X1 U1008 ( .A(n198), .ZN(n196) );
  NAND2_X1 U1009 ( .A1(n164), .A2(n188), .ZN(n162) );
  NAND2_X1 U1010 ( .A1(n188), .A2(n175), .ZN(n173) );
  OAI21_X1 U1011 ( .B1(n196), .B2(n190), .A(n191), .ZN(n185) );
  OAI21_X1 U1012 ( .B1(n196), .B2(n173), .A(n174), .ZN(n172) );
  AOI21_X1 U1013 ( .B1(n189), .B2(n175), .A(n176), .ZN(n174) );
  INV_X1 U1014 ( .A(n178), .ZN(n176) );
  INV_X1 U1015 ( .A(n268), .ZN(n267) );
  INV_X1 U1016 ( .A(n124), .ZN(n122) );
  INV_X1 U1017 ( .A(n992), .ZN(n177) );
  INV_X1 U1018 ( .A(n180), .ZN(n178) );
  NAND2_X1 U1019 ( .A1(n1027), .A2(n250), .ZN(n241) );
  NAND2_X1 U1020 ( .A1(n122), .A2(n976), .ZN(n109) );
  INV_X1 U1021 ( .A(n251), .ZN(n249) );
  INV_X1 U1022 ( .A(n233), .ZN(n231) );
  INV_X1 U1023 ( .A(n205), .ZN(n203) );
  INV_X1 U1024 ( .A(n983), .ZN(n148) );
  INV_X1 U1025 ( .A(n988), .ZN(n230) );
  NAND2_X1 U1026 ( .A1(n982), .A2(n261), .ZN(n73) );
  NAND2_X1 U1027 ( .A1(n978), .A2(n272), .ZN(n75) );
  INV_X1 U1028 ( .A(n272), .ZN(n270) );
  XOR2_X1 U1029 ( .A(n254), .B(n72), .Z(product[12]) );
  XNOR2_X1 U1030 ( .A(n267), .B(n74), .ZN(product[10]) );
  NAND2_X1 U1031 ( .A1(n968), .A2(n266), .ZN(n74) );
  NOR2_X1 U1032 ( .A1(n459), .A2(n470), .ZN(n238) );
  INV_X1 U1033 ( .A(n157), .ZN(n308) );
  INV_X1 U1034 ( .A(n199), .ZN(n312) );
  NAND2_X1 U1035 ( .A1(n445), .A2(n458), .ZN(n233) );
  OAI21_X1 U1036 ( .B1(n256), .B2(n268), .A(n257), .ZN(n255) );
  NAND2_X1 U1037 ( .A1(n982), .A2(n968), .ZN(n256) );
  AOI21_X1 U1038 ( .B1(n982), .B2(n264), .A(n259), .ZN(n257) );
  NOR2_X1 U1039 ( .A1(n393), .A2(n404), .ZN(n204) );
  NOR2_X1 U1040 ( .A1(n445), .A2(n458), .ZN(n232) );
  OAI21_X1 U1041 ( .B1(n196), .B2(n162), .A(n163), .ZN(n161) );
  AOI21_X1 U1042 ( .B1(n164), .B2(n189), .A(n165), .ZN(n163) );
  OAI21_X1 U1043 ( .B1(n178), .B2(n166), .A(n169), .ZN(n165) );
  NOR2_X1 U1044 ( .A1(n190), .A2(n153), .ZN(n151) );
  NAND2_X1 U1045 ( .A1(n135), .A2(n972), .ZN(n124) );
  XNOR2_X1 U1046 ( .A(n247), .B(n71), .ZN(product[13]) );
  OAI21_X1 U1047 ( .B1(n254), .B2(n252), .A(n249), .ZN(n247) );
  INV_X1 U1048 ( .A(n136), .ZN(n134) );
  AOI21_X1 U1049 ( .B1(n123), .B2(n976), .A(n114), .ZN(n110) );
  INV_X1 U1050 ( .A(n99), .ZN(n97) );
  INV_X1 U1051 ( .A(n125), .ZN(n123) );
  NAND2_X1 U1052 ( .A1(n393), .A2(n404), .ZN(n205) );
  INV_X1 U1053 ( .A(n190), .ZN(n188) );
  INV_X1 U1054 ( .A(n191), .ZN(n189) );
  INV_X1 U1055 ( .A(n135), .ZN(n133) );
  INV_X1 U1056 ( .A(n182), .ZN(n180) );
  NAND2_X1 U1057 ( .A1(n431), .A2(n444), .ZN(n228) );
  NAND2_X1 U1058 ( .A1(n405), .A2(n416), .ZN(n212) );
  NAND2_X1 U1059 ( .A1(n976), .A2(n971), .ZN(n100) );
  INV_X1 U1060 ( .A(n167), .ZN(n166) );
  INV_X1 U1061 ( .A(n266), .ZN(n264) );
  NAND2_X1 U1062 ( .A1(n98), .A2(n973), .ZN(n87) );
  INV_X1 U1063 ( .A(n261), .ZN(n259) );
  INV_X1 U1064 ( .A(n144), .ZN(n143) );
  NAND2_X1 U1065 ( .A1(n326), .A2(n283), .ZN(n78) );
  NAND2_X1 U1066 ( .A1(n324), .A2(n275), .ZN(n76) );
  INV_X1 U1067 ( .A(n274), .ZN(n324) );
  NAND2_X1 U1068 ( .A1(n977), .A2(n288), .ZN(n79) );
  NAND2_X1 U1069 ( .A1(n979), .A2(n280), .ZN(n77) );
  XOR2_X1 U1070 ( .A(n117), .B(n56), .Z(product[28]) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n116), .ZN(n56) );
  INV_X1 U1072 ( .A(n280), .ZN(n278) );
  OAI21_X1 U1073 ( .B1(n125), .B2(n100), .A(n101), .ZN(n99) );
  AOI21_X1 U1074 ( .B1(n114), .B2(n971), .A(n103), .ZN(n101) );
  INV_X1 U1075 ( .A(n105), .ZN(n103) );
  INV_X1 U1076 ( .A(n288), .ZN(n286) );
  NOR2_X1 U1077 ( .A1(n351), .A2(n356), .ZN(n157) );
  AOI21_X1 U1078 ( .B1(n136), .B2(n972), .A(n127), .ZN(n125) );
  INV_X1 U1079 ( .A(n129), .ZN(n127) );
  INV_X1 U1080 ( .A(n137), .ZN(n306) );
  XOR2_X1 U1081 ( .A(n93), .B(n54), .Z(product[30]) );
  NAND2_X1 U1082 ( .A1(n973), .A2(n92), .ZN(n54) );
  NOR2_X1 U1083 ( .A1(n357), .A2(n364), .ZN(n168) );
  OAI21_X1 U1084 ( .B1(n276), .B2(n274), .A(n275), .ZN(n273) );
  NAND2_X1 U1085 ( .A1(n373), .A2(n382), .ZN(n191) );
  AOI21_X1 U1086 ( .B1(n99), .B2(n973), .A(n90), .ZN(n88) );
  INV_X1 U1087 ( .A(n92), .ZN(n90) );
  NAND2_X1 U1088 ( .A1(n357), .A2(n364), .ZN(n169) );
  NAND2_X1 U1089 ( .A1(n503), .A2(n510), .ZN(n266) );
  NAND2_X1 U1090 ( .A1(n493), .A2(n502), .ZN(n261) );
  NAND2_X1 U1091 ( .A1(n511), .A2(n518), .ZN(n272) );
  NAND2_X1 U1092 ( .A1(n345), .A2(n350), .ZN(n145) );
  INV_X1 U1093 ( .A(n116), .ZN(n114) );
  NAND2_X1 U1094 ( .A1(n330), .A2(n299), .ZN(n82) );
  INV_X1 U1095 ( .A(n298), .ZN(n330) );
  NAND2_X1 U1096 ( .A1(n328), .A2(n291), .ZN(n80) );
  INV_X1 U1097 ( .A(n290), .ZN(n328) );
  NAND2_X1 U1098 ( .A1(n574), .A2(n332), .ZN(n92) );
  NAND2_X1 U1099 ( .A1(n525), .A2(n530), .ZN(n280) );
  NOR2_X1 U1100 ( .A1(n341), .A2(n344), .ZN(n137) );
  NOR2_X1 U1101 ( .A1(n519), .A2(n524), .ZN(n274) );
  INV_X1 U1102 ( .A(n332), .ZN(n333) );
  XNOR2_X1 U1103 ( .A(n643), .B(n601), .ZN(n443) );
  OR2_X1 U1104 ( .A1(n643), .A2(n601), .ZN(n442) );
  INV_X1 U1105 ( .A(n428), .ZN(n429) );
  NAND2_X1 U1106 ( .A1(n700), .A2(n685), .ZN(n299) );
  NAND2_X1 U1107 ( .A1(n535), .A2(n538), .ZN(n288) );
  NAND2_X1 U1108 ( .A1(n337), .A2(n340), .ZN(n129) );
  NAND2_X1 U1109 ( .A1(n336), .A2(n335), .ZN(n116) );
  NAND2_X1 U1110 ( .A1(n334), .A2(n333), .ZN(n105) );
  NAND2_X1 U1111 ( .A1(n519), .A2(n524), .ZN(n275) );
  NAND2_X1 U1112 ( .A1(n341), .A2(n344), .ZN(n138) );
  NAND2_X1 U1113 ( .A1(n531), .A2(n534), .ZN(n283) );
  OAI22_X1 U1114 ( .A1(n5), .A2(n835), .B1(n834), .B2(n877), .ZN(n700) );
  OAI22_X1 U1115 ( .A1(n12), .A2(n805), .B1(n10), .B2(n804), .ZN(n428) );
  OAI22_X1 U1116 ( .A1(n17), .A2(n788), .B1(n16), .B2(n787), .ZN(n402) );
  OAI22_X1 U1117 ( .A1(n24), .A2(n771), .B1(n22), .B2(n770), .ZN(n380) );
  OAI22_X1 U1118 ( .A1(n42), .A2(n720), .B1(n40), .B2(n719), .ZN(n338) );
  OAI22_X1 U1119 ( .A1(n41), .A2(n731), .B1(n39), .B2(n730), .ZN(n601) );
  OAI22_X1 U1120 ( .A1(n29), .A2(n754), .B1(n28), .B2(n753), .ZN(n362) );
  OAI22_X1 U1121 ( .A1(n24), .A2(n776), .B1(n22), .B2(n775), .ZN(n643) );
  OAI22_X1 U1122 ( .A1(n5), .A2(n832), .B1(n831), .B2(n877), .ZN(n697) );
  OAI22_X1 U1123 ( .A1(n11), .A2(n817), .B1(n10), .B2(n816), .ZN(n682) );
  OAI22_X1 U1124 ( .A1(n48), .A2(n705), .B1(n46), .B2(n704), .ZN(n576) );
  INV_X1 U1125 ( .A(n338), .ZN(n339) );
  OAI22_X1 U1126 ( .A1(n48), .A2(n706), .B1(n46), .B2(n705), .ZN(n577) );
  AND2_X1 U1127 ( .A1(n1032), .A2(n558), .ZN(n669) );
  OAI22_X1 U1128 ( .A1(n5), .A2(n833), .B1(n832), .B2(n877), .ZN(n698) );
  OAI22_X1 U1129 ( .A1(n11), .A2(n818), .B1(n10), .B2(n817), .ZN(n683) );
  AOI21_X1 U1130 ( .B1(n29), .B2(n28), .A(n753), .ZN(n551) );
  OAI22_X1 U1131 ( .A1(n29), .A2(n764), .B1(n27), .B2(n763), .ZN(n632) );
  OAI22_X1 U1132 ( .A1(n18), .A2(n794), .B1(n16), .B2(n793), .ZN(n660) );
  OAI22_X1 U1133 ( .A1(n35), .A2(n749), .B1(n33), .B2(n748), .ZN(n618) );
  OAI22_X1 U1134 ( .A1(n48), .A2(n878), .B1(n718), .B2(n46), .ZN(n566) );
  OAI22_X1 U1135 ( .A1(n47), .A2(n717), .B1(n45), .B2(n716), .ZN(n588) );
  OR2_X1 U1136 ( .A1(n1032), .A2(n878), .ZN(n718) );
  OAI22_X1 U1137 ( .A1(n18), .A2(n792), .B1(n16), .B2(n791), .ZN(n658) );
  OAI22_X1 U1138 ( .A1(n6), .A2(n822), .B1(n821), .B2(n4), .ZN(n687) );
  OAI22_X1 U1139 ( .A1(n5), .A2(n830), .B1(n829), .B2(n4), .ZN(n695) );
  OAI22_X1 U1140 ( .A1(n11), .A2(n815), .B1(n10), .B2(n814), .ZN(n680) );
  OAI22_X1 U1141 ( .A1(n18), .A2(n800), .B1(n15), .B2(n799), .ZN(n666) );
  OAI22_X1 U1142 ( .A1(n6), .A2(n826), .B1(n825), .B2(n4), .ZN(n691) );
  OAI22_X1 U1143 ( .A1(n29), .A2(n766), .B1(n27), .B2(n765), .ZN(n634) );
  OAI22_X1 U1144 ( .A1(n30), .A2(n758), .B1(n28), .B2(n757), .ZN(n626) );
  OAI22_X1 U1145 ( .A1(n773), .A2(n24), .B1(n22), .B2(n772), .ZN(n640) );
  OAI22_X1 U1146 ( .A1(n35), .A2(n743), .B1(n34), .B2(n742), .ZN(n612) );
  OAI22_X1 U1147 ( .A1(n18), .A2(n801), .B1(n15), .B2(n800), .ZN(n667) );
  OAI22_X1 U1148 ( .A1(n47), .A2(n712), .B1(n45), .B2(n711), .ZN(n583) );
  INV_X1 U1149 ( .A(n557), .ZN(n654) );
  AOI21_X1 U1150 ( .B1(n18), .B2(n16), .A(n787), .ZN(n557) );
  AOI21_X1 U1151 ( .B1(n24), .B2(n22), .A(n770), .ZN(n554) );
  INV_X1 U1152 ( .A(n542), .ZN(n574) );
  AOI21_X1 U1153 ( .B1(n48), .B2(n46), .A(n702), .ZN(n542) );
  AOI21_X1 U1154 ( .B1(n6), .B2(n4), .A(n821), .ZN(n563) );
  AND2_X1 U1155 ( .A1(n956), .A2(n561), .ZN(n685) );
  INV_X1 U1156 ( .A(n10), .ZN(n561) );
  AND2_X1 U1157 ( .A1(n1032), .A2(a[0]), .ZN(product[0]) );
  OAI22_X1 U1158 ( .A1(n48), .A2(n707), .B1(n46), .B2(n706), .ZN(n578) );
  OAI22_X1 U1159 ( .A1(n42), .A2(n722), .B1(n40), .B2(n721), .ZN(n592) );
  OAI22_X1 U1160 ( .A1(n29), .A2(n759), .B1(n28), .B2(n758), .ZN(n627) );
  OAI22_X1 U1161 ( .A1(n35), .A2(n744), .B1(n33), .B2(n743), .ZN(n613) );
  OAI22_X1 U1162 ( .A1(n47), .A2(n711), .B1(n45), .B2(n710), .ZN(n582) );
  OAI22_X1 U1163 ( .A1(n29), .A2(n756), .B1(n28), .B2(n755), .ZN(n624) );
  OAI22_X1 U1164 ( .A1(n42), .A2(n726), .B1(n40), .B2(n725), .ZN(n596) );
  OAI22_X1 U1165 ( .A1(n23), .A2(n780), .B1(n21), .B2(n779), .ZN(n647) );
  OAI22_X1 U1166 ( .A1(n12), .A2(n810), .B1(n10), .B2(n809), .ZN(n675) );
  OAI22_X1 U1167 ( .A1(n35), .A2(n750), .B1(n33), .B2(n749), .ZN(n619) );
  OAI22_X1 U1168 ( .A1(n23), .A2(n779), .B1(n21), .B2(n778), .ZN(n646) );
  OAI22_X1 U1169 ( .A1(n6), .A2(n987), .B1(n823), .B2(n4), .ZN(n689) );
  OAI22_X1 U1170 ( .A1(n12), .A2(n809), .B1(n10), .B2(n808), .ZN(n674) );
  OAI22_X1 U1171 ( .A1(n30), .A2(n760), .B1(n28), .B2(n759), .ZN(n628) );
  OAI22_X1 U1172 ( .A1(n775), .A2(n24), .B1(n22), .B2(n774), .ZN(n642) );
  OAI22_X1 U1173 ( .A1(n41), .A2(n730), .B1(n39), .B2(n729), .ZN(n600) );
  OAI22_X1 U1174 ( .A1(n24), .A2(n774), .B1(n22), .B2(n773), .ZN(n641) );
  OAI22_X1 U1175 ( .A1(n18), .A2(n789), .B1(n16), .B2(n788), .ZN(n655) );
  OAI22_X1 U1176 ( .A1(n41), .A2(n729), .B1(n39), .B2(n728), .ZN(n599) );
  OAI22_X1 U1177 ( .A1(n35), .A2(n740), .B1(n34), .B2(n739), .ZN(n609) );
  OAI22_X1 U1178 ( .A1(n42), .A2(n725), .B1(n40), .B2(n724), .ZN(n595) );
  OAI22_X1 U1179 ( .A1(n17), .A2(n791), .B1(n16), .B2(n790), .ZN(n657) );
  OAI22_X1 U1180 ( .A1(n12), .A2(n806), .B1(n10), .B2(n805), .ZN(n671) );
  OAI22_X1 U1181 ( .A1(n36), .A2(n746), .B1(n33), .B2(n745), .ZN(n615) );
  OAI22_X1 U1182 ( .A1(n23), .A2(n781), .B1(n21), .B2(n780), .ZN(n648) );
  OAI22_X1 U1183 ( .A1(n12), .A2(n811), .B1(n10), .B2(n810), .ZN(n676) );
  OAI22_X1 U1184 ( .A1(n35), .A2(n741), .B1(n34), .B2(n740), .ZN(n610) );
  INV_X1 U1185 ( .A(n380), .ZN(n381) );
  OAI22_X1 U1186 ( .A1(n35), .A2(n742), .B1(n34), .B2(n741), .ZN(n611) );
  OAI22_X1 U1187 ( .A1(n24), .A2(n772), .B1(n22), .B2(n771), .ZN(n639) );
  OAI22_X1 U1188 ( .A1(n41), .A2(n727), .B1(n39), .B2(n726), .ZN(n597) );
  OAI22_X1 U1189 ( .A1(n11), .A2(n813), .B1(n10), .B2(n812), .ZN(n678) );
  OAI22_X1 U1190 ( .A1(n18), .A2(n798), .B1(n15), .B2(n797), .ZN(n664) );
  OAI22_X1 U1191 ( .A1(n23), .A2(n783), .B1(n21), .B2(n782), .ZN(n650) );
  OAI22_X1 U1192 ( .A1(n18), .A2(n797), .B1(n15), .B2(n796), .ZN(n663) );
  OAI22_X1 U1193 ( .A1(n29), .A2(n767), .B1(n27), .B2(n766), .ZN(n635) );
  OAI22_X1 U1194 ( .A1(n11), .A2(n812), .B1(n10), .B2(n811), .ZN(n677) );
  OAI22_X1 U1195 ( .A1(n23), .A2(n778), .B1(n21), .B2(n777), .ZN(n645) );
  OAI22_X1 U1196 ( .A1(n18), .A2(n793), .B1(n16), .B2(n792), .ZN(n659) );
  OAI22_X1 U1197 ( .A1(n47), .A2(n710), .B1(n45), .B2(n709), .ZN(n581) );
  OAI22_X1 U1198 ( .A1(n29), .A2(n755), .B1(n28), .B2(n754), .ZN(n623) );
  INV_X1 U1199 ( .A(n554), .ZN(n638) );
  OAI22_X1 U1200 ( .A1(n42), .A2(n721), .B1(n40), .B2(n720), .ZN(n591) );
  INV_X1 U1201 ( .A(n548), .ZN(n606) );
  AOI21_X1 U1202 ( .B1(n35), .B2(n34), .A(n736), .ZN(n548) );
  OAI22_X1 U1203 ( .A1(n23), .A2(n784), .B1(n21), .B2(n783), .ZN(n651) );
  OAI22_X1 U1204 ( .A1(n11), .A2(n814), .B1(n10), .B2(n813), .ZN(n679) );
  OAI22_X1 U1205 ( .A1(n6), .A2(n828), .B1(n827), .B2(n4), .ZN(n693) );
  OAI22_X1 U1206 ( .A1(n12), .A2(n807), .B1(n10), .B2(n806), .ZN(n672) );
  OAI22_X1 U1207 ( .A1(n6), .A2(n827), .B1(n826), .B2(n4), .ZN(n692) );
  OAI22_X1 U1208 ( .A1(n23), .A2(n782), .B1(n21), .B2(n781), .ZN(n649) );
  AND2_X1 U1209 ( .A1(n956), .A2(n549), .ZN(n621) );
  OAI22_X1 U1210 ( .A1(n6), .A2(n823), .B1(n822), .B2(n4), .ZN(n688) );
  AND2_X1 U1211 ( .A1(n1032), .A2(n543), .ZN(n589) );
  OAI22_X1 U1212 ( .A1(n36), .A2(n748), .B1(n33), .B2(n747), .ZN(n617) );
  OAI22_X1 U1213 ( .A1(n715), .A2(n47), .B1(n45), .B2(n714), .ZN(n586) );
  OAI22_X1 U1214 ( .A1(n17), .A2(n790), .B1(n16), .B2(n789), .ZN(n656) );
  OAI22_X1 U1215 ( .A1(n36), .A2(n993), .B1(n33), .B2(n744), .ZN(n614) );
  OAI22_X1 U1216 ( .A1(n5), .A2(n831), .B1(n830), .B2(n4), .ZN(n696) );
  AND2_X1 U1217 ( .A1(n1032), .A2(n555), .ZN(n653) );
  OAI22_X1 U1218 ( .A1(n11), .A2(n816), .B1(n10), .B2(n815), .ZN(n681) );
  OAI22_X1 U1219 ( .A1(n29), .A2(n763), .B1(n27), .B2(n762), .ZN(n631) );
  OAI22_X1 U1220 ( .A1(n12), .A2(n808), .B1(n10), .B2(n807), .ZN(n673) );
  OAI22_X1 U1221 ( .A1(n41), .A2(n733), .B1(n39), .B2(n732), .ZN(n603) );
  OAI22_X1 U1222 ( .A1(n47), .A2(n714), .B1(n45), .B2(n713), .ZN(n585) );
  INV_X1 U1223 ( .A(n560), .ZN(n670) );
  AOI21_X1 U1224 ( .B1(n12), .B2(n10), .A(n804), .ZN(n560) );
  OAI22_X1 U1225 ( .A1(n48), .A2(n708), .B1(n46), .B2(n707), .ZN(n579) );
  OAI22_X1 U1226 ( .A1(n42), .A2(n723), .B1(n40), .B2(n722), .ZN(n593) );
  INV_X1 U1227 ( .A(n551), .ZN(n622) );
  OAI22_X1 U1228 ( .A1(n24), .A2(n777), .B1(n22), .B2(n776), .ZN(n644) );
  OAI22_X1 U1229 ( .A1(n35), .A2(n747), .B1(n33), .B2(n746), .ZN(n616) );
  OAI22_X1 U1230 ( .A1(n41), .A2(n732), .B1(n39), .B2(n731), .ZN(n602) );
  OAI22_X1 U1231 ( .A1(n29), .A2(n757), .B1(n28), .B2(n756), .ZN(n625) );
  OAI22_X1 U1232 ( .A1(n18), .A2(n795), .B1(n15), .B2(n794), .ZN(n661) );
  OAI22_X1 U1233 ( .A1(n35), .A2(n738), .B1(n34), .B2(n737), .ZN(n607) );
  OAI22_X1 U1234 ( .A1(n5), .A2(n829), .B1(n828), .B2(n877), .ZN(n694) );
  AND2_X1 U1235 ( .A1(n1032), .A2(n552), .ZN(n637) );
  OAI22_X1 U1236 ( .A1(n18), .A2(n799), .B1(n15), .B2(n798), .ZN(n665) );
  OAI22_X1 U1237 ( .A1(n35), .A2(n739), .B1(n34), .B2(n738), .ZN(n608) );
  OAI22_X1 U1238 ( .A1(n48), .A2(n709), .B1(n46), .B2(n708), .ZN(n580) );
  OAI22_X1 U1239 ( .A1(n42), .A2(n724), .B1(n40), .B2(n723), .ZN(n594) );
  NAND2_X1 U1240 ( .A1(n701), .A2(n573), .ZN(n301) );
  OAI22_X1 U1241 ( .A1(n36), .A2(n880), .B1(n752), .B2(n34), .ZN(n568) );
  OAI22_X1 U1242 ( .A1(n751), .A2(n36), .B1(n33), .B2(n750), .ZN(n620) );
  OR2_X1 U1243 ( .A1(n1033), .A2(n880), .ZN(n752) );
  NAND2_X1 U1244 ( .A1(n539), .A2(n540), .ZN(n291) );
  OAI22_X1 U1245 ( .A1(n42), .A2(n879), .B1(n735), .B2(n40), .ZN(n567) );
  OAI22_X1 U1246 ( .A1(n734), .A2(n41), .B1(n39), .B2(n733), .ZN(n604) );
  OR2_X1 U1247 ( .A1(n1032), .A2(n879), .ZN(n735) );
  OAI22_X1 U1248 ( .A1(n47), .A2(n713), .B1(n45), .B2(n712), .ZN(n584) );
  OAI22_X1 U1249 ( .A1(n41), .A2(n728), .B1(n39), .B2(n727), .ZN(n598) );
  INV_X1 U1250 ( .A(n402), .ZN(n403) );
  OAI22_X1 U1251 ( .A1(n6), .A2(n825), .B1(n824), .B2(n4), .ZN(n690) );
  OAI22_X1 U1252 ( .A1(n30), .A2(n765), .B1(n27), .B2(n764), .ZN(n633) );
  AND2_X1 U1253 ( .A1(n956), .A2(n546), .ZN(n605) );
  OR2_X1 U1254 ( .A1(n956), .A2(n883), .ZN(n803) );
  OR2_X1 U1255 ( .A1(n1032), .A2(n881), .ZN(n769) );
  OR2_X1 U1256 ( .A1(n956), .A2(n882), .ZN(n786) );
  INV_X1 U1257 ( .A(n15), .ZN(n558) );
  INV_X1 U1258 ( .A(n27), .ZN(n552) );
  OAI22_X1 U1259 ( .A1(n47), .A2(n716), .B1(n45), .B2(n715), .ZN(n587) );
  OAI22_X1 U1260 ( .A1(n30), .A2(n761), .B1(n27), .B2(n760), .ZN(n629) );
  INV_X1 U1261 ( .A(n563), .ZN(n686) );
  OAI22_X1 U1262 ( .A1(n48), .A2(n704), .B1(n46), .B2(n703), .ZN(n575) );
  INV_X1 U1263 ( .A(n545), .ZN(n590) );
  AOI21_X1 U1264 ( .B1(n42), .B2(n40), .A(n719), .ZN(n545) );
  INV_X1 U1265 ( .A(n21), .ZN(n555) );
  INV_X1 U1266 ( .A(n39), .ZN(n546) );
  INV_X1 U1267 ( .A(n33), .ZN(n549) );
  INV_X1 U1268 ( .A(n45), .ZN(n543) );
  BUF_X1 U1269 ( .A(n877), .Z(n4) );
  OAI22_X1 U1270 ( .A1(n11), .A2(n819), .B1(n10), .B2(n818), .ZN(n684) );
  OAI22_X1 U1271 ( .A1(n5), .A2(n834), .B1(n833), .B2(n4), .ZN(n699) );
  OAI22_X1 U1272 ( .A1(n6), .A2(n885), .B1(n837), .B2(n4), .ZN(n573) );
  OR2_X1 U1273 ( .A1(n956), .A2(n885), .ZN(n837) );
  INV_X1 U1274 ( .A(n1), .ZN(n885) );
  OAI22_X1 U1275 ( .A1(n12), .A2(n884), .B1(n820), .B2(n10), .ZN(n572) );
  OR2_X1 U1276 ( .A1(n956), .A2(n884), .ZN(n820) );
  OAI22_X1 U1277 ( .A1(n5), .A2(n836), .B1(n835), .B2(n4), .ZN(n701) );
  OAI22_X1 U1278 ( .A1(n29), .A2(n768), .B1(n27), .B2(n767), .ZN(n636) );
  OAI22_X1 U1279 ( .A1(n29), .A2(n881), .B1(n769), .B2(n28), .ZN(n569) );
  XNOR2_X1 U1280 ( .A(n989), .B(n851), .ZN(n732) );
  XNOR2_X1 U1281 ( .A(n989), .B(n850), .ZN(n731) );
  XNOR2_X1 U1282 ( .A(n989), .B(n1009), .ZN(n723) );
  OAI22_X1 U1283 ( .A1(n23), .A2(n785), .B1(n21), .B2(n784), .ZN(n652) );
  OAI22_X1 U1284 ( .A1(n24), .A2(n882), .B1(n786), .B2(n22), .ZN(n570) );
  XNOR2_X1 U1285 ( .A(n989), .B(n838), .ZN(n719) );
  XNOR2_X1 U1286 ( .A(n848), .B(n37), .ZN(n729) );
  XNOR2_X1 U1287 ( .A(n37), .B(n847), .ZN(n728) );
  XNOR2_X1 U1288 ( .A(n37), .B(n852), .ZN(n733) );
  XNOR2_X1 U1289 ( .A(n989), .B(n846), .ZN(n727) );
  XNOR2_X1 U1290 ( .A(n989), .B(n849), .ZN(n730) );
  XNOR2_X1 U1291 ( .A(n989), .B(n1005), .ZN(n725) );
  XNOR2_X1 U1292 ( .A(n989), .B(n843), .ZN(n724) );
  XNOR2_X1 U1293 ( .A(n989), .B(n845), .ZN(n726) );
  XNOR2_X1 U1294 ( .A(n989), .B(n840), .ZN(n721) );
  XNOR2_X1 U1295 ( .A(n989), .B(n1030), .ZN(n722) );
  XNOR2_X1 U1296 ( .A(n989), .B(n995), .ZN(n720) );
  OAI22_X1 U1297 ( .A1(n17), .A2(n802), .B1(n15), .B2(n801), .ZN(n668) );
  OAI22_X1 U1298 ( .A1(n17), .A2(n883), .B1(n803), .B2(n16), .ZN(n571) );
  BUF_X1 U1299 ( .A(n871), .Z(n39) );
  BUF_X1 U1300 ( .A(n872), .Z(n33) );
  BUF_X1 U1301 ( .A(n871), .Z(n40) );
  BUF_X1 U1302 ( .A(n870), .Z(n46) );
  BUF_X1 U1303 ( .A(n862), .Z(n48) );
  XNOR2_X1 U1304 ( .A(n37), .B(n1032), .ZN(n734) );
  BUF_X1 U1305 ( .A(n868), .Z(n11) );
  INV_X1 U1306 ( .A(n25), .ZN(n881) );
  INV_X1 U1307 ( .A(n13), .ZN(n883) );
  INV_X1 U1308 ( .A(n19), .ZN(n882) );
  INV_X1 U1309 ( .A(n43), .ZN(n878) );
  INV_X1 U1310 ( .A(n31), .ZN(n880) );
  XNOR2_X1 U1311 ( .A(a[12]), .B(a[11]), .ZN(n871) );
  XNOR2_X1 U1312 ( .A(a[10]), .B(a[9]), .ZN(n872) );
  XNOR2_X1 U1313 ( .A(a[14]), .B(a[13]), .ZN(n870) );
  BUF_X2 U1314 ( .A(a[11]), .Z(n31) );
  NAND2_X1 U1315 ( .A1(n860), .A2(n876), .ZN(n868) );
  NAND2_X1 U1316 ( .A1(n855), .A2(n871), .ZN(n863) );
  XNOR2_X1 U1317 ( .A(a[6]), .B(a[5]), .ZN(n874) );
  OAI22_X1 U1318 ( .A1(n35), .A2(n737), .B1(n34), .B2(n736), .ZN(n348) );
  INV_X1 U1319 ( .A(n348), .ZN(n349) );
  INV_X1 U1320 ( .A(n7), .ZN(n884) );
  XNOR2_X1 U1321 ( .A(n7), .B(n844), .ZN(n810) );
  XNOR2_X1 U1322 ( .A(n7), .B(n840), .ZN(n806) );
  XNOR2_X1 U1323 ( .A(n7), .B(n1029), .ZN(n807) );
  XNOR2_X1 U1324 ( .A(n7), .B(n843), .ZN(n809) );
  XNOR2_X1 U1325 ( .A(n7), .B(n1008), .ZN(n808) );
  XNOR2_X1 U1326 ( .A(n7), .B(n1032), .ZN(n819) );
  XNOR2_X1 U1327 ( .A(n7), .B(n847), .ZN(n813) );
  XNOR2_X1 U1328 ( .A(n7), .B(n849), .ZN(n815) );
  XNOR2_X1 U1329 ( .A(n7), .B(n848), .ZN(n814) );
  XNOR2_X1 U1330 ( .A(n7), .B(n846), .ZN(n812) );
  XNOR2_X1 U1331 ( .A(n7), .B(n845), .ZN(n811) );
  XNOR2_X1 U1332 ( .A(n7), .B(n852), .ZN(n818) );
  XNOR2_X1 U1333 ( .A(n7), .B(n850), .ZN(n816) );
  XNOR2_X1 U1334 ( .A(n7), .B(n839), .ZN(n805) );
  XNOR2_X1 U1335 ( .A(n7), .B(n851), .ZN(n817) );
  XNOR2_X1 U1336 ( .A(n7), .B(n838), .ZN(n804) );
  NAND2_X1 U1337 ( .A1(n856), .A2(n872), .ZN(n864) );
  XNOR2_X1 U1338 ( .A(a[8]), .B(a[7]), .ZN(n873) );
  NOR2_X1 U1339 ( .A1(n144), .A2(n137), .ZN(n135) );
  OAI21_X1 U1340 ( .B1(n145), .B2(n137), .A(n138), .ZN(n136) );
  INV_X1 U1341 ( .A(n252), .ZN(n250) );
  NOR2_X1 U1342 ( .A1(n492), .A2(n483), .ZN(n252) );
  NAND2_X1 U1343 ( .A1(n417), .A2(n430), .ZN(n219) );
  NAND2_X1 U1344 ( .A1(n861), .A2(n877), .ZN(n869) );
  AOI21_X1 U1345 ( .B1(n974), .B2(n297), .A(n294), .ZN(n292) );
  INV_X1 U1346 ( .A(n296), .ZN(n294) );
  NAND2_X1 U1347 ( .A1(n974), .A2(n296), .ZN(n81) );
  OAI21_X1 U1348 ( .B1(n224), .B2(n1000), .A(n985), .ZN(n215) );
  INV_X1 U1349 ( .A(n990), .ZN(n224) );
  INV_X1 U1350 ( .A(n362), .ZN(n363) );
  INV_X1 U1351 ( .A(a[0]), .ZN(n877) );
  INV_X1 U1352 ( .A(n282), .ZN(n326) );
  NOR2_X1 U1353 ( .A1(n531), .A2(n534), .ZN(n282) );
  OAI21_X1 U1354 ( .B1(n290), .B2(n292), .A(n291), .ZN(n289) );
  NAND2_X1 U1355 ( .A1(n541), .A2(n572), .ZN(n296) );
  NAND2_X1 U1356 ( .A1(n858), .A2(n874), .ZN(n866) );
  NAND2_X1 U1357 ( .A1(n365), .A2(n372), .ZN(n182) );
  INV_X1 U1358 ( .A(n37), .ZN(n879) );
  NAND2_X1 U1359 ( .A1(n459), .A2(n470), .ZN(n239) );
  OAI21_X1 U1360 ( .B1(n227), .B2(n233), .A(n228), .ZN(n226) );
  XNOR2_X1 U1361 ( .A(n19), .B(n1032), .ZN(n785) );
  XNOR2_X1 U1362 ( .A(n19), .B(n844), .ZN(n776) );
  XNOR2_X1 U1363 ( .A(n19), .B(n845), .ZN(n777) );
  XNOR2_X1 U1364 ( .A(n19), .B(n852), .ZN(n784) );
  XNOR2_X1 U1365 ( .A(n19), .B(n848), .ZN(n780) );
  XNOR2_X1 U1366 ( .A(n19), .B(n846), .ZN(n778) );
  XNOR2_X1 U1367 ( .A(n19), .B(n843), .ZN(n775) );
  XNOR2_X1 U1368 ( .A(n19), .B(n847), .ZN(n779) );
  XNOR2_X1 U1369 ( .A(n19), .B(n851), .ZN(n783) );
  XNOR2_X1 U1370 ( .A(n19), .B(n842), .ZN(n774) );
  XNOR2_X1 U1371 ( .A(n19), .B(n839), .ZN(n771) );
  XNOR2_X1 U1372 ( .A(n19), .B(n850), .ZN(n782) );
  XNOR2_X1 U1373 ( .A(n19), .B(n849), .ZN(n781) );
  XNOR2_X1 U1374 ( .A(n19), .B(n838), .ZN(n770) );
  XNOR2_X1 U1375 ( .A(n19), .B(n1030), .ZN(n773) );
  XNOR2_X1 U1376 ( .A(n19), .B(n840), .ZN(n772) );
  AOI21_X1 U1377 ( .B1(n209), .B2(n226), .A(n210), .ZN(n208) );
  XNOR2_X1 U1378 ( .A(n43), .B(n840), .ZN(n704) );
  XNOR2_X1 U1379 ( .A(n43), .B(n1029), .ZN(n705) );
  XNOR2_X1 U1380 ( .A(n43), .B(n995), .ZN(n703) );
  XNOR2_X1 U1381 ( .A(n43), .B(n838), .ZN(n702) );
  XNOR2_X1 U1382 ( .A(n43), .B(n843), .ZN(n707) );
  XNOR2_X1 U1383 ( .A(n43), .B(n1008), .ZN(n706) );
  XNOR2_X1 U1384 ( .A(n43), .B(n1005), .ZN(n708) );
  XNOR2_X1 U1385 ( .A(n43), .B(n847), .ZN(n711) );
  XNOR2_X1 U1386 ( .A(n43), .B(n846), .ZN(n710) );
  XNOR2_X1 U1387 ( .A(n43), .B(n851), .ZN(n715) );
  XNOR2_X1 U1388 ( .A(n43), .B(n956), .ZN(n717) );
  XNOR2_X1 U1389 ( .A(n43), .B(n845), .ZN(n709) );
  XNOR2_X1 U1390 ( .A(n43), .B(n852), .ZN(n716) );
  XNOR2_X1 U1391 ( .A(n43), .B(n850), .ZN(n714) );
  XNOR2_X1 U1392 ( .A(n43), .B(n849), .ZN(n713) );
  XNOR2_X1 U1393 ( .A(n43), .B(n848), .ZN(n712) );
  XNOR2_X1 U1394 ( .A(n25), .B(n1029), .ZN(n756) );
  XNOR2_X1 U1395 ( .A(n25), .B(n956), .ZN(n768) );
  XNOR2_X1 U1396 ( .A(n25), .B(n840), .ZN(n755) );
  XNOR2_X1 U1397 ( .A(n25), .B(n845), .ZN(n760) );
  XNOR2_X1 U1398 ( .A(n25), .B(n847), .ZN(n762) );
  XNOR2_X1 U1399 ( .A(n25), .B(n849), .ZN(n764) );
  XNOR2_X1 U1400 ( .A(n25), .B(n848), .ZN(n763) );
  XNOR2_X1 U1401 ( .A(n25), .B(n852), .ZN(n767) );
  XNOR2_X1 U1402 ( .A(n25), .B(n844), .ZN(n759) );
  XNOR2_X1 U1403 ( .A(n25), .B(n846), .ZN(n761) );
  XNOR2_X1 U1404 ( .A(n25), .B(n843), .ZN(n758) );
  XNOR2_X1 U1405 ( .A(n25), .B(n851), .ZN(n766) );
  XNOR2_X1 U1406 ( .A(n25), .B(n850), .ZN(n765) );
  XNOR2_X1 U1407 ( .A(n25), .B(n1008), .ZN(n757) );
  XNOR2_X1 U1408 ( .A(n25), .B(n839), .ZN(n754) );
  XNOR2_X1 U1409 ( .A(n25), .B(n838), .ZN(n753) );
  XNOR2_X1 U1410 ( .A(n81), .B(n297), .ZN(product[3]) );
  XOR2_X1 U1411 ( .A(n82), .B(n301), .Z(product[2]) );
  OAI21_X1 U1412 ( .B1(n298), .B2(n301), .A(n299), .ZN(n297) );
  XNOR2_X1 U1413 ( .A(n1), .B(n845), .ZN(n828) );
  XNOR2_X1 U1414 ( .A(n1), .B(n956), .ZN(n836) );
  XNOR2_X1 U1415 ( .A(n1), .B(n846), .ZN(n829) );
  XNOR2_X1 U1416 ( .A(n1), .B(n1029), .ZN(n824) );
  XNOR2_X1 U1417 ( .A(n1), .B(n842), .ZN(n825) );
  XNOR2_X1 U1418 ( .A(n1), .B(n840), .ZN(n823) );
  XNOR2_X1 U1419 ( .A(n1), .B(n839), .ZN(n822) );
  XNOR2_X1 U1420 ( .A(n1), .B(n849), .ZN(n832) );
  XNOR2_X1 U1421 ( .A(n1), .B(n847), .ZN(n830) );
  XNOR2_X1 U1422 ( .A(n1), .B(n844), .ZN(n827) );
  XNOR2_X1 U1423 ( .A(n1), .B(n848), .ZN(n831) );
  XNOR2_X1 U1424 ( .A(n1), .B(n843), .ZN(n826) );
  XNOR2_X1 U1425 ( .A(n1), .B(n838), .ZN(n821) );
  XNOR2_X1 U1426 ( .A(n1), .B(n850), .ZN(n833) );
  XNOR2_X1 U1427 ( .A(n1), .B(n851), .ZN(n834) );
  XNOR2_X1 U1428 ( .A(n1), .B(n852), .ZN(n835) );
  XNOR2_X1 U1429 ( .A(a[2]), .B(a[1]), .ZN(n876) );
  OAI21_X1 U1430 ( .B1(n282), .B2(n284), .A(n283), .ZN(n281) );
  XOR2_X1 U1431 ( .A(n262), .B(n73), .Z(product[11]) );
  AOI21_X1 U1432 ( .B1(n267), .B2(n968), .A(n264), .ZN(n262) );
  OAI21_X1 U1433 ( .B1(n254), .B2(n241), .A(n994), .ZN(n240) );
  AOI21_X1 U1434 ( .B1(n1027), .B2(n251), .A(n244), .ZN(n242) );
  XNOR2_X1 U1435 ( .A(n1001), .B(n840), .ZN(n738) );
  XNOR2_X1 U1436 ( .A(n1001), .B(n843), .ZN(n741) );
  XNOR2_X1 U1437 ( .A(n1001), .B(n848), .ZN(n746) );
  XNOR2_X1 U1438 ( .A(n1001), .B(n842), .ZN(n740) );
  XNOR2_X1 U1439 ( .A(n1001), .B(n1030), .ZN(n739) );
  XNOR2_X1 U1440 ( .A(n31), .B(n847), .ZN(n745) );
  XNOR2_X1 U1441 ( .A(n31), .B(n846), .ZN(n744) );
  XNOR2_X1 U1442 ( .A(n1001), .B(n851), .ZN(n749) );
  XNOR2_X1 U1443 ( .A(n1001), .B(n1033), .ZN(n751) );
  XNOR2_X1 U1444 ( .A(n1001), .B(n850), .ZN(n748) );
  XNOR2_X1 U1445 ( .A(n31), .B(n849), .ZN(n747) );
  XNOR2_X1 U1446 ( .A(n31), .B(n852), .ZN(n750) );
  XNOR2_X1 U1447 ( .A(n1001), .B(n845), .ZN(n743) );
  XNOR2_X1 U1448 ( .A(n31), .B(n1005), .ZN(n742) );
  XNOR2_X1 U1449 ( .A(n1001), .B(n995), .ZN(n737) );
  XNOR2_X1 U1450 ( .A(n1001), .B(n838), .ZN(n736) );
  AOI21_X1 U1451 ( .B1(n970), .B2(n151), .A(n152), .ZN(n150) );
  NAND2_X1 U1452 ( .A1(n383), .A2(n392), .ZN(n200) );
  NAND2_X1 U1453 ( .A1(n857), .A2(n873), .ZN(n865) );
  OAI22_X1 U1454 ( .A1(n30), .A2(n762), .B1(n27), .B2(n761), .ZN(n630) );
  INV_X1 U1455 ( .A(n246), .ZN(n244) );
  NAND2_X1 U1456 ( .A1(n1027), .A2(n246), .ZN(n71) );
  NAND2_X1 U1457 ( .A1(n483), .A2(n492), .ZN(n253) );
  INV_X1 U1458 ( .A(n253), .ZN(n251) );
  NAND2_X1 U1459 ( .A1(n250), .A2(n253), .ZN(n72) );
  NOR2_X1 U1460 ( .A1(n1031), .A2(n87), .ZN(n85) );
  NOR2_X1 U1461 ( .A1(n1031), .A2(n96), .ZN(n94) );
  NOR2_X1 U1462 ( .A1(n1031), .A2(n133), .ZN(n131) );
  NOR2_X1 U1463 ( .A1(n1031), .A2(n144), .ZN(n140) );
  NOR2_X1 U1464 ( .A1(n1031), .A2(n109), .ZN(n107) );
  NOR2_X1 U1465 ( .A1(n1031), .A2(n124), .ZN(n118) );
  AOI21_X1 U1466 ( .B1(n234), .B2(n230), .A(n231), .ZN(n229) );
  XNOR2_X1 U1467 ( .A(n234), .B(n69), .ZN(product[15]) );
  AOI21_X1 U1468 ( .B1(n214), .B2(n234), .A(n215), .ZN(n213) );
  AOI21_X1 U1469 ( .B1(n234), .B2(n221), .A(n990), .ZN(n220) );
  INV_X1 U1470 ( .A(n997), .ZN(n234) );
  XNOR2_X1 U1471 ( .A(n79), .B(n289), .ZN(product[5]) );
  AOI21_X1 U1472 ( .B1(n255), .B2(n236), .A(n237), .ZN(n235) );
  AOI21_X1 U1473 ( .B1(n289), .B2(n977), .A(n286), .ZN(n284) );
  AOI21_X1 U1474 ( .B1(n155), .B2(n180), .A(n156), .ZN(n154) );
  NAND2_X1 U1475 ( .A1(n155), .A2(n992), .ZN(n153) );
  INV_X1 U1476 ( .A(n1000), .ZN(n315) );
  NOR2_X1 U1477 ( .A1(n417), .A2(n430), .ZN(n218) );
  NAND2_X1 U1478 ( .A1(n209), .A2(n225), .ZN(n207) );
  OAI21_X1 U1479 ( .B1(n984), .B2(n87), .A(n88), .ZN(n86) );
  OAI21_X1 U1480 ( .B1(n984), .B2(n96), .A(n97), .ZN(n95) );
  OAI21_X1 U1481 ( .B1(n150), .B2(n144), .A(n145), .ZN(n141) );
  OAI21_X1 U1482 ( .B1(n984), .B2(n109), .A(n110), .ZN(n108) );
  OAI21_X1 U1483 ( .B1(n983), .B2(n124), .A(n125), .ZN(n119) );
  OAI21_X1 U1484 ( .B1(n150), .B2(n133), .A(n134), .ZN(n132) );
  OAI21_X1 U1485 ( .B1(n153), .B2(n191), .A(n154), .ZN(n152) );
  NAND2_X1 U1486 ( .A1(n859), .A2(n875), .ZN(n867) );
  OAI21_X1 U1487 ( .B1(n207), .B2(n235), .A(n208), .ZN(n206) );
  INV_X1 U1488 ( .A(n168), .ZN(n167) );
  NOR2_X1 U1489 ( .A1(n168), .A2(n157), .ZN(n155) );
  NAND2_X1 U1490 ( .A1(n854), .A2(n870), .ZN(n862) );
  NOR2_X1 U1491 ( .A1(n227), .A2(n232), .ZN(n225) );
  AOI21_X1 U1492 ( .B1(n273), .B2(n978), .A(n270), .ZN(n268) );
  NOR2_X1 U1493 ( .A1(n991), .A2(n218), .ZN(n209) );
  OAI21_X1 U1494 ( .B1(n211), .B2(n219), .A(n212), .ZN(n210) );
  OAI21_X1 U1495 ( .B1(n157), .B2(n169), .A(n158), .ZN(n156) );
  NAND2_X1 U1496 ( .A1(n351), .A2(n356), .ZN(n158) );
  XNOR2_X1 U1497 ( .A(n273), .B(n75), .ZN(product[9]) );
  XNOR2_X1 U1498 ( .A(n13), .B(n845), .ZN(n794) );
  XNOR2_X1 U1499 ( .A(n13), .B(n851), .ZN(n800) );
  XNOR2_X1 U1500 ( .A(n13), .B(n1005), .ZN(n793) );
  XNOR2_X1 U1501 ( .A(n13), .B(n843), .ZN(n792) );
  XNOR2_X1 U1502 ( .A(n13), .B(n848), .ZN(n797) );
  XNOR2_X1 U1503 ( .A(n13), .B(n1028), .ZN(n790) );
  XNOR2_X1 U1504 ( .A(n13), .B(n1009), .ZN(n791) );
  XNOR2_X1 U1505 ( .A(n13), .B(n840), .ZN(n789) );
  XNOR2_X1 U1506 ( .A(n13), .B(n850), .ZN(n799) );
  XNOR2_X1 U1507 ( .A(n13), .B(n849), .ZN(n798) );
  XNOR2_X1 U1508 ( .A(n13), .B(n847), .ZN(n796) );
  XNOR2_X1 U1509 ( .A(n13), .B(n846), .ZN(n795) );
  XNOR2_X1 U1510 ( .A(n13), .B(n1033), .ZN(n802) );
  XNOR2_X1 U1511 ( .A(n13), .B(n839), .ZN(n788) );
  XNOR2_X1 U1512 ( .A(n13), .B(n852), .ZN(n801) );
  XNOR2_X1 U1513 ( .A(n13), .B(n838), .ZN(n787) );
  XOR2_X1 U1514 ( .A(a[14]), .B(a[15]), .Z(n854) );
  XOR2_X1 U1515 ( .A(a[6]), .B(a[7]), .Z(n858) );
  NOR2_X1 U1516 ( .A1(n241), .A2(n238), .ZN(n236) );
  OAI21_X1 U1517 ( .B1(n242), .B2(n238), .A(n239), .ZN(n237) );
  XOR2_X1 U1518 ( .A(a[12]), .B(a[13]), .Z(n855) );
  XOR2_X1 U1519 ( .A(a[10]), .B(a[11]), .Z(n856) );
  XOR2_X1 U1520 ( .A(n80), .B(n292), .Z(product[4]) );
  XOR2_X1 U1521 ( .A(a[8]), .B(a[9]), .Z(n857) );
  AOI21_X1 U1522 ( .B1(n1026), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U1523 ( .B1(n1026), .B2(n94), .A(n95), .ZN(n93) );
  AOI21_X1 U1524 ( .B1(n1026), .B2(n118), .A(n119), .ZN(n117) );
  AOI21_X1 U1525 ( .B1(n1026), .B2(n107), .A(n108), .ZN(n106) );
  AOI21_X1 U1526 ( .B1(n1026), .B2(n160), .A(n161), .ZN(n159) );
  AOI21_X1 U1527 ( .B1(n1026), .B2(n140), .A(n141), .ZN(n139) );
  AOI21_X1 U1528 ( .B1(n1026), .B2(n131), .A(n132), .ZN(n130) );
  AOI21_X1 U1529 ( .B1(n51), .B2(n193), .A(n970), .ZN(n192) );
  XNOR2_X1 U1530 ( .A(n1026), .B(n65), .ZN(product[19]) );
  AOI21_X1 U1531 ( .B1(n51), .B2(n313), .A(n203), .ZN(n201) );
  AOI21_X1 U1532 ( .B1(n51), .B2(n184), .A(n185), .ZN(n183) );
  AOI21_X1 U1533 ( .B1(n51), .B2(n171), .A(n172), .ZN(n170) );
  XOR2_X1 U1534 ( .A(a[0]), .B(a[1]), .Z(n861) );
  NOR2_X1 U1535 ( .A1(n204), .A2(n199), .ZN(n197) );
  NAND2_X1 U1536 ( .A1(n471), .A2(n482), .ZN(n246) );
  XNOR2_X1 U1537 ( .A(a[4]), .B(a[3]), .ZN(n875) );
  XOR2_X1 U1538 ( .A(a[2]), .B(a[3]), .Z(n860) );
  AOI21_X1 U1539 ( .B1(n51), .B2(n147), .A(n148), .ZN(n146) );
  XOR2_X1 U1540 ( .A(n953), .B(n76), .Z(product[8]) );
  XNOR2_X1 U1541 ( .A(n986), .B(n77), .ZN(product[7]) );
  AOI21_X1 U1542 ( .B1(n281), .B2(n979), .A(n278), .ZN(n276) );
  XOR2_X1 U1543 ( .A(a[4]), .B(a[5]), .Z(n859) );
  XOR2_X1 U1544 ( .A(n78), .B(n1004), .Z(product[6]) );
endmodule


module datapath_DW_mult_tc_9 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n15, n16, n17, n18,
         n19, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34, n35,
         n36, n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n51, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n84, n85, n86, n87, n88, n90, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n103, n105, n106, n107, n108, n109, n110,
         n114, n116, n117, n118, n119, n122, n123, n124, n125, n127, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n177, n182, n183, n184, n185, n186, n188, n189, n190, n191,
         n192, n194, n195, n196, n197, n198, n199, n200, n201, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n217, n218, n219, n220, n221, n224, n225, n226, n227, n228, n229,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n247, n249, n251, n252, n253, n254, n255, n256, n257, n259,
         n261, n262, n264, n266, n267, n268, n270, n272, n273, n274, n275,
         n276, n278, n280, n281, n282, n283, n284, n286, n288, n289, n290,
         n291, n292, n294, n296, n297, n298, n299, n301, n306, n308, n312,
         n313, n316, n317, n318, n320, n324, n326, n328, n330, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n545, n546, n548, n549, n551, n552, n554, n555, n557, n558, n560,
         n561, n563, n564, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1056, n1057, n1058;
  assign product[31] = n84;

  FA_X1 U364 ( .A(n575), .B(n338), .CI(n590), .CO(n334), .S(n335) );
  FA_X1 U365 ( .A(n339), .B(n576), .CI(n342), .CO(n336), .S(n337) );
  FA_X1 U367 ( .A(n346), .B(n577), .CI(n343), .CO(n340), .S(n341) );
  FA_X1 U368 ( .A(n591), .B(n348), .CI(n606), .CO(n342), .S(n343) );
  FA_X1 U369 ( .A(n347), .B(n354), .CI(n352), .CO(n344), .S(n345) );
  FA_X1 U370 ( .A(n578), .B(n592), .CI(n349), .CO(n346), .S(n347) );
  FA_X1 U372 ( .A(n358), .B(n355), .CI(n353), .CO(n350), .S(n351) );
  FA_X1 U373 ( .A(n362), .B(n607), .CI(n360), .CO(n352), .S(n353) );
  FA_X1 U374 ( .A(n593), .B(n579), .CI(n622), .CO(n354), .S(n355) );
  FA_X1 U375 ( .A(n359), .B(n361), .CI(n366), .CO(n356), .S(n357) );
  FA_X1 U376 ( .A(n370), .B(n363), .CI(n368), .CO(n358), .S(n359) );
  FA_X1 U377 ( .A(n580), .B(n594), .CI(n608), .CO(n360), .S(n361) );
  FA_X1 U379 ( .A(n367), .B(n376), .CI(n374), .CO(n364), .S(n365) );
  FA_X1 U380 ( .A(n369), .B(n378), .CI(n371), .CO(n366), .S(n367) );
  FA_X1 U381 ( .A(n595), .B(n609), .CI(n380), .CO(n368), .S(n369) );
  FA_X1 U382 ( .A(n623), .B(n581), .CI(n638), .CO(n370), .S(n371) );
  FA_X1 U383 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  FA_X1 U384 ( .A(n379), .B(n388), .CI(n386), .CO(n374), .S(n375) );
  FA_X1 U385 ( .A(n381), .B(n610), .CI(n390), .CO(n376), .S(n377) );
  FA_X1 U386 ( .A(n624), .B(n596), .CI(n582), .CO(n378), .S(n379) );
  FA_X1 U388 ( .A(n394), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U389 ( .A(n391), .B(n389), .CI(n396), .CO(n384), .S(n385) );
  FA_X1 U390 ( .A(n400), .B(n625), .CI(n398), .CO(n386), .S(n387) );
  FA_X1 U391 ( .A(n597), .B(n639), .CI(n611), .CO(n388), .S(n389) );
  FA_X1 U392 ( .A(n1033), .B(n583), .CI(n654), .CO(n390), .S(n391) );
  FA_X1 U395 ( .A(n412), .B(n414), .CI(n401), .CO(n396), .S(n397) );
  FA_X1 U396 ( .A(n584), .B(n598), .CI(n403), .CO(n398), .S(n399) );
  FA_X1 U397 ( .A(n612), .B(n626), .CI(n640), .CO(n400), .S(n401) );
  FA_X1 U400 ( .A(n411), .B(n420), .CI(n422), .CO(n406), .S(n407) );
  FA_X1 U401 ( .A(n413), .B(n424), .CI(n415), .CO(n408), .S(n409) );
  FA_X1 U402 ( .A(n613), .B(n627), .CI(n426), .CO(n410), .S(n411) );
  FA_X1 U403 ( .A(n641), .B(n655), .CI(n599), .CO(n412), .S(n413) );
  FA_X1 U404 ( .A(n428), .B(n585), .CI(n670), .CO(n414), .S(n415) );
  FA_X1 U405 ( .A(n432), .B(n421), .CI(n419), .CO(n416), .S(n417) );
  FA_X1 U406 ( .A(n423), .B(n436), .CI(n434), .CO(n418), .S(n419) );
  FA_X1 U407 ( .A(n425), .B(n438), .CI(n427), .CO(n420), .S(n421) );
  FA_X1 U409 ( .A(n600), .B(n628), .CI(n642), .CO(n424), .S(n425) );
  FA_X1 U410 ( .A(n656), .B(n586), .CI(n614), .CO(n426), .S(n427) );
  FA_X1 U413 ( .A(n437), .B(n450), .CI(n448), .CO(n432), .S(n433) );
  FA_X1 U414 ( .A(n439), .B(n452), .CI(n441), .CO(n434), .S(n435) );
  FA_X1 U415 ( .A(n443), .B(n456), .CI(n454), .CO(n436), .S(n437) );
  FA_X1 U416 ( .A(n671), .B(n657), .CI(n615), .CO(n438), .S(n439) );
  FA_X1 U417 ( .A(n686), .B(n629), .CI(n587), .CO(n440), .S(n441) );
  FA_X1 U421 ( .A(n462), .B(n455), .CI(n451), .CO(n446), .S(n447) );
  FA_X1 U422 ( .A(n464), .B(n466), .CI(n453), .CO(n448), .S(n449) );
  FA_X1 U423 ( .A(n457), .B(n672), .CI(n468), .CO(n450), .S(n451) );
  FA_X1 U424 ( .A(n687), .B(n630), .CI(n658), .CO(n452), .S(n453) );
  FA_X1 U425 ( .A(n602), .B(n644), .CI(n616), .CO(n454), .S(n455) );
  HA_X1 U426 ( .A(n566), .B(n588), .CO(n456), .S(n457) );
  FA_X1 U427 ( .A(n463), .B(n472), .CI(n461), .CO(n458), .S(n459) );
  FA_X1 U428 ( .A(n465), .B(n467), .CI(n474), .CO(n460), .S(n461) );
  FA_X1 U429 ( .A(n476), .B(n478), .CI(n469), .CO(n462), .S(n463) );
  FA_X1 U430 ( .A(n645), .B(n659), .CI(n480), .CO(n464), .S(n465) );
  FA_X1 U431 ( .A(n603), .B(n673), .CI(n631), .CO(n466), .S(n467) );
  FA_X1 U432 ( .A(n617), .B(n589), .CI(n688), .CO(n468), .S(n469) );
  FA_X1 U434 ( .A(n479), .B(n477), .CI(n486), .CO(n472), .S(n473) );
  FA_X1 U435 ( .A(n490), .B(n481), .CI(n488), .CO(n474), .S(n475) );
  FA_X1 U436 ( .A(n618), .B(n660), .CI(n632), .CO(n476), .S(n477) );
  FA_X1 U437 ( .A(n689), .B(n674), .CI(n646), .CO(n478), .S(n479) );
  HA_X1 U438 ( .A(n604), .B(n567), .CO(n480), .S(n481) );
  FA_X1 U440 ( .A(n491), .B(n489), .CI(n496), .CO(n484), .S(n485) );
  FA_X1 U441 ( .A(n958), .B(n661), .CI(n498), .CO(n486), .S(n487) );
  FA_X1 U442 ( .A(n619), .B(n675), .CI(n647), .CO(n488), .S(n489) );
  FA_X1 U443 ( .A(n690), .B(n605), .CI(n633), .CO(n490), .S(n491) );
  FA_X1 U444 ( .A(n504), .B(n497), .CI(n495), .CO(n492), .S(n493) );
  FA_X1 U445 ( .A(n506), .B(n508), .CI(n499), .CO(n494), .S(n495) );
  FA_X1 U446 ( .A(n648), .B(n676), .CI(n501), .CO(n496), .S(n497) );
  FA_X1 U447 ( .A(n634), .B(n662), .CI(n691), .CO(n498), .S(n499) );
  FA_X1 U449 ( .A(n512), .B(n507), .CI(n505), .CO(n502), .S(n503) );
  FA_X1 U450 ( .A(n514), .B(n516), .CI(n509), .CO(n504), .S(n505) );
  FA_X1 U451 ( .A(n635), .B(n663), .CI(n677), .CO(n506), .S(n507) );
  FA_X1 U452 ( .A(n692), .B(n621), .CI(n649), .CO(n508), .S(n509) );
  FA_X1 U453 ( .A(n515), .B(n520), .CI(n513), .CO(n510), .S(n511) );
  FA_X1 U454 ( .A(n517), .B(n693), .CI(n522), .CO(n512), .S(n513) );
  FA_X1 U455 ( .A(n650), .B(n664), .CI(n678), .CO(n514), .S(n515) );
  HA_X1 U456 ( .A(n569), .B(n636), .CO(n516), .S(n517) );
  FA_X1 U457 ( .A(n523), .B(n526), .CI(n521), .CO(n518), .S(n519) );
  FA_X1 U458 ( .A(n651), .B(n679), .CI(n528), .CO(n520), .S(n521) );
  FA_X1 U459 ( .A(n665), .B(n637), .CI(n694), .CO(n522), .S(n523) );
  FA_X1 U460 ( .A(n532), .B(n529), .CI(n527), .CO(n524), .S(n525) );
  FA_X1 U461 ( .A(n666), .B(n695), .CI(n680), .CO(n526), .S(n527) );
  HA_X1 U462 ( .A(n570), .B(n652), .CO(n528), .S(n529) );
  FA_X1 U463 ( .A(n536), .B(n667), .CI(n533), .CO(n530), .S(n531) );
  FA_X1 U464 ( .A(n696), .B(n653), .CI(n681), .CO(n532), .S(n533) );
  FA_X1 U465 ( .A(n682), .B(n697), .CI(n537), .CO(n534), .S(n535) );
  HA_X1 U466 ( .A(n668), .B(n571), .CO(n536), .S(n537) );
  FA_X1 U467 ( .A(n698), .B(n669), .CI(n683), .CO(n538), .S(n539) );
  HA_X1 U468 ( .A(n684), .B(n699), .CO(n540), .S(n541) );
  AOI21_X1 U822 ( .B1(n273), .B2(n982), .A(n270), .ZN(n953) );
  AOI21_X2 U823 ( .B1(n980), .B2(n297), .A(n294), .ZN(n292) );
  BUF_X1 U824 ( .A(n150), .Z(n954) );
  CLKBUF_X3 U825 ( .A(b[4]), .Z(n849) );
  XNOR2_X1 U826 ( .A(n407), .B(n1006), .ZN(n955) );
  CLKBUF_X1 U827 ( .A(n418), .Z(n956) );
  BUF_X2 U828 ( .A(b[13]), .Z(n840) );
  CLKBUF_X1 U829 ( .A(n417), .Z(n957) );
  CLKBUF_X3 U830 ( .A(b[12]), .Z(n841) );
  BUF_X1 U831 ( .A(b[9]), .Z(n844) );
  BUF_X4 U832 ( .A(a[3]), .Z(n7) );
  BUF_X4 U833 ( .A(a[1]), .Z(n1) );
  CLKBUF_X1 U834 ( .A(n868), .Z(n12) );
  BUF_X1 U835 ( .A(n875), .Z(n16) );
  BUF_X1 U836 ( .A(n49), .Z(n1045) );
  AND2_X1 U837 ( .A1(n968), .A2(n568), .ZN(n958) );
  OR2_X1 U838 ( .A1(n503), .A2(n510), .ZN(n959) );
  BUF_X1 U839 ( .A(n1057), .Z(n1015) );
  XOR2_X1 U840 ( .A(n494), .B(n487), .Z(n960) );
  XOR2_X1 U841 ( .A(n485), .B(n960), .Z(n483) );
  NAND2_X1 U842 ( .A1(n485), .A2(n494), .ZN(n961) );
  NAND2_X1 U843 ( .A1(n485), .A2(n487), .ZN(n962) );
  NAND2_X1 U844 ( .A1(n494), .A2(n487), .ZN(n963) );
  NAND3_X1 U845 ( .A1(n961), .A2(n962), .A3(n963), .ZN(n482) );
  AOI21_X2 U846 ( .B1(n198), .B2(n151), .A(n152), .ZN(n150) );
  NOR2_X1 U847 ( .A1(n459), .A2(n470), .ZN(n964) );
  NOR2_X1 U848 ( .A1(n459), .A2(n470), .ZN(n238) );
  OAI21_X1 U849 ( .B1(n953), .B2(n256), .A(n257), .ZN(n965) );
  CLKBUF_X1 U850 ( .A(n281), .Z(n966) );
  CLKBUF_X1 U851 ( .A(n18), .Z(n967) );
  CLKBUF_X1 U852 ( .A(b[15]), .Z(n1021) );
  XOR2_X1 U853 ( .A(n620), .B(n568), .Z(n501) );
  CLKBUF_X1 U854 ( .A(n620), .Z(n968) );
  CLKBUF_X1 U855 ( .A(n871), .Z(n40) );
  XNOR2_X1 U856 ( .A(n433), .B(n969), .ZN(n431) );
  XNOR2_X1 U857 ( .A(n446), .B(n435), .ZN(n969) );
  BUF_X1 U858 ( .A(n49), .Z(n1058) );
  XOR2_X1 U859 ( .A(n484), .B(n475), .Z(n970) );
  XOR2_X1 U860 ( .A(n473), .B(n970), .Z(n471) );
  NAND2_X1 U861 ( .A1(n473), .A2(n484), .ZN(n971) );
  NAND2_X1 U862 ( .A1(n473), .A2(n475), .ZN(n972) );
  NAND2_X1 U863 ( .A1(n484), .A2(n475), .ZN(n973) );
  NAND3_X1 U864 ( .A1(n971), .A2(n972), .A3(n973), .ZN(n470) );
  BUF_X2 U865 ( .A(a[5]), .Z(n974) );
  CLKBUF_X1 U866 ( .A(a[5]), .Z(n13) );
  BUF_X1 U867 ( .A(b[8]), .Z(n845) );
  XNOR2_X1 U868 ( .A(n440), .B(n975), .ZN(n423) );
  XNOR2_X1 U869 ( .A(n429), .B(n442), .ZN(n975) );
  BUF_X2 U870 ( .A(n871), .Z(n39) );
  BUF_X2 U871 ( .A(a[9]), .Z(n1030) );
  BUF_X2 U872 ( .A(n846), .Z(n1038) );
  BUF_X2 U873 ( .A(b[11]), .Z(n842) );
  OAI22_X1 U874 ( .A1(n48), .A2(n703), .B1(n46), .B2(n702), .ZN(n332) );
  OR2_X1 U875 ( .A1(n337), .A2(n340), .ZN(n976) );
  OR2_X1 U876 ( .A1(n334), .A2(n333), .ZN(n977) );
  OR2_X1 U877 ( .A1(n493), .A2(n502), .ZN(n978) );
  OR2_X1 U878 ( .A1(n574), .A2(n332), .ZN(n979) );
  OR2_X1 U879 ( .A1(n541), .A2(n572), .ZN(n980) );
  OR2_X1 U880 ( .A1(n336), .A2(n335), .ZN(n981) );
  OR2_X1 U881 ( .A1(n511), .A2(n518), .ZN(n982) );
  OR2_X1 U882 ( .A1(n525), .A2(n530), .ZN(n983) );
  OR2_X1 U883 ( .A1(n535), .A2(n538), .ZN(n984) );
  OR2_X1 U884 ( .A1(n471), .A2(n482), .ZN(n985) );
  BUF_X1 U885 ( .A(n226), .Z(n1034) );
  OR2_X1 U886 ( .A1(n701), .A2(n573), .ZN(n986) );
  NOR2_X1 U887 ( .A1(n345), .A2(n350), .ZN(n144) );
  NOR2_X1 U888 ( .A1(n373), .A2(n382), .ZN(n190) );
  OR2_X2 U889 ( .A1(n643), .A2(n601), .ZN(n442) );
  CLKBUF_X2 U890 ( .A(b[3]), .Z(n850) );
  CLKBUF_X1 U891 ( .A(n1019), .Z(n987) );
  AND2_X1 U892 ( .A1(n471), .A2(n482), .ZN(n1019) );
  CLKBUF_X1 U893 ( .A(n847), .Z(n988) );
  BUF_X2 U894 ( .A(b[6]), .Z(n847) );
  BUF_X1 U895 ( .A(b[0]), .Z(n49) );
  NAND2_X1 U896 ( .A1(n433), .A2(n446), .ZN(n989) );
  NAND2_X1 U897 ( .A1(n433), .A2(n435), .ZN(n990) );
  NAND2_X1 U898 ( .A1(n446), .A2(n435), .ZN(n991) );
  NAND3_X1 U899 ( .A1(n989), .A2(n990), .A3(n991), .ZN(n430) );
  BUF_X1 U900 ( .A(n846), .Z(n1037) );
  BUF_X1 U901 ( .A(n867), .Z(n17) );
  XNOR2_X1 U902 ( .A(n992), .B(n395), .ZN(n393) );
  XNOR2_X1 U903 ( .A(n397), .B(n406), .ZN(n992) );
  XOR2_X1 U904 ( .A(n410), .B(n399), .Z(n993) );
  XOR2_X1 U905 ( .A(n993), .B(n408), .Z(n395) );
  NAND2_X1 U906 ( .A1(n410), .A2(n399), .ZN(n994) );
  NAND2_X1 U907 ( .A1(n410), .A2(n408), .ZN(n995) );
  NAND2_X1 U908 ( .A1(n399), .A2(n408), .ZN(n996) );
  NAND3_X1 U909 ( .A1(n994), .A2(n995), .A3(n996), .ZN(n394) );
  NAND2_X1 U910 ( .A1(n397), .A2(n406), .ZN(n997) );
  NAND2_X1 U911 ( .A1(n397), .A2(n395), .ZN(n998) );
  NAND2_X1 U912 ( .A1(n406), .A2(n395), .ZN(n999) );
  NAND3_X1 U913 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n392) );
  CLKBUF_X1 U914 ( .A(n24), .Z(n23) );
  BUF_X2 U915 ( .A(n866), .Z(n24) );
  NAND2_X1 U916 ( .A1(n440), .A2(n429), .ZN(n1000) );
  NAND2_X1 U917 ( .A1(n440), .A2(n442), .ZN(n1001) );
  NAND2_X1 U918 ( .A1(n429), .A2(n442), .ZN(n1002) );
  NAND3_X1 U919 ( .A1(n1000), .A2(n1001), .A3(n1002), .ZN(n422) );
  OR2_X1 U920 ( .A1(n365), .A2(n372), .ZN(n1003) );
  NOR2_X1 U921 ( .A1(n483), .A2(n492), .ZN(n252) );
  CLKBUF_X1 U922 ( .A(n219), .Z(n1004) );
  CLKBUF_X1 U923 ( .A(n42), .Z(n1005) );
  XNOR2_X1 U924 ( .A(n407), .B(n1006), .ZN(n405) );
  XNOR2_X1 U925 ( .A(n418), .B(n409), .ZN(n1006) );
  NAND2_X1 U926 ( .A1(n407), .A2(n956), .ZN(n1007) );
  NAND2_X1 U927 ( .A1(n407), .A2(n409), .ZN(n1008) );
  NAND2_X1 U928 ( .A1(n956), .A2(n409), .ZN(n1009) );
  NAND3_X1 U929 ( .A1(n1007), .A2(n1008), .A3(n1009), .ZN(n404) );
  XNOR2_X1 U930 ( .A(n850), .B(n25), .ZN(n1010) );
  CLKBUF_X2 U931 ( .A(n872), .Z(n34) );
  BUF_X1 U932 ( .A(n872), .Z(n33) );
  CLKBUF_X3 U933 ( .A(a[11]), .Z(n1011) );
  CLKBUF_X1 U934 ( .A(a[11]), .Z(n31) );
  XNOR2_X1 U935 ( .A(n25), .B(n851), .ZN(n1012) );
  BUF_X1 U936 ( .A(n865), .Z(n29) );
  BUF_X1 U937 ( .A(n874), .Z(n22) );
  CLKBUF_X2 U938 ( .A(n874), .Z(n21) );
  CLKBUF_X3 U939 ( .A(b[1]), .Z(n852) );
  OR2_X1 U940 ( .A1(n955), .A2(n416), .ZN(n1013) );
  CLKBUF_X1 U941 ( .A(n276), .Z(n1014) );
  BUF_X2 U942 ( .A(n49), .Z(n1057) );
  INV_X1 U943 ( .A(n884), .ZN(n1016) );
  NOR2_X1 U944 ( .A1(n957), .A2(n430), .ZN(n1017) );
  NOR2_X1 U945 ( .A1(n417), .A2(n430), .ZN(n218) );
  OR2_X1 U946 ( .A1(n471), .A2(n482), .ZN(n1018) );
  BUF_X1 U947 ( .A(n873), .Z(n28) );
  CLKBUF_X2 U948 ( .A(n873), .Z(n27) );
  CLKBUF_X1 U949 ( .A(n1031), .Z(n1020) );
  CLKBUF_X1 U950 ( .A(b[15]), .Z(n838) );
  CLKBUF_X1 U951 ( .A(n284), .Z(n1022) );
  INV_X1 U952 ( .A(n987), .ZN(n1023) );
  NOR2_X1 U953 ( .A1(n393), .A2(n404), .ZN(n204) );
  XNOR2_X1 U954 ( .A(n146), .B(n1024), .ZN(product[25]) );
  AND2_X1 U955 ( .A1(n143), .A2(n145), .ZN(n1024) );
  NOR2_X1 U956 ( .A1(n218), .A2(n211), .ZN(n1025) );
  NOR2_X1 U957 ( .A1(n955), .A2(n416), .ZN(n1026) );
  BUF_X2 U958 ( .A(b[10]), .Z(n843) );
  OR2_X1 U959 ( .A1(n227), .A2(n232), .ZN(n1027) );
  BUF_X2 U960 ( .A(n866), .Z(n1028) );
  XNOR2_X1 U961 ( .A(n139), .B(n1029), .ZN(product[26]) );
  AND2_X1 U962 ( .A1(n306), .A2(n138), .ZN(n1029) );
  CLKBUF_X1 U963 ( .A(a[9]), .Z(n25) );
  BUF_X1 U964 ( .A(n206), .Z(n1031) );
  NOR2_X1 U965 ( .A1(n431), .A2(n444), .ZN(n1032) );
  BUF_X1 U966 ( .A(n206), .Z(n51) );
  OAI22_X1 U967 ( .A1(n18), .A2(n788), .B1(n16), .B2(n787), .ZN(n1033) );
  CLKBUF_X1 U968 ( .A(n839), .Z(n1035) );
  BUF_X2 U969 ( .A(n206), .Z(n1036) );
  BUF_X1 U970 ( .A(b[5]), .Z(n848) );
  BUF_X1 U971 ( .A(b[7]), .Z(n846) );
  NOR2_X1 U972 ( .A1(n357), .A2(n364), .ZN(n168) );
  CLKBUF_X3 U973 ( .A(b[2]), .Z(n851) );
  XNOR2_X1 U974 ( .A(n201), .B(n1039), .ZN(product[20]) );
  AND2_X1 U975 ( .A1(n312), .A2(n200), .ZN(n1039) );
  AOI21_X1 U976 ( .B1(n985), .B2(n251), .A(n987), .ZN(n1040) );
  XOR2_X1 U977 ( .A(n460), .B(n449), .Z(n1041) );
  XOR2_X1 U978 ( .A(n447), .B(n1041), .Z(n445) );
  NAND2_X1 U979 ( .A1(n447), .A2(n460), .ZN(n1042) );
  NAND2_X1 U980 ( .A1(n447), .A2(n449), .ZN(n1043) );
  NAND2_X1 U981 ( .A1(n460), .A2(n449), .ZN(n1044) );
  NAND3_X1 U982 ( .A1(n1042), .A2(n1043), .A3(n1044), .ZN(n444) );
  NOR2_X1 U983 ( .A1(n431), .A2(n444), .ZN(n227) );
  XNOR2_X1 U984 ( .A(n192), .B(n1046), .ZN(product[21]) );
  AND2_X1 U985 ( .A1(n188), .A2(n191), .ZN(n1046) );
  BUF_X1 U986 ( .A(n867), .Z(n1047) );
  INV_X1 U987 ( .A(n198), .ZN(n196) );
  INV_X1 U988 ( .A(n197), .ZN(n195) );
  NAND2_X1 U989 ( .A1(n188), .A2(n175), .ZN(n173) );
  XNOR2_X1 U990 ( .A(n170), .B(n1048), .ZN(product[23]) );
  AND2_X1 U991 ( .A1(n167), .A2(n169), .ZN(n1048) );
  XNOR2_X1 U992 ( .A(n159), .B(n1049), .ZN(product[24]) );
  AND2_X1 U993 ( .A1(n308), .A2(n158), .ZN(n1049) );
  AOI21_X1 U994 ( .B1(n1018), .B2(n251), .A(n1019), .ZN(n242) );
  XNOR2_X1 U995 ( .A(n130), .B(n1050), .ZN(product[27]) );
  AND2_X1 U996 ( .A1(n976), .A2(n129), .ZN(n1050) );
  XNOR2_X1 U997 ( .A(n183), .B(n1051), .ZN(product[22]) );
  AND2_X1 U998 ( .A1(n175), .A2(n182), .ZN(n1051) );
  XNOR2_X1 U999 ( .A(n117), .B(n1052), .ZN(product[28]) );
  AND2_X1 U1000 ( .A1(n981), .A2(n116), .ZN(n1052) );
  XNOR2_X1 U1001 ( .A(n106), .B(n1053), .ZN(product[29]) );
  AND2_X1 U1002 ( .A1(n977), .A2(n105), .ZN(n1053) );
  XNOR2_X1 U1003 ( .A(n93), .B(n1054), .ZN(product[30]) );
  AND2_X1 U1004 ( .A1(n979), .A2(n92), .ZN(n1054) );
  NAND2_X1 U1005 ( .A1(n417), .A2(n430), .ZN(n219) );
  NAND2_X1 U1006 ( .A1(n483), .A2(n492), .ZN(n253) );
  NOR2_X1 U1007 ( .A1(n341), .A2(n344), .ZN(n137) );
  NOR2_X1 U1008 ( .A1(n700), .A2(n685), .ZN(n298) );
  NOR2_X1 U1009 ( .A1(n531), .A2(n534), .ZN(n282) );
  AND2_X1 U1010 ( .A1(n986), .A2(n301), .ZN(product[1]) );
  XOR2_X1 U1011 ( .A(a[14]), .B(a[15]), .Z(n854) );
  NOR2_X1 U1012 ( .A1(n195), .A2(n173), .ZN(n171) );
  NOR2_X1 U1013 ( .A1(n195), .A2(n186), .ZN(n184) );
  NOR2_X1 U1014 ( .A1(n195), .A2(n162), .ZN(n160) );
  NOR2_X1 U1015 ( .A1(n149), .A2(n124), .ZN(n118) );
  NOR2_X1 U1016 ( .A1(n149), .A2(n96), .ZN(n94) );
  NOR2_X1 U1017 ( .A1(n149), .A2(n109), .ZN(n107) );
  INV_X1 U1018 ( .A(n177), .ZN(n175) );
  INV_X1 U1019 ( .A(n1027), .ZN(n221) );
  INV_X1 U1020 ( .A(n98), .ZN(n96) );
  INV_X1 U1021 ( .A(n196), .ZN(n194) );
  INV_X1 U1022 ( .A(n149), .ZN(n147) );
  NOR2_X1 U1023 ( .A1(n177), .A2(n166), .ZN(n164) );
  NOR2_X1 U1024 ( .A1(n124), .A2(n100), .ZN(n98) );
  OAI21_X1 U1025 ( .B1(n196), .B2(n173), .A(n174), .ZN(n172) );
  AOI21_X1 U1026 ( .B1(n189), .B2(n175), .A(n1056), .ZN(n174) );
  INV_X1 U1027 ( .A(n1034), .ZN(n224) );
  XNOR2_X1 U1028 ( .A(n240), .B(n70), .ZN(product[14]) );
  NAND2_X1 U1029 ( .A1(n318), .A2(n239), .ZN(n70) );
  OAI21_X1 U1030 ( .B1(n254), .B2(n241), .A(n1040), .ZN(n240) );
  INV_X1 U1031 ( .A(n964), .ZN(n318) );
  INV_X1 U1032 ( .A(n953), .ZN(n267) );
  NOR2_X1 U1033 ( .A1(n1027), .A2(n1017), .ZN(n214) );
  OAI21_X1 U1034 ( .B1(n196), .B2(n186), .A(n191), .ZN(n185) );
  NAND2_X1 U1035 ( .A1(n164), .A2(n188), .ZN(n162) );
  INV_X1 U1036 ( .A(n188), .ZN(n186) );
  INV_X1 U1037 ( .A(n1003), .ZN(n177) );
  NAND2_X1 U1038 ( .A1(n985), .A2(n320), .ZN(n241) );
  NOR2_X1 U1039 ( .A1(n149), .A2(n133), .ZN(n131) );
  NOR2_X1 U1040 ( .A1(n149), .A2(n144), .ZN(n140) );
  INV_X1 U1041 ( .A(n124), .ZN(n122) );
  NAND2_X1 U1042 ( .A1(n122), .A2(n981), .ZN(n109) );
  INV_X1 U1043 ( .A(n251), .ZN(n249) );
  NAND2_X1 U1044 ( .A1(n313), .A2(n205), .ZN(n65) );
  INV_X1 U1045 ( .A(n204), .ZN(n313) );
  NAND2_X1 U1046 ( .A1(n982), .A2(n272), .ZN(n75) );
  XOR2_X1 U1047 ( .A(n254), .B(n72), .Z(product[12]) );
  NAND2_X1 U1048 ( .A1(n320), .A2(n253), .ZN(n72) );
  INV_X1 U1049 ( .A(n252), .ZN(n320) );
  XNOR2_X1 U1050 ( .A(n234), .B(n69), .ZN(product[15]) );
  NAND2_X1 U1051 ( .A1(n317), .A2(n233), .ZN(n69) );
  XNOR2_X1 U1052 ( .A(n247), .B(n71), .ZN(product[13]) );
  NAND2_X1 U1053 ( .A1(n985), .A2(n1023), .ZN(n71) );
  OAI21_X1 U1054 ( .B1(n254), .B2(n252), .A(n249), .ZN(n247) );
  XNOR2_X1 U1055 ( .A(n267), .B(n74), .ZN(product[10]) );
  NAND2_X1 U1056 ( .A1(n959), .A2(n266), .ZN(n74) );
  XOR2_X1 U1057 ( .A(n229), .B(n68), .Z(product[16]) );
  NAND2_X1 U1058 ( .A1(n316), .A2(n228), .ZN(n68) );
  INV_X1 U1059 ( .A(n1032), .ZN(n316) );
  INV_X1 U1060 ( .A(n157), .ZN(n308) );
  XOR2_X1 U1061 ( .A(n262), .B(n73), .Z(product[11]) );
  NAND2_X1 U1062 ( .A1(n978), .A2(n261), .ZN(n73) );
  AOI21_X1 U1063 ( .B1(n267), .B2(n959), .A(n264), .ZN(n262) );
  NAND2_X1 U1064 ( .A1(n978), .A2(n959), .ZN(n256) );
  AOI21_X1 U1065 ( .B1(n978), .B2(n264), .A(n259), .ZN(n257) );
  XOR2_X1 U1066 ( .A(n220), .B(n67), .Z(product[17]) );
  NAND2_X1 U1067 ( .A1(n217), .A2(n1004), .ZN(n67) );
  AOI21_X1 U1068 ( .B1(n234), .B2(n221), .A(n1034), .ZN(n220) );
  XOR2_X1 U1069 ( .A(n213), .B(n66), .Z(product[18]) );
  NAND2_X1 U1070 ( .A1(n1013), .A2(n212), .ZN(n66) );
  AOI21_X1 U1071 ( .B1(n214), .B2(n234), .A(n215), .ZN(n213) );
  AOI21_X1 U1072 ( .B1(n273), .B2(n982), .A(n270), .ZN(n268) );
  INV_X1 U1073 ( .A(n272), .ZN(n270) );
  OAI21_X1 U1074 ( .B1(n196), .B2(n162), .A(n163), .ZN(n161) );
  AOI21_X1 U1075 ( .B1(n164), .B2(n189), .A(n165), .ZN(n163) );
  OAI21_X1 U1076 ( .B1(n182), .B2(n166), .A(n169), .ZN(n165) );
  INV_X1 U1077 ( .A(n136), .ZN(n134) );
  INV_X1 U1078 ( .A(n99), .ZN(n97) );
  AOI21_X1 U1079 ( .B1(n123), .B2(n981), .A(n114), .ZN(n110) );
  OAI21_X1 U1080 ( .B1(n224), .B2(n1017), .A(n1004), .ZN(n215) );
  INV_X1 U1081 ( .A(n190), .ZN(n188) );
  INV_X1 U1082 ( .A(n191), .ZN(n189) );
  NAND2_X1 U1083 ( .A1(n98), .A2(n979), .ZN(n87) );
  NAND2_X1 U1084 ( .A1(n981), .A2(n977), .ZN(n100) );
  NAND2_X1 U1085 ( .A1(n135), .A2(n976), .ZN(n124) );
  NAND2_X1 U1086 ( .A1(n459), .A2(n470), .ZN(n239) );
  NOR2_X1 U1087 ( .A1(n149), .A2(n87), .ZN(n85) );
  OAI21_X1 U1088 ( .B1(n954), .B2(n87), .A(n88), .ZN(n86) );
  INV_X1 U1089 ( .A(n253), .ZN(n251) );
  INV_X1 U1090 ( .A(n1017), .ZN(n217) );
  INV_X1 U1091 ( .A(n167), .ZN(n166) );
  INV_X1 U1092 ( .A(n168), .ZN(n167) );
  INV_X1 U1093 ( .A(n266), .ZN(n264) );
  INV_X1 U1094 ( .A(n125), .ZN(n123) );
  INV_X1 U1095 ( .A(n135), .ZN(n133) );
  INV_X1 U1096 ( .A(n144), .ZN(n143) );
  INV_X1 U1097 ( .A(n261), .ZN(n259) );
  INV_X1 U1098 ( .A(n205), .ZN(n203) );
  INV_X1 U1099 ( .A(n233), .ZN(n231) );
  NAND2_X1 U1100 ( .A1(n326), .A2(n283), .ZN(n78) );
  INV_X1 U1101 ( .A(n282), .ZN(n326) );
  NAND2_X1 U1102 ( .A1(n324), .A2(n275), .ZN(n76) );
  INV_X1 U1103 ( .A(n274), .ZN(n324) );
  NAND2_X1 U1104 ( .A1(n983), .A2(n280), .ZN(n77) );
  NAND2_X1 U1105 ( .A1(n984), .A2(n288), .ZN(n79) );
  INV_X1 U1106 ( .A(n137), .ZN(n306) );
  NOR2_X1 U1107 ( .A1(n351), .A2(n356), .ZN(n157) );
  AOI21_X1 U1108 ( .B1(n136), .B2(n976), .A(n127), .ZN(n125) );
  INV_X1 U1109 ( .A(n129), .ZN(n127) );
  OAI21_X1 U1110 ( .B1(n145), .B2(n137), .A(n138), .ZN(n136) );
  OAI21_X1 U1111 ( .B1(n125), .B2(n100), .A(n101), .ZN(n99) );
  AOI21_X1 U1112 ( .B1(n114), .B2(n977), .A(n103), .ZN(n101) );
  INV_X1 U1113 ( .A(n105), .ZN(n103) );
  OAI21_X1 U1114 ( .B1(n282), .B2(n284), .A(n283), .ZN(n281) );
  AOI21_X1 U1115 ( .B1(n281), .B2(n983), .A(n278), .ZN(n276) );
  INV_X1 U1116 ( .A(n280), .ZN(n278) );
  NAND2_X1 U1117 ( .A1(n393), .A2(n404), .ZN(n205) );
  NOR2_X1 U1118 ( .A1(n445), .A2(n458), .ZN(n232) );
  NOR2_X1 U1119 ( .A1(n144), .A2(n137), .ZN(n135) );
  AOI21_X1 U1120 ( .B1(n99), .B2(n979), .A(n90), .ZN(n88) );
  INV_X1 U1121 ( .A(n92), .ZN(n90) );
  NAND2_X1 U1122 ( .A1(n345), .A2(n350), .ZN(n145) );
  NAND2_X1 U1123 ( .A1(n373), .A2(n382), .ZN(n191) );
  NAND2_X1 U1124 ( .A1(n357), .A2(n364), .ZN(n169) );
  NAND2_X1 U1125 ( .A1(n445), .A2(n458), .ZN(n233) );
  NAND2_X1 U1126 ( .A1(n511), .A2(n518), .ZN(n272) );
  NAND2_X1 U1127 ( .A1(n503), .A2(n510), .ZN(n266) );
  NAND2_X1 U1128 ( .A1(n493), .A2(n502), .ZN(n261) );
  NAND2_X1 U1129 ( .A1(n431), .A2(n444), .ZN(n228) );
  NAND2_X1 U1130 ( .A1(n955), .A2(n416), .ZN(n212) );
  NAND2_X1 U1131 ( .A1(n383), .A2(n392), .ZN(n200) );
  INV_X1 U1132 ( .A(n116), .ZN(n114) );
  AOI21_X1 U1133 ( .B1(n984), .B2(n289), .A(n286), .ZN(n284) );
  INV_X1 U1134 ( .A(n288), .ZN(n286) );
  XOR2_X1 U1135 ( .A(n82), .B(n301), .Z(product[2]) );
  NAND2_X1 U1136 ( .A1(n330), .A2(n299), .ZN(n82) );
  INV_X1 U1137 ( .A(n298), .ZN(n330) );
  XNOR2_X1 U1138 ( .A(n81), .B(n297), .ZN(product[3]) );
  OAI21_X1 U1139 ( .B1(n292), .B2(n290), .A(n291), .ZN(n289) );
  OAI21_X1 U1140 ( .B1(n298), .B2(n301), .A(n299), .ZN(n297) );
  NAND2_X1 U1141 ( .A1(n574), .A2(n332), .ZN(n92) );
  NAND2_X1 U1142 ( .A1(n535), .A2(n538), .ZN(n288) );
  INV_X1 U1143 ( .A(n296), .ZN(n294) );
  INV_X1 U1144 ( .A(n332), .ZN(n333) );
  NOR2_X1 U1145 ( .A1(n519), .A2(n524), .ZN(n274) );
  NAND2_X1 U1146 ( .A1(n700), .A2(n685), .ZN(n299) );
  NAND2_X1 U1147 ( .A1(n337), .A2(n340), .ZN(n129) );
  NAND2_X1 U1148 ( .A1(n341), .A2(n344), .ZN(n138) );
  NAND2_X1 U1149 ( .A1(n336), .A2(n335), .ZN(n116) );
  NAND2_X1 U1150 ( .A1(n525), .A2(n530), .ZN(n280) );
  NAND2_X1 U1151 ( .A1(n334), .A2(n333), .ZN(n105) );
  NAND2_X1 U1152 ( .A1(n531), .A2(n534), .ZN(n283) );
  NAND2_X1 U1153 ( .A1(n519), .A2(n524), .ZN(n275) );
  NAND2_X1 U1154 ( .A1(n328), .A2(n291), .ZN(n80) );
  INV_X1 U1155 ( .A(n290), .ZN(n328) );
  OAI22_X1 U1156 ( .A1(n1005), .A2(n720), .B1(n40), .B2(n719), .ZN(n338) );
  OAI22_X1 U1157 ( .A1(n5), .A2(n835), .B1(n834), .B2(n3), .ZN(n700) );
  OAI22_X1 U1158 ( .A1(n12), .A2(n805), .B1(n10), .B2(n804), .ZN(n428) );
  OAI22_X1 U1159 ( .A1(n42), .A2(n731), .B1(n39), .B2(n730), .ZN(n601) );
  OAI22_X1 U1160 ( .A1(n30), .A2(n754), .B1(n27), .B2(n753), .ZN(n362) );
  OAI22_X1 U1161 ( .A1(n18), .A2(n788), .B1(n16), .B2(n787), .ZN(n402) );
  OAI22_X1 U1162 ( .A1(n48), .A2(n704), .B1(n46), .B2(n703), .ZN(n575) );
  INV_X1 U1163 ( .A(n545), .ZN(n590) );
  AOI21_X1 U1164 ( .B1(n1005), .B2(n40), .A(n719), .ZN(n545) );
  OAI22_X1 U1165 ( .A1(n48), .A2(n705), .B1(n46), .B2(n704), .ZN(n576) );
  INV_X1 U1166 ( .A(n338), .ZN(n339) );
  OAI22_X1 U1167 ( .A1(n48), .A2(n706), .B1(n46), .B2(n705), .ZN(n577) );
  OAI22_X1 U1168 ( .A1(n5), .A2(n833), .B1(n832), .B2(n3), .ZN(n698) );
  OAI22_X1 U1169 ( .A1(n11), .A2(n818), .B1(n9), .B2(n817), .ZN(n683) );
  AND2_X1 U1170 ( .A1(n1015), .A2(n558), .ZN(n669) );
  OAI22_X1 U1171 ( .A1(n48), .A2(n878), .B1(n718), .B2(n46), .ZN(n566) );
  OAI22_X1 U1172 ( .A1(n47), .A2(n717), .B1(n45), .B2(n716), .ZN(n588) );
  OR2_X1 U1173 ( .A1(n1058), .A2(n878), .ZN(n718) );
  OAI22_X1 U1174 ( .A1(n11), .A2(n813), .B1(n9), .B2(n812), .ZN(n678) );
  OAI22_X1 U1175 ( .A1(n24), .A2(n783), .B1(n21), .B2(n782), .ZN(n650) );
  OAI22_X1 U1176 ( .A1(n47), .A2(n711), .B1(n45), .B2(n710), .ZN(n582) );
  OAI22_X1 U1177 ( .A1(n42), .A2(n726), .B1(n40), .B2(n725), .ZN(n596) );
  OAI22_X1 U1178 ( .A1(n5), .A2(n832), .B1(n831), .B2(n3), .ZN(n697) );
  OAI22_X1 U1179 ( .A1(n11), .A2(n817), .B1(n9), .B2(n816), .ZN(n682) );
  NAND2_X1 U1180 ( .A1(n701), .A2(n573), .ZN(n301) );
  NOR2_X1 U1181 ( .A1(n539), .A2(n540), .ZN(n290) );
  AND2_X1 U1182 ( .A1(n1045), .A2(n561), .ZN(n685) );
  INV_X1 U1183 ( .A(n9), .ZN(n561) );
  OAI22_X1 U1184 ( .A1(n47), .A2(n712), .B1(n45), .B2(n711), .ZN(n583) );
  INV_X1 U1185 ( .A(n557), .ZN(n654) );
  OAI22_X1 U1186 ( .A1(n48), .A2(n707), .B1(n46), .B2(n706), .ZN(n578) );
  OAI22_X1 U1187 ( .A1(n1005), .A2(n722), .B1(n40), .B2(n721), .ZN(n592) );
  INV_X1 U1188 ( .A(n428), .ZN(n429) );
  OAI22_X1 U1189 ( .A1(n35), .A2(n744), .B1(n33), .B2(n743), .ZN(n613) );
  OAI22_X1 U1190 ( .A1(n11), .A2(n810), .B1(n10), .B2(n809), .ZN(n675) );
  OAI22_X1 U1191 ( .A1(n35), .A2(n750), .B1(n33), .B2(n749), .ZN(n619) );
  OAI22_X1 U1192 ( .A1(n24), .A2(n780), .B1(n21), .B2(n779), .ZN(n647) );
  OAI22_X1 U1193 ( .A1(n6), .A2(n824), .B1(n823), .B2(n4), .ZN(n689) );
  OAI22_X1 U1194 ( .A1(n11), .A2(n809), .B1(n10), .B2(n808), .ZN(n674) );
  OAI22_X1 U1195 ( .A1(n24), .A2(n779), .B1(n21), .B2(n778), .ZN(n646) );
  OAI22_X1 U1196 ( .A1(n17), .A2(n791), .B1(n16), .B2(n790), .ZN(n657) );
  OAI22_X1 U1197 ( .A1(n36), .A2(n746), .B1(n33), .B2(n745), .ZN(n615) );
  OAI22_X1 U1198 ( .A1(n12), .A2(n806), .B1(n805), .B2(n10), .ZN(n671) );
  OAI22_X1 U1199 ( .A1(n35), .A2(n740), .B1(n34), .B2(n739), .ZN(n609) );
  OAI22_X1 U1200 ( .A1(n48), .A2(n708), .B1(n46), .B2(n707), .ZN(n579) );
  OAI22_X1 U1201 ( .A1(n1005), .A2(n723), .B1(n40), .B2(n722), .ZN(n593) );
  INV_X1 U1202 ( .A(n551), .ZN(n622) );
  OAI22_X1 U1203 ( .A1(n825), .A2(n6), .B1(n824), .B2(n4), .ZN(n690) );
  OAI22_X1 U1204 ( .A1(n1010), .A2(n30), .B1(n28), .B2(n764), .ZN(n633) );
  AND2_X1 U1205 ( .A1(n1015), .A2(n546), .ZN(n605) );
  OAI22_X1 U1206 ( .A1(n18), .A2(n794), .B1(n16), .B2(n793), .ZN(n660) );
  OAI22_X1 U1207 ( .A1(n35), .A2(n749), .B1(n33), .B2(n748), .ZN(n618) );
  OAI22_X1 U1208 ( .A1(n30), .A2(n764), .B1(n27), .B2(n763), .ZN(n632) );
  OAI22_X1 U1209 ( .A1(n11), .A2(n812), .B1(n9), .B2(n811), .ZN(n677) );
  OAI22_X1 U1210 ( .A1(n30), .A2(n767), .B1(n27), .B2(n1012), .ZN(n635) );
  OAI22_X1 U1211 ( .A1(n18), .A2(n793), .B1(n16), .B2(n792), .ZN(n659) );
  OAI22_X1 U1212 ( .A1(n24), .A2(n778), .B1(n21), .B2(n777), .ZN(n645) );
  OAI22_X1 U1213 ( .A1(n47), .A2(n710), .B1(n45), .B2(n709), .ZN(n581) );
  OAI22_X1 U1214 ( .A1(n1005), .A2(n721), .B1(n40), .B2(n720), .ZN(n591) );
  INV_X1 U1215 ( .A(n548), .ZN(n606) );
  AOI21_X1 U1216 ( .B1(n35), .B2(n34), .A(n736), .ZN(n548) );
  OAI22_X1 U1217 ( .A1(n11), .A2(n814), .B1(n9), .B2(n813), .ZN(n679) );
  OAI22_X1 U1218 ( .A1(n23), .A2(n784), .B1(n21), .B2(n783), .ZN(n651) );
  OAI22_X1 U1219 ( .A1(n47), .A2(n714), .B1(n45), .B2(n713), .ZN(n585) );
  OAI22_X1 U1220 ( .A1(n47), .A2(n716), .B1(n45), .B2(n715), .ZN(n587) );
  OAI22_X1 U1221 ( .A1(n11), .A2(n807), .B1(n10), .B2(n806), .ZN(n672) );
  XNOR2_X1 U1222 ( .A(n643), .B(n601), .ZN(n443) );
  OAI22_X1 U1223 ( .A1(n35), .A2(n738), .B1(n34), .B2(n737), .ZN(n607) );
  OAI22_X1 U1224 ( .A1(n6), .A2(n828), .B1(n827), .B2(n4), .ZN(n693) );
  OAI22_X1 U1225 ( .A1(n6), .A2(n823), .B1(n822), .B2(n4), .ZN(n688) );
  OAI22_X1 U1226 ( .A1(n36), .A2(n748), .B1(n33), .B2(n747), .ZN(n617) );
  AND2_X1 U1227 ( .A1(n1045), .A2(n543), .ZN(n589) );
  OAI22_X1 U1228 ( .A1(n6), .A2(n827), .B1(n826), .B2(n4), .ZN(n692) );
  AND2_X1 U1229 ( .A1(n1015), .A2(n549), .ZN(n621) );
  OAI22_X1 U1230 ( .A1(n24), .A2(n782), .B1(n21), .B2(n781), .ZN(n649) );
  OAI22_X1 U1231 ( .A1(n18), .A2(n790), .B1(n16), .B2(n789), .ZN(n656) );
  OAI22_X1 U1232 ( .A1(n47), .A2(n715), .B1(n45), .B2(n714), .ZN(n586) );
  OAI22_X1 U1233 ( .A1(n11), .A2(n815), .B1(n9), .B2(n814), .ZN(n680) );
  OAI22_X1 U1234 ( .A1(n5), .A2(n830), .B1(n829), .B2(n3), .ZN(n695) );
  OAI22_X1 U1235 ( .A1(n5), .A2(n831), .B1(n830), .B2(n3), .ZN(n696) );
  OAI22_X1 U1236 ( .A1(n11), .A2(n816), .B1(n9), .B2(n815), .ZN(n681) );
  AND2_X1 U1237 ( .A1(n1045), .A2(n555), .ZN(n653) );
  OAI22_X1 U1238 ( .A1(n30), .A2(n763), .B1(n27), .B2(n762), .ZN(n631) );
  OAI22_X1 U1239 ( .A1(n11), .A2(n808), .B1(n10), .B2(n807), .ZN(n673) );
  OAI22_X1 U1240 ( .A1(n42), .A2(n733), .B1(n39), .B2(n732), .ZN(n603) );
  OAI22_X1 U1241 ( .A1(n18), .A2(n792), .B1(n16), .B2(n791), .ZN(n658) );
  OAI22_X1 U1242 ( .A1(n30), .A2(n762), .B1(n761), .B2(n27), .ZN(n630) );
  OAI22_X1 U1243 ( .A1(n6), .A2(n822), .B1(n821), .B2(n4), .ZN(n687) );
  OAI22_X1 U1244 ( .A1(n35), .A2(n741), .B1(n34), .B2(n740), .ZN(n610) );
  INV_X1 U1245 ( .A(n380), .ZN(n381) );
  OAI22_X1 U1246 ( .A1(n11), .A2(n811), .B1(n10), .B2(n810), .ZN(n676) );
  OAI22_X1 U1247 ( .A1(n24), .A2(n781), .B1(n21), .B2(n780), .ZN(n648) );
  OAI22_X1 U1248 ( .A1(n6), .A2(n826), .B1(n825), .B2(n4), .ZN(n691) );
  OAI22_X1 U1249 ( .A1(n766), .A2(n29), .B1(n765), .B2(n28), .ZN(n634) );
  OAI22_X1 U1250 ( .A1(n35), .A2(n739), .B1(n34), .B2(n738), .ZN(n608) );
  OAI22_X1 U1251 ( .A1(n48), .A2(n709), .B1(n46), .B2(n708), .ZN(n580) );
  OAI22_X1 U1252 ( .A1(n5), .A2(n829), .B1(n828), .B2(n3), .ZN(n694) );
  AND2_X1 U1253 ( .A1(n1058), .A2(n552), .ZN(n637) );
  NAND2_X1 U1254 ( .A1(n539), .A2(n540), .ZN(n291) );
  OAI22_X1 U1255 ( .A1(n42), .A2(n879), .B1(n735), .B2(n39), .ZN(n567) );
  OAI22_X1 U1256 ( .A1(n734), .A2(n42), .B1(n39), .B2(n733), .ZN(n604) );
  OR2_X1 U1257 ( .A1(n1058), .A2(n879), .ZN(n735) );
  INV_X1 U1258 ( .A(n542), .ZN(n574) );
  AOI21_X1 U1259 ( .B1(n48), .B2(n46), .A(n702), .ZN(n542) );
  AND2_X1 U1260 ( .A1(n1015), .A2(n564), .ZN(product[0]) );
  INV_X1 U1261 ( .A(n3), .ZN(n564) );
  OR2_X1 U1262 ( .A1(n1058), .A2(n880), .ZN(n752) );
  OR2_X1 U1263 ( .A1(n1045), .A2(n883), .ZN(n803) );
  OR2_X1 U1264 ( .A1(n1058), .A2(n882), .ZN(n786) );
  OR2_X1 U1265 ( .A1(n1057), .A2(n881), .ZN(n769) );
  INV_X1 U1266 ( .A(n15), .ZN(n558) );
  INV_X1 U1267 ( .A(n21), .ZN(n555) );
  INV_X1 U1268 ( .A(n45), .ZN(n543) );
  INV_X1 U1269 ( .A(n33), .ZN(n549) );
  INV_X1 U1270 ( .A(n27), .ZN(n552) );
  INV_X1 U1271 ( .A(n39), .ZN(n546) );
  OAI22_X1 U1272 ( .A1(n1028), .A2(n771), .B1(n22), .B2(n770), .ZN(n380) );
  BUF_X1 U1273 ( .A(n877), .Z(n3) );
  OAI22_X1 U1274 ( .A1(n1028), .A2(n776), .B1(n22), .B2(n775), .ZN(n643) );
  OAI22_X1 U1275 ( .A1(n6), .A2(n885), .B1(n837), .B2(n4), .ZN(n573) );
  OR2_X1 U1276 ( .A1(n1058), .A2(n885), .ZN(n837) );
  INV_X1 U1277 ( .A(n1), .ZN(n885) );
  OAI22_X1 U1278 ( .A1(n5), .A2(n836), .B1(n835), .B2(n3), .ZN(n701) );
  OAI22_X1 U1279 ( .A1(n30), .A2(n768), .B1(n27), .B2(n767), .ZN(n636) );
  OAI22_X1 U1280 ( .A1(n5), .A2(n834), .B1(n833), .B2(n3), .ZN(n699) );
  OAI22_X1 U1281 ( .A1(n11), .A2(n819), .B1(n9), .B2(n818), .ZN(n684) );
  OAI22_X1 U1282 ( .A1(n35), .A2(n747), .B1(n33), .B2(n746), .ZN(n616) );
  OAI22_X1 U1283 ( .A1(n1028), .A2(n777), .B1(n22), .B2(n776), .ZN(n644) );
  OAI22_X1 U1284 ( .A1(n42), .A2(n732), .B1(n39), .B2(n731), .ZN(n602) );
  BUF_X1 U1285 ( .A(n877), .Z(n4) );
  CLKBUF_X3 U1286 ( .A(n863), .Z(n42) );
  OAI22_X1 U1287 ( .A1(n1047), .A2(n883), .B1(n803), .B2(n16), .ZN(n571) );
  OAI22_X1 U1288 ( .A1(n36), .A2(n751), .B1(n33), .B2(n750), .ZN(n620) );
  OAI22_X1 U1289 ( .A1(n36), .A2(n880), .B1(n752), .B2(n34), .ZN(n568) );
  BUF_X1 U1290 ( .A(n869), .Z(n5) );
  BUF_X2 U1291 ( .A(n862), .Z(n47) );
  BUF_X2 U1292 ( .A(n10), .Z(n9) );
  BUF_X1 U1293 ( .A(n870), .Z(n45) );
  BUF_X2 U1294 ( .A(b[14]), .Z(n839) );
  BUF_X2 U1295 ( .A(n875), .Z(n15) );
  BUF_X1 U1296 ( .A(n870), .Z(n46) );
  BUF_X2 U1297 ( .A(n862), .Z(n48) );
  BUF_X2 U1298 ( .A(n876), .Z(n10) );
  OAI22_X1 U1299 ( .A1(n1028), .A2(n774), .B1(n22), .B2(n773), .ZN(n641) );
  OAI22_X1 U1300 ( .A1(n35), .A2(n742), .B1(n34), .B2(n741), .ZN(n611) );
  OAI22_X1 U1301 ( .A1(n1028), .A2(n775), .B1(n22), .B2(n774), .ZN(n642) );
  INV_X1 U1302 ( .A(n13), .ZN(n883) );
  BUF_X1 U1303 ( .A(n863), .Z(n41) );
  OAI22_X1 U1304 ( .A1(n24), .A2(n785), .B1(n21), .B2(n784), .ZN(n652) );
  OAI22_X1 U1305 ( .A1(n1028), .A2(n882), .B1(n786), .B2(n22), .ZN(n570) );
  OAI22_X1 U1306 ( .A1(n11), .A2(n884), .B1(n820), .B2(n10), .ZN(n572) );
  OR2_X1 U1307 ( .A1(n1058), .A2(n884), .ZN(n820) );
  INV_X1 U1308 ( .A(n7), .ZN(n884) );
  INV_X1 U1309 ( .A(n37), .ZN(n879) );
  INV_X1 U1310 ( .A(n31), .ZN(n880) );
  INV_X1 U1311 ( .A(n1030), .ZN(n881) );
  INV_X1 U1312 ( .A(n19), .ZN(n882) );
  XNOR2_X1 U1313 ( .A(a[10]), .B(a[9]), .ZN(n872) );
  XNOR2_X1 U1314 ( .A(a[14]), .B(a[13]), .ZN(n870) );
  XNOR2_X1 U1315 ( .A(a[12]), .B(a[11]), .ZN(n871) );
  XNOR2_X1 U1316 ( .A(a[7]), .B(a[8]), .ZN(n873) );
  BUF_X4 U1317 ( .A(a[7]), .Z(n19) );
  INV_X1 U1318 ( .A(a[0]), .ZN(n877) );
  OAI21_X1 U1319 ( .B1(n219), .B2(n1026), .A(n212), .ZN(n210) );
  NOR2_X1 U1320 ( .A1(n218), .A2(n211), .ZN(n209) );
  NOR2_X1 U1321 ( .A1(n405), .A2(n416), .ZN(n211) );
  XOR2_X1 U1322 ( .A(n1014), .B(n76), .Z(product[8]) );
  OAI21_X1 U1323 ( .B1(n276), .B2(n274), .A(n275), .ZN(n273) );
  INV_X1 U1324 ( .A(n235), .ZN(n234) );
  OAI22_X1 U1325 ( .A1(n35), .A2(n737), .B1(n34), .B2(n736), .ZN(n348) );
  INV_X1 U1326 ( .A(n348), .ZN(n349) );
  NAND2_X1 U1327 ( .A1(n209), .A2(n225), .ZN(n207) );
  NOR2_X1 U1328 ( .A1(n227), .A2(n232), .ZN(n225) );
  OAI22_X1 U1329 ( .A1(n1047), .A2(n801), .B1(n15), .B2(n800), .ZN(n667) );
  OAI22_X1 U1330 ( .A1(n967), .A2(n795), .B1(n15), .B2(n794), .ZN(n661) );
  OAI22_X1 U1331 ( .A1(n1047), .A2(n799), .B1(n15), .B2(n798), .ZN(n665) );
  OAI22_X1 U1332 ( .A1(n18), .A2(n800), .B1(n15), .B2(n799), .ZN(n666) );
  OAI22_X1 U1333 ( .A1(n18), .A2(n797), .B1(n15), .B2(n796), .ZN(n663) );
  OAI22_X1 U1334 ( .A1(n18), .A2(n798), .B1(n15), .B2(n797), .ZN(n664) );
  OAI22_X1 U1335 ( .A1(n18), .A2(n802), .B1(n15), .B2(n801), .ZN(n668) );
  OAI22_X1 U1336 ( .A1(n796), .A2(n17), .B1(n15), .B2(n795), .ZN(n662) );
  INV_X1 U1337 ( .A(n965), .ZN(n254) );
  AOI21_X1 U1338 ( .B1(n255), .B2(n236), .A(n237), .ZN(n235) );
  XNOR2_X1 U1339 ( .A(n966), .B(n77), .ZN(product[7]) );
  INV_X1 U1340 ( .A(n150), .ZN(n148) );
  OAI21_X1 U1341 ( .B1(n150), .B2(n133), .A(n134), .ZN(n132) );
  OAI21_X1 U1342 ( .B1(n150), .B2(n144), .A(n145), .ZN(n141) );
  OAI21_X1 U1343 ( .B1(n150), .B2(n124), .A(n125), .ZN(n119) );
  OAI21_X1 U1344 ( .B1(n954), .B2(n96), .A(n97), .ZN(n95) );
  OAI21_X1 U1345 ( .B1(n150), .B2(n109), .A(n110), .ZN(n108) );
  OAI22_X1 U1346 ( .A1(n42), .A2(n724), .B1(n40), .B2(n723), .ZN(n594) );
  OAI22_X1 U1347 ( .A1(n41), .A2(n725), .B1(n40), .B2(n724), .ZN(n595) );
  OAI22_X1 U1348 ( .A1(n1028), .A2(n772), .B1(n22), .B2(n771), .ZN(n639) );
  NAND2_X1 U1349 ( .A1(n857), .A2(n873), .ZN(n865) );
  XNOR2_X1 U1350 ( .A(a[6]), .B(a[5]), .ZN(n874) );
  OAI22_X1 U1351 ( .A1(n41), .A2(n729), .B1(n39), .B2(n728), .ZN(n599) );
  OAI22_X1 U1352 ( .A1(n41), .A2(n730), .B1(n39), .B2(n729), .ZN(n600) );
  OAI22_X1 U1353 ( .A1(n42), .A2(n727), .B1(n39), .B2(n726), .ZN(n597) );
  OAI22_X1 U1354 ( .A1(n41), .A2(n728), .B1(n39), .B2(n727), .ZN(n598) );
  AND2_X1 U1355 ( .A1(n365), .A2(n372), .ZN(n1056) );
  NAND2_X1 U1356 ( .A1(n856), .A2(n872), .ZN(n864) );
  INV_X1 U1357 ( .A(n554), .ZN(n638) );
  AOI21_X1 U1358 ( .B1(n1028), .B2(n22), .A(n770), .ZN(n554) );
  INV_X1 U1359 ( .A(n402), .ZN(n403) );
  BUF_X2 U1360 ( .A(n867), .Z(n18) );
  XOR2_X1 U1361 ( .A(n80), .B(n292), .Z(product[4]) );
  XOR2_X1 U1362 ( .A(n78), .B(n1022), .Z(product[6]) );
  XNOR2_X1 U1363 ( .A(n7), .B(n848), .ZN(n814) );
  XNOR2_X1 U1364 ( .A(n7), .B(n842), .ZN(n808) );
  XNOR2_X1 U1365 ( .A(n1016), .B(n988), .ZN(n813) );
  XNOR2_X1 U1366 ( .A(n7), .B(n841), .ZN(n807) );
  XNOR2_X1 U1367 ( .A(n7), .B(n844), .ZN(n810) );
  XNOR2_X1 U1368 ( .A(n7), .B(n843), .ZN(n809) );
  XNOR2_X1 U1369 ( .A(n1016), .B(n1038), .ZN(n812) );
  XNOR2_X1 U1370 ( .A(n7), .B(n845), .ZN(n811) );
  XNOR2_X1 U1371 ( .A(n7), .B(n851), .ZN(n817) );
  XNOR2_X1 U1372 ( .A(n7), .B(n1045), .ZN(n819) );
  XNOR2_X1 U1373 ( .A(n7), .B(n850), .ZN(n816) );
  XNOR2_X1 U1374 ( .A(n7), .B(n849), .ZN(n815) );
  XNOR2_X1 U1375 ( .A(n7), .B(n852), .ZN(n818) );
  XNOR2_X1 U1376 ( .A(n7), .B(n840), .ZN(n806) );
  XNOR2_X1 U1377 ( .A(n43), .B(n988), .ZN(n711) );
  XNOR2_X1 U1378 ( .A(n43), .B(n849), .ZN(n713) );
  XNOR2_X1 U1379 ( .A(n43), .B(n850), .ZN(n714) );
  XNOR2_X1 U1380 ( .A(n43), .B(n851), .ZN(n715) );
  XNOR2_X1 U1381 ( .A(n43), .B(n852), .ZN(n716) );
  XNOR2_X1 U1382 ( .A(n43), .B(n1057), .ZN(n717) );
  INV_X1 U1383 ( .A(n43), .ZN(n878) );
  XNOR2_X1 U1384 ( .A(n43), .B(n1038), .ZN(n710) );
  XNOR2_X1 U1385 ( .A(n43), .B(n845), .ZN(n709) );
  XNOR2_X1 U1386 ( .A(n43), .B(n844), .ZN(n708) );
  XNOR2_X1 U1387 ( .A(n43), .B(n843), .ZN(n707) );
  XNOR2_X1 U1388 ( .A(n43), .B(n842), .ZN(n706) );
  XNOR2_X1 U1389 ( .A(n43), .B(n841), .ZN(n705) );
  XNOR2_X1 U1390 ( .A(n43), .B(n840), .ZN(n704) );
  XNOR2_X1 U1391 ( .A(n43), .B(n848), .ZN(n712) );
  XNOR2_X1 U1392 ( .A(n43), .B(n1035), .ZN(n703) );
  XNOR2_X1 U1393 ( .A(n7), .B(n839), .ZN(n805) );
  INV_X1 U1394 ( .A(n563), .ZN(n686) );
  AOI21_X1 U1395 ( .B1(n6), .B2(n4), .A(n821), .ZN(n563) );
  OAI22_X1 U1396 ( .A1(n1047), .A2(n789), .B1(n16), .B2(n788), .ZN(n655) );
  XNOR2_X1 U1397 ( .A(n43), .B(n1021), .ZN(n702) );
  XNOR2_X1 U1398 ( .A(n7), .B(n838), .ZN(n804) );
  AOI21_X1 U1399 ( .B1(n967), .B2(n16), .A(n787), .ZN(n557) );
  NAND2_X1 U1400 ( .A1(n854), .A2(n870), .ZN(n862) );
  XNOR2_X1 U1401 ( .A(n19), .B(n1058), .ZN(n785) );
  XNOR2_X1 U1402 ( .A(n19), .B(n852), .ZN(n784) );
  XNOR2_X1 U1403 ( .A(n19), .B(n848), .ZN(n780) );
  XNOR2_X1 U1404 ( .A(n19), .B(n1038), .ZN(n778) );
  XNOR2_X1 U1405 ( .A(n847), .B(n19), .ZN(n779) );
  XNOR2_X1 U1406 ( .A(n19), .B(n851), .ZN(n783) );
  XNOR2_X1 U1407 ( .A(n19), .B(n850), .ZN(n782) );
  XNOR2_X1 U1408 ( .A(n19), .B(n849), .ZN(n781) );
  XNOR2_X1 U1409 ( .A(n19), .B(n845), .ZN(n777) );
  XNOR2_X1 U1410 ( .A(n19), .B(n844), .ZN(n776) );
  XNOR2_X1 U1411 ( .A(n19), .B(n843), .ZN(n775) );
  XNOR2_X1 U1412 ( .A(n19), .B(n842), .ZN(n774) );
  XNOR2_X1 U1413 ( .A(n19), .B(n839), .ZN(n771) );
  XNOR2_X1 U1414 ( .A(n19), .B(n841), .ZN(n773) );
  XNOR2_X1 U1415 ( .A(n19), .B(n840), .ZN(n772) );
  XNOR2_X1 U1416 ( .A(n19), .B(n1021), .ZN(n770) );
  INV_X1 U1417 ( .A(n232), .ZN(n317) );
  XNOR2_X1 U1418 ( .A(n1030), .B(n1058), .ZN(n768) );
  XNOR2_X1 U1419 ( .A(n1030), .B(n848), .ZN(n763) );
  XNOR2_X1 U1420 ( .A(n1030), .B(n849), .ZN(n764) );
  XNOR2_X1 U1421 ( .A(n1030), .B(n852), .ZN(n767) );
  XNOR2_X1 U1422 ( .A(n25), .B(n851), .ZN(n766) );
  XNOR2_X1 U1423 ( .A(n850), .B(n25), .ZN(n765) );
  XNOR2_X1 U1424 ( .A(n1030), .B(n847), .ZN(n762) );
  XNOR2_X1 U1425 ( .A(n1030), .B(n1038), .ZN(n761) );
  XNOR2_X1 U1426 ( .A(n1030), .B(n1021), .ZN(n753) );
  XNOR2_X1 U1427 ( .A(n1030), .B(n841), .ZN(n756) );
  XNOR2_X1 U1428 ( .A(n1030), .B(n839), .ZN(n754) );
  XNOR2_X1 U1429 ( .A(n1030), .B(n840), .ZN(n755) );
  XNOR2_X1 U1430 ( .A(n1030), .B(n845), .ZN(n760) );
  XNOR2_X1 U1431 ( .A(n25), .B(n844), .ZN(n759) );
  XNOR2_X1 U1432 ( .A(n1030), .B(n843), .ZN(n758) );
  XNOR2_X1 U1433 ( .A(n1030), .B(n842), .ZN(n757) );
  OAI22_X1 U1434 ( .A1(n761), .A2(n29), .B1(n27), .B2(n760), .ZN(n629) );
  NOR2_X1 U1435 ( .A1(n241), .A2(n964), .ZN(n236) );
  OAI21_X1 U1436 ( .B1(n242), .B2(n238), .A(n239), .ZN(n237) );
  XNOR2_X1 U1437 ( .A(n37), .B(n840), .ZN(n721) );
  XNOR2_X1 U1438 ( .A(n37), .B(n1035), .ZN(n720) );
  XNOR2_X1 U1439 ( .A(n37), .B(n1021), .ZN(n719) );
  XNOR2_X1 U1440 ( .A(n37), .B(n841), .ZN(n722) );
  XNOR2_X1 U1441 ( .A(n37), .B(n1057), .ZN(n734) );
  XNOR2_X1 U1442 ( .A(n37), .B(n852), .ZN(n733) );
  XNOR2_X1 U1443 ( .A(n37), .B(n851), .ZN(n732) );
  XNOR2_X1 U1444 ( .A(n37), .B(n842), .ZN(n723) );
  XNOR2_X1 U1445 ( .A(n37), .B(n850), .ZN(n731) );
  XNOR2_X1 U1446 ( .A(n37), .B(n849), .ZN(n730) );
  XNOR2_X1 U1447 ( .A(n37), .B(n845), .ZN(n726) );
  XNOR2_X1 U1448 ( .A(n37), .B(n844), .ZN(n725) );
  XNOR2_X1 U1449 ( .A(n37), .B(n843), .ZN(n724) );
  XNOR2_X1 U1450 ( .A(n37), .B(n848), .ZN(n729) );
  XNOR2_X1 U1451 ( .A(n37), .B(n847), .ZN(n728) );
  XNOR2_X1 U1452 ( .A(n37), .B(n1038), .ZN(n727) );
  BUF_X2 U1453 ( .A(n864), .Z(n35) );
  OAI22_X1 U1454 ( .A1(n35), .A2(n745), .B1(n744), .B2(n33), .ZN(n614) );
  AOI21_X1 U1455 ( .B1(n226), .B2(n1025), .A(n210), .ZN(n208) );
  OAI21_X1 U1456 ( .B1(n1032), .B2(n233), .A(n228), .ZN(n226) );
  XNOR2_X1 U1457 ( .A(a[2]), .B(a[1]), .ZN(n876) );
  BUF_X2 U1458 ( .A(n868), .Z(n11) );
  NAND2_X1 U1459 ( .A1(n860), .A2(n876), .ZN(n868) );
  OAI22_X1 U1460 ( .A1(n47), .A2(n713), .B1(n45), .B2(n712), .ZN(n584) );
  XNOR2_X1 U1461 ( .A(n1011), .B(n849), .ZN(n747) );
  XNOR2_X1 U1462 ( .A(n1011), .B(n840), .ZN(n738) );
  XNOR2_X1 U1463 ( .A(n1011), .B(n851), .ZN(n749) );
  XNOR2_X1 U1464 ( .A(n1011), .B(n843), .ZN(n741) );
  XNOR2_X1 U1465 ( .A(n1011), .B(n1057), .ZN(n751) );
  XNOR2_X1 U1466 ( .A(n1011), .B(n850), .ZN(n748) );
  XNOR2_X1 U1467 ( .A(n1011), .B(n852), .ZN(n750) );
  XNOR2_X1 U1468 ( .A(n1011), .B(n1035), .ZN(n737) );
  XNOR2_X1 U1469 ( .A(n1011), .B(n1021), .ZN(n736) );
  XNOR2_X1 U1470 ( .A(n31), .B(n848), .ZN(n746) );
  XNOR2_X1 U1471 ( .A(n1011), .B(n842), .ZN(n740) );
  XNOR2_X1 U1472 ( .A(n847), .B(n31), .ZN(n745) );
  XNOR2_X1 U1473 ( .A(n1011), .B(n1038), .ZN(n744) );
  XNOR2_X1 U1474 ( .A(n1011), .B(n841), .ZN(n739) );
  XNOR2_X1 U1475 ( .A(n1011), .B(n845), .ZN(n743) );
  XNOR2_X1 U1476 ( .A(n31), .B(n844), .ZN(n742) );
  XNOR2_X1 U1477 ( .A(n1), .B(n845), .ZN(n828) );
  XNOR2_X1 U1478 ( .A(n1), .B(n1038), .ZN(n829) );
  XNOR2_X1 U1479 ( .A(n1), .B(n844), .ZN(n827) );
  XNOR2_X1 U1480 ( .A(n1), .B(n849), .ZN(n832) );
  XNOR2_X1 U1481 ( .A(n1), .B(n839), .ZN(n822) );
  XNOR2_X1 U1482 ( .A(n1), .B(n848), .ZN(n831) );
  XNOR2_X1 U1483 ( .A(n1), .B(n1045), .ZN(n836) );
  XNOR2_X1 U1484 ( .A(n1), .B(n847), .ZN(n830) );
  XNOR2_X1 U1485 ( .A(n1), .B(n841), .ZN(n824) );
  XNOR2_X1 U1486 ( .A(n1), .B(n850), .ZN(n833) );
  XNOR2_X1 U1487 ( .A(n1), .B(n840), .ZN(n823) );
  XNOR2_X1 U1488 ( .A(n1), .B(n852), .ZN(n835) );
  XNOR2_X1 U1489 ( .A(n1), .B(n851), .ZN(n834) );
  XNOR2_X1 U1490 ( .A(n1), .B(n842), .ZN(n825) );
  XNOR2_X1 U1491 ( .A(n1), .B(n843), .ZN(n826) );
  XNOR2_X1 U1492 ( .A(n1), .B(n838), .ZN(n821) );
  OAI22_X1 U1493 ( .A1(n36), .A2(n743), .B1(n34), .B2(n742), .ZN(n612) );
  BUF_X2 U1494 ( .A(n864), .Z(n36) );
  NAND2_X1 U1495 ( .A1(n858), .A2(n874), .ZN(n866) );
  AOI21_X1 U1496 ( .B1(n12), .B2(n10), .A(n804), .ZN(n560) );
  INV_X1 U1497 ( .A(n560), .ZN(n670) );
  NAND2_X1 U1498 ( .A1(n365), .A2(n372), .ZN(n182) );
  OAI22_X1 U1499 ( .A1(n24), .A2(n773), .B1(n22), .B2(n772), .ZN(n640) );
  OAI21_X1 U1500 ( .B1(n268), .B2(n256), .A(n257), .ZN(n255) );
  XNOR2_X1 U1501 ( .A(n974), .B(n848), .ZN(n797) );
  XNOR2_X1 U1502 ( .A(n974), .B(n849), .ZN(n798) );
  XNOR2_X1 U1503 ( .A(n974), .B(n843), .ZN(n792) );
  XNOR2_X1 U1504 ( .A(n974), .B(n851), .ZN(n800) );
  XNOR2_X1 U1505 ( .A(n974), .B(n850), .ZN(n799) );
  XNOR2_X1 U1506 ( .A(n974), .B(n845), .ZN(n794) );
  XNOR2_X1 U1507 ( .A(n974), .B(n844), .ZN(n793) );
  XNOR2_X1 U1508 ( .A(n13), .B(n842), .ZN(n791) );
  XNOR2_X1 U1509 ( .A(n847), .B(n13), .ZN(n796) );
  XNOR2_X1 U1510 ( .A(n13), .B(n1037), .ZN(n795) );
  XNOR2_X1 U1511 ( .A(n13), .B(n841), .ZN(n790) );
  XNOR2_X1 U1512 ( .A(n974), .B(n1057), .ZN(n802) );
  XNOR2_X1 U1513 ( .A(n974), .B(n852), .ZN(n801) );
  XNOR2_X1 U1514 ( .A(n974), .B(n840), .ZN(n789) );
  XNOR2_X1 U1515 ( .A(n974), .B(n839), .ZN(n788) );
  XNOR2_X1 U1516 ( .A(n974), .B(n838), .ZN(n787) );
  NAND2_X1 U1517 ( .A1(n861), .A2(n877), .ZN(n869) );
  BUF_X2 U1518 ( .A(n869), .Z(n6) );
  AOI21_X1 U1519 ( .B1(n234), .B2(n317), .A(n231), .ZN(n229) );
  INV_X1 U1520 ( .A(n362), .ZN(n363) );
  OAI22_X1 U1521 ( .A1(n30), .A2(n881), .B1(n769), .B2(n27), .ZN(n569) );
  AOI21_X1 U1522 ( .B1(n30), .B2(n27), .A(n753), .ZN(n551) );
  OAI22_X1 U1523 ( .A1(n30), .A2(n759), .B1(n27), .B2(n758), .ZN(n627) );
  OAI22_X1 U1524 ( .A1(n30), .A2(n757), .B1(n27), .B2(n756), .ZN(n625) );
  OAI22_X1 U1525 ( .A1(n30), .A2(n756), .B1(n27), .B2(n755), .ZN(n624) );
  OAI22_X1 U1526 ( .A1(n30), .A2(n755), .B1(n27), .B2(n754), .ZN(n623) );
  OAI22_X1 U1527 ( .A1(n29), .A2(n760), .B1(n28), .B2(n759), .ZN(n628) );
  OAI22_X1 U1528 ( .A1(n29), .A2(n758), .B1(n28), .B2(n757), .ZN(n626) );
  NAND2_X1 U1529 ( .A1(n859), .A2(n875), .ZN(n867) );
  NAND2_X1 U1530 ( .A1(n197), .A2(n151), .ZN(n149) );
  NAND2_X1 U1531 ( .A1(n855), .A2(n871), .ZN(n863) );
  XNOR2_X1 U1532 ( .A(n79), .B(n289), .ZN(product[5]) );
  XNOR2_X1 U1533 ( .A(n273), .B(n75), .ZN(product[9]) );
  BUF_X4 U1534 ( .A(a[15]), .Z(n43) );
  NOR2_X1 U1535 ( .A1(n204), .A2(n199), .ZN(n197) );
  OAI21_X1 U1536 ( .B1(n199), .B2(n205), .A(n200), .ZN(n198) );
  INV_X1 U1537 ( .A(n199), .ZN(n312) );
  NOR2_X1 U1538 ( .A1(n383), .A2(n392), .ZN(n199) );
  AOI21_X1 U1539 ( .B1(n1020), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U1540 ( .B1(n1036), .B2(n94), .A(n95), .ZN(n93) );
  AOI21_X1 U1541 ( .B1(n1031), .B2(n118), .A(n119), .ZN(n117) );
  AOI21_X1 U1542 ( .B1(n1036), .B2(n107), .A(n108), .ZN(n106) );
  AOI21_X1 U1543 ( .B1(n1031), .B2(n131), .A(n132), .ZN(n130) );
  AOI21_X1 U1544 ( .B1(n1036), .B2(n140), .A(n141), .ZN(n139) );
  AOI21_X1 U1545 ( .B1(n51), .B2(n184), .A(n185), .ZN(n183) );
  XNOR2_X1 U1546 ( .A(n1031), .B(n65), .ZN(product[19]) );
  AOI21_X1 U1547 ( .B1(n51), .B2(n171), .A(n172), .ZN(n170) );
  AOI21_X1 U1548 ( .B1(n1036), .B2(n313), .A(n203), .ZN(n201) );
  AOI21_X1 U1549 ( .B1(n1036), .B2(n147), .A(n148), .ZN(n146) );
  AOI21_X1 U1550 ( .B1(n51), .B2(n197), .A(n194), .ZN(n192) );
  OAI21_X1 U1551 ( .B1(n157), .B2(n169), .A(n158), .ZN(n156) );
  NOR2_X1 U1552 ( .A1(n168), .A2(n157), .ZN(n155) );
  NAND2_X1 U1553 ( .A1(n351), .A2(n356), .ZN(n158) );
  XOR2_X1 U1554 ( .A(a[7]), .B(a[6]), .Z(n858) );
  BUF_X4 U1555 ( .A(a[13]), .Z(n37) );
  XOR2_X1 U1556 ( .A(a[12]), .B(a[13]), .Z(n855) );
  XOR2_X1 U1557 ( .A(a[8]), .B(a[9]), .Z(n857) );
  AOI21_X1 U1558 ( .B1(n155), .B2(n1056), .A(n156), .ZN(n154) );
  NOR2_X1 U1559 ( .A1(n190), .A2(n153), .ZN(n151) );
  NAND2_X1 U1560 ( .A1(n155), .A2(n1003), .ZN(n153) );
  OAI21_X1 U1561 ( .B1(n235), .B2(n207), .A(n208), .ZN(n206) );
  XOR2_X1 U1562 ( .A(a[10]), .B(a[11]), .Z(n856) );
  AOI21_X1 U1563 ( .B1(n1036), .B2(n160), .A(n161), .ZN(n159) );
  OAI21_X1 U1564 ( .B1(n153), .B2(n191), .A(n154), .ZN(n152) );
  BUF_X2 U1565 ( .A(n865), .Z(n30) );
  NAND2_X1 U1566 ( .A1(n980), .A2(n296), .ZN(n81) );
  XOR2_X1 U1567 ( .A(a[2]), .B(a[3]), .Z(n860) );
  XNOR2_X1 U1568 ( .A(a[4]), .B(a[3]), .ZN(n875) );
  NAND2_X1 U1569 ( .A1(n541), .A2(n572), .ZN(n296) );
  XOR2_X1 U1570 ( .A(a[4]), .B(a[5]), .Z(n859) );
  XOR2_X1 U1571 ( .A(a[0]), .B(a[1]), .Z(n861) );
endmodule


module datapath_DW_mult_tc_10 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n4, n5, n6, n7, n10, n11, n12, n13, n15, n16, n17, n18, n19, n21,
         n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34, n35, n36, n37,
         n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n51, n54, n55, n56,
         n59, n60, n65, n66, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n84, n85, n86, n87, n88, n90, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n103, n105, n106, n107, n108,
         n109, n110, n114, n116, n117, n118, n119, n122, n123, n124, n125,
         n127, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n143, n144, n145, n146, n147, n148, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n180, n182, n183, n184, n185, n188,
         n189, n190, n191, n192, n193, n195, n196, n197, n198, n199, n200,
         n201, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n217, n218, n219, n220, n222, n223, n224, n225,
         n226, n227, n228, n229, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n244, n246, n247, n248, n253, n254,
         n255, n256, n257, n259, n261, n262, n264, n266, n267, n268, n270,
         n272, n273, n274, n275, n276, n278, n280, n281, n282, n283, n284,
         n286, n288, n289, n290, n291, n292, n294, n296, n297, n298, n299,
         n301, n306, n308, n312, n313, n314, n316, n317, n324, n326, n328,
         n330, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n545, n546, n548, n549, n551, n552, n554,
         n555, n557, n558, n560, n561, n563, n564, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1064, n1065;
  assign product[31] = n84;

  FA_X1 U364 ( .A(n575), .B(n338), .CI(n590), .CO(n334), .S(n335) );
  FA_X1 U365 ( .A(n339), .B(n576), .CI(n342), .CO(n336), .S(n337) );
  FA_X1 U367 ( .A(n346), .B(n577), .CI(n343), .CO(n340), .S(n341) );
  FA_X1 U368 ( .A(n591), .B(n348), .CI(n606), .CO(n342), .S(n343) );
  FA_X1 U369 ( .A(n347), .B(n354), .CI(n352), .CO(n344), .S(n345) );
  FA_X1 U370 ( .A(n578), .B(n592), .CI(n349), .CO(n346), .S(n347) );
  FA_X1 U372 ( .A(n358), .B(n355), .CI(n353), .CO(n350), .S(n351) );
  FA_X1 U373 ( .A(n362), .B(n607), .CI(n360), .CO(n352), .S(n353) );
  FA_X1 U374 ( .A(n593), .B(n579), .CI(n622), .CO(n354), .S(n355) );
  FA_X1 U375 ( .A(n359), .B(n361), .CI(n366), .CO(n356), .S(n357) );
  FA_X1 U376 ( .A(n370), .B(n363), .CI(n368), .CO(n358), .S(n359) );
  FA_X1 U377 ( .A(n580), .B(n594), .CI(n608), .CO(n360), .S(n361) );
  FA_X1 U379 ( .A(n374), .B(n376), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U380 ( .A(n369), .B(n378), .CI(n371), .CO(n366), .S(n367) );
  FA_X1 U381 ( .A(n595), .B(n380), .CI(n609), .CO(n368), .S(n369) );
  FA_X1 U382 ( .A(n623), .B(n581), .CI(n638), .CO(n370), .S(n371) );
  FA_X1 U383 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  FA_X1 U385 ( .A(n381), .B(n610), .CI(n390), .CO(n376), .S(n377) );
  FA_X1 U386 ( .A(n624), .B(n596), .CI(n582), .CO(n378), .S(n379) );
  FA_X1 U388 ( .A(n394), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U389 ( .A(n391), .B(n389), .CI(n396), .CO(n384), .S(n385) );
  FA_X1 U390 ( .A(n400), .B(n625), .CI(n398), .CO(n386), .S(n387) );
  FA_X1 U391 ( .A(n597), .B(n639), .CI(n611), .CO(n388), .S(n389) );
  FA_X1 U392 ( .A(n1040), .B(n583), .CI(n654), .CO(n390), .S(n391) );
  FA_X1 U393 ( .A(n406), .B(n397), .CI(n395), .CO(n392), .S(n393) );
  FA_X1 U394 ( .A(n410), .B(n399), .CI(n408), .CO(n394), .S(n395) );
  FA_X1 U395 ( .A(n412), .B(n414), .CI(n401), .CO(n396), .S(n397) );
  FA_X1 U396 ( .A(n584), .B(n598), .CI(n403), .CO(n398), .S(n399) );
  FA_X1 U397 ( .A(n640), .B(n626), .CI(n612), .CO(n400), .S(n401) );
  FA_X1 U399 ( .A(n418), .B(n409), .CI(n407), .CO(n404), .S(n405) );
  FA_X1 U400 ( .A(n411), .B(n422), .CI(n420), .CO(n406), .S(n407) );
  FA_X1 U401 ( .A(n413), .B(n424), .CI(n415), .CO(n408), .S(n409) );
  FA_X1 U403 ( .A(n599), .B(n655), .CI(n641), .CO(n412), .S(n413) );
  FA_X1 U404 ( .A(n954), .B(n585), .CI(n670), .CO(n414), .S(n415) );
  FA_X1 U405 ( .A(n432), .B(n421), .CI(n419), .CO(n416), .S(n417) );
  FA_X1 U406 ( .A(n423), .B(n436), .CI(n434), .CO(n418), .S(n419) );
  FA_X1 U409 ( .A(n600), .B(n642), .CI(n628), .CO(n424), .S(n425) );
  FA_X1 U410 ( .A(n586), .B(n614), .CI(n656), .CO(n426), .S(n427) );
  FA_X1 U415 ( .A(n443), .B(n456), .CI(n454), .CO(n436), .S(n437) );
  FA_X1 U416 ( .A(n615), .B(n657), .CI(n671), .CO(n438), .S(n439) );
  FA_X1 U417 ( .A(n587), .B(n629), .CI(n686), .CO(n440), .S(n441) );
  FA_X1 U421 ( .A(n462), .B(n455), .CI(n451), .CO(n446), .S(n447) );
  FA_X1 U422 ( .A(n464), .B(n466), .CI(n453), .CO(n448), .S(n449) );
  FA_X1 U423 ( .A(n457), .B(n672), .CI(n468), .CO(n450), .S(n451) );
  FA_X1 U424 ( .A(n687), .B(n630), .CI(n658), .CO(n452), .S(n453) );
  FA_X1 U425 ( .A(n602), .B(n644), .CI(n616), .CO(n454), .S(n455) );
  HA_X1 U426 ( .A(n566), .B(n588), .CO(n456), .S(n457) );
  FA_X1 U428 ( .A(n465), .B(n467), .CI(n474), .CO(n460), .S(n461) );
  FA_X1 U429 ( .A(n476), .B(n478), .CI(n469), .CO(n462), .S(n463) );
  FA_X1 U430 ( .A(n645), .B(n659), .CI(n480), .CO(n464), .S(n465) );
  FA_X1 U431 ( .A(n603), .B(n673), .CI(n631), .CO(n466), .S(n467) );
  FA_X1 U432 ( .A(n688), .B(n589), .CI(n617), .CO(n468), .S(n469) );
  FA_X1 U435 ( .A(n490), .B(n481), .CI(n488), .CO(n474), .S(n475) );
  FA_X1 U436 ( .A(n618), .B(n660), .CI(n632), .CO(n476), .S(n477) );
  FA_X1 U437 ( .A(n689), .B(n646), .CI(n674), .CO(n478), .S(n479) );
  HA_X1 U438 ( .A(n604), .B(n567), .CO(n480), .S(n481) );
  FA_X1 U440 ( .A(n489), .B(n491), .CI(n496), .CO(n484), .S(n485) );
  FA_X1 U441 ( .A(n500), .B(n661), .CI(n498), .CO(n486), .S(n487) );
  FA_X1 U442 ( .A(n619), .B(n647), .CI(n675), .CO(n488), .S(n489) );
  FA_X1 U443 ( .A(n690), .B(n605), .CI(n633), .CO(n490), .S(n491) );
  FA_X1 U444 ( .A(n504), .B(n497), .CI(n495), .CO(n492), .S(n493) );
  FA_X1 U445 ( .A(n506), .B(n508), .CI(n499), .CO(n494), .S(n495) );
  FA_X1 U447 ( .A(n634), .B(n662), .CI(n691), .CO(n498), .S(n499) );
  HA_X1 U448 ( .A(n620), .B(n568), .CO(n500), .S(n501) );
  FA_X1 U449 ( .A(n512), .B(n507), .CI(n505), .CO(n502), .S(n503) );
  FA_X1 U450 ( .A(n514), .B(n516), .CI(n509), .CO(n504), .S(n505) );
  FA_X1 U451 ( .A(n635), .B(n677), .CI(n663), .CO(n506), .S(n507) );
  FA_X1 U452 ( .A(n649), .B(n621), .CI(n692), .CO(n508), .S(n509) );
  FA_X1 U453 ( .A(n515), .B(n520), .CI(n513), .CO(n510), .S(n511) );
  FA_X1 U454 ( .A(n517), .B(n693), .CI(n522), .CO(n512), .S(n513) );
  FA_X1 U455 ( .A(n650), .B(n678), .CI(n664), .CO(n514), .S(n515) );
  HA_X1 U456 ( .A(n569), .B(n636), .CO(n516), .S(n517) );
  FA_X1 U457 ( .A(n523), .B(n526), .CI(n521), .CO(n518), .S(n519) );
  FA_X1 U458 ( .A(n651), .B(n679), .CI(n528), .CO(n520), .S(n521) );
  FA_X1 U459 ( .A(n665), .B(n637), .CI(n694), .CO(n522), .S(n523) );
  FA_X1 U460 ( .A(n532), .B(n529), .CI(n527), .CO(n524), .S(n525) );
  FA_X1 U461 ( .A(n666), .B(n695), .CI(n680), .CO(n526), .S(n527) );
  HA_X1 U462 ( .A(n570), .B(n652), .CO(n528), .S(n529) );
  FA_X1 U463 ( .A(n536), .B(n667), .CI(n533), .CO(n530), .S(n531) );
  FA_X1 U464 ( .A(n696), .B(n653), .CI(n681), .CO(n532), .S(n533) );
  HA_X1 U466 ( .A(n571), .B(n668), .CO(n536), .S(n537) );
  FA_X1 U467 ( .A(n698), .B(n669), .CI(n683), .CO(n538), .S(n539) );
  HA_X1 U468 ( .A(n684), .B(n699), .CO(n540), .S(n541) );
  OAI22_X1 U822 ( .A1(n12), .A2(n811), .B1(n10), .B2(n810), .ZN(n676) );
  CLKBUF_X3 U823 ( .A(b[4]), .Z(n849) );
  BUF_X1 U824 ( .A(n427), .Z(n953) );
  OR2_X2 U825 ( .A1(n643), .A2(n601), .ZN(n442) );
  OAI22_X1 U826 ( .A1(n12), .A2(n805), .B1(n10), .B2(n804), .ZN(n954) );
  AND2_X1 U827 ( .A1(n483), .A2(n492), .ZN(n957) );
  INV_X1 U828 ( .A(n957), .ZN(n253) );
  BUF_X1 U829 ( .A(n822), .Z(n955) );
  CLKBUF_X1 U830 ( .A(n839), .Z(n956) );
  CLKBUF_X2 U831 ( .A(b[1]), .Z(n852) );
  BUF_X1 U832 ( .A(n867), .Z(n17) );
  BUF_X2 U833 ( .A(n875), .Z(n15) );
  BUF_X2 U834 ( .A(b[2]), .Z(n851) );
  CLKBUF_X3 U835 ( .A(b[11]), .Z(n842) );
  XOR2_X1 U836 ( .A(n441), .B(n452), .Z(n958) );
  XOR2_X1 U837 ( .A(n439), .B(n958), .Z(n435) );
  NAND2_X1 U838 ( .A1(n439), .A2(n441), .ZN(n959) );
  NAND2_X1 U839 ( .A1(n439), .A2(n452), .ZN(n960) );
  NAND2_X1 U840 ( .A1(n441), .A2(n452), .ZN(n961) );
  NAND3_X1 U841 ( .A1(n959), .A2(n960), .A3(n961), .ZN(n434) );
  XOR2_X1 U842 ( .A(n676), .B(n648), .Z(n962) );
  XOR2_X1 U843 ( .A(n501), .B(n962), .Z(n497) );
  NAND2_X1 U844 ( .A1(n501), .A2(n676), .ZN(n963) );
  NAND2_X1 U845 ( .A1(n501), .A2(n648), .ZN(n964) );
  NAND2_X4 U846 ( .A1(n676), .A2(n648), .ZN(n965) );
  NAND3_X1 U847 ( .A1(n963), .A2(n964), .A3(n965), .ZN(n496) );
  OAI22_X2 U848 ( .A1(n24), .A2(n781), .B1(n21), .B2(n780), .ZN(n648) );
  XOR2_X1 U849 ( .A(n682), .B(n697), .Z(n966) );
  XOR2_X1 U850 ( .A(n537), .B(n966), .Z(n535) );
  NAND2_X1 U851 ( .A1(n537), .A2(n682), .ZN(n967) );
  NAND2_X1 U852 ( .A1(n537), .A2(n697), .ZN(n968) );
  NAND2_X1 U853 ( .A1(n682), .A2(n697), .ZN(n969) );
  NAND3_X1 U854 ( .A1(n967), .A2(n968), .A3(n969), .ZN(n534) );
  BUF_X2 U855 ( .A(b[15]), .Z(n838) );
  BUF_X2 U856 ( .A(n867), .Z(n1058) );
  NOR2_X2 U857 ( .A1(n373), .A2(n382), .ZN(n190) );
  BUF_X2 U858 ( .A(n866), .Z(n23) );
  NOR2_X2 U859 ( .A1(n190), .A2(n153), .ZN(n151) );
  BUF_X1 U860 ( .A(n848), .Z(n1026) );
  BUF_X2 U861 ( .A(n876), .Z(n10) );
  BUF_X2 U862 ( .A(n868), .Z(n12) );
  XNOR2_X1 U863 ( .A(n220), .B(n970), .ZN(product[17]) );
  AND2_X1 U864 ( .A1(n217), .A2(n1044), .ZN(n970) );
  BUF_X1 U865 ( .A(n872), .Z(n33) );
  OAI21_X1 U866 ( .B1(n199), .B2(n205), .A(n200), .ZN(n971) );
  CLKBUF_X3 U867 ( .A(b[13]), .Z(n840) );
  XNOR2_X1 U868 ( .A(n448), .B(n972), .ZN(n433) );
  XNOR2_X1 U869 ( .A(n437), .B(n450), .ZN(n972) );
  CLKBUF_X1 U870 ( .A(b[0]), .Z(n49) );
  BUF_X4 U871 ( .A(a[3]), .Z(n7) );
  BUF_X2 U872 ( .A(b[8]), .Z(n845) );
  BUF_X2 U873 ( .A(n865), .Z(n29) );
  BUF_X1 U874 ( .A(n867), .Z(n18) );
  BUF_X2 U875 ( .A(n862), .Z(n47) );
  OAI21_X1 U876 ( .B1(n199), .B2(n205), .A(n200), .ZN(n198) );
  OAI22_X1 U877 ( .A1(n48), .A2(n703), .B1(n46), .B2(n702), .ZN(n332) );
  BUF_X2 U878 ( .A(n49), .Z(n1064) );
  AOI21_X1 U879 ( .B1(n1008), .B2(n289), .A(n286), .ZN(n284) );
  XOR2_X1 U880 ( .A(n442), .B(n429), .Z(n973) );
  XOR2_X1 U881 ( .A(n440), .B(n973), .Z(n423) );
  NAND2_X1 U882 ( .A1(n440), .A2(n442), .ZN(n974) );
  NAND2_X1 U883 ( .A1(n440), .A2(n429), .ZN(n975) );
  NAND2_X1 U884 ( .A1(n442), .A2(n429), .ZN(n976) );
  NAND3_X1 U885 ( .A1(n974), .A2(n975), .A3(n976), .ZN(n422) );
  XOR2_X1 U886 ( .A(n460), .B(n449), .Z(n977) );
  XOR2_X1 U887 ( .A(n447), .B(n977), .Z(n445) );
  NAND2_X1 U888 ( .A1(n447), .A2(n460), .ZN(n978) );
  NAND2_X1 U889 ( .A1(n447), .A2(n449), .ZN(n979) );
  NAND2_X1 U890 ( .A1(n460), .A2(n449), .ZN(n980) );
  NAND3_X1 U891 ( .A1(n978), .A2(n979), .A3(n980), .ZN(n444) );
  XOR2_X1 U892 ( .A(n472), .B(n463), .Z(n981) );
  XOR2_X1 U893 ( .A(n461), .B(n981), .Z(n459) );
  NAND2_X1 U894 ( .A1(n461), .A2(n472), .ZN(n982) );
  NAND2_X1 U895 ( .A1(n461), .A2(n463), .ZN(n983) );
  NAND2_X1 U896 ( .A1(n472), .A2(n463), .ZN(n984) );
  NAND3_X1 U897 ( .A1(n982), .A2(n983), .A3(n984), .ZN(n458) );
  NAND2_X1 U898 ( .A1(n448), .A2(n437), .ZN(n985) );
  NAND2_X1 U899 ( .A1(n448), .A2(n450), .ZN(n986) );
  NAND2_X1 U900 ( .A1(n437), .A2(n450), .ZN(n987) );
  NAND3_X1 U901 ( .A1(n985), .A2(n986), .A3(n987), .ZN(n432) );
  XOR2_X1 U902 ( .A(n613), .B(n627), .Z(n988) );
  XOR2_X1 U903 ( .A(n426), .B(n988), .Z(n411) );
  NAND2_X1 U904 ( .A1(n426), .A2(n613), .ZN(n989) );
  NAND2_X1 U905 ( .A1(n426), .A2(n627), .ZN(n990) );
  NAND2_X1 U906 ( .A1(n613), .A2(n627), .ZN(n991) );
  NAND3_X1 U907 ( .A1(n989), .A2(n990), .A3(n991), .ZN(n410) );
  XOR2_X1 U908 ( .A(n379), .B(n388), .Z(n992) );
  XOR2_X1 U909 ( .A(n386), .B(n992), .Z(n375) );
  NAND2_X1 U910 ( .A1(n386), .A2(n379), .ZN(n993) );
  NAND2_X1 U911 ( .A1(n386), .A2(n388), .ZN(n994) );
  NAND2_X1 U912 ( .A1(n379), .A2(n388), .ZN(n995) );
  NAND3_X1 U913 ( .A1(n993), .A2(n994), .A3(n995), .ZN(n374) );
  XOR2_X1 U914 ( .A(n953), .B(n438), .Z(n996) );
  XOR2_X1 U915 ( .A(n425), .B(n996), .Z(n421) );
  NAND2_X1 U916 ( .A1(n425), .A2(n427), .ZN(n997) );
  NAND2_X1 U917 ( .A1(n425), .A2(n438), .ZN(n998) );
  NAND2_X1 U918 ( .A1(n427), .A2(n438), .ZN(n999) );
  NAND3_X1 U919 ( .A1(n997), .A2(n998), .A3(n999), .ZN(n420) );
  OR2_X1 U920 ( .A1(n483), .A2(n492), .ZN(n1000) );
  OR2_X1 U921 ( .A1(n503), .A2(n510), .ZN(n1001) );
  OR2_X1 U922 ( .A1(n334), .A2(n333), .ZN(n1002) );
  OR2_X1 U923 ( .A1(n337), .A2(n340), .ZN(n1003) );
  OR2_X1 U924 ( .A1(n574), .A2(n332), .ZN(n1004) );
  OR2_X1 U925 ( .A1(n511), .A2(n518), .ZN(n1005) );
  OR2_X1 U926 ( .A1(n471), .A2(n482), .ZN(n1006) );
  OR2_X1 U927 ( .A1(n493), .A2(n502), .ZN(n1007) );
  OR2_X1 U928 ( .A1(n535), .A2(n538), .ZN(n1008) );
  OR2_X1 U929 ( .A1(n541), .A2(n572), .ZN(n1009) );
  OR2_X1 U930 ( .A1(n336), .A2(n335), .ZN(n1010) );
  OR2_X1 U931 ( .A1(n525), .A2(n530), .ZN(n1011) );
  BUF_X1 U932 ( .A(n225), .Z(n1060) );
  OR2_X1 U933 ( .A1(n701), .A2(n573), .ZN(n1012) );
  CLKBUF_X2 U934 ( .A(b[3]), .Z(n850) );
  AOI21_X1 U935 ( .B1(n971), .B2(n151), .A(n152), .ZN(n1013) );
  AOI21_X1 U936 ( .B1(n971), .B2(n151), .A(n152), .ZN(n1014) );
  AOI21_X1 U937 ( .B1(n971), .B2(n151), .A(n152), .ZN(n150) );
  BUF_X1 U938 ( .A(n875), .Z(n16) );
  CLKBUF_X1 U939 ( .A(n871), .Z(n39) );
  CLKBUF_X3 U940 ( .A(n871), .Z(n40) );
  XOR2_X1 U941 ( .A(n494), .B(n487), .Z(n1015) );
  XOR2_X1 U942 ( .A(n1015), .B(n485), .Z(n483) );
  NAND2_X1 U943 ( .A1(n485), .A2(n494), .ZN(n1016) );
  NAND2_X1 U944 ( .A1(n485), .A2(n487), .ZN(n1017) );
  NAND2_X1 U945 ( .A1(n494), .A2(n487), .ZN(n1018) );
  NAND3_X1 U946 ( .A1(n1016), .A2(n1017), .A3(n1018), .ZN(n482) );
  CLKBUF_X1 U947 ( .A(n211), .Z(n1019) );
  BUF_X2 U948 ( .A(b[12]), .Z(n841) );
  AOI21_X1 U949 ( .B1(n273), .B2(n1005), .A(n270), .ZN(n1020) );
  AOI21_X1 U950 ( .B1(n273), .B2(n1005), .A(n270), .ZN(n268) );
  BUF_X4 U951 ( .A(a[7]), .Z(n19) );
  BUF_X2 U952 ( .A(n874), .Z(n22) );
  INV_X1 U953 ( .A(n148), .ZN(n1021) );
  NOR2_X2 U954 ( .A1(n383), .A2(n392), .ZN(n199) );
  XNOR2_X1 U955 ( .A(n1022), .B(n473), .ZN(n471) );
  XNOR2_X1 U956 ( .A(n484), .B(n475), .ZN(n1022) );
  CLKBUF_X1 U957 ( .A(n218), .Z(n1023) );
  XNOR2_X1 U958 ( .A(n139), .B(n1024), .ZN(product[26]) );
  AND2_X1 U959 ( .A1(n306), .A2(n138), .ZN(n1024) );
  XNOR2_X1 U960 ( .A(n201), .B(n1025), .ZN(product[20]) );
  AND2_X1 U961 ( .A1(n312), .A2(n200), .ZN(n1025) );
  CLKBUF_X1 U962 ( .A(n273), .Z(n1027) );
  XNOR2_X1 U963 ( .A(n433), .B(n1028), .ZN(n431) );
  XNOR2_X1 U964 ( .A(n446), .B(n435), .ZN(n1028) );
  BUF_X2 U965 ( .A(n866), .Z(n24) );
  OR2_X1 U966 ( .A1(n459), .A2(n470), .ZN(n1029) );
  CLKBUF_X1 U967 ( .A(n242), .Z(n1030) );
  BUF_X2 U968 ( .A(n872), .Z(n34) );
  XNOR2_X1 U969 ( .A(n1), .B(n838), .ZN(n1031) );
  BUF_X4 U970 ( .A(a[1]), .Z(n1) );
  OR2_X1 U971 ( .A1(n365), .A2(n372), .ZN(n1032) );
  CLKBUF_X1 U972 ( .A(n843), .Z(n1033) );
  CLKBUF_X2 U973 ( .A(n206), .Z(n1039) );
  XNOR2_X1 U974 ( .A(n183), .B(n1034), .ZN(product[22]) );
  AND2_X1 U975 ( .A1(n175), .A2(n182), .ZN(n1034) );
  XNOR2_X1 U976 ( .A(n1035), .B(n486), .ZN(n473) );
  XNOR2_X1 U977 ( .A(n479), .B(n477), .ZN(n1035) );
  BUF_X2 U978 ( .A(b[6]), .Z(n1036) );
  OAI21_X1 U979 ( .B1(n256), .B2(n1020), .A(n257), .ZN(n1037) );
  XNOR2_X1 U980 ( .A(n31), .B(n847), .ZN(n1038) );
  BUF_X2 U981 ( .A(b[6]), .Z(n847) );
  BUF_X2 U982 ( .A(n865), .Z(n30) );
  OAI22_X1 U983 ( .A1(n1058), .A2(n788), .B1(n16), .B2(n787), .ZN(n1040) );
  NOR2_X1 U984 ( .A1(n405), .A2(n416), .ZN(n1041) );
  XNOR2_X1 U985 ( .A(n130), .B(n1042), .ZN(product[27]) );
  AND2_X1 U986 ( .A1(n1003), .A2(n129), .ZN(n1042) );
  XNOR2_X1 U987 ( .A(n192), .B(n1043), .ZN(product[21]) );
  AND2_X1 U988 ( .A1(n188), .A2(n191), .ZN(n1043) );
  CLKBUF_X1 U989 ( .A(n219), .Z(n1044) );
  BUF_X4 U990 ( .A(a[11]), .Z(n31) );
  BUF_X2 U991 ( .A(n864), .Z(n36) );
  NAND2_X1 U992 ( .A1(n433), .A2(n446), .ZN(n1045) );
  NAND2_X1 U993 ( .A1(n433), .A2(n435), .ZN(n1046) );
  NAND2_X1 U994 ( .A1(n446), .A2(n435), .ZN(n1047) );
  NAND3_X1 U995 ( .A1(n1045), .A2(n1046), .A3(n1047), .ZN(n430) );
  NOR2_X1 U996 ( .A1(n531), .A2(n534), .ZN(n282) );
  CLKBUF_X2 U997 ( .A(b[7]), .Z(n846) );
  NAND2_X1 U998 ( .A1(n479), .A2(n477), .ZN(n1048) );
  NAND2_X1 U999 ( .A1(n479), .A2(n486), .ZN(n1049) );
  NAND2_X1 U1000 ( .A1(n477), .A2(n486), .ZN(n1050) );
  NAND3_X1 U1001 ( .A1(n1048), .A2(n1049), .A3(n1050), .ZN(n472) );
  NAND2_X1 U1002 ( .A1(n484), .A2(n475), .ZN(n1051) );
  NAND2_X1 U1003 ( .A1(n484), .A2(n473), .ZN(n1052) );
  NAND2_X1 U1004 ( .A1(n475), .A2(n473), .ZN(n1053) );
  NAND3_X1 U1005 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n470) );
  OR2_X1 U1006 ( .A1(n6), .A2(n826), .ZN(n1054) );
  OR2_X1 U1007 ( .A1(n825), .A2(n4), .ZN(n1055) );
  NAND2_X1 U1008 ( .A1(n1054), .A2(n1055), .ZN(n691) );
  BUF_X2 U1009 ( .A(n869), .Z(n6) );
  BUF_X2 U1010 ( .A(n877), .Z(n4) );
  CLKBUF_X1 U1011 ( .A(n233), .Z(n1056) );
  NOR2_X1 U1012 ( .A1(n431), .A2(n444), .ZN(n1057) );
  BUF_X4 U1013 ( .A(a[9]), .Z(n25) );
  BUF_X4 U1014 ( .A(a[5]), .Z(n13) );
  OAI21_X1 U1015 ( .B1(n282), .B2(n284), .A(n283), .ZN(n281) );
  OAI21_X1 U1016 ( .B1(n276), .B2(n274), .A(n275), .ZN(n273) );
  XNOR2_X1 U1017 ( .A(n170), .B(n1059), .ZN(product[23]) );
  AND2_X1 U1018 ( .A1(n167), .A2(n169), .ZN(n1059) );
  BUF_X2 U1019 ( .A(n863), .Z(n41) );
  BUF_X4 U1020 ( .A(a[13]), .Z(n37) );
  BUF_X2 U1021 ( .A(b[14]), .Z(n839) );
  BUF_X2 U1022 ( .A(b[9]), .Z(n844) );
  BUF_X2 U1023 ( .A(b[5]), .Z(n848) );
  BUF_X2 U1024 ( .A(n49), .Z(n1065) );
  BUF_X2 U1025 ( .A(b[10]), .Z(n843) );
  AOI21_X1 U1026 ( .B1(n236), .B2(n1037), .A(n237), .ZN(n1061) );
  NAND2_X1 U1027 ( .A1(n197), .A2(n151), .ZN(n1062) );
  NOR2_X1 U1028 ( .A1(n345), .A2(n350), .ZN(n144) );
  NOR2_X1 U1029 ( .A1(n341), .A2(n344), .ZN(n137) );
  NOR2_X1 U1030 ( .A1(n700), .A2(n685), .ZN(n298) );
  NOR2_X1 U1031 ( .A1(n539), .A2(n540), .ZN(n290) );
  AND2_X1 U1032 ( .A1(n1012), .A2(n301), .ZN(product[1]) );
  BUF_X1 U1033 ( .A(n874), .Z(n21) );
  INV_X1 U1034 ( .A(n224), .ZN(n222) );
  INV_X1 U1035 ( .A(n1060), .ZN(n223) );
  INV_X1 U1036 ( .A(n226), .ZN(n224) );
  NOR2_X1 U1037 ( .A1(n195), .A2(n162), .ZN(n160) );
  NOR2_X1 U1038 ( .A1(n195), .A2(n190), .ZN(n184) );
  NOR2_X1 U1039 ( .A1(n195), .A2(n173), .ZN(n171) );
  INV_X1 U1040 ( .A(n177), .ZN(n175) );
  NOR2_X1 U1041 ( .A1(n223), .A2(n1023), .ZN(n214) );
  INV_X1 U1042 ( .A(n195), .ZN(n193) );
  INV_X1 U1043 ( .A(n98), .ZN(n96) );
  XNOR2_X1 U1044 ( .A(n240), .B(n70), .ZN(product[14]) );
  NAND2_X1 U1045 ( .A1(n1029), .A2(n239), .ZN(n70) );
  NAND2_X1 U1046 ( .A1(n313), .A2(n205), .ZN(n65) );
  NAND2_X1 U1047 ( .A1(n317), .A2(n1056), .ZN(n69) );
  INV_X1 U1048 ( .A(n232), .ZN(n317) );
  XOR2_X1 U1049 ( .A(n229), .B(n68), .Z(product[16]) );
  NAND2_X1 U1050 ( .A1(n316), .A2(n228), .ZN(n68) );
  INV_X1 U1051 ( .A(n1057), .ZN(n316) );
  INV_X1 U1052 ( .A(n197), .ZN(n195) );
  XOR2_X1 U1053 ( .A(n213), .B(n66), .Z(product[18]) );
  NAND2_X1 U1054 ( .A1(n314), .A2(n212), .ZN(n66) );
  INV_X1 U1055 ( .A(n1019), .ZN(n314) );
  NOR2_X1 U1056 ( .A1(n177), .A2(n166), .ZN(n164) );
  NOR2_X1 U1057 ( .A1(n124), .A2(n100), .ZN(n98) );
  OAI21_X1 U1058 ( .B1(n196), .B2(n173), .A(n174), .ZN(n172) );
  AOI21_X1 U1059 ( .B1(n189), .B2(n175), .A(n176), .ZN(n174) );
  INV_X1 U1060 ( .A(n178), .ZN(n176) );
  INV_X1 U1061 ( .A(n198), .ZN(n196) );
  INV_X1 U1062 ( .A(n1020), .ZN(n267) );
  INV_X1 U1063 ( .A(n1037), .ZN(n254) );
  NAND2_X1 U1064 ( .A1(n164), .A2(n188), .ZN(n162) );
  OAI21_X1 U1065 ( .B1(n196), .B2(n190), .A(n191), .ZN(n185) );
  NAND2_X1 U1066 ( .A1(n188), .A2(n175), .ZN(n173) );
  OAI21_X1 U1067 ( .B1(n224), .B2(n1023), .A(n1044), .ZN(n215) );
  INV_X1 U1068 ( .A(n1032), .ZN(n177) );
  INV_X1 U1069 ( .A(n1023), .ZN(n217) );
  INV_X1 U1070 ( .A(n180), .ZN(n178) );
  INV_X1 U1071 ( .A(n124), .ZN(n122) );
  NAND2_X1 U1072 ( .A1(n1006), .A2(n1000), .ZN(n241) );
  NAND2_X1 U1073 ( .A1(n122), .A2(n1010), .ZN(n109) );
  INV_X1 U1074 ( .A(n1000), .ZN(n248) );
  INV_X1 U1075 ( .A(n1056), .ZN(n231) );
  INV_X1 U1076 ( .A(n205), .ZN(n203) );
  NAND2_X1 U1077 ( .A1(n1005), .A2(n272), .ZN(n75) );
  XOR2_X1 U1078 ( .A(n254), .B(n72), .Z(product[12]) );
  NAND2_X1 U1079 ( .A1(n1000), .A2(n253), .ZN(n72) );
  XNOR2_X1 U1080 ( .A(n267), .B(n74), .ZN(product[10]) );
  NAND2_X1 U1081 ( .A1(n1001), .A2(n266), .ZN(n74) );
  INV_X1 U1082 ( .A(n272), .ZN(n270) );
  AOI21_X1 U1083 ( .B1(n1007), .B2(n264), .A(n259), .ZN(n257) );
  NAND2_X1 U1084 ( .A1(n1007), .A2(n1001), .ZN(n256) );
  NOR2_X1 U1085 ( .A1(n417), .A2(n430), .ZN(n218) );
  NOR2_X1 U1086 ( .A1(n445), .A2(n458), .ZN(n232) );
  NOR2_X1 U1087 ( .A1(n431), .A2(n444), .ZN(n227) );
  NOR2_X1 U1088 ( .A1(n405), .A2(n416), .ZN(n211) );
  INV_X1 U1089 ( .A(n199), .ZN(n312) );
  NAND2_X1 U1090 ( .A1(n308), .A2(n158), .ZN(n60) );
  INV_X1 U1091 ( .A(n157), .ZN(n308) );
  INV_X1 U1092 ( .A(n190), .ZN(n188) );
  XOR2_X1 U1093 ( .A(n146), .B(n59), .Z(product[25]) );
  NAND2_X1 U1094 ( .A1(n143), .A2(n145), .ZN(n59) );
  NAND2_X1 U1095 ( .A1(n445), .A2(n458), .ZN(n233) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n246), .ZN(n71) );
  NOR2_X1 U1097 ( .A1(n459), .A2(n470), .ZN(n238) );
  INV_X1 U1098 ( .A(n136), .ZN(n134) );
  AOI21_X1 U1099 ( .B1(n123), .B2(n1010), .A(n114), .ZN(n110) );
  INV_X1 U1100 ( .A(n99), .ZN(n97) );
  XOR2_X1 U1101 ( .A(n262), .B(n73), .Z(product[11]) );
  NAND2_X1 U1102 ( .A1(n1007), .A2(n261), .ZN(n73) );
  AOI21_X1 U1103 ( .B1(n267), .B2(n1001), .A(n264), .ZN(n262) );
  AOI21_X1 U1104 ( .B1(n1006), .B2(n957), .A(n244), .ZN(n242) );
  INV_X1 U1105 ( .A(n246), .ZN(n244) );
  OAI21_X1 U1106 ( .B1(n196), .B2(n162), .A(n163), .ZN(n161) );
  AOI21_X1 U1107 ( .B1(n164), .B2(n189), .A(n165), .ZN(n163) );
  OAI21_X1 U1108 ( .B1(n178), .B2(n166), .A(n169), .ZN(n165) );
  NAND2_X1 U1109 ( .A1(n417), .A2(n430), .ZN(n219) );
  NAND2_X1 U1110 ( .A1(n393), .A2(n404), .ZN(n205) );
  INV_X1 U1111 ( .A(n191), .ZN(n189) );
  INV_X1 U1112 ( .A(n266), .ZN(n264) );
  NAND2_X1 U1113 ( .A1(n1010), .A2(n1002), .ZN(n100) );
  NAND2_X1 U1114 ( .A1(n135), .A2(n1003), .ZN(n124) );
  NAND2_X1 U1115 ( .A1(n459), .A2(n470), .ZN(n239) );
  NAND2_X1 U1116 ( .A1(n431), .A2(n444), .ZN(n228) );
  NAND2_X1 U1117 ( .A1(n405), .A2(n416), .ZN(n212) );
  INV_X1 U1118 ( .A(n167), .ZN(n166) );
  INV_X1 U1119 ( .A(n168), .ZN(n167) );
  INV_X1 U1120 ( .A(n125), .ZN(n123) );
  NAND2_X1 U1121 ( .A1(n98), .A2(n1004), .ZN(n87) );
  INV_X1 U1122 ( .A(n261), .ZN(n259) );
  INV_X1 U1123 ( .A(n135), .ZN(n133) );
  INV_X1 U1124 ( .A(n144), .ZN(n143) );
  NAND2_X1 U1125 ( .A1(n326), .A2(n283), .ZN(n78) );
  INV_X1 U1126 ( .A(n282), .ZN(n326) );
  NAND2_X1 U1127 ( .A1(n324), .A2(n275), .ZN(n76) );
  INV_X1 U1128 ( .A(n274), .ZN(n324) );
  NAND2_X1 U1129 ( .A1(n1011), .A2(n280), .ZN(n77) );
  XNOR2_X1 U1130 ( .A(n79), .B(n289), .ZN(product[5]) );
  NAND2_X1 U1131 ( .A1(n1008), .A2(n288), .ZN(n79) );
  NOR2_X1 U1132 ( .A1(n357), .A2(n364), .ZN(n168) );
  INV_X1 U1133 ( .A(n280), .ZN(n278) );
  NAND2_X1 U1134 ( .A1(n1004), .A2(n92), .ZN(n54) );
  AOI21_X1 U1135 ( .B1(n136), .B2(n1003), .A(n127), .ZN(n125) );
  INV_X1 U1136 ( .A(n129), .ZN(n127) );
  INV_X1 U1137 ( .A(n137), .ZN(n306) );
  XOR2_X1 U1138 ( .A(n106), .B(n55), .Z(product[29]) );
  NAND2_X1 U1139 ( .A1(n1002), .A2(n105), .ZN(n55) );
  OAI21_X1 U1140 ( .B1(n145), .B2(n137), .A(n138), .ZN(n136) );
  OAI21_X1 U1141 ( .B1(n125), .B2(n100), .A(n101), .ZN(n99) );
  AOI21_X1 U1142 ( .B1(n114), .B2(n1002), .A(n103), .ZN(n101) );
  INV_X1 U1143 ( .A(n105), .ZN(n103) );
  XOR2_X1 U1144 ( .A(n117), .B(n56), .Z(product[28]) );
  NAND2_X1 U1145 ( .A1(n1010), .A2(n116), .ZN(n56) );
  NOR2_X1 U1146 ( .A1(n144), .A2(n137), .ZN(n135) );
  INV_X1 U1147 ( .A(n288), .ZN(n286) );
  NOR2_X1 U1148 ( .A1(n351), .A2(n356), .ZN(n157) );
  NAND2_X1 U1149 ( .A1(n471), .A2(n482), .ZN(n246) );
  NAND2_X1 U1150 ( .A1(n345), .A2(n350), .ZN(n145) );
  AOI21_X1 U1151 ( .B1(n99), .B2(n1004), .A(n90), .ZN(n88) );
  INV_X1 U1152 ( .A(n92), .ZN(n90) );
  NAND2_X1 U1153 ( .A1(n373), .A2(n382), .ZN(n191) );
  NAND2_X1 U1154 ( .A1(n493), .A2(n502), .ZN(n261) );
  NAND2_X1 U1155 ( .A1(n351), .A2(n356), .ZN(n158) );
  INV_X1 U1156 ( .A(n116), .ZN(n114) );
  NAND2_X1 U1157 ( .A1(n328), .A2(n291), .ZN(n80) );
  INV_X1 U1158 ( .A(n290), .ZN(n328) );
  XOR2_X1 U1159 ( .A(n82), .B(n301), .Z(product[2]) );
  NAND2_X1 U1160 ( .A1(n330), .A2(n299), .ZN(n82) );
  INV_X1 U1161 ( .A(n298), .ZN(n330) );
  XNOR2_X1 U1162 ( .A(n81), .B(n297), .ZN(product[3]) );
  NAND2_X1 U1163 ( .A1(n1009), .A2(n296), .ZN(n81) );
  OAI21_X1 U1164 ( .B1(n290), .B2(n292), .A(n291), .ZN(n289) );
  NAND2_X1 U1165 ( .A1(n574), .A2(n332), .ZN(n92) );
  OAI21_X1 U1166 ( .B1(n298), .B2(n301), .A(n299), .ZN(n297) );
  INV_X1 U1167 ( .A(n332), .ZN(n333) );
  NAND2_X1 U1168 ( .A1(n700), .A2(n685), .ZN(n299) );
  INV_X1 U1169 ( .A(n428), .ZN(n429) );
  XNOR2_X1 U1170 ( .A(n643), .B(n601), .ZN(n443) );
  NAND2_X1 U1171 ( .A1(n525), .A2(n530), .ZN(n280) );
  NAND2_X1 U1172 ( .A1(n535), .A2(n538), .ZN(n288) );
  NAND2_X1 U1173 ( .A1(n337), .A2(n340), .ZN(n129) );
  NAND2_X1 U1174 ( .A1(n341), .A2(n344), .ZN(n138) );
  NAND2_X1 U1175 ( .A1(n336), .A2(n335), .ZN(n116) );
  NAND2_X1 U1176 ( .A1(n334), .A2(n333), .ZN(n105) );
  NAND2_X1 U1177 ( .A1(n531), .A2(n534), .ZN(n283) );
  OAI22_X1 U1178 ( .A1(n23), .A2(n771), .B1(n22), .B2(n770), .ZN(n380) );
  OAI22_X1 U1179 ( .A1(n42), .A2(n720), .B1(n40), .B2(n719), .ZN(n338) );
  OAI22_X1 U1180 ( .A1(n5), .A2(n835), .B1(n834), .B2(n4), .ZN(n700) );
  OAI22_X1 U1181 ( .A1(n1058), .A2(n788), .B1(n16), .B2(n787), .ZN(n402) );
  OAI22_X1 U1182 ( .A1(n12), .A2(n805), .B1(n10), .B2(n804), .ZN(n428) );
  OAI22_X1 U1183 ( .A1(n23), .A2(n776), .B1(n22), .B2(n775), .ZN(n643) );
  OAI22_X1 U1184 ( .A1(n41), .A2(n731), .B1(n40), .B2(n730), .ZN(n601) );
  AND2_X1 U1185 ( .A1(n1065), .A2(n552), .ZN(n637) );
  OAI22_X1 U1186 ( .A1(n5), .A2(n829), .B1(n828), .B2(n4), .ZN(n694) );
  OAI22_X1 U1187 ( .A1(n1058), .A2(n799), .B1(n15), .B2(n798), .ZN(n665) );
  OAI22_X1 U1188 ( .A1(n35), .A2(n1038), .B1(n33), .B2(n744), .ZN(n614) );
  OAI22_X1 U1189 ( .A1(n47), .A2(n715), .B1(n45), .B2(n714), .ZN(n586) );
  OAI22_X1 U1190 ( .A1(n1058), .A2(n790), .B1(n16), .B2(n789), .ZN(n656) );
  OAI22_X1 U1191 ( .A1(n48), .A2(n704), .B1(n46), .B2(n703), .ZN(n575) );
  INV_X1 U1192 ( .A(n545), .ZN(n590) );
  AOI21_X1 U1193 ( .B1(n42), .B2(n40), .A(n719), .ZN(n545) );
  OAI22_X1 U1194 ( .A1(n48), .A2(n705), .B1(n46), .B2(n704), .ZN(n576) );
  INV_X1 U1195 ( .A(n338), .ZN(n339) );
  OAI22_X1 U1196 ( .A1(n11), .A2(n817), .B1(n10), .B2(n816), .ZN(n682) );
  OAI22_X1 U1197 ( .A1(n5), .A2(n832), .B1(n831), .B2(n4), .ZN(n697) );
  OAI22_X1 U1198 ( .A1(n48), .A2(n706), .B1(n46), .B2(n705), .ZN(n577) );
  OAI22_X1 U1199 ( .A1(n11), .A2(n818), .B1(n10), .B2(n817), .ZN(n683) );
  OAI22_X1 U1200 ( .A1(n5), .A2(n833), .B1(n832), .B2(n4), .ZN(n698) );
  AND2_X1 U1201 ( .A1(n1065), .A2(n558), .ZN(n669) );
  AOI21_X1 U1202 ( .B1(n23), .B2(n22), .A(n770), .ZN(n554) );
  OAI22_X1 U1203 ( .A1(n48), .A2(n878), .B1(n718), .B2(n46), .ZN(n566) );
  OAI22_X1 U1204 ( .A1(n47), .A2(n717), .B1(n45), .B2(n716), .ZN(n588) );
  OR2_X1 U1205 ( .A1(n1064), .A2(n878), .ZN(n718) );
  OAI22_X1 U1206 ( .A1(n24), .A2(n779), .B1(n21), .B2(n778), .ZN(n646) );
  OAI22_X1 U1207 ( .A1(n12), .A2(n809), .B1(n10), .B2(n808), .ZN(n674) );
  OAI22_X1 U1208 ( .A1(n6), .A2(n824), .B1(n823), .B2(n4), .ZN(n689) );
  OAI22_X1 U1209 ( .A1(n36), .A2(n742), .B1(n34), .B2(n741), .ZN(n611) );
  OAI22_X1 U1210 ( .A1(n23), .A2(n772), .B1(n22), .B2(n771), .ZN(n639) );
  OAI22_X1 U1211 ( .A1(n42), .A2(n727), .B1(n40), .B2(n726), .ZN(n597) );
  OAI22_X1 U1212 ( .A1(n30), .A2(n760), .B1(n28), .B2(n759), .ZN(n628) );
  OAI22_X1 U1213 ( .A1(n24), .A2(n775), .B1(n22), .B2(n774), .ZN(n642) );
  OAI22_X1 U1214 ( .A1(n41), .A2(n730), .B1(n39), .B2(n729), .ZN(n600) );
  INV_X1 U1215 ( .A(n542), .ZN(n574) );
  AOI21_X1 U1216 ( .B1(n48), .B2(n46), .A(n702), .ZN(n542) );
  AOI21_X1 U1217 ( .B1(n6), .B2(n4), .A(n821), .ZN(n563) );
  AOI21_X1 U1218 ( .B1(n30), .B2(n28), .A(n753), .ZN(n551) );
  OAI22_X1 U1219 ( .A1(n1058), .A2(n801), .B1(n15), .B2(n800), .ZN(n667) );
  NAND2_X1 U1220 ( .A1(n701), .A2(n573), .ZN(n301) );
  AND2_X1 U1221 ( .A1(n1065), .A2(n561), .ZN(n685) );
  INV_X1 U1222 ( .A(n10), .ZN(n561) );
  OAI22_X1 U1223 ( .A1(n47), .A2(n712), .B1(n45), .B2(n711), .ZN(n583) );
  INV_X1 U1224 ( .A(n557), .ZN(n654) );
  AOI21_X1 U1225 ( .B1(n1058), .B2(n16), .A(n787), .ZN(n557) );
  OAI22_X1 U1226 ( .A1(n48), .A2(n707), .B1(n46), .B2(n706), .ZN(n578) );
  OAI22_X1 U1227 ( .A1(n42), .A2(n722), .B1(n40), .B2(n721), .ZN(n592) );
  OAI22_X1 U1228 ( .A1(n30), .A2(n759), .B1(n28), .B2(n758), .ZN(n627) );
  OAI22_X1 U1229 ( .A1(n36), .A2(n744), .B1(n33), .B2(n743), .ZN(n613) );
  OAI22_X1 U1230 ( .A1(n864), .A2(n746), .B1(n33), .B2(n745), .ZN(n615) );
  OAI22_X1 U1231 ( .A1(n18), .A2(n791), .B1(n790), .B2(n16), .ZN(n657) );
  OAI22_X1 U1232 ( .A1(n12), .A2(n806), .B1(n10), .B2(n805), .ZN(n671) );
  OAI22_X1 U1233 ( .A1(n47), .A2(n711), .B1(n45), .B2(n710), .ZN(n582) );
  OAI22_X1 U1234 ( .A1(n30), .A2(n756), .B1(n28), .B2(n755), .ZN(n624) );
  OAI22_X1 U1235 ( .A1(n42), .A2(n726), .B1(n40), .B2(n725), .ZN(n596) );
  OAI22_X1 U1236 ( .A1(n36), .A2(n750), .B1(n33), .B2(n749), .ZN(n619) );
  OAI22_X1 U1237 ( .A1(n23), .A2(n780), .B1(n21), .B2(n779), .ZN(n647) );
  OAI22_X1 U1238 ( .A1(n12), .A2(n810), .B1(n10), .B2(n809), .ZN(n675) );
  OAI22_X1 U1239 ( .A1(n36), .A2(n740), .B1(n34), .B2(n739), .ZN(n609) );
  OAI22_X1 U1240 ( .A1(n42), .A2(n725), .B1(n40), .B2(n724), .ZN(n595) );
  OAI22_X1 U1241 ( .A1(n23), .A2(n774), .B1(n22), .B2(n773), .ZN(n641) );
  OAI22_X1 U1242 ( .A1(n41), .A2(n729), .B1(n39), .B2(n728), .ZN(n599) );
  OAI22_X1 U1243 ( .A1(n17), .A2(n789), .B1(n16), .B2(n788), .ZN(n655) );
  OAI22_X1 U1244 ( .A1(n36), .A2(n741), .B1(n34), .B2(n740), .ZN(n610) );
  INV_X1 U1245 ( .A(n380), .ZN(n381) );
  OAI22_X1 U1246 ( .A1(n36), .A2(n749), .B1(n33), .B2(n748), .ZN(n618) );
  OAI22_X1 U1247 ( .A1(n1058), .A2(n794), .B1(n16), .B2(n793), .ZN(n660) );
  OAI22_X1 U1248 ( .A1(n6), .A2(n825), .B1(n824), .B2(n4), .ZN(n690) );
  AND2_X1 U1249 ( .A1(n1065), .A2(n546), .ZN(n605) );
  OAI22_X1 U1250 ( .A1(n6), .A2(n828), .B1(n827), .B2(n4), .ZN(n693) );
  OAI22_X1 U1251 ( .A1(n1058), .A2(n797), .B1(n15), .B2(n796), .ZN(n663) );
  OAI22_X1 U1252 ( .A1(n11), .A2(n812), .B1(n10), .B2(n811), .ZN(n677) );
  OAI22_X1 U1253 ( .A1(n24), .A2(n783), .B1(n21), .B2(n782), .ZN(n650) );
  OAI22_X1 U1254 ( .A1(n11), .A2(n813), .B1(n10), .B2(n812), .ZN(n678) );
  OAI22_X1 U1255 ( .A1(n1058), .A2(n798), .B1(n15), .B2(n797), .ZN(n664) );
  OAI22_X1 U1256 ( .A1(n30), .A2(n758), .B1(n28), .B2(n757), .ZN(n626) );
  OAI22_X1 U1257 ( .A1(n773), .A2(n23), .B1(n22), .B2(n772), .ZN(n640) );
  OAI22_X1 U1258 ( .A1(n36), .A2(n743), .B1(n34), .B2(n742), .ZN(n612) );
  OAI22_X1 U1259 ( .A1(n24), .A2(n778), .B1(n21), .B2(n777), .ZN(n645) );
  OAI22_X1 U1260 ( .A1(n1058), .A2(n793), .B1(n16), .B2(n792), .ZN(n659) );
  OAI22_X1 U1261 ( .A1(n30), .A2(n755), .B1(n28), .B2(n754), .ZN(n623) );
  OAI22_X1 U1262 ( .A1(n47), .A2(n710), .B1(n45), .B2(n709), .ZN(n581) );
  INV_X1 U1263 ( .A(n554), .ZN(n638) );
  OAI22_X1 U1264 ( .A1(n47), .A2(n714), .B1(n45), .B2(n713), .ZN(n585) );
  INV_X1 U1265 ( .A(n560), .ZN(n670) );
  AOI21_X1 U1266 ( .B1(n12), .B2(n10), .A(n804), .ZN(n560) );
  OAI22_X1 U1267 ( .A1(n42), .A2(n721), .B1(n40), .B2(n720), .ZN(n591) );
  INV_X1 U1268 ( .A(n548), .ZN(n606) );
  AOI21_X1 U1269 ( .B1(n36), .B2(n34), .A(n736), .ZN(n548) );
  OAI22_X1 U1270 ( .A1(n24), .A2(n784), .B1(n21), .B2(n783), .ZN(n651) );
  OAI22_X1 U1271 ( .A1(n11), .A2(n814), .B1(n10), .B2(n813), .ZN(n679) );
  OAI22_X1 U1272 ( .A1(n12), .A2(n807), .B1(n10), .B2(n806), .ZN(n672) );
  OAI22_X1 U1273 ( .A1(n6), .A2(n955), .B1(n1031), .B2(n4), .ZN(n687) );
  OAI22_X1 U1274 ( .A1(n1058), .A2(n792), .B1(n16), .B2(n791), .ZN(n658) );
  OAI22_X1 U1275 ( .A1(n17), .A2(n800), .B1(n15), .B2(n799), .ZN(n666) );
  OAI22_X1 U1276 ( .A1(n5), .A2(n830), .B1(n829), .B2(n4), .ZN(n695) );
  OAI22_X1 U1277 ( .A1(n11), .A2(n815), .B1(n10), .B2(n814), .ZN(n680) );
  OAI22_X1 U1278 ( .A1(n11), .A2(n816), .B1(n10), .B2(n815), .ZN(n681) );
  AND2_X1 U1279 ( .A1(n1065), .A2(n555), .ZN(n653) );
  OAI22_X1 U1280 ( .A1(n5), .A2(n831), .B1(n830), .B2(n4), .ZN(n696) );
  OAI22_X1 U1281 ( .A1(n41), .A2(n733), .B1(n40), .B2(n732), .ZN(n603) );
  OAI22_X1 U1282 ( .A1(n12), .A2(n808), .B1(n10), .B2(n807), .ZN(n673) );
  OAI22_X1 U1283 ( .A1(n42), .A2(n723), .B1(n40), .B2(n722), .ZN(n593) );
  OAI22_X1 U1284 ( .A1(n48), .A2(n708), .B1(n46), .B2(n707), .ZN(n579) );
  INV_X1 U1285 ( .A(n551), .ZN(n622) );
  OAI22_X1 U1286 ( .A1(n30), .A2(n757), .B1(n28), .B2(n756), .ZN(n625) );
  OAI22_X1 U1287 ( .A1(n17), .A2(n795), .B1(n15), .B2(n794), .ZN(n661) );
  OAI22_X1 U1288 ( .A1(n47), .A2(n713), .B1(n45), .B2(n712), .ZN(n584) );
  OAI22_X1 U1289 ( .A1(n41), .A2(n728), .B1(n39), .B2(n727), .ZN(n598) );
  INV_X1 U1290 ( .A(n402), .ZN(n403) );
  OAI22_X1 U1291 ( .A1(n36), .A2(n738), .B1(n34), .B2(n737), .ZN(n607) );
  OAI22_X1 U1292 ( .A1(n47), .A2(n716), .B1(n45), .B2(n715), .ZN(n587) );
  INV_X1 U1293 ( .A(n563), .ZN(n686) );
  OAI22_X1 U1294 ( .A1(n36), .A2(n747), .B1(n33), .B2(n746), .ZN(n616) );
  OAI22_X1 U1295 ( .A1(n41), .A2(n732), .B1(n40), .B2(n731), .ZN(n602) );
  OAI22_X1 U1296 ( .A1(n24), .A2(n777), .B1(n22), .B2(n776), .ZN(n644) );
  OAI22_X1 U1297 ( .A1(n17), .A2(n796), .B1(n15), .B2(n795), .ZN(n662) );
  OAI22_X1 U1298 ( .A1(n6), .A2(n823), .B1(n822), .B2(n4), .ZN(n688) );
  OAI22_X1 U1299 ( .A1(n35), .A2(n748), .B1(n747), .B2(n33), .ZN(n617) );
  AND2_X1 U1300 ( .A1(n1065), .A2(n543), .ZN(n589) );
  OAI22_X1 U1301 ( .A1(n36), .A2(n739), .B1(n34), .B2(n738), .ZN(n608) );
  OAI22_X1 U1302 ( .A1(n48), .A2(n709), .B1(n46), .B2(n708), .ZN(n580) );
  OAI22_X1 U1303 ( .A1(n42), .A2(n724), .B1(n40), .B2(n723), .ZN(n594) );
  INV_X1 U1304 ( .A(n15), .ZN(n558) );
  NAND2_X1 U1305 ( .A1(n539), .A2(n540), .ZN(n291) );
  INV_X1 U1306 ( .A(n27), .ZN(n552) );
  OAI22_X1 U1307 ( .A1(n41), .A2(n879), .B1(n735), .B2(n39), .ZN(n567) );
  OR2_X1 U1308 ( .A1(n1064), .A2(n879), .ZN(n735) );
  OAI22_X1 U1309 ( .A1(n6), .A2(n827), .B1(n826), .B2(n4), .ZN(n692) );
  OAI22_X1 U1310 ( .A1(n24), .A2(n782), .B1(n21), .B2(n781), .ZN(n649) );
  AND2_X1 U1311 ( .A1(n1065), .A2(n549), .ZN(n621) );
  OR2_X1 U1312 ( .A1(n1064), .A2(n880), .ZN(n752) );
  OR2_X1 U1313 ( .A1(n1065), .A2(n882), .ZN(n786) );
  OR2_X1 U1314 ( .A1(n1065), .A2(n881), .ZN(n769) );
  AND2_X1 U1315 ( .A1(n1065), .A2(n564), .ZN(product[0]) );
  INV_X1 U1316 ( .A(n4), .ZN(n564) );
  INV_X1 U1317 ( .A(n33), .ZN(n549) );
  INV_X1 U1318 ( .A(n21), .ZN(n555) );
  INV_X1 U1319 ( .A(n45), .ZN(n543) );
  INV_X1 U1320 ( .A(n39), .ZN(n546) );
  OR2_X1 U1321 ( .A1(n1065), .A2(n884), .ZN(n820) );
  INV_X1 U1322 ( .A(n7), .ZN(n884) );
  BUF_X1 U1323 ( .A(n873), .Z(n28) );
  OAI22_X1 U1324 ( .A1(n6), .A2(n885), .B1(n837), .B2(n4), .ZN(n573) );
  OR2_X1 U1325 ( .A1(n1064), .A2(n885), .ZN(n837) );
  INV_X1 U1326 ( .A(n1), .ZN(n885) );
  OAI22_X1 U1327 ( .A1(n5), .A2(n836), .B1(n835), .B2(n4), .ZN(n701) );
  XNOR2_X1 U1328 ( .A(n13), .B(n842), .ZN(n791) );
  OAI22_X1 U1329 ( .A1(n23), .A2(n785), .B1(n21), .B2(n784), .ZN(n652) );
  OAI22_X1 U1330 ( .A1(n24), .A2(n882), .B1(n786), .B2(n22), .ZN(n570) );
  XNOR2_X1 U1331 ( .A(n13), .B(n838), .ZN(n787) );
  OAI22_X1 U1332 ( .A1(n5), .A2(n834), .B1(n833), .B2(n4), .ZN(n699) );
  OAI22_X1 U1333 ( .A1(n11), .A2(n819), .B1(n10), .B2(n818), .ZN(n684) );
  OAI22_X1 U1334 ( .A1(n35), .A2(n751), .B1(n33), .B2(n750), .ZN(n620) );
  OAI22_X1 U1335 ( .A1(n35), .A2(n880), .B1(n752), .B2(n34), .ZN(n568) );
  XNOR2_X1 U1336 ( .A(n13), .B(n847), .ZN(n796) );
  XNOR2_X1 U1337 ( .A(n13), .B(n846), .ZN(n795) );
  XNOR2_X1 U1338 ( .A(n13), .B(n839), .ZN(n788) );
  XNOR2_X1 U1339 ( .A(n13), .B(n844), .ZN(n793) );
  XNOR2_X1 U1340 ( .A(n13), .B(n1026), .ZN(n797) );
  XNOR2_X1 U1341 ( .A(n13), .B(n845), .ZN(n794) );
  XNOR2_X1 U1342 ( .A(n849), .B(n13), .ZN(n798) );
  XNOR2_X1 U1343 ( .A(n13), .B(n840), .ZN(n789) );
  XNOR2_X1 U1344 ( .A(n13), .B(n841), .ZN(n790) );
  XNOR2_X1 U1345 ( .A(n13), .B(n850), .ZN(n799) );
  XNOR2_X1 U1346 ( .A(n13), .B(n851), .ZN(n800) );
  XNOR2_X1 U1347 ( .A(n13), .B(n843), .ZN(n792) );
  XNOR2_X1 U1348 ( .A(n13), .B(n852), .ZN(n801) );
  BUF_X1 U1349 ( .A(n870), .Z(n45) );
  BUF_X1 U1350 ( .A(n870), .Z(n46) );
  BUF_X1 U1351 ( .A(n863), .Z(n42) );
  BUF_X1 U1352 ( .A(n864), .Z(n35) );
  BUF_X1 U1353 ( .A(n868), .Z(n11) );
  BUF_X1 U1354 ( .A(n869), .Z(n5) );
  XNOR2_X1 U1355 ( .A(n13), .B(n1064), .ZN(n802) );
  OAI22_X1 U1356 ( .A1(n30), .A2(n881), .B1(n769), .B2(n28), .ZN(n569) );
  INV_X1 U1357 ( .A(n31), .ZN(n880) );
  INV_X1 U1358 ( .A(n37), .ZN(n879) );
  INV_X1 U1359 ( .A(n19), .ZN(n882) );
  INV_X1 U1360 ( .A(n25), .ZN(n881) );
  INV_X1 U1361 ( .A(n43), .ZN(n878) );
  XNOR2_X1 U1362 ( .A(a[2]), .B(a[1]), .ZN(n876) );
  XNOR2_X1 U1363 ( .A(a[11]), .B(a[12]), .ZN(n871) );
  XNOR2_X1 U1364 ( .A(a[14]), .B(a[13]), .ZN(n870) );
  BUF_X2 U1365 ( .A(a[15]), .Z(n43) );
  NAND2_X1 U1366 ( .A1(n861), .A2(n877), .ZN(n869) );
  NAND2_X1 U1367 ( .A1(n860), .A2(n876), .ZN(n868) );
  NAND2_X1 U1368 ( .A1(n855), .A2(n871), .ZN(n863) );
  INV_X1 U1369 ( .A(a[0]), .ZN(n877) );
  XOR2_X1 U1370 ( .A(n80), .B(n292), .Z(product[4]) );
  AOI21_X1 U1371 ( .B1(n1009), .B2(n297), .A(n294), .ZN(n292) );
  BUF_X2 U1372 ( .A(n206), .Z(n51) );
  CLKBUF_X1 U1373 ( .A(n873), .Z(n27) );
  XNOR2_X1 U1374 ( .A(a[8]), .B(a[7]), .ZN(n873) );
  OAI22_X1 U1375 ( .A1(n36), .A2(n737), .B1(n34), .B2(n736), .ZN(n348) );
  INV_X1 U1376 ( .A(n348), .ZN(n349) );
  NAND2_X1 U1377 ( .A1(n858), .A2(n874), .ZN(n866) );
  XNOR2_X1 U1378 ( .A(a[5]), .B(a[6]), .ZN(n874) );
  INV_X1 U1379 ( .A(n1014), .ZN(n148) );
  NAND2_X1 U1380 ( .A1(n357), .A2(n364), .ZN(n169) );
  XOR2_X1 U1381 ( .A(n159), .B(n60), .Z(product[24]) );
  NAND2_X1 U1382 ( .A1(n854), .A2(n870), .ZN(n862) );
  BUF_X2 U1383 ( .A(n862), .Z(n48) );
  OAI22_X1 U1384 ( .A1(n41), .A2(n734), .B1(n39), .B2(n733), .ZN(n604) );
  INV_X1 U1385 ( .A(n182), .ZN(n180) );
  NAND2_X1 U1386 ( .A1(n365), .A2(n372), .ZN(n182) );
  NAND2_X1 U1387 ( .A1(n859), .A2(n875), .ZN(n867) );
  XNOR2_X1 U1388 ( .A(n7), .B(n841), .ZN(n807) );
  XNOR2_X1 U1389 ( .A(n7), .B(n845), .ZN(n811) );
  XNOR2_X1 U1390 ( .A(n7), .B(n847), .ZN(n813) );
  XNOR2_X1 U1391 ( .A(n7), .B(n846), .ZN(n812) );
  XNOR2_X1 U1392 ( .A(n7), .B(n842), .ZN(n808) );
  XNOR2_X1 U1393 ( .A(n7), .B(n840), .ZN(n806) );
  XNOR2_X1 U1394 ( .A(n7), .B(n850), .ZN(n816) );
  XNOR2_X1 U1395 ( .A(n7), .B(n849), .ZN(n815) );
  XNOR2_X1 U1396 ( .A(n7), .B(n844), .ZN(n810) );
  XNOR2_X1 U1397 ( .A(n7), .B(n1026), .ZN(n814) );
  XNOR2_X1 U1398 ( .A(n7), .B(n843), .ZN(n809) );
  XNOR2_X1 U1399 ( .A(n7), .B(n839), .ZN(n805) );
  XNOR2_X1 U1400 ( .A(n7), .B(n851), .ZN(n817) );
  XNOR2_X1 U1401 ( .A(n7), .B(n1064), .ZN(n819) );
  XNOR2_X1 U1402 ( .A(n7), .B(n852), .ZN(n818) );
  XNOR2_X1 U1403 ( .A(n7), .B(n838), .ZN(n804) );
  XNOR2_X1 U1404 ( .A(n25), .B(n838), .ZN(n753) );
  XNOR2_X1 U1405 ( .A(n25), .B(n1065), .ZN(n768) );
  XNOR2_X1 U1406 ( .A(n25), .B(n841), .ZN(n756) );
  XNOR2_X1 U1407 ( .A(n25), .B(n852), .ZN(n767) );
  XNOR2_X1 U1408 ( .A(n25), .B(n840), .ZN(n755) );
  XNOR2_X1 U1409 ( .A(n25), .B(n1036), .ZN(n762) );
  XNOR2_X1 U1410 ( .A(n25), .B(n839), .ZN(n754) );
  XNOR2_X1 U1411 ( .A(n25), .B(n848), .ZN(n763) );
  XNOR2_X1 U1412 ( .A(n25), .B(n846), .ZN(n761) );
  XNOR2_X1 U1413 ( .A(n25), .B(n845), .ZN(n760) );
  XNOR2_X1 U1414 ( .A(n25), .B(n844), .ZN(n759) );
  XNOR2_X1 U1415 ( .A(n849), .B(n25), .ZN(n764) );
  XNOR2_X1 U1416 ( .A(n25), .B(n843), .ZN(n758) );
  XNOR2_X1 U1417 ( .A(n25), .B(n851), .ZN(n766) );
  XNOR2_X1 U1418 ( .A(n25), .B(n842), .ZN(n757) );
  XNOR2_X1 U1419 ( .A(n25), .B(n850), .ZN(n765) );
  NOR2_X1 U1420 ( .A1(n218), .A2(n211), .ZN(n209) );
  XNOR2_X1 U1421 ( .A(n43), .B(n840), .ZN(n704) );
  XNOR2_X1 U1422 ( .A(n43), .B(n841), .ZN(n705) );
  XNOR2_X1 U1423 ( .A(n43), .B(n956), .ZN(n703) );
  XNOR2_X1 U1424 ( .A(n43), .B(n838), .ZN(n702) );
  XNOR2_X1 U1425 ( .A(n43), .B(n1033), .ZN(n707) );
  XNOR2_X1 U1426 ( .A(n43), .B(n842), .ZN(n706) );
  XNOR2_X1 U1427 ( .A(n43), .B(n844), .ZN(n708) );
  XNOR2_X1 U1428 ( .A(n43), .B(n1036), .ZN(n711) );
  XNOR2_X1 U1429 ( .A(n43), .B(n846), .ZN(n710) );
  XNOR2_X1 U1430 ( .A(n43), .B(n1064), .ZN(n717) );
  XNOR2_X1 U1431 ( .A(n43), .B(n845), .ZN(n709) );
  XNOR2_X1 U1432 ( .A(n43), .B(n850), .ZN(n714) );
  XNOR2_X1 U1433 ( .A(n43), .B(n849), .ZN(n713) );
  XNOR2_X1 U1434 ( .A(n43), .B(n848), .ZN(n712) );
  XNOR2_X1 U1435 ( .A(n43), .B(n852), .ZN(n716) );
  XNOR2_X1 U1436 ( .A(n43), .B(n851), .ZN(n715) );
  NAND2_X1 U1437 ( .A1(n503), .A2(n510), .ZN(n266) );
  NAND2_X1 U1438 ( .A1(n519), .A2(n524), .ZN(n275) );
  NOR2_X1 U1439 ( .A1(n519), .A2(n524), .ZN(n274) );
  XNOR2_X1 U1440 ( .A(n19), .B(n1065), .ZN(n785) );
  XNOR2_X1 U1441 ( .A(n19), .B(n852), .ZN(n784) );
  XNOR2_X1 U1442 ( .A(n19), .B(n848), .ZN(n780) );
  XNOR2_X1 U1443 ( .A(n19), .B(n846), .ZN(n778) );
  XNOR2_X1 U1444 ( .A(n19), .B(n1036), .ZN(n779) );
  XNOR2_X1 U1445 ( .A(n19), .B(n843), .ZN(n775) );
  XNOR2_X1 U1446 ( .A(n19), .B(n842), .ZN(n774) );
  XNOR2_X1 U1447 ( .A(n19), .B(n845), .ZN(n777) );
  XNOR2_X1 U1448 ( .A(n19), .B(n851), .ZN(n783) );
  XNOR2_X1 U1449 ( .A(n19), .B(n844), .ZN(n776) );
  XNOR2_X1 U1450 ( .A(n19), .B(n841), .ZN(n773) );
  XNOR2_X1 U1451 ( .A(n19), .B(n840), .ZN(n772) );
  XNOR2_X1 U1452 ( .A(n19), .B(n850), .ZN(n782) );
  XNOR2_X1 U1453 ( .A(n19), .B(n849), .ZN(n781) );
  XNOR2_X1 U1454 ( .A(n19), .B(n839), .ZN(n771) );
  XNOR2_X1 U1455 ( .A(n19), .B(n838), .ZN(n770) );
  NAND2_X1 U1456 ( .A1(n383), .A2(n392), .ZN(n200) );
  INV_X1 U1457 ( .A(n362), .ZN(n363) );
  OAI22_X1 U1458 ( .A1(n30), .A2(n754), .B1(n28), .B2(n753), .ZN(n362) );
  INV_X1 U1459 ( .A(n296), .ZN(n294) );
  OAI22_X1 U1460 ( .A1(n12), .A2(n884), .B1(n820), .B2(n10), .ZN(n572) );
  NAND2_X1 U1461 ( .A1(n511), .A2(n518), .ZN(n272) );
  OAI22_X1 U1462 ( .A1(n29), .A2(n763), .B1(n27), .B2(n762), .ZN(n631) );
  OAI22_X1 U1463 ( .A1(n29), .A2(n764), .B1(n27), .B2(n763), .ZN(n632) );
  OAI22_X1 U1464 ( .A1(n29), .A2(n768), .B1(n27), .B2(n767), .ZN(n636) );
  OAI22_X1 U1465 ( .A1(n29), .A2(n762), .B1(n27), .B2(n761), .ZN(n630) );
  OAI22_X1 U1466 ( .A1(n29), .A2(n767), .B1(n27), .B2(n766), .ZN(n635) );
  OAI22_X1 U1467 ( .A1(n29), .A2(n761), .B1(n27), .B2(n760), .ZN(n629) );
  OAI22_X1 U1468 ( .A1(n29), .A2(n766), .B1(n27), .B2(n765), .ZN(n634) );
  OAI21_X1 U1469 ( .B1(n254), .B2(n241), .A(n1030), .ZN(n240) );
  XNOR2_X1 U1470 ( .A(n31), .B(n840), .ZN(n738) );
  XNOR2_X1 U1471 ( .A(n31), .B(n1033), .ZN(n741) );
  XNOR2_X1 U1472 ( .A(n31), .B(n842), .ZN(n740) );
  XNOR2_X1 U1473 ( .A(n31), .B(n841), .ZN(n739) );
  XNOR2_X1 U1474 ( .A(n31), .B(n850), .ZN(n748) );
  XNOR2_X1 U1475 ( .A(n31), .B(n846), .ZN(n744) );
  XNOR2_X1 U1476 ( .A(n849), .B(n31), .ZN(n747) );
  XNOR2_X1 U1477 ( .A(n31), .B(n851), .ZN(n749) );
  XNOR2_X1 U1478 ( .A(n31), .B(n845), .ZN(n743) );
  XNOR2_X1 U1479 ( .A(n31), .B(n848), .ZN(n746) );
  XNOR2_X1 U1480 ( .A(n31), .B(n1064), .ZN(n751) );
  XNOR2_X1 U1481 ( .A(n31), .B(n844), .ZN(n742) );
  XNOR2_X1 U1482 ( .A(n31), .B(n847), .ZN(n745) );
  XNOR2_X1 U1483 ( .A(n31), .B(n852), .ZN(n750) );
  XNOR2_X1 U1484 ( .A(n31), .B(n956), .ZN(n737) );
  XNOR2_X1 U1485 ( .A(n31), .B(n838), .ZN(n736) );
  INV_X1 U1486 ( .A(n13), .ZN(n883) );
  OAI22_X1 U1487 ( .A1(n18), .A2(n802), .B1(n15), .B2(n801), .ZN(n668) );
  OAI22_X1 U1488 ( .A1(n18), .A2(n883), .B1(n803), .B2(n16), .ZN(n571) );
  OR2_X1 U1489 ( .A1(n1064), .A2(n883), .ZN(n803) );
  NOR2_X1 U1490 ( .A1(n241), .A2(n238), .ZN(n236) );
  XNOR2_X1 U1491 ( .A(n37), .B(n841), .ZN(n722) );
  XNOR2_X1 U1492 ( .A(n37), .B(n840), .ZN(n721) );
  XNOR2_X1 U1493 ( .A(n37), .B(n842), .ZN(n723) );
  XNOR2_X1 U1494 ( .A(n37), .B(n845), .ZN(n726) );
  XNOR2_X1 U1495 ( .A(n37), .B(n844), .ZN(n725) );
  XNOR2_X1 U1496 ( .A(n37), .B(n956), .ZN(n720) );
  XNOR2_X1 U1497 ( .A(n37), .B(n843), .ZN(n724) );
  XNOR2_X1 U1498 ( .A(n37), .B(n851), .ZN(n732) );
  XNOR2_X1 U1499 ( .A(n37), .B(n850), .ZN(n731) );
  XNOR2_X1 U1500 ( .A(n37), .B(n838), .ZN(n719) );
  XNOR2_X1 U1501 ( .A(n37), .B(n846), .ZN(n727) );
  XNOR2_X1 U1502 ( .A(n849), .B(n37), .ZN(n730) );
  XNOR2_X1 U1503 ( .A(n37), .B(n1064), .ZN(n734) );
  XNOR2_X1 U1504 ( .A(n848), .B(n37), .ZN(n729) );
  XNOR2_X1 U1505 ( .A(n37), .B(n1036), .ZN(n728) );
  XNOR2_X1 U1506 ( .A(n37), .B(n852), .ZN(n733) );
  XNOR2_X1 U1507 ( .A(n247), .B(n71), .ZN(product[13]) );
  OAI21_X1 U1508 ( .B1(n254), .B2(n248), .A(n253), .ZN(n247) );
  NOR2_X1 U1509 ( .A1(n1062), .A2(n87), .ZN(n85) );
  XOR2_X1 U1510 ( .A(n93), .B(n54), .Z(product[30]) );
  NOR2_X1 U1511 ( .A1(n1062), .A2(n144), .ZN(n140) );
  NOR2_X1 U1512 ( .A1(n1062), .A2(n133), .ZN(n131) );
  NOR2_X1 U1513 ( .A1(n1062), .A2(n109), .ZN(n107) );
  NOR2_X1 U1514 ( .A1(n1062), .A2(n124), .ZN(n118) );
  NOR2_X1 U1515 ( .A1(n1062), .A2(n96), .ZN(n94) );
  XNOR2_X1 U1516 ( .A(n1), .B(n845), .ZN(n828) );
  XNOR2_X1 U1517 ( .A(n1), .B(n840), .ZN(n823) );
  XNOR2_X1 U1518 ( .A(n1), .B(n848), .ZN(n831) );
  XNOR2_X1 U1519 ( .A(n1), .B(n846), .ZN(n829) );
  XNOR2_X1 U1520 ( .A(n1), .B(n847), .ZN(n830) );
  XNOR2_X1 U1521 ( .A(n1), .B(n844), .ZN(n827) );
  XNOR2_X1 U1522 ( .A(n1), .B(n841), .ZN(n824) );
  XNOR2_X1 U1523 ( .A(n1), .B(n839), .ZN(n822) );
  XNOR2_X1 U1524 ( .A(n1), .B(n849), .ZN(n832) );
  XNOR2_X1 U1525 ( .A(n1), .B(n843), .ZN(n826) );
  XNOR2_X1 U1526 ( .A(n1), .B(n842), .ZN(n825) );
  XNOR2_X1 U1527 ( .A(n1), .B(n1065), .ZN(n836) );
  XNOR2_X1 U1528 ( .A(n1), .B(n852), .ZN(n835) );
  XNOR2_X1 U1529 ( .A(n1), .B(n851), .ZN(n834) );
  XNOR2_X1 U1530 ( .A(n1), .B(n850), .ZN(n833) );
  XNOR2_X1 U1531 ( .A(n1), .B(n838), .ZN(n821) );
  AOI21_X1 U1532 ( .B1(n281), .B2(n1011), .A(n278), .ZN(n276) );
  OAI22_X1 U1533 ( .A1(n29), .A2(n765), .B1(n27), .B2(n764), .ZN(n633) );
  OAI21_X1 U1534 ( .B1(n242), .B2(n238), .A(n239), .ZN(n237) );
  NAND2_X1 U1535 ( .A1(n857), .A2(n873), .ZN(n865) );
  XNOR2_X1 U1536 ( .A(n234), .B(n69), .ZN(product[15]) );
  AOI21_X1 U1537 ( .B1(n214), .B2(n234), .A(n215), .ZN(n213) );
  AOI21_X1 U1538 ( .B1(n234), .B2(n317), .A(n231), .ZN(n229) );
  AOI21_X1 U1539 ( .B1(n234), .B2(n1060), .A(n222), .ZN(n220) );
  NAND2_X1 U1540 ( .A1(n209), .A2(n225), .ZN(n207) );
  OAI21_X1 U1541 ( .B1(n227), .B2(n233), .A(n228), .ZN(n226) );
  NOR2_X1 U1542 ( .A1(n1057), .A2(n232), .ZN(n225) );
  INV_X1 U1543 ( .A(n1061), .ZN(n234) );
  AOI21_X1 U1544 ( .B1(n209), .B2(n226), .A(n210), .ZN(n208) );
  OAI21_X1 U1545 ( .B1(n219), .B2(n1041), .A(n212), .ZN(n210) );
  OAI21_X1 U1546 ( .B1(n1021), .B2(n87), .A(n88), .ZN(n86) );
  OAI21_X1 U1547 ( .B1(n1013), .B2(n133), .A(n134), .ZN(n132) );
  OAI21_X1 U1548 ( .B1(n1014), .B2(n144), .A(n145), .ZN(n141) );
  OAI21_X1 U1549 ( .B1(n150), .B2(n109), .A(n110), .ZN(n108) );
  OAI21_X1 U1550 ( .B1(n1013), .B2(n96), .A(n97), .ZN(n95) );
  OAI21_X1 U1551 ( .B1(n150), .B2(n124), .A(n125), .ZN(n119) );
  OAI21_X1 U1552 ( .B1(n153), .B2(n191), .A(n154), .ZN(n152) );
  OAI21_X1 U1553 ( .B1(n157), .B2(n169), .A(n158), .ZN(n156) );
  XOR2_X1 U1554 ( .A(a[14]), .B(a[15]), .Z(n854) );
  XNOR2_X1 U1555 ( .A(a[9]), .B(a[10]), .ZN(n872) );
  XOR2_X1 U1556 ( .A(a[8]), .B(a[9]), .Z(n857) );
  AOI21_X1 U1557 ( .B1(n155), .B2(n180), .A(n156), .ZN(n154) );
  NAND2_X1 U1558 ( .A1(n1032), .A2(n155), .ZN(n153) );
  XOR2_X1 U1559 ( .A(a[6]), .B(a[7]), .Z(n858) );
  OAI21_X1 U1560 ( .B1(n207), .B2(n235), .A(n208), .ZN(n206) );
  AOI21_X1 U1561 ( .B1(n236), .B2(n255), .A(n237), .ZN(n235) );
  XOR2_X1 U1562 ( .A(a[12]), .B(a[13]), .Z(n855) );
  NOR2_X1 U1563 ( .A1(n168), .A2(n157), .ZN(n155) );
  NAND2_X1 U1564 ( .A1(n856), .A2(n872), .ZN(n864) );
  OAI21_X1 U1565 ( .B1(n256), .B2(n268), .A(n257), .ZN(n255) );
  XOR2_X1 U1566 ( .A(a[10]), .B(a[11]), .Z(n856) );
  INV_X1 U1567 ( .A(n1062), .ZN(n147) );
  NOR2_X1 U1568 ( .A1(n204), .A2(n199), .ZN(n197) );
  INV_X1 U1569 ( .A(n204), .ZN(n313) );
  NOR2_X1 U1570 ( .A1(n393), .A2(n404), .ZN(n204) );
  AOI21_X1 U1571 ( .B1(n1039), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U1572 ( .B1(n51), .B2(n131), .A(n132), .ZN(n130) );
  AOI21_X1 U1573 ( .B1(n1039), .B2(n94), .A(n95), .ZN(n93) );
  AOI21_X1 U1574 ( .B1(n1039), .B2(n118), .A(n119), .ZN(n117) );
  AOI21_X1 U1575 ( .B1(n1039), .B2(n140), .A(n141), .ZN(n139) );
  AOI21_X1 U1576 ( .B1(n1039), .B2(n107), .A(n108), .ZN(n106) );
  AOI21_X1 U1577 ( .B1(n1039), .B2(n160), .A(n161), .ZN(n159) );
  AOI21_X1 U1578 ( .B1(n51), .B2(n147), .A(n148), .ZN(n146) );
  XNOR2_X1 U1579 ( .A(n1039), .B(n65), .ZN(product[19]) );
  AOI21_X1 U1580 ( .B1(n51), .B2(n313), .A(n203), .ZN(n201) );
  AOI21_X1 U1581 ( .B1(n51), .B2(n171), .A(n172), .ZN(n170) );
  AOI21_X1 U1582 ( .B1(n51), .B2(n184), .A(n185), .ZN(n183) );
  AOI21_X1 U1583 ( .B1(n51), .B2(n193), .A(n198), .ZN(n192) );
  XNOR2_X1 U1584 ( .A(n1027), .B(n75), .ZN(product[9]) );
  NAND2_X1 U1585 ( .A1(n541), .A2(n572), .ZN(n296) );
  XNOR2_X1 U1586 ( .A(a[3]), .B(a[4]), .ZN(n875) );
  XOR2_X1 U1587 ( .A(a[3]), .B(a[2]), .Z(n860) );
  XOR2_X1 U1588 ( .A(a[0]), .B(a[1]), .Z(n861) );
  XOR2_X1 U1589 ( .A(n276), .B(n76), .Z(product[8]) );
  XOR2_X1 U1590 ( .A(a[4]), .B(a[5]), .Z(n859) );
  XNOR2_X1 U1591 ( .A(n281), .B(n77), .ZN(product[7]) );
  XOR2_X1 U1592 ( .A(n78), .B(n284), .Z(product[6]) );
endmodule


module datapath_DW_mult_tc_11 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n4, n5, n6, n7, n9, n10, n11, n12, n13, n15, n16, n17, n18, n19,
         n21, n22, n23, n24, n25, n27, n29, n30, n31, n33, n34, n35, n36, n37,
         n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n51, n54, n55, n56,
         n57, n58, n59, n61, n65, n67, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n84, n85, n86, n87, n88, n90, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n103, n105, n106, n107,
         n108, n109, n110, n114, n116, n117, n118, n119, n122, n123, n124,
         n125, n127, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n143, n144, n145, n146, n147, n148, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n180, n182, n183, n184, n185,
         n188, n189, n190, n191, n192, n194, n195, n196, n197, n198, n199,
         n200, n201, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n246, n247, n248,
         n249, n251, n253, n254, n255, n256, n257, n259, n261, n262, n264,
         n266, n267, n268, n270, n272, n273, n274, n275, n276, n278, n280,
         n281, n282, n283, n284, n286, n288, n289, n290, n291, n292, n294,
         n296, n297, n298, n299, n301, n306, n308, n312, n313, n314, n316,
         n317, n318, n324, n326, n328, n330, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n545, n546,
         n548, n549, n551, n552, n554, n555, n557, n558, n560, n561, n563,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1010, n1011, n1012, n1013, n1014;
  assign product[31] = n84;

  FA_X1 U364 ( .A(n575), .B(n338), .CI(n590), .CO(n334), .S(n335) );
  FA_X1 U365 ( .A(n339), .B(n576), .CI(n342), .CO(n336), .S(n337) );
  FA_X1 U367 ( .A(n346), .B(n577), .CI(n343), .CO(n340), .S(n341) );
  FA_X1 U368 ( .A(n591), .B(n348), .CI(n606), .CO(n342), .S(n343) );
  FA_X1 U369 ( .A(n347), .B(n354), .CI(n352), .CO(n344), .S(n345) );
  FA_X1 U370 ( .A(n578), .B(n592), .CI(n349), .CO(n346), .S(n347) );
  FA_X1 U372 ( .A(n358), .B(n355), .CI(n353), .CO(n350), .S(n351) );
  FA_X1 U373 ( .A(n362), .B(n607), .CI(n360), .CO(n352), .S(n353) );
  FA_X1 U374 ( .A(n593), .B(n579), .CI(n622), .CO(n354), .S(n355) );
  FA_X1 U375 ( .A(n359), .B(n361), .CI(n366), .CO(n356), .S(n357) );
  FA_X1 U376 ( .A(n370), .B(n363), .CI(n368), .CO(n358), .S(n359) );
  FA_X1 U377 ( .A(n580), .B(n594), .CI(n608), .CO(n360), .S(n361) );
  FA_X1 U379 ( .A(n374), .B(n376), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U380 ( .A(n369), .B(n378), .CI(n371), .CO(n366), .S(n367) );
  FA_X1 U381 ( .A(n595), .B(n609), .CI(n380), .CO(n368), .S(n369) );
  FA_X1 U382 ( .A(n623), .B(n581), .CI(n638), .CO(n370), .S(n371) );
  FA_X1 U383 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  FA_X1 U384 ( .A(n379), .B(n388), .CI(n386), .CO(n374), .S(n375) );
  FA_X1 U385 ( .A(n381), .B(n610), .CI(n390), .CO(n376), .S(n377) );
  FA_X1 U386 ( .A(n624), .B(n596), .CI(n582), .CO(n378), .S(n379) );
  FA_X1 U388 ( .A(n394), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U389 ( .A(n391), .B(n389), .CI(n396), .CO(n384), .S(n385) );
  FA_X1 U390 ( .A(n400), .B(n625), .CI(n398), .CO(n386), .S(n387) );
  FA_X1 U391 ( .A(n597), .B(n639), .CI(n611), .CO(n388), .S(n389) );
  FA_X1 U392 ( .A(n402), .B(n583), .CI(n654), .CO(n390), .S(n391) );
  FA_X1 U393 ( .A(n406), .B(n397), .CI(n395), .CO(n392), .S(n393) );
  FA_X1 U394 ( .A(n410), .B(n399), .CI(n408), .CO(n394), .S(n395) );
  FA_X1 U395 ( .A(n412), .B(n414), .CI(n401), .CO(n396), .S(n397) );
  FA_X1 U396 ( .A(n584), .B(n598), .CI(n403), .CO(n398), .S(n399) );
  FA_X1 U397 ( .A(n640), .B(n626), .CI(n612), .CO(n400), .S(n401) );
  FA_X1 U399 ( .A(n418), .B(n409), .CI(n407), .CO(n404), .S(n405) );
  FA_X1 U400 ( .A(n411), .B(n422), .CI(n420), .CO(n406), .S(n407) );
  FA_X1 U401 ( .A(n413), .B(n424), .CI(n415), .CO(n408), .S(n409) );
  FA_X1 U403 ( .A(n599), .B(n655), .CI(n641), .CO(n412), .S(n413) );
  FA_X1 U404 ( .A(n428), .B(n585), .CI(n670), .CO(n414), .S(n415) );
  FA_X1 U405 ( .A(n432), .B(n421), .CI(n419), .CO(n416), .S(n417) );
  FA_X1 U406 ( .A(n423), .B(n436), .CI(n434), .CO(n418), .S(n419) );
  FA_X1 U407 ( .A(n425), .B(n438), .CI(n427), .CO(n420), .S(n421) );
  FA_X1 U408 ( .A(n442), .B(n429), .CI(n440), .CO(n422), .S(n423) );
  FA_X1 U409 ( .A(n628), .B(n642), .CI(n600), .CO(n424), .S(n425) );
  FA_X1 U410 ( .A(n656), .B(n614), .CI(n586), .CO(n426), .S(n427) );
  FA_X1 U412 ( .A(n446), .B(n435), .CI(n433), .CO(n430), .S(n431) );
  FA_X1 U413 ( .A(n448), .B(n450), .CI(n437), .CO(n432), .S(n433) );
  FA_X1 U414 ( .A(n439), .B(n452), .CI(n441), .CO(n434), .S(n435) );
  FA_X1 U415 ( .A(n443), .B(n456), .CI(n454), .CO(n436), .S(n437) );
  FA_X1 U416 ( .A(n615), .B(n671), .CI(n657), .CO(n438), .S(n439) );
  FA_X1 U417 ( .A(n587), .B(n629), .CI(n686), .CO(n440), .S(n441) );
  FA_X1 U420 ( .A(n449), .B(n460), .CI(n447), .CO(n444), .S(n445) );
  FA_X1 U421 ( .A(n462), .B(n455), .CI(n451), .CO(n446), .S(n447) );
  FA_X1 U422 ( .A(n464), .B(n466), .CI(n453), .CO(n448), .S(n449) );
  FA_X1 U423 ( .A(n457), .B(n672), .CI(n468), .CO(n450), .S(n451) );
  FA_X1 U424 ( .A(n687), .B(n630), .CI(n658), .CO(n452), .S(n453) );
  FA_X1 U425 ( .A(n602), .B(n644), .CI(n616), .CO(n454), .S(n455) );
  HA_X1 U426 ( .A(n566), .B(n588), .CO(n456), .S(n457) );
  FA_X1 U427 ( .A(n463), .B(n472), .CI(n461), .CO(n458), .S(n459) );
  FA_X1 U428 ( .A(n465), .B(n467), .CI(n474), .CO(n460), .S(n461) );
  FA_X1 U429 ( .A(n476), .B(n478), .CI(n469), .CO(n462), .S(n463) );
  FA_X1 U430 ( .A(n645), .B(n659), .CI(n480), .CO(n464), .S(n465) );
  FA_X1 U431 ( .A(n603), .B(n673), .CI(n631), .CO(n466), .S(n467) );
  FA_X1 U432 ( .A(n617), .B(n589), .CI(n688), .CO(n468), .S(n469) );
  FA_X1 U433 ( .A(n484), .B(n475), .CI(n473), .CO(n470), .S(n471) );
  FA_X1 U434 ( .A(n479), .B(n477), .CI(n486), .CO(n472), .S(n473) );
  FA_X1 U435 ( .A(n490), .B(n481), .CI(n488), .CO(n474), .S(n475) );
  FA_X1 U436 ( .A(n618), .B(n632), .CI(n660), .CO(n476), .S(n477) );
  FA_X1 U437 ( .A(n689), .B(n646), .CI(n674), .CO(n478), .S(n479) );
  HA_X1 U438 ( .A(n604), .B(n567), .CO(n480), .S(n481) );
  FA_X1 U439 ( .A(n487), .B(n494), .CI(n485), .CO(n482), .S(n483) );
  FA_X1 U440 ( .A(n489), .B(n491), .CI(n496), .CO(n484), .S(n485) );
  FA_X1 U441 ( .A(n500), .B(n661), .CI(n498), .CO(n486), .S(n487) );
  FA_X1 U442 ( .A(n619), .B(n675), .CI(n647), .CO(n488), .S(n489) );
  FA_X1 U443 ( .A(n633), .B(n605), .CI(n690), .CO(n490), .S(n491) );
  FA_X1 U444 ( .A(n504), .B(n497), .CI(n495), .CO(n492), .S(n493) );
  FA_X1 U445 ( .A(n506), .B(n508), .CI(n499), .CO(n494), .S(n495) );
  FA_X1 U446 ( .A(n648), .B(n676), .CI(n501), .CO(n496), .S(n497) );
  FA_X1 U449 ( .A(n512), .B(n507), .CI(n505), .CO(n502), .S(n503) );
  FA_X1 U450 ( .A(n514), .B(n516), .CI(n509), .CO(n504), .S(n505) );
  FA_X1 U451 ( .A(n635), .B(n677), .CI(n663), .CO(n506), .S(n507) );
  FA_X1 U452 ( .A(n649), .B(n621), .CI(n692), .CO(n508), .S(n509) );
  FA_X1 U453 ( .A(n515), .B(n520), .CI(n513), .CO(n510), .S(n511) );
  FA_X1 U454 ( .A(n517), .B(n693), .CI(n522), .CO(n512), .S(n513) );
  FA_X1 U455 ( .A(n650), .B(n664), .CI(n678), .CO(n514), .S(n515) );
  HA_X1 U456 ( .A(n569), .B(n636), .CO(n516), .S(n517) );
  FA_X1 U457 ( .A(n523), .B(n526), .CI(n521), .CO(n518), .S(n519) );
  FA_X1 U458 ( .A(n651), .B(n679), .CI(n528), .CO(n520), .S(n521) );
  FA_X1 U459 ( .A(n665), .B(n637), .CI(n694), .CO(n522), .S(n523) );
  FA_X1 U460 ( .A(n532), .B(n529), .CI(n527), .CO(n524), .S(n525) );
  FA_X1 U461 ( .A(n666), .B(n695), .CI(n680), .CO(n526), .S(n527) );
  HA_X1 U462 ( .A(n570), .B(n652), .CO(n528), .S(n529) );
  FA_X1 U463 ( .A(n536), .B(n667), .CI(n533), .CO(n530), .S(n531) );
  FA_X1 U464 ( .A(n696), .B(n653), .CI(n681), .CO(n532), .S(n533) );
  FA_X1 U465 ( .A(n682), .B(n697), .CI(n537), .CO(n534), .S(n535) );
  HA_X1 U466 ( .A(n571), .B(n668), .CO(n536), .S(n537) );
  FA_X1 U467 ( .A(n698), .B(n669), .CI(n683), .CO(n538), .S(n539) );
  HA_X1 U468 ( .A(n684), .B(n699), .CO(n540), .S(n541) );
  BUF_X1 U822 ( .A(b[15]), .Z(n953) );
  BUF_X1 U823 ( .A(n234), .Z(n986) );
  CLKBUF_X2 U824 ( .A(b[4]), .Z(n849) );
  CLKBUF_X3 U825 ( .A(n865), .Z(n29) );
  CLKBUF_X1 U826 ( .A(n276), .Z(n954) );
  NOR2_X2 U827 ( .A1(n373), .A2(n382), .ZN(n190) );
  CLKBUF_X3 U828 ( .A(n864), .Z(n36) );
  CLKBUF_X3 U829 ( .A(n49), .Z(n1012) );
  AOI21_X2 U830 ( .B1(n972), .B2(n289), .A(n286), .ZN(n284) );
  BUF_X2 U831 ( .A(n864), .Z(n35) );
  BUF_X4 U832 ( .A(a[11]), .Z(n31) );
  INV_X1 U833 ( .A(n879), .ZN(n955) );
  CLKBUF_X3 U834 ( .A(a[13]), .Z(n37) );
  BUF_X2 U835 ( .A(n871), .Z(n39) );
  XOR2_X1 U836 ( .A(n568), .B(n620), .Z(n501) );
  INV_X1 U837 ( .A(n956), .ZN(n500) );
  NAND2_X1 U838 ( .A1(n568), .A2(n620), .ZN(n956) );
  XOR2_X1 U839 ( .A(n613), .B(n627), .Z(n957) );
  XOR2_X1 U840 ( .A(n426), .B(n957), .Z(n411) );
  NAND2_X1 U841 ( .A1(n426), .A2(n613), .ZN(n958) );
  NAND2_X1 U842 ( .A1(n426), .A2(n627), .ZN(n959) );
  NAND2_X1 U843 ( .A1(n613), .A2(n627), .ZN(n960) );
  NAND3_X1 U844 ( .A1(n958), .A2(n959), .A3(n960), .ZN(n410) );
  CLKBUF_X1 U845 ( .A(n842), .Z(n961) );
  BUF_X1 U846 ( .A(n842), .Z(n962) );
  BUF_X2 U847 ( .A(n842), .Z(n963) );
  BUF_X1 U848 ( .A(b[11]), .Z(n842) );
  BUF_X2 U849 ( .A(n867), .Z(n17) );
  BUF_X1 U850 ( .A(b[0]), .Z(n49) );
  BUF_X1 U851 ( .A(b[7]), .Z(n846) );
  BUF_X1 U852 ( .A(b[15]), .Z(n838) );
  BUF_X2 U853 ( .A(n863), .Z(n41) );
  BUF_X2 U854 ( .A(n871), .Z(n40) );
  NAND2_X1 U855 ( .A1(n198), .A2(n151), .ZN(n964) );
  INV_X1 U856 ( .A(n152), .ZN(n965) );
  AND2_X2 U857 ( .A1(n964), .A2(n965), .ZN(n150) );
  AND2_X1 U858 ( .A1(n471), .A2(n482), .ZN(n1001) );
  OAI22_X1 U859 ( .A1(n6), .A2(n826), .B1(n825), .B2(n4), .ZN(n691) );
  BUF_X2 U860 ( .A(n867), .Z(n18) );
  OAI22_X1 U861 ( .A1(n48), .A2(n703), .B1(n46), .B2(n702), .ZN(n332) );
  BUF_X1 U862 ( .A(n206), .Z(n1007) );
  INV_X1 U863 ( .A(n1001), .ZN(n246) );
  OR2_X1 U864 ( .A1(n503), .A2(n510), .ZN(n966) );
  OR2_X1 U865 ( .A1(n337), .A2(n340), .ZN(n967) );
  OR2_X1 U866 ( .A1(n334), .A2(n333), .ZN(n968) );
  OR2_X1 U867 ( .A1(n574), .A2(n332), .ZN(n969) );
  OR2_X1 U868 ( .A1(n483), .A2(n492), .ZN(n970) );
  OR2_X1 U869 ( .A1(n493), .A2(n502), .ZN(n971) );
  OR2_X1 U870 ( .A1(n535), .A2(n538), .ZN(n972) );
  OR2_X1 U871 ( .A1(n541), .A2(n572), .ZN(n973) );
  OR2_X1 U872 ( .A1(n365), .A2(n372), .ZN(n974) );
  OR2_X1 U873 ( .A1(n336), .A2(n335), .ZN(n975) );
  OR2_X1 U874 ( .A1(n525), .A2(n530), .ZN(n976) );
  OR2_X1 U875 ( .A1(n511), .A2(n518), .ZN(n977) );
  NOR2_X1 U876 ( .A1(n357), .A2(n364), .ZN(n168) );
  OR2_X1 U877 ( .A1(n701), .A2(n573), .ZN(n978) );
  CLKBUF_X2 U878 ( .A(b[1]), .Z(n852) );
  CLKBUF_X1 U879 ( .A(n251), .Z(n979) );
  NOR2_X1 U880 ( .A1(n405), .A2(n416), .ZN(n980) );
  XOR2_X1 U881 ( .A(n691), .B(n662), .Z(n981) );
  XOR2_X1 U882 ( .A(n634), .B(n981), .Z(n499) );
  NAND2_X1 U883 ( .A1(n634), .A2(n691), .ZN(n982) );
  NAND2_X1 U884 ( .A1(n634), .A2(n662), .ZN(n983) );
  NAND2_X1 U885 ( .A1(n691), .A2(n662), .ZN(n984) );
  NAND3_X1 U886 ( .A1(n982), .A2(n983), .A3(n984), .ZN(n498) );
  BUF_X1 U887 ( .A(n206), .Z(n51) );
  BUF_X2 U888 ( .A(n49), .Z(n1014) );
  CLKBUF_X2 U889 ( .A(b[12]), .Z(n841) );
  BUF_X1 U890 ( .A(n206), .Z(n1011) );
  BUF_X2 U891 ( .A(n869), .Z(n6) );
  BUF_X4 U892 ( .A(a[5]), .Z(n13) );
  BUF_X2 U893 ( .A(n873), .Z(n27) );
  BUF_X1 U894 ( .A(b[9]), .Z(n844) );
  BUF_X2 U895 ( .A(n863), .Z(n42) );
  BUF_X1 U896 ( .A(n206), .Z(n1010) );
  XNOR2_X1 U897 ( .A(n201), .B(n985), .ZN(product[20]) );
  AND2_X1 U898 ( .A1(n312), .A2(n200), .ZN(n985) );
  XNOR2_X1 U899 ( .A(n213), .B(n987), .ZN(product[18]) );
  AND2_X1 U900 ( .A1(n314), .A2(n212), .ZN(n987) );
  XNOR2_X1 U901 ( .A(n159), .B(n988), .ZN(product[24]) );
  AND2_X1 U902 ( .A1(n308), .A2(n158), .ZN(n988) );
  XNOR2_X1 U903 ( .A(n183), .B(n989), .ZN(product[22]) );
  AND2_X1 U904 ( .A1(n175), .A2(n182), .ZN(n989) );
  XNOR2_X1 U905 ( .A(n192), .B(n990), .ZN(product[21]) );
  AND2_X1 U906 ( .A1(n188), .A2(n191), .ZN(n990) );
  XNOR2_X1 U907 ( .A(n1), .B(n963), .ZN(n991) );
  BUF_X1 U908 ( .A(b[3]), .Z(n850) );
  BUF_X2 U909 ( .A(n839), .Z(n992) );
  CLKBUF_X1 U910 ( .A(b[14]), .Z(n839) );
  NOR2_X1 U911 ( .A1(n431), .A2(n444), .ZN(n993) );
  BUF_X1 U912 ( .A(n844), .Z(n994) );
  BUF_X1 U913 ( .A(n844), .Z(n995) );
  BUF_X1 U914 ( .A(n844), .Z(n996) );
  BUF_X1 U915 ( .A(n845), .Z(n997) );
  BUF_X1 U916 ( .A(n845), .Z(n998) );
  BUF_X1 U917 ( .A(n845), .Z(n999) );
  CLKBUF_X1 U918 ( .A(b[8]), .Z(n845) );
  AOI21_X1 U919 ( .B1(n1002), .B2(n979), .A(n1001), .ZN(n1000) );
  CLKBUF_X2 U920 ( .A(b[5]), .Z(n848) );
  OR2_X2 U921 ( .A1(n471), .A2(n482), .ZN(n1002) );
  BUF_X1 U922 ( .A(b[2]), .Z(n851) );
  CLKBUF_X2 U923 ( .A(b[10]), .Z(n843) );
  NAND2_X1 U924 ( .A1(n25), .A2(n850), .ZN(n1004) );
  NAND2_X1 U925 ( .A1(n881), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U926 ( .A1(n1004), .A2(n1005), .ZN(n765) );
  INV_X1 U927 ( .A(n850), .ZN(n1003) );
  BUF_X4 U928 ( .A(a[9]), .Z(n25) );
  XNOR2_X1 U929 ( .A(n229), .B(n1006), .ZN(product[16]) );
  AND2_X1 U930 ( .A1(n316), .A2(n228), .ZN(n1006) );
  BUF_X2 U931 ( .A(b[6]), .Z(n847) );
  NAND2_X1 U932 ( .A1(n197), .A2(n151), .ZN(n1008) );
  NOR2_X1 U933 ( .A1(n345), .A2(n350), .ZN(n144) );
  NOR2_X1 U934 ( .A1(n351), .A2(n356), .ZN(n157) );
  NOR2_X1 U935 ( .A1(n341), .A2(n344), .ZN(n137) );
  NOR2_X1 U936 ( .A1(n531), .A2(n534), .ZN(n282) );
  AND2_X1 U937 ( .A1(n978), .A2(n301), .ZN(product[1]) );
  BUF_X1 U938 ( .A(n49), .Z(n1013) );
  INV_X1 U939 ( .A(n224), .ZN(n222) );
  INV_X1 U940 ( .A(n223), .ZN(n221) );
  INV_X1 U941 ( .A(n226), .ZN(n224) );
  INV_X1 U942 ( .A(n225), .ZN(n223) );
  INV_X1 U943 ( .A(n177), .ZN(n175) );
  NOR2_X1 U944 ( .A1(n195), .A2(n162), .ZN(n160) );
  NOR2_X1 U945 ( .A1(n195), .A2(n173), .ZN(n171) );
  NOR2_X1 U946 ( .A1(n195), .A2(n190), .ZN(n184) );
  INV_X1 U947 ( .A(n196), .ZN(n194) );
  INV_X1 U948 ( .A(n98), .ZN(n96) );
  INV_X1 U949 ( .A(n1008), .ZN(n147) );
  INV_X1 U950 ( .A(n198), .ZN(n196) );
  NAND2_X1 U951 ( .A1(n313), .A2(n205), .ZN(n65) );
  INV_X1 U952 ( .A(n204), .ZN(n313) );
  NAND2_X1 U953 ( .A1(n217), .A2(n219), .ZN(n67) );
  INV_X1 U954 ( .A(n211), .ZN(n314) );
  NOR2_X1 U955 ( .A1(n177), .A2(n166), .ZN(n164) );
  NOR2_X1 U956 ( .A1(n124), .A2(n100), .ZN(n98) );
  OAI21_X1 U957 ( .B1(n196), .B2(n173), .A(n174), .ZN(n172) );
  AOI21_X1 U958 ( .B1(n189), .B2(n175), .A(n176), .ZN(n174) );
  INV_X1 U959 ( .A(n178), .ZN(n176) );
  NOR2_X1 U960 ( .A1(n227), .A2(n232), .ZN(n225) );
  XNOR2_X1 U961 ( .A(n240), .B(n70), .ZN(product[14]) );
  NAND2_X1 U962 ( .A1(n318), .A2(n239), .ZN(n70) );
  XNOR2_X1 U963 ( .A(n986), .B(n69), .ZN(product[15]) );
  NAND2_X1 U964 ( .A1(n317), .A2(n233), .ZN(n69) );
  INV_X1 U965 ( .A(n232), .ZN(n317) );
  INV_X1 U966 ( .A(n197), .ZN(n195) );
  NOR2_X1 U967 ( .A1(n218), .A2(n211), .ZN(n209) );
  NAND2_X1 U968 ( .A1(n155), .A2(n974), .ZN(n153) );
  INV_X1 U969 ( .A(n268), .ZN(n267) );
  OAI21_X1 U970 ( .B1(n196), .B2(n190), .A(n191), .ZN(n185) );
  NAND2_X1 U971 ( .A1(n164), .A2(n188), .ZN(n162) );
  NAND2_X1 U972 ( .A1(n188), .A2(n175), .ZN(n173) );
  INV_X1 U973 ( .A(n974), .ZN(n177) );
  INV_X1 U974 ( .A(n124), .ZN(n122) );
  NAND2_X1 U975 ( .A1(n1002), .A2(n970), .ZN(n241) );
  INV_X1 U976 ( .A(n180), .ZN(n178) );
  INV_X1 U977 ( .A(n217), .ZN(n216) );
  INV_X1 U978 ( .A(n979), .ZN(n249) );
  NAND2_X1 U979 ( .A1(n122), .A2(n975), .ZN(n109) );
  INV_X1 U980 ( .A(n970), .ZN(n248) );
  INV_X1 U981 ( .A(n205), .ZN(n203) );
  INV_X1 U982 ( .A(n233), .ZN(n231) );
  NOR2_X1 U983 ( .A1(n405), .A2(n416), .ZN(n211) );
  NAND2_X1 U984 ( .A1(n143), .A2(n145), .ZN(n59) );
  INV_X1 U985 ( .A(n199), .ZN(n312) );
  NAND2_X1 U986 ( .A1(n324), .A2(n275), .ZN(n76) );
  INV_X1 U987 ( .A(n274), .ZN(n324) );
  NOR2_X1 U988 ( .A1(n204), .A2(n199), .ZN(n197) );
  AOI21_X1 U989 ( .B1(n971), .B2(n264), .A(n259), .ZN(n257) );
  NAND2_X1 U990 ( .A1(n971), .A2(n966), .ZN(n256) );
  INV_X1 U991 ( .A(n261), .ZN(n259) );
  OAI21_X1 U992 ( .B1(n153), .B2(n191), .A(n154), .ZN(n152) );
  AOI21_X1 U993 ( .B1(n155), .B2(n180), .A(n156), .ZN(n154) );
  AOI21_X1 U994 ( .B1(n273), .B2(n977), .A(n270), .ZN(n268) );
  INV_X1 U995 ( .A(n272), .ZN(n270) );
  NOR2_X1 U996 ( .A1(n417), .A2(n430), .ZN(n218) );
  INV_X1 U997 ( .A(n190), .ZN(n188) );
  OAI21_X1 U998 ( .B1(n276), .B2(n274), .A(n275), .ZN(n273) );
  NOR2_X1 U999 ( .A1(n393), .A2(n404), .ZN(n204) );
  NAND2_X1 U1000 ( .A1(n393), .A2(n404), .ZN(n205) );
  XOR2_X1 U1001 ( .A(n262), .B(n73), .Z(product[11]) );
  NAND2_X1 U1002 ( .A1(n971), .A2(n261), .ZN(n73) );
  AOI21_X1 U1003 ( .B1(n267), .B2(n966), .A(n264), .ZN(n262) );
  INV_X1 U1004 ( .A(n157), .ZN(n308) );
  XOR2_X1 U1005 ( .A(n254), .B(n72), .Z(product[12]) );
  XOR2_X1 U1006 ( .A(n170), .B(n61), .Z(product[23]) );
  AOI21_X1 U1007 ( .B1(n1002), .B2(n251), .A(n1001), .ZN(n242) );
  OAI21_X1 U1008 ( .B1(n196), .B2(n162), .A(n163), .ZN(n161) );
  AOI21_X1 U1009 ( .B1(n164), .B2(n189), .A(n165), .ZN(n163) );
  XNOR2_X1 U1010 ( .A(n267), .B(n74), .ZN(product[10]) );
  NAND2_X1 U1011 ( .A1(n966), .A2(n266), .ZN(n74) );
  INV_X1 U1012 ( .A(n99), .ZN(n97) );
  INV_X1 U1013 ( .A(n136), .ZN(n134) );
  AOI21_X1 U1014 ( .B1(n123), .B2(n975), .A(n114), .ZN(n110) );
  INV_X1 U1015 ( .A(n125), .ZN(n123) );
  NAND2_X1 U1016 ( .A1(n417), .A2(n430), .ZN(n219) );
  XNOR2_X1 U1017 ( .A(n247), .B(n71), .ZN(product[13]) );
  OAI21_X1 U1018 ( .B1(n254), .B2(n248), .A(n249), .ZN(n247) );
  INV_X1 U1019 ( .A(n191), .ZN(n189) );
  NAND2_X1 U1020 ( .A1(n445), .A2(n458), .ZN(n233) );
  INV_X1 U1021 ( .A(n182), .ZN(n180) );
  INV_X1 U1022 ( .A(n266), .ZN(n264) );
  NAND2_X1 U1023 ( .A1(n135), .A2(n967), .ZN(n124) );
  NAND2_X1 U1024 ( .A1(n459), .A2(n470), .ZN(n239) );
  NAND2_X1 U1025 ( .A1(n975), .A2(n968), .ZN(n100) );
  INV_X1 U1026 ( .A(n167), .ZN(n166) );
  NAND2_X1 U1027 ( .A1(n98), .A2(n969), .ZN(n87) );
  INV_X1 U1028 ( .A(n135), .ZN(n133) );
  INV_X1 U1029 ( .A(n144), .ZN(n143) );
  AOI21_X1 U1030 ( .B1(n114), .B2(n968), .A(n103), .ZN(n101) );
  INV_X1 U1031 ( .A(n105), .ZN(n103) );
  INV_X1 U1032 ( .A(n288), .ZN(n286) );
  NOR2_X1 U1033 ( .A1(n383), .A2(n392), .ZN(n199) );
  NAND2_X1 U1034 ( .A1(n968), .A2(n105), .ZN(n55) );
  NAND2_X1 U1035 ( .A1(n972), .A2(n288), .ZN(n79) );
  NAND2_X1 U1036 ( .A1(n976), .A2(n280), .ZN(n77) );
  NAND2_X1 U1037 ( .A1(n373), .A2(n382), .ZN(n191) );
  AOI21_X1 U1038 ( .B1(n281), .B2(n976), .A(n278), .ZN(n276) );
  INV_X1 U1039 ( .A(n280), .ZN(n278) );
  XOR2_X1 U1040 ( .A(n117), .B(n56), .Z(product[28]) );
  NAND2_X1 U1041 ( .A1(n975), .A2(n116), .ZN(n56) );
  AOI21_X1 U1042 ( .B1(n136), .B2(n967), .A(n127), .ZN(n125) );
  INV_X1 U1043 ( .A(n129), .ZN(n127) );
  NAND2_X1 U1044 ( .A1(n967), .A2(n129), .ZN(n57) );
  OAI21_X1 U1045 ( .B1(n282), .B2(n284), .A(n283), .ZN(n281) );
  XOR2_X1 U1046 ( .A(n139), .B(n58), .Z(product[26]) );
  NAND2_X1 U1047 ( .A1(n306), .A2(n138), .ZN(n58) );
  INV_X1 U1048 ( .A(n137), .ZN(n306) );
  XOR2_X1 U1049 ( .A(n93), .B(n54), .Z(product[30]) );
  NAND2_X1 U1050 ( .A1(n969), .A2(n92), .ZN(n54) );
  NOR2_X1 U1051 ( .A1(n144), .A2(n137), .ZN(n135) );
  NAND2_X1 U1052 ( .A1(n493), .A2(n502), .ZN(n261) );
  AOI21_X1 U1053 ( .B1(n99), .B2(n969), .A(n90), .ZN(n88) );
  INV_X1 U1054 ( .A(n92), .ZN(n90) );
  NAND2_X1 U1055 ( .A1(n345), .A2(n350), .ZN(n145) );
  INV_X1 U1056 ( .A(n116), .ZN(n114) );
  NAND2_X1 U1057 ( .A1(n326), .A2(n283), .ZN(n78) );
  INV_X1 U1058 ( .A(n282), .ZN(n326) );
  NAND2_X1 U1059 ( .A1(n328), .A2(n291), .ZN(n80) );
  XOR2_X1 U1060 ( .A(n82), .B(n301), .Z(product[2]) );
  NAND2_X1 U1061 ( .A1(n330), .A2(n299), .ZN(n82) );
  INV_X1 U1062 ( .A(n298), .ZN(n330) );
  NAND2_X1 U1063 ( .A1(n574), .A2(n332), .ZN(n92) );
  NAND2_X1 U1064 ( .A1(n535), .A2(n538), .ZN(n288) );
  INV_X1 U1065 ( .A(n332), .ZN(n333) );
  NOR2_X1 U1066 ( .A1(n700), .A2(n685), .ZN(n298) );
  XNOR2_X1 U1067 ( .A(n643), .B(n601), .ZN(n443) );
  OR2_X1 U1068 ( .A1(n643), .A2(n601), .ZN(n442) );
  NAND2_X1 U1069 ( .A1(n700), .A2(n685), .ZN(n299) );
  NAND2_X1 U1070 ( .A1(n337), .A2(n340), .ZN(n129) );
  NAND2_X1 U1071 ( .A1(n525), .A2(n530), .ZN(n280) );
  NAND2_X1 U1072 ( .A1(n336), .A2(n335), .ZN(n116) );
  NAND2_X1 U1073 ( .A1(n334), .A2(n333), .ZN(n105) );
  NAND2_X1 U1074 ( .A1(n531), .A2(n534), .ZN(n283) );
  NAND2_X1 U1075 ( .A1(n341), .A2(n344), .ZN(n138) );
  OAI22_X1 U1076 ( .A1(n5), .A2(n835), .B1(n834), .B2(n877), .ZN(n700) );
  OAI22_X1 U1077 ( .A1(n18), .A2(n788), .B1(n16), .B2(n787), .ZN(n402) );
  OAI22_X1 U1078 ( .A1(n24), .A2(n771), .B1(n22), .B2(n770), .ZN(n380) );
  OAI22_X1 U1079 ( .A1(n42), .A2(n720), .B1(n40), .B2(n719), .ZN(n338) );
  OAI22_X1 U1080 ( .A1(n42), .A2(n731), .B1(n39), .B2(n730), .ZN(n601) );
  OAI22_X1 U1081 ( .A1(n24), .A2(n776), .B1(n22), .B2(n775), .ZN(n643) );
  OAI22_X1 U1082 ( .A1(n30), .A2(n754), .B1(n27), .B2(n753), .ZN(n362) );
  OAI22_X1 U1083 ( .A1(n48), .A2(n704), .B1(n46), .B2(n703), .ZN(n575) );
  INV_X1 U1084 ( .A(n545), .ZN(n590) );
  AOI21_X1 U1085 ( .B1(n42), .B2(n40), .A(n719), .ZN(n545) );
  OAI22_X1 U1086 ( .A1(n48), .A2(n706), .B1(n46), .B2(n705), .ZN(n577) );
  OAI22_X1 U1087 ( .A1(n48), .A2(n705), .B1(n46), .B2(n704), .ZN(n576) );
  INV_X1 U1088 ( .A(n338), .ZN(n339) );
  OAI22_X1 U1089 ( .A1(n17), .A2(n801), .B1(n15), .B2(n800), .ZN(n667) );
  OAI22_X1 U1090 ( .A1(n48), .A2(n878), .B1(n718), .B2(n46), .ZN(n566) );
  OAI22_X1 U1091 ( .A1(n47), .A2(n717), .B1(n45), .B2(n716), .ZN(n588) );
  OR2_X1 U1092 ( .A1(n1013), .A2(n878), .ZN(n718) );
  OAI22_X1 U1093 ( .A1(n11), .A2(n813), .B1(n9), .B2(n812), .ZN(n678) );
  OAI22_X1 U1094 ( .A1(n17), .A2(n798), .B1(n15), .B2(n797), .ZN(n664) );
  OAI22_X1 U1095 ( .A1(n23), .A2(n783), .B1(n21), .B2(n782), .ZN(n650) );
  OAI22_X1 U1096 ( .A1(n11), .A2(n815), .B1(n9), .B2(n814), .ZN(n680) );
  OAI22_X1 U1097 ( .A1(n5), .A2(n830), .B1(n829), .B2(n877), .ZN(n695) );
  OAI22_X1 U1098 ( .A1(n17), .A2(n800), .B1(n15), .B2(n799), .ZN(n666) );
  OAI22_X1 U1099 ( .A1(n35), .A2(n747), .B1(n33), .B2(n746), .ZN(n616) );
  OAI22_X1 U1100 ( .A1(n24), .A2(n777), .B1(n22), .B2(n776), .ZN(n644) );
  OAI22_X1 U1101 ( .A1(n41), .A2(n732), .B1(n39), .B2(n731), .ZN(n602) );
  OAI22_X1 U1102 ( .A1(n24), .A2(n882), .B1(n786), .B2(n22), .ZN(n570) );
  OAI22_X1 U1103 ( .A1(n23), .A2(n785), .B1(n21), .B2(n784), .ZN(n652) );
  OR2_X1 U1104 ( .A1(n1013), .A2(n882), .ZN(n786) );
  OAI22_X1 U1105 ( .A1(n12), .A2(n809), .B1(n10), .B2(n808), .ZN(n674) );
  OAI22_X1 U1106 ( .A1(n6), .A2(n824), .B1(n823), .B2(n4), .ZN(n689) );
  OAI22_X1 U1107 ( .A1(n23), .A2(n779), .B1(n21), .B2(n778), .ZN(n646) );
  OAI22_X1 U1108 ( .A1(n5), .A2(n832), .B1(n831), .B2(n877), .ZN(n697) );
  OAI22_X1 U1109 ( .A1(n11), .A2(n817), .B1(n9), .B2(n816), .ZN(n682) );
  AOI21_X1 U1110 ( .B1(n24), .B2(n22), .A(n770), .ZN(n554) );
  AOI21_X1 U1111 ( .B1(n30), .B2(n27), .A(n753), .ZN(n551) );
  INV_X1 U1112 ( .A(n542), .ZN(n574) );
  AOI21_X1 U1113 ( .B1(n48), .B2(n46), .A(n702), .ZN(n542) );
  AOI21_X1 U1114 ( .B1(n6), .B2(n4), .A(n821), .ZN(n563) );
  OAI22_X1 U1115 ( .A1(n11), .A2(n818), .B1(n9), .B2(n817), .ZN(n683) );
  OAI22_X1 U1116 ( .A1(n5), .A2(n833), .B1(n832), .B2(n4), .ZN(n698) );
  AND2_X1 U1117 ( .A1(n1014), .A2(n558), .ZN(n669) );
  NAND2_X1 U1118 ( .A1(n701), .A2(n573), .ZN(n301) );
  OAI22_X1 U1119 ( .A1(n47), .A2(n712), .B1(n45), .B2(n711), .ZN(n583) );
  INV_X1 U1120 ( .A(n557), .ZN(n654) );
  AOI21_X1 U1121 ( .B1(n18), .B2(n16), .A(n787), .ZN(n557) );
  OAI22_X1 U1122 ( .A1(n48), .A2(n707), .B1(n46), .B2(n706), .ZN(n578) );
  OAI22_X1 U1123 ( .A1(n42), .A2(n722), .B1(n40), .B2(n721), .ZN(n592) );
  OAI22_X1 U1124 ( .A1(n30), .A2(n759), .B1(n27), .B2(n758), .ZN(n627) );
  OAI22_X1 U1125 ( .A1(n35), .A2(n744), .B1(n33), .B2(n743), .ZN(n613) );
  OAI22_X1 U1126 ( .A1(n30), .A2(n760), .B1(n759), .B2(n27), .ZN(n628) );
  OAI22_X1 U1127 ( .A1(n24), .A2(n775), .B1(n22), .B2(n774), .ZN(n642) );
  OAI22_X1 U1128 ( .A1(n41), .A2(n730), .B1(n39), .B2(n729), .ZN(n600) );
  OAI22_X1 U1129 ( .A1(n47), .A2(n711), .B1(n45), .B2(n710), .ZN(n582) );
  OAI22_X1 U1130 ( .A1(n30), .A2(n756), .B1(n27), .B2(n755), .ZN(n624) );
  OAI22_X1 U1131 ( .A1(n42), .A2(n726), .B1(n40), .B2(n725), .ZN(n596) );
  OAI22_X1 U1132 ( .A1(n36), .A2(n740), .B1(n34), .B2(n739), .ZN(n609) );
  OAI22_X1 U1133 ( .A1(n42), .A2(n725), .B1(n40), .B2(n724), .ZN(n595) );
  OAI22_X1 U1134 ( .A1(n24), .A2(n774), .B1(n22), .B2(n773), .ZN(n641) );
  OAI22_X1 U1135 ( .A1(n18), .A2(n789), .B1(n16), .B2(n788), .ZN(n655) );
  OAI22_X1 U1136 ( .A1(n42), .A2(n729), .B1(n39), .B2(n728), .ZN(n599) );
  OAI22_X1 U1137 ( .A1(n23), .A2(n780), .B1(n21), .B2(n779), .ZN(n647) );
  OAI22_X1 U1138 ( .A1(n35), .A2(n750), .B1(n33), .B2(n749), .ZN(n619) );
  OAI22_X1 U1139 ( .A1(n12), .A2(n810), .B1(n10), .B2(n809), .ZN(n675) );
  OAI22_X1 U1140 ( .A1(n18), .A2(n791), .B1(n16), .B2(n790), .ZN(n657) );
  OAI22_X1 U1141 ( .A1(n12), .A2(n806), .B1(n10), .B2(n805), .ZN(n671) );
  OAI22_X1 U1142 ( .A1(n35), .A2(n746), .B1(n33), .B2(n745), .ZN(n615) );
  OAI22_X1 U1143 ( .A1(n48), .A2(n708), .B1(n46), .B2(n707), .ZN(n579) );
  OAI22_X1 U1144 ( .A1(n42), .A2(n723), .B1(n40), .B2(n722), .ZN(n593) );
  INV_X1 U1145 ( .A(n551), .ZN(n622) );
  OAI22_X1 U1146 ( .A1(n18), .A2(n794), .B1(n16), .B2(n793), .ZN(n660) );
  OAI22_X1 U1147 ( .A1(n35), .A2(n749), .B1(n33), .B2(n748), .ZN(n618) );
  OAI22_X1 U1148 ( .A1(n36), .A2(n742), .B1(n34), .B2(n741), .ZN(n611) );
  OAI22_X1 U1149 ( .A1(n24), .A2(n772), .B1(n22), .B2(n771), .ZN(n639) );
  OAI22_X1 U1150 ( .A1(n42), .A2(n727), .B1(n39), .B2(n726), .ZN(n597) );
  OAI22_X1 U1151 ( .A1(n6), .A2(n991), .B1(n824), .B2(n4), .ZN(n690) );
  AND2_X1 U1152 ( .A1(n1014), .A2(n546), .ZN(n605) );
  OAI22_X1 U1153 ( .A1(n6), .A2(n828), .B1(n827), .B2(n4), .ZN(n693) );
  OAI22_X1 U1154 ( .A1(n30), .A2(n758), .B1(n27), .B2(n757), .ZN(n626) );
  OAI22_X1 U1155 ( .A1(n24), .A2(n773), .B1(n22), .B2(n772), .ZN(n640) );
  OAI22_X1 U1156 ( .A1(n36), .A2(n743), .B1(n34), .B2(n742), .ZN(n612) );
  OAI22_X1 U1157 ( .A1(n17), .A2(n797), .B1(n15), .B2(n796), .ZN(n663) );
  OAI22_X1 U1158 ( .A1(n11), .A2(n812), .B1(n9), .B2(n811), .ZN(n677) );
  OAI22_X1 U1159 ( .A1(n30), .A2(n755), .B1(n27), .B2(n754), .ZN(n623) );
  OAI22_X1 U1160 ( .A1(n47), .A2(n710), .B1(n45), .B2(n709), .ZN(n581) );
  INV_X1 U1161 ( .A(n554), .ZN(n638) );
  OAI22_X1 U1162 ( .A1(n23), .A2(n778), .B1(n21), .B2(n777), .ZN(n645) );
  OAI22_X1 U1163 ( .A1(n18), .A2(n793), .B1(n16), .B2(n792), .ZN(n659) );
  OAI22_X1 U1164 ( .A1(n42), .A2(n721), .B1(n40), .B2(n720), .ZN(n591) );
  INV_X1 U1165 ( .A(n548), .ZN(n606) );
  AOI21_X1 U1166 ( .B1(n36), .B2(n34), .A(n736), .ZN(n548) );
  OAI22_X1 U1167 ( .A1(n11), .A2(n814), .B1(n9), .B2(n813), .ZN(n679) );
  OAI22_X1 U1168 ( .A1(n23), .A2(n784), .B1(n21), .B2(n783), .ZN(n651) );
  OAI22_X1 U1169 ( .A1(n12), .A2(n807), .B1(n10), .B2(n806), .ZN(n672) );
  OAI22_X1 U1170 ( .A1(n36), .A2(n738), .B1(n34), .B2(n737), .ZN(n607) );
  OAI22_X1 U1171 ( .A1(n6), .A2(n827), .B1(n826), .B2(n4), .ZN(n692) );
  OAI22_X1 U1172 ( .A1(n23), .A2(n782), .B1(n21), .B2(n781), .ZN(n649) );
  AND2_X1 U1173 ( .A1(n1013), .A2(n549), .ZN(n621) );
  OAI22_X1 U1174 ( .A1(n18), .A2(n792), .B1(n16), .B2(n791), .ZN(n658) );
  OAI22_X1 U1175 ( .A1(n6), .A2(n822), .B1(n821), .B2(n4), .ZN(n687) );
  OAI22_X1 U1176 ( .A1(n6), .A2(n823), .B1(n822), .B2(n4), .ZN(n688) );
  AND2_X1 U1177 ( .A1(n1013), .A2(n543), .ZN(n589) );
  OAI22_X1 U1178 ( .A1(n11), .A2(n816), .B1(n9), .B2(n815), .ZN(n681) );
  OAI22_X1 U1179 ( .A1(n5), .A2(n831), .B1(n830), .B2(n4), .ZN(n696) );
  AND2_X1 U1180 ( .A1(n1013), .A2(n555), .ZN(n653) );
  OAI22_X1 U1181 ( .A1(n47), .A2(n715), .B1(n45), .B2(n714), .ZN(n586) );
  OAI22_X1 U1182 ( .A1(n18), .A2(n790), .B1(n16), .B2(n789), .ZN(n656) );
  OAI22_X1 U1183 ( .A1(n35), .A2(n745), .B1(n33), .B2(n744), .ZN(n614) );
  OAI22_X1 U1184 ( .A1(n36), .A2(n741), .B1(n34), .B2(n740), .ZN(n610) );
  INV_X1 U1185 ( .A(n380), .ZN(n381) );
  OAI22_X1 U1186 ( .A1(n12), .A2(n808), .B1(n10), .B2(n807), .ZN(n673) );
  OAI22_X1 U1187 ( .A1(n42), .A2(n733), .B1(n39), .B2(n732), .ZN(n603) );
  OAI22_X1 U1188 ( .A1(n47), .A2(n714), .B1(n45), .B2(n713), .ZN(n585) );
  OAI22_X1 U1189 ( .A1(n30), .A2(n757), .B1(n27), .B2(n756), .ZN(n625) );
  OAI22_X1 U1190 ( .A1(n23), .A2(n781), .B1(n21), .B2(n780), .ZN(n648) );
  OAI22_X1 U1191 ( .A1(n12), .A2(n811), .B1(n10), .B2(n810), .ZN(n676) );
  OAI22_X1 U1192 ( .A1(n47), .A2(n713), .B1(n45), .B2(n712), .ZN(n584) );
  OAI22_X1 U1193 ( .A1(n41), .A2(n728), .B1(n39), .B2(n727), .ZN(n598) );
  INV_X1 U1194 ( .A(n402), .ZN(n403) );
  OAI22_X1 U1195 ( .A1(n17), .A2(n795), .B1(n15), .B2(n794), .ZN(n661) );
  OAI22_X1 U1196 ( .A1(n17), .A2(n796), .B1(n15), .B2(n795), .ZN(n662) );
  AND2_X1 U1197 ( .A1(n1012), .A2(n552), .ZN(n637) );
  OAI22_X1 U1198 ( .A1(n5), .A2(n829), .B1(n828), .B2(n877), .ZN(n694) );
  OAI22_X1 U1199 ( .A1(n17), .A2(n799), .B1(n15), .B2(n798), .ZN(n665) );
  OAI22_X1 U1200 ( .A1(n36), .A2(n739), .B1(n34), .B2(n738), .ZN(n608) );
  OAI22_X1 U1201 ( .A1(n48), .A2(n709), .B1(n46), .B2(n708), .ZN(n580) );
  OAI22_X1 U1202 ( .A1(n42), .A2(n724), .B1(n40), .B2(n723), .ZN(n594) );
  INV_X1 U1203 ( .A(n27), .ZN(n552) );
  OAI22_X1 U1204 ( .A1(n41), .A2(n734), .B1(n39), .B2(n733), .ZN(n604) );
  NAND2_X1 U1205 ( .A1(n539), .A2(n540), .ZN(n291) );
  AND2_X1 U1206 ( .A1(n1012), .A2(n561), .ZN(n685) );
  INV_X1 U1207 ( .A(n9), .ZN(n561) );
  AND2_X1 U1208 ( .A1(n1013), .A2(a[0]), .ZN(product[0]) );
  OR2_X1 U1209 ( .A1(n1013), .A2(n883), .ZN(n803) );
  OR2_X1 U1210 ( .A1(n1013), .A2(n880), .ZN(n752) );
  OR2_X1 U1211 ( .A1(n1013), .A2(n881), .ZN(n769) );
  OAI22_X1 U1212 ( .A1(n47), .A2(n716), .B1(n45), .B2(n715), .ZN(n587) );
  INV_X1 U1213 ( .A(n563), .ZN(n686) );
  INV_X1 U1214 ( .A(n15), .ZN(n558) );
  INV_X1 U1215 ( .A(n21), .ZN(n555) );
  INV_X1 U1216 ( .A(n39), .ZN(n546) );
  INV_X1 U1217 ( .A(n45), .ZN(n543) );
  INV_X1 U1218 ( .A(n33), .ZN(n549) );
  BUF_X1 U1219 ( .A(n876), .Z(n9) );
  BUF_X1 U1220 ( .A(n865), .Z(n30) );
  OAI22_X1 U1221 ( .A1(n5), .A2(n834), .B1(n833), .B2(n4), .ZN(n699) );
  OAI22_X1 U1222 ( .A1(n12), .A2(n884), .B1(n820), .B2(n10), .ZN(n572) );
  OR2_X1 U1223 ( .A1(n1012), .A2(n884), .ZN(n820) );
  INV_X1 U1224 ( .A(n7), .ZN(n884) );
  BUF_X1 U1225 ( .A(n868), .Z(n12) );
  OAI22_X1 U1226 ( .A1(n6), .A2(n885), .B1(n837), .B2(n4), .ZN(n573) );
  OR2_X1 U1227 ( .A1(n1013), .A2(n885), .ZN(n837) );
  INV_X1 U1228 ( .A(n1), .ZN(n885) );
  OAI22_X1 U1229 ( .A1(n5), .A2(n836), .B1(n835), .B2(n4), .ZN(n701) );
  BUF_X1 U1230 ( .A(n868), .Z(n11) );
  XNOR2_X1 U1231 ( .A(n37), .B(n852), .ZN(n733) );
  XNOR2_X1 U1232 ( .A(n37), .B(n851), .ZN(n732) );
  XNOR2_X1 U1233 ( .A(n37), .B(n850), .ZN(n731) );
  XNOR2_X1 U1234 ( .A(n955), .B(n838), .ZN(n719) );
  OAI22_X1 U1235 ( .A1(n17), .A2(n802), .B1(n15), .B2(n801), .ZN(n668) );
  OAI22_X1 U1236 ( .A1(n18), .A2(n883), .B1(n803), .B2(n16), .ZN(n571) );
  XNOR2_X1 U1237 ( .A(n37), .B(n963), .ZN(n723) );
  XNOR2_X1 U1238 ( .A(n37), .B(n848), .ZN(n729) );
  XNOR2_X1 U1239 ( .A(n37), .B(n849), .ZN(n730) );
  XNOR2_X1 U1240 ( .A(n37), .B(n847), .ZN(n728) );
  XNOR2_X1 U1241 ( .A(n37), .B(n996), .ZN(n725) );
  XNOR2_X1 U1242 ( .A(n37), .B(n846), .ZN(n727) );
  XNOR2_X1 U1243 ( .A(n37), .B(n843), .ZN(n724) );
  XNOR2_X1 U1244 ( .A(n37), .B(n999), .ZN(n726) );
  XNOR2_X1 U1245 ( .A(n955), .B(n841), .ZN(n722) );
  XNOR2_X1 U1246 ( .A(n955), .B(n840), .ZN(n721) );
  XNOR2_X1 U1247 ( .A(n955), .B(n992), .ZN(n720) );
  OAI22_X1 U1248 ( .A1(n35), .A2(n751), .B1(n33), .B2(n750), .ZN(n620) );
  OAI22_X1 U1249 ( .A1(n36), .A2(n880), .B1(n752), .B2(n34), .ZN(n568) );
  BUF_X1 U1250 ( .A(n875), .Z(n15) );
  BUF_X1 U1251 ( .A(n874), .Z(n21) );
  BUF_X1 U1252 ( .A(n870), .Z(n45) );
  BUF_X1 U1253 ( .A(n872), .Z(n33) );
  BUF_X1 U1254 ( .A(n877), .Z(n4) );
  BUF_X1 U1255 ( .A(n875), .Z(n16) );
  BUF_X1 U1256 ( .A(n874), .Z(n22) );
  BUF_X1 U1257 ( .A(n870), .Z(n46) );
  BUF_X1 U1258 ( .A(n866), .Z(n24) );
  BUF_X1 U1259 ( .A(n862), .Z(n48) );
  BUF_X1 U1260 ( .A(n872), .Z(n34) );
  XNOR2_X1 U1261 ( .A(n37), .B(n1014), .ZN(n734) );
  BUF_X1 U1262 ( .A(n869), .Z(n5) );
  BUF_X1 U1263 ( .A(n866), .Z(n23) );
  BUF_X1 U1264 ( .A(n862), .Z(n47) );
  BUF_X1 U1265 ( .A(b[13]), .Z(n840) );
  OAI22_X1 U1266 ( .A1(n30), .A2(n881), .B1(n769), .B2(n27), .ZN(n569) );
  INV_X1 U1267 ( .A(n13), .ZN(n883) );
  INV_X1 U1268 ( .A(n25), .ZN(n881) );
  INV_X1 U1269 ( .A(n19), .ZN(n882) );
  INV_X1 U1270 ( .A(n43), .ZN(n878) );
  INV_X1 U1271 ( .A(n31), .ZN(n880) );
  XNOR2_X1 U1272 ( .A(a[6]), .B(a[5]), .ZN(n874) );
  XNOR2_X1 U1273 ( .A(a[10]), .B(a[9]), .ZN(n872) );
  XNOR2_X1 U1274 ( .A(a[14]), .B(a[13]), .ZN(n870) );
  XNOR2_X1 U1275 ( .A(a[12]), .B(a[11]), .ZN(n871) );
  BUF_X2 U1276 ( .A(a[1]), .Z(n1) );
  BUF_X2 U1277 ( .A(a[3]), .Z(n7) );
  BUF_X2 U1278 ( .A(a[7]), .Z(n19) );
  BUF_X2 U1279 ( .A(a[15]), .Z(n43) );
  NAND2_X1 U1280 ( .A1(n858), .A2(n874), .ZN(n866) );
  NAND2_X1 U1281 ( .A1(n855), .A2(n871), .ZN(n863) );
  NAND2_X1 U1282 ( .A1(n854), .A2(n870), .ZN(n862) );
  NAND2_X1 U1283 ( .A1(n856), .A2(n872), .ZN(n864) );
  INV_X1 U1284 ( .A(a[0]), .ZN(n877) );
  OAI22_X1 U1285 ( .A1(n36), .A2(n737), .B1(n34), .B2(n736), .ZN(n348) );
  INV_X1 U1286 ( .A(n348), .ZN(n349) );
  XNOR2_X1 U1287 ( .A(a[8]), .B(a[7]), .ZN(n873) );
  NAND2_X1 U1288 ( .A1(n860), .A2(n876), .ZN(n868) );
  XNOR2_X1 U1289 ( .A(a[2]), .B(a[1]), .ZN(n876) );
  INV_X1 U1290 ( .A(n290), .ZN(n328) );
  NOR2_X1 U1291 ( .A1(n539), .A2(n540), .ZN(n290) );
  INV_X1 U1292 ( .A(n296), .ZN(n294) );
  NAND2_X1 U1293 ( .A1(n973), .A2(n296), .ZN(n81) );
  OAI22_X1 U1294 ( .A1(n35), .A2(n748), .B1(n33), .B2(n747), .ZN(n617) );
  NAND2_X1 U1295 ( .A1(n861), .A2(n877), .ZN(n869) );
  XNOR2_X1 U1296 ( .A(n7), .B(n841), .ZN(n807) );
  XNOR2_X1 U1297 ( .A(n7), .B(n840), .ZN(n806) );
  XNOR2_X1 U1298 ( .A(n7), .B(n847), .ZN(n813) );
  XNOR2_X1 U1299 ( .A(n7), .B(n996), .ZN(n810) );
  XNOR2_X1 U1300 ( .A(n7), .B(n962), .ZN(n808) );
  XNOR2_X1 U1301 ( .A(n7), .B(n846), .ZN(n812) );
  XNOR2_X1 U1302 ( .A(n7), .B(n998), .ZN(n811) );
  XNOR2_X1 U1303 ( .A(n7), .B(n843), .ZN(n809) );
  XNOR2_X1 U1304 ( .A(n7), .B(n848), .ZN(n814) );
  XNOR2_X1 U1305 ( .A(n7), .B(n851), .ZN(n817) );
  XNOR2_X1 U1306 ( .A(n7), .B(n839), .ZN(n805) );
  XNOR2_X1 U1307 ( .A(n7), .B(n1012), .ZN(n819) );
  XNOR2_X1 U1308 ( .A(n7), .B(n850), .ZN(n816) );
  XNOR2_X1 U1309 ( .A(n7), .B(n838), .ZN(n804) );
  XNOR2_X1 U1310 ( .A(n7), .B(n849), .ZN(n815) );
  XNOR2_X1 U1311 ( .A(n7), .B(n852), .ZN(n818) );
  NAND2_X1 U1312 ( .A1(n977), .A2(n272), .ZN(n75) );
  XNOR2_X1 U1313 ( .A(n25), .B(n1012), .ZN(n768) );
  XNOR2_X1 U1314 ( .A(n25), .B(n847), .ZN(n762) );
  XNOR2_X1 U1315 ( .A(n25), .B(n841), .ZN(n756) );
  XNOR2_X1 U1316 ( .A(n25), .B(n997), .ZN(n760) );
  XNOR2_X1 U1317 ( .A(n25), .B(n846), .ZN(n761) );
  XNOR2_X1 U1318 ( .A(n25), .B(n838), .ZN(n753) );
  XNOR2_X1 U1319 ( .A(n25), .B(n852), .ZN(n767) );
  XNOR2_X1 U1320 ( .A(n25), .B(n994), .ZN(n759) );
  XNOR2_X1 U1321 ( .A(n25), .B(n849), .ZN(n764) );
  XNOR2_X1 U1322 ( .A(n25), .B(n848), .ZN(n763) );
  XNOR2_X1 U1323 ( .A(n25), .B(n840), .ZN(n755) );
  XNOR2_X1 U1324 ( .A(n25), .B(n992), .ZN(n754) );
  XNOR2_X1 U1325 ( .A(n25), .B(n843), .ZN(n758) );
  XNOR2_X1 U1326 ( .A(n25), .B(n851), .ZN(n766) );
  XNOR2_X1 U1327 ( .A(n25), .B(n963), .ZN(n757) );
  OAI21_X1 U1328 ( .B1(n125), .B2(n100), .A(n101), .ZN(n99) );
  NAND2_X1 U1329 ( .A1(n511), .A2(n518), .ZN(n272) );
  INV_X1 U1330 ( .A(n37), .ZN(n879) );
  OR2_X1 U1331 ( .A1(n1014), .A2(n879), .ZN(n735) );
  OAI22_X1 U1332 ( .A1(n41), .A2(n879), .B1(n735), .B2(n40), .ZN(n567) );
  NAND2_X1 U1333 ( .A1(n431), .A2(n444), .ZN(n228) );
  INV_X1 U1334 ( .A(n238), .ZN(n318) );
  NOR2_X1 U1335 ( .A1(n459), .A2(n470), .ZN(n238) );
  NOR2_X1 U1336 ( .A1(n168), .A2(n157), .ZN(n155) );
  INV_X1 U1337 ( .A(n168), .ZN(n167) );
  INV_X1 U1338 ( .A(n560), .ZN(n670) );
  AOI21_X1 U1339 ( .B1(n12), .B2(n10), .A(n804), .ZN(n560) );
  CLKBUF_X1 U1340 ( .A(n876), .Z(n10) );
  NAND2_X1 U1341 ( .A1(n519), .A2(n524), .ZN(n275) );
  NOR2_X1 U1342 ( .A1(n519), .A2(n524), .ZN(n274) );
  XNOR2_X1 U1343 ( .A(n19), .B(n1014), .ZN(n785) );
  XNOR2_X1 U1344 ( .A(n19), .B(n997), .ZN(n777) );
  XNOR2_X1 U1345 ( .A(n19), .B(n994), .ZN(n776) );
  XNOR2_X1 U1346 ( .A(n19), .B(n848), .ZN(n780) );
  XNOR2_X1 U1347 ( .A(n19), .B(n851), .ZN(n783) );
  XNOR2_X1 U1348 ( .A(n19), .B(n852), .ZN(n784) );
  XNOR2_X1 U1349 ( .A(n19), .B(n843), .ZN(n775) );
  XNOR2_X1 U1350 ( .A(n19), .B(n847), .ZN(n779) );
  XNOR2_X1 U1351 ( .A(n19), .B(n846), .ZN(n778) );
  XNOR2_X1 U1352 ( .A(n19), .B(n961), .ZN(n774) );
  XNOR2_X1 U1353 ( .A(n19), .B(n850), .ZN(n782) );
  XNOR2_X1 U1354 ( .A(n19), .B(n849), .ZN(n781) );
  XNOR2_X1 U1355 ( .A(n19), .B(n992), .ZN(n771) );
  XNOR2_X1 U1356 ( .A(n19), .B(n841), .ZN(n773) );
  XNOR2_X1 U1357 ( .A(n19), .B(n840), .ZN(n772) );
  XNOR2_X1 U1358 ( .A(n19), .B(n953), .ZN(n770) );
  AOI21_X1 U1359 ( .B1(n973), .B2(n297), .A(n294), .ZN(n292) );
  XNOR2_X1 U1360 ( .A(n81), .B(n297), .ZN(product[3]) );
  OAI21_X1 U1361 ( .B1(n298), .B2(n301), .A(n299), .ZN(n297) );
  NOR2_X1 U1362 ( .A1(n190), .A2(n153), .ZN(n151) );
  NAND2_X1 U1363 ( .A1(n365), .A2(n372), .ZN(n182) );
  NAND2_X1 U1364 ( .A1(n503), .A2(n510), .ZN(n266) );
  OAI22_X1 U1365 ( .A1(n29), .A2(n763), .B1(n27), .B2(n762), .ZN(n631) );
  OAI22_X1 U1366 ( .A1(n29), .A2(n761), .B1(n27), .B2(n760), .ZN(n629) );
  OAI22_X1 U1367 ( .A1(n29), .A2(n765), .B1(n27), .B2(n764), .ZN(n633) );
  OAI22_X1 U1368 ( .A1(n29), .A2(n764), .B1(n27), .B2(n763), .ZN(n632) );
  OAI22_X1 U1369 ( .A1(n29), .A2(n767), .B1(n27), .B2(n766), .ZN(n635) );
  OAI22_X1 U1370 ( .A1(n29), .A2(n768), .B1(n27), .B2(n767), .ZN(n636) );
  OAI22_X1 U1371 ( .A1(n766), .A2(n29), .B1(n27), .B2(n765), .ZN(n634) );
  XNOR2_X1 U1372 ( .A(n31), .B(n848), .ZN(n746) );
  XNOR2_X1 U1373 ( .A(n31), .B(n843), .ZN(n741) );
  XNOR2_X1 U1374 ( .A(n31), .B(n847), .ZN(n745) );
  XNOR2_X1 U1375 ( .A(n31), .B(n846), .ZN(n744) );
  XNOR2_X1 U1376 ( .A(n31), .B(n840), .ZN(n738) );
  XNOR2_X1 U1377 ( .A(n31), .B(n851), .ZN(n749) );
  XNOR2_X1 U1378 ( .A(n31), .B(n1013), .ZN(n751) );
  XNOR2_X1 U1379 ( .A(n31), .B(n962), .ZN(n740) );
  XNOR2_X1 U1380 ( .A(n31), .B(n850), .ZN(n748) );
  XNOR2_X1 U1381 ( .A(n31), .B(n852), .ZN(n750) );
  XNOR2_X1 U1382 ( .A(n31), .B(n841), .ZN(n739) );
  XNOR2_X1 U1383 ( .A(n31), .B(n849), .ZN(n747) );
  XNOR2_X1 U1384 ( .A(n31), .B(n998), .ZN(n743) );
  XNOR2_X1 U1385 ( .A(n31), .B(n996), .ZN(n742) );
  XNOR2_X1 U1386 ( .A(n31), .B(n992), .ZN(n737) );
  XNOR2_X1 U1387 ( .A(n31), .B(n953), .ZN(n736) );
  NAND2_X1 U1388 ( .A1(n1002), .A2(n246), .ZN(n71) );
  OAI21_X1 U1389 ( .B1(n199), .B2(n205), .A(n200), .ZN(n198) );
  NAND2_X1 U1390 ( .A1(n383), .A2(n392), .ZN(n200) );
  NAND2_X1 U1391 ( .A1(n209), .A2(n225), .ZN(n207) );
  NOR2_X1 U1392 ( .A1(n445), .A2(n458), .ZN(n232) );
  XNOR2_X1 U1393 ( .A(n43), .B(n840), .ZN(n704) );
  XNOR2_X1 U1394 ( .A(n43), .B(n841), .ZN(n705) );
  XNOR2_X1 U1395 ( .A(n43), .B(n992), .ZN(n703) );
  XNOR2_X1 U1396 ( .A(n43), .B(n953), .ZN(n702) );
  XNOR2_X1 U1397 ( .A(n43), .B(n962), .ZN(n706) );
  XNOR2_X1 U1398 ( .A(n43), .B(n843), .ZN(n707) );
  XNOR2_X1 U1399 ( .A(n43), .B(n847), .ZN(n711) );
  XNOR2_X1 U1400 ( .A(n43), .B(n995), .ZN(n708) );
  XNOR2_X1 U1401 ( .A(n43), .B(n846), .ZN(n710) );
  XNOR2_X1 U1402 ( .A(n43), .B(n999), .ZN(n709) );
  XNOR2_X1 U1403 ( .A(n43), .B(n851), .ZN(n715) );
  XNOR2_X1 U1404 ( .A(n43), .B(n848), .ZN(n712) );
  XNOR2_X1 U1405 ( .A(n43), .B(n850), .ZN(n714) );
  XNOR2_X1 U1406 ( .A(n43), .B(n849), .ZN(n713) );
  XNOR2_X1 U1407 ( .A(n43), .B(n1014), .ZN(n717) );
  XNOR2_X1 U1408 ( .A(n43), .B(n852), .ZN(n716) );
  INV_X1 U1409 ( .A(n253), .ZN(n251) );
  NAND2_X1 U1410 ( .A1(n970), .A2(n253), .ZN(n72) );
  NAND2_X1 U1411 ( .A1(n167), .A2(n169), .ZN(n61) );
  OAI21_X1 U1412 ( .B1(n178), .B2(n166), .A(n169), .ZN(n165) );
  OAI21_X1 U1413 ( .B1(n157), .B2(n169), .A(n158), .ZN(n156) );
  NAND2_X1 U1414 ( .A1(n357), .A2(n364), .ZN(n169) );
  NAND2_X1 U1415 ( .A1(n859), .A2(n875), .ZN(n867) );
  XNOR2_X1 U1416 ( .A(n1), .B(n998), .ZN(n828) );
  XNOR2_X1 U1417 ( .A(n1), .B(n1012), .ZN(n836) );
  XNOR2_X1 U1418 ( .A(n1), .B(n846), .ZN(n829) );
  XNOR2_X1 U1419 ( .A(n1), .B(n852), .ZN(n835) );
  XNOR2_X1 U1420 ( .A(n1), .B(n849), .ZN(n832) );
  XNOR2_X1 U1421 ( .A(n1), .B(n841), .ZN(n824) );
  XNOR2_X1 U1422 ( .A(n1), .B(n848), .ZN(n831) );
  XNOR2_X1 U1423 ( .A(n1), .B(n847), .ZN(n830) );
  XNOR2_X1 U1424 ( .A(n1), .B(n840), .ZN(n823) );
  XNOR2_X1 U1425 ( .A(n1), .B(n838), .ZN(n821) );
  XNOR2_X1 U1426 ( .A(n1), .B(n839), .ZN(n822) );
  XNOR2_X1 U1427 ( .A(n1), .B(n962), .ZN(n825) );
  XNOR2_X1 U1428 ( .A(n1), .B(n995), .ZN(n827) );
  XNOR2_X1 U1429 ( .A(n843), .B(n1), .ZN(n826) );
  XNOR2_X1 U1430 ( .A(n1), .B(n851), .ZN(n834) );
  XNOR2_X1 U1431 ( .A(n1), .B(n850), .ZN(n833) );
  OAI22_X1 U1432 ( .A1(n29), .A2(n762), .B1(n27), .B2(n761), .ZN(n630) );
  NAND2_X1 U1433 ( .A1(n857), .A2(n873), .ZN(n865) );
  OAI21_X1 U1434 ( .B1(n224), .B2(n216), .A(n219), .ZN(n215) );
  NOR2_X1 U1435 ( .A1(n223), .A2(n216), .ZN(n214) );
  INV_X1 U1436 ( .A(n150), .ZN(n148) );
  INV_X1 U1437 ( .A(n255), .ZN(n254) );
  AOI21_X1 U1438 ( .B1(n214), .B2(n234), .A(n215), .ZN(n213) );
  AOI21_X1 U1439 ( .B1(n234), .B2(n317), .A(n231), .ZN(n229) );
  INV_X1 U1440 ( .A(n428), .ZN(n429) );
  OAI22_X1 U1441 ( .A1(n12), .A2(n805), .B1(n10), .B2(n804), .ZN(n428) );
  OAI21_X1 U1442 ( .B1(n145), .B2(n137), .A(n138), .ZN(n136) );
  NAND2_X1 U1443 ( .A1(n483), .A2(n492), .ZN(n253) );
  INV_X1 U1444 ( .A(n235), .ZN(n234) );
  OAI21_X1 U1445 ( .B1(n207), .B2(n235), .A(n208), .ZN(n206) );
  INV_X1 U1446 ( .A(n362), .ZN(n363) );
  OAI21_X1 U1447 ( .B1(n268), .B2(n256), .A(n257), .ZN(n255) );
  AOI21_X1 U1448 ( .B1(n255), .B2(n236), .A(n237), .ZN(n235) );
  NOR2_X1 U1449 ( .A1(n1008), .A2(n87), .ZN(n85) );
  NOR2_X1 U1450 ( .A1(n1008), .A2(n133), .ZN(n131) );
  NOR2_X1 U1451 ( .A1(n1008), .A2(n124), .ZN(n118) );
  NOR2_X1 U1452 ( .A1(n1008), .A2(n144), .ZN(n140) );
  NOR2_X1 U1453 ( .A1(n1008), .A2(n96), .ZN(n94) );
  NOR2_X1 U1454 ( .A1(n1008), .A2(n109), .ZN(n107) );
  XOR2_X1 U1455 ( .A(n146), .B(n59), .Z(product[25]) );
  XOR2_X1 U1456 ( .A(n130), .B(n57), .Z(product[27]) );
  AOI21_X1 U1457 ( .B1(n226), .B2(n209), .A(n210), .ZN(n208) );
  NAND2_X1 U1458 ( .A1(n351), .A2(n356), .ZN(n158) );
  XNOR2_X1 U1459 ( .A(n273), .B(n75), .ZN(product[9]) );
  OAI21_X1 U1460 ( .B1(n993), .B2(n233), .A(n228), .ZN(n226) );
  INV_X1 U1461 ( .A(n993), .ZN(n316) );
  NOR2_X1 U1462 ( .A1(n431), .A2(n444), .ZN(n227) );
  OAI21_X1 U1463 ( .B1(n980), .B2(n219), .A(n212), .ZN(n210) );
  NAND2_X1 U1464 ( .A1(n405), .A2(n416), .ZN(n212) );
  OAI21_X1 U1465 ( .B1(n150), .B2(n87), .A(n88), .ZN(n86) );
  OAI21_X1 U1466 ( .B1(n150), .B2(n124), .A(n125), .ZN(n119) );
  OAI21_X1 U1467 ( .B1(n150), .B2(n144), .A(n145), .ZN(n141) );
  OAI21_X1 U1468 ( .B1(n150), .B2(n96), .A(n97), .ZN(n95) );
  OAI21_X1 U1469 ( .B1(n150), .B2(n133), .A(n134), .ZN(n132) );
  OAI21_X1 U1470 ( .B1(n150), .B2(n109), .A(n110), .ZN(n108) );
  INV_X1 U1471 ( .A(n218), .ZN(n217) );
  OAI22_X1 U1472 ( .A1(n11), .A2(n819), .B1(n9), .B2(n818), .ZN(n684) );
  XOR2_X1 U1473 ( .A(n954), .B(n76), .Z(product[8]) );
  XNOR2_X1 U1474 ( .A(n281), .B(n77), .ZN(product[7]) );
  XNOR2_X1 U1475 ( .A(n13), .B(n999), .ZN(n794) );
  XNOR2_X1 U1476 ( .A(n13), .B(n848), .ZN(n797) );
  XNOR2_X1 U1477 ( .A(n13), .B(n995), .ZN(n793) );
  XNOR2_X1 U1478 ( .A(n13), .B(n841), .ZN(n790) );
  XNOR2_X1 U1479 ( .A(n13), .B(n843), .ZN(n792) );
  XNOR2_X1 U1480 ( .A(n13), .B(n840), .ZN(n789) );
  XNOR2_X1 U1481 ( .A(n13), .B(n849), .ZN(n798) );
  XNOR2_X1 U1482 ( .A(n13), .B(n847), .ZN(n796) );
  XNOR2_X1 U1483 ( .A(n13), .B(n963), .ZN(n791) );
  XNOR2_X1 U1484 ( .A(n13), .B(n846), .ZN(n795) );
  XNOR2_X1 U1485 ( .A(n13), .B(n851), .ZN(n800) );
  XNOR2_X1 U1486 ( .A(n13), .B(n850), .ZN(n799) );
  XNOR2_X1 U1487 ( .A(n13), .B(n839), .ZN(n788) );
  XNOR2_X1 U1488 ( .A(n13), .B(n953), .ZN(n787) );
  XNOR2_X1 U1489 ( .A(n13), .B(n1012), .ZN(n802) );
  XNOR2_X1 U1490 ( .A(n13), .B(n852), .ZN(n801) );
  XOR2_X1 U1491 ( .A(n106), .B(n55), .Z(product[29]) );
  XOR2_X1 U1492 ( .A(a[14]), .B(a[15]), .Z(n854) );
  XOR2_X1 U1493 ( .A(a[10]), .B(a[11]), .Z(n856) );
  NOR2_X1 U1494 ( .A1(n241), .A2(n238), .ZN(n236) );
  OAI21_X1 U1495 ( .B1(n242), .B2(n238), .A(n239), .ZN(n237) );
  XOR2_X1 U1496 ( .A(a[12]), .B(a[13]), .Z(n855) );
  XOR2_X1 U1497 ( .A(n220), .B(n67), .Z(product[17]) );
  AOI21_X1 U1498 ( .B1(n234), .B2(n221), .A(n222), .ZN(n220) );
  AOI21_X1 U1499 ( .B1(n1010), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U1500 ( .B1(n1007), .B2(n94), .A(n95), .ZN(n93) );
  AOI21_X1 U1501 ( .B1(n1010), .B2(n118), .A(n119), .ZN(n117) );
  AOI21_X1 U1502 ( .B1(n1010), .B2(n140), .A(n141), .ZN(n139) );
  AOI21_X1 U1503 ( .B1(n1010), .B2(n131), .A(n132), .ZN(n130) );
  AOI21_X1 U1504 ( .B1(n1007), .B2(n197), .A(n194), .ZN(n192) );
  AOI21_X1 U1505 ( .B1(n51), .B2(n313), .A(n203), .ZN(n201) );
  AOI21_X1 U1506 ( .B1(n51), .B2(n171), .A(n172), .ZN(n170) );
  AOI21_X1 U1507 ( .B1(n1007), .B2(n147), .A(n148), .ZN(n146) );
  AOI21_X1 U1508 ( .B1(n1007), .B2(n184), .A(n185), .ZN(n183) );
  AOI21_X1 U1509 ( .B1(n51), .B2(n107), .A(n108), .ZN(n106) );
  AOI21_X1 U1510 ( .B1(n1007), .B2(n160), .A(n161), .ZN(n159) );
  XNOR2_X1 U1511 ( .A(n1011), .B(n65), .ZN(product[19]) );
  OAI21_X1 U1512 ( .B1(n254), .B2(n241), .A(n1000), .ZN(n240) );
  XOR2_X1 U1513 ( .A(a[8]), .B(a[9]), .Z(n857) );
  XOR2_X1 U1514 ( .A(n78), .B(n284), .Z(product[6]) );
  XNOR2_X1 U1515 ( .A(n79), .B(n289), .ZN(product[5]) );
  XOR2_X1 U1516 ( .A(a[6]), .B(a[7]), .Z(n858) );
  XOR2_X1 U1517 ( .A(n80), .B(n292), .Z(product[4]) );
  OAI21_X1 U1518 ( .B1(n290), .B2(n292), .A(n291), .ZN(n289) );
  NAND2_X1 U1519 ( .A1(n541), .A2(n572), .ZN(n296) );
  XNOR2_X1 U1520 ( .A(a[4]), .B(a[3]), .ZN(n875) );
  XOR2_X1 U1521 ( .A(a[2]), .B(a[3]), .Z(n860) );
  XOR2_X1 U1522 ( .A(a[4]), .B(a[5]), .Z(n859) );
  XOR2_X1 U1523 ( .A(a[0]), .B(a[1]), .Z(n861) );
endmodule


module datapath_DW_mult_tc_12 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n3, n4, n5, n7, n9, n10, n11, n12, n13, n15, n16, n17, n18, n19,
         n21, n22, n23, n24, n25, n28, n29, n31, n33, n34, n35, n36, n37, n39,
         n40, n41, n42, n43, n47, n48, n49, n51, n54, n55, n56, n60, n65, n66,
         n67, n68, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n84, n85, n86, n87, n88, n90, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n103, n105, n106, n107, n108, n109, n110, n114, n116,
         n117, n118, n119, n122, n123, n124, n125, n127, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n143,
         n144, n145, n146, n147, n148, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n180, n182, n183, n184, n185, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n218, n219, n220, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n244, n246, n247, n249, n252, n254, n255, n256, n257, n259,
         n261, n262, n264, n266, n267, n268, n270, n272, n273, n274, n275,
         n276, n278, n280, n281, n282, n283, n284, n286, n288, n289, n290,
         n291, n292, n294, n296, n297, n298, n299, n301, n306, n308, n312,
         n313, n314, n315, n318, n324, n326, n328, n330, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n545,
         n546, n548, n549, n551, n552, n554, n555, n557, n558, n560, n561,
         n563, n564, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1065, n1066,
         n1067, n1068;
  assign product[31] = n84;

  FA_X1 U364 ( .A(n575), .B(n338), .CI(n590), .CO(n334), .S(n335) );
  FA_X1 U365 ( .A(n339), .B(n576), .CI(n342), .CO(n336), .S(n337) );
  FA_X1 U367 ( .A(n346), .B(n577), .CI(n343), .CO(n340), .S(n341) );
  FA_X1 U368 ( .A(n591), .B(n348), .CI(n606), .CO(n342), .S(n343) );
  FA_X1 U369 ( .A(n347), .B(n354), .CI(n352), .CO(n344), .S(n345) );
  FA_X1 U370 ( .A(n578), .B(n592), .CI(n349), .CO(n346), .S(n347) );
  FA_X1 U372 ( .A(n358), .B(n355), .CI(n353), .CO(n350), .S(n351) );
  FA_X1 U373 ( .A(n362), .B(n607), .CI(n360), .CO(n352), .S(n353) );
  FA_X1 U374 ( .A(n593), .B(n579), .CI(n622), .CO(n354), .S(n355) );
  FA_X1 U375 ( .A(n359), .B(n361), .CI(n366), .CO(n356), .S(n357) );
  FA_X1 U376 ( .A(n370), .B(n363), .CI(n368), .CO(n358), .S(n359) );
  FA_X1 U377 ( .A(n580), .B(n594), .CI(n608), .CO(n360), .S(n361) );
  FA_X1 U379 ( .A(n367), .B(n376), .CI(n374), .CO(n364), .S(n365) );
  FA_X1 U380 ( .A(n369), .B(n378), .CI(n371), .CO(n366), .S(n367) );
  FA_X1 U381 ( .A(n595), .B(n380), .CI(n609), .CO(n368), .S(n369) );
  FA_X1 U382 ( .A(n623), .B(n581), .CI(n638), .CO(n370), .S(n371) );
  FA_X1 U383 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  FA_X1 U384 ( .A(n379), .B(n388), .CI(n386), .CO(n374), .S(n375) );
  FA_X1 U385 ( .A(n381), .B(n610), .CI(n390), .CO(n376), .S(n377) );
  FA_X1 U386 ( .A(n624), .B(n596), .CI(n582), .CO(n378), .S(n379) );
  FA_X1 U388 ( .A(n394), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U389 ( .A(n391), .B(n389), .CI(n396), .CO(n384), .S(n385) );
  FA_X1 U390 ( .A(n400), .B(n625), .CI(n398), .CO(n386), .S(n387) );
  FA_X1 U391 ( .A(n597), .B(n639), .CI(n611), .CO(n388), .S(n389) );
  FA_X1 U392 ( .A(n1030), .B(n583), .CI(n654), .CO(n390), .S(n391) );
  FA_X1 U394 ( .A(n410), .B(n399), .CI(n408), .CO(n394), .S(n395) );
  FA_X1 U396 ( .A(n584), .B(n598), .CI(n403), .CO(n398), .S(n399) );
  FA_X1 U397 ( .A(n640), .B(n612), .CI(n626), .CO(n400), .S(n401) );
  FA_X1 U399 ( .A(n418), .B(n409), .CI(n407), .CO(n404), .S(n405) );
  FA_X1 U400 ( .A(n411), .B(n422), .CI(n420), .CO(n406), .S(n407) );
  FA_X1 U401 ( .A(n413), .B(n424), .CI(n415), .CO(n408), .S(n409) );
  FA_X1 U403 ( .A(n599), .B(n655), .CI(n641), .CO(n412), .S(n413) );
  FA_X1 U404 ( .A(n428), .B(n585), .CI(n670), .CO(n414), .S(n415) );
  FA_X1 U405 ( .A(n432), .B(n421), .CI(n419), .CO(n416), .S(n417) );
  FA_X1 U406 ( .A(n423), .B(n436), .CI(n434), .CO(n418), .S(n419) );
  FA_X1 U408 ( .A(n442), .B(n429), .CI(n440), .CO(n422), .S(n423) );
  FA_X1 U409 ( .A(n600), .B(n642), .CI(n628), .CO(n424), .S(n425) );
  FA_X1 U410 ( .A(n656), .B(n586), .CI(n614), .CO(n426), .S(n427) );
  FA_X1 U413 ( .A(n448), .B(n450), .CI(n437), .CO(n432), .S(n433) );
  FA_X1 U415 ( .A(n443), .B(n456), .CI(n454), .CO(n436), .S(n437) );
  FA_X1 U416 ( .A(n671), .B(n657), .CI(n615), .CO(n438), .S(n439) );
  FA_X1 U417 ( .A(n587), .B(n686), .CI(n629), .CO(n440), .S(n441) );
  FA_X1 U420 ( .A(n449), .B(n460), .CI(n447), .CO(n444), .S(n445) );
  FA_X1 U421 ( .A(n462), .B(n455), .CI(n451), .CO(n446), .S(n447) );
  FA_X1 U423 ( .A(n457), .B(n672), .CI(n468), .CO(n450), .S(n451) );
  FA_X1 U424 ( .A(n687), .B(n630), .CI(n658), .CO(n452), .S(n453) );
  FA_X1 U425 ( .A(n616), .B(n644), .CI(n602), .CO(n454), .S(n455) );
  HA_X1 U426 ( .A(n566), .B(n588), .CO(n456), .S(n457) );
  FA_X1 U428 ( .A(n465), .B(n467), .CI(n474), .CO(n460), .S(n461) );
  FA_X1 U429 ( .A(n476), .B(n478), .CI(n469), .CO(n462), .S(n463) );
  FA_X1 U430 ( .A(n645), .B(n659), .CI(n480), .CO(n464), .S(n465) );
  FA_X1 U431 ( .A(n603), .B(n673), .CI(n631), .CO(n466), .S(n467) );
  FA_X1 U432 ( .A(n589), .B(n688), .CI(n617), .CO(n468), .S(n469) );
  FA_X1 U434 ( .A(n479), .B(n477), .CI(n486), .CO(n472), .S(n473) );
  FA_X1 U435 ( .A(n490), .B(n481), .CI(n488), .CO(n474), .S(n475) );
  FA_X1 U436 ( .A(n618), .B(n660), .CI(n632), .CO(n476), .S(n477) );
  FA_X1 U437 ( .A(n646), .B(n689), .CI(n674), .CO(n478), .S(n479) );
  HA_X1 U438 ( .A(n604), .B(n567), .CO(n480), .S(n481) );
  FA_X1 U439 ( .A(n487), .B(n494), .CI(n485), .CO(n482), .S(n483) );
  FA_X1 U440 ( .A(n489), .B(n491), .CI(n496), .CO(n484), .S(n485) );
  FA_X1 U441 ( .A(n974), .B(n661), .CI(n498), .CO(n486), .S(n487) );
  FA_X1 U442 ( .A(n619), .B(n675), .CI(n647), .CO(n488), .S(n489) );
  FA_X1 U443 ( .A(n690), .B(n605), .CI(n633), .CO(n490), .S(n491) );
  FA_X1 U444 ( .A(n504), .B(n497), .CI(n495), .CO(n492), .S(n493) );
  FA_X1 U445 ( .A(n506), .B(n508), .CI(n499), .CO(n494), .S(n495) );
  FA_X1 U446 ( .A(n648), .B(n676), .CI(n501), .CO(n496), .S(n497) );
  FA_X1 U447 ( .A(n691), .B(n662), .CI(n634), .CO(n498), .S(n499) );
  FA_X1 U449 ( .A(n512), .B(n507), .CI(n505), .CO(n502), .S(n503) );
  FA_X1 U450 ( .A(n514), .B(n516), .CI(n509), .CO(n504), .S(n505) );
  FA_X1 U451 ( .A(n635), .B(n677), .CI(n663), .CO(n506), .S(n507) );
  FA_X1 U452 ( .A(n649), .B(n621), .CI(n692), .CO(n508), .S(n509) );
  FA_X1 U453 ( .A(n515), .B(n520), .CI(n513), .CO(n510), .S(n511) );
  FA_X1 U454 ( .A(n517), .B(n693), .CI(n522), .CO(n512), .S(n513) );
  FA_X1 U455 ( .A(n650), .B(n664), .CI(n678), .CO(n514), .S(n515) );
  HA_X1 U456 ( .A(n569), .B(n636), .CO(n516), .S(n517) );
  FA_X1 U457 ( .A(n523), .B(n526), .CI(n521), .CO(n518), .S(n519) );
  FA_X1 U458 ( .A(n651), .B(n679), .CI(n528), .CO(n520), .S(n521) );
  FA_X1 U459 ( .A(n665), .B(n637), .CI(n694), .CO(n522), .S(n523) );
  FA_X1 U460 ( .A(n532), .B(n529), .CI(n527), .CO(n524), .S(n525) );
  FA_X1 U461 ( .A(n666), .B(n695), .CI(n680), .CO(n526), .S(n527) );
  HA_X1 U462 ( .A(n570), .B(n652), .CO(n528), .S(n529) );
  FA_X1 U464 ( .A(n653), .B(n696), .CI(n681), .CO(n532), .S(n533) );
  FA_X1 U465 ( .A(n682), .B(n697), .CI(n537), .CO(n534), .S(n535) );
  HA_X1 U466 ( .A(n668), .B(n571), .CO(n536), .S(n537) );
  FA_X1 U467 ( .A(n698), .B(n669), .CI(n683), .CO(n538), .S(n539) );
  HA_X1 U468 ( .A(n684), .B(n699), .CO(n540), .S(n541) );
  CLKBUF_X1 U822 ( .A(b[13]), .Z(n961) );
  CLKBUF_X1 U823 ( .A(n1022), .Z(n953) );
  XNOR2_X1 U824 ( .A(n461), .B(n954), .ZN(n459) );
  XNOR2_X1 U825 ( .A(n472), .B(n463), .ZN(n954) );
  CLKBUF_X1 U826 ( .A(n10), .Z(n955) );
  BUF_X1 U827 ( .A(n10), .Z(n956) );
  BUF_X1 U828 ( .A(n10), .Z(n957) );
  CLKBUF_X1 U829 ( .A(n427), .Z(n958) );
  BUF_X1 U830 ( .A(n864), .Z(n36) );
  CLKBUF_X3 U831 ( .A(n864), .Z(n35) );
  BUF_X4 U832 ( .A(a[15]), .Z(n43) );
  NOR2_X2 U833 ( .A1(n373), .A2(n382), .ZN(n190) );
  AOI21_X2 U834 ( .B1(n198), .B2(n151), .A(n152), .ZN(n150) );
  CLKBUF_X1 U835 ( .A(n242), .Z(n959) );
  BUF_X1 U836 ( .A(n850), .Z(n1017) );
  CLKBUF_X1 U837 ( .A(n1028), .Z(n960) );
  CLKBUF_X1 U838 ( .A(b[3]), .Z(n850) );
  BUF_X2 U839 ( .A(b[15]), .Z(n1065) );
  CLKBUF_X1 U840 ( .A(b[13]), .Z(n840) );
  BUF_X2 U841 ( .A(n867), .Z(n18) );
  AOI21_X1 U842 ( .B1(n273), .B2(n1011), .A(n270), .ZN(n962) );
  CLKBUF_X1 U843 ( .A(n276), .Z(n963) );
  AOI21_X1 U844 ( .B1(n273), .B2(n1011), .A(n270), .ZN(n268) );
  CLKBUF_X1 U845 ( .A(n225), .Z(n1056) );
  BUF_X2 U846 ( .A(b[2]), .Z(n851) );
  CLKBUF_X1 U847 ( .A(n1022), .Z(n964) );
  CLKBUF_X3 U848 ( .A(n25), .Z(n983) );
  BUF_X1 U849 ( .A(n821), .Z(n965) );
  CLKBUF_X3 U850 ( .A(b[11]), .Z(n842) );
  XOR2_X1 U851 ( .A(n401), .B(n412), .Z(n966) );
  XOR2_X1 U852 ( .A(n414), .B(n966), .Z(n397) );
  NAND2_X1 U853 ( .A1(n414), .A2(n401), .ZN(n967) );
  NAND2_X1 U854 ( .A1(n414), .A2(n412), .ZN(n968) );
  NAND2_X1 U855 ( .A1(n401), .A2(n412), .ZN(n969) );
  NAND3_X1 U856 ( .A1(n967), .A2(n968), .A3(n969), .ZN(n396) );
  XOR2_X1 U857 ( .A(n453), .B(n466), .Z(n970) );
  XOR2_X1 U858 ( .A(n464), .B(n970), .Z(n449) );
  NAND2_X1 U859 ( .A1(n464), .A2(n453), .ZN(n971) );
  NAND2_X1 U860 ( .A1(n464), .A2(n466), .ZN(n972) );
  NAND2_X1 U861 ( .A1(n453), .A2(n466), .ZN(n973) );
  NAND3_X1 U862 ( .A1(n971), .A2(n972), .A3(n973), .ZN(n448) );
  OR2_X1 U863 ( .A1(n483), .A2(n492), .ZN(n976) );
  BUF_X2 U864 ( .A(n25), .Z(n984) );
  BUF_X2 U865 ( .A(a[13]), .Z(n37) );
  BUF_X2 U866 ( .A(n49), .Z(n1068) );
  BUF_X1 U867 ( .A(n863), .Z(n42) );
  INV_X1 U868 ( .A(n976), .ZN(n252) );
  AND2_X1 U869 ( .A1(n568), .A2(n620), .ZN(n974) );
  XOR2_X1 U870 ( .A(n568), .B(n620), .Z(n501) );
  CLKBUF_X2 U871 ( .A(b[7]), .Z(n846) );
  CLKBUF_X1 U872 ( .A(n219), .Z(n975) );
  NAND2_X1 U873 ( .A1(n461), .A2(n472), .ZN(n977) );
  NAND2_X1 U874 ( .A1(n461), .A2(n463), .ZN(n978) );
  NAND2_X1 U875 ( .A1(n472), .A2(n463), .ZN(n979) );
  NAND3_X1 U876 ( .A1(n977), .A2(n978), .A3(n979), .ZN(n458) );
  CLKBUF_X3 U877 ( .A(n871), .Z(n39) );
  OAI21_X1 U878 ( .B1(n227), .B2(n233), .A(n228), .ZN(n980) );
  NOR2_X1 U879 ( .A1(n211), .A2(n218), .ZN(n981) );
  CLKBUF_X1 U880 ( .A(n25), .Z(n982) );
  BUF_X1 U881 ( .A(a[9]), .Z(n25) );
  BUF_X1 U882 ( .A(a[1]), .Z(n1) );
  BUF_X1 U883 ( .A(n865), .Z(n29) );
  BUF_X1 U884 ( .A(n867), .Z(n1060) );
  OAI22_X1 U885 ( .A1(n48), .A2(n703), .B1(n1039), .B2(n702), .ZN(n332) );
  XOR2_X1 U886 ( .A(n536), .B(n667), .Z(n985) );
  XOR2_X1 U887 ( .A(n533), .B(n985), .Z(n531) );
  NAND2_X1 U888 ( .A1(n533), .A2(n536), .ZN(n986) );
  NAND2_X1 U889 ( .A1(n533), .A2(n667), .ZN(n987) );
  NAND2_X1 U890 ( .A1(n536), .A2(n667), .ZN(n988) );
  NAND3_X1 U891 ( .A1(n986), .A2(n987), .A3(n988), .ZN(n530) );
  XOR2_X1 U892 ( .A(n613), .B(n627), .Z(n989) );
  XOR2_X1 U893 ( .A(n426), .B(n989), .Z(n411) );
  NAND2_X1 U894 ( .A1(n426), .A2(n613), .ZN(n990) );
  NAND2_X1 U895 ( .A1(n426), .A2(n627), .ZN(n991) );
  NAND2_X1 U896 ( .A1(n613), .A2(n627), .ZN(n992) );
  NAND3_X1 U897 ( .A1(n990), .A2(n991), .A3(n992), .ZN(n410) );
  NAND2_X1 U898 ( .A1(n31), .A2(n846), .ZN(n995) );
  NAND2_X1 U899 ( .A1(n993), .A2(n994), .ZN(n996) );
  NAND2_X1 U900 ( .A1(n995), .A2(n996), .ZN(n744) );
  INV_X1 U901 ( .A(n31), .ZN(n993) );
  INV_X1 U902 ( .A(n846), .ZN(n994) );
  XOR2_X1 U903 ( .A(n406), .B(n397), .Z(n997) );
  XOR2_X1 U904 ( .A(n395), .B(n997), .Z(n393) );
  NAND2_X1 U905 ( .A1(n395), .A2(n406), .ZN(n998) );
  NAND2_X1 U906 ( .A1(n395), .A2(n397), .ZN(n999) );
  NAND2_X1 U907 ( .A1(n406), .A2(n397), .ZN(n1000) );
  NAND3_X1 U908 ( .A1(n998), .A2(n999), .A3(n1000), .ZN(n392) );
  XOR2_X1 U909 ( .A(n441), .B(n452), .Z(n1001) );
  XOR2_X1 U910 ( .A(n439), .B(n1001), .Z(n435) );
  NAND2_X1 U911 ( .A1(n439), .A2(n441), .ZN(n1002) );
  NAND2_X1 U912 ( .A1(n439), .A2(n452), .ZN(n1003) );
  NAND2_X1 U913 ( .A1(n441), .A2(n452), .ZN(n1004) );
  NAND3_X1 U914 ( .A1(n1002), .A2(n1003), .A3(n1004), .ZN(n434) );
  OR2_X1 U915 ( .A1(n503), .A2(n510), .ZN(n1005) );
  OR2_X1 U916 ( .A1(n334), .A2(n333), .ZN(n1006) );
  OR2_X1 U917 ( .A1(n337), .A2(n340), .ZN(n1007) );
  OR2_X1 U918 ( .A1(n574), .A2(n332), .ZN(n1008) );
  OR2_X1 U919 ( .A1(n471), .A2(n482), .ZN(n1009) );
  OR2_X1 U920 ( .A1(n493), .A2(n502), .ZN(n1010) );
  OR2_X1 U921 ( .A1(n511), .A2(n518), .ZN(n1011) );
  OR2_X1 U922 ( .A1(n541), .A2(n572), .ZN(n1012) );
  OR2_X1 U923 ( .A1(n336), .A2(n335), .ZN(n1013) );
  OR2_X1 U924 ( .A1(n525), .A2(n530), .ZN(n1014) );
  OR2_X1 U925 ( .A1(n535), .A2(n538), .ZN(n1015) );
  OR2_X1 U926 ( .A1(n701), .A2(n573), .ZN(n1016) );
  AND2_X1 U927 ( .A1(n483), .A2(n492), .ZN(n1028) );
  CLKBUF_X3 U928 ( .A(b[1]), .Z(n852) );
  BUF_X2 U929 ( .A(n850), .Z(n1018) );
  CLKBUF_X1 U930 ( .A(n871), .Z(n40) );
  CLKBUF_X2 U931 ( .A(a[1]), .Z(n1023) );
  NOR2_X2 U932 ( .A1(n383), .A2(n392), .ZN(n199) );
  CLKBUF_X1 U933 ( .A(n284), .Z(n1019) );
  CLKBUF_X1 U934 ( .A(n1061), .Z(n1020) );
  NOR2_X2 U935 ( .A1(n459), .A2(n470), .ZN(n238) );
  XNOR2_X1 U936 ( .A(n1020), .B(n1021), .ZN(product[15]) );
  AND2_X1 U937 ( .A1(n230), .A2(n233), .ZN(n1021) );
  NAND2_X1 U938 ( .A1(n877), .A2(n861), .ZN(n1022) );
  BUF_X1 U939 ( .A(b[12]), .Z(n841) );
  XOR2_X1 U940 ( .A(n425), .B(n438), .Z(n1024) );
  XOR2_X1 U941 ( .A(n958), .B(n1024), .Z(n421) );
  NAND2_X1 U942 ( .A1(n427), .A2(n425), .ZN(n1025) );
  NAND2_X1 U943 ( .A1(n427), .A2(n438), .ZN(n1026) );
  NAND2_X1 U944 ( .A1(n425), .A2(n438), .ZN(n1027) );
  NAND3_X1 U945 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n420) );
  CLKBUF_X1 U946 ( .A(n211), .Z(n1029) );
  CLKBUF_X2 U947 ( .A(n872), .Z(n33) );
  INV_X1 U948 ( .A(n403), .ZN(n1030) );
  INV_X1 U949 ( .A(n879), .ZN(n1031) );
  BUF_X2 U950 ( .A(n49), .Z(n1067) );
  BUF_X1 U951 ( .A(b[0]), .Z(n49) );
  BUF_X2 U952 ( .A(n869), .Z(n5) );
  BUF_X1 U953 ( .A(n876), .Z(n10) );
  BUF_X2 U954 ( .A(n868), .Z(n12) );
  CLKBUF_X1 U955 ( .A(n872), .Z(n34) );
  BUF_X2 U956 ( .A(n873), .Z(n28) );
  OR2_X1 U957 ( .A1(n365), .A2(n372), .ZN(n1032) );
  BUF_X1 U958 ( .A(n206), .Z(n51) );
  XNOR2_X1 U959 ( .A(n139), .B(n1033), .ZN(product[26]) );
  AND2_X1 U960 ( .A1(n306), .A2(n138), .ZN(n1033) );
  BUF_X2 U961 ( .A(n206), .Z(n1034) );
  BUF_X1 U962 ( .A(n206), .Z(n1035) );
  XNOR2_X1 U963 ( .A(n146), .B(n1036), .ZN(product[25]) );
  AND2_X1 U964 ( .A1(n143), .A2(n145), .ZN(n1036) );
  XNOR2_X1 U965 ( .A(n201), .B(n1037), .ZN(product[20]) );
  AND2_X1 U966 ( .A1(n312), .A2(n200), .ZN(n1037) );
  CLKBUF_X1 U967 ( .A(n843), .Z(n1038) );
  BUF_X2 U968 ( .A(n862), .Z(n47) );
  CLKBUF_X3 U969 ( .A(n870), .Z(n1039) );
  CLKBUF_X1 U970 ( .A(n273), .Z(n1040) );
  XNOR2_X1 U971 ( .A(n183), .B(n1041), .ZN(product[22]) );
  AND2_X1 U972 ( .A1(n175), .A2(n182), .ZN(n1041) );
  OAI21_X1 U973 ( .B1(n256), .B2(n962), .A(n257), .ZN(n1042) );
  BUF_X1 U974 ( .A(n865), .Z(n1043) );
  BUF_X1 U975 ( .A(n865), .Z(n1044) );
  BUF_X2 U976 ( .A(n866), .Z(n23) );
  XNOR2_X1 U977 ( .A(n130), .B(n1045), .ZN(product[27]) );
  AND2_X1 U978 ( .A1(n1007), .A2(n129), .ZN(n1045) );
  BUF_X2 U979 ( .A(a[7]), .Z(n1046) );
  CLKBUF_X1 U980 ( .A(a[7]), .Z(n19) );
  XNOR2_X1 U981 ( .A(n433), .B(n1047), .ZN(n431) );
  XNOR2_X1 U982 ( .A(n446), .B(n435), .ZN(n1047) );
  CLKBUF_X1 U983 ( .A(n218), .Z(n1048) );
  XNOR2_X1 U984 ( .A(n170), .B(n1049), .ZN(product[23]) );
  AND2_X1 U985 ( .A1(n167), .A2(n169), .ZN(n1049) );
  NOR2_X1 U986 ( .A1(n405), .A2(n416), .ZN(n1050) );
  BUF_X2 U987 ( .A(n866), .Z(n24) );
  NOR2_X1 U988 ( .A1(n405), .A2(n416), .ZN(n211) );
  NAND2_X1 U989 ( .A1(n433), .A2(n446), .ZN(n1051) );
  NAND2_X1 U990 ( .A1(n433), .A2(n435), .ZN(n1052) );
  NAND2_X1 U991 ( .A1(n446), .A2(n435), .ZN(n1053) );
  NAND3_X1 U992 ( .A1(n1051), .A2(n1052), .A3(n1053), .ZN(n430) );
  BUF_X4 U993 ( .A(a[11]), .Z(n31) );
  BUF_X1 U994 ( .A(n867), .Z(n17) );
  BUF_X4 U995 ( .A(a[5]), .Z(n13) );
  XNOR2_X1 U996 ( .A(n473), .B(n1054), .ZN(n471) );
  XNOR2_X1 U997 ( .A(n484), .B(n475), .ZN(n1054) );
  XNOR2_X1 U998 ( .A(n192), .B(n1055), .ZN(product[21]) );
  AND2_X1 U999 ( .A1(n188), .A2(n191), .ZN(n1055) );
  NAND2_X1 U1000 ( .A1(n473), .A2(n484), .ZN(n1057) );
  NAND2_X1 U1001 ( .A1(n473), .A2(n475), .ZN(n1058) );
  NAND2_X1 U1002 ( .A1(n484), .A2(n475), .ZN(n1059) );
  NAND3_X1 U1003 ( .A1(n1057), .A2(n1058), .A3(n1059), .ZN(n470) );
  BUF_X2 U1004 ( .A(b[5]), .Z(n848) );
  BUF_X2 U1005 ( .A(b[4]), .Z(n849) );
  BUF_X2 U1006 ( .A(n863), .Z(n41) );
  BUF_X2 U1007 ( .A(b[10]), .Z(n843) );
  AOI21_X1 U1008 ( .B1(n236), .B2(n1042), .A(n237), .ZN(n1061) );
  BUF_X2 U1009 ( .A(b[6]), .Z(n847) );
  OR2_X1 U1010 ( .A1(n431), .A2(n444), .ZN(n1062) );
  NAND2_X1 U1011 ( .A1(n197), .A2(n151), .ZN(n1063) );
  NOR2_X1 U1012 ( .A1(n345), .A2(n350), .ZN(n144) );
  NOR2_X1 U1013 ( .A1(n341), .A2(n344), .ZN(n137) );
  NOR2_X1 U1014 ( .A1(n531), .A2(n534), .ZN(n282) );
  NOR2_X1 U1015 ( .A1(n539), .A2(n540), .ZN(n290) );
  AND2_X1 U1016 ( .A1(n1016), .A2(n301), .ZN(product[1]) );
  BUF_X1 U1017 ( .A(n875), .Z(n15) );
  BUF_X1 U1018 ( .A(n876), .Z(n9) );
  BUF_X2 U1019 ( .A(a[3]), .Z(n7) );
  XNOR2_X1 U1020 ( .A(n13), .B(n1065), .ZN(n787) );
  INV_X1 U1021 ( .A(n980), .ZN(n224) );
  INV_X1 U1022 ( .A(n1056), .ZN(n223) );
  NOR2_X1 U1023 ( .A1(n195), .A2(n190), .ZN(n184) );
  NOR2_X1 U1024 ( .A1(n195), .A2(n162), .ZN(n160) );
  NOR2_X1 U1025 ( .A1(n195), .A2(n173), .ZN(n171) );
  NOR2_X1 U1026 ( .A1(n1063), .A2(n124), .ZN(n118) );
  NOR2_X1 U1027 ( .A1(n1063), .A2(n109), .ZN(n107) );
  NOR2_X1 U1028 ( .A1(n1063), .A2(n96), .ZN(n94) );
  INV_X1 U1029 ( .A(n98), .ZN(n96) );
  NOR2_X1 U1030 ( .A1(n223), .A2(n1048), .ZN(n214) );
  INV_X1 U1031 ( .A(n177), .ZN(n175) );
  INV_X1 U1032 ( .A(n1063), .ZN(n147) );
  INV_X1 U1033 ( .A(n195), .ZN(n193) );
  INV_X1 U1034 ( .A(n196), .ZN(n194) );
  NAND2_X1 U1035 ( .A1(n313), .A2(n205), .ZN(n65) );
  INV_X1 U1036 ( .A(n204), .ZN(n313) );
  XOR2_X1 U1037 ( .A(n213), .B(n66), .Z(product[18]) );
  NAND2_X1 U1038 ( .A1(n314), .A2(n212), .ZN(n66) );
  INV_X1 U1039 ( .A(n1029), .ZN(n314) );
  XNOR2_X1 U1040 ( .A(n240), .B(n70), .ZN(product[14]) );
  NAND2_X1 U1041 ( .A1(n318), .A2(n239), .ZN(n70) );
  INV_X1 U1042 ( .A(n238), .ZN(n318) );
  XOR2_X1 U1043 ( .A(n220), .B(n67), .Z(product[17]) );
  NAND2_X1 U1044 ( .A1(n315), .A2(n975), .ZN(n67) );
  OAI21_X1 U1045 ( .B1(n227), .B2(n233), .A(n228), .ZN(n226) );
  XOR2_X1 U1046 ( .A(n229), .B(n68), .Z(product[16]) );
  NAND2_X1 U1047 ( .A1(n1062), .A2(n228), .ZN(n68) );
  NOR2_X1 U1048 ( .A1(n177), .A2(n166), .ZN(n164) );
  NOR2_X1 U1049 ( .A1(n124), .A2(n100), .ZN(n98) );
  OAI21_X1 U1050 ( .B1(n196), .B2(n173), .A(n174), .ZN(n172) );
  AOI21_X1 U1051 ( .B1(n189), .B2(n175), .A(n176), .ZN(n174) );
  INV_X1 U1052 ( .A(n178), .ZN(n176) );
  INV_X1 U1053 ( .A(n197), .ZN(n195) );
  INV_X1 U1054 ( .A(n198), .ZN(n196) );
  INV_X1 U1055 ( .A(n962), .ZN(n267) );
  NAND2_X1 U1056 ( .A1(n164), .A2(n188), .ZN(n162) );
  NAND2_X1 U1057 ( .A1(n188), .A2(n175), .ZN(n173) );
  OAI21_X1 U1058 ( .B1(n196), .B2(n190), .A(n191), .ZN(n185) );
  OAI21_X1 U1059 ( .B1(n224), .B2(n1048), .A(n975), .ZN(n215) );
  INV_X1 U1060 ( .A(n1032), .ZN(n177) );
  INV_X1 U1061 ( .A(n180), .ZN(n178) );
  NOR2_X1 U1062 ( .A1(n1063), .A2(n144), .ZN(n140) );
  NOR2_X1 U1063 ( .A1(n1063), .A2(n133), .ZN(n131) );
  INV_X1 U1064 ( .A(n124), .ZN(n122) );
  NAND2_X1 U1065 ( .A1(n122), .A2(n1013), .ZN(n109) );
  NAND2_X1 U1066 ( .A1(n1009), .A2(n976), .ZN(n241) );
  INV_X1 U1067 ( .A(n150), .ZN(n148) );
  INV_X1 U1068 ( .A(n205), .ZN(n203) );
  INV_X1 U1069 ( .A(n233), .ZN(n231) );
  INV_X1 U1070 ( .A(n960), .ZN(n249) );
  INV_X1 U1071 ( .A(n232), .ZN(n230) );
  NAND2_X1 U1072 ( .A1(n1011), .A2(n272), .ZN(n75) );
  XOR2_X1 U1073 ( .A(n254), .B(n72), .Z(product[12]) );
  NAND2_X1 U1074 ( .A1(n976), .A2(n249), .ZN(n72) );
  XNOR2_X1 U1075 ( .A(n267), .B(n74), .ZN(product[10]) );
  NAND2_X1 U1076 ( .A1(n1005), .A2(n266), .ZN(n74) );
  INV_X1 U1077 ( .A(n272), .ZN(n270) );
  XOR2_X1 U1078 ( .A(n159), .B(n60), .Z(product[24]) );
  NAND2_X1 U1079 ( .A1(n308), .A2(n158), .ZN(n60) );
  NOR2_X1 U1080 ( .A1(n431), .A2(n444), .ZN(n227) );
  INV_X1 U1081 ( .A(n199), .ZN(n312) );
  OAI21_X1 U1082 ( .B1(n199), .B2(n205), .A(n200), .ZN(n198) );
  NAND2_X1 U1083 ( .A1(n1010), .A2(n1005), .ZN(n256) );
  AOI21_X1 U1084 ( .B1(n1010), .B2(n264), .A(n259), .ZN(n257) );
  XOR2_X1 U1085 ( .A(n262), .B(n73), .Z(product[11]) );
  NAND2_X1 U1086 ( .A1(n1010), .A2(n261), .ZN(n73) );
  AOI21_X1 U1087 ( .B1(n267), .B2(n1005), .A(n264), .ZN(n262) );
  NAND2_X1 U1088 ( .A1(n445), .A2(n458), .ZN(n233) );
  NAND2_X1 U1089 ( .A1(n393), .A2(n404), .ZN(n205) );
  INV_X1 U1090 ( .A(n190), .ZN(n188) );
  XNOR2_X1 U1091 ( .A(n247), .B(n71), .ZN(product[13]) );
  OAI21_X1 U1092 ( .B1(n254), .B2(n252), .A(n249), .ZN(n247) );
  NOR2_X1 U1093 ( .A1(n393), .A2(n404), .ZN(n204) );
  NOR2_X1 U1094 ( .A1(n445), .A2(n458), .ZN(n232) );
  AOI21_X1 U1095 ( .B1(n123), .B2(n1013), .A(n114), .ZN(n110) );
  INV_X1 U1096 ( .A(n136), .ZN(n134) );
  NAND2_X1 U1097 ( .A1(n417), .A2(n430), .ZN(n219) );
  INV_X1 U1098 ( .A(n191), .ZN(n189) );
  NAND2_X1 U1099 ( .A1(n98), .A2(n1008), .ZN(n87) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1006), .ZN(n100) );
  NAND2_X1 U1101 ( .A1(n135), .A2(n1007), .ZN(n124) );
  OAI21_X1 U1102 ( .B1(n150), .B2(n96), .A(n97), .ZN(n95) );
  INV_X1 U1103 ( .A(n99), .ZN(n97) );
  NAND2_X1 U1104 ( .A1(n405), .A2(n416), .ZN(n212) );
  OAI21_X1 U1105 ( .B1(n196), .B2(n162), .A(n163), .ZN(n161) );
  AOI21_X1 U1106 ( .B1(n164), .B2(n189), .A(n165), .ZN(n163) );
  OAI21_X1 U1107 ( .B1(n178), .B2(n166), .A(n169), .ZN(n165) );
  NOR2_X1 U1108 ( .A1(n1063), .A2(n87), .ZN(n85) );
  OAI21_X1 U1109 ( .B1(n150), .B2(n87), .A(n88), .ZN(n86) );
  INV_X1 U1110 ( .A(n167), .ZN(n166) );
  INV_X1 U1111 ( .A(n266), .ZN(n264) );
  INV_X1 U1112 ( .A(n125), .ZN(n123) );
  INV_X1 U1113 ( .A(n135), .ZN(n133) );
  INV_X1 U1114 ( .A(n144), .ZN(n143) );
  INV_X1 U1115 ( .A(n261), .ZN(n259) );
  NAND2_X1 U1116 ( .A1(n326), .A2(n283), .ZN(n78) );
  INV_X1 U1117 ( .A(n282), .ZN(n326) );
  NAND2_X1 U1118 ( .A1(n324), .A2(n275), .ZN(n76) );
  INV_X1 U1119 ( .A(n274), .ZN(n324) );
  NAND2_X1 U1120 ( .A1(n1014), .A2(n280), .ZN(n77) );
  INV_X1 U1121 ( .A(n137), .ZN(n306) );
  NAND2_X1 U1122 ( .A1(n1008), .A2(n92), .ZN(n54) );
  INV_X1 U1123 ( .A(n280), .ZN(n278) );
  NAND2_X1 U1124 ( .A1(n1013), .A2(n116), .ZN(n56) );
  NAND2_X1 U1125 ( .A1(n1006), .A2(n105), .ZN(n55) );
  AOI21_X1 U1126 ( .B1(n136), .B2(n1007), .A(n127), .ZN(n125) );
  INV_X1 U1127 ( .A(n129), .ZN(n127) );
  OAI21_X1 U1128 ( .B1(n145), .B2(n137), .A(n138), .ZN(n136) );
  OAI21_X1 U1129 ( .B1(n125), .B2(n100), .A(n101), .ZN(n99) );
  AOI21_X1 U1130 ( .B1(n114), .B2(n1006), .A(n103), .ZN(n101) );
  INV_X1 U1131 ( .A(n105), .ZN(n103) );
  NOR2_X1 U1132 ( .A1(n144), .A2(n137), .ZN(n135) );
  NOR2_X1 U1133 ( .A1(n351), .A2(n356), .ZN(n157) );
  AOI21_X1 U1134 ( .B1(n99), .B2(n1008), .A(n90), .ZN(n88) );
  INV_X1 U1135 ( .A(n92), .ZN(n90) );
  AOI21_X1 U1136 ( .B1(n1015), .B2(n289), .A(n286), .ZN(n284) );
  INV_X1 U1137 ( .A(n288), .ZN(n286) );
  NAND2_X1 U1138 ( .A1(n345), .A2(n350), .ZN(n145) );
  NAND2_X1 U1139 ( .A1(n373), .A2(n382), .ZN(n191) );
  NAND2_X1 U1140 ( .A1(n503), .A2(n510), .ZN(n266) );
  NAND2_X1 U1141 ( .A1(n511), .A2(n518), .ZN(n272) );
  NAND2_X1 U1142 ( .A1(n493), .A2(n502), .ZN(n261) );
  NAND2_X1 U1143 ( .A1(n383), .A2(n392), .ZN(n200) );
  INV_X1 U1144 ( .A(n116), .ZN(n114) );
  XNOR2_X1 U1145 ( .A(n79), .B(n289), .ZN(product[5]) );
  NAND2_X1 U1146 ( .A1(n1015), .A2(n288), .ZN(n79) );
  XOR2_X1 U1147 ( .A(n80), .B(n292), .Z(product[4]) );
  NAND2_X1 U1148 ( .A1(n328), .A2(n291), .ZN(n80) );
  INV_X1 U1149 ( .A(n290), .ZN(n328) );
  NOR2_X1 U1150 ( .A1(n700), .A2(n685), .ZN(n298) );
  XNOR2_X1 U1151 ( .A(n81), .B(n297), .ZN(product[3]) );
  NAND2_X1 U1152 ( .A1(n1012), .A2(n296), .ZN(n81) );
  AOI21_X1 U1153 ( .B1(n1012), .B2(n297), .A(n294), .ZN(n292) );
  NOR2_X1 U1154 ( .A1(n519), .A2(n524), .ZN(n274) );
  OAI21_X1 U1155 ( .B1(n290), .B2(n292), .A(n291), .ZN(n289) );
  NAND2_X1 U1156 ( .A1(n574), .A2(n332), .ZN(n92) );
  OAI21_X1 U1157 ( .B1(n298), .B2(n301), .A(n299), .ZN(n297) );
  XNOR2_X1 U1158 ( .A(n643), .B(n601), .ZN(n443) );
  INV_X1 U1159 ( .A(n332), .ZN(n333) );
  NAND2_X1 U1160 ( .A1(n700), .A2(n685), .ZN(n299) );
  INV_X1 U1161 ( .A(n428), .ZN(n429) );
  OR2_X1 U1162 ( .A1(n643), .A2(n601), .ZN(n442) );
  NAND2_X1 U1163 ( .A1(n535), .A2(n538), .ZN(n288) );
  NAND2_X1 U1164 ( .A1(n337), .A2(n340), .ZN(n129) );
  NAND2_X1 U1165 ( .A1(n341), .A2(n344), .ZN(n138) );
  NAND2_X1 U1166 ( .A1(n336), .A2(n335), .ZN(n116) );
  NAND2_X1 U1167 ( .A1(n334), .A2(n333), .ZN(n105) );
  NAND2_X1 U1168 ( .A1(n525), .A2(n530), .ZN(n280) );
  NAND2_X1 U1169 ( .A1(n531), .A2(n534), .ZN(n283) );
  XOR2_X1 U1170 ( .A(n82), .B(n301), .Z(product[2]) );
  NAND2_X1 U1171 ( .A1(n330), .A2(n299), .ZN(n82) );
  INV_X1 U1172 ( .A(n298), .ZN(n330) );
  OAI22_X1 U1173 ( .A1(n41), .A2(n720), .B1(n39), .B2(n719), .ZN(n338) );
  OAI22_X1 U1174 ( .A1(n5), .A2(n835), .B1(n834), .B2(n3), .ZN(n700) );
  OAI22_X1 U1175 ( .A1(n12), .A2(n805), .B1(n957), .B2(n804), .ZN(n428) );
  OAI22_X1 U1176 ( .A1(n24), .A2(n771), .B1(n22), .B2(n770), .ZN(n380) );
  OAI22_X1 U1177 ( .A1(n11), .A2(n813), .B1(n9), .B2(n812), .ZN(n678) );
  OAI22_X1 U1178 ( .A1(n48), .A2(n704), .B1(n1039), .B2(n703), .ZN(n575) );
  INV_X1 U1179 ( .A(n545), .ZN(n590) );
  AOI21_X1 U1180 ( .B1(n41), .B2(n39), .A(n719), .ZN(n545) );
  OAI22_X1 U1181 ( .A1(n48), .A2(n705), .B1(n1039), .B2(n704), .ZN(n576) );
  INV_X1 U1182 ( .A(n338), .ZN(n339) );
  OAI22_X1 U1183 ( .A1(n11), .A2(n817), .B1(n9), .B2(n816), .ZN(n682) );
  OAI22_X1 U1184 ( .A1(n5), .A2(n832), .B1(n831), .B2(n3), .ZN(n697) );
  OAI22_X1 U1185 ( .A1(n48), .A2(n706), .B1(n1039), .B2(n705), .ZN(n577) );
  OAI22_X1 U1186 ( .A1(n11), .A2(n818), .B1(n9), .B2(n817), .ZN(n683) );
  AND2_X1 U1187 ( .A1(n1067), .A2(n558), .ZN(n669) );
  OAI22_X1 U1188 ( .A1(n5), .A2(n833), .B1(n832), .B2(n3), .ZN(n698) );
  OAI22_X1 U1189 ( .A1(n48), .A2(n878), .B1(n718), .B2(n1039), .ZN(n566) );
  OAI22_X1 U1190 ( .A1(n47), .A2(n717), .B1(n1039), .B2(n716), .ZN(n588) );
  OR2_X1 U1191 ( .A1(n1067), .A2(n878), .ZN(n718) );
  AND2_X1 U1192 ( .A1(n1067), .A2(n555), .ZN(n653) );
  OAI22_X1 U1193 ( .A1(n12), .A2(n816), .B1(n9), .B2(n815), .ZN(n681) );
  OAI22_X1 U1194 ( .A1(n5), .A2(n831), .B1(n830), .B2(n3), .ZN(n696) );
  OAI22_X1 U1195 ( .A1(n12), .A2(n806), .B1(n956), .B2(n805), .ZN(n671) );
  OAI22_X1 U1196 ( .A1(n36), .A2(n746), .B1(n33), .B2(n745), .ZN(n615) );
  OAI22_X1 U1197 ( .A1(n35), .A2(n739), .B1(n34), .B2(n738), .ZN(n608) );
  OAI22_X1 U1198 ( .A1(n41), .A2(n724), .B1(n39), .B2(n723), .ZN(n594) );
  OAI22_X1 U1199 ( .A1(n5), .A2(n822), .B1(n4), .B2(n965), .ZN(n687) );
  OAI22_X1 U1200 ( .A1(n29), .A2(n762), .B1(n28), .B2(n761), .ZN(n630) );
  OAI22_X1 U1201 ( .A1(n47), .A2(n715), .B1(n1039), .B2(n714), .ZN(n586) );
  OAI22_X1 U1202 ( .A1(n35), .A2(n745), .B1(n744), .B2(n33), .ZN(n614) );
  INV_X1 U1203 ( .A(n542), .ZN(n574) );
  AOI21_X1 U1204 ( .B1(n48), .B2(n1039), .A(n702), .ZN(n542) );
  OAI22_X1 U1205 ( .A1(n36), .A2(n880), .B1(n752), .B2(n33), .ZN(n568) );
  OAI22_X1 U1206 ( .A1(n751), .A2(n36), .B1(n33), .B2(n750), .ZN(n620) );
  OR2_X1 U1207 ( .A1(n1068), .A2(n880), .ZN(n752) );
  NAND2_X1 U1208 ( .A1(n701), .A2(n573), .ZN(n301) );
  AND2_X1 U1209 ( .A1(n1067), .A2(n561), .ZN(n685) );
  INV_X1 U1210 ( .A(n9), .ZN(n561) );
  AND2_X1 U1211 ( .A1(n1067), .A2(n564), .ZN(product[0]) );
  INV_X1 U1212 ( .A(n3), .ZN(n564) );
  OAI22_X1 U1213 ( .A1(n41), .A2(n722), .B1(n39), .B2(n721), .ZN(n592) );
  OAI22_X1 U1214 ( .A1(n48), .A2(n707), .B1(n1039), .B2(n706), .ZN(n578) );
  OAI22_X1 U1215 ( .A1(n35), .A2(n744), .B1(n34), .B2(n743), .ZN(n613) );
  OAI22_X1 U1216 ( .A1(n48), .A2(n711), .B1(n1039), .B2(n710), .ZN(n582) );
  OAI22_X1 U1217 ( .A1(n41), .A2(n726), .B1(n39), .B2(n725), .ZN(n596) );
  OAI22_X1 U1218 ( .A1(n35), .A2(n740), .B1(n34), .B2(n739), .ZN(n609) );
  OAI22_X1 U1219 ( .A1(n41), .A2(n725), .B1(n39), .B2(n724), .ZN(n595) );
  OAI22_X1 U1220 ( .A1(n35), .A2(n750), .B1(n33), .B2(n749), .ZN(n619) );
  OAI22_X1 U1221 ( .A1(n12), .A2(n810), .B1(n957), .B2(n809), .ZN(n675) );
  OAI22_X1 U1222 ( .A1(n35), .A2(n741), .B1(n34), .B2(n740), .ZN(n610) );
  INV_X1 U1223 ( .A(n380), .ZN(n381) );
  OAI22_X1 U1224 ( .A1(n953), .A2(n825), .B1(n824), .B2(n4), .ZN(n690) );
  OAI22_X1 U1225 ( .A1(n1044), .A2(n765), .B1(n28), .B2(n764), .ZN(n633) );
  AND2_X1 U1226 ( .A1(n1067), .A2(n546), .ZN(n605) );
  OAI22_X1 U1227 ( .A1(n35), .A2(n742), .B1(n34), .B2(n741), .ZN(n611) );
  OAI22_X1 U1228 ( .A1(n11), .A2(n812), .B1(n9), .B2(n811), .ZN(n677) );
  OAI22_X1 U1229 ( .A1(n29), .A2(n767), .B1(n28), .B2(n766), .ZN(n635) );
  OAI22_X1 U1230 ( .A1(n35), .A2(n749), .B1(n33), .B2(n748), .ZN(n618) );
  OAI22_X1 U1231 ( .A1(n1043), .A2(n764), .B1(n28), .B2(n763), .ZN(n632) );
  OAI22_X1 U1232 ( .A1(n36), .A2(n743), .B1(n33), .B2(n742), .ZN(n612) );
  OAI22_X1 U1233 ( .A1(n41), .A2(n721), .B1(n39), .B2(n720), .ZN(n591) );
  INV_X1 U1234 ( .A(n548), .ZN(n606) );
  AOI21_X1 U1235 ( .B1(n35), .B2(n34), .A(n736), .ZN(n548) );
  OAI22_X1 U1236 ( .A1(n11), .A2(n814), .B1(n9), .B2(n813), .ZN(n679) );
  OAI22_X1 U1237 ( .A1(n48), .A2(n710), .B1(n1039), .B2(n709), .ZN(n581) );
  INV_X1 U1238 ( .A(n554), .ZN(n638) );
  OAI22_X1 U1239 ( .A1(n5), .A2(n828), .B1(n827), .B2(n4), .ZN(n693) );
  OAI22_X1 U1240 ( .A1(n11), .A2(n807), .B1(n957), .B2(n806), .ZN(n672) );
  OAI22_X1 U1241 ( .A1(n5), .A2(n827), .B1(n826), .B2(n4), .ZN(n692) );
  AND2_X1 U1242 ( .A1(n1067), .A2(n549), .ZN(n621) );
  OAI22_X1 U1243 ( .A1(n5), .A2(n830), .B1(n829), .B2(n3), .ZN(n695) );
  OAI22_X1 U1244 ( .A1(n11), .A2(n815), .B1(n9), .B2(n814), .ZN(n680) );
  OAI22_X1 U1245 ( .A1(n1044), .A2(n763), .B1(n28), .B2(n762), .ZN(n631) );
  OAI22_X1 U1246 ( .A1(n11), .A2(n808), .B1(n957), .B2(n807), .ZN(n673) );
  OAI22_X1 U1247 ( .A1(n953), .A2(n824), .B1(n823), .B2(n4), .ZN(n689) );
  OAI22_X1 U1248 ( .A1(n12), .A2(n809), .B1(n955), .B2(n808), .ZN(n674) );
  AOI21_X1 U1249 ( .B1(n12), .B2(n956), .A(n804), .ZN(n560) );
  OAI22_X1 U1250 ( .A1(n41), .A2(n723), .B1(n39), .B2(n722), .ZN(n593) );
  OAI22_X1 U1251 ( .A1(n48), .A2(n708), .B1(n1039), .B2(n707), .ZN(n579) );
  INV_X1 U1252 ( .A(n551), .ZN(n622) );
  OAI22_X1 U1253 ( .A1(n11), .A2(n811), .B1(n956), .B2(n810), .ZN(n676) );
  OAI22_X1 U1254 ( .A1(n35), .A2(n747), .B1(n33), .B2(n746), .ZN(n616) );
  OAI22_X1 U1255 ( .A1(n823), .A2(n1022), .B1(n822), .B2(n4), .ZN(n688) );
  OAI22_X1 U1256 ( .A1(n36), .A2(n748), .B1(n33), .B2(n747), .ZN(n617) );
  AND2_X1 U1257 ( .A1(n1067), .A2(n543), .ZN(n589) );
  OAI22_X1 U1258 ( .A1(n35), .A2(n738), .B1(n34), .B2(n737), .ZN(n607) );
  OAI22_X1 U1259 ( .A1(n47), .A2(n716), .B1(n1039), .B2(n715), .ZN(n587) );
  OAI22_X1 U1260 ( .A1(n761), .A2(n1043), .B1(n28), .B2(n760), .ZN(n629) );
  INV_X1 U1261 ( .A(n563), .ZN(n686) );
  OAI22_X1 U1262 ( .A1(n5), .A2(n826), .B1(n825), .B2(n4), .ZN(n691) );
  OAI22_X1 U1263 ( .A1(n5), .A2(n829), .B1(n828), .B2(n3), .ZN(n694) );
  AND2_X1 U1264 ( .A1(n1067), .A2(n552), .ZN(n637) );
  NAND2_X1 U1265 ( .A1(n539), .A2(n540), .ZN(n291) );
  OAI22_X1 U1266 ( .A1(n42), .A2(n879), .B1(n735), .B2(n40), .ZN(n567) );
  OR2_X1 U1267 ( .A1(n1068), .A2(n879), .ZN(n735) );
  INV_X1 U1268 ( .A(n870), .ZN(n543) );
  OR2_X1 U1269 ( .A1(n1067), .A2(n881), .ZN(n769) );
  INV_X1 U1270 ( .A(n33), .ZN(n549) );
  INV_X1 U1271 ( .A(n28), .ZN(n552) );
  INV_X1 U1272 ( .A(n15), .ZN(n558) );
  INV_X1 U1273 ( .A(n40), .ZN(n546) );
  BUF_X1 U1274 ( .A(n877), .Z(n3) );
  BUF_X1 U1275 ( .A(n877), .Z(n4) );
  OAI22_X1 U1276 ( .A1(n11), .A2(n884), .B1(n820), .B2(n956), .ZN(n572) );
  OR2_X1 U1277 ( .A1(n1067), .A2(n884), .ZN(n820) );
  INV_X1 U1278 ( .A(n7), .ZN(n884) );
  OAI22_X1 U1279 ( .A1(n11), .A2(n819), .B1(n9), .B2(n818), .ZN(n684) );
  OAI22_X1 U1280 ( .A1(n1043), .A2(n768), .B1(n28), .B2(n767), .ZN(n636) );
  OAI22_X1 U1281 ( .A1(n18), .A2(n788), .B1(n16), .B2(n787), .ZN(n402) );
  OAI22_X1 U1282 ( .A1(n5), .A2(n885), .B1(n837), .B2(n4), .ZN(n573) );
  OR2_X1 U1283 ( .A1(n1067), .A2(n885), .ZN(n837) );
  INV_X1 U1284 ( .A(n1023), .ZN(n885) );
  OAI22_X1 U1285 ( .A1(n5), .A2(n836), .B1(n835), .B2(n3), .ZN(n701) );
  BUF_X1 U1286 ( .A(n874), .Z(n22) );
  BUF_X1 U1287 ( .A(n875), .Z(n16) );
  BUF_X1 U1288 ( .A(n868), .Z(n11) );
  BUF_X1 U1289 ( .A(n874), .Z(n21) );
  OAI22_X1 U1290 ( .A1(n48), .A2(n712), .B1(n1039), .B2(n711), .ZN(n583) );
  INV_X1 U1291 ( .A(n557), .ZN(n654) );
  INV_X1 U1292 ( .A(n31), .ZN(n880) );
  INV_X1 U1293 ( .A(n37), .ZN(n879) );
  INV_X1 U1294 ( .A(n43), .ZN(n878) );
  INV_X1 U1295 ( .A(n983), .ZN(n881) );
  INV_X1 U1296 ( .A(n1046), .ZN(n882) );
  XNOR2_X1 U1297 ( .A(a[9]), .B(a[10]), .ZN(n872) );
  XNOR2_X1 U1298 ( .A(a[12]), .B(a[11]), .ZN(n871) );
  XNOR2_X1 U1299 ( .A(a[14]), .B(a[13]), .ZN(n870) );
  XNOR2_X1 U1300 ( .A(a[8]), .B(a[7]), .ZN(n873) );
  BUF_X1 U1301 ( .A(b[14]), .Z(n839) );
  BUF_X1 U1302 ( .A(b[9]), .Z(n844) );
  BUF_X1 U1303 ( .A(b[8]), .Z(n845) );
  INV_X1 U1304 ( .A(a[0]), .ZN(n877) );
  OAI22_X1 U1305 ( .A1(n35), .A2(n737), .B1(n34), .B2(n736), .ZN(n348) );
  INV_X1 U1306 ( .A(n348), .ZN(n349) );
  INV_X1 U1307 ( .A(n168), .ZN(n167) );
  NOR2_X1 U1308 ( .A1(n364), .A2(n357), .ZN(n168) );
  INV_X1 U1309 ( .A(n402), .ZN(n403) );
  INV_X1 U1310 ( .A(n13), .ZN(n883) );
  OAI22_X1 U1311 ( .A1(n17), .A2(n799), .B1(n15), .B2(n798), .ZN(n665) );
  OAI22_X1 U1312 ( .A1(n18), .A2(n798), .B1(n15), .B2(n797), .ZN(n664) );
  OAI22_X1 U1313 ( .A1(n17), .A2(n797), .B1(n15), .B2(n796), .ZN(n663) );
  OAI22_X1 U1314 ( .A1(n18), .A2(n801), .B1(n15), .B2(n800), .ZN(n667) );
  OAI22_X1 U1315 ( .A1(n18), .A2(n800), .B1(n15), .B2(n799), .ZN(n666) );
  OAI22_X1 U1316 ( .A1(n17), .A2(n795), .B1(n15), .B2(n794), .ZN(n661) );
  OAI22_X1 U1317 ( .A1(n18), .A2(n802), .B1(n15), .B2(n801), .ZN(n668) );
  OR2_X1 U1318 ( .A1(n1068), .A2(n883), .ZN(n803) );
  OAI22_X1 U1319 ( .A1(n18), .A2(n796), .B1(n15), .B2(n795), .ZN(n662) );
  OAI22_X1 U1320 ( .A1(n23), .A2(n778), .B1(n21), .B2(n777), .ZN(n645) );
  OAI22_X1 U1321 ( .A1(n23), .A2(n779), .B1(n21), .B2(n778), .ZN(n646) );
  OAI22_X1 U1322 ( .A1(n23), .A2(n780), .B1(n21), .B2(n779), .ZN(n647) );
  OAI22_X1 U1323 ( .A1(n23), .A2(n781), .B1(n21), .B2(n780), .ZN(n648) );
  OAI22_X1 U1324 ( .A1(n23), .A2(n782), .B1(n21), .B2(n781), .ZN(n649) );
  OAI22_X1 U1325 ( .A1(n23), .A2(n783), .B1(n21), .B2(n782), .ZN(n650) );
  OAI22_X1 U1326 ( .A1(n23), .A2(n784), .B1(n21), .B2(n783), .ZN(n651) );
  OAI22_X1 U1327 ( .A1(n23), .A2(n785), .B1(n21), .B2(n784), .ZN(n652) );
  INV_X1 U1328 ( .A(n21), .ZN(n555) );
  AOI21_X1 U1329 ( .B1(n24), .B2(n22), .A(n770), .ZN(n554) );
  OAI22_X1 U1330 ( .A1(n24), .A2(n772), .B1(n22), .B2(n771), .ZN(n639) );
  OAI22_X1 U1331 ( .A1(n24), .A2(n773), .B1(n22), .B2(n772), .ZN(n640) );
  OAI22_X1 U1332 ( .A1(n24), .A2(n774), .B1(n22), .B2(n773), .ZN(n641) );
  OAI22_X1 U1333 ( .A1(n24), .A2(n775), .B1(n22), .B2(n774), .ZN(n642) );
  OAI22_X1 U1334 ( .A1(n24), .A2(n776), .B1(n22), .B2(n775), .ZN(n643) );
  OAI22_X1 U1335 ( .A1(n24), .A2(n777), .B1(n22), .B2(n776), .ZN(n644) );
  CLKBUF_X1 U1336 ( .A(b[15]), .Z(n1066) );
  NOR2_X1 U1337 ( .A1(n190), .A2(n153), .ZN(n151) );
  OAI22_X1 U1338 ( .A1(n41), .A2(n733), .B1(n39), .B2(n732), .ZN(n603) );
  OAI22_X1 U1339 ( .A1(n41), .A2(n732), .B1(n39), .B2(n731), .ZN(n602) );
  OAI22_X1 U1340 ( .A1(n734), .A2(n42), .B1(n40), .B2(n733), .ZN(n604) );
  OAI22_X1 U1341 ( .A1(n41), .A2(n731), .B1(n39), .B2(n730), .ZN(n601) );
  OAI22_X1 U1342 ( .A1(n41), .A2(n727), .B1(n39), .B2(n726), .ZN(n597) );
  OAI22_X1 U1343 ( .A1(n42), .A2(n730), .B1(n729), .B2(n39), .ZN(n600) );
  OAI22_X1 U1344 ( .A1(n42), .A2(n729), .B1(n40), .B2(n728), .ZN(n599) );
  XNOR2_X1 U1345 ( .A(a[6]), .B(a[5]), .ZN(n874) );
  INV_X1 U1346 ( .A(n560), .ZN(n670) );
  XNOR2_X1 U1347 ( .A(a[1]), .B(a[2]), .ZN(n876) );
  INV_X1 U1348 ( .A(n182), .ZN(n180) );
  OAI22_X1 U1349 ( .A1(n17), .A2(n793), .B1(n16), .B2(n792), .ZN(n659) );
  OAI22_X1 U1350 ( .A1(n17), .A2(n792), .B1(n16), .B2(n791), .ZN(n658) );
  OAI22_X1 U1351 ( .A1(n1060), .A2(n794), .B1(n16), .B2(n793), .ZN(n660) );
  OAI22_X1 U1352 ( .A1(n1060), .A2(n791), .B1(n16), .B2(n790), .ZN(n657) );
  OAI22_X1 U1353 ( .A1(n1060), .A2(n790), .B1(n16), .B2(n789), .ZN(n656) );
  OAI22_X1 U1354 ( .A1(n17), .A2(n883), .B1(n803), .B2(n16), .ZN(n571) );
  AOI21_X1 U1355 ( .B1(n18), .B2(n16), .A(n787), .ZN(n557) );
  OAI22_X1 U1356 ( .A1(n1060), .A2(n789), .B1(n16), .B2(n788), .ZN(n655) );
  AOI21_X1 U1357 ( .B1(n1022), .B2(n4), .A(n821), .ZN(n563) );
  OAI22_X1 U1358 ( .A1(n48), .A2(n709), .B1(n1039), .B2(n708), .ZN(n580) );
  INV_X1 U1359 ( .A(n296), .ZN(n294) );
  OAI22_X1 U1360 ( .A1(n964), .A2(n834), .B1(n833), .B2(n3), .ZN(n699) );
  INV_X1 U1361 ( .A(n157), .ZN(n308) );
  AOI21_X1 U1362 ( .B1(n1009), .B2(n1028), .A(n244), .ZN(n242) );
  OAI21_X1 U1363 ( .B1(n276), .B2(n274), .A(n275), .ZN(n273) );
  NAND2_X1 U1364 ( .A1(n519), .A2(n524), .ZN(n275) );
  OAI22_X1 U1365 ( .A1(n24), .A2(n882), .B1(n786), .B2(n22), .ZN(n570) );
  XNOR2_X1 U1366 ( .A(n1046), .B(n1067), .ZN(n785) );
  OR2_X1 U1367 ( .A1(n1067), .A2(n882), .ZN(n786) );
  XNOR2_X1 U1368 ( .A(n1046), .B(n852), .ZN(n784) );
  XNOR2_X1 U1369 ( .A(n1046), .B(n845), .ZN(n777) );
  XNOR2_X1 U1370 ( .A(n1046), .B(n851), .ZN(n783) );
  XNOR2_X1 U1371 ( .A(n1046), .B(n844), .ZN(n776) );
  XNOR2_X1 U1372 ( .A(n1046), .B(n848), .ZN(n780) );
  XNOR2_X1 U1373 ( .A(n1046), .B(n846), .ZN(n778) );
  XNOR2_X1 U1374 ( .A(n1046), .B(n1018), .ZN(n782) );
  XNOR2_X1 U1375 ( .A(n1046), .B(n847), .ZN(n779) );
  XNOR2_X1 U1376 ( .A(n1046), .B(n849), .ZN(n781) );
  XNOR2_X1 U1377 ( .A(n1046), .B(n843), .ZN(n775) );
  XNOR2_X1 U1378 ( .A(n19), .B(n842), .ZN(n774) );
  XNOR2_X1 U1379 ( .A(n1046), .B(n839), .ZN(n771) );
  XNOR2_X1 U1380 ( .A(n19), .B(n841), .ZN(n773) );
  XNOR2_X1 U1381 ( .A(n19), .B(n840), .ZN(n772) );
  XNOR2_X1 U1382 ( .A(n1046), .B(n1065), .ZN(n770) );
  XNOR2_X1 U1383 ( .A(n43), .B(n961), .ZN(n704) );
  XNOR2_X1 U1384 ( .A(n43), .B(n841), .ZN(n705) );
  XNOR2_X1 U1385 ( .A(n43), .B(n839), .ZN(n703) );
  XNOR2_X1 U1386 ( .A(n43), .B(n1065), .ZN(n702) );
  XNOR2_X1 U1387 ( .A(n43), .B(n842), .ZN(n706) );
  XNOR2_X1 U1388 ( .A(n43), .B(n1038), .ZN(n707) );
  XNOR2_X1 U1389 ( .A(n43), .B(n1068), .ZN(n717) );
  XNOR2_X1 U1390 ( .A(n43), .B(n844), .ZN(n708) );
  XNOR2_X1 U1391 ( .A(n43), .B(n852), .ZN(n716) );
  XNOR2_X1 U1392 ( .A(n43), .B(n851), .ZN(n715) );
  XNOR2_X1 U1393 ( .A(n43), .B(n847), .ZN(n711) );
  XNOR2_X1 U1394 ( .A(n43), .B(n846), .ZN(n710) );
  XNOR2_X1 U1395 ( .A(n43), .B(n845), .ZN(n709) );
  XNOR2_X1 U1396 ( .A(n43), .B(n1017), .ZN(n714) );
  XNOR2_X1 U1397 ( .A(n43), .B(n849), .ZN(n713) );
  XNOR2_X1 U1398 ( .A(n43), .B(n848), .ZN(n712) );
  INV_X1 U1399 ( .A(n1042), .ZN(n254) );
  XNOR2_X1 U1400 ( .A(n984), .B(n1067), .ZN(n768) );
  XNOR2_X1 U1401 ( .A(n984), .B(n852), .ZN(n767) );
  XNOR2_X1 U1402 ( .A(n983), .B(n847), .ZN(n762) );
  XNOR2_X1 U1403 ( .A(n984), .B(n848), .ZN(n763) );
  XNOR2_X1 U1404 ( .A(n983), .B(n1065), .ZN(n753) );
  XNOR2_X1 U1405 ( .A(n982), .B(n846), .ZN(n761) );
  XNOR2_X1 U1406 ( .A(n984), .B(n849), .ZN(n764) );
  XNOR2_X1 U1407 ( .A(n983), .B(n851), .ZN(n766) );
  XNOR2_X1 U1408 ( .A(n983), .B(n845), .ZN(n760) );
  XNOR2_X1 U1409 ( .A(n984), .B(n1018), .ZN(n765) );
  XNOR2_X1 U1410 ( .A(n983), .B(n841), .ZN(n756) );
  XNOR2_X1 U1411 ( .A(n982), .B(n844), .ZN(n759) );
  XNOR2_X1 U1412 ( .A(n983), .B(n839), .ZN(n754) );
  XNOR2_X1 U1413 ( .A(n984), .B(n961), .ZN(n755) );
  XNOR2_X1 U1414 ( .A(n984), .B(n843), .ZN(n758) );
  XNOR2_X1 U1415 ( .A(n982), .B(n842), .ZN(n757) );
  XNOR2_X1 U1416 ( .A(n1031), .B(n961), .ZN(n721) );
  XNOR2_X1 U1417 ( .A(n1031), .B(n839), .ZN(n720) );
  XNOR2_X1 U1418 ( .A(n1031), .B(n1066), .ZN(n719) );
  XNOR2_X1 U1419 ( .A(n1031), .B(n841), .ZN(n722) );
  XNOR2_X1 U1420 ( .A(n37), .B(n851), .ZN(n732) );
  XNOR2_X1 U1421 ( .A(n37), .B(n1068), .ZN(n734) );
  XNOR2_X1 U1422 ( .A(n37), .B(n1018), .ZN(n731) );
  XNOR2_X1 U1423 ( .A(n37), .B(n842), .ZN(n723) );
  XNOR2_X1 U1424 ( .A(n37), .B(n852), .ZN(n733) );
  XNOR2_X1 U1425 ( .A(n37), .B(n845), .ZN(n726) );
  XNOR2_X1 U1426 ( .A(n849), .B(n37), .ZN(n730) );
  XNOR2_X1 U1427 ( .A(n37), .B(n844), .ZN(n725) );
  XNOR2_X1 U1428 ( .A(n37), .B(n843), .ZN(n724) );
  XNOR2_X1 U1429 ( .A(n37), .B(n848), .ZN(n729) );
  XNOR2_X1 U1430 ( .A(n37), .B(n847), .ZN(n728) );
  XNOR2_X1 U1431 ( .A(n37), .B(n846), .ZN(n727) );
  NAND2_X1 U1432 ( .A1(n459), .A2(n470), .ZN(n239) );
  AOI21_X1 U1433 ( .B1(n234), .B2(n230), .A(n231), .ZN(n229) );
  AOI21_X1 U1434 ( .B1(n234), .B2(n1056), .A(n980), .ZN(n220) );
  XNOR2_X1 U1435 ( .A(n7), .B(n841), .ZN(n807) );
  XNOR2_X1 U1436 ( .A(n7), .B(n848), .ZN(n814) );
  XNOR2_X1 U1437 ( .A(n7), .B(n847), .ZN(n813) );
  XNOR2_X1 U1438 ( .A(n7), .B(n846), .ZN(n812) );
  XNOR2_X1 U1439 ( .A(n7), .B(n845), .ZN(n811) );
  XNOR2_X1 U1440 ( .A(n7), .B(n1018), .ZN(n816) );
  XNOR2_X1 U1441 ( .A(n7), .B(n849), .ZN(n815) );
  XNOR2_X1 U1442 ( .A(n7), .B(n842), .ZN(n808) );
  XNOR2_X1 U1443 ( .A(n7), .B(n844), .ZN(n810) );
  XNOR2_X1 U1444 ( .A(n7), .B(n961), .ZN(n806) );
  XNOR2_X1 U1445 ( .A(n7), .B(n843), .ZN(n809) );
  XNOR2_X1 U1446 ( .A(n7), .B(n851), .ZN(n817) );
  XNOR2_X1 U1447 ( .A(n7), .B(n1067), .ZN(n819) );
  XNOR2_X1 U1448 ( .A(n7), .B(n852), .ZN(n818) );
  XNOR2_X1 U1449 ( .A(n7), .B(n839), .ZN(n805) );
  XNOR2_X1 U1450 ( .A(n7), .B(n1066), .ZN(n804) );
  OAI21_X1 U1451 ( .B1(n1050), .B2(n219), .A(n212), .ZN(n210) );
  NAND2_X1 U1452 ( .A1(n861), .A2(n877), .ZN(n869) );
  NAND2_X1 U1453 ( .A1(n855), .A2(n871), .ZN(n863) );
  OAI22_X1 U1454 ( .A1(n41), .A2(n728), .B1(n727), .B2(n39), .ZN(n598) );
  AOI21_X1 U1455 ( .B1(n236), .B2(n255), .A(n237), .ZN(n235) );
  OAI21_X1 U1456 ( .B1(n256), .B2(n268), .A(n257), .ZN(n255) );
  NOR2_X1 U1457 ( .A1(n218), .A2(n211), .ZN(n209) );
  INV_X1 U1458 ( .A(n1048), .ZN(n315) );
  AOI21_X1 U1459 ( .B1(n214), .B2(n234), .A(n215), .ZN(n213) );
  NOR2_X1 U1460 ( .A1(n417), .A2(n430), .ZN(n218) );
  NAND2_X1 U1461 ( .A1(n858), .A2(n874), .ZN(n866) );
  NOR2_X1 U1462 ( .A1(n241), .A2(n238), .ZN(n236) );
  OAI22_X1 U1463 ( .A1(n47), .A2(n713), .B1(n1039), .B2(n712), .ZN(n584) );
  AOI21_X1 U1464 ( .B1(n1044), .B2(n28), .A(n753), .ZN(n551) );
  OAI22_X1 U1465 ( .A1(n29), .A2(n759), .B1(n28), .B2(n758), .ZN(n627) );
  OAI22_X1 U1466 ( .A1(n1044), .A2(n757), .B1(n28), .B2(n756), .ZN(n625) );
  OAI22_X1 U1467 ( .A1(n1043), .A2(n881), .B1(n769), .B2(n28), .ZN(n569) );
  OAI22_X1 U1468 ( .A1(n1044), .A2(n756), .B1(n28), .B2(n755), .ZN(n624) );
  OAI22_X1 U1469 ( .A1(n1044), .A2(n755), .B1(n28), .B2(n754), .ZN(n623) );
  OAI22_X1 U1470 ( .A1(n1044), .A2(n760), .B1(n28), .B2(n759), .ZN(n628) );
  OAI22_X1 U1471 ( .A1(n29), .A2(n758), .B1(n28), .B2(n757), .ZN(n626) );
  OAI21_X1 U1472 ( .B1(n254), .B2(n241), .A(n959), .ZN(n240) );
  OAI21_X1 U1473 ( .B1(n242), .B2(n238), .A(n239), .ZN(n237) );
  XNOR2_X1 U1474 ( .A(n31), .B(n961), .ZN(n738) );
  XNOR2_X1 U1475 ( .A(n31), .B(n1038), .ZN(n741) );
  XNOR2_X1 U1476 ( .A(n849), .B(n31), .ZN(n747) );
  XNOR2_X1 U1477 ( .A(n31), .B(n842), .ZN(n740) );
  XNOR2_X1 U1478 ( .A(n848), .B(n31), .ZN(n746) );
  XNOR2_X1 U1479 ( .A(n31), .B(n839), .ZN(n737) );
  XNOR2_X1 U1480 ( .A(n31), .B(n841), .ZN(n739) );
  XNOR2_X1 U1481 ( .A(n31), .B(n847), .ZN(n745) );
  XNOR2_X1 U1482 ( .A(n31), .B(n851), .ZN(n749) );
  XNOR2_X1 U1483 ( .A(n31), .B(n1017), .ZN(n748) );
  XNOR2_X1 U1484 ( .A(n31), .B(n1066), .ZN(n736) );
  XNOR2_X1 U1485 ( .A(n31), .B(n1068), .ZN(n751) );
  XNOR2_X1 U1486 ( .A(n31), .B(n852), .ZN(n750) );
  XNOR2_X1 U1487 ( .A(n31), .B(n845), .ZN(n743) );
  XNOR2_X1 U1488 ( .A(n31), .B(n844), .ZN(n742) );
  OAI22_X1 U1489 ( .A1(n1043), .A2(n766), .B1(n28), .B2(n765), .ZN(n634) );
  INV_X1 U1490 ( .A(n246), .ZN(n244) );
  NAND2_X1 U1491 ( .A1(n1009), .A2(n246), .ZN(n71) );
  AOI21_X1 U1492 ( .B1(n981), .B2(n226), .A(n210), .ZN(n208) );
  XNOR2_X1 U1493 ( .A(a[4]), .B(a[3]), .ZN(n875) );
  NAND2_X1 U1494 ( .A1(n859), .A2(n875), .ZN(n867) );
  NAND2_X1 U1495 ( .A1(n857), .A2(n873), .ZN(n865) );
  INV_X1 U1496 ( .A(n1061), .ZN(n234) );
  NAND2_X1 U1497 ( .A1(n357), .A2(n364), .ZN(n169) );
  NOR2_X1 U1498 ( .A1(n227), .A2(n232), .ZN(n225) );
  NAND2_X1 U1499 ( .A1(n431), .A2(n444), .ZN(n228) );
  XNOR2_X1 U1500 ( .A(n1023), .B(n845), .ZN(n828) );
  XNOR2_X1 U1501 ( .A(n1), .B(n840), .ZN(n823) );
  XNOR2_X1 U1502 ( .A(n1), .B(n839), .ZN(n822) );
  XNOR2_X1 U1503 ( .A(n1), .B(n841), .ZN(n824) );
  XNOR2_X1 U1504 ( .A(n1023), .B(n1067), .ZN(n836) );
  XNOR2_X1 U1505 ( .A(n1023), .B(n844), .ZN(n827) );
  XNOR2_X1 U1506 ( .A(n1023), .B(n848), .ZN(n831) );
  XNOR2_X1 U1507 ( .A(n1), .B(n842), .ZN(n825) );
  XNOR2_X1 U1508 ( .A(n1023), .B(n843), .ZN(n826) );
  XNOR2_X1 U1509 ( .A(n1), .B(n1065), .ZN(n821) );
  XNOR2_X1 U1510 ( .A(n1023), .B(n846), .ZN(n829) );
  XNOR2_X1 U1511 ( .A(n1023), .B(n847), .ZN(n830) );
  XNOR2_X1 U1512 ( .A(n1023), .B(n849), .ZN(n832) );
  XNOR2_X1 U1513 ( .A(n1023), .B(n852), .ZN(n835) );
  XNOR2_X1 U1514 ( .A(n1023), .B(n1018), .ZN(n833) );
  XNOR2_X1 U1515 ( .A(n1023), .B(n851), .ZN(n834) );
  BUF_X2 U1516 ( .A(n862), .Z(n48) );
  OAI22_X1 U1517 ( .A1(n47), .A2(n714), .B1(n1039), .B2(n713), .ZN(n585) );
  NAND2_X1 U1518 ( .A1(n854), .A2(n870), .ZN(n862) );
  INV_X1 U1519 ( .A(n362), .ZN(n363) );
  OAI22_X1 U1520 ( .A1(n1043), .A2(n754), .B1(n28), .B2(n753), .ZN(n362) );
  XOR2_X1 U1521 ( .A(n93), .B(n54), .Z(product[30]) );
  OAI21_X1 U1522 ( .B1(n150), .B2(n109), .A(n110), .ZN(n108) );
  XNOR2_X1 U1523 ( .A(n1040), .B(n75), .ZN(product[9]) );
  XNOR2_X1 U1524 ( .A(n13), .B(n849), .ZN(n798) );
  XNOR2_X1 U1525 ( .A(n13), .B(n848), .ZN(n797) );
  XNOR2_X1 U1526 ( .A(n13), .B(n843), .ZN(n792) );
  XNOR2_X1 U1527 ( .A(n13), .B(n841), .ZN(n790) );
  XNOR2_X1 U1528 ( .A(n13), .B(n842), .ZN(n791) );
  XNOR2_X1 U1529 ( .A(n13), .B(n840), .ZN(n789) );
  XNOR2_X1 U1530 ( .A(n13), .B(n851), .ZN(n800) );
  XNOR2_X1 U1531 ( .A(n13), .B(n1018), .ZN(n799) );
  XNOR2_X1 U1532 ( .A(n13), .B(n845), .ZN(n794) );
  XNOR2_X1 U1533 ( .A(n13), .B(n844), .ZN(n793) );
  XNOR2_X1 U1534 ( .A(n13), .B(n1068), .ZN(n802) );
  XNOR2_X1 U1535 ( .A(n13), .B(n852), .ZN(n801) );
  XNOR2_X1 U1536 ( .A(n13), .B(n847), .ZN(n796) );
  XNOR2_X1 U1537 ( .A(n13), .B(n846), .ZN(n795) );
  XNOR2_X1 U1538 ( .A(n13), .B(n839), .ZN(n788) );
  OAI21_X1 U1539 ( .B1(n150), .B2(n133), .A(n134), .ZN(n132) );
  XOR2_X1 U1540 ( .A(n117), .B(n56), .Z(product[28]) );
  OAI21_X1 U1541 ( .B1(n150), .B2(n124), .A(n125), .ZN(n119) );
  OAI21_X1 U1542 ( .B1(n150), .B2(n144), .A(n145), .ZN(n141) );
  NOR2_X1 U1543 ( .A1(n204), .A2(n199), .ZN(n197) );
  NAND2_X1 U1544 ( .A1(n856), .A2(n872), .ZN(n864) );
  NAND2_X1 U1545 ( .A1(n365), .A2(n372), .ZN(n182) );
  NOR2_X1 U1546 ( .A1(n168), .A2(n157), .ZN(n155) );
  OAI21_X1 U1547 ( .B1(n157), .B2(n169), .A(n158), .ZN(n156) );
  NAND2_X1 U1548 ( .A1(n351), .A2(n356), .ZN(n158) );
  XOR2_X1 U1549 ( .A(a[14]), .B(a[15]), .Z(n854) );
  AOI21_X1 U1550 ( .B1(n1035), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U1551 ( .B1(n1034), .B2(n118), .A(n119), .ZN(n117) );
  AOI21_X1 U1552 ( .B1(n1034), .B2(n94), .A(n95), .ZN(n93) );
  AOI21_X1 U1553 ( .B1(n1034), .B2(n140), .A(n141), .ZN(n139) );
  AOI21_X1 U1554 ( .B1(n1034), .B2(n131), .A(n132), .ZN(n130) );
  AOI21_X1 U1555 ( .B1(n1034), .B2(n160), .A(n161), .ZN(n159) );
  AOI21_X1 U1556 ( .B1(n1034), .B2(n313), .A(n203), .ZN(n201) );
  AOI21_X1 U1557 ( .B1(n51), .B2(n184), .A(n185), .ZN(n183) );
  AOI21_X1 U1558 ( .B1(n51), .B2(n171), .A(n172), .ZN(n170) );
  AOI21_X1 U1559 ( .B1(n51), .B2(n193), .A(n194), .ZN(n192) );
  XNOR2_X1 U1560 ( .A(n1035), .B(n65), .ZN(product[19]) );
  XOR2_X1 U1561 ( .A(a[12]), .B(a[13]), .Z(n855) );
  XOR2_X1 U1562 ( .A(a[6]), .B(a[7]), .Z(n858) );
  NAND2_X1 U1563 ( .A1(n860), .A2(n876), .ZN(n868) );
  NAND2_X1 U1564 ( .A1(n155), .A2(n1032), .ZN(n153) );
  AOI21_X1 U1565 ( .B1(n155), .B2(n180), .A(n156), .ZN(n154) );
  AOI21_X1 U1566 ( .B1(n1035), .B2(n147), .A(n148), .ZN(n146) );
  OAI21_X1 U1567 ( .B1(n207), .B2(n235), .A(n208), .ZN(n206) );
  NAND2_X1 U1568 ( .A1(n209), .A2(n225), .ZN(n207) );
  XOR2_X1 U1569 ( .A(a[8]), .B(a[9]), .Z(n857) );
  XOR2_X1 U1570 ( .A(a[11]), .B(a[10]), .Z(n856) );
  NAND2_X1 U1571 ( .A1(n471), .A2(n482), .ZN(n246) );
  XOR2_X1 U1572 ( .A(a[2]), .B(a[3]), .Z(n860) );
  OAI21_X1 U1573 ( .B1(n153), .B2(n191), .A(n154), .ZN(n152) );
  XOR2_X1 U1574 ( .A(n106), .B(n55), .Z(product[29]) );
  AOI21_X1 U1575 ( .B1(n1035), .B2(n107), .A(n108), .ZN(n106) );
  NAND2_X1 U1576 ( .A1(n541), .A2(n572), .ZN(n296) );
  XOR2_X1 U1577 ( .A(a[4]), .B(a[5]), .Z(n859) );
  XOR2_X1 U1578 ( .A(n963), .B(n76), .Z(product[8]) );
  XNOR2_X1 U1579 ( .A(n281), .B(n77), .ZN(product[7]) );
  AOI21_X1 U1580 ( .B1(n281), .B2(n1014), .A(n278), .ZN(n276) );
  XOR2_X1 U1581 ( .A(n78), .B(n1019), .Z(product[6]) );
  OAI21_X1 U1582 ( .B1(n284), .B2(n282), .A(n283), .ZN(n281) );
  XOR2_X1 U1583 ( .A(a[1]), .B(a[0]), .Z(n861) );
endmodule


module datapath_DW_mult_tc_13 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n16, n17, n18, n19,
         n21, n22, n23, n24, n25, n28, n29, n30, n31, n33, n34, n35, n37, n39,
         n40, n41, n42, n43, n45, n46, n47, n48, n49, n51, n54, n55, n56, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n84, n85, n86, n87, n88, n90, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n103, n105, n106, n107, n108, n109, n110,
         n114, n116, n117, n118, n119, n122, n123, n124, n125, n127, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n168, n169, n170, n171, n172, n173, n174, n175,
         n177, n178, n180, n182, n183, n184, n185, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n223, n224, n225, n226, n227,
         n228, n229, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n246, n247, n248, n249, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n264, n266, n267, n268, n270, n272,
         n273, n274, n275, n276, n278, n280, n281, n282, n283, n284, n286,
         n288, n289, n290, n291, n292, n294, n296, n297, n298, n299, n301,
         n306, n308, n312, n313, n316, n317, n321, n324, n326, n328, n330,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n545, n546, n548, n549, n551, n552, n554, n555, n557,
         n558, n560, n561, n563, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1068, n1069;
  assign product[31] = n84;

  FA_X1 U364 ( .A(n575), .B(n338), .CI(n590), .CO(n334), .S(n335) );
  FA_X1 U365 ( .A(n339), .B(n576), .CI(n342), .CO(n336), .S(n337) );
  FA_X1 U367 ( .A(n346), .B(n577), .CI(n343), .CO(n340), .S(n341) );
  FA_X1 U368 ( .A(n591), .B(n348), .CI(n606), .CO(n342), .S(n343) );
  FA_X1 U369 ( .A(n347), .B(n354), .CI(n352), .CO(n344), .S(n345) );
  FA_X1 U370 ( .A(n578), .B(n592), .CI(n349), .CO(n346), .S(n347) );
  FA_X1 U372 ( .A(n358), .B(n355), .CI(n353), .CO(n350), .S(n351) );
  FA_X1 U373 ( .A(n362), .B(n607), .CI(n360), .CO(n352), .S(n353) );
  FA_X1 U374 ( .A(n593), .B(n579), .CI(n622), .CO(n354), .S(n355) );
  FA_X1 U375 ( .A(n359), .B(n361), .CI(n366), .CO(n356), .S(n357) );
  FA_X1 U376 ( .A(n370), .B(n363), .CI(n368), .CO(n358), .S(n359) );
  FA_X1 U377 ( .A(n580), .B(n594), .CI(n608), .CO(n360), .S(n361) );
  FA_X1 U379 ( .A(n374), .B(n376), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U380 ( .A(n369), .B(n378), .CI(n371), .CO(n366), .S(n367) );
  FA_X1 U381 ( .A(n595), .B(n380), .CI(n609), .CO(n368), .S(n369) );
  FA_X1 U382 ( .A(n623), .B(n581), .CI(n638), .CO(n370), .S(n371) );
  FA_X1 U383 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  FA_X1 U384 ( .A(n379), .B(n388), .CI(n386), .CO(n374), .S(n375) );
  FA_X1 U385 ( .A(n381), .B(n610), .CI(n390), .CO(n376), .S(n377) );
  FA_X1 U386 ( .A(n624), .B(n596), .CI(n582), .CO(n378), .S(n379) );
  FA_X1 U388 ( .A(n394), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U390 ( .A(n400), .B(n625), .CI(n398), .CO(n386), .S(n387) );
  FA_X1 U391 ( .A(n597), .B(n639), .CI(n611), .CO(n388), .S(n389) );
  FA_X1 U392 ( .A(n654), .B(n583), .CI(n1026), .CO(n390), .S(n391) );
  FA_X1 U394 ( .A(n410), .B(n399), .CI(n408), .CO(n394), .S(n395) );
  FA_X1 U395 ( .A(n412), .B(n414), .CI(n401), .CO(n396), .S(n397) );
  FA_X1 U396 ( .A(n584), .B(n598), .CI(n403), .CO(n398), .S(n399) );
  FA_X1 U397 ( .A(n640), .B(n626), .CI(n612), .CO(n400), .S(n401) );
  FA_X1 U399 ( .A(n418), .B(n409), .CI(n407), .CO(n404), .S(n405) );
  FA_X1 U400 ( .A(n411), .B(n422), .CI(n420), .CO(n406), .S(n407) );
  FA_X1 U401 ( .A(n413), .B(n424), .CI(n415), .CO(n408), .S(n409) );
  FA_X1 U403 ( .A(n599), .B(n641), .CI(n655), .CO(n412), .S(n413) );
  FA_X1 U404 ( .A(n670), .B(n585), .CI(n428), .CO(n414), .S(n415) );
  FA_X1 U405 ( .A(n432), .B(n421), .CI(n419), .CO(n416), .S(n417) );
  FA_X1 U406 ( .A(n423), .B(n436), .CI(n434), .CO(n418), .S(n419) );
  FA_X1 U409 ( .A(n642), .B(n628), .CI(n600), .CO(n424), .S(n425) );
  FA_X1 U410 ( .A(n614), .B(n586), .CI(n656), .CO(n426), .S(n427) );
  FA_X1 U413 ( .A(n437), .B(n450), .CI(n448), .CO(n432), .S(n433) );
  FA_X1 U415 ( .A(n443), .B(n456), .CI(n454), .CO(n436), .S(n437) );
  FA_X1 U416 ( .A(n657), .B(n615), .CI(n671), .CO(n438), .S(n439) );
  FA_X1 U417 ( .A(n629), .B(n587), .CI(n686), .CO(n440), .S(n441) );
  FA_X1 U421 ( .A(n455), .B(n462), .CI(n451), .CO(n446), .S(n447) );
  FA_X1 U422 ( .A(n453), .B(n466), .CI(n464), .CO(n448), .S(n449) );
  FA_X1 U423 ( .A(n457), .B(n672), .CI(n468), .CO(n450), .S(n451) );
  FA_X1 U424 ( .A(n687), .B(n630), .CI(n658), .CO(n452), .S(n453) );
  FA_X1 U425 ( .A(n602), .B(n644), .CI(n616), .CO(n454), .S(n455) );
  HA_X1 U426 ( .A(n566), .B(n588), .CO(n456), .S(n457) );
  FA_X1 U427 ( .A(n463), .B(n472), .CI(n461), .CO(n458), .S(n459) );
  FA_X1 U428 ( .A(n465), .B(n467), .CI(n474), .CO(n460), .S(n461) );
  FA_X1 U430 ( .A(n645), .B(n659), .CI(n480), .CO(n464), .S(n465) );
  FA_X1 U431 ( .A(n603), .B(n673), .CI(n631), .CO(n466), .S(n467) );
  FA_X1 U432 ( .A(n617), .B(n589), .CI(n688), .CO(n468), .S(n469) );
  FA_X1 U434 ( .A(n479), .B(n477), .CI(n486), .CO(n472), .S(n473) );
  FA_X1 U435 ( .A(n490), .B(n481), .CI(n488), .CO(n474), .S(n475) );
  FA_X1 U437 ( .A(n689), .B(n646), .CI(n674), .CO(n478), .S(n479) );
  HA_X1 U438 ( .A(n604), .B(n567), .CO(n480), .S(n481) );
  FA_X1 U439 ( .A(n487), .B(n494), .CI(n485), .CO(n482), .S(n483) );
  FA_X1 U440 ( .A(n489), .B(n491), .CI(n496), .CO(n484), .S(n485) );
  FA_X1 U441 ( .A(n1003), .B(n661), .CI(n498), .CO(n486), .S(n487) );
  FA_X1 U442 ( .A(n619), .B(n647), .CI(n675), .CO(n488), .S(n489) );
  FA_X1 U443 ( .A(n690), .B(n605), .CI(n633), .CO(n490), .S(n491) );
  FA_X1 U444 ( .A(n504), .B(n497), .CI(n495), .CO(n492), .S(n493) );
  FA_X1 U445 ( .A(n506), .B(n508), .CI(n499), .CO(n494), .S(n495) );
  FA_X1 U446 ( .A(n648), .B(n676), .CI(n501), .CO(n496), .S(n497) );
  FA_X1 U447 ( .A(n662), .B(n634), .CI(n691), .CO(n498), .S(n499) );
  FA_X1 U449 ( .A(n512), .B(n507), .CI(n505), .CO(n502), .S(n503) );
  FA_X1 U450 ( .A(n514), .B(n516), .CI(n509), .CO(n504), .S(n505) );
  FA_X1 U451 ( .A(n635), .B(n677), .CI(n663), .CO(n506), .S(n507) );
  FA_X1 U452 ( .A(n649), .B(n621), .CI(n692), .CO(n508), .S(n509) );
  FA_X1 U453 ( .A(n515), .B(n520), .CI(n513), .CO(n510), .S(n511) );
  FA_X1 U454 ( .A(n517), .B(n693), .CI(n522), .CO(n512), .S(n513) );
  FA_X1 U455 ( .A(n650), .B(n664), .CI(n678), .CO(n514), .S(n515) );
  HA_X1 U456 ( .A(n569), .B(n636), .CO(n516), .S(n517) );
  FA_X1 U457 ( .A(n523), .B(n526), .CI(n521), .CO(n518), .S(n519) );
  FA_X1 U458 ( .A(n651), .B(n679), .CI(n528), .CO(n520), .S(n521) );
  FA_X1 U459 ( .A(n665), .B(n637), .CI(n694), .CO(n522), .S(n523) );
  FA_X1 U460 ( .A(n532), .B(n529), .CI(n527), .CO(n524), .S(n525) );
  FA_X1 U461 ( .A(n666), .B(n695), .CI(n680), .CO(n526), .S(n527) );
  HA_X1 U462 ( .A(n570), .B(n652), .CO(n528), .S(n529) );
  FA_X1 U463 ( .A(n536), .B(n667), .CI(n533), .CO(n530), .S(n531) );
  FA_X1 U464 ( .A(n696), .B(n653), .CI(n681), .CO(n532), .S(n533) );
  FA_X1 U465 ( .A(n682), .B(n697), .CI(n537), .CO(n534), .S(n535) );
  HA_X1 U466 ( .A(n668), .B(n571), .CO(n536), .S(n537) );
  FA_X1 U467 ( .A(n698), .B(n669), .CI(n683), .CO(n538), .S(n539) );
  HA_X1 U468 ( .A(n684), .B(n699), .CO(n540), .S(n541) );
  CLKBUF_X1 U822 ( .A(n459), .Z(n953) );
  BUF_X4 U823 ( .A(a[15]), .Z(n43) );
  CLKBUF_X3 U824 ( .A(n871), .Z(n39) );
  BUF_X2 U825 ( .A(n31), .Z(n954) );
  NOR2_X2 U826 ( .A1(n373), .A2(n382), .ZN(n190) );
  CLKBUF_X1 U827 ( .A(n425), .Z(n955) );
  NOR2_X1 U828 ( .A1(n459), .A2(n470), .ZN(n956) );
  CLKBUF_X3 U829 ( .A(b[3]), .Z(n850) );
  CLKBUF_X3 U830 ( .A(b[1]), .Z(n852) );
  BUF_X2 U831 ( .A(b[2]), .Z(n851) );
  CLKBUF_X3 U832 ( .A(b[11]), .Z(n842) );
  OAI21_X2 U833 ( .B1(n268), .B2(n256), .A(n257), .ZN(n255) );
  BUF_X2 U834 ( .A(b[10]), .Z(n843) );
  BUF_X2 U835 ( .A(n19), .Z(n1032) );
  OAI21_X1 U836 ( .B1(n282), .B2(n284), .A(n283), .ZN(n281) );
  BUF_X1 U837 ( .A(n866), .Z(n23) );
  AND2_X1 U838 ( .A1(n1007), .A2(n1008), .ZN(n150) );
  CLKBUF_X1 U839 ( .A(n225), .Z(n1063) );
  BUF_X1 U840 ( .A(n875), .Z(n16) );
  BUF_X2 U841 ( .A(n873), .Z(n1022) );
  BUF_X2 U842 ( .A(n872), .Z(n33) );
  AND2_X2 U843 ( .A1(n1007), .A2(n1008), .ZN(n957) );
  BUF_X2 U844 ( .A(n49), .Z(n1029) );
  BUF_X1 U845 ( .A(b[0]), .Z(n49) );
  XNOR2_X1 U846 ( .A(n440), .B(n958), .ZN(n423) );
  XNOR2_X1 U847 ( .A(n442), .B(n429), .ZN(n958) );
  XNOR2_X1 U848 ( .A(n146), .B(n959), .ZN(product[25]) );
  AND2_X1 U849 ( .A1(n143), .A2(n145), .ZN(n959) );
  BUF_X1 U850 ( .A(b[8]), .Z(n845) );
  XNOR2_X1 U851 ( .A(n473), .B(n960), .ZN(n471) );
  XNOR2_X1 U852 ( .A(n484), .B(n475), .ZN(n960) );
  AND2_X1 U853 ( .A1(n483), .A2(n492), .ZN(n1058) );
  BUF_X2 U854 ( .A(n864), .Z(n1023) );
  BUF_X1 U855 ( .A(a[7]), .Z(n19) );
  BUF_X2 U856 ( .A(n49), .Z(n1068) );
  BUF_X2 U857 ( .A(n863), .Z(n41) );
  BUF_X1 U858 ( .A(n864), .Z(n35) );
  OAI22_X1 U859 ( .A1(n48), .A2(n703), .B1(n46), .B2(n702), .ZN(n332) );
  NAND3_X1 U860 ( .A1(n970), .A2(n971), .A3(n972), .ZN(n476) );
  XOR2_X1 U861 ( .A(n391), .B(n389), .Z(n961) );
  XOR2_X1 U862 ( .A(n396), .B(n961), .Z(n385) );
  NAND2_X1 U863 ( .A1(n396), .A2(n391), .ZN(n962) );
  NAND2_X1 U864 ( .A1(n396), .A2(n389), .ZN(n963) );
  NAND2_X1 U865 ( .A1(n391), .A2(n389), .ZN(n964) );
  NAND3_X1 U866 ( .A1(n962), .A2(n963), .A3(n964), .ZN(n384) );
  XOR2_X1 U867 ( .A(n406), .B(n397), .Z(n965) );
  XOR2_X1 U868 ( .A(n395), .B(n965), .Z(n393) );
  NAND2_X1 U869 ( .A1(n395), .A2(n406), .ZN(n966) );
  NAND2_X1 U870 ( .A1(n395), .A2(n397), .ZN(n967) );
  NAND2_X1 U871 ( .A1(n406), .A2(n397), .ZN(n968) );
  NAND3_X1 U872 ( .A1(n966), .A2(n967), .A3(n968), .ZN(n392) );
  XOR2_X1 U873 ( .A(n618), .B(n660), .Z(n969) );
  XOR2_X1 U874 ( .A(n969), .B(n632), .Z(n477) );
  NAND2_X1 U875 ( .A1(n618), .A2(n660), .ZN(n970) );
  NAND2_X1 U876 ( .A1(n618), .A2(n632), .ZN(n971) );
  NAND2_X1 U877 ( .A1(n660), .A2(n632), .ZN(n972) );
  XOR2_X1 U878 ( .A(n478), .B(n469), .Z(n973) );
  XOR2_X1 U879 ( .A(n973), .B(n476), .Z(n463) );
  NAND2_X1 U880 ( .A1(n478), .A2(n469), .ZN(n974) );
  NAND2_X1 U881 ( .A1(n478), .A2(n476), .ZN(n975) );
  NAND2_X1 U882 ( .A1(n469), .A2(n476), .ZN(n976) );
  NAND3_X1 U883 ( .A1(n974), .A2(n975), .A3(n976), .ZN(n462) );
  XOR2_X1 U884 ( .A(n460), .B(n449), .Z(n977) );
  XOR2_X1 U885 ( .A(n447), .B(n977), .Z(n445) );
  NAND2_X1 U886 ( .A1(n447), .A2(n460), .ZN(n978) );
  NAND2_X1 U887 ( .A1(n447), .A2(n449), .ZN(n979) );
  NAND2_X1 U888 ( .A1(n460), .A2(n449), .ZN(n980) );
  NAND3_X1 U889 ( .A1(n978), .A2(n979), .A3(n980), .ZN(n444) );
  XOR2_X1 U890 ( .A(n627), .B(n613), .Z(n981) );
  XOR2_X1 U891 ( .A(n426), .B(n981), .Z(n411) );
  NAND2_X1 U892 ( .A1(n426), .A2(n627), .ZN(n982) );
  NAND2_X1 U893 ( .A1(n426), .A2(n613), .ZN(n983) );
  NAND2_X1 U894 ( .A1(n627), .A2(n613), .ZN(n984) );
  NAND3_X1 U895 ( .A1(n982), .A2(n983), .A3(n984), .ZN(n410) );
  NAND2_X1 U896 ( .A1(n440), .A2(n442), .ZN(n985) );
  NAND2_X1 U897 ( .A1(n440), .A2(n429), .ZN(n986) );
  NAND2_X1 U898 ( .A1(n442), .A2(n429), .ZN(n987) );
  NAND3_X1 U899 ( .A1(n985), .A2(n986), .A3(n987), .ZN(n422) );
  OR2_X2 U900 ( .A1(n643), .A2(n601), .ZN(n442) );
  NAND2_X1 U901 ( .A1(n473), .A2(n484), .ZN(n988) );
  NAND2_X1 U902 ( .A1(n473), .A2(n475), .ZN(n989) );
  NAND2_X1 U903 ( .A1(n484), .A2(n475), .ZN(n990) );
  NAND3_X1 U904 ( .A1(n988), .A2(n989), .A3(n990), .ZN(n470) );
  XOR2_X1 U905 ( .A(n441), .B(n452), .Z(n991) );
  XOR2_X1 U906 ( .A(n439), .B(n991), .Z(n435) );
  NAND2_X1 U907 ( .A1(n439), .A2(n441), .ZN(n992) );
  NAND2_X1 U908 ( .A1(n439), .A2(n452), .ZN(n993) );
  NAND2_X1 U909 ( .A1(n441), .A2(n452), .ZN(n994) );
  NAND3_X1 U910 ( .A1(n992), .A2(n993), .A3(n994), .ZN(n434) );
  OR2_X1 U911 ( .A1(n334), .A2(n333), .ZN(n995) );
  OR2_X1 U912 ( .A1(n337), .A2(n340), .ZN(n996) );
  OR2_X1 U913 ( .A1(n574), .A2(n332), .ZN(n997) );
  OR2_X1 U914 ( .A1(n541), .A2(n572), .ZN(n998) );
  OR2_X1 U915 ( .A1(n336), .A2(n335), .ZN(n999) );
  OR2_X1 U916 ( .A1(n511), .A2(n518), .ZN(n1000) );
  OR2_X1 U917 ( .A1(n525), .A2(n530), .ZN(n1001) );
  OR2_X1 U918 ( .A1(n535), .A2(n538), .ZN(n1002) );
  AND2_X1 U919 ( .A1(n568), .A2(n620), .ZN(n1003) );
  OR2_X1 U920 ( .A1(n701), .A2(n573), .ZN(n1004) );
  CLKBUF_X1 U921 ( .A(n276), .Z(n1005) );
  CLKBUF_X1 U922 ( .A(n11), .Z(n1006) );
  BUF_X1 U923 ( .A(n868), .Z(n11) );
  CLKBUF_X1 U924 ( .A(n876), .Z(n9) );
  NAND2_X1 U925 ( .A1(n198), .A2(n151), .ZN(n1007) );
  INV_X1 U926 ( .A(n152), .ZN(n1008) );
  CLKBUF_X1 U927 ( .A(n219), .Z(n1009) );
  BUF_X2 U928 ( .A(b[6]), .Z(n847) );
  FA_X1 U929 ( .A(n418), .B(n409), .CI(n407), .S(n1010) );
  OR2_X1 U930 ( .A1(n483), .A2(n492), .ZN(n1011) );
  BUF_X2 U931 ( .A(b[15]), .Z(n838) );
  OR2_X1 U932 ( .A1(n503), .A2(n510), .ZN(n1012) );
  XOR2_X1 U933 ( .A(n955), .B(n438), .Z(n1013) );
  XOR2_X1 U934 ( .A(n427), .B(n1013), .Z(n421) );
  NAND2_X1 U935 ( .A1(n427), .A2(n425), .ZN(n1014) );
  NAND2_X1 U936 ( .A1(n427), .A2(n438), .ZN(n1015) );
  NAND2_X1 U937 ( .A1(n425), .A2(n438), .ZN(n1016) );
  NAND3_X1 U938 ( .A1(n1014), .A2(n1015), .A3(n1016), .ZN(n420) );
  CLKBUF_X1 U939 ( .A(n875), .Z(n1024) );
  CLKBUF_X1 U940 ( .A(n875), .Z(n1025) );
  BUF_X2 U941 ( .A(b[4]), .Z(n849) );
  BUF_X2 U942 ( .A(n19), .Z(n1031) );
  BUF_X2 U943 ( .A(a[5]), .Z(n1019) );
  BUF_X1 U944 ( .A(n206), .Z(n51) );
  BUF_X2 U945 ( .A(b[12]), .Z(n841) );
  CLKBUF_X3 U946 ( .A(a[13]), .Z(n1043) );
  CLKBUF_X1 U947 ( .A(a[13]), .Z(n37) );
  BUF_X2 U948 ( .A(n863), .Z(n42) );
  BUF_X1 U949 ( .A(n865), .Z(n1034) );
  CLKBUF_X1 U950 ( .A(n865), .Z(n1033) );
  CLKBUF_X1 U951 ( .A(n865), .Z(n29) );
  OR2_X1 U952 ( .A1(n365), .A2(n372), .ZN(n1017) );
  AOI21_X1 U953 ( .B1(n255), .B2(n236), .A(n237), .ZN(n1018) );
  CLKBUF_X3 U954 ( .A(n862), .Z(n47) );
  CLKBUF_X1 U955 ( .A(a[5]), .Z(n13) );
  BUF_X2 U956 ( .A(b[9]), .Z(n844) );
  BUF_X2 U957 ( .A(n866), .Z(n24) );
  BUF_X1 U958 ( .A(n868), .Z(n1020) );
  BUF_X1 U959 ( .A(n868), .Z(n1021) );
  CLKBUF_X1 U960 ( .A(n868), .Z(n12) );
  OAI22_X1 U961 ( .A1(n18), .A2(n788), .B1(n1025), .B2(n787), .ZN(n1026) );
  XNOR2_X1 U962 ( .A(n25), .B(n851), .ZN(n1027) );
  CLKBUF_X3 U963 ( .A(a[1]), .Z(n1028) );
  CLKBUF_X1 U964 ( .A(a[1]), .Z(n1) );
  OR2_X2 U965 ( .A1(n471), .A2(n482), .ZN(n1066) );
  CLKBUF_X1 U966 ( .A(n19), .Z(n1030) );
  INV_X1 U967 ( .A(n1059), .ZN(n246) );
  AND2_X1 U968 ( .A1(n471), .A2(n482), .ZN(n1059) );
  NOR2_X1 U969 ( .A1(n218), .A2(n211), .ZN(n1035) );
  CLKBUF_X1 U970 ( .A(n841), .Z(n1036) );
  OR2_X1 U971 ( .A1(n953), .A2(n470), .ZN(n1037) );
  CLKBUF_X1 U972 ( .A(n284), .Z(n1038) );
  XNOR2_X1 U973 ( .A(n201), .B(n1039), .ZN(product[20]) );
  AND2_X1 U974 ( .A1(n312), .A2(n200), .ZN(n1039) );
  XNOR2_X1 U975 ( .A(n433), .B(n1040), .ZN(n431) );
  XNOR2_X1 U976 ( .A(n446), .B(n435), .ZN(n1040) );
  XNOR2_X1 U977 ( .A(n159), .B(n1041), .ZN(product[24]) );
  AND2_X1 U978 ( .A1(n308), .A2(n158), .ZN(n1041) );
  NOR2_X1 U979 ( .A1(n405), .A2(n416), .ZN(n1042) );
  XNOR2_X1 U980 ( .A(n130), .B(n1044), .ZN(product[27]) );
  AND2_X1 U981 ( .A1(n996), .A2(n129), .ZN(n1044) );
  XNOR2_X1 U982 ( .A(n139), .B(n1045), .ZN(product[26]) );
  AND2_X1 U983 ( .A1(n306), .A2(n138), .ZN(n1045) );
  AOI21_X1 U984 ( .B1(n1066), .B2(n1058), .A(n1059), .ZN(n1046) );
  XNOR2_X1 U985 ( .A(n192), .B(n1047), .ZN(product[21]) );
  AND2_X1 U986 ( .A1(n188), .A2(n191), .ZN(n1047) );
  BUF_X1 U987 ( .A(n869), .Z(n1048) );
  BUF_X1 U988 ( .A(n869), .Z(n1049) );
  BUF_X4 U989 ( .A(a[11]), .Z(n31) );
  XNOR2_X1 U990 ( .A(n183), .B(n1050), .ZN(product[22]) );
  AND2_X1 U991 ( .A1(n175), .A2(n182), .ZN(n1050) );
  OR2_X1 U992 ( .A1(n357), .A2(n364), .ZN(n1051) );
  BUF_X2 U993 ( .A(n206), .Z(n1052) );
  CLKBUF_X1 U994 ( .A(n843), .Z(n1053) );
  CLKBUF_X1 U995 ( .A(n273), .Z(n1054) );
  NAND2_X1 U996 ( .A1(n433), .A2(n446), .ZN(n1055) );
  NAND2_X1 U997 ( .A1(n433), .A2(n435), .ZN(n1056) );
  NAND2_X1 U998 ( .A1(n446), .A2(n435), .ZN(n1057) );
  NAND3_X1 U999 ( .A1(n1055), .A2(n1056), .A3(n1057), .ZN(n430) );
  CLKBUF_X3 U1000 ( .A(b[13]), .Z(n840) );
  BUF_X2 U1001 ( .A(n867), .Z(n17) );
  XOR2_X1 U1002 ( .A(n620), .B(n568), .Z(n501) );
  NOR2_X1 U1003 ( .A1(n431), .A2(n444), .ZN(n1060) );
  OAI21_X1 U1004 ( .B1(n227), .B2(n233), .A(n228), .ZN(n1061) );
  NOR2_X1 U1005 ( .A1(n431), .A2(n444), .ZN(n227) );
  BUF_X2 U1006 ( .A(n867), .Z(n18) );
  CLKBUF_X3 U1007 ( .A(b[7]), .Z(n846) );
  XNOR2_X1 U1008 ( .A(n170), .B(n1062), .ZN(product[23]) );
  AND2_X1 U1009 ( .A1(n1051), .A2(n169), .ZN(n1062) );
  XNOR2_X1 U1010 ( .A(n25), .B(n850), .ZN(n1064) );
  BUF_X4 U1011 ( .A(a[9]), .Z(n25) );
  BUF_X2 U1012 ( .A(b[5]), .Z(n848) );
  OR2_X1 U1013 ( .A1(n1010), .A2(n416), .ZN(n1065) );
  BUF_X2 U1014 ( .A(b[14]), .Z(n839) );
  NOR2_X1 U1015 ( .A1(n1010), .A2(n416), .ZN(n211) );
  NOR2_X1 U1016 ( .A1(n341), .A2(n344), .ZN(n137) );
  NOR2_X1 U1017 ( .A1(n700), .A2(n685), .ZN(n298) );
  NOR2_X1 U1018 ( .A1(n519), .A2(n524), .ZN(n274) );
  NOR2_X1 U1019 ( .A1(n539), .A2(n540), .ZN(n290) );
  AND2_X1 U1020 ( .A1(n1004), .A2(n301), .ZN(product[1]) );
  CLKBUF_X1 U1021 ( .A(n49), .Z(n1069) );
  BUF_X1 U1022 ( .A(n862), .Z(n48) );
  BUF_X1 U1023 ( .A(n871), .Z(n40) );
  BUF_X1 U1024 ( .A(n876), .Z(n10) );
  INV_X1 U1025 ( .A(n1018), .ZN(n234) );
  INV_X1 U1026 ( .A(n1061), .ZN(n224) );
  INV_X1 U1027 ( .A(n1063), .ZN(n223) );
  NOR2_X1 U1028 ( .A1(n195), .A2(n162), .ZN(n160) );
  NOR2_X1 U1029 ( .A1(n195), .A2(n190), .ZN(n184) );
  NOR2_X1 U1030 ( .A1(n195), .A2(n173), .ZN(n171) );
  NOR2_X1 U1031 ( .A1(n149), .A2(n96), .ZN(n94) );
  NOR2_X1 U1032 ( .A1(n149), .A2(n124), .ZN(n118) );
  NOR2_X1 U1033 ( .A1(n149), .A2(n109), .ZN(n107) );
  INV_X1 U1034 ( .A(n98), .ZN(n96) );
  INV_X1 U1035 ( .A(n177), .ZN(n175) );
  INV_X1 U1036 ( .A(n149), .ZN(n147) );
  INV_X1 U1037 ( .A(n196), .ZN(n194) );
  INV_X1 U1038 ( .A(n195), .ZN(n193) );
  NAND2_X1 U1039 ( .A1(n317), .A2(n233), .ZN(n69) );
  INV_X1 U1040 ( .A(n232), .ZN(n317) );
  XNOR2_X1 U1041 ( .A(n240), .B(n70), .ZN(product[14]) );
  NAND2_X1 U1042 ( .A1(n1037), .A2(n239), .ZN(n70) );
  NAND2_X1 U1043 ( .A1(n1065), .A2(n212), .ZN(n66) );
  NOR2_X1 U1044 ( .A1(n223), .A2(n216), .ZN(n214) );
  NAND2_X1 U1045 ( .A1(n313), .A2(n205), .ZN(n65) );
  INV_X1 U1046 ( .A(n204), .ZN(n313) );
  XOR2_X1 U1047 ( .A(n229), .B(n68), .Z(product[16]) );
  NAND2_X1 U1048 ( .A1(n316), .A2(n228), .ZN(n68) );
  INV_X1 U1049 ( .A(n227), .ZN(n316) );
  OAI21_X1 U1050 ( .B1(n227), .B2(n233), .A(n228), .ZN(n226) );
  NOR2_X1 U1051 ( .A1(n232), .A2(n1060), .ZN(n225) );
  AOI21_X1 U1052 ( .B1(n255), .B2(n236), .A(n237), .ZN(n235) );
  XOR2_X1 U1053 ( .A(n220), .B(n67), .Z(product[17]) );
  NAND2_X1 U1054 ( .A1(n217), .A2(n1009), .ZN(n67) );
  NOR2_X1 U1055 ( .A1(n124), .A2(n100), .ZN(n98) );
  NOR2_X1 U1056 ( .A1(n177), .A2(n166), .ZN(n164) );
  INV_X1 U1057 ( .A(n197), .ZN(n195) );
  INV_X1 U1058 ( .A(n198), .ZN(n196) );
  OAI21_X1 U1059 ( .B1(n150), .B2(n124), .A(n125), .ZN(n119) );
  NAND2_X1 U1060 ( .A1(n164), .A2(n188), .ZN(n162) );
  OAI21_X1 U1061 ( .B1(n196), .B2(n190), .A(n191), .ZN(n185) );
  OAI21_X1 U1062 ( .B1(n196), .B2(n173), .A(n174), .ZN(n172) );
  AOI21_X1 U1063 ( .B1(n189), .B2(n175), .A(n180), .ZN(n174) );
  NAND2_X1 U1064 ( .A1(n188), .A2(n175), .ZN(n173) );
  NAND2_X1 U1065 ( .A1(n122), .A2(n999), .ZN(n109) );
  OAI21_X1 U1066 ( .B1(n224), .B2(n216), .A(n1009), .ZN(n215) );
  INV_X1 U1067 ( .A(n255), .ZN(n254) );
  INV_X1 U1068 ( .A(n124), .ZN(n122) );
  INV_X1 U1069 ( .A(n217), .ZN(n216) );
  INV_X1 U1070 ( .A(n218), .ZN(n217) );
  INV_X1 U1071 ( .A(n1017), .ZN(n177) );
  NOR2_X1 U1072 ( .A1(n149), .A2(n144), .ZN(n140) );
  NOR2_X1 U1073 ( .A1(n149), .A2(n133), .ZN(n131) );
  INV_X1 U1074 ( .A(n180), .ZN(n178) );
  NAND2_X1 U1075 ( .A1(n1066), .A2(n1011), .ZN(n241) );
  INV_X1 U1076 ( .A(n957), .ZN(n148) );
  INV_X1 U1077 ( .A(n1011), .ZN(n248) );
  INV_X1 U1078 ( .A(n233), .ZN(n231) );
  INV_X1 U1079 ( .A(n205), .ZN(n203) );
  INV_X1 U1080 ( .A(n1058), .ZN(n249) );
  NAND2_X1 U1081 ( .A1(n1011), .A2(n249), .ZN(n72) );
  NAND2_X1 U1082 ( .A1(n1000), .A2(n272), .ZN(n75) );
  NAND2_X1 U1083 ( .A1(n258), .A2(n1012), .ZN(n256) );
  AOI21_X1 U1084 ( .B1(n258), .B2(n264), .A(n259), .ZN(n257) );
  XNOR2_X1 U1085 ( .A(n267), .B(n74), .ZN(product[10]) );
  NAND2_X1 U1086 ( .A1(n1012), .A2(n266), .ZN(n74) );
  INV_X1 U1087 ( .A(n157), .ZN(n308) );
  INV_X1 U1088 ( .A(n272), .ZN(n270) );
  XOR2_X1 U1089 ( .A(n262), .B(n73), .Z(product[11]) );
  NAND2_X1 U1090 ( .A1(n321), .A2(n261), .ZN(n73) );
  AOI21_X1 U1091 ( .B1(n267), .B2(n1012), .A(n264), .ZN(n262) );
  INV_X1 U1092 ( .A(n199), .ZN(n312) );
  NOR2_X1 U1093 ( .A1(n458), .A2(n445), .ZN(n232) );
  XNOR2_X1 U1094 ( .A(n247), .B(n71), .ZN(product[13]) );
  NAND2_X1 U1095 ( .A1(n1066), .A2(n246), .ZN(n71) );
  NOR2_X1 U1096 ( .A1(n393), .A2(n404), .ZN(n204) );
  INV_X1 U1097 ( .A(n136), .ZN(n134) );
  NOR2_X1 U1098 ( .A1(n459), .A2(n470), .ZN(n238) );
  NAND2_X1 U1099 ( .A1(n135), .A2(n996), .ZN(n124) );
  AOI21_X1 U1100 ( .B1(n1066), .B2(n1058), .A(n1059), .ZN(n242) );
  OAI21_X1 U1101 ( .B1(n196), .B2(n162), .A(n163), .ZN(n161) );
  AOI21_X1 U1102 ( .B1(n164), .B2(n189), .A(n165), .ZN(n163) );
  OAI21_X1 U1103 ( .B1(n178), .B2(n166), .A(n169), .ZN(n165) );
  NAND2_X1 U1104 ( .A1(n445), .A2(n458), .ZN(n233) );
  NOR2_X1 U1105 ( .A1(n190), .A2(n153), .ZN(n151) );
  NAND2_X1 U1106 ( .A1(n393), .A2(n404), .ZN(n205) );
  OAI21_X1 U1107 ( .B1(n957), .B2(n96), .A(n97), .ZN(n95) );
  INV_X1 U1108 ( .A(n99), .ZN(n97) );
  OAI21_X1 U1109 ( .B1(n957), .B2(n109), .A(n110), .ZN(n108) );
  AOI21_X1 U1110 ( .B1(n123), .B2(n999), .A(n114), .ZN(n110) );
  NAND2_X1 U1111 ( .A1(n417), .A2(n430), .ZN(n219) );
  INV_X1 U1112 ( .A(n135), .ZN(n133) );
  INV_X1 U1113 ( .A(n190), .ZN(n188) );
  INV_X1 U1114 ( .A(n191), .ZN(n189) );
  NAND2_X1 U1115 ( .A1(n98), .A2(n997), .ZN(n87) );
  NAND2_X1 U1116 ( .A1(n999), .A2(n995), .ZN(n100) );
  NAND2_X1 U1117 ( .A1(n459), .A2(n470), .ZN(n239) );
  NAND2_X1 U1118 ( .A1(n405), .A2(n416), .ZN(n212) );
  INV_X1 U1119 ( .A(n182), .ZN(n180) );
  NOR2_X1 U1120 ( .A1(n149), .A2(n87), .ZN(n85) );
  OAI21_X1 U1121 ( .B1(n957), .B2(n87), .A(n88), .ZN(n86) );
  INV_X1 U1122 ( .A(n266), .ZN(n264) );
  INV_X1 U1123 ( .A(n125), .ZN(n123) );
  INV_X1 U1124 ( .A(n1051), .ZN(n166) );
  INV_X1 U1125 ( .A(n144), .ZN(n143) );
  INV_X1 U1126 ( .A(n261), .ZN(n259) );
  NAND2_X1 U1127 ( .A1(n326), .A2(n283), .ZN(n78) );
  NAND2_X1 U1128 ( .A1(n324), .A2(n275), .ZN(n76) );
  INV_X1 U1129 ( .A(n274), .ZN(n324) );
  NAND2_X1 U1130 ( .A1(n1001), .A2(n280), .ZN(n77) );
  XOR2_X1 U1131 ( .A(n93), .B(n54), .Z(product[30]) );
  NAND2_X1 U1132 ( .A1(n997), .A2(n92), .ZN(n54) );
  XOR2_X1 U1133 ( .A(n106), .B(n55), .Z(product[29]) );
  NAND2_X1 U1134 ( .A1(n995), .A2(n105), .ZN(n55) );
  INV_X1 U1135 ( .A(n280), .ZN(n278) );
  INV_X1 U1136 ( .A(n137), .ZN(n306) );
  AOI21_X1 U1137 ( .B1(n136), .B2(n996), .A(n127), .ZN(n125) );
  INV_X1 U1138 ( .A(n129), .ZN(n127) );
  XOR2_X1 U1139 ( .A(n117), .B(n56), .Z(product[28]) );
  NAND2_X1 U1140 ( .A1(n999), .A2(n116), .ZN(n56) );
  OAI21_X1 U1141 ( .B1(n125), .B2(n100), .A(n101), .ZN(n99) );
  AOI21_X1 U1142 ( .B1(n114), .B2(n995), .A(n103), .ZN(n101) );
  INV_X1 U1143 ( .A(n105), .ZN(n103) );
  OAI21_X1 U1144 ( .B1(n145), .B2(n137), .A(n138), .ZN(n136) );
  NOR2_X1 U1145 ( .A1(n357), .A2(n364), .ZN(n168) );
  NOR2_X1 U1146 ( .A1(n345), .A2(n350), .ZN(n144) );
  NOR2_X1 U1147 ( .A1(n383), .A2(n392), .ZN(n199) );
  NOR2_X1 U1148 ( .A1(n351), .A2(n356), .ZN(n157) );
  AOI21_X1 U1149 ( .B1(n99), .B2(n997), .A(n90), .ZN(n88) );
  INV_X1 U1150 ( .A(n92), .ZN(n90) );
  NAND2_X1 U1151 ( .A1(n345), .A2(n350), .ZN(n145) );
  NAND2_X1 U1152 ( .A1(n373), .A2(n382), .ZN(n191) );
  NAND2_X1 U1153 ( .A1(n357), .A2(n364), .ZN(n169) );
  NAND2_X1 U1154 ( .A1(n503), .A2(n510), .ZN(n266) );
  NAND2_X1 U1155 ( .A1(n493), .A2(n502), .ZN(n261) );
  NAND2_X1 U1156 ( .A1(n511), .A2(n518), .ZN(n272) );
  NAND2_X1 U1157 ( .A1(n383), .A2(n392), .ZN(n200) );
  NAND2_X1 U1158 ( .A1(n351), .A2(n356), .ZN(n158) );
  INV_X1 U1159 ( .A(n116), .ZN(n114) );
  XOR2_X1 U1160 ( .A(n82), .B(n301), .Z(product[2]) );
  NAND2_X1 U1161 ( .A1(n330), .A2(n299), .ZN(n82) );
  INV_X1 U1162 ( .A(n298), .ZN(n330) );
  XNOR2_X1 U1163 ( .A(n81), .B(n297), .ZN(product[3]) );
  NAND2_X1 U1164 ( .A1(n998), .A2(n296), .ZN(n81) );
  OAI21_X1 U1165 ( .B1(n298), .B2(n301), .A(n299), .ZN(n297) );
  OAI21_X1 U1166 ( .B1(n292), .B2(n290), .A(n291), .ZN(n289) );
  NAND2_X1 U1167 ( .A1(n574), .A2(n332), .ZN(n92) );
  AOI21_X1 U1168 ( .B1(n998), .B2(n297), .A(n294), .ZN(n292) );
  INV_X1 U1169 ( .A(n296), .ZN(n294) );
  NAND2_X1 U1170 ( .A1(n525), .A2(n530), .ZN(n280) );
  XNOR2_X1 U1171 ( .A(n643), .B(n601), .ZN(n443) );
  INV_X1 U1172 ( .A(n332), .ZN(n333) );
  NAND2_X1 U1173 ( .A1(n700), .A2(n685), .ZN(n299) );
  INV_X1 U1174 ( .A(n362), .ZN(n363) );
  INV_X1 U1175 ( .A(n428), .ZN(n429) );
  NAND2_X1 U1176 ( .A1(n337), .A2(n340), .ZN(n129) );
  NAND2_X1 U1177 ( .A1(n341), .A2(n344), .ZN(n138) );
  NAND2_X1 U1178 ( .A1(n336), .A2(n335), .ZN(n116) );
  NAND2_X1 U1179 ( .A1(n334), .A2(n333), .ZN(n105) );
  NAND2_X1 U1180 ( .A1(n519), .A2(n524), .ZN(n275) );
  NAND2_X1 U1181 ( .A1(n328), .A2(n291), .ZN(n80) );
  INV_X1 U1182 ( .A(n290), .ZN(n328) );
  OAI22_X1 U1183 ( .A1(n41), .A2(n720), .B1(n40), .B2(n719), .ZN(n338) );
  OAI22_X1 U1184 ( .A1(n5), .A2(n835), .B1(n834), .B2(n3), .ZN(n700) );
  OAI22_X1 U1185 ( .A1(n1021), .A2(n805), .B1(n10), .B2(n804), .ZN(n428) );
  OAI22_X1 U1186 ( .A1(n788), .A2(n17), .B1(n16), .B2(n787), .ZN(n402) );
  OAI22_X1 U1187 ( .A1(n29), .A2(n754), .B1(n1022), .B2(n753), .ZN(n362) );
  OAI22_X1 U1188 ( .A1(n1023), .A2(n737), .B1(n34), .B2(n736), .ZN(n348) );
  OAI22_X1 U1189 ( .A1(n41), .A2(n731), .B1(n39), .B2(n730), .ZN(n601) );
  OAI22_X1 U1190 ( .A1(n23), .A2(n776), .B1(n22), .B2(n775), .ZN(n643) );
  OAI22_X1 U1191 ( .A1(n48), .A2(n704), .B1(n46), .B2(n703), .ZN(n575) );
  INV_X1 U1192 ( .A(n545), .ZN(n590) );
  AOI21_X1 U1193 ( .B1(n41), .B2(n40), .A(n719), .ZN(n545) );
  OAI22_X1 U1194 ( .A1(n48), .A2(n706), .B1(n46), .B2(n705), .ZN(n577) );
  OAI22_X1 U1195 ( .A1(n11), .A2(n818), .B1(n9), .B2(n817), .ZN(n683) );
  OAI22_X1 U1196 ( .A1(n1049), .A2(n833), .B1(n832), .B2(n3), .ZN(n698) );
  AND2_X1 U1197 ( .A1(n1029), .A2(n558), .ZN(n669) );
  OAI22_X1 U1198 ( .A1(n48), .A2(n878), .B1(n718), .B2(n45), .ZN(n566) );
  OAI22_X1 U1199 ( .A1(n47), .A2(n717), .B1(n45), .B2(n716), .ZN(n588) );
  OR2_X1 U1200 ( .A1(n1069), .A2(n878), .ZN(n718) );
  OAI22_X1 U1201 ( .A1(n1023), .A2(n739), .B1(n34), .B2(n738), .ZN(n608) );
  OAI22_X1 U1202 ( .A1(n41), .A2(n724), .B1(n40), .B2(n723), .ZN(n594) );
  OAI22_X1 U1203 ( .A1(n48), .A2(n709), .B1(n46), .B2(n708), .ZN(n580) );
  OAI22_X1 U1204 ( .A1(n758), .A2(n30), .B1(n28), .B2(n757), .ZN(n626) );
  OAI22_X1 U1205 ( .A1(n773), .A2(n24), .B1(n22), .B2(n772), .ZN(n640) );
  OAI22_X1 U1206 ( .A1(n35), .A2(n743), .B1(n33), .B2(n742), .ZN(n612) );
  OAI22_X1 U1207 ( .A1(n1023), .A2(n749), .B1(n34), .B2(n748), .ZN(n618) );
  OAI22_X1 U1208 ( .A1(n29), .A2(n764), .B1(n1022), .B2(n763), .ZN(n632) );
  OAI22_X1 U1209 ( .A1(n18), .A2(n794), .B1(n1025), .B2(n793), .ZN(n660) );
  AOI21_X1 U1210 ( .B1(n1033), .B2(n28), .A(n753), .ZN(n551) );
  AOI21_X1 U1211 ( .B1(n1048), .B2(n4), .A(n821), .ZN(n563) );
  AOI21_X1 U1212 ( .B1(n24), .B2(n22), .A(n770), .ZN(n554) );
  OAI22_X1 U1213 ( .A1(n17), .A2(n802), .B1(n1025), .B2(n801), .ZN(n668) );
  OAI22_X1 U1214 ( .A1(n1006), .A2(n817), .B1(n9), .B2(n816), .ZN(n682) );
  OAI22_X1 U1215 ( .A1(n1049), .A2(n832), .B1(n831), .B2(n3), .ZN(n697) );
  NAND2_X1 U1216 ( .A1(n701), .A2(n573), .ZN(n301) );
  AND2_X1 U1217 ( .A1(n1029), .A2(n561), .ZN(n685) );
  INV_X1 U1218 ( .A(n9), .ZN(n561) );
  OAI22_X1 U1219 ( .A1(n47), .A2(n712), .B1(n46), .B2(n711), .ZN(n583) );
  INV_X1 U1220 ( .A(n557), .ZN(n654) );
  AOI21_X1 U1221 ( .B1(n18), .B2(n16), .A(n787), .ZN(n557) );
  OAI22_X1 U1222 ( .A1(n1023), .A2(n744), .B1(n34), .B2(n743), .ZN(n613) );
  OAI22_X1 U1223 ( .A1(n1033), .A2(n759), .B1(n28), .B2(n758), .ZN(n627) );
  OAI22_X1 U1224 ( .A1(n23), .A2(n774), .B1(n22), .B2(n773), .ZN(n641) );
  OAI22_X1 U1225 ( .A1(n18), .A2(n789), .B1(n788), .B2(n1024), .ZN(n655) );
  OAI22_X1 U1226 ( .A1(n42), .A2(n729), .B1(n39), .B2(n728), .ZN(n599) );
  OAI22_X1 U1227 ( .A1(n47), .A2(n711), .B1(n46), .B2(n710), .ZN(n582) );
  OAI22_X1 U1228 ( .A1(n1034), .A2(n756), .B1(n1022), .B2(n755), .ZN(n624) );
  OAI22_X1 U1229 ( .A1(n41), .A2(n726), .B1(n40), .B2(n725), .ZN(n596) );
  OAI22_X1 U1230 ( .A1(n1023), .A2(n740), .B1(n34), .B2(n739), .ZN(n609) );
  OAI22_X1 U1231 ( .A1(n41), .A2(n725), .B1(n40), .B2(n724), .ZN(n595) );
  OAI22_X1 U1232 ( .A1(n1020), .A2(n809), .B1(n10), .B2(n808), .ZN(n674) );
  OAI22_X1 U1233 ( .A1(n23), .A2(n779), .B1(n21), .B2(n778), .ZN(n646) );
  OAI22_X1 U1234 ( .A1(n6), .A2(n824), .B1(n823), .B2(n4), .ZN(n689) );
  OAI22_X1 U1235 ( .A1(n1023), .A2(n750), .B1(n33), .B2(n749), .ZN(n619) );
  OAI22_X1 U1236 ( .A1(n24), .A2(n780), .B1(n21), .B2(n779), .ZN(n647) );
  OAI22_X1 U1237 ( .A1(n1020), .A2(n810), .B1(n10), .B2(n809), .ZN(n675) );
  OAI22_X1 U1238 ( .A1(n42), .A2(n730), .B1(n39), .B2(n729), .ZN(n600) );
  OAI22_X1 U1239 ( .A1(n1023), .A2(n741), .B1(n34), .B2(n740), .ZN(n610) );
  OAI22_X1 U1240 ( .A1(n1023), .A2(n742), .B1(n34), .B2(n741), .ZN(n611) );
  OAI22_X1 U1241 ( .A1(n24), .A2(n772), .B1(n22), .B2(n771), .ZN(n639) );
  OAI22_X1 U1242 ( .A1(n41), .A2(n727), .B1(n39), .B2(n726), .ZN(n597) );
  OAI22_X1 U1243 ( .A1(n18), .A2(n801), .B1(n1024), .B2(n800), .ZN(n667) );
  OAI22_X1 U1244 ( .A1(n5), .A2(n828), .B1(n827), .B2(n4), .ZN(n693) );
  OAI22_X1 U1245 ( .A1(n18), .A2(n797), .B1(n1024), .B2(n796), .ZN(n663) );
  OAI22_X1 U1246 ( .A1(n29), .A2(n767), .B1(n1022), .B2(n1027), .ZN(n635) );
  OAI22_X1 U1247 ( .A1(n11), .A2(n812), .B1(n9), .B2(n811), .ZN(n677) );
  OAI22_X1 U1248 ( .A1(n1020), .A2(n813), .B1(n9), .B2(n812), .ZN(n678) );
  OAI22_X1 U1249 ( .A1(n24), .A2(n783), .B1(n21), .B2(n782), .ZN(n650) );
  OAI22_X1 U1250 ( .A1(n18), .A2(n798), .B1(n1024), .B2(n797), .ZN(n664) );
  OAI22_X1 U1251 ( .A1(n1021), .A2(n816), .B1(n9), .B2(n815), .ZN(n681) );
  OAI22_X1 U1252 ( .A1(n1048), .A2(n831), .B1(n830), .B2(n3), .ZN(n696) );
  AND2_X1 U1253 ( .A1(n1069), .A2(n555), .ZN(n653) );
  OAI22_X1 U1254 ( .A1(n24), .A2(n778), .B1(n21), .B2(n777), .ZN(n645) );
  OAI22_X1 U1255 ( .A1(n18), .A2(n793), .B1(n16), .B2(n792), .ZN(n659) );
  OAI22_X1 U1256 ( .A1(n23), .A2(n784), .B1(n21), .B2(n783), .ZN(n651) );
  OAI22_X1 U1257 ( .A1(n1006), .A2(n814), .B1(n9), .B2(n813), .ZN(n679) );
  OAI22_X1 U1258 ( .A1(n18), .A2(n792), .B1(n16), .B2(n791), .ZN(n658) );
  OAI22_X1 U1259 ( .A1(n5), .A2(n822), .B1(n821), .B2(n4), .ZN(n687) );
  OAI22_X1 U1260 ( .A1(n1034), .A2(n762), .B1(n1022), .B2(n761), .ZN(n630) );
  OAI22_X1 U1261 ( .A1(n1021), .A2(n807), .B1(n10), .B2(n806), .ZN(n672) );
  OAI22_X1 U1262 ( .A1(n6), .A2(n827), .B1(n826), .B2(n4), .ZN(n692) );
  AND2_X1 U1263 ( .A1(n1029), .A2(n549), .ZN(n621) );
  OAI22_X1 U1264 ( .A1(n6), .A2(n830), .B1(n829), .B2(n3), .ZN(n695) );
  OAI22_X1 U1265 ( .A1(n18), .A2(n800), .B1(n1025), .B2(n799), .ZN(n666) );
  OAI22_X1 U1266 ( .A1(n1021), .A2(n815), .B1(n9), .B2(n814), .ZN(n680) );
  OAI22_X1 U1267 ( .A1(n1034), .A2(n763), .B1(n1022), .B2(n762), .ZN(n631) );
  OAI22_X1 U1268 ( .A1(n41), .A2(n733), .B1(n39), .B2(n732), .ZN(n603) );
  OAI22_X1 U1269 ( .A1(n1021), .A2(n808), .B1(n10), .B2(n807), .ZN(n673) );
  OAI22_X1 U1270 ( .A1(n35), .A2(n746), .B1(n34), .B2(n745), .ZN(n615) );
  OAI22_X1 U1271 ( .A1(n17), .A2(n791), .B1(n790), .B2(n1024), .ZN(n657) );
  OAI22_X1 U1272 ( .A1(n11), .A2(n806), .B1(n10), .B2(n805), .ZN(n671) );
  OAI22_X1 U1273 ( .A1(n47), .A2(n714), .B1(n45), .B2(n713), .ZN(n585) );
  INV_X1 U1274 ( .A(n560), .ZN(n670) );
  AOI21_X1 U1275 ( .B1(n12), .B2(n10), .A(n804), .ZN(n560) );
  OAI22_X1 U1276 ( .A1(n48), .A2(n708), .B1(n46), .B2(n707), .ZN(n579) );
  OAI22_X1 U1277 ( .A1(n41), .A2(n723), .B1(n40), .B2(n722), .ZN(n593) );
  INV_X1 U1278 ( .A(n551), .ZN(n622) );
  OAI22_X1 U1279 ( .A1(n48), .A2(n705), .B1(n46), .B2(n704), .ZN(n576) );
  INV_X1 U1280 ( .A(n338), .ZN(n339) );
  OAI22_X1 U1281 ( .A1(n1034), .A2(n757), .B1(n1022), .B2(n756), .ZN(n625) );
  OAI22_X1 U1282 ( .A1(n18), .A2(n795), .B1(n16), .B2(n794), .ZN(n661) );
  OAI22_X1 U1283 ( .A1(n1023), .A2(n738), .B1(n34), .B2(n737), .ZN(n607) );
  OAI22_X1 U1284 ( .A1(n24), .A2(n781), .B1(n21), .B2(n780), .ZN(n648) );
  OAI22_X1 U1285 ( .A1(n1020), .A2(n811), .B1(n10), .B2(n810), .ZN(n676) );
  OAI22_X1 U1286 ( .A1(n1023), .A2(n747), .B1(n34), .B2(n746), .ZN(n616) );
  OAI22_X1 U1287 ( .A1(n42), .A2(n732), .B1(n39), .B2(n731), .ZN(n602) );
  OAI22_X1 U1288 ( .A1(n23), .A2(n777), .B1(n22), .B2(n776), .ZN(n644) );
  OAI22_X1 U1289 ( .A1(n1048), .A2(n826), .B1(n825), .B2(n4), .ZN(n691) );
  OAI22_X1 U1290 ( .A1(n796), .A2(n17), .B1(n795), .B2(n1024), .ZN(n662) );
  OAI22_X1 U1291 ( .A1(n47), .A2(n716), .B1(n45), .B2(n715), .ZN(n587) );
  OAI22_X1 U1292 ( .A1(n1034), .A2(n761), .B1(n28), .B2(n760), .ZN(n629) );
  INV_X1 U1293 ( .A(n563), .ZN(n686) );
  OAI22_X1 U1294 ( .A1(n6), .A2(n829), .B1(n828), .B2(n3), .ZN(n694) );
  OAI22_X1 U1295 ( .A1(n18), .A2(n799), .B1(n1025), .B2(n798), .ZN(n665) );
  AND2_X1 U1296 ( .A1(n1069), .A2(n552), .ZN(n637) );
  OAI22_X1 U1297 ( .A1(n5), .A2(n823), .B1(n822), .B2(n4), .ZN(n688) );
  OAI22_X1 U1298 ( .A1(n35), .A2(n748), .B1(n747), .B2(n33), .ZN(n617) );
  AND2_X1 U1299 ( .A1(n1029), .A2(n543), .ZN(n589) );
  OAI22_X1 U1300 ( .A1(n47), .A2(n715), .B1(n45), .B2(n714), .ZN(n586) );
  OAI22_X1 U1301 ( .A1(n35), .A2(n745), .B1(n33), .B2(n744), .ZN(n614) );
  OAI22_X1 U1302 ( .A1(n17), .A2(n790), .B1(n16), .B2(n789), .ZN(n656) );
  NAND2_X1 U1303 ( .A1(n539), .A2(n540), .ZN(n291) );
  OAI22_X1 U1304 ( .A1(n42), .A2(n879), .B1(n735), .B2(n40), .ZN(n567) );
  OAI22_X1 U1305 ( .A1(n734), .A2(n42), .B1(n39), .B2(n733), .ZN(n604) );
  OR2_X1 U1306 ( .A1(n1068), .A2(n879), .ZN(n735) );
  INV_X1 U1307 ( .A(n542), .ZN(n574) );
  AOI21_X1 U1308 ( .B1(n48), .B2(n46), .A(n702), .ZN(n542) );
  OAI22_X1 U1309 ( .A1(n41), .A2(n728), .B1(n39), .B2(n727), .ZN(n598) );
  OAI22_X1 U1310 ( .A1(n47), .A2(n713), .B1(n46), .B2(n712), .ZN(n584) );
  INV_X1 U1311 ( .A(n402), .ZN(n403) );
  OAI22_X1 U1312 ( .A1(n48), .A2(n707), .B1(n46), .B2(n706), .ZN(n578) );
  OAI22_X1 U1313 ( .A1(n41), .A2(n722), .B1(n40), .B2(n721), .ZN(n592) );
  INV_X1 U1314 ( .A(n348), .ZN(n349) );
  AND2_X1 U1315 ( .A1(n1069), .A2(a[0]), .ZN(product[0]) );
  OAI22_X1 U1316 ( .A1(n1049), .A2(n825), .B1(n824), .B2(n4), .ZN(n690) );
  OAI22_X1 U1317 ( .A1(n1033), .A2(n1064), .B1(n28), .B2(n764), .ZN(n633) );
  AND2_X1 U1318 ( .A1(n1069), .A2(n546), .ZN(n605) );
  OR2_X1 U1319 ( .A1(n1068), .A2(n880), .ZN(n752) );
  OR2_X1 U1320 ( .A1(n1029), .A2(n882), .ZN(n786) );
  OR2_X1 U1321 ( .A1(n1029), .A2(n881), .ZN(n769) );
  OAI22_X1 U1322 ( .A1(n41), .A2(n721), .B1(n40), .B2(n720), .ZN(n591) );
  INV_X1 U1323 ( .A(n548), .ZN(n606) );
  AOI21_X1 U1324 ( .B1(n35), .B2(n34), .A(n736), .ZN(n548) );
  OAI22_X1 U1325 ( .A1(n1033), .A2(n755), .B1(n1022), .B2(n754), .ZN(n623) );
  OAI22_X1 U1326 ( .A1(n47), .A2(n710), .B1(n46), .B2(n709), .ZN(n581) );
  INV_X1 U1327 ( .A(n554), .ZN(n638) );
  INV_X1 U1328 ( .A(n39), .ZN(n546) );
  INV_X1 U1329 ( .A(n16), .ZN(n558) );
  INV_X1 U1330 ( .A(n33), .ZN(n549) );
  INV_X1 U1331 ( .A(n45), .ZN(n543) );
  INV_X1 U1332 ( .A(n1022), .ZN(n552) );
  INV_X1 U1333 ( .A(n21), .ZN(n555) );
  BUF_X1 U1334 ( .A(n877), .Z(n3) );
  OAI22_X1 U1335 ( .A1(n6), .A2(n834), .B1(n833), .B2(n3), .ZN(n699) );
  OAI22_X1 U1336 ( .A1(n11), .A2(n819), .B1(n9), .B2(n818), .ZN(n684) );
  BUF_X1 U1337 ( .A(n865), .Z(n30) );
  BUF_X1 U1338 ( .A(n874), .Z(n22) );
  OAI22_X1 U1339 ( .A1(n1049), .A2(n836), .B1(n835), .B2(n3), .ZN(n701) );
  OAI22_X1 U1340 ( .A1(n29), .A2(n768), .B1(n1022), .B2(n767), .ZN(n636) );
  OAI22_X1 U1341 ( .A1(n1033), .A2(n881), .B1(n769), .B2(n1022), .ZN(n569) );
  BUF_X1 U1342 ( .A(n870), .Z(n46) );
  XNOR2_X1 U1343 ( .A(n1019), .B(n839), .ZN(n788) );
  XNOR2_X1 U1344 ( .A(n847), .B(n13), .ZN(n796) );
  XNOR2_X1 U1345 ( .A(n1019), .B(n840), .ZN(n789) );
  XNOR2_X1 U1346 ( .A(n13), .B(n846), .ZN(n795) );
  XNOR2_X1 U1347 ( .A(n1019), .B(n844), .ZN(n793) );
  XNOR2_X1 U1348 ( .A(n1019), .B(n845), .ZN(n794) );
  XNOR2_X1 U1349 ( .A(n1019), .B(n841), .ZN(n790) );
  XNOR2_X1 U1350 ( .A(n1019), .B(n852), .ZN(n801) );
  XNOR2_X1 U1351 ( .A(n1019), .B(n848), .ZN(n797) );
  XNOR2_X1 U1352 ( .A(n1019), .B(n849), .ZN(n798) );
  XNOR2_X1 U1353 ( .A(n1019), .B(n843), .ZN(n792) );
  XNOR2_X1 U1354 ( .A(n1019), .B(n842), .ZN(n791) );
  XNOR2_X1 U1355 ( .A(n1019), .B(n851), .ZN(n800) );
  XNOR2_X1 U1356 ( .A(n1019), .B(n850), .ZN(n799) );
  OAI22_X1 U1357 ( .A1(n1023), .A2(n751), .B1(n33), .B2(n750), .ZN(n620) );
  OAI22_X1 U1358 ( .A1(n35), .A2(n880), .B1(n752), .B2(n33), .ZN(n568) );
  BUF_X1 U1359 ( .A(n870), .Z(n45) );
  BUF_X1 U1360 ( .A(n874), .Z(n21) );
  BUF_X1 U1361 ( .A(n877), .Z(n4) );
  BUF_X1 U1362 ( .A(n872), .Z(n34) );
  BUF_X1 U1363 ( .A(n869), .Z(n6) );
  BUF_X1 U1364 ( .A(n873), .Z(n28) );
  XNOR2_X1 U1365 ( .A(n1019), .B(n1068), .ZN(n802) );
  BUF_X1 U1366 ( .A(n869), .Z(n5) );
  OAI22_X1 U1367 ( .A1(n24), .A2(n785), .B1(n21), .B2(n784), .ZN(n652) );
  OAI22_X1 U1368 ( .A1(n23), .A2(n882), .B1(n786), .B2(n22), .ZN(n570) );
  OAI22_X1 U1369 ( .A1(n5), .A2(n885), .B1(n837), .B2(n4), .ZN(n573) );
  INV_X1 U1370 ( .A(n1028), .ZN(n885) );
  OAI22_X1 U1371 ( .A1(n1020), .A2(n884), .B1(n820), .B2(n10), .ZN(n572) );
  OR2_X1 U1372 ( .A1(n1029), .A2(n884), .ZN(n820) );
  INV_X1 U1373 ( .A(n7), .ZN(n884) );
  INV_X1 U1374 ( .A(n1032), .ZN(n882) );
  INV_X1 U1375 ( .A(n25), .ZN(n881) );
  INV_X1 U1376 ( .A(n37), .ZN(n879) );
  INV_X1 U1377 ( .A(n31), .ZN(n880) );
  INV_X1 U1378 ( .A(n43), .ZN(n878) );
  XNOR2_X1 U1379 ( .A(a[8]), .B(a[7]), .ZN(n873) );
  XNOR2_X1 U1380 ( .A(a[6]), .B(a[5]), .ZN(n874) );
  XNOR2_X1 U1381 ( .A(a[10]), .B(a[9]), .ZN(n872) );
  BUF_X2 U1382 ( .A(a[3]), .Z(n7) );
  XNOR2_X1 U1383 ( .A(a[14]), .B(a[13]), .ZN(n870) );
  NAND2_X1 U1384 ( .A1(n855), .A2(n871), .ZN(n863) );
  NAND2_X1 U1385 ( .A1(n860), .A2(n876), .ZN(n868) );
  NAND2_X1 U1386 ( .A1(n857), .A2(n873), .ZN(n865) );
  NAND2_X1 U1387 ( .A1(n858), .A2(n874), .ZN(n866) );
  INV_X1 U1388 ( .A(a[0]), .ZN(n877) );
  XNOR2_X1 U1389 ( .A(n13), .B(n838), .ZN(n787) );
  OAI22_X1 U1390 ( .A1(n24), .A2(n771), .B1(n22), .B2(n770), .ZN(n380) );
  INV_X1 U1391 ( .A(n380), .ZN(n381) );
  NAND2_X1 U1392 ( .A1(n531), .A2(n534), .ZN(n283) );
  NAND2_X1 U1393 ( .A1(n854), .A2(n870), .ZN(n862) );
  OAI22_X1 U1394 ( .A1(n766), .A2(n30), .B1(n765), .B2(n28), .ZN(n634) );
  NAND2_X1 U1395 ( .A1(n209), .A2(n225), .ZN(n207) );
  NAND2_X1 U1396 ( .A1(n856), .A2(n872), .ZN(n864) );
  OAI22_X1 U1397 ( .A1(n24), .A2(n782), .B1(n21), .B2(n781), .ZN(n649) );
  XNOR2_X1 U1398 ( .A(n25), .B(n1069), .ZN(n768) );
  XNOR2_X1 U1399 ( .A(n25), .B(n838), .ZN(n753) );
  XNOR2_X1 U1400 ( .A(n25), .B(n841), .ZN(n756) );
  XNOR2_X1 U1401 ( .A(n25), .B(n840), .ZN(n755) );
  XNOR2_X1 U1402 ( .A(n25), .B(n852), .ZN(n767) );
  XNOR2_X1 U1403 ( .A(n25), .B(n839), .ZN(n754) );
  XNOR2_X1 U1404 ( .A(n25), .B(n847), .ZN(n762) );
  XNOR2_X1 U1405 ( .A(n846), .B(n25), .ZN(n761) );
  XNOR2_X1 U1406 ( .A(n25), .B(n848), .ZN(n763) );
  XNOR2_X1 U1407 ( .A(n25), .B(n845), .ZN(n760) );
  XNOR2_X1 U1408 ( .A(n25), .B(n843), .ZN(n758) );
  XNOR2_X1 U1409 ( .A(n25), .B(n849), .ZN(n764) );
  XNOR2_X1 U1410 ( .A(n25), .B(n842), .ZN(n757) );
  XNOR2_X1 U1411 ( .A(n25), .B(n844), .ZN(n759) );
  XNOR2_X1 U1412 ( .A(n25), .B(n851), .ZN(n766) );
  XNOR2_X1 U1413 ( .A(n25), .B(n850), .ZN(n765) );
  INV_X1 U1414 ( .A(n282), .ZN(n326) );
  NOR2_X1 U1415 ( .A1(n531), .A2(n534), .ZN(n282) );
  OAI21_X1 U1416 ( .B1(n219), .B2(n1042), .A(n212), .ZN(n210) );
  OAI22_X1 U1417 ( .A1(n30), .A2(n760), .B1(n759), .B2(n1022), .ZN(n628) );
  XNOR2_X1 U1418 ( .A(n1031), .B(n1029), .ZN(n785) );
  XNOR2_X1 U1419 ( .A(n1031), .B(n851), .ZN(n783) );
  XNOR2_X1 U1420 ( .A(n1032), .B(n852), .ZN(n784) );
  XNOR2_X1 U1421 ( .A(n1032), .B(n845), .ZN(n777) );
  XNOR2_X1 U1422 ( .A(n1032), .B(n844), .ZN(n776) );
  XNOR2_X1 U1423 ( .A(n1031), .B(n848), .ZN(n780) );
  XNOR2_X1 U1424 ( .A(n1032), .B(n850), .ZN(n782) );
  XNOR2_X1 U1425 ( .A(n1032), .B(n849), .ZN(n781) );
  XNOR2_X1 U1426 ( .A(n1031), .B(n847), .ZN(n779) );
  XNOR2_X1 U1427 ( .A(n1031), .B(n846), .ZN(n778) );
  XNOR2_X1 U1428 ( .A(n1032), .B(n843), .ZN(n775) );
  XNOR2_X1 U1429 ( .A(n1030), .B(n841), .ZN(n773) );
  XNOR2_X1 U1430 ( .A(n1030), .B(n840), .ZN(n772) );
  XNOR2_X1 U1431 ( .A(n1030), .B(n842), .ZN(n774) );
  XNOR2_X1 U1432 ( .A(n1031), .B(n839), .ZN(n771) );
  XNOR2_X1 U1433 ( .A(n1031), .B(n838), .ZN(n770) );
  AOI21_X1 U1434 ( .B1(n1035), .B2(n226), .A(n210), .ZN(n208) );
  XNOR2_X1 U1435 ( .A(a[12]), .B(a[11]), .ZN(n871) );
  XNOR2_X1 U1436 ( .A(n79), .B(n289), .ZN(product[5]) );
  AOI21_X1 U1437 ( .B1(n1002), .B2(n289), .A(n286), .ZN(n284) );
  XNOR2_X1 U1438 ( .A(n7), .B(n847), .ZN(n813) );
  XNOR2_X1 U1439 ( .A(n7), .B(n846), .ZN(n812) );
  XNOR2_X1 U1440 ( .A(n7), .B(n845), .ZN(n811) );
  XNOR2_X1 U1441 ( .A(n7), .B(n850), .ZN(n816) );
  XNOR2_X1 U1442 ( .A(n7), .B(n849), .ZN(n815) );
  XNOR2_X1 U1443 ( .A(n7), .B(n848), .ZN(n814) );
  XNOR2_X1 U1444 ( .A(n7), .B(n844), .ZN(n810) );
  XNOR2_X1 U1445 ( .A(n7), .B(n851), .ZN(n817) );
  XNOR2_X1 U1446 ( .A(n7), .B(n841), .ZN(n807) );
  XNOR2_X1 U1447 ( .A(n7), .B(n842), .ZN(n808) );
  XNOR2_X1 U1448 ( .A(n7), .B(n843), .ZN(n809) );
  XNOR2_X1 U1449 ( .A(n7), .B(n840), .ZN(n806) );
  XNOR2_X1 U1450 ( .A(n7), .B(n839), .ZN(n805) );
  XNOR2_X1 U1451 ( .A(n7), .B(n1068), .ZN(n819) );
  XNOR2_X1 U1452 ( .A(n7), .B(n852), .ZN(n818) );
  XNOR2_X1 U1453 ( .A(n7), .B(n838), .ZN(n804) );
  XNOR2_X1 U1454 ( .A(a[4]), .B(a[3]), .ZN(n875) );
  XOR2_X1 U1455 ( .A(n80), .B(n292), .Z(product[4]) );
  NOR2_X1 U1456 ( .A1(n218), .A2(n211), .ZN(n209) );
  NOR2_X1 U1457 ( .A1(n417), .A2(n430), .ZN(n218) );
  NAND2_X1 U1458 ( .A1(n861), .A2(n877), .ZN(n869) );
  NAND2_X1 U1459 ( .A1(n431), .A2(n444), .ZN(n228) );
  XNOR2_X1 U1460 ( .A(n43), .B(n840), .ZN(n704) );
  XNOR2_X1 U1461 ( .A(n43), .B(n1036), .ZN(n705) );
  XNOR2_X1 U1462 ( .A(n43), .B(n839), .ZN(n703) );
  XNOR2_X1 U1463 ( .A(n43), .B(n838), .ZN(n702) );
  XNOR2_X1 U1464 ( .A(n43), .B(n1053), .ZN(n707) );
  XNOR2_X1 U1465 ( .A(n43), .B(n842), .ZN(n706) );
  XNOR2_X1 U1466 ( .A(n43), .B(n844), .ZN(n708) );
  XNOR2_X1 U1467 ( .A(n43), .B(n847), .ZN(n711) );
  XNOR2_X1 U1468 ( .A(n43), .B(n846), .ZN(n710) );
  XNOR2_X1 U1469 ( .A(n43), .B(n845), .ZN(n709) );
  XNOR2_X1 U1470 ( .A(n43), .B(n849), .ZN(n713) );
  XNOR2_X1 U1471 ( .A(n848), .B(n43), .ZN(n712) );
  XNOR2_X1 U1472 ( .A(n43), .B(n1029), .ZN(n717) );
  XNOR2_X1 U1473 ( .A(n43), .B(n851), .ZN(n715) );
  XNOR2_X1 U1474 ( .A(n43), .B(n852), .ZN(n716) );
  XNOR2_X1 U1475 ( .A(n43), .B(n850), .ZN(n714) );
  INV_X1 U1476 ( .A(n13), .ZN(n883) );
  OAI21_X1 U1477 ( .B1(n254), .B2(n248), .A(n249), .ZN(n247) );
  OAI21_X1 U1478 ( .B1(n254), .B2(n241), .A(n1046), .ZN(n240) );
  XOR2_X1 U1479 ( .A(n254), .B(n72), .Z(product[12]) );
  NAND2_X1 U1480 ( .A1(n859), .A2(n875), .ZN(n867) );
  OAI21_X1 U1481 ( .B1(n150), .B2(n144), .A(n145), .ZN(n141) );
  OAI21_X1 U1482 ( .B1(n150), .B2(n133), .A(n134), .ZN(n132) );
  AOI21_X1 U1483 ( .B1(n281), .B2(n1001), .A(n278), .ZN(n276) );
  OAI21_X1 U1484 ( .B1(n276), .B2(n274), .A(n275), .ZN(n273) );
  OAI22_X1 U1485 ( .A1(n17), .A2(n883), .B1(n803), .B2(n1025), .ZN(n571) );
  OR2_X1 U1486 ( .A1(n1068), .A2(n883), .ZN(n803) );
  XNOR2_X1 U1487 ( .A(n954), .B(n839), .ZN(n737) );
  XNOR2_X1 U1488 ( .A(n954), .B(n838), .ZN(n736) );
  XNOR2_X1 U1489 ( .A(n954), .B(n840), .ZN(n738) );
  XNOR2_X1 U1490 ( .A(n954), .B(n1053), .ZN(n741) );
  XNOR2_X1 U1491 ( .A(n31), .B(n842), .ZN(n740) );
  XNOR2_X1 U1492 ( .A(n31), .B(n841), .ZN(n739) );
  XNOR2_X1 U1493 ( .A(n31), .B(n1068), .ZN(n751) );
  XNOR2_X1 U1494 ( .A(n31), .B(n851), .ZN(n749) );
  XNOR2_X1 U1495 ( .A(n31), .B(n852), .ZN(n750) );
  XNOR2_X1 U1496 ( .A(n31), .B(n845), .ZN(n743) );
  XNOR2_X1 U1497 ( .A(n31), .B(n850), .ZN(n748) );
  XNOR2_X1 U1498 ( .A(n31), .B(n844), .ZN(n742) );
  XNOR2_X1 U1499 ( .A(n31), .B(n848), .ZN(n746) );
  XNOR2_X1 U1500 ( .A(n31), .B(n849), .ZN(n747) );
  XNOR2_X1 U1501 ( .A(n31), .B(n846), .ZN(n744) );
  XNOR2_X1 U1502 ( .A(n847), .B(n31), .ZN(n745) );
  OAI22_X1 U1503 ( .A1(n23), .A2(n775), .B1(n22), .B2(n774), .ZN(n642) );
  NAND2_X1 U1504 ( .A1(n365), .A2(n372), .ZN(n182) );
  INV_X1 U1505 ( .A(n288), .ZN(n286) );
  NAND2_X1 U1506 ( .A1(n1002), .A2(n288), .ZN(n79) );
  INV_X1 U1507 ( .A(n260), .ZN(n258) );
  INV_X1 U1508 ( .A(n260), .ZN(n321) );
  NOR2_X1 U1509 ( .A1(n493), .A2(n502), .ZN(n260) );
  NAND2_X1 U1510 ( .A1(n535), .A2(n538), .ZN(n288) );
  NOR2_X1 U1511 ( .A1(n204), .A2(n199), .ZN(n197) );
  OAI21_X1 U1512 ( .B1(n199), .B2(n205), .A(n200), .ZN(n198) );
  AOI21_X1 U1513 ( .B1(n214), .B2(n234), .A(n215), .ZN(n213) );
  XNOR2_X1 U1514 ( .A(n234), .B(n69), .ZN(product[15]) );
  AOI21_X1 U1515 ( .B1(n234), .B2(n317), .A(n231), .ZN(n229) );
  AOI21_X1 U1516 ( .B1(n234), .B2(n1063), .A(n1061), .ZN(n220) );
  XNOR2_X1 U1517 ( .A(n1028), .B(n845), .ZN(n828) );
  XNOR2_X1 U1518 ( .A(n1028), .B(n848), .ZN(n831) );
  XNOR2_X1 U1519 ( .A(n1028), .B(n846), .ZN(n829) );
  XNOR2_X1 U1520 ( .A(n1), .B(n847), .ZN(n830) );
  XNOR2_X1 U1521 ( .A(n1028), .B(n841), .ZN(n824) );
  XNOR2_X1 U1522 ( .A(n1028), .B(n849), .ZN(n832) );
  XNOR2_X1 U1523 ( .A(n1028), .B(n840), .ZN(n823) );
  XNOR2_X1 U1524 ( .A(n1028), .B(n844), .ZN(n827) );
  XNOR2_X1 U1525 ( .A(n1028), .B(n1029), .ZN(n836) );
  XNOR2_X1 U1526 ( .A(n1), .B(n842), .ZN(n825) );
  XNOR2_X1 U1527 ( .A(n1), .B(n843), .ZN(n826) );
  XNOR2_X1 U1528 ( .A(n1), .B(n839), .ZN(n822) );
  XNOR2_X1 U1529 ( .A(n1028), .B(n852), .ZN(n835) );
  XNOR2_X1 U1530 ( .A(n1028), .B(n851), .ZN(n834) );
  XNOR2_X1 U1531 ( .A(n1), .B(n850), .ZN(n833) );
  XNOR2_X1 U1532 ( .A(n1), .B(n838), .ZN(n821) );
  NOR2_X1 U1533 ( .A1(n144), .A2(n137), .ZN(n135) );
  NOR2_X1 U1534 ( .A1(n241), .A2(n956), .ZN(n236) );
  OAI21_X1 U1535 ( .B1(n242), .B2(n238), .A(n239), .ZN(n237) );
  XNOR2_X1 U1536 ( .A(n1043), .B(n1036), .ZN(n722) );
  XNOR2_X1 U1537 ( .A(n1043), .B(n840), .ZN(n721) );
  XNOR2_X1 U1538 ( .A(n1043), .B(n842), .ZN(n723) );
  XNOR2_X1 U1539 ( .A(n1043), .B(n845), .ZN(n726) );
  XNOR2_X1 U1540 ( .A(n1043), .B(n839), .ZN(n720) );
  XNOR2_X1 U1541 ( .A(n1043), .B(n844), .ZN(n725) );
  XNOR2_X1 U1542 ( .A(n1043), .B(n838), .ZN(n719) );
  XNOR2_X1 U1543 ( .A(n1043), .B(n843), .ZN(n724) );
  XNOR2_X1 U1544 ( .A(n1043), .B(n846), .ZN(n727) );
  XNOR2_X1 U1545 ( .A(n1043), .B(n851), .ZN(n732) );
  XNOR2_X1 U1546 ( .A(n1043), .B(n850), .ZN(n731) );
  XNOR2_X1 U1547 ( .A(n37), .B(n849), .ZN(n730) );
  XNOR2_X1 U1548 ( .A(n37), .B(n847), .ZN(n728) );
  XNOR2_X1 U1549 ( .A(n848), .B(n37), .ZN(n729) );
  XNOR2_X1 U1550 ( .A(n1043), .B(n1029), .ZN(n734) );
  XNOR2_X1 U1551 ( .A(n37), .B(n852), .ZN(n733) );
  XOR2_X1 U1552 ( .A(n213), .B(n66), .Z(product[18]) );
  NAND2_X1 U1553 ( .A1(n197), .A2(n151), .ZN(n149) );
  OAI21_X1 U1554 ( .B1(n153), .B2(n191), .A(n154), .ZN(n152) );
  XOR2_X1 U1555 ( .A(a[6]), .B(a[7]), .Z(n858) );
  OAI21_X1 U1556 ( .B1(n207), .B2(n235), .A(n208), .ZN(n206) );
  XOR2_X1 U1557 ( .A(a[14]), .B(a[15]), .Z(n854) );
  INV_X1 U1558 ( .A(n268), .ZN(n267) );
  AOI21_X1 U1559 ( .B1(n273), .B2(n1000), .A(n270), .ZN(n268) );
  XOR2_X1 U1560 ( .A(a[2]), .B(a[3]), .Z(n860) );
  XOR2_X1 U1561 ( .A(a[12]), .B(a[13]), .Z(n855) );
  AOI21_X1 U1562 ( .B1(n155), .B2(n180), .A(n156), .ZN(n154) );
  NAND2_X1 U1563 ( .A1(n1017), .A2(n155), .ZN(n153) );
  XOR2_X1 U1564 ( .A(a[10]), .B(a[11]), .Z(n856) );
  XNOR2_X1 U1565 ( .A(n1054), .B(n75), .ZN(product[9]) );
  XOR2_X1 U1566 ( .A(a[4]), .B(a[5]), .Z(n859) );
  XOR2_X1 U1567 ( .A(a[0]), .B(a[1]), .Z(n861) );
  XNOR2_X1 U1568 ( .A(a[2]), .B(a[1]), .ZN(n876) );
  XOR2_X1 U1569 ( .A(a[8]), .B(a[9]), .Z(n857) );
  AOI21_X1 U1570 ( .B1(n1052), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U1571 ( .B1(n1052), .B2(n94), .A(n95), .ZN(n93) );
  AOI21_X1 U1572 ( .B1(n51), .B2(n147), .A(n148), .ZN(n146) );
  AOI21_X1 U1573 ( .B1(n1052), .B2(n131), .A(n132), .ZN(n130) );
  AOI21_X1 U1574 ( .B1(n1052), .B2(n160), .A(n161), .ZN(n159) );
  AOI21_X1 U1575 ( .B1(n1052), .B2(n140), .A(n141), .ZN(n139) );
  AOI21_X1 U1576 ( .B1(n1052), .B2(n118), .A(n119), .ZN(n117) );
  AOI21_X1 U1577 ( .B1(n51), .B2(n193), .A(n194), .ZN(n192) );
  AOI21_X1 U1578 ( .B1(n1052), .B2(n107), .A(n108), .ZN(n106) );
  XNOR2_X1 U1579 ( .A(n1052), .B(n65), .ZN(product[19]) );
  AOI21_X1 U1580 ( .B1(n51), .B2(n184), .A(n185), .ZN(n183) );
  XOR2_X1 U1581 ( .A(n1005), .B(n76), .Z(product[8]) );
  AOI21_X1 U1582 ( .B1(n1052), .B2(n313), .A(n203), .ZN(n201) );
  OAI21_X1 U1583 ( .B1(n157), .B2(n169), .A(n158), .ZN(n156) );
  XNOR2_X1 U1584 ( .A(n281), .B(n77), .ZN(product[7]) );
  NOR2_X1 U1585 ( .A1(n168), .A2(n157), .ZN(n155) );
  XOR2_X1 U1586 ( .A(n78), .B(n1038), .Z(product[6]) );
  AOI21_X1 U1587 ( .B1(n51), .B2(n171), .A(n172), .ZN(n170) );
  OR2_X1 U1588 ( .A1(n1069), .A2(n885), .ZN(n837) );
  NAND2_X1 U1589 ( .A1(n541), .A2(n572), .ZN(n296) );
endmodule


module datapath_DW_mult_tc_14 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n3, n4, n5, n6, n7, n10, n11, n12, n15, n17, n18, n19, n22, n23,
         n24, n25, n27, n28, n29, n30, n34, n35, n36, n37, n39, n40, n41, n42,
         n43, n45, n46, n47, n48, n49, n65, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n84, n85, n86, n87, n88, n90, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n103, n105, n106, n107,
         n108, n109, n110, n114, n116, n117, n118, n119, n122, n123, n124,
         n125, n127, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n143, n144, n145, n146, n147, n148, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n180, n182, n183, n184, n185,
         n188, n189, n190, n191, n192, n193, n195, n196, n197, n198, n199,
         n200, n201, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n217, n218, n219, n220, n221, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n246, n247, n249, n250, n252,
         n253, n254, n255, n256, n257, n259, n261, n262, n264, n266, n267,
         n268, n270, n272, n273, n274, n275, n276, n278, n280, n281, n282,
         n283, n284, n286, n288, n289, n290, n291, n292, n294, n296, n297,
         n298, n299, n301, n306, n308, n312, n313, n316, n318, n320, n324,
         n326, n328, n330, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n545, n546, n548, n549, n551, n552, n554,
         n555, n557, n558, n560, n561, n563, n564, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n884, n885, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066;
  assign product[31] = n84;

  FA_X1 U364 ( .A(n575), .B(n338), .CI(n590), .CO(n334), .S(n335) );
  FA_X1 U365 ( .A(n339), .B(n576), .CI(n342), .CO(n336), .S(n337) );
  FA_X1 U367 ( .A(n346), .B(n577), .CI(n343), .CO(n340), .S(n341) );
  FA_X1 U368 ( .A(n591), .B(n348), .CI(n606), .CO(n342), .S(n343) );
  FA_X1 U369 ( .A(n347), .B(n354), .CI(n352), .CO(n344), .S(n345) );
  FA_X1 U370 ( .A(n578), .B(n592), .CI(n349), .CO(n346), .S(n347) );
  FA_X1 U372 ( .A(n358), .B(n355), .CI(n353), .CO(n350), .S(n351) );
  FA_X1 U373 ( .A(n362), .B(n607), .CI(n360), .CO(n352), .S(n353) );
  FA_X1 U374 ( .A(n593), .B(n579), .CI(n622), .CO(n354), .S(n355) );
  FA_X1 U375 ( .A(n359), .B(n361), .CI(n366), .CO(n356), .S(n357) );
  FA_X1 U376 ( .A(n370), .B(n363), .CI(n368), .CO(n358), .S(n359) );
  FA_X1 U377 ( .A(n580), .B(n594), .CI(n608), .CO(n360), .S(n361) );
  FA_X1 U379 ( .A(n367), .B(n376), .CI(n374), .CO(n364), .S(n365) );
  FA_X1 U380 ( .A(n369), .B(n378), .CI(n371), .CO(n366), .S(n367) );
  FA_X1 U381 ( .A(n595), .B(n380), .CI(n609), .CO(n368), .S(n369) );
  FA_X1 U382 ( .A(n623), .B(n581), .CI(n638), .CO(n370), .S(n371) );
  FA_X1 U383 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  FA_X1 U384 ( .A(n379), .B(n388), .CI(n386), .CO(n374), .S(n375) );
  FA_X1 U385 ( .A(n381), .B(n610), .CI(n390), .CO(n376), .S(n377) );
  FA_X1 U386 ( .A(n624), .B(n596), .CI(n582), .CO(n378), .S(n379) );
  FA_X1 U388 ( .A(n394), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U391 ( .A(n597), .B(n639), .CI(n611), .CO(n388), .S(n389) );
  FA_X1 U392 ( .A(n1026), .B(n583), .CI(n654), .CO(n390), .S(n391) );
  FA_X1 U393 ( .A(n406), .B(n397), .CI(n395), .CO(n392), .S(n393) );
  FA_X1 U394 ( .A(n410), .B(n399), .CI(n408), .CO(n394), .S(n395) );
  FA_X1 U396 ( .A(n584), .B(n598), .CI(n403), .CO(n398), .S(n399) );
  FA_X1 U397 ( .A(n612), .B(n626), .CI(n640), .CO(n400), .S(n401) );
  FA_X1 U400 ( .A(n411), .B(n422), .CI(n420), .CO(n406), .S(n407) );
  FA_X1 U401 ( .A(n413), .B(n424), .CI(n415), .CO(n408), .S(n409) );
  FA_X1 U402 ( .A(n613), .B(n627), .CI(n426), .CO(n410), .S(n411) );
  FA_X1 U403 ( .A(n655), .B(n641), .CI(n599), .CO(n412), .S(n413) );
  FA_X1 U404 ( .A(n670), .B(n585), .CI(n428), .CO(n414), .S(n415) );
  FA_X1 U405 ( .A(n432), .B(n421), .CI(n419), .CO(n416), .S(n417) );
  FA_X1 U406 ( .A(n423), .B(n436), .CI(n434), .CO(n418), .S(n419) );
  FA_X1 U407 ( .A(n425), .B(n438), .CI(n427), .CO(n420), .S(n421) );
  FA_X1 U408 ( .A(n442), .B(n429), .CI(n440), .CO(n422), .S(n423) );
  FA_X1 U409 ( .A(n600), .B(n642), .CI(n628), .CO(n424), .S(n425) );
  FA_X1 U410 ( .A(n586), .B(n614), .CI(n656), .CO(n426), .S(n427) );
  FA_X1 U413 ( .A(n448), .B(n450), .CI(n437), .CO(n432), .S(n433) );
  FA_X1 U415 ( .A(n443), .B(n971), .CI(n454), .CO(n436), .S(n437) );
  FA_X1 U416 ( .A(n671), .B(n657), .CI(n615), .CO(n438), .S(n439) );
  FA_X1 U417 ( .A(n587), .B(n629), .CI(n686), .CO(n440), .S(n441) );
  FA_X1 U420 ( .A(n449), .B(n460), .CI(n447), .CO(n444), .S(n445) );
  FA_X1 U421 ( .A(n462), .B(n455), .CI(n451), .CO(n446), .S(n447) );
  FA_X1 U423 ( .A(n457), .B(n672), .CI(n468), .CO(n450), .S(n451) );
  FA_X1 U424 ( .A(n687), .B(n630), .CI(n658), .CO(n452), .S(n453) );
  FA_X1 U425 ( .A(n602), .B(n644), .CI(n616), .CO(n454), .S(n455) );
  FA_X1 U427 ( .A(n463), .B(n472), .CI(n461), .CO(n458), .S(n459) );
  FA_X1 U428 ( .A(n465), .B(n467), .CI(n474), .CO(n460), .S(n461) );
  FA_X1 U429 ( .A(n476), .B(n478), .CI(n469), .CO(n462), .S(n463) );
  FA_X1 U430 ( .A(n645), .B(n659), .CI(n480), .CO(n464), .S(n465) );
  FA_X1 U431 ( .A(n603), .B(n673), .CI(n631), .CO(n466), .S(n467) );
  FA_X1 U432 ( .A(n589), .B(n688), .CI(n617), .CO(n468), .S(n469) );
  FA_X1 U434 ( .A(n479), .B(n477), .CI(n486), .CO(n472), .S(n473) );
  FA_X1 U435 ( .A(n490), .B(n481), .CI(n488), .CO(n474), .S(n475) );
  FA_X1 U436 ( .A(n618), .B(n660), .CI(n632), .CO(n476), .S(n477) );
  FA_X1 U437 ( .A(n674), .B(n689), .CI(n646), .CO(n478), .S(n479) );
  HA_X1 U438 ( .A(n567), .B(n604), .CO(n480), .S(n481) );
  FA_X1 U439 ( .A(n487), .B(n494), .CI(n485), .CO(n482), .S(n483) );
  FA_X1 U440 ( .A(n489), .B(n491), .CI(n496), .CO(n484), .S(n485) );
  FA_X1 U441 ( .A(n500), .B(n661), .CI(n498), .CO(n486), .S(n487) );
  FA_X1 U442 ( .A(n619), .B(n675), .CI(n647), .CO(n488), .S(n489) );
  FA_X1 U443 ( .A(n690), .B(n605), .CI(n633), .CO(n490), .S(n491) );
  FA_X1 U444 ( .A(n504), .B(n495), .CI(n497), .CO(n492), .S(n493) );
  FA_X1 U445 ( .A(n506), .B(n508), .CI(n499), .CO(n494), .S(n495) );
  FA_X1 U446 ( .A(n648), .B(n676), .CI(n501), .CO(n496), .S(n497) );
  FA_X1 U447 ( .A(n634), .B(n691), .CI(n662), .CO(n498), .S(n499) );
  HA_X1 U448 ( .A(n568), .B(n620), .CO(n500), .S(n501) );
  FA_X1 U450 ( .A(n514), .B(n516), .CI(n509), .CO(n504), .S(n505) );
  FA_X1 U451 ( .A(n635), .B(n677), .CI(n663), .CO(n506), .S(n507) );
  FA_X1 U452 ( .A(n649), .B(n621), .CI(n692), .CO(n508), .S(n509) );
  FA_X1 U453 ( .A(n515), .B(n520), .CI(n513), .CO(n510), .S(n511) );
  FA_X1 U454 ( .A(n517), .B(n693), .CI(n522), .CO(n512), .S(n513) );
  FA_X1 U455 ( .A(n650), .B(n664), .CI(n678), .CO(n514), .S(n515) );
  HA_X1 U456 ( .A(n569), .B(n636), .CO(n516), .S(n517) );
  FA_X1 U457 ( .A(n523), .B(n526), .CI(n521), .CO(n518), .S(n519) );
  FA_X1 U458 ( .A(n651), .B(n679), .CI(n528), .CO(n520), .S(n521) );
  FA_X1 U459 ( .A(n665), .B(n637), .CI(n694), .CO(n522), .S(n523) );
  FA_X1 U460 ( .A(n532), .B(n529), .CI(n527), .CO(n524), .S(n525) );
  FA_X1 U461 ( .A(n666), .B(n695), .CI(n680), .CO(n526), .S(n527) );
  HA_X1 U462 ( .A(n570), .B(n652), .CO(n528), .S(n529) );
  FA_X1 U463 ( .A(n536), .B(n667), .CI(n533), .CO(n530), .S(n531) );
  FA_X1 U464 ( .A(n696), .B(n653), .CI(n681), .CO(n532), .S(n533) );
  FA_X1 U465 ( .A(n682), .B(n697), .CI(n537), .CO(n534), .S(n535) );
  HA_X1 U466 ( .A(n571), .B(n668), .CO(n536), .S(n537) );
  FA_X1 U467 ( .A(n698), .B(n669), .CI(n683), .CO(n538), .S(n539) );
  HA_X1 U468 ( .A(n684), .B(n699), .CO(n540), .S(n541) );
  INV_X1 U822 ( .A(n879), .ZN(n953) );
  CLKBUF_X3 U823 ( .A(a[13]), .Z(n37) );
  OAI22_X1 U824 ( .A1(n47), .A2(n717), .B1(n45), .B2(n716), .ZN(n954) );
  INV_X1 U825 ( .A(n878), .ZN(n955) );
  CLKBUF_X3 U826 ( .A(a[15]), .Z(n43) );
  AND2_X2 U827 ( .A1(n483), .A2(n492), .ZN(n956) );
  INV_X4 U828 ( .A(n956), .ZN(n253) );
  BUF_X1 U829 ( .A(n863), .Z(n41) );
  NOR2_X2 U830 ( .A1(n373), .A2(n382), .ZN(n190) );
  AOI21_X2 U831 ( .B1(n198), .B2(n151), .A(n152), .ZN(n150) );
  BUF_X2 U832 ( .A(a[5]), .Z(n1057) );
  BUF_X2 U833 ( .A(a[11]), .Z(n957) );
  CLKBUF_X1 U834 ( .A(a[11]), .Z(n1058) );
  NOR2_X1 U835 ( .A1(n974), .A2(n416), .ZN(n958) );
  NOR2_X1 U836 ( .A1(n974), .A2(n416), .ZN(n211) );
  OR2_X1 U837 ( .A1(n227), .A2(n232), .ZN(n959) );
  NOR2_X2 U838 ( .A1(n459), .A2(n470), .ZN(n238) );
  BUF_X1 U839 ( .A(n865), .Z(n29) );
  CLKBUF_X1 U840 ( .A(n398), .Z(n960) );
  CLKBUF_X1 U841 ( .A(n845), .Z(n961) );
  CLKBUF_X3 U842 ( .A(b[2]), .Z(n851) );
  BUF_X4 U843 ( .A(n872), .Z(n34) );
  XOR2_X1 U844 ( .A(n441), .B(n452), .Z(n962) );
  XOR2_X1 U845 ( .A(n439), .B(n962), .Z(n435) );
  NAND2_X1 U846 ( .A1(n439), .A2(n441), .ZN(n963) );
  NAND2_X1 U847 ( .A1(n439), .A2(n452), .ZN(n964) );
  NAND2_X1 U848 ( .A1(n441), .A2(n452), .ZN(n965) );
  NAND3_X1 U849 ( .A1(n963), .A2(n964), .A3(n965), .ZN(n434) );
  XOR2_X1 U850 ( .A(n453), .B(n466), .Z(n966) );
  XOR2_X1 U851 ( .A(n464), .B(n966), .Z(n449) );
  NAND2_X1 U852 ( .A1(n464), .A2(n453), .ZN(n967) );
  NAND2_X1 U853 ( .A1(n464), .A2(n466), .ZN(n968) );
  NAND2_X1 U854 ( .A1(n453), .A2(n466), .ZN(n969) );
  NAND3_X1 U855 ( .A1(n967), .A2(n968), .A3(n969), .ZN(n448) );
  BUF_X1 U856 ( .A(n866), .Z(n24) );
  OR2_X1 U857 ( .A1(n503), .A2(n510), .ZN(n970) );
  AND2_X1 U858 ( .A1(n566), .A2(n954), .ZN(n971) );
  NAND2_X1 U859 ( .A1(n197), .A2(n151), .ZN(n972) );
  CLKBUF_X2 U860 ( .A(b[7]), .Z(n846) );
  CLKBUF_X1 U861 ( .A(n205), .Z(n973) );
  XNOR2_X1 U862 ( .A(n407), .B(n1027), .ZN(n974) );
  XOR2_X1 U863 ( .A(n512), .B(n507), .Z(n975) );
  XOR2_X1 U864 ( .A(n505), .B(n975), .Z(n503) );
  NAND2_X1 U865 ( .A1(n505), .A2(n512), .ZN(n976) );
  NAND2_X1 U866 ( .A1(n505), .A2(n507), .ZN(n977) );
  NAND2_X1 U867 ( .A1(n512), .A2(n507), .ZN(n978) );
  NAND3_X1 U868 ( .A1(n976), .A2(n977), .A3(n978), .ZN(n502) );
  BUF_X1 U869 ( .A(n850), .Z(n979) );
  OR2_X2 U870 ( .A1(n493), .A2(n502), .ZN(n1063) );
  CLKBUF_X2 U871 ( .A(n873), .Z(n27) );
  CLKBUF_X3 U872 ( .A(n873), .Z(n28) );
  BUF_X1 U873 ( .A(b[15]), .Z(n838) );
  NOR2_X1 U874 ( .A1(n218), .A2(n958), .ZN(n980) );
  XOR2_X1 U875 ( .A(n588), .B(n566), .Z(n457) );
  CLKBUF_X3 U876 ( .A(b[1]), .Z(n852) );
  CLKBUF_X1 U877 ( .A(b[13]), .Z(n1019) );
  CLKBUF_X1 U878 ( .A(b[13]), .Z(n1020) );
  BUF_X2 U879 ( .A(n841), .Z(n1004) );
  BUF_X2 U880 ( .A(n863), .Z(n42) );
  BUF_X2 U881 ( .A(b[8]), .Z(n845) );
  BUF_X2 U882 ( .A(b[4]), .Z(n849) );
  BUF_X2 U883 ( .A(n870), .Z(n45) );
  BUF_X2 U884 ( .A(n870), .Z(n46) );
  OAI22_X1 U885 ( .A1(n48), .A2(n703), .B1(n46), .B2(n702), .ZN(n332) );
  NOR2_X1 U886 ( .A1(n144), .A2(n137), .ZN(n135) );
  BUF_X1 U887 ( .A(n877), .Z(n4) );
  INV_X1 U888 ( .A(a[0]), .ZN(n877) );
  INV_X1 U889 ( .A(n137), .ZN(n306) );
  XOR2_X1 U890 ( .A(n412), .B(n414), .Z(n981) );
  XOR2_X1 U891 ( .A(n401), .B(n981), .Z(n397) );
  NAND2_X1 U892 ( .A1(n401), .A2(n412), .ZN(n982) );
  NAND2_X1 U893 ( .A1(n401), .A2(n414), .ZN(n983) );
  NAND2_X1 U894 ( .A1(n412), .A2(n414), .ZN(n984) );
  NAND3_X1 U895 ( .A1(n982), .A2(n983), .A3(n984), .ZN(n396) );
  XOR2_X1 U896 ( .A(n960), .B(n625), .Z(n985) );
  XOR2_X1 U897 ( .A(n400), .B(n985), .Z(n387) );
  NAND2_X1 U898 ( .A1(n400), .A2(n398), .ZN(n986) );
  NAND2_X1 U899 ( .A1(n400), .A2(n625), .ZN(n987) );
  NAND2_X1 U900 ( .A1(n398), .A2(n625), .ZN(n988) );
  NAND3_X1 U901 ( .A1(n986), .A2(n987), .A3(n988), .ZN(n386) );
  XOR2_X1 U902 ( .A(n484), .B(n475), .Z(n989) );
  XOR2_X1 U903 ( .A(n473), .B(n989), .Z(n471) );
  NAND2_X1 U904 ( .A1(n473), .A2(n484), .ZN(n990) );
  NAND2_X1 U905 ( .A1(n473), .A2(n475), .ZN(n991) );
  NAND2_X1 U906 ( .A1(n484), .A2(n475), .ZN(n992) );
  NAND3_X1 U907 ( .A1(n990), .A2(n991), .A3(n992), .ZN(n470) );
  OR2_X1 U908 ( .A1(n337), .A2(n340), .ZN(n993) );
  OR2_X1 U909 ( .A1(n334), .A2(n333), .ZN(n994) );
  OR2_X1 U910 ( .A1(n574), .A2(n332), .ZN(n995) );
  OR2_X1 U911 ( .A1(n541), .A2(n572), .ZN(n996) );
  AND2_X1 U912 ( .A1(n1002), .A2(n301), .ZN(product[1]) );
  OR2_X1 U913 ( .A1(n336), .A2(n335), .ZN(n998) );
  OR2_X1 U914 ( .A1(n511), .A2(n518), .ZN(n999) );
  OR2_X1 U915 ( .A1(n525), .A2(n530), .ZN(n1000) );
  OR2_X1 U916 ( .A1(n535), .A2(n538), .ZN(n1001) );
  BUF_X2 U917 ( .A(b[9]), .Z(n844) );
  OR2_X1 U918 ( .A1(n701), .A2(n573), .ZN(n1002) );
  NOR2_X1 U919 ( .A1(n364), .A2(n357), .ZN(n168) );
  NOR2_X1 U920 ( .A1(n345), .A2(n350), .ZN(n144) );
  BUF_X1 U921 ( .A(n850), .Z(n1003) );
  BUF_X1 U922 ( .A(b[3]), .Z(n850) );
  CLKBUF_X1 U923 ( .A(n843), .Z(n1005) );
  BUF_X2 U924 ( .A(b[10]), .Z(n843) );
  CLKBUF_X3 U925 ( .A(b[11]), .Z(n842) );
  CLKBUF_X1 U926 ( .A(n839), .Z(n1006) );
  XOR2_X1 U927 ( .A(n391), .B(n389), .Z(n1007) );
  XOR2_X1 U928 ( .A(n396), .B(n1007), .Z(n385) );
  NAND2_X1 U929 ( .A1(n396), .A2(n391), .ZN(n1008) );
  NAND2_X1 U930 ( .A1(n396), .A2(n389), .ZN(n1009) );
  NAND2_X1 U931 ( .A1(n391), .A2(n389), .ZN(n1010) );
  NAND3_X1 U932 ( .A1(n1008), .A2(n1009), .A3(n1010), .ZN(n384) );
  CLKBUF_X1 U933 ( .A(n838), .Z(n1011) );
  OAI22_X1 U934 ( .A1(n30), .A2(n754), .B1(n28), .B2(n753), .ZN(n362) );
  AOI21_X1 U935 ( .B1(n273), .B2(n999), .A(n270), .ZN(n268) );
  OAI21_X1 U936 ( .B1(n199), .B2(n205), .A(n200), .ZN(n1012) );
  NOR2_X2 U937 ( .A1(n383), .A2(n392), .ZN(n199) );
  CLKBUF_X3 U938 ( .A(n869), .Z(n1013) );
  CLKBUF_X1 U939 ( .A(n869), .Z(n6) );
  XOR2_X1 U940 ( .A(n1050), .B(n838), .Z(n787) );
  BUF_X1 U941 ( .A(n1047), .Z(n1014) );
  CLKBUF_X1 U942 ( .A(n1047), .Z(n1015) );
  BUF_X1 U943 ( .A(n1047), .Z(n1060) );
  CLKBUF_X2 U944 ( .A(n49), .Z(n1016) );
  XNOR2_X1 U945 ( .A(n159), .B(n1017), .ZN(product[24]) );
  AND2_X1 U946 ( .A1(n308), .A2(n158), .ZN(n1017) );
  CLKBUF_X1 U947 ( .A(n276), .Z(n1018) );
  CLKBUF_X1 U948 ( .A(b[13]), .Z(n840) );
  CLKBUF_X1 U949 ( .A(n232), .Z(n1021) );
  OAI22_X1 U950 ( .A1(n12), .A2(n805), .B1(n10), .B2(n804), .ZN(n428) );
  OAI21_X1 U951 ( .B1(n1034), .B2(n233), .A(n228), .ZN(n1022) );
  CLKBUF_X1 U952 ( .A(n284), .Z(n1023) );
  NOR2_X1 U953 ( .A1(n241), .A2(n238), .ZN(n236) );
  XNOR2_X1 U954 ( .A(n433), .B(n1024), .ZN(n431) );
  XNOR2_X1 U955 ( .A(n446), .B(n435), .ZN(n1024) );
  OAI21_X1 U956 ( .B1(n256), .B2(n268), .A(n257), .ZN(n1025) );
  OAI22_X1 U957 ( .A1(n17), .A2(n788), .B1(n15), .B2(n787), .ZN(n1026) );
  XNOR2_X1 U958 ( .A(n418), .B(n409), .ZN(n1027) );
  CLKBUF_X2 U959 ( .A(n49), .Z(n1065) );
  BUF_X2 U960 ( .A(n49), .Z(n1066) );
  NAND2_X1 U961 ( .A1(n407), .A2(n418), .ZN(n1028) );
  NAND2_X1 U962 ( .A1(n407), .A2(n409), .ZN(n1029) );
  NAND2_X1 U963 ( .A1(n418), .A2(n409), .ZN(n1030) );
  NAND3_X1 U964 ( .A1(n1028), .A2(n1029), .A3(n1030), .ZN(n404) );
  XNOR2_X1 U965 ( .A(n117), .B(n1031), .ZN(product[28]) );
  AND2_X1 U966 ( .A1(n998), .A2(n116), .ZN(n1031) );
  CLKBUF_X1 U967 ( .A(n218), .Z(n1032) );
  OR2_X1 U968 ( .A1(n974), .A2(n416), .ZN(n1033) );
  NOR2_X1 U969 ( .A1(n431), .A2(n444), .ZN(n1034) );
  NOR2_X1 U970 ( .A1(n431), .A2(n444), .ZN(n227) );
  XNOR2_X1 U971 ( .A(n201), .B(n1035), .ZN(product[20]) );
  AND2_X1 U972 ( .A1(n312), .A2(n200), .ZN(n1035) );
  XNOR2_X1 U973 ( .A(n183), .B(n1036), .ZN(product[22]) );
  AND2_X1 U974 ( .A1(n175), .A2(n182), .ZN(n1036) );
  CLKBUF_X1 U975 ( .A(n273), .Z(n1037) );
  XNOR2_X1 U976 ( .A(n192), .B(n1038), .ZN(product[21]) );
  AND2_X1 U977 ( .A1(n188), .A2(n191), .ZN(n1038) );
  BUF_X2 U978 ( .A(n867), .Z(n17) );
  OR2_X2 U979 ( .A1(n471), .A2(n482), .ZN(n1039) );
  NAND2_X1 U980 ( .A1(n433), .A2(n446), .ZN(n1040) );
  NAND2_X1 U981 ( .A1(n433), .A2(n435), .ZN(n1041) );
  NAND2_X1 U982 ( .A1(n446), .A2(n435), .ZN(n1042) );
  NAND3_X1 U983 ( .A1(n1040), .A2(n1041), .A3(n1042), .ZN(n430) );
  XNOR2_X1 U984 ( .A(n170), .B(n1043), .ZN(product[23]) );
  AND2_X1 U985 ( .A1(n167), .A2(n169), .ZN(n1043) );
  BUF_X1 U986 ( .A(n1060), .Z(n1059) );
  XNOR2_X1 U987 ( .A(n146), .B(n1044), .ZN(product[25]) );
  AND2_X1 U988 ( .A1(n143), .A2(n145), .ZN(n1044) );
  XOR2_X1 U989 ( .A(a[4]), .B(a[5]), .Z(n859) );
  OAI21_X1 U990 ( .B1(n1034), .B2(n233), .A(n228), .ZN(n226) );
  OR2_X1 U991 ( .A1(n365), .A2(n372), .ZN(n1045) );
  XNOR2_X1 U992 ( .A(n130), .B(n1046), .ZN(product[27]) );
  AND2_X1 U993 ( .A1(n993), .A2(n129), .ZN(n1046) );
  OAI21_X1 U994 ( .B1(n235), .B2(n207), .A(n208), .ZN(n1047) );
  AOI21_X1 U995 ( .B1(n236), .B2(n255), .A(n237), .ZN(n1048) );
  AOI21_X1 U996 ( .B1(n236), .B2(n1025), .A(n237), .ZN(n1049) );
  INV_X1 U997 ( .A(a[5]), .ZN(n1050) );
  XNOR2_X1 U998 ( .A(n213), .B(n1051), .ZN(product[18]) );
  AND2_X1 U999 ( .A1(n1033), .A2(n212), .ZN(n1051) );
  XNOR2_X1 U1000 ( .A(n220), .B(n1052), .ZN(product[17]) );
  AND2_X1 U1001 ( .A1(n217), .A2(n219), .ZN(n1052) );
  XNOR2_X1 U1002 ( .A(n229), .B(n1053), .ZN(product[16]) );
  AND2_X1 U1003 ( .A1(n316), .A2(n228), .ZN(n1053) );
  NAND2_X1 U1004 ( .A1(n188), .A2(n175), .ZN(n173) );
  INV_X1 U1005 ( .A(n1045), .ZN(n177) );
  NOR2_X1 U1006 ( .A1(n393), .A2(n404), .ZN(n204) );
  INV_X1 U1007 ( .A(n190), .ZN(n188) );
  NAND2_X1 U1008 ( .A1(n135), .A2(n993), .ZN(n124) );
  XNOR2_X1 U1009 ( .A(n93), .B(n1054), .ZN(product[30]) );
  AND2_X1 U1010 ( .A1(n995), .A2(n92), .ZN(n1054) );
  XNOR2_X1 U1011 ( .A(n106), .B(n1055), .ZN(product[29]) );
  AND2_X1 U1012 ( .A1(n994), .A2(n105), .ZN(n1055) );
  NOR2_X1 U1013 ( .A1(n351), .A2(n356), .ZN(n157) );
  NOR2_X1 U1014 ( .A1(n519), .A2(n524), .ZN(n274) );
  NAND2_X1 U1015 ( .A1(n373), .A2(n382), .ZN(n191) );
  NOR2_X1 U1016 ( .A1(n700), .A2(n685), .ZN(n298) );
  NOR2_X1 U1017 ( .A1(n539), .A2(n540), .ZN(n290) );
  BUF_X1 U1018 ( .A(n877), .Z(n3) );
  BUF_X2 U1019 ( .A(b[12]), .Z(n841) );
  BUF_X2 U1020 ( .A(b[5]), .Z(n848) );
  INV_X1 U1021 ( .A(n98), .ZN(n96) );
  INV_X1 U1022 ( .A(n177), .ZN(n175) );
  NOR2_X1 U1023 ( .A1(n972), .A2(n96), .ZN(n94) );
  NOR2_X1 U1024 ( .A1(n972), .A2(n124), .ZN(n118) );
  NOR2_X1 U1025 ( .A1(n959), .A2(n1032), .ZN(n214) );
  NOR2_X1 U1026 ( .A1(n195), .A2(n173), .ZN(n171) );
  NOR2_X1 U1027 ( .A1(n195), .A2(n190), .ZN(n184) );
  NOR2_X1 U1028 ( .A1(n195), .A2(n162), .ZN(n160) );
  INV_X1 U1029 ( .A(n1022), .ZN(n224) );
  INV_X1 U1030 ( .A(n972), .ZN(n147) );
  NAND2_X1 U1031 ( .A1(n313), .A2(n973), .ZN(n65) );
  INV_X1 U1032 ( .A(n204), .ZN(n313) );
  XNOR2_X1 U1033 ( .A(n240), .B(n70), .ZN(product[14]) );
  NAND2_X1 U1034 ( .A1(n318), .A2(n239), .ZN(n70) );
  INV_X1 U1035 ( .A(n238), .ZN(n318) );
  INV_X1 U1036 ( .A(n1012), .ZN(n196) );
  NOR2_X1 U1037 ( .A1(n177), .A2(n166), .ZN(n164) );
  NOR2_X1 U1038 ( .A1(n124), .A2(n100), .ZN(n98) );
  INV_X1 U1039 ( .A(n197), .ZN(n195) );
  OAI21_X1 U1040 ( .B1(n150), .B2(n124), .A(n125), .ZN(n119) );
  OAI21_X1 U1041 ( .B1(n196), .B2(n173), .A(n174), .ZN(n172) );
  AOI21_X1 U1042 ( .B1(n189), .B2(n175), .A(n176), .ZN(n174) );
  INV_X1 U1043 ( .A(n178), .ZN(n176) );
  OAI21_X1 U1044 ( .B1(n196), .B2(n190), .A(n191), .ZN(n185) );
  NAND2_X1 U1045 ( .A1(n164), .A2(n188), .ZN(n162) );
  OAI21_X1 U1046 ( .B1(n224), .B2(n1032), .A(n219), .ZN(n215) );
  INV_X1 U1047 ( .A(n124), .ZN(n122) );
  NOR2_X1 U1048 ( .A1(n972), .A2(n144), .ZN(n140) );
  NOR2_X1 U1049 ( .A1(n972), .A2(n133), .ZN(n131) );
  INV_X1 U1050 ( .A(n180), .ZN(n178) );
  INV_X1 U1051 ( .A(n150), .ZN(n148) );
  INV_X1 U1052 ( .A(n233), .ZN(n231) );
  NAND2_X1 U1053 ( .A1(n122), .A2(n998), .ZN(n109) );
  INV_X1 U1054 ( .A(n973), .ZN(n203) );
  NAND2_X1 U1055 ( .A1(n324), .A2(n275), .ZN(n76) );
  INV_X1 U1056 ( .A(n274), .ZN(n324) );
  NAND2_X1 U1057 ( .A1(n999), .A2(n272), .ZN(n75) );
  XOR2_X1 U1058 ( .A(n254), .B(n72), .Z(product[12]) );
  XNOR2_X1 U1059 ( .A(n267), .B(n74), .ZN(product[10]) );
  NAND2_X1 U1060 ( .A1(n970), .A2(n266), .ZN(n74) );
  INV_X1 U1061 ( .A(n195), .ZN(n193) );
  INV_X1 U1062 ( .A(n272), .ZN(n270) );
  NAND2_X1 U1063 ( .A1(n1063), .A2(n970), .ZN(n256) );
  NOR2_X1 U1064 ( .A1(n204), .A2(n199), .ZN(n197) );
  XOR2_X1 U1065 ( .A(n262), .B(n73), .Z(product[11]) );
  NAND2_X1 U1066 ( .A1(n1063), .A2(n261), .ZN(n73) );
  AOI21_X1 U1067 ( .B1(n267), .B2(n970), .A(n264), .ZN(n262) );
  INV_X1 U1068 ( .A(n157), .ZN(n308) );
  INV_X1 U1069 ( .A(n199), .ZN(n312) );
  NAND2_X1 U1070 ( .A1(n393), .A2(n404), .ZN(n205) );
  NAND2_X1 U1071 ( .A1(n1039), .A2(n246), .ZN(n71) );
  AOI21_X1 U1072 ( .B1(n123), .B2(n998), .A(n114), .ZN(n110) );
  OAI21_X1 U1073 ( .B1(n196), .B2(n162), .A(n163), .ZN(n161) );
  AOI21_X1 U1074 ( .B1(n164), .B2(n189), .A(n165), .ZN(n163) );
  OAI21_X1 U1075 ( .B1(n178), .B2(n166), .A(n169), .ZN(n165) );
  OAI21_X1 U1076 ( .B1(n276), .B2(n274), .A(n275), .ZN(n273) );
  INV_X1 U1077 ( .A(n125), .ZN(n123) );
  OAI21_X1 U1078 ( .B1(n150), .B2(n96), .A(n97), .ZN(n95) );
  INV_X1 U1079 ( .A(n99), .ZN(n97) );
  OAI21_X1 U1080 ( .B1(n150), .B2(n133), .A(n134), .ZN(n132) );
  INV_X1 U1081 ( .A(n136), .ZN(n134) );
  NAND2_X1 U1082 ( .A1(n417), .A2(n430), .ZN(n219) );
  INV_X1 U1083 ( .A(n191), .ZN(n189) );
  NAND2_X1 U1084 ( .A1(n98), .A2(n995), .ZN(n87) );
  INV_X1 U1085 ( .A(n182), .ZN(n180) );
  NAND2_X1 U1086 ( .A1(n459), .A2(n470), .ZN(n239) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n994), .ZN(n100) );
  INV_X1 U1088 ( .A(n135), .ZN(n133) );
  NOR2_X1 U1089 ( .A1(n972), .A2(n87), .ZN(n85) );
  OAI21_X1 U1090 ( .B1(n150), .B2(n87), .A(n88), .ZN(n86) );
  INV_X1 U1091 ( .A(n167), .ZN(n166) );
  INV_X1 U1092 ( .A(n168), .ZN(n167) );
  INV_X1 U1093 ( .A(n144), .ZN(n143) );
  INV_X1 U1094 ( .A(n1061), .ZN(n246) );
  NAND2_X1 U1095 ( .A1(n326), .A2(n283), .ZN(n78) );
  NAND2_X1 U1096 ( .A1(n1001), .A2(n288), .ZN(n79) );
  NAND2_X1 U1097 ( .A1(n1000), .A2(n280), .ZN(n77) );
  INV_X1 U1098 ( .A(n280), .ZN(n278) );
  OAI21_X1 U1099 ( .B1(n125), .B2(n100), .A(n101), .ZN(n99) );
  AOI21_X1 U1100 ( .B1(n114), .B2(n994), .A(n103), .ZN(n101) );
  INV_X1 U1101 ( .A(n105), .ZN(n103) );
  XNOR2_X1 U1102 ( .A(n139), .B(n1056), .ZN(product[26]) );
  AND2_X1 U1103 ( .A1(n306), .A2(n138), .ZN(n1056) );
  AOI21_X1 U1104 ( .B1(n136), .B2(n993), .A(n127), .ZN(n125) );
  INV_X1 U1105 ( .A(n129), .ZN(n127) );
  AOI21_X1 U1106 ( .B1(n99), .B2(n995), .A(n90), .ZN(n88) );
  INV_X1 U1107 ( .A(n92), .ZN(n90) );
  NAND2_X1 U1108 ( .A1(n511), .A2(n518), .ZN(n272) );
  NAND2_X1 U1109 ( .A1(n357), .A2(n364), .ZN(n169) );
  NAND2_X1 U1110 ( .A1(n345), .A2(n350), .ZN(n145) );
  NAND2_X1 U1111 ( .A1(n351), .A2(n356), .ZN(n158) );
  NAND2_X1 U1112 ( .A1(n493), .A2(n502), .ZN(n261) );
  NAND2_X1 U1113 ( .A1(n503), .A2(n510), .ZN(n266) );
  INV_X1 U1114 ( .A(n116), .ZN(n114) );
  NAND2_X1 U1115 ( .A1(n328), .A2(n291), .ZN(n80) );
  INV_X1 U1116 ( .A(n290), .ZN(n328) );
  NAND2_X1 U1117 ( .A1(n330), .A2(n299), .ZN(n82) );
  INV_X1 U1118 ( .A(n298), .ZN(n330) );
  XNOR2_X1 U1119 ( .A(n81), .B(n297), .ZN(product[3]) );
  NAND2_X1 U1120 ( .A1(n996), .A2(n296), .ZN(n81) );
  NOR2_X1 U1121 ( .A1(n341), .A2(n344), .ZN(n137) );
  NAND2_X1 U1122 ( .A1(n574), .A2(n332), .ZN(n92) );
  INV_X1 U1123 ( .A(n332), .ZN(n333) );
  INV_X1 U1124 ( .A(n362), .ZN(n363) );
  NAND2_X1 U1125 ( .A1(n700), .A2(n685), .ZN(n299) );
  XNOR2_X1 U1126 ( .A(n643), .B(n601), .ZN(n443) );
  INV_X1 U1127 ( .A(n428), .ZN(n429) );
  OR2_X1 U1128 ( .A1(n643), .A2(n601), .ZN(n442) );
  NAND2_X1 U1129 ( .A1(n535), .A2(n538), .ZN(n288) );
  NAND2_X1 U1130 ( .A1(n337), .A2(n340), .ZN(n129) );
  NAND2_X1 U1131 ( .A1(n336), .A2(n335), .ZN(n116) );
  NAND2_X1 U1132 ( .A1(n334), .A2(n333), .ZN(n105) );
  NAND2_X1 U1133 ( .A1(n525), .A2(n530), .ZN(n280) );
  NAND2_X1 U1134 ( .A1(n341), .A2(n344), .ZN(n138) );
  AOI21_X1 U1135 ( .B1(n996), .B2(n297), .A(n294), .ZN(n292) );
  INV_X1 U1136 ( .A(n296), .ZN(n294) );
  OAI22_X1 U1137 ( .A1(n24), .A2(n771), .B1(n22), .B2(n770), .ZN(n380) );
  OAI22_X1 U1138 ( .A1(n42), .A2(n720), .B1(n40), .B2(n719), .ZN(n338) );
  OAI22_X1 U1139 ( .A1(n5), .A2(n835), .B1(n834), .B2(n3), .ZN(n700) );
  OAI22_X1 U1140 ( .A1(n36), .A2(n737), .B1(n34), .B2(n736), .ZN(n348) );
  OAI22_X1 U1141 ( .A1(n42), .A2(n731), .B1(n39), .B2(n730), .ZN(n601) );
  OAI22_X1 U1142 ( .A1(n23), .A2(n776), .B1(n22), .B2(n775), .ZN(n643) );
  OAI22_X1 U1143 ( .A1(n35), .A2(n745), .B1(n34), .B2(n744), .ZN(n614) );
  OAI22_X1 U1144 ( .A1(n47), .A2(n715), .B1(n45), .B2(n714), .ZN(n586) );
  OAI22_X1 U1145 ( .A1(n48), .A2(n704), .B1(n46), .B2(n703), .ZN(n575) );
  INV_X1 U1146 ( .A(n545), .ZN(n590) );
  AOI21_X1 U1147 ( .B1(n42), .B2(n40), .A(n719), .ZN(n545) );
  OAI22_X1 U1148 ( .A1(n48), .A2(n705), .B1(n46), .B2(n704), .ZN(n576) );
  INV_X1 U1149 ( .A(n338), .ZN(n339) );
  OAI22_X1 U1150 ( .A1(n48), .A2(n706), .B1(n46), .B2(n705), .ZN(n577) );
  AND2_X1 U1151 ( .A1(n1066), .A2(n558), .ZN(n669) );
  OAI22_X1 U1152 ( .A1(n11), .A2(n818), .B1(n10), .B2(n817), .ZN(n683) );
  OAI22_X1 U1153 ( .A1(n5), .A2(n833), .B1(n832), .B2(n3), .ZN(n698) );
  OAI22_X1 U1154 ( .A1(n30), .A2(n768), .B1(n27), .B2(n767), .ZN(n636) );
  OAI22_X1 U1155 ( .A1(n47), .A2(n717), .B1(n45), .B2(n716), .ZN(n588) );
  OR2_X1 U1156 ( .A1(n1066), .A2(n878), .ZN(n718) );
  OAI22_X1 U1157 ( .A1(n35), .A2(n747), .B1(n34), .B2(n746), .ZN(n616) );
  OAI22_X1 U1158 ( .A1(n23), .A2(n777), .B1(n22), .B2(n776), .ZN(n644) );
  OAI22_X1 U1159 ( .A1(n42), .A2(n732), .B1(n39), .B2(n731), .ZN(n602) );
  OAI22_X1 U1160 ( .A1(n29), .A2(n758), .B1(n28), .B2(n757), .ZN(n626) );
  OAI22_X1 U1161 ( .A1(n23), .A2(n773), .B1(n22), .B2(n772), .ZN(n640) );
  OAI22_X1 U1162 ( .A1(n36), .A2(n743), .B1(n34), .B2(n742), .ZN(n612) );
  OAI22_X1 U1163 ( .A1(n11), .A2(n813), .B1(n10), .B2(n812), .ZN(n678) );
  OAI22_X1 U1164 ( .A1(n23), .A2(n783), .B1(n22), .B2(n782), .ZN(n650) );
  OAI22_X1 U1165 ( .A1(n17), .A2(n798), .B1(n15), .B2(n797), .ZN(n664) );
  AOI21_X1 U1166 ( .B1(n24), .B2(n22), .A(n770), .ZN(n554) );
  XNOR2_X1 U1167 ( .A(n844), .B(n1058), .ZN(n742) );
  XNOR2_X1 U1168 ( .A(n957), .B(n845), .ZN(n743) );
  XNOR2_X1 U1169 ( .A(n1058), .B(n849), .ZN(n747) );
  OAI22_X1 U1170 ( .A1(n24), .A2(n775), .B1(n22), .B2(n774), .ZN(n642) );
  OAI22_X1 U1171 ( .A1(n41), .A2(n730), .B1(n39), .B2(n729), .ZN(n600) );
  OAI22_X1 U1172 ( .A1(n30), .A2(n760), .B1(n28), .B2(n759), .ZN(n628) );
  OAI22_X1 U1173 ( .A1(n47), .A2(n714), .B1(n45), .B2(n713), .ZN(n585) );
  INV_X1 U1174 ( .A(n560), .ZN(n670) );
  AOI21_X1 U1175 ( .B1(n12), .B2(n10), .A(n804), .ZN(n560) );
  AOI21_X1 U1176 ( .B1(n6), .B2(n4), .A(n821), .ZN(n563) );
  AOI21_X1 U1177 ( .B1(n30), .B2(n28), .A(n753), .ZN(n551) );
  XNOR2_X1 U1178 ( .A(n957), .B(n1006), .ZN(n737) );
  OAI22_X1 U1179 ( .A1(n35), .A2(n751), .B1(n34), .B2(n750), .ZN(n620) );
  XNOR2_X1 U1180 ( .A(n957), .B(n1065), .ZN(n751) );
  OAI22_X1 U1181 ( .A1(n18), .A2(n802), .B1(n15), .B2(n801), .ZN(n668) );
  OR2_X1 U1182 ( .A1(n1016), .A2(n1050), .ZN(n803) );
  XNOR2_X1 U1183 ( .A(n1057), .B(n848), .ZN(n797) );
  XNOR2_X1 U1184 ( .A(n1057), .B(n849), .ZN(n798) );
  XNOR2_X1 U1185 ( .A(n957), .B(n1005), .ZN(n741) );
  XNOR2_X1 U1186 ( .A(n957), .B(n1019), .ZN(n738) );
  XNOR2_X1 U1187 ( .A(n957), .B(n841), .ZN(n739) );
  XNOR2_X1 U1188 ( .A(n957), .B(n848), .ZN(n746) );
  XNOR2_X1 U1189 ( .A(n957), .B(n847), .ZN(n745) );
  OAI22_X1 U1190 ( .A1(n17), .A2(n801), .B1(n15), .B2(n800), .ZN(n667) );
  XNOR2_X1 U1191 ( .A(n1057), .B(n845), .ZN(n794) );
  XNOR2_X1 U1192 ( .A(n1057), .B(n844), .ZN(n793) );
  XNOR2_X1 U1193 ( .A(n1057), .B(n843), .ZN(n792) );
  XNOR2_X1 U1194 ( .A(n1057), .B(n1066), .ZN(n802) );
  AND2_X1 U1195 ( .A1(n1016), .A2(n561), .ZN(n685) );
  INV_X1 U1196 ( .A(n10), .ZN(n561) );
  OAI22_X1 U1197 ( .A1(n11), .A2(n817), .B1(n10), .B2(n816), .ZN(n682) );
  OAI22_X1 U1198 ( .A1(n1013), .A2(n832), .B1(n831), .B2(n3), .ZN(n697) );
  OAI22_X1 U1199 ( .A1(n48), .A2(n707), .B1(n46), .B2(n706), .ZN(n578) );
  OAI22_X1 U1200 ( .A1(n42), .A2(n722), .B1(n40), .B2(n721), .ZN(n592) );
  INV_X1 U1201 ( .A(n348), .ZN(n349) );
  OAI22_X1 U1202 ( .A1(n36), .A2(n740), .B1(n34), .B2(n739), .ZN(n609) );
  OAI22_X1 U1203 ( .A1(n42), .A2(n725), .B1(n40), .B2(n724), .ZN(n595) );
  OAI22_X1 U1204 ( .A1(n12), .A2(n806), .B1(n10), .B2(n805), .ZN(n671) );
  OAI22_X1 U1205 ( .A1(n35), .A2(n746), .B1(n34), .B2(n745), .ZN(n615) );
  OAI22_X1 U1206 ( .A1(n30), .A2(n759), .B1(n28), .B2(n758), .ZN(n627) );
  OAI22_X1 U1207 ( .A1(n35), .A2(n744), .B1(n34), .B2(n743), .ZN(n613) );
  OAI22_X1 U1208 ( .A1(n47), .A2(n711), .B1(n45), .B2(n710), .ZN(n582) );
  OAI22_X1 U1209 ( .A1(n42), .A2(n726), .B1(n40), .B2(n725), .ZN(n596) );
  OAI22_X1 U1210 ( .A1(n30), .A2(n756), .B1(n28), .B2(n755), .ZN(n624) );
  OAI22_X1 U1211 ( .A1(n48), .A2(n708), .B1(n46), .B2(n707), .ZN(n579) );
  OAI22_X1 U1212 ( .A1(n42), .A2(n723), .B1(n40), .B2(n722), .ZN(n593) );
  INV_X1 U1213 ( .A(n551), .ZN(n622) );
  OAI22_X1 U1214 ( .A1(n36), .A2(n742), .B1(n34), .B2(n741), .ZN(n611) );
  OAI22_X1 U1215 ( .A1(n23), .A2(n772), .B1(n22), .B2(n771), .ZN(n639) );
  OAI22_X1 U1216 ( .A1(n42), .A2(n727), .B1(n39), .B2(n726), .ZN(n597) );
  OAI22_X1 U1217 ( .A1(n36), .A2(n741), .B1(n34), .B2(n740), .ZN(n610) );
  INV_X1 U1218 ( .A(n380), .ZN(n381) );
  OAI22_X1 U1219 ( .A1(n24), .A2(n774), .B1(n773), .B2(n22), .ZN(n641) );
  OAI22_X1 U1220 ( .A1(n30), .A2(n764), .B1(n27), .B2(n763), .ZN(n632) );
  OAI22_X1 U1221 ( .A1(n35), .A2(n749), .B1(n34), .B2(n748), .ZN(n618) );
  AND2_X1 U1222 ( .A1(n1016), .A2(n546), .ZN(n605) );
  OAI22_X1 U1223 ( .A1(n29), .A2(n765), .B1(n27), .B2(n764), .ZN(n633) );
  OAI22_X1 U1224 ( .A1(n1013), .A2(n825), .B1(n824), .B2(n4), .ZN(n690) );
  OAI22_X1 U1225 ( .A1(n29), .A2(n766), .B1(n27), .B2(n765), .ZN(n634) );
  OAI22_X1 U1226 ( .A1(n18), .A2(n796), .B1(n795), .B2(n15), .ZN(n662) );
  OAI22_X1 U1227 ( .A1(n826), .A2(n6), .B1(n825), .B2(n4), .ZN(n691) );
  OAI22_X1 U1228 ( .A1(n11), .A2(n812), .B1(n10), .B2(n811), .ZN(n677) );
  OAI22_X1 U1229 ( .A1(n30), .A2(n767), .B1(n27), .B2(n766), .ZN(n635) );
  OAI22_X1 U1230 ( .A1(n17), .A2(n797), .B1(n15), .B2(n796), .ZN(n663) );
  OAI22_X1 U1231 ( .A1(n11), .A2(n816), .B1(n10), .B2(n815), .ZN(n681) );
  AND2_X1 U1232 ( .A1(n1066), .A2(n555), .ZN(n653) );
  OAI22_X1 U1233 ( .A1(n5), .A2(n831), .B1(n830), .B2(n3), .ZN(n696) );
  OAI22_X1 U1234 ( .A1(n47), .A2(n710), .B1(n45), .B2(n709), .ZN(n581) );
  OAI22_X1 U1235 ( .A1(n29), .A2(n755), .B1(n28), .B2(n754), .ZN(n623) );
  INV_X1 U1236 ( .A(n554), .ZN(n638) );
  OAI22_X1 U1237 ( .A1(n23), .A2(n778), .B1(n22), .B2(n777), .ZN(n645) );
  OAI22_X1 U1238 ( .A1(n42), .A2(n721), .B1(n40), .B2(n720), .ZN(n591) );
  INV_X1 U1239 ( .A(n548), .ZN(n606) );
  AOI21_X1 U1240 ( .B1(n36), .B2(n34), .A(n736), .ZN(n548) );
  OAI22_X1 U1241 ( .A1(n11), .A2(n814), .B1(n10), .B2(n813), .ZN(n679) );
  OAI22_X1 U1242 ( .A1(n23), .A2(n784), .B1(n22), .B2(n783), .ZN(n651) );
  AND2_X1 U1243 ( .A1(n1066), .A2(n549), .ZN(n621) );
  OAI22_X1 U1244 ( .A1(n23), .A2(n782), .B1(n22), .B2(n781), .ZN(n649) );
  OAI22_X1 U1245 ( .A1(n5), .A2(n827), .B1(n826), .B2(n4), .ZN(n692) );
  OAI22_X1 U1246 ( .A1(n30), .A2(n762), .B1(n27), .B2(n761), .ZN(n630) );
  OAI22_X1 U1247 ( .A1(n5), .A2(n822), .B1(n821), .B2(n4), .ZN(n687) );
  OAI22_X1 U1248 ( .A1(n12), .A2(n807), .B1(n10), .B2(n806), .ZN(n672) );
  OAI22_X1 U1249 ( .A1(n36), .A2(n738), .B1(n34), .B2(n737), .ZN(n607) );
  OAI22_X1 U1250 ( .A1(n5), .A2(n828), .B1(n827), .B2(n4), .ZN(n693) );
  OAI22_X1 U1251 ( .A1(n11), .A2(n815), .B1(n10), .B2(n814), .ZN(n680) );
  OAI22_X1 U1252 ( .A1(n17), .A2(n800), .B1(n15), .B2(n799), .ZN(n666) );
  OAI22_X1 U1253 ( .A1(n1013), .A2(n830), .B1(n829), .B2(n3), .ZN(n695) );
  OAI22_X1 U1254 ( .A1(n30), .A2(n763), .B1(n27), .B2(n762), .ZN(n631) );
  OAI22_X1 U1255 ( .A1(n12), .A2(n808), .B1(n10), .B2(n807), .ZN(n673) );
  OAI22_X1 U1256 ( .A1(n42), .A2(n733), .B1(n39), .B2(n732), .ZN(n603) );
  OAI22_X1 U1257 ( .A1(n12), .A2(n809), .B1(n10), .B2(n808), .ZN(n674) );
  OAI22_X1 U1258 ( .A1(n23), .A2(n779), .B1(n22), .B2(n778), .ZN(n646) );
  OAI22_X1 U1259 ( .A1(n1013), .A2(n824), .B1(n823), .B2(n4), .ZN(n689) );
  OAI22_X1 U1260 ( .A1(n30), .A2(n757), .B1(n28), .B2(n756), .ZN(n625) );
  OAI22_X1 U1261 ( .A1(n42), .A2(n728), .B1(n39), .B2(n727), .ZN(n598) );
  OAI22_X1 U1262 ( .A1(n47), .A2(n713), .B1(n45), .B2(n712), .ZN(n584) );
  AND2_X1 U1263 ( .A1(n1016), .A2(n543), .ZN(n589) );
  OAI22_X1 U1264 ( .A1(n35), .A2(n748), .B1(n34), .B2(n747), .ZN(n617) );
  OAI22_X1 U1265 ( .A1(n6), .A2(n823), .B1(n822), .B2(n4), .ZN(n688) );
  OAI22_X1 U1266 ( .A1(n17), .A2(n795), .B1(n15), .B2(n794), .ZN(n661) );
  OAI22_X1 U1267 ( .A1(n42), .A2(n724), .B1(n40), .B2(n723), .ZN(n594) );
  OAI22_X1 U1268 ( .A1(n36), .A2(n739), .B1(n34), .B2(n738), .ZN(n608) );
  OAI22_X1 U1269 ( .A1(n48), .A2(n709), .B1(n46), .B2(n708), .ZN(n580) );
  OAI22_X1 U1270 ( .A1(n23), .A2(n780), .B1(n22), .B2(n779), .ZN(n647) );
  OAI22_X1 U1271 ( .A1(n12), .A2(n810), .B1(n10), .B2(n809), .ZN(n675) );
  OAI22_X1 U1272 ( .A1(n35), .A2(n750), .B1(n34), .B2(n749), .ZN(n619) );
  OAI22_X1 U1273 ( .A1(n23), .A2(n781), .B1(n22), .B2(n780), .ZN(n648) );
  OAI22_X1 U1274 ( .A1(n12), .A2(n811), .B1(n10), .B2(n810), .ZN(n676) );
  AND2_X1 U1275 ( .A1(n1016), .A2(n552), .ZN(n637) );
  OAI22_X1 U1276 ( .A1(n17), .A2(n799), .B1(n15), .B2(n798), .ZN(n665) );
  OAI22_X1 U1277 ( .A1(n5), .A2(n829), .B1(n828), .B2(n3), .ZN(n694) );
  INV_X1 U1278 ( .A(n22), .ZN(n555) );
  NAND2_X1 U1279 ( .A1(n539), .A2(n540), .ZN(n291) );
  OAI22_X1 U1280 ( .A1(n23), .A2(n882), .B1(n786), .B2(n22), .ZN(n570) );
  OAI22_X1 U1281 ( .A1(n23), .A2(n785), .B1(n22), .B2(n784), .ZN(n652) );
  OR2_X1 U1282 ( .A1(n1066), .A2(n882), .ZN(n786) );
  OAI22_X1 U1283 ( .A1(n41), .A2(n879), .B1(n735), .B2(n39), .ZN(n567) );
  OAI22_X1 U1284 ( .A1(n734), .A2(n41), .B1(n39), .B2(n733), .ZN(n604) );
  OR2_X1 U1285 ( .A1(n1065), .A2(n879), .ZN(n735) );
  INV_X1 U1286 ( .A(n542), .ZN(n574) );
  AOI21_X1 U1287 ( .B1(n48), .B2(n46), .A(n702), .ZN(n542) );
  OAI22_X1 U1288 ( .A1(n47), .A2(n712), .B1(n45), .B2(n711), .ZN(n583) );
  INV_X1 U1289 ( .A(n557), .ZN(n654) );
  OAI22_X1 U1290 ( .A1(n29), .A2(n761), .B1(n27), .B2(n760), .ZN(n629) );
  OAI22_X1 U1291 ( .A1(n47), .A2(n716), .B1(n45), .B2(n715), .ZN(n587) );
  INV_X1 U1292 ( .A(n563), .ZN(n686) );
  INV_X1 U1293 ( .A(n45), .ZN(n543) );
  INV_X1 U1294 ( .A(n34), .ZN(n549) );
  INV_X1 U1295 ( .A(n15), .ZN(n558) );
  INV_X1 U1296 ( .A(n27), .ZN(n552) );
  INV_X1 U1297 ( .A(n39), .ZN(n546) );
  AND2_X1 U1298 ( .A1(n1066), .A2(n564), .ZN(product[0]) );
  INV_X1 U1299 ( .A(n3), .ZN(n564) );
  XNOR2_X1 U1300 ( .A(n957), .B(n851), .ZN(n749) );
  XNOR2_X1 U1301 ( .A(n25), .B(n851), .ZN(n766) );
  XNOR2_X1 U1302 ( .A(n1057), .B(n851), .ZN(n800) );
  XNOR2_X1 U1303 ( .A(n1), .B(n851), .ZN(n834) );
  XNOR2_X1 U1304 ( .A(n25), .B(n850), .ZN(n765) );
  XNOR2_X1 U1305 ( .A(n957), .B(n850), .ZN(n748) );
  XNOR2_X1 U1306 ( .A(n1057), .B(n979), .ZN(n799) );
  OAI22_X1 U1307 ( .A1(n11), .A2(n819), .B1(n10), .B2(n818), .ZN(n684) );
  OAI22_X1 U1308 ( .A1(n1013), .A2(n834), .B1(n833), .B2(n3), .ZN(n699) );
  OAI22_X1 U1309 ( .A1(n1013), .A2(n836), .B1(n835), .B2(n3), .ZN(n701) );
  XNOR2_X1 U1310 ( .A(n1), .B(n1066), .ZN(n836) );
  XNOR2_X1 U1311 ( .A(n25), .B(n838), .ZN(n753) );
  XNOR2_X1 U1312 ( .A(n957), .B(n1011), .ZN(n736) );
  OAI22_X1 U1313 ( .A1(n1013), .A2(n885), .B1(n837), .B2(n4), .ZN(n573) );
  OR2_X1 U1314 ( .A1(n1016), .A2(n885), .ZN(n837) );
  BUF_X2 U1315 ( .A(n874), .Z(n22) );
  XNOR2_X1 U1316 ( .A(n1058), .B(n852), .ZN(n750) );
  XNOR2_X1 U1317 ( .A(n25), .B(n852), .ZN(n767) );
  XNOR2_X1 U1318 ( .A(n1057), .B(n852), .ZN(n801) );
  XNOR2_X1 U1319 ( .A(n1), .B(n852), .ZN(n835) );
  XNOR2_X1 U1320 ( .A(n957), .B(n842), .ZN(n740) );
  XNOR2_X1 U1321 ( .A(n25), .B(n842), .ZN(n757) );
  XNOR2_X1 U1322 ( .A(n25), .B(n1004), .ZN(n756) );
  XNOR2_X1 U1323 ( .A(n25), .B(n843), .ZN(n758) );
  XNOR2_X1 U1324 ( .A(n25), .B(n1020), .ZN(n755) );
  XNOR2_X1 U1325 ( .A(n25), .B(n839), .ZN(n754) );
  XNOR2_X1 U1326 ( .A(n25), .B(n844), .ZN(n759) );
  XNOR2_X1 U1327 ( .A(n25), .B(n845), .ZN(n760) );
  XNOR2_X1 U1328 ( .A(n25), .B(n846), .ZN(n761) );
  XNOR2_X1 U1329 ( .A(n25), .B(n848), .ZN(n763) );
  XNOR2_X1 U1330 ( .A(n25), .B(n847), .ZN(n762) );
  XNOR2_X1 U1331 ( .A(n25), .B(n849), .ZN(n764) );
  XNOR2_X1 U1332 ( .A(n957), .B(n846), .ZN(n744) );
  XNOR2_X1 U1333 ( .A(n1), .B(n842), .ZN(n825) );
  XNOR2_X1 U1334 ( .A(n1), .B(n839), .ZN(n822) );
  XNOR2_X1 U1335 ( .A(n1), .B(n846), .ZN(n829) );
  XNOR2_X1 U1336 ( .A(n1), .B(n840), .ZN(n823) );
  XNOR2_X1 U1337 ( .A(n1), .B(n841), .ZN(n824) );
  XNOR2_X1 U1338 ( .A(n1), .B(n844), .ZN(n827) );
  XNOR2_X1 U1339 ( .A(n1), .B(n843), .ZN(n826) );
  XNOR2_X1 U1340 ( .A(n1), .B(n961), .ZN(n828) );
  XNOR2_X1 U1341 ( .A(n1), .B(n849), .ZN(n832) );
  XNOR2_X1 U1342 ( .A(n1), .B(n847), .ZN(n830) );
  XNOR2_X1 U1343 ( .A(n1), .B(n848), .ZN(n831) );
  BUF_X2 U1344 ( .A(b[14]), .Z(n839) );
  BUF_X2 U1345 ( .A(n875), .Z(n15) );
  BUF_X2 U1346 ( .A(n871), .Z(n39) );
  BUF_X2 U1347 ( .A(n876), .Z(n10) );
  BUF_X2 U1348 ( .A(n868), .Z(n12) );
  BUF_X2 U1349 ( .A(b[6]), .Z(n847) );
  BUF_X2 U1350 ( .A(n864), .Z(n36) );
  BUF_X2 U1351 ( .A(n862), .Z(n48) );
  XNOR2_X1 U1352 ( .A(n1057), .B(n842), .ZN(n791) );
  XNOR2_X1 U1353 ( .A(n25), .B(n1016), .ZN(n768) );
  BUF_X2 U1354 ( .A(n862), .Z(n47) );
  BUF_X2 U1355 ( .A(n864), .Z(n35) );
  BUF_X1 U1356 ( .A(n868), .Z(n11) );
  BUF_X1 U1357 ( .A(n869), .Z(n5) );
  BUF_X2 U1358 ( .A(n866), .Z(n23) );
  INV_X1 U1359 ( .A(n1058), .ZN(n880) );
  OAI22_X1 U1360 ( .A1(n12), .A2(n884), .B1(n820), .B2(n10), .ZN(n572) );
  OR2_X1 U1361 ( .A1(n1016), .A2(n884), .ZN(n820) );
  INV_X1 U1362 ( .A(n7), .ZN(n884) );
  INV_X1 U1363 ( .A(n37), .ZN(n879) );
  INV_X1 U1364 ( .A(n19), .ZN(n882) );
  INV_X1 U1365 ( .A(n43), .ZN(n878) );
  CLKBUF_X1 U1366 ( .A(b[0]), .Z(n49) );
  INV_X1 U1367 ( .A(n1021), .ZN(n230) );
  NOR2_X1 U1368 ( .A1(n445), .A2(n458), .ZN(n232) );
  XOR2_X1 U1369 ( .A(n80), .B(n292), .Z(product[4]) );
  NOR2_X1 U1370 ( .A1(n218), .A2(n958), .ZN(n209) );
  AOI21_X1 U1371 ( .B1(n1001), .B2(n289), .A(n286), .ZN(n284) );
  XNOR2_X1 U1372 ( .A(n79), .B(n289), .ZN(product[5]) );
  BUF_X1 U1373 ( .A(n871), .Z(n40) );
  XNOR2_X1 U1374 ( .A(a[12]), .B(a[11]), .ZN(n871) );
  NAND2_X1 U1375 ( .A1(n858), .A2(n874), .ZN(n866) );
  XNOR2_X1 U1376 ( .A(a[6]), .B(a[5]), .ZN(n874) );
  XNOR2_X1 U1377 ( .A(n247), .B(n71), .ZN(product[13]) );
  OAI21_X1 U1378 ( .B1(n254), .B2(n252), .A(n249), .ZN(n247) );
  NAND2_X1 U1379 ( .A1(n974), .A2(n416), .ZN(n212) );
  INV_X1 U1380 ( .A(n1), .ZN(n885) );
  INV_X1 U1381 ( .A(n25), .ZN(n881) );
  OAI22_X1 U1382 ( .A1(n30), .A2(n881), .B1(n769), .B2(n28), .ZN(n569) );
  OR2_X1 U1383 ( .A1(n1066), .A2(n881), .ZN(n769) );
  INV_X1 U1384 ( .A(n402), .ZN(n403) );
  XNOR2_X1 U1385 ( .A(n7), .B(n847), .ZN(n813) );
  XNOR2_X1 U1386 ( .A(n7), .B(n846), .ZN(n812) );
  XNOR2_X1 U1387 ( .A(n7), .B(n844), .ZN(n810) );
  XNOR2_X1 U1388 ( .A(n7), .B(n845), .ZN(n811) );
  XNOR2_X1 U1389 ( .A(n7), .B(n979), .ZN(n816) );
  XNOR2_X1 U1390 ( .A(n7), .B(n843), .ZN(n809) );
  XNOR2_X1 U1391 ( .A(n7), .B(n849), .ZN(n815) );
  XNOR2_X1 U1392 ( .A(n7), .B(n842), .ZN(n808) );
  XNOR2_X1 U1393 ( .A(n7), .B(n841), .ZN(n807) );
  XNOR2_X1 U1394 ( .A(n7), .B(n848), .ZN(n814) );
  XNOR2_X1 U1395 ( .A(n7), .B(n851), .ZN(n817) );
  XNOR2_X1 U1396 ( .A(n7), .B(n1066), .ZN(n819) );
  XNOR2_X1 U1397 ( .A(n7), .B(n1020), .ZN(n806) );
  XNOR2_X1 U1398 ( .A(n7), .B(n852), .ZN(n818) );
  XNOR2_X1 U1399 ( .A(n7), .B(n839), .ZN(n805) );
  XNOR2_X1 U1400 ( .A(n7), .B(n838), .ZN(n804) );
  AND2_X1 U1401 ( .A1(n471), .A2(n482), .ZN(n1061) );
  CLKBUF_X1 U1402 ( .A(n956), .Z(n1062) );
  BUF_X2 U1403 ( .A(n867), .Z(n18) );
  NAND2_X1 U1404 ( .A1(n861), .A2(n877), .ZN(n869) );
  AOI21_X1 U1405 ( .B1(n1063), .B2(n264), .A(n259), .ZN(n257) );
  INV_X1 U1406 ( .A(n266), .ZN(n264) );
  INV_X1 U1407 ( .A(n261), .ZN(n259) );
  NAND2_X1 U1408 ( .A1(n519), .A2(n524), .ZN(n275) );
  XNOR2_X1 U1409 ( .A(n19), .B(n848), .ZN(n780) );
  XNOR2_X1 U1410 ( .A(n19), .B(n1066), .ZN(n785) );
  XNOR2_X1 U1411 ( .A(n19), .B(n852), .ZN(n784) );
  XNOR2_X1 U1412 ( .A(n19), .B(n845), .ZN(n777) );
  XNOR2_X1 U1413 ( .A(n19), .B(n844), .ZN(n776) );
  XNOR2_X1 U1414 ( .A(n19), .B(n847), .ZN(n779) );
  XNOR2_X1 U1415 ( .A(n19), .B(n846), .ZN(n778) );
  XNOR2_X1 U1416 ( .A(n19), .B(n851), .ZN(n783) );
  XNOR2_X1 U1417 ( .A(n19), .B(n1003), .ZN(n782) );
  XNOR2_X1 U1418 ( .A(n19), .B(n849), .ZN(n781) );
  XNOR2_X1 U1419 ( .A(n19), .B(n841), .ZN(n773) );
  XNOR2_X1 U1420 ( .A(n19), .B(n843), .ZN(n775) );
  XNOR2_X1 U1421 ( .A(n19), .B(n840), .ZN(n772) );
  XNOR2_X1 U1422 ( .A(n19), .B(n842), .ZN(n774) );
  XNOR2_X1 U1423 ( .A(n19), .B(n839), .ZN(n771) );
  XNOR2_X1 U1424 ( .A(n19), .B(n838), .ZN(n770) );
  AOI21_X1 U1425 ( .B1(n1039), .B2(n1062), .A(n1061), .ZN(n1064) );
  XNOR2_X1 U1426 ( .A(n953), .B(n1004), .ZN(n722) );
  XNOR2_X1 U1427 ( .A(n953), .B(n1020), .ZN(n721) );
  XNOR2_X1 U1428 ( .A(n37), .B(n845), .ZN(n726) );
  XNOR2_X1 U1429 ( .A(n37), .B(n842), .ZN(n723) );
  XNOR2_X1 U1430 ( .A(n37), .B(n851), .ZN(n732) );
  XNOR2_X1 U1431 ( .A(n37), .B(n844), .ZN(n725) );
  XNOR2_X1 U1432 ( .A(n37), .B(n850), .ZN(n731) );
  XNOR2_X1 U1433 ( .A(n37), .B(n843), .ZN(n724) );
  XNOR2_X1 U1434 ( .A(n37), .B(n1065), .ZN(n734) );
  XNOR2_X1 U1435 ( .A(n37), .B(n846), .ZN(n727) );
  XNOR2_X1 U1436 ( .A(n953), .B(n1006), .ZN(n720) );
  XNOR2_X1 U1437 ( .A(n37), .B(n852), .ZN(n733) );
  XNOR2_X1 U1438 ( .A(n37), .B(n847), .ZN(n728) );
  XNOR2_X1 U1439 ( .A(n37), .B(n849), .ZN(n730) );
  XNOR2_X1 U1440 ( .A(n953), .B(n1011), .ZN(n719) );
  XNOR2_X1 U1441 ( .A(n37), .B(n848), .ZN(n729) );
  XNOR2_X1 U1442 ( .A(a[13]), .B(a[14]), .ZN(n870) );
  OAI21_X1 U1443 ( .B1(n199), .B2(n205), .A(n200), .ZN(n198) );
  NAND2_X1 U1444 ( .A1(n383), .A2(n392), .ZN(n200) );
  INV_X1 U1445 ( .A(n1062), .ZN(n249) );
  AOI21_X1 U1446 ( .B1(n1039), .B2(n956), .A(n1061), .ZN(n242) );
  NOR2_X1 U1447 ( .A1(n531), .A2(n534), .ZN(n282) );
  NAND2_X1 U1448 ( .A1(n531), .A2(n534), .ZN(n283) );
  INV_X1 U1449 ( .A(n282), .ZN(n326) );
  NAND2_X1 U1450 ( .A1(n1039), .A2(n250), .ZN(n241) );
  INV_X1 U1451 ( .A(n252), .ZN(n250) );
  OAI22_X1 U1452 ( .A1(n17), .A2(n793), .B1(n15), .B2(n792), .ZN(n659) );
  OAI22_X1 U1453 ( .A1(n17), .A2(n1050), .B1(n803), .B2(n15), .ZN(n571) );
  OAI22_X1 U1454 ( .A1(n18), .A2(n794), .B1(n15), .B2(n793), .ZN(n660) );
  OAI22_X1 U1455 ( .A1(n17), .A2(n792), .B1(n15), .B2(n791), .ZN(n658) );
  OAI22_X1 U1456 ( .A1(n18), .A2(n791), .B1(n790), .B2(n15), .ZN(n657) );
  AOI21_X1 U1457 ( .B1(n17), .B2(n15), .A(n787), .ZN(n557) );
  OAI22_X1 U1458 ( .A1(n17), .A2(n790), .B1(n15), .B2(n789), .ZN(n656) );
  OAI22_X1 U1459 ( .A1(n18), .A2(n789), .B1(n788), .B2(n15), .ZN(n655) );
  OAI22_X1 U1460 ( .A1(n18), .A2(n788), .B1(n15), .B2(n787), .ZN(n402) );
  NAND2_X1 U1461 ( .A1(n859), .A2(n875), .ZN(n867) );
  XNOR2_X1 U1462 ( .A(n955), .B(n1004), .ZN(n705) );
  XNOR2_X1 U1463 ( .A(n955), .B(n1019), .ZN(n704) );
  XNOR2_X1 U1464 ( .A(n955), .B(n1006), .ZN(n703) );
  XNOR2_X1 U1465 ( .A(n43), .B(n1005), .ZN(n707) );
  XNOR2_X1 U1466 ( .A(n955), .B(n1011), .ZN(n702) );
  XNOR2_X1 U1467 ( .A(n43), .B(n842), .ZN(n706) );
  XNOR2_X1 U1468 ( .A(n43), .B(n844), .ZN(n708) );
  XNOR2_X1 U1469 ( .A(n43), .B(n1016), .ZN(n717) );
  XNOR2_X1 U1470 ( .A(n43), .B(n846), .ZN(n710) );
  XNOR2_X1 U1471 ( .A(n43), .B(n845), .ZN(n709) );
  XNOR2_X1 U1472 ( .A(n43), .B(n847), .ZN(n711) );
  XNOR2_X1 U1473 ( .A(n43), .B(n852), .ZN(n716) );
  XNOR2_X1 U1474 ( .A(n43), .B(n848), .ZN(n712) );
  XNOR2_X1 U1475 ( .A(n43), .B(n851), .ZN(n715) );
  XNOR2_X1 U1476 ( .A(n43), .B(n850), .ZN(n714) );
  XNOR2_X1 U1477 ( .A(n43), .B(n849), .ZN(n713) );
  OAI21_X1 U1478 ( .B1(n254), .B2(n241), .A(n1064), .ZN(n240) );
  XOR2_X1 U1479 ( .A(n82), .B(n301), .Z(product[2]) );
  OAI21_X1 U1480 ( .B1(n298), .B2(n301), .A(n299), .ZN(n297) );
  NAND2_X1 U1481 ( .A1(n701), .A2(n573), .ZN(n301) );
  INV_X1 U1482 ( .A(n959), .ZN(n221) );
  BUF_X2 U1483 ( .A(n865), .Z(n30) );
  NAND2_X1 U1484 ( .A1(n857), .A2(n873), .ZN(n865) );
  NAND2_X1 U1485 ( .A1(n856), .A2(n872), .ZN(n864) );
  NAND2_X1 U1486 ( .A1(n445), .A2(n458), .ZN(n233) );
  AOI21_X1 U1487 ( .B1(n155), .B2(n180), .A(n156), .ZN(n154) );
  XNOR2_X1 U1488 ( .A(a[4]), .B(a[3]), .ZN(n875) );
  NAND2_X1 U1489 ( .A1(n320), .A2(n253), .ZN(n72) );
  OAI22_X1 U1490 ( .A1(n48), .A2(n878), .B1(n718), .B2(n46), .ZN(n566) );
  OAI21_X1 U1491 ( .B1(n150), .B2(n144), .A(n145), .ZN(n141) );
  OAI22_X1 U1492 ( .A1(n41), .A2(n729), .B1(n39), .B2(n728), .ZN(n599) );
  OAI21_X1 U1493 ( .B1(n282), .B2(n284), .A(n283), .ZN(n281) );
  INV_X1 U1494 ( .A(n288), .ZN(n286) );
  AOI21_X1 U1495 ( .B1(n980), .B2(n226), .A(n210), .ZN(n208) );
  OAI21_X1 U1496 ( .B1(n211), .B2(n219), .A(n212), .ZN(n210) );
  OAI22_X1 U1497 ( .A1(n36), .A2(n880), .B1(n752), .B2(n34), .ZN(n568) );
  OR2_X1 U1498 ( .A1(n1065), .A2(n880), .ZN(n752) );
  NAND2_X1 U1499 ( .A1(n860), .A2(n876), .ZN(n868) );
  OAI21_X1 U1500 ( .B1(n290), .B2(n292), .A(n291), .ZN(n289) );
  XNOR2_X1 U1501 ( .A(n1057), .B(n839), .ZN(n788) );
  XNOR2_X1 U1502 ( .A(n1057), .B(n846), .ZN(n795) );
  XNOR2_X1 U1503 ( .A(n1057), .B(n847), .ZN(n796) );
  XNOR2_X1 U1504 ( .A(n1057), .B(n1019), .ZN(n789) );
  XNOR2_X1 U1505 ( .A(n1057), .B(n841), .ZN(n790) );
  INV_X1 U1506 ( .A(n1034), .ZN(n316) );
  NAND2_X1 U1507 ( .A1(n431), .A2(n444), .ZN(n228) );
  INV_X1 U1508 ( .A(n252), .ZN(n320) );
  NOR2_X1 U1509 ( .A1(n483), .A2(n492), .ZN(n252) );
  XNOR2_X1 U1510 ( .A(a[2]), .B(a[1]), .ZN(n876) );
  XNOR2_X1 U1511 ( .A(n1), .B(n838), .ZN(n821) );
  XNOR2_X1 U1512 ( .A(n1), .B(n850), .ZN(n833) );
  AOI21_X1 U1513 ( .B1(n236), .B2(n255), .A(n237), .ZN(n235) );
  INV_X1 U1514 ( .A(n1025), .ZN(n254) );
  OAI21_X1 U1515 ( .B1(n256), .B2(n268), .A(n257), .ZN(n255) );
  INV_X1 U1516 ( .A(n1049), .ZN(n234) );
  OAI21_X1 U1517 ( .B1(n150), .B2(n109), .A(n110), .ZN(n108) );
  OAI21_X1 U1518 ( .B1(n145), .B2(n137), .A(n138), .ZN(n136) );
  AOI21_X1 U1519 ( .B1(n214), .B2(n234), .A(n215), .ZN(n213) );
  AOI21_X1 U1520 ( .B1(n234), .B2(n230), .A(n231), .ZN(n229) );
  AOI21_X1 U1521 ( .B1(n234), .B2(n221), .A(n1022), .ZN(n220) );
  OAI21_X1 U1522 ( .B1(n153), .B2(n191), .A(n154), .ZN(n152) );
  NAND2_X1 U1523 ( .A1(n854), .A2(n870), .ZN(n862) );
  NOR2_X1 U1524 ( .A1(n417), .A2(n430), .ZN(n218) );
  INV_X1 U1525 ( .A(n1032), .ZN(n217) );
  NAND2_X1 U1526 ( .A1(n365), .A2(n372), .ZN(n182) );
  NAND2_X1 U1527 ( .A1(n855), .A2(n871), .ZN(n863) );
  NOR2_X1 U1528 ( .A1(n168), .A2(n157), .ZN(n155) );
  OAI21_X1 U1529 ( .B1(n157), .B2(n169), .A(n158), .ZN(n156) );
  AOI21_X1 U1530 ( .B1(n1059), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U1531 ( .B1(n1014), .B2(n94), .A(n95), .ZN(n93) );
  XNOR2_X1 U1532 ( .A(n1015), .B(n65), .ZN(product[19]) );
  AOI21_X1 U1533 ( .B1(n1060), .B2(n131), .A(n132), .ZN(n130) );
  AOI21_X1 U1534 ( .B1(n1059), .B2(n118), .A(n119), .ZN(n117) );
  AOI21_X1 U1535 ( .B1(n1014), .B2(n147), .A(n148), .ZN(n146) );
  AOI21_X1 U1536 ( .B1(n206), .B2(n184), .A(n185), .ZN(n183) );
  AOI21_X1 U1537 ( .B1(n206), .B2(n313), .A(n203), .ZN(n201) );
  AOI21_X1 U1538 ( .B1(n1014), .B2(n160), .A(n161), .ZN(n159) );
  AOI21_X1 U1539 ( .B1(n193), .B2(n206), .A(n1012), .ZN(n192) );
  AOI21_X1 U1540 ( .B1(n1060), .B2(n140), .A(n141), .ZN(n139) );
  AOI21_X1 U1541 ( .B1(n171), .B2(n206), .A(n172), .ZN(n170) );
  AOI21_X1 U1542 ( .B1(n1015), .B2(n107), .A(n108), .ZN(n106) );
  XOR2_X1 U1543 ( .A(a[14]), .B(a[15]), .Z(n854) );
  NOR2_X1 U1544 ( .A1(n972), .A2(n109), .ZN(n107) );
  NOR2_X1 U1545 ( .A1(n190), .A2(n153), .ZN(n151) );
  XNOR2_X1 U1546 ( .A(n234), .B(n69), .ZN(product[15]) );
  NAND2_X1 U1547 ( .A1(n230), .A2(n233), .ZN(n69) );
  OAI21_X1 U1548 ( .B1(n1048), .B2(n207), .A(n208), .ZN(n206) );
  NAND2_X1 U1549 ( .A1(n209), .A2(n225), .ZN(n207) );
  NOR2_X1 U1550 ( .A1(n227), .A2(n232), .ZN(n225) );
  BUF_X4 U1551 ( .A(a[7]), .Z(n19) );
  XOR2_X1 U1552 ( .A(a[6]), .B(a[7]), .Z(n858) );
  XNOR2_X1 U1553 ( .A(a[7]), .B(a[8]), .ZN(n873) );
  BUF_X4 U1554 ( .A(a[3]), .Z(n7) );
  XOR2_X1 U1555 ( .A(a[2]), .B(a[3]), .Z(n860) );
  INV_X1 U1556 ( .A(n268), .ZN(n267) );
  XOR2_X1 U1557 ( .A(a[12]), .B(a[13]), .Z(n855) );
  OAI21_X1 U1558 ( .B1(n242), .B2(n238), .A(n239), .ZN(n237) );
  BUF_X4 U1559 ( .A(a[9]), .Z(n25) );
  XOR2_X1 U1560 ( .A(a[8]), .B(a[9]), .Z(n857) );
  XNOR2_X1 U1561 ( .A(a[10]), .B(a[9]), .ZN(n872) );
  XNOR2_X1 U1562 ( .A(n1037), .B(n75), .ZN(product[9]) );
  NAND2_X1 U1563 ( .A1(n155), .A2(n1045), .ZN(n153) );
  XOR2_X1 U1564 ( .A(a[10]), .B(a[11]), .Z(n856) );
  XOR2_X1 U1565 ( .A(n1018), .B(n76), .Z(product[8]) );
  NAND2_X1 U1566 ( .A1(n541), .A2(n572), .ZN(n296) );
  XNOR2_X1 U1567 ( .A(n281), .B(n77), .ZN(product[7]) );
  AOI21_X1 U1568 ( .B1(n281), .B2(n1000), .A(n278), .ZN(n276) );
  BUF_X4 U1569 ( .A(a[1]), .Z(n1) );
  XOR2_X1 U1570 ( .A(a[0]), .B(a[1]), .Z(n861) );
  XOR2_X1 U1571 ( .A(n78), .B(n1023), .Z(product[6]) );
endmodule


module datapath_DW_mult_tc_15 ( a, b, product );
  input [15:0] a;
  input [15:0] b;
  output [31:0] product;
  wire   n1, n3, n5, n6, n7, n9, n10, n11, n12, n13, n15, n16, n17, n18, n19,
         n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34, n35, n36,
         n37, n39, n40, n41, n42, n43, n45, n46, n47, n48, n49, n51, n54, n65,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n84, n85, n86, n87, n88, n90, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n103, n105, n106, n107, n108, n109, n110, n114, n116,
         n117, n118, n119, n122, n123, n124, n125, n127, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n143,
         n144, n145, n146, n147, n148, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n180, n182, n183, n184, n185, n188, n189, n190, n191, n192,
         n194, n195, n196, n197, n198, n199, n200, n201, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n217,
         n218, n219, n220, n224, n225, n226, n227, n228, n229, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n246,
         n247, n251, n252, n253, n254, n255, n256, n257, n259, n261, n262,
         n264, n266, n267, n268, n270, n272, n273, n274, n275, n276, n278,
         n280, n281, n282, n283, n284, n286, n288, n289, n290, n291, n292,
         n294, n296, n297, n298, n299, n301, n306, n308, n312, n313, n314,
         n316, n317, n318, n320, n324, n326, n328, n330, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n545,
         n546, n548, n549, n551, n552, n554, n555, n557, n558, n560, n561,
         n563, n564, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1032, n1033;
  assign product[31] = n84;

  FA_X1 U364 ( .A(n575), .B(n338), .CI(n590), .CO(n334), .S(n335) );
  FA_X1 U365 ( .A(n339), .B(n576), .CI(n342), .CO(n336), .S(n337) );
  FA_X1 U367 ( .A(n346), .B(n577), .CI(n343), .CO(n340), .S(n341) );
  FA_X1 U368 ( .A(n591), .B(n348), .CI(n606), .CO(n342), .S(n343) );
  FA_X1 U369 ( .A(n347), .B(n354), .CI(n352), .CO(n344), .S(n345) );
  FA_X1 U370 ( .A(n578), .B(n592), .CI(n349), .CO(n346), .S(n347) );
  FA_X1 U372 ( .A(n358), .B(n355), .CI(n353), .CO(n350), .S(n351) );
  FA_X1 U373 ( .A(n362), .B(n607), .CI(n360), .CO(n352), .S(n353) );
  FA_X1 U374 ( .A(n593), .B(n579), .CI(n622), .CO(n354), .S(n355) );
  FA_X1 U375 ( .A(n359), .B(n361), .CI(n366), .CO(n356), .S(n357) );
  FA_X1 U376 ( .A(n370), .B(n363), .CI(n368), .CO(n358), .S(n359) );
  FA_X1 U377 ( .A(n580), .B(n594), .CI(n608), .CO(n360), .S(n361) );
  FA_X1 U379 ( .A(n374), .B(n376), .CI(n367), .CO(n364), .S(n365) );
  FA_X1 U380 ( .A(n369), .B(n378), .CI(n371), .CO(n366), .S(n367) );
  FA_X1 U381 ( .A(n595), .B(n380), .CI(n609), .CO(n368), .S(n369) );
  FA_X1 U382 ( .A(n623), .B(n581), .CI(n638), .CO(n370), .S(n371) );
  FA_X1 U383 ( .A(n384), .B(n377), .CI(n375), .CO(n372), .S(n373) );
  FA_X1 U384 ( .A(n379), .B(n388), .CI(n386), .CO(n374), .S(n375) );
  FA_X1 U385 ( .A(n381), .B(n610), .CI(n390), .CO(n376), .S(n377) );
  FA_X1 U386 ( .A(n624), .B(n596), .CI(n582), .CO(n378), .S(n379) );
  FA_X1 U388 ( .A(n394), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FA_X1 U389 ( .A(n391), .B(n389), .CI(n396), .CO(n384), .S(n385) );
  FA_X1 U390 ( .A(n400), .B(n625), .CI(n398), .CO(n386), .S(n387) );
  FA_X1 U391 ( .A(n597), .B(n639), .CI(n611), .CO(n388), .S(n389) );
  FA_X1 U392 ( .A(n1004), .B(n583), .CI(n654), .CO(n390), .S(n391) );
  FA_X1 U393 ( .A(n406), .B(n397), .CI(n395), .CO(n392), .S(n393) );
  FA_X1 U394 ( .A(n410), .B(n399), .CI(n408), .CO(n394), .S(n395) );
  FA_X1 U395 ( .A(n412), .B(n414), .CI(n401), .CO(n396), .S(n397) );
  FA_X1 U396 ( .A(n584), .B(n598), .CI(n403), .CO(n398), .S(n399) );
  FA_X1 U397 ( .A(n612), .B(n626), .CI(n640), .CO(n400), .S(n401) );
  FA_X1 U399 ( .A(n418), .B(n409), .CI(n407), .CO(n404), .S(n405) );
  FA_X1 U400 ( .A(n411), .B(n422), .CI(n420), .CO(n406), .S(n407) );
  FA_X1 U401 ( .A(n413), .B(n424), .CI(n415), .CO(n408), .S(n409) );
  FA_X1 U402 ( .A(n613), .B(n627), .CI(n426), .CO(n410), .S(n411) );
  FA_X1 U403 ( .A(n599), .B(n655), .CI(n641), .CO(n412), .S(n413) );
  FA_X1 U404 ( .A(n428), .B(n585), .CI(n670), .CO(n414), .S(n415) );
  FA_X1 U405 ( .A(n432), .B(n421), .CI(n419), .CO(n416), .S(n417) );
  FA_X1 U406 ( .A(n423), .B(n436), .CI(n434), .CO(n418), .S(n419) );
  FA_X1 U407 ( .A(n427), .B(n438), .CI(n425), .CO(n420), .S(n421) );
  FA_X1 U408 ( .A(n442), .B(n429), .CI(n440), .CO(n422), .S(n423) );
  FA_X1 U409 ( .A(n642), .B(n628), .CI(n600), .CO(n424), .S(n425) );
  FA_X1 U410 ( .A(n586), .B(n614), .CI(n656), .CO(n426), .S(n427) );
  FA_X1 U413 ( .A(n437), .B(n450), .CI(n448), .CO(n432), .S(n433) );
  FA_X1 U414 ( .A(n439), .B(n452), .CI(n441), .CO(n434), .S(n435) );
  FA_X1 U415 ( .A(n443), .B(n456), .CI(n454), .CO(n436), .S(n437) );
  FA_X1 U416 ( .A(n671), .B(n615), .CI(n657), .CO(n438), .S(n439) );
  FA_X1 U417 ( .A(n629), .B(n587), .CI(n686), .CO(n440), .S(n441) );
  FA_X1 U420 ( .A(n449), .B(n460), .CI(n447), .CO(n444), .S(n445) );
  FA_X1 U421 ( .A(n455), .B(n462), .CI(n451), .CO(n446), .S(n447) );
  FA_X1 U422 ( .A(n464), .B(n466), .CI(n453), .CO(n448), .S(n449) );
  FA_X1 U423 ( .A(n457), .B(n672), .CI(n468), .CO(n450), .S(n451) );
  FA_X1 U424 ( .A(n687), .B(n630), .CI(n658), .CO(n452), .S(n453) );
  FA_X1 U425 ( .A(n602), .B(n644), .CI(n616), .CO(n454), .S(n455) );
  HA_X1 U426 ( .A(n566), .B(n588), .CO(n456), .S(n457) );
  FA_X1 U428 ( .A(n465), .B(n467), .CI(n474), .CO(n460), .S(n461) );
  FA_X1 U429 ( .A(n476), .B(n478), .CI(n469), .CO(n462), .S(n463) );
  FA_X1 U430 ( .A(n645), .B(n659), .CI(n480), .CO(n464), .S(n465) );
  FA_X1 U431 ( .A(n603), .B(n673), .CI(n631), .CO(n466), .S(n467) );
  FA_X1 U432 ( .A(n688), .B(n589), .CI(n617), .CO(n468), .S(n469) );
  FA_X1 U434 ( .A(n479), .B(n477), .CI(n486), .CO(n472), .S(n473) );
  FA_X1 U435 ( .A(n490), .B(n481), .CI(n488), .CO(n474), .S(n475) );
  FA_X1 U436 ( .A(n618), .B(n632), .CI(n660), .CO(n476), .S(n477) );
  FA_X1 U437 ( .A(n689), .B(n646), .CI(n674), .CO(n478), .S(n479) );
  HA_X1 U438 ( .A(n604), .B(n567), .CO(n480), .S(n481) );
  FA_X1 U441 ( .A(n976), .B(n661), .CI(n498), .CO(n486), .S(n487) );
  FA_X1 U442 ( .A(n619), .B(n675), .CI(n647), .CO(n488), .S(n489) );
  FA_X1 U443 ( .A(n633), .B(n605), .CI(n690), .CO(n490), .S(n491) );
  FA_X1 U444 ( .A(n504), .B(n497), .CI(n495), .CO(n492), .S(n493) );
  FA_X1 U445 ( .A(n506), .B(n508), .CI(n499), .CO(n494), .S(n495) );
  FA_X1 U446 ( .A(n648), .B(n676), .CI(n501), .CO(n496), .S(n497) );
  FA_X1 U447 ( .A(n691), .B(n634), .CI(n662), .CO(n498), .S(n499) );
  FA_X1 U449 ( .A(n512), .B(n507), .CI(n505), .CO(n502), .S(n503) );
  FA_X1 U450 ( .A(n514), .B(n516), .CI(n509), .CO(n504), .S(n505) );
  FA_X1 U451 ( .A(n635), .B(n677), .CI(n663), .CO(n506), .S(n507) );
  FA_X1 U452 ( .A(n649), .B(n621), .CI(n692), .CO(n508), .S(n509) );
  FA_X1 U453 ( .A(n515), .B(n520), .CI(n513), .CO(n510), .S(n511) );
  FA_X1 U454 ( .A(n517), .B(n693), .CI(n522), .CO(n512), .S(n513) );
  FA_X1 U455 ( .A(n650), .B(n664), .CI(n678), .CO(n514), .S(n515) );
  HA_X1 U456 ( .A(n569), .B(n636), .CO(n516), .S(n517) );
  FA_X1 U457 ( .A(n523), .B(n526), .CI(n521), .CO(n518), .S(n519) );
  FA_X1 U458 ( .A(n651), .B(n679), .CI(n528), .CO(n520), .S(n521) );
  FA_X1 U459 ( .A(n665), .B(n637), .CI(n694), .CO(n522), .S(n523) );
  FA_X1 U460 ( .A(n532), .B(n529), .CI(n527), .CO(n524), .S(n525) );
  FA_X1 U461 ( .A(n666), .B(n695), .CI(n680), .CO(n526), .S(n527) );
  HA_X1 U462 ( .A(n570), .B(n652), .CO(n528), .S(n529) );
  FA_X1 U463 ( .A(n536), .B(n667), .CI(n533), .CO(n530), .S(n531) );
  FA_X1 U464 ( .A(n696), .B(n653), .CI(n681), .CO(n532), .S(n533) );
  FA_X1 U465 ( .A(n682), .B(n697), .CI(n537), .CO(n534), .S(n535) );
  HA_X1 U466 ( .A(n668), .B(n571), .CO(n536), .S(n537) );
  FA_X1 U467 ( .A(n698), .B(n669), .CI(n683), .CO(n538), .S(n539) );
  HA_X1 U468 ( .A(n684), .B(n699), .CO(n540), .S(n541) );
  CLKBUF_X1 U822 ( .A(n850), .Z(n959) );
  BUF_X2 U823 ( .A(b[7]), .Z(n846) );
  CLKBUF_X3 U824 ( .A(b[4]), .Z(n849) );
  BUF_X4 U825 ( .A(a[1]), .Z(n1) );
  OR2_X2 U826 ( .A1(n471), .A2(n482), .ZN(n1028) );
  BUF_X2 U827 ( .A(n868), .Z(n12) );
  NOR2_X2 U828 ( .A1(n383), .A2(n392), .ZN(n199) );
  XNOR2_X1 U829 ( .A(n473), .B(n953), .ZN(n471) );
  XNOR2_X1 U830 ( .A(n484), .B(n475), .ZN(n953) );
  BUF_X2 U831 ( .A(n866), .Z(n23) );
  CLKBUF_X1 U832 ( .A(n845), .Z(n954) );
  BUF_X2 U833 ( .A(n864), .Z(n36) );
  CLKBUF_X1 U834 ( .A(n226), .Z(n955) );
  CLKBUF_X3 U835 ( .A(b[2]), .Z(n851) );
  XNOR2_X1 U836 ( .A(n433), .B(n956), .ZN(n431) );
  XNOR2_X1 U837 ( .A(n446), .B(n435), .ZN(n956) );
  BUF_X2 U838 ( .A(n877), .Z(n3) );
  CLKBUF_X3 U839 ( .A(b[11]), .Z(n842) );
  CLKBUF_X3 U840 ( .A(b[13]), .Z(n840) );
  NAND2_X1 U841 ( .A1(n198), .A2(n151), .ZN(n957) );
  INV_X1 U842 ( .A(n152), .ZN(n958) );
  AND2_X2 U843 ( .A1(n957), .A2(n958), .ZN(n150) );
  BUF_X2 U844 ( .A(n850), .Z(n960) );
  BUF_X1 U845 ( .A(b[3]), .Z(n850) );
  BUF_X2 U846 ( .A(b[15]), .Z(n838) );
  BUF_X2 U847 ( .A(b[8]), .Z(n845) );
  BUF_X2 U848 ( .A(b[10]), .Z(n843) );
  CLKBUF_X1 U849 ( .A(n218), .Z(n961) );
  XOR2_X1 U850 ( .A(n472), .B(n463), .Z(n962) );
  XOR2_X1 U851 ( .A(n461), .B(n962), .Z(n459) );
  NAND2_X1 U852 ( .A1(n461), .A2(n472), .ZN(n963) );
  NAND2_X1 U853 ( .A1(n461), .A2(n463), .ZN(n964) );
  NAND2_X1 U854 ( .A1(n472), .A2(n463), .ZN(n965) );
  NAND3_X1 U855 ( .A1(n963), .A2(n964), .A3(n965), .ZN(n458) );
  CLKBUF_X1 U856 ( .A(b[0]), .Z(n49) );
  BUF_X1 U857 ( .A(b[9]), .Z(n844) );
  OR2_X1 U858 ( .A1(n503), .A2(n510), .ZN(n966) );
  OR2_X1 U859 ( .A1(n337), .A2(n340), .ZN(n967) );
  OR2_X1 U860 ( .A1(n334), .A2(n333), .ZN(n968) );
  OR2_X1 U861 ( .A1(n574), .A2(n332), .ZN(n969) );
  OR2_X1 U862 ( .A1(n493), .A2(n502), .ZN(n970) );
  OR2_X1 U863 ( .A1(n541), .A2(n572), .ZN(n971) );
  OR2_X1 U864 ( .A1(n336), .A2(n335), .ZN(n972) );
  OR2_X1 U865 ( .A1(n511), .A2(n518), .ZN(n973) );
  OR2_X1 U866 ( .A1(n525), .A2(n530), .ZN(n974) );
  OR2_X1 U867 ( .A1(n535), .A2(n538), .ZN(n975) );
  AND2_X1 U868 ( .A1(n568), .A2(n620), .ZN(n976) );
  OR2_X1 U869 ( .A1(n701), .A2(n573), .ZN(n977) );
  CLKBUF_X2 U870 ( .A(n862), .Z(n48) );
  OAI22_X1 U871 ( .A1(n48), .A2(n703), .B1(n45), .B2(n702), .ZN(n332) );
  CLKBUF_X2 U872 ( .A(b[1]), .Z(n852) );
  CLKBUF_X1 U873 ( .A(n1005), .Z(n978) );
  BUF_X1 U874 ( .A(n235), .Z(n1001) );
  XOR2_X1 U875 ( .A(n620), .B(n568), .Z(n501) );
  BUF_X2 U876 ( .A(b[9]), .Z(n979) );
  XNOR2_X1 U877 ( .A(n159), .B(n980), .ZN(product[24]) );
  AND2_X1 U878 ( .A1(n308), .A2(n158), .ZN(n980) );
  XNOR2_X1 U879 ( .A(n106), .B(n981), .ZN(product[29]) );
  AND2_X1 U880 ( .A1(n968), .A2(n105), .ZN(n981) );
  XNOR2_X1 U881 ( .A(n183), .B(n982), .ZN(product[22]) );
  AND2_X1 U882 ( .A1(n175), .A2(n182), .ZN(n982) );
  XNOR2_X1 U883 ( .A(n117), .B(n983), .ZN(product[28]) );
  AND2_X1 U884 ( .A1(n972), .A2(n116), .ZN(n983) );
  CLKBUF_X1 U885 ( .A(n211), .Z(n984) );
  NAND2_X1 U886 ( .A1(n473), .A2(n484), .ZN(n985) );
  NAND2_X1 U887 ( .A1(n473), .A2(n475), .ZN(n986) );
  NAND2_X1 U888 ( .A1(n484), .A2(n475), .ZN(n987) );
  NAND3_X1 U889 ( .A1(n985), .A2(n986), .A3(n987), .ZN(n470) );
  CLKBUF_X3 U890 ( .A(n865), .Z(n29) );
  CLKBUF_X3 U891 ( .A(n870), .Z(n45) );
  CLKBUF_X3 U892 ( .A(n864), .Z(n35) );
  BUF_X2 U893 ( .A(b[12]), .Z(n841) );
  BUF_X2 U894 ( .A(n862), .Z(n47) );
  BUF_X4 U895 ( .A(a[15]), .Z(n43) );
  XNOR2_X1 U896 ( .A(n146), .B(n988), .ZN(product[25]) );
  AND2_X1 U897 ( .A1(n143), .A2(n145), .ZN(n988) );
  XNOR2_X1 U898 ( .A(n213), .B(n989), .ZN(product[18]) );
  AND2_X1 U899 ( .A1(n314), .A2(n212), .ZN(n989) );
  BUF_X2 U900 ( .A(n866), .Z(n24) );
  XNOR2_X1 U901 ( .A(n25), .B(n960), .ZN(n990) );
  BUF_X2 U902 ( .A(n871), .Z(n39) );
  BUF_X1 U903 ( .A(n869), .Z(n991) );
  BUF_X1 U904 ( .A(n864), .Z(n992) );
  OR2_X1 U905 ( .A1(n365), .A2(n372), .ZN(n993) );
  XNOR2_X1 U906 ( .A(n139), .B(n994), .ZN(product[26]) );
  AND2_X1 U907 ( .A1(n306), .A2(n138), .ZN(n994) );
  BUF_X2 U908 ( .A(a[11]), .Z(n995) );
  BUF_X2 U909 ( .A(n49), .Z(n1032) );
  BUF_X2 U910 ( .A(n49), .Z(n1033) );
  CLKBUF_X1 U911 ( .A(n839), .Z(n996) );
  BUF_X2 U912 ( .A(n865), .Z(n30) );
  XNOR2_X1 U913 ( .A(n229), .B(n997), .ZN(product[16]) );
  AND2_X1 U914 ( .A1(n316), .A2(n228), .ZN(n997) );
  XNOR2_X1 U915 ( .A(n220), .B(n998), .ZN(product[17]) );
  AND2_X1 U916 ( .A1(n217), .A2(n219), .ZN(n998) );
  XNOR2_X1 U917 ( .A(n201), .B(n999), .ZN(product[20]) );
  AND2_X1 U918 ( .A1(n312), .A2(n200), .ZN(n999) );
  XNOR2_X1 U919 ( .A(n130), .B(n1000), .ZN(product[27]) );
  AND2_X1 U920 ( .A1(n967), .A2(n129), .ZN(n1000) );
  BUF_X1 U921 ( .A(n863), .Z(n1002) );
  CLKBUF_X1 U922 ( .A(n242), .Z(n1003) );
  BUF_X1 U923 ( .A(n402), .Z(n1004) );
  BUF_X2 U924 ( .A(n206), .Z(n1005) );
  NOR2_X1 U925 ( .A1(n405), .A2(n416), .ZN(n1006) );
  XNOR2_X1 U926 ( .A(n170), .B(n1007), .ZN(product[23]) );
  AND2_X1 U927 ( .A1(n167), .A2(n169), .ZN(n1007) );
  XNOR2_X1 U928 ( .A(n192), .B(n1008), .ZN(product[21]) );
  AND2_X1 U929 ( .A1(n188), .A2(n191), .ZN(n1008) );
  NOR2_X2 U930 ( .A1(n459), .A2(n470), .ZN(n238) );
  INV_X1 U931 ( .A(n1018), .ZN(n246) );
  AND2_X1 U932 ( .A1(n471), .A2(n482), .ZN(n1018) );
  CLKBUF_X1 U933 ( .A(n276), .Z(n1009) );
  CLKBUF_X1 U934 ( .A(n284), .Z(n1010) );
  NAND2_X1 U935 ( .A1(n433), .A2(n446), .ZN(n1011) );
  NAND2_X1 U936 ( .A1(n433), .A2(n435), .ZN(n1012) );
  NAND2_X1 U937 ( .A1(n446), .A2(n435), .ZN(n1013) );
  NAND3_X1 U938 ( .A1(n1011), .A2(n1012), .A3(n1013), .ZN(n430) );
  NAND2_X1 U939 ( .A1(n37), .A2(n1032), .ZN(n1015) );
  NAND2_X1 U940 ( .A1(n879), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U941 ( .A1(n1015), .A2(n1016), .ZN(n734) );
  INV_X1 U942 ( .A(n1032), .ZN(n1014) );
  BUF_X4 U943 ( .A(a[13]), .Z(n37) );
  OR2_X1 U944 ( .A1(n227), .A2(n232), .ZN(n1017) );
  XOR2_X1 U945 ( .A(n489), .B(n491), .Z(n1019) );
  XOR2_X1 U946 ( .A(n1019), .B(n496), .Z(n485) );
  XOR2_X1 U947 ( .A(n487), .B(n494), .Z(n1020) );
  XOR2_X1 U948 ( .A(n1020), .B(n485), .Z(n483) );
  NAND2_X1 U949 ( .A1(n489), .A2(n491), .ZN(n1021) );
  NAND2_X1 U950 ( .A1(n489), .A2(n496), .ZN(n1022) );
  NAND2_X1 U951 ( .A1(n491), .A2(n496), .ZN(n1023) );
  NAND3_X1 U952 ( .A1(n1021), .A2(n1022), .A3(n1023), .ZN(n484) );
  NAND2_X1 U953 ( .A1(n487), .A2(n494), .ZN(n1024) );
  NAND2_X1 U954 ( .A1(n487), .A2(n485), .ZN(n1025) );
  NAND2_X1 U955 ( .A1(n494), .A2(n485), .ZN(n1026) );
  NAND3_X1 U956 ( .A1(n1024), .A2(n1025), .A3(n1026), .ZN(n482) );
  BUF_X2 U957 ( .A(b[14]), .Z(n839) );
  BUF_X2 U958 ( .A(b[6]), .Z(n1027) );
  CLKBUF_X1 U959 ( .A(n867), .Z(n17) );
  BUF_X2 U960 ( .A(n867), .Z(n18) );
  BUF_X2 U961 ( .A(b[5]), .Z(n848) );
  BUF_X4 U962 ( .A(a[9]), .Z(n25) );
  BUF_X4 U963 ( .A(a[5]), .Z(n13) );
  BUF_X2 U964 ( .A(b[6]), .Z(n847) );
  NOR2_X1 U965 ( .A1(n431), .A2(n444), .ZN(n1029) );
  NAND2_X1 U966 ( .A1(n197), .A2(n151), .ZN(n1030) );
  NOR2_X1 U967 ( .A1(n345), .A2(n350), .ZN(n144) );
  NOR2_X1 U968 ( .A1(n341), .A2(n344), .ZN(n137) );
  NOR2_X1 U969 ( .A1(n700), .A2(n685), .ZN(n298) );
  NOR2_X1 U970 ( .A1(n531), .A2(n534), .ZN(n282) );
  NOR2_X1 U971 ( .A1(n539), .A2(n540), .ZN(n290) );
  AND2_X1 U972 ( .A1(n977), .A2(n301), .ZN(product[1]) );
  BUF_X1 U973 ( .A(n876), .Z(n9) );
  BUF_X1 U974 ( .A(n875), .Z(n15) );
  BUF_X1 U975 ( .A(n873), .Z(n27) );
  BUF_X1 U976 ( .A(n874), .Z(n21) );
  BUF_X1 U977 ( .A(n875), .Z(n16) );
  BUF_X1 U978 ( .A(n876), .Z(n10) );
  BUF_X2 U979 ( .A(a[11]), .Z(n31) );
  NOR2_X1 U980 ( .A1(n1017), .A2(n961), .ZN(n214) );
  NOR2_X1 U981 ( .A1(n195), .A2(n162), .ZN(n160) );
  NOR2_X1 U982 ( .A1(n195), .A2(n190), .ZN(n184) );
  NOR2_X1 U983 ( .A1(n195), .A2(n173), .ZN(n171) );
  INV_X1 U984 ( .A(n177), .ZN(n175) );
  INV_X1 U985 ( .A(n98), .ZN(n96) );
  INV_X1 U986 ( .A(n196), .ZN(n194) );
  INV_X1 U987 ( .A(n1030), .ZN(n147) );
  NAND2_X1 U988 ( .A1(n313), .A2(n205), .ZN(n65) );
  XNOR2_X1 U989 ( .A(n234), .B(n69), .ZN(product[15]) );
  NAND2_X1 U990 ( .A1(n317), .A2(n233), .ZN(n69) );
  AOI21_X1 U991 ( .B1(n214), .B2(n234), .A(n215), .ZN(n213) );
  INV_X1 U992 ( .A(n984), .ZN(n314) );
  INV_X1 U993 ( .A(n1001), .ZN(n234) );
  AOI21_X1 U994 ( .B1(n234), .B2(n225), .A(n955), .ZN(n220) );
  AOI21_X1 U995 ( .B1(n234), .B2(n317), .A(n231), .ZN(n229) );
  INV_X1 U996 ( .A(n227), .ZN(n316) );
  NOR2_X1 U997 ( .A1(n124), .A2(n100), .ZN(n98) );
  OAI21_X1 U998 ( .B1(n196), .B2(n173), .A(n174), .ZN(n172) );
  AOI21_X1 U999 ( .B1(n189), .B2(n175), .A(n176), .ZN(n174) );
  INV_X1 U1000 ( .A(n178), .ZN(n176) );
  NAND2_X1 U1001 ( .A1(n188), .A2(n175), .ZN(n173) );
  NOR2_X1 U1002 ( .A1(n227), .A2(n232), .ZN(n225) );
  BUF_X2 U1003 ( .A(n206), .Z(n51) );
  INV_X1 U1004 ( .A(n197), .ZN(n195) );
  INV_X1 U1005 ( .A(n198), .ZN(n196) );
  NOR2_X1 U1006 ( .A1(n211), .A2(n218), .ZN(n209) );
  NOR2_X1 U1007 ( .A1(n177), .A2(n166), .ZN(n164) );
  OAI21_X1 U1008 ( .B1(n196), .B2(n190), .A(n191), .ZN(n185) );
  INV_X1 U1009 ( .A(n993), .ZN(n177) );
  INV_X1 U1010 ( .A(n124), .ZN(n122) );
  NAND2_X1 U1011 ( .A1(n155), .A2(n993), .ZN(n153) );
  INV_X1 U1012 ( .A(n180), .ZN(n178) );
  INV_X1 U1013 ( .A(n961), .ZN(n217) );
  NAND2_X1 U1014 ( .A1(n1028), .A2(n320), .ZN(n241) );
  NAND2_X1 U1015 ( .A1(n122), .A2(n972), .ZN(n109) );
  INV_X1 U1016 ( .A(n150), .ZN(n148) );
  INV_X1 U1017 ( .A(n233), .ZN(n231) );
  INV_X1 U1018 ( .A(n205), .ZN(n203) );
  NAND2_X1 U1019 ( .A1(n320), .A2(n253), .ZN(n72) );
  INV_X1 U1020 ( .A(n252), .ZN(n320) );
  NAND2_X1 U1021 ( .A1(n973), .A2(n272), .ZN(n75) );
  XNOR2_X1 U1022 ( .A(n240), .B(n70), .ZN(product[14]) );
  NAND2_X1 U1023 ( .A1(n318), .A2(n239), .ZN(n70) );
  INV_X1 U1024 ( .A(n238), .ZN(n318) );
  XNOR2_X1 U1025 ( .A(n267), .B(n74), .ZN(product[10]) );
  NAND2_X1 U1026 ( .A1(n966), .A2(n266), .ZN(n74) );
  NOR2_X1 U1027 ( .A1(n431), .A2(n444), .ZN(n227) );
  XOR2_X1 U1028 ( .A(n262), .B(n73), .Z(product[11]) );
  NOR2_X1 U1029 ( .A1(n393), .A2(n404), .ZN(n204) );
  INV_X1 U1030 ( .A(n272), .ZN(n270) );
  XNOR2_X1 U1031 ( .A(n247), .B(n71), .ZN(product[13]) );
  OAI21_X1 U1032 ( .B1(n199), .B2(n205), .A(n200), .ZN(n198) );
  NOR2_X1 U1033 ( .A1(n445), .A2(n458), .ZN(n232) );
  AOI21_X1 U1034 ( .B1(n236), .B2(n255), .A(n237), .ZN(n235) );
  INV_X1 U1035 ( .A(n199), .ZN(n312) );
  NOR2_X1 U1036 ( .A1(n417), .A2(n430), .ZN(n218) );
  NOR2_X1 U1037 ( .A1(n405), .A2(n416), .ZN(n211) );
  NOR2_X1 U1038 ( .A1(n168), .A2(n157), .ZN(n155) );
  INV_X1 U1039 ( .A(n99), .ZN(n97) );
  AOI21_X1 U1040 ( .B1(n123), .B2(n972), .A(n114), .ZN(n110) );
  INV_X1 U1041 ( .A(n136), .ZN(n134) );
  AOI21_X1 U1042 ( .B1(n1028), .B2(n251), .A(n1018), .ZN(n242) );
  NAND2_X1 U1043 ( .A1(n393), .A2(n404), .ZN(n205) );
  NAND2_X1 U1044 ( .A1(n445), .A2(n458), .ZN(n233) );
  OAI21_X1 U1045 ( .B1(n196), .B2(n162), .A(n163), .ZN(n161) );
  AOI21_X1 U1046 ( .B1(n164), .B2(n189), .A(n165), .ZN(n163) );
  NAND2_X1 U1047 ( .A1(n417), .A2(n430), .ZN(n219) );
  NAND2_X1 U1048 ( .A1(n972), .A2(n968), .ZN(n100) );
  INV_X1 U1049 ( .A(n190), .ZN(n188) );
  NAND2_X1 U1050 ( .A1(n135), .A2(n967), .ZN(n124) );
  NAND2_X1 U1051 ( .A1(n405), .A2(n416), .ZN(n212) );
  INV_X1 U1052 ( .A(n191), .ZN(n189) );
  INV_X1 U1053 ( .A(n253), .ZN(n251) );
  INV_X1 U1054 ( .A(n125), .ZN(n123) );
  INV_X1 U1055 ( .A(n167), .ZN(n166) );
  INV_X1 U1056 ( .A(n168), .ZN(n167) );
  NAND2_X1 U1057 ( .A1(n98), .A2(n969), .ZN(n87) );
  INV_X1 U1058 ( .A(n135), .ZN(n133) );
  INV_X1 U1059 ( .A(n266), .ZN(n264) );
  INV_X1 U1060 ( .A(n144), .ZN(n143) );
  INV_X1 U1061 ( .A(n261), .ZN(n259) );
  NAND2_X1 U1062 ( .A1(n326), .A2(n283), .ZN(n78) );
  INV_X1 U1063 ( .A(n282), .ZN(n326) );
  NAND2_X1 U1064 ( .A1(n324), .A2(n275), .ZN(n76) );
  INV_X1 U1065 ( .A(n274), .ZN(n324) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n280), .ZN(n77) );
  XOR2_X1 U1067 ( .A(n93), .B(n54), .Z(product[30]) );
  NAND2_X1 U1068 ( .A1(n969), .A2(n92), .ZN(n54) );
  XNOR2_X1 U1069 ( .A(n79), .B(n289), .ZN(product[5]) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n288), .ZN(n79) );
  NOR2_X1 U1071 ( .A1(n357), .A2(n364), .ZN(n168) );
  INV_X1 U1072 ( .A(n137), .ZN(n306) );
  AOI21_X1 U1073 ( .B1(n136), .B2(n967), .A(n127), .ZN(n125) );
  INV_X1 U1074 ( .A(n129), .ZN(n127) );
  NOR2_X1 U1075 ( .A1(n351), .A2(n356), .ZN(n157) );
  OAI21_X1 U1076 ( .B1(n145), .B2(n137), .A(n138), .ZN(n136) );
  OAI21_X1 U1077 ( .B1(n125), .B2(n100), .A(n101), .ZN(n99) );
  AOI21_X1 U1078 ( .B1(n114), .B2(n968), .A(n103), .ZN(n101) );
  INV_X1 U1079 ( .A(n105), .ZN(n103) );
  OAI21_X1 U1080 ( .B1(n282), .B2(n284), .A(n283), .ZN(n281) );
  AOI21_X1 U1081 ( .B1(n281), .B2(n974), .A(n278), .ZN(n276) );
  INV_X1 U1082 ( .A(n280), .ZN(n278) );
  NOR2_X1 U1083 ( .A1(n373), .A2(n382), .ZN(n190) );
  NOR2_X1 U1084 ( .A1(n144), .A2(n137), .ZN(n135) );
  AOI21_X1 U1085 ( .B1(n975), .B2(n289), .A(n286), .ZN(n284) );
  INV_X1 U1086 ( .A(n288), .ZN(n286) );
  NOR2_X1 U1087 ( .A1(n483), .A2(n492), .ZN(n252) );
  NAND2_X1 U1088 ( .A1(n345), .A2(n350), .ZN(n145) );
  NAND2_X1 U1089 ( .A1(n373), .A2(n382), .ZN(n191) );
  AOI21_X1 U1090 ( .B1(n99), .B2(n969), .A(n90), .ZN(n88) );
  INV_X1 U1091 ( .A(n92), .ZN(n90) );
  NAND2_X1 U1092 ( .A1(n483), .A2(n492), .ZN(n253) );
  NAND2_X1 U1093 ( .A1(n503), .A2(n510), .ZN(n266) );
  NAND2_X1 U1094 ( .A1(n511), .A2(n518), .ZN(n272) );
  NAND2_X1 U1095 ( .A1(n383), .A2(n392), .ZN(n200) );
  NAND2_X1 U1096 ( .A1(n357), .A2(n364), .ZN(n169) );
  NAND2_X1 U1097 ( .A1(n493), .A2(n502), .ZN(n261) );
  NAND2_X1 U1098 ( .A1(n459), .A2(n470), .ZN(n239) );
  NAND2_X1 U1099 ( .A1(n351), .A2(n356), .ZN(n158) );
  INV_X1 U1100 ( .A(n116), .ZN(n114) );
  XOR2_X1 U1101 ( .A(n80), .B(n292), .Z(product[4]) );
  NAND2_X1 U1102 ( .A1(n328), .A2(n291), .ZN(n80) );
  INV_X1 U1103 ( .A(n290), .ZN(n328) );
  XOR2_X1 U1104 ( .A(n82), .B(n301), .Z(product[2]) );
  NAND2_X1 U1105 ( .A1(n330), .A2(n299), .ZN(n82) );
  INV_X1 U1106 ( .A(n298), .ZN(n330) );
  XNOR2_X1 U1107 ( .A(n81), .B(n297), .ZN(product[3]) );
  AOI21_X1 U1108 ( .B1(n971), .B2(n297), .A(n294), .ZN(n292) );
  INV_X1 U1109 ( .A(n296), .ZN(n294) );
  OAI21_X1 U1110 ( .B1(n298), .B2(n301), .A(n299), .ZN(n297) );
  OAI21_X1 U1111 ( .B1(n290), .B2(n292), .A(n291), .ZN(n289) );
  NAND2_X1 U1112 ( .A1(n700), .A2(n685), .ZN(n299) );
  NAND2_X1 U1113 ( .A1(n574), .A2(n332), .ZN(n92) );
  INV_X1 U1114 ( .A(n332), .ZN(n333) );
  NOR2_X1 U1115 ( .A1(n519), .A2(n524), .ZN(n274) );
  INV_X1 U1116 ( .A(n428), .ZN(n429) );
  OR2_X1 U1117 ( .A1(n643), .A2(n601), .ZN(n442) );
  INV_X1 U1118 ( .A(n362), .ZN(n363) );
  XNOR2_X1 U1119 ( .A(n643), .B(n601), .ZN(n443) );
  NAND2_X1 U1120 ( .A1(n535), .A2(n538), .ZN(n288) );
  NAND2_X1 U1121 ( .A1(n525), .A2(n530), .ZN(n280) );
  NAND2_X1 U1122 ( .A1(n337), .A2(n340), .ZN(n129) );
  NAND2_X1 U1123 ( .A1(n341), .A2(n344), .ZN(n138) );
  NAND2_X1 U1124 ( .A1(n336), .A2(n335), .ZN(n116) );
  NAND2_X1 U1125 ( .A1(n334), .A2(n333), .ZN(n105) );
  NAND2_X1 U1126 ( .A1(n531), .A2(n534), .ZN(n283) );
  NAND2_X1 U1127 ( .A1(n519), .A2(n524), .ZN(n275) );
  OAI22_X1 U1128 ( .A1(n41), .A2(n720), .B1(n40), .B2(n719), .ZN(n338) );
  OAI22_X1 U1129 ( .A1(n12), .A2(n805), .B1(n10), .B2(n804), .ZN(n428) );
  OAI22_X1 U1130 ( .A1(n18), .A2(n788), .B1(n16), .B2(n787), .ZN(n402) );
  OAI22_X1 U1131 ( .A1(n30), .A2(n754), .B1(n28), .B2(n753), .ZN(n362) );
  OAI22_X1 U1132 ( .A1(n24), .A2(n771), .B1(n22), .B2(n770), .ZN(n380) );
  OAI22_X1 U1133 ( .A1(n1002), .A2(n731), .B1(n39), .B2(n730), .ZN(n601) );
  OAI22_X1 U1134 ( .A1(n24), .A2(n776), .B1(n22), .B2(n775), .ZN(n643) );
  OAI22_X1 U1135 ( .A1(n48), .A2(n704), .B1(n45), .B2(n703), .ZN(n575) );
  INV_X1 U1136 ( .A(n545), .ZN(n590) );
  AOI21_X1 U1137 ( .B1(n42), .B2(n40), .A(n719), .ZN(n545) );
  OAI22_X1 U1138 ( .A1(n48), .A2(n705), .B1(n45), .B2(n704), .ZN(n576) );
  INV_X1 U1139 ( .A(n338), .ZN(n339) );
  OAI22_X1 U1140 ( .A1(n48), .A2(n706), .B1(n45), .B2(n705), .ZN(n577) );
  OAI22_X1 U1141 ( .A1(n11), .A2(n817), .B1(n9), .B2(n816), .ZN(n682) );
  OAI22_X1 U1142 ( .A1(n6), .A2(n832), .B1(n831), .B2(n3), .ZN(n697) );
  OAI22_X1 U1143 ( .A1(n18), .A2(n801), .B1(n15), .B2(n800), .ZN(n667) );
  OAI22_X1 U1144 ( .A1(n11), .A2(n818), .B1(n9), .B2(n817), .ZN(n683) );
  OAI22_X1 U1145 ( .A1(n991), .A2(n833), .B1(n832), .B2(n3), .ZN(n698) );
  AND2_X1 U1146 ( .A1(n1033), .A2(n558), .ZN(n669) );
  OAI22_X1 U1147 ( .A1(n48), .A2(n878), .B1(n718), .B2(n45), .ZN(n566) );
  OAI22_X1 U1148 ( .A1(n47), .A2(n717), .B1(n45), .B2(n716), .ZN(n588) );
  OR2_X1 U1149 ( .A1(n1032), .A2(n878), .ZN(n718) );
  OAI22_X1 U1150 ( .A1(n5), .A2(n829), .B1(n828), .B2(n3), .ZN(n694) );
  AND2_X1 U1151 ( .A1(n1033), .A2(n552), .ZN(n637) );
  OAI22_X1 U1152 ( .A1(n18), .A2(n799), .B1(n15), .B2(n798), .ZN(n665) );
  OAI22_X1 U1153 ( .A1(n18), .A2(n792), .B1(n16), .B2(n791), .ZN(n658) );
  OAI22_X1 U1154 ( .A1(n29), .A2(n762), .B1(n27), .B2(n761), .ZN(n630) );
  OAI22_X1 U1155 ( .A1(n6), .A2(n822), .B1(n821), .B2(n877), .ZN(n687) );
  OAI22_X1 U1156 ( .A1(n11), .A2(n816), .B1(n9), .B2(n815), .ZN(n681) );
  AND2_X1 U1157 ( .A1(n1033), .A2(n555), .ZN(n653) );
  OAI22_X1 U1158 ( .A1(n5), .A2(n831), .B1(n830), .B2(n3), .ZN(n696) );
  OAI22_X1 U1159 ( .A1(n5), .A2(n825), .B1(n824), .B2(n877), .ZN(n690) );
  AND2_X1 U1160 ( .A1(n1033), .A2(n546), .ZN(n605) );
  OAI22_X1 U1161 ( .A1(n29), .A2(n990), .B1(n27), .B2(n764), .ZN(n633) );
  OAI22_X1 U1162 ( .A1(n24), .A2(n775), .B1(n22), .B2(n774), .ZN(n642) );
  OAI22_X1 U1163 ( .A1(n30), .A2(n760), .B1(n759), .B2(n28), .ZN(n628) );
  OAI22_X1 U1164 ( .A1(n41), .A2(n730), .B1(n39), .B2(n729), .ZN(n600) );
  OAI22_X1 U1165 ( .A1(n18), .A2(n791), .B1(n16), .B2(n790), .ZN(n657) );
  OAI22_X1 U1166 ( .A1(n746), .A2(n992), .B1(n33), .B2(n745), .ZN(n615) );
  OAI22_X1 U1167 ( .A1(n12), .A2(n806), .B1(n10), .B2(n805), .ZN(n671) );
  OAI22_X1 U1168 ( .A1(n35), .A2(n747), .B1(n33), .B2(n746), .ZN(n616) );
  OAI22_X1 U1169 ( .A1(n1002), .A2(n732), .B1(n39), .B2(n731), .ZN(n602) );
  OAI22_X1 U1170 ( .A1(n24), .A2(n777), .B1(n22), .B2(n776), .ZN(n644) );
  OAI22_X1 U1171 ( .A1(n47), .A2(n712), .B1(n45), .B2(n711), .ZN(n583) );
  INV_X1 U1172 ( .A(n557), .ZN(n654) );
  AOI21_X1 U1173 ( .B1(n18), .B2(n16), .A(n787), .ZN(n557) );
  AOI21_X1 U1174 ( .B1(n24), .B2(n22), .A(n770), .ZN(n554) );
  AOI21_X1 U1175 ( .B1(n30), .B2(n28), .A(n753), .ZN(n551) );
  AOI21_X1 U1176 ( .B1(n991), .B2(n3), .A(n821), .ZN(n563) );
  OAI22_X1 U1177 ( .A1(n17), .A2(n883), .B1(n803), .B2(n16), .ZN(n571) );
  OAI22_X1 U1178 ( .A1(n17), .A2(n802), .B1(n15), .B2(n801), .ZN(n668) );
  OR2_X1 U1179 ( .A1(n1032), .A2(n883), .ZN(n803) );
  NAND2_X1 U1180 ( .A1(n701), .A2(n573), .ZN(n301) );
  AND2_X1 U1181 ( .A1(n1033), .A2(n561), .ZN(n685) );
  INV_X1 U1182 ( .A(n9), .ZN(n561) );
  OAI22_X1 U1183 ( .A1(n48), .A2(n707), .B1(n45), .B2(n706), .ZN(n578) );
  OAI22_X1 U1184 ( .A1(n1002), .A2(n722), .B1(n40), .B2(n721), .ZN(n592) );
  OAI22_X1 U1185 ( .A1(n992), .A2(n744), .B1(n33), .B2(n743), .ZN(n613) );
  OAI22_X1 U1186 ( .A1(n30), .A2(n759), .B1(n28), .B2(n758), .ZN(n627) );
  OAI22_X1 U1187 ( .A1(n35), .A2(n750), .B1(n33), .B2(n749), .ZN(n619) );
  OAI22_X1 U1188 ( .A1(n23), .A2(n780), .B1(n21), .B2(n779), .ZN(n647) );
  OAI22_X1 U1189 ( .A1(n12), .A2(n810), .B1(n10), .B2(n809), .ZN(n675) );
  OAI22_X1 U1190 ( .A1(n12), .A2(n809), .B1(n10), .B2(n808), .ZN(n674) );
  OAI22_X1 U1191 ( .A1(n23), .A2(n779), .B1(n21), .B2(n778), .ZN(n646) );
  OAI22_X1 U1192 ( .A1(n6), .A2(n824), .B1(n823), .B2(n877), .ZN(n689) );
  OAI22_X1 U1193 ( .A1(n992), .A2(n740), .B1(n34), .B2(n739), .ZN(n609) );
  OAI22_X1 U1194 ( .A1(n1002), .A2(n725), .B1(n40), .B2(n724), .ZN(n595) );
  OAI22_X1 U1195 ( .A1(n36), .A2(n741), .B1(n34), .B2(n740), .ZN(n610) );
  INV_X1 U1196 ( .A(n380), .ZN(n381) );
  OAI22_X1 U1197 ( .A1(n35), .A2(n742), .B1(n34), .B2(n741), .ZN(n611) );
  OAI22_X1 U1198 ( .A1(n24), .A2(n772), .B1(n22), .B2(n771), .ZN(n639) );
  OAI22_X1 U1199 ( .A1(n1002), .A2(n727), .B1(n39), .B2(n726), .ZN(n597) );
  OAI22_X1 U1200 ( .A1(n29), .A2(n764), .B1(n27), .B2(n763), .ZN(n632) );
  OAI22_X1 U1201 ( .A1(n35), .A2(n749), .B1(n33), .B2(n748), .ZN(n618) );
  OAI22_X1 U1202 ( .A1(n18), .A2(n794), .B1(n16), .B2(n793), .ZN(n660) );
  OAI22_X1 U1203 ( .A1(n11), .A2(n813), .B1(n9), .B2(n812), .ZN(n678) );
  OAI22_X1 U1204 ( .A1(n23), .A2(n783), .B1(n21), .B2(n782), .ZN(n650) );
  OAI22_X1 U1205 ( .A1(n18), .A2(n798), .B1(n15), .B2(n797), .ZN(n664) );
  OAI22_X1 U1206 ( .A1(n29), .A2(n767), .B1(n27), .B2(n766), .ZN(n635) );
  OAI22_X1 U1207 ( .A1(n18), .A2(n797), .B1(n796), .B2(n15), .ZN(n663) );
  OAI22_X1 U1208 ( .A1(n11), .A2(n812), .B1(n9), .B2(n811), .ZN(n677) );
  OAI22_X1 U1209 ( .A1(n24), .A2(n774), .B1(n22), .B2(n773), .ZN(n641) );
  OAI22_X1 U1210 ( .A1(n42), .A2(n729), .B1(n39), .B2(n728), .ZN(n599) );
  OAI22_X1 U1211 ( .A1(n18), .A2(n789), .B1(n16), .B2(n788), .ZN(n655) );
  OAI22_X1 U1212 ( .A1(n30), .A2(n758), .B1(n28), .B2(n757), .ZN(n626) );
  OAI22_X1 U1213 ( .A1(n773), .A2(n24), .B1(n22), .B2(n772), .ZN(n640) );
  OAI22_X1 U1214 ( .A1(n992), .A2(n743), .B1(n34), .B2(n742), .ZN(n612) );
  OAI22_X1 U1215 ( .A1(n23), .A2(n778), .B1(n21), .B2(n777), .ZN(n645) );
  OAI22_X1 U1216 ( .A1(n18), .A2(n793), .B1(n16), .B2(n792), .ZN(n659) );
  OAI22_X1 U1217 ( .A1(n47), .A2(n710), .B1(n45), .B2(n709), .ZN(n581) );
  OAI22_X1 U1218 ( .A1(n30), .A2(n755), .B1(n28), .B2(n754), .ZN(n623) );
  INV_X1 U1219 ( .A(n554), .ZN(n638) );
  OAI22_X1 U1220 ( .A1(n42), .A2(n721), .B1(n40), .B2(n720), .ZN(n591) );
  INV_X1 U1221 ( .A(n548), .ZN(n606) );
  AOI21_X1 U1222 ( .B1(n35), .B2(n34), .A(n736), .ZN(n548) );
  OAI22_X1 U1223 ( .A1(n23), .A2(n784), .B1(n21), .B2(n783), .ZN(n651) );
  OAI22_X1 U1224 ( .A1(n11), .A2(n814), .B1(n9), .B2(n813), .ZN(n679) );
  OAI22_X1 U1225 ( .A1(n12), .A2(n807), .B1(n10), .B2(n806), .ZN(n672) );
  OAI22_X1 U1226 ( .A1(n5), .A2(n828), .B1(n827), .B2(n877), .ZN(n693) );
  OAI22_X1 U1227 ( .A1(n6), .A2(n830), .B1(n829), .B2(n3), .ZN(n695) );
  OAI22_X1 U1228 ( .A1(n11), .A2(n815), .B1(n9), .B2(n814), .ZN(n680) );
  OAI22_X1 U1229 ( .A1(n18), .A2(n800), .B1(n15), .B2(n799), .ZN(n666) );
  OAI22_X1 U1230 ( .A1(n991), .A2(n827), .B1(n826), .B2(n877), .ZN(n692) );
  OAI22_X1 U1231 ( .A1(n23), .A2(n782), .B1(n21), .B2(n781), .ZN(n649) );
  AND2_X1 U1232 ( .A1(n1033), .A2(n549), .ZN(n621) );
  OAI22_X1 U1233 ( .A1(n47), .A2(n711), .B1(n45), .B2(n710), .ZN(n582) );
  OAI22_X1 U1234 ( .A1(n30), .A2(n756), .B1(n28), .B2(n755), .ZN(n624) );
  OAI22_X1 U1235 ( .A1(n42), .A2(n726), .B1(n40), .B2(n725), .ZN(n596) );
  OAI22_X1 U1236 ( .A1(n29), .A2(n763), .B1(n27), .B2(n762), .ZN(n631) );
  OAI22_X1 U1237 ( .A1(n42), .A2(n733), .B1(n39), .B2(n732), .ZN(n603) );
  OAI22_X1 U1238 ( .A1(n12), .A2(n808), .B1(n10), .B2(n807), .ZN(n673) );
  INV_X1 U1239 ( .A(n560), .ZN(n670) );
  AOI21_X1 U1240 ( .B1(n12), .B2(n10), .A(n804), .ZN(n560) );
  OAI22_X1 U1241 ( .A1(n42), .A2(n723), .B1(n40), .B2(n722), .ZN(n593) );
  OAI22_X1 U1242 ( .A1(n48), .A2(n708), .B1(n45), .B2(n707), .ZN(n579) );
  INV_X1 U1243 ( .A(n551), .ZN(n622) );
  OAI22_X1 U1244 ( .A1(n30), .A2(n757), .B1(n28), .B2(n756), .ZN(n625) );
  OAI22_X1 U1245 ( .A1(n18), .A2(n795), .B1(n15), .B2(n794), .ZN(n661) );
  OAI22_X1 U1246 ( .A1(n23), .A2(n781), .B1(n21), .B2(n780), .ZN(n648) );
  OAI22_X1 U1247 ( .A1(n12), .A2(n811), .B1(n10), .B2(n810), .ZN(n676) );
  OAI22_X1 U1248 ( .A1(n36), .A2(n738), .B1(n34), .B2(n737), .ZN(n607) );
  OAI22_X1 U1249 ( .A1(n47), .A2(n716), .B1(n46), .B2(n715), .ZN(n587) );
  OAI22_X1 U1250 ( .A1(n29), .A2(n761), .B1(n27), .B2(n760), .ZN(n629) );
  INV_X1 U1251 ( .A(n563), .ZN(n686) );
  OAI22_X1 U1252 ( .A1(n826), .A2(n5), .B1(n825), .B2(n3), .ZN(n691) );
  OAI22_X1 U1253 ( .A1(n796), .A2(n17), .B1(n795), .B2(n15), .ZN(n662) );
  OAI22_X1 U1254 ( .A1(n47), .A2(n715), .B1(n46), .B2(n714), .ZN(n586) );
  OAI22_X1 U1255 ( .A1(n35), .A2(n745), .B1(n33), .B2(n744), .ZN(n614) );
  OAI22_X1 U1256 ( .A1(n17), .A2(n790), .B1(n16), .B2(n789), .ZN(n656) );
  OAI22_X1 U1257 ( .A1(n36), .A2(n739), .B1(n34), .B2(n738), .ZN(n608) );
  OAI22_X1 U1258 ( .A1(n41), .A2(n724), .B1(n40), .B2(n723), .ZN(n594) );
  OAI22_X1 U1259 ( .A1(n48), .A2(n709), .B1(n45), .B2(n708), .ZN(n580) );
  INV_X1 U1260 ( .A(n46), .ZN(n543) );
  NAND2_X1 U1261 ( .A1(n539), .A2(n540), .ZN(n291) );
  INV_X1 U1262 ( .A(n542), .ZN(n574) );
  AOI21_X1 U1263 ( .B1(n48), .B2(n45), .A(n702), .ZN(n542) );
  OAI22_X1 U1264 ( .A1(n1002), .A2(n728), .B1(n39), .B2(n727), .ZN(n598) );
  OAI22_X1 U1265 ( .A1(n47), .A2(n713), .B1(n45), .B2(n712), .ZN(n584) );
  INV_X1 U1266 ( .A(n402), .ZN(n403) );
  OAI22_X1 U1267 ( .A1(n6), .A2(n823), .B1(n822), .B2(n3), .ZN(n688) );
  OAI22_X1 U1268 ( .A1(n36), .A2(n748), .B1(n33), .B2(n747), .ZN(n617) );
  AND2_X1 U1269 ( .A1(n1033), .A2(n543), .ZN(n589) );
  AND2_X1 U1270 ( .A1(n1033), .A2(n564), .ZN(product[0]) );
  INV_X1 U1271 ( .A(n3), .ZN(n564) );
  OR2_X1 U1272 ( .A1(n1032), .A2(n880), .ZN(n752) );
  OR2_X1 U1273 ( .A1(n1033), .A2(n881), .ZN(n769) );
  OR2_X1 U1274 ( .A1(n1032), .A2(n879), .ZN(n735) );
  OR2_X1 U1275 ( .A1(n1033), .A2(n882), .ZN(n786) );
  INV_X1 U1276 ( .A(n15), .ZN(n558) );
  INV_X1 U1277 ( .A(n21), .ZN(n555) );
  INV_X1 U1278 ( .A(n39), .ZN(n546) );
  INV_X1 U1279 ( .A(n33), .ZN(n549) );
  INV_X1 U1280 ( .A(n27), .ZN(n552) );
  OR2_X1 U1281 ( .A1(n1032), .A2(n885), .ZN(n837) );
  INV_X1 U1282 ( .A(n1), .ZN(n885) );
  BUF_X1 U1283 ( .A(n863), .Z(n42) );
  OAI22_X1 U1284 ( .A1(n41), .A2(n734), .B1(n39), .B2(n733), .ZN(n604) );
  OAI22_X1 U1285 ( .A1(n41), .A2(n879), .B1(n735), .B2(n39), .ZN(n567) );
  OAI22_X1 U1286 ( .A1(n5), .A2(n836), .B1(n835), .B2(n3), .ZN(n701) );
  BUF_X1 U1287 ( .A(n869), .Z(n5) );
  OAI22_X1 U1288 ( .A1(n29), .A2(n768), .B1(n27), .B2(n767), .ZN(n636) );
  OAI22_X1 U1289 ( .A1(n30), .A2(n881), .B1(n769), .B2(n28), .ZN(n569) );
  OAI22_X1 U1290 ( .A1(n991), .A2(n834), .B1(n833), .B2(n3), .ZN(n699) );
  OAI22_X1 U1291 ( .A1(n11), .A2(n819), .B1(n9), .B2(n818), .ZN(n684) );
  OAI22_X1 U1292 ( .A1(n36), .A2(n751), .B1(n33), .B2(n750), .ZN(n620) );
  OAI22_X1 U1293 ( .A1(n36), .A2(n880), .B1(n752), .B2(n34), .ZN(n568) );
  BUF_X1 U1294 ( .A(n872), .Z(n33) );
  BUF_X1 U1295 ( .A(n874), .Z(n22) );
  BUF_X1 U1296 ( .A(n873), .Z(n28) );
  BUF_X1 U1297 ( .A(n872), .Z(n34) );
  BUF_X1 U1298 ( .A(n869), .Z(n6) );
  BUF_X1 U1299 ( .A(n868), .Z(n11) );
  OAI22_X1 U1300 ( .A1(n23), .A2(n785), .B1(n21), .B2(n784), .ZN(n652) );
  OAI22_X1 U1301 ( .A1(n24), .A2(n882), .B1(n786), .B2(n22), .ZN(n570) );
  OAI22_X1 U1302 ( .A1(n12), .A2(n884), .B1(n820), .B2(n10), .ZN(n572) );
  OR2_X1 U1303 ( .A1(n1033), .A2(n884), .ZN(n820) );
  INV_X1 U1304 ( .A(n7), .ZN(n884) );
  INV_X1 U1305 ( .A(n25), .ZN(n881) );
  INV_X1 U1306 ( .A(n31), .ZN(n880) );
  INV_X1 U1307 ( .A(n37), .ZN(n879) );
  INV_X1 U1308 ( .A(n19), .ZN(n882) );
  INV_X1 U1309 ( .A(n13), .ZN(n883) );
  INV_X1 U1310 ( .A(n43), .ZN(n878) );
  XNOR2_X1 U1311 ( .A(a[10]), .B(a[9]), .ZN(n872) );
  BUF_X2 U1312 ( .A(a[3]), .Z(n7) );
  BUF_X2 U1313 ( .A(a[7]), .Z(n19) );
  NAND2_X1 U1314 ( .A1(n856), .A2(n872), .ZN(n864) );
  NAND2_X1 U1315 ( .A1(n861), .A2(n877), .ZN(n869) );
  INV_X1 U1316 ( .A(a[0]), .ZN(n877) );
  XNOR2_X1 U1317 ( .A(a[12]), .B(a[11]), .ZN(n871) );
  OAI22_X1 U1318 ( .A1(n992), .A2(n737), .B1(n34), .B2(n736), .ZN(n348) );
  INV_X1 U1319 ( .A(n348), .ZN(n349) );
  OAI22_X1 U1320 ( .A1(n6), .A2(n885), .B1(n837), .B2(n877), .ZN(n573) );
  BUF_X1 U1321 ( .A(n863), .Z(n41) );
  NAND2_X1 U1322 ( .A1(n855), .A2(n871), .ZN(n863) );
  CLKBUF_X1 U1323 ( .A(n871), .Z(n40) );
  NAND2_X1 U1324 ( .A1(n854), .A2(n870), .ZN(n862) );
  OAI22_X1 U1325 ( .A1(n47), .A2(n714), .B1(n45), .B2(n713), .ZN(n585) );
  NAND2_X1 U1326 ( .A1(n164), .A2(n188), .ZN(n162) );
  NOR2_X1 U1327 ( .A1(n190), .A2(n153), .ZN(n151) );
  OAI21_X1 U1328 ( .B1(n224), .B2(n961), .A(n219), .ZN(n215) );
  NAND2_X1 U1329 ( .A1(n431), .A2(n444), .ZN(n228) );
  INV_X1 U1330 ( .A(n182), .ZN(n180) );
  OAI21_X1 U1331 ( .B1(n178), .B2(n166), .A(n169), .ZN(n165) );
  OAI21_X1 U1332 ( .B1(n254), .B2(n241), .A(n1003), .ZN(n240) );
  XOR2_X1 U1333 ( .A(n254), .B(n72), .Z(product[12]) );
  OAI21_X1 U1334 ( .B1(n254), .B2(n252), .A(n253), .ZN(n247) );
  CLKBUF_X1 U1335 ( .A(n870), .Z(n46) );
  INV_X1 U1336 ( .A(n204), .ZN(n313) );
  NAND2_X1 U1337 ( .A1(n858), .A2(n874), .ZN(n866) );
  NAND2_X1 U1338 ( .A1(n857), .A2(n873), .ZN(n865) );
  OAI22_X1 U1339 ( .A1(n766), .A2(n29), .B1(n27), .B2(n765), .ZN(n634) );
  NOR2_X1 U1340 ( .A1(n1030), .A2(n87), .ZN(n85) );
  NOR2_X1 U1341 ( .A1(n1030), .A2(n96), .ZN(n94) );
  NOR2_X1 U1342 ( .A1(n1030), .A2(n144), .ZN(n140) );
  NOR2_X1 U1343 ( .A1(n1030), .A2(n133), .ZN(n131) );
  NOR2_X1 U1344 ( .A1(n1030), .A2(n109), .ZN(n107) );
  NOR2_X1 U1345 ( .A1(n1030), .A2(n124), .ZN(n118) );
  INV_X1 U1346 ( .A(n255), .ZN(n254) );
  XNOR2_X1 U1347 ( .A(n7), .B(n841), .ZN(n807) );
  XNOR2_X1 U1348 ( .A(n7), .B(n847), .ZN(n813) );
  XNOR2_X1 U1349 ( .A(n7), .B(n848), .ZN(n814) );
  XNOR2_X1 U1350 ( .A(n7), .B(n840), .ZN(n806) );
  XNOR2_X1 U1351 ( .A(n7), .B(n960), .ZN(n816) );
  XNOR2_X1 U1352 ( .A(n7), .B(n842), .ZN(n808) );
  XNOR2_X1 U1353 ( .A(n7), .B(n849), .ZN(n815) );
  XNOR2_X1 U1354 ( .A(n7), .B(n846), .ZN(n812) );
  XNOR2_X1 U1355 ( .A(n7), .B(n845), .ZN(n811) );
  XNOR2_X1 U1356 ( .A(n7), .B(n851), .ZN(n817) );
  XNOR2_X1 U1357 ( .A(n7), .B(n979), .ZN(n810) );
  XNOR2_X1 U1358 ( .A(n7), .B(n843), .ZN(n809) );
  XNOR2_X1 U1359 ( .A(n7), .B(n839), .ZN(n805) );
  XNOR2_X1 U1360 ( .A(n7), .B(n1032), .ZN(n819) );
  XNOR2_X1 U1361 ( .A(n7), .B(n838), .ZN(n804) );
  XNOR2_X1 U1362 ( .A(n7), .B(n852), .ZN(n818) );
  OAI21_X1 U1363 ( .B1(n276), .B2(n274), .A(n275), .ZN(n273) );
  XNOR2_X1 U1364 ( .A(n19), .B(n1033), .ZN(n785) );
  XNOR2_X1 U1365 ( .A(n19), .B(n979), .ZN(n776) );
  XNOR2_X1 U1366 ( .A(n19), .B(n845), .ZN(n777) );
  XNOR2_X1 U1367 ( .A(n19), .B(n852), .ZN(n784) );
  XNOR2_X1 U1368 ( .A(n19), .B(n851), .ZN(n783) );
  XNOR2_X1 U1369 ( .A(n19), .B(n839), .ZN(n771) );
  XNOR2_X1 U1370 ( .A(n19), .B(n843), .ZN(n775) );
  XNOR2_X1 U1371 ( .A(n19), .B(n846), .ZN(n778) );
  XNOR2_X1 U1372 ( .A(n19), .B(n960), .ZN(n782) );
  XNOR2_X1 U1373 ( .A(n19), .B(n848), .ZN(n780) );
  XNOR2_X1 U1374 ( .A(n19), .B(n842), .ZN(n774) );
  XNOR2_X1 U1375 ( .A(n19), .B(n840), .ZN(n772) );
  XNOR2_X1 U1376 ( .A(n19), .B(n849), .ZN(n781) );
  XNOR2_X1 U1377 ( .A(n19), .B(n847), .ZN(n779) );
  XNOR2_X1 U1378 ( .A(n19), .B(n841), .ZN(n773) );
  XNOR2_X1 U1379 ( .A(n19), .B(n838), .ZN(n770) );
  NAND2_X1 U1380 ( .A1(n209), .A2(n225), .ZN(n207) );
  XNOR2_X1 U1381 ( .A(n43), .B(n840), .ZN(n704) );
  XNOR2_X1 U1382 ( .A(n43), .B(n841), .ZN(n705) );
  XNOR2_X1 U1383 ( .A(n43), .B(n996), .ZN(n703) );
  XNOR2_X1 U1384 ( .A(n43), .B(n838), .ZN(n702) );
  XNOR2_X1 U1385 ( .A(n43), .B(n843), .ZN(n707) );
  XNOR2_X1 U1386 ( .A(n43), .B(n842), .ZN(n706) );
  XNOR2_X1 U1387 ( .A(n43), .B(n979), .ZN(n708) );
  XNOR2_X1 U1388 ( .A(n43), .B(n1027), .ZN(n711) );
  XNOR2_X1 U1389 ( .A(n43), .B(n846), .ZN(n710) );
  XNOR2_X1 U1390 ( .A(n43), .B(n1032), .ZN(n717) );
  XNOR2_X1 U1391 ( .A(n43), .B(n845), .ZN(n709) );
  XNOR2_X1 U1392 ( .A(n43), .B(n848), .ZN(n712) );
  XNOR2_X1 U1393 ( .A(n43), .B(n852), .ZN(n716) );
  XNOR2_X1 U1394 ( .A(n43), .B(n851), .ZN(n715) );
  XNOR2_X1 U1395 ( .A(n43), .B(n850), .ZN(n714) );
  XNOR2_X1 U1396 ( .A(n43), .B(n849), .ZN(n713) );
  NAND2_X1 U1397 ( .A1(n1028), .A2(n246), .ZN(n71) );
  OAI21_X1 U1398 ( .B1(n256), .B2(n268), .A(n257), .ZN(n255) );
  NAND2_X1 U1399 ( .A1(n970), .A2(n966), .ZN(n256) );
  AOI21_X1 U1400 ( .B1(n970), .B2(n264), .A(n259), .ZN(n257) );
  XNOR2_X1 U1401 ( .A(n25), .B(n841), .ZN(n756) );
  XNOR2_X1 U1402 ( .A(n25), .B(n838), .ZN(n753) );
  XNOR2_X1 U1403 ( .A(n25), .B(n1033), .ZN(n768) );
  XNOR2_X1 U1404 ( .A(n25), .B(n840), .ZN(n755) );
  XNOR2_X1 U1405 ( .A(n25), .B(n839), .ZN(n754) );
  XNOR2_X1 U1406 ( .A(n25), .B(n843), .ZN(n758) );
  XNOR2_X1 U1407 ( .A(n25), .B(n845), .ZN(n760) );
  XNOR2_X1 U1408 ( .A(n25), .B(n842), .ZN(n757) );
  XNOR2_X1 U1409 ( .A(n1027), .B(n25), .ZN(n762) );
  XNOR2_X1 U1410 ( .A(n25), .B(n844), .ZN(n759) );
  XNOR2_X1 U1411 ( .A(n25), .B(n848), .ZN(n763) );
  XNOR2_X1 U1412 ( .A(n25), .B(n846), .ZN(n761) );
  XNOR2_X1 U1413 ( .A(n25), .B(n852), .ZN(n767) );
  XNOR2_X1 U1414 ( .A(n25), .B(n849), .ZN(n764) );
  XNOR2_X1 U1415 ( .A(n25), .B(n851), .ZN(n766) );
  XNOR2_X1 U1416 ( .A(n25), .B(n960), .ZN(n765) );
  NAND2_X1 U1417 ( .A1(n970), .A2(n261), .ZN(n73) );
  AOI21_X1 U1418 ( .B1(n267), .B2(n966), .A(n264), .ZN(n262) );
  OAI22_X1 U1419 ( .A1(n991), .A2(n835), .B1(n834), .B2(n3), .ZN(n700) );
  OAI21_X1 U1420 ( .B1(n150), .B2(n87), .A(n88), .ZN(n86) );
  OAI21_X1 U1421 ( .B1(n150), .B2(n96), .A(n97), .ZN(n95) );
  OAI21_X1 U1422 ( .B1(n150), .B2(n109), .A(n110), .ZN(n108) );
  OAI21_X1 U1423 ( .B1(n150), .B2(n124), .A(n125), .ZN(n119) );
  OAI21_X1 U1424 ( .B1(n150), .B2(n133), .A(n134), .ZN(n132) );
  OAI21_X1 U1425 ( .B1(n150), .B2(n144), .A(n145), .ZN(n141) );
  AOI21_X1 U1426 ( .B1(n209), .B2(n226), .A(n210), .ZN(n208) );
  INV_X1 U1427 ( .A(n955), .ZN(n224) );
  OAI21_X1 U1428 ( .B1(n1029), .B2(n233), .A(n228), .ZN(n226) );
  NOR2_X1 U1429 ( .A1(n204), .A2(n199), .ZN(n197) );
  NAND2_X1 U1430 ( .A1(n971), .A2(n296), .ZN(n81) );
  OAI21_X1 U1431 ( .B1(n153), .B2(n191), .A(n154), .ZN(n152) );
  OAI21_X1 U1432 ( .B1(n1006), .B2(n219), .A(n212), .ZN(n210) );
  NOR2_X1 U1433 ( .A1(n241), .A2(n238), .ZN(n236) );
  OAI21_X1 U1434 ( .B1(n242), .B2(n238), .A(n239), .ZN(n237) );
  XNOR2_X1 U1435 ( .A(n37), .B(n840), .ZN(n721) );
  XNOR2_X1 U1436 ( .A(n37), .B(n841), .ZN(n722) );
  XNOR2_X1 U1437 ( .A(n37), .B(n842), .ZN(n723) );
  XNOR2_X1 U1438 ( .A(n37), .B(n996), .ZN(n720) );
  XNOR2_X1 U1439 ( .A(n37), .B(n838), .ZN(n719) );
  XNOR2_X1 U1440 ( .A(n37), .B(n954), .ZN(n726) );
  XNOR2_X1 U1441 ( .A(n37), .B(n851), .ZN(n732) );
  XNOR2_X1 U1442 ( .A(n37), .B(n960), .ZN(n731) );
  XNOR2_X1 U1443 ( .A(n37), .B(n979), .ZN(n725) );
  XNOR2_X1 U1444 ( .A(n37), .B(n843), .ZN(n724) );
  XNOR2_X1 U1445 ( .A(n37), .B(n852), .ZN(n733) );
  XNOR2_X1 U1446 ( .A(n37), .B(n1027), .ZN(n728) );
  XNOR2_X1 U1447 ( .A(n37), .B(n846), .ZN(n727) );
  XNOR2_X1 U1448 ( .A(n37), .B(n849), .ZN(n730) );
  XNOR2_X1 U1449 ( .A(n848), .B(n37), .ZN(n729) );
  XNOR2_X1 U1450 ( .A(n1), .B(n954), .ZN(n828) );
  XNOR2_X1 U1451 ( .A(n1), .B(n846), .ZN(n829) );
  XNOR2_X1 U1452 ( .A(n1), .B(n847), .ZN(n830) );
  XNOR2_X1 U1453 ( .A(n1), .B(n848), .ZN(n831) );
  XNOR2_X1 U1454 ( .A(n1), .B(n1033), .ZN(n836) );
  XNOR2_X1 U1455 ( .A(n1), .B(n979), .ZN(n827) );
  XNOR2_X1 U1456 ( .A(n1), .B(n839), .ZN(n822) );
  XNOR2_X1 U1457 ( .A(n1), .B(n849), .ZN(n832) );
  XNOR2_X1 U1458 ( .A(n1), .B(n852), .ZN(n835) );
  XNOR2_X1 U1459 ( .A(n1), .B(n840), .ZN(n823) );
  XNOR2_X1 U1460 ( .A(n1), .B(n841), .ZN(n824) );
  XNOR2_X1 U1461 ( .A(n1), .B(n959), .ZN(n833) );
  XNOR2_X1 U1462 ( .A(n1), .B(n851), .ZN(n834) );
  XNOR2_X1 U1463 ( .A(n1), .B(n842), .ZN(n825) );
  XNOR2_X1 U1464 ( .A(n1), .B(n838), .ZN(n821) );
  XNOR2_X1 U1465 ( .A(n1), .B(n843), .ZN(n826) );
  INV_X1 U1466 ( .A(n268), .ZN(n267) );
  OAI21_X1 U1467 ( .B1(n207), .B2(n235), .A(n208), .ZN(n206) );
  XNOR2_X1 U1468 ( .A(n13), .B(n851), .ZN(n800) );
  XNOR2_X1 U1469 ( .A(n13), .B(n843), .ZN(n792) );
  XNOR2_X1 U1470 ( .A(n13), .B(n842), .ZN(n791) );
  XNOR2_X1 U1471 ( .A(n13), .B(n960), .ZN(n799) );
  XNOR2_X1 U1472 ( .A(n13), .B(n849), .ZN(n798) );
  XNOR2_X1 U1473 ( .A(n13), .B(n848), .ZN(n797) );
  XNOR2_X1 U1474 ( .A(n13), .B(n841), .ZN(n790) );
  XNOR2_X1 U1475 ( .A(n13), .B(n840), .ZN(n789) );
  XNOR2_X1 U1476 ( .A(n13), .B(n1032), .ZN(n802) );
  XNOR2_X1 U1477 ( .A(n13), .B(n845), .ZN(n794) );
  XNOR2_X1 U1478 ( .A(n13), .B(n839), .ZN(n788) );
  XNOR2_X1 U1479 ( .A(n13), .B(n979), .ZN(n793) );
  XNOR2_X1 U1480 ( .A(n13), .B(n852), .ZN(n801) );
  XNOR2_X1 U1481 ( .A(n13), .B(n838), .ZN(n787) );
  XNOR2_X1 U1482 ( .A(n13), .B(n847), .ZN(n796) );
  XNOR2_X1 U1483 ( .A(n13), .B(n846), .ZN(n795) );
  OAI21_X1 U1484 ( .B1(n157), .B2(n169), .A(n158), .ZN(n156) );
  INV_X1 U1485 ( .A(n157), .ZN(n308) );
  XNOR2_X1 U1486 ( .A(n995), .B(n843), .ZN(n741) );
  XNOR2_X1 U1487 ( .A(n849), .B(n31), .ZN(n747) );
  XNOR2_X1 U1488 ( .A(n995), .B(n842), .ZN(n740) );
  XNOR2_X1 U1489 ( .A(n995), .B(n840), .ZN(n738) );
  XNOR2_X1 U1490 ( .A(n995), .B(n996), .ZN(n737) );
  XNOR2_X1 U1491 ( .A(n995), .B(n841), .ZN(n739) );
  XNOR2_X1 U1492 ( .A(n995), .B(n851), .ZN(n749) );
  XNOR2_X1 U1493 ( .A(n995), .B(n838), .ZN(n736) );
  XNOR2_X1 U1494 ( .A(n31), .B(n959), .ZN(n748) );
  XNOR2_X1 U1495 ( .A(n995), .B(n848), .ZN(n746) );
  XNOR2_X1 U1496 ( .A(n995), .B(n1032), .ZN(n751) );
  XNOR2_X1 U1497 ( .A(n31), .B(n1027), .ZN(n745) );
  XNOR2_X1 U1498 ( .A(n995), .B(n852), .ZN(n750) );
  XNOR2_X1 U1499 ( .A(n846), .B(n31), .ZN(n744) );
  XNOR2_X1 U1500 ( .A(n995), .B(n845), .ZN(n743) );
  XNOR2_X1 U1501 ( .A(n31), .B(n844), .ZN(n742) );
  AOI21_X1 U1502 ( .B1(n155), .B2(n180), .A(n156), .ZN(n154) );
  NAND2_X1 U1503 ( .A1(n365), .A2(n372), .ZN(n182) );
  NAND2_X1 U1504 ( .A1(n860), .A2(n876), .ZN(n868) );
  XOR2_X1 U1505 ( .A(a[14]), .B(a[15]), .Z(n854) );
  INV_X1 U1506 ( .A(n232), .ZN(n317) );
  NAND2_X1 U1507 ( .A1(n859), .A2(n875), .ZN(n867) );
  XOR2_X1 U1508 ( .A(a[6]), .B(a[7]), .Z(n858) );
  XNOR2_X1 U1509 ( .A(a[8]), .B(a[7]), .ZN(n873) );
  XOR2_X1 U1510 ( .A(a[12]), .B(a[13]), .Z(n855) );
  XNOR2_X1 U1511 ( .A(a[14]), .B(a[13]), .ZN(n870) );
  XOR2_X1 U1512 ( .A(a[8]), .B(a[9]), .Z(n857) );
  XOR2_X1 U1513 ( .A(a[10]), .B(a[11]), .Z(n856) );
  XNOR2_X1 U1514 ( .A(n273), .B(n75), .ZN(product[9]) );
  AOI21_X1 U1515 ( .B1(n273), .B2(n973), .A(n270), .ZN(n268) );
  XOR2_X1 U1516 ( .A(a[1]), .B(a[0]), .Z(n861) );
  XNOR2_X1 U1517 ( .A(a[1]), .B(a[2]), .ZN(n876) );
  AOI21_X1 U1518 ( .B1(n978), .B2(n85), .A(n86), .ZN(n84) );
  AOI21_X1 U1519 ( .B1(n1005), .B2(n94), .A(n95), .ZN(n93) );
  AOI21_X1 U1520 ( .B1(n1005), .B2(n140), .A(n141), .ZN(n139) );
  AOI21_X1 U1521 ( .B1(n1005), .B2(n131), .A(n132), .ZN(n130) );
  AOI21_X1 U1522 ( .B1(n1005), .B2(n147), .A(n148), .ZN(n146) );
  AOI21_X1 U1523 ( .B1(n51), .B2(n160), .A(n161), .ZN(n159) );
  AOI21_X1 U1524 ( .B1(n1005), .B2(n118), .A(n119), .ZN(n117) );
  AOI21_X1 U1525 ( .B1(n1005), .B2(n107), .A(n108), .ZN(n106) );
  AOI21_X1 U1526 ( .B1(n51), .B2(n184), .A(n185), .ZN(n183) );
  AOI21_X1 U1527 ( .B1(n51), .B2(n197), .A(n194), .ZN(n192) );
  XNOR2_X1 U1528 ( .A(n1005), .B(n65), .ZN(product[19]) );
  AOI21_X1 U1529 ( .B1(n51), .B2(n171), .A(n172), .ZN(n170) );
  XNOR2_X1 U1530 ( .A(a[6]), .B(a[5]), .ZN(n874) );
  XOR2_X1 U1531 ( .A(a[4]), .B(a[5]), .Z(n859) );
  NAND2_X1 U1532 ( .A1(n541), .A2(n572), .ZN(n296) );
  XNOR2_X1 U1533 ( .A(a[4]), .B(a[3]), .ZN(n875) );
  XOR2_X1 U1534 ( .A(a[2]), .B(a[3]), .Z(n860) );
  AOI21_X1 U1535 ( .B1(n51), .B2(n313), .A(n203), .ZN(n201) );
  XOR2_X1 U1536 ( .A(n1009), .B(n76), .Z(product[8]) );
  XNOR2_X1 U1537 ( .A(n281), .B(n77), .ZN(product[7]) );
  XOR2_X1 U1538 ( .A(n78), .B(n1010), .Z(product[6]) );
endmodule


module datapath_DW01_add_8 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n40, n41, n42, n43, n44, n45, n46,
         n47, n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n88, n89, n90, n91,
         n92, n93, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n193, n194, n195, n196, n197, n198,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n234, n237, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n281, n284, n286, n290, n292,
         n294, n296, n297, n298, n300, n302, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n440, n441;

  BUF_X2 U349 ( .A(n178), .Z(n2) );
  BUF_X2 U350 ( .A(n178), .Z(n1) );
  NOR2_X1 U351 ( .A1(B[25]), .A2(A[25]), .ZN(n416) );
  OR2_X1 U352 ( .A1(A[26]), .A2(n424), .ZN(n429) );
  OR2_X1 U353 ( .A1(A[30]), .A2(B[30]), .ZN(n417) );
  CLKBUF_X1 U354 ( .A(n436), .Z(n418) );
  INV_X1 U355 ( .A(n105), .ZN(n419) );
  OAI21_X1 U356 ( .B1(n416), .B2(n107), .A(n100), .ZN(n420) );
  NOR2_X1 U357 ( .A1(n151), .A2(n113), .ZN(n421) );
  CLKBUF_X1 U358 ( .A(n136), .Z(n422) );
  NOR2_X1 U359 ( .A1(A[22]), .A2(B[22]), .ZN(n423) );
  CLKBUF_X1 U360 ( .A(B[26]), .Z(n424) );
  CLKBUF_X1 U361 ( .A(n432), .Z(n425) );
  NOR2_X1 U362 ( .A1(A[19]), .A2(B[19]), .ZN(n426) );
  CLKBUF_X1 U363 ( .A(n61), .Z(n427) );
  CLKBUF_X1 U364 ( .A(B[25]), .Z(n428) );
  NOR2_X1 U365 ( .A1(n423), .A2(n117), .ZN(n430) );
  OR2_X1 U366 ( .A1(A[25]), .A2(n428), .ZN(n431) );
  NOR2_X1 U367 ( .A1(B[23]), .A2(A[23]), .ZN(n432) );
  NOR2_X1 U368 ( .A1(B[21]), .A2(A[21]), .ZN(n433) );
  NAND2_X1 U369 ( .A1(n77), .A2(n98), .ZN(n434) );
  INV_X1 U370 ( .A(n78), .ZN(n435) );
  AND2_X2 U371 ( .A1(n434), .A2(n435), .ZN(n5) );
  NOR2_X1 U372 ( .A1(B[27]), .A2(A[27]), .ZN(n436) );
  OR2_X1 U373 ( .A1(n144), .A2(n433), .ZN(n437) );
  BUF_X1 U374 ( .A(n112), .Z(n438) );
  NOR2_X1 U375 ( .A1(A[10]), .A2(B[10]), .ZN(n230) );
  NOR2_X1 U376 ( .A1(A[12]), .A2(B[12]), .ZN(n212) );
  NOR2_X1 U377 ( .A1(A[4]), .A2(B[4]), .ZN(n265) );
  NOR2_X1 U378 ( .A1(A[3]), .A2(B[3]), .ZN(n271) );
  NOR2_X1 U379 ( .A1(A[5]), .A2(B[5]), .ZN(n260) );
  NOR2_X1 U380 ( .A1(A[7]), .A2(B[7]), .ZN(n252) );
  NOR2_X1 U381 ( .A1(A[8]), .A2(B[8]), .ZN(n244) );
  NOR2_X1 U382 ( .A1(A[11]), .A2(B[11]), .ZN(n223) );
  NOR2_X1 U383 ( .A1(A[2]), .A2(B[2]), .ZN(n274) );
  NOR2_X1 U384 ( .A1(A[6]), .A2(B[6]), .ZN(n255) );
  NOR2_X1 U385 ( .A1(A[1]), .A2(B[1]), .ZN(n278) );
  INV_X1 U386 ( .A(n150), .ZN(n148) );
  AOI21_X1 U387 ( .B1(n150), .B2(n131), .A(n132), .ZN(n130) );
  INV_X1 U388 ( .A(n437), .ZN(n131) );
  INV_X1 U389 ( .A(n219), .ZN(n217) );
  OAI21_X1 U390 ( .B1(n246), .B2(n197), .A(n198), .ZN(n196) );
  AOI21_X1 U391 ( .B1(n218), .B2(n203), .A(n204), .ZN(n198) );
  NAND2_X1 U392 ( .A1(n217), .A2(n203), .ZN(n197) );
  OAI21_X1 U393 ( .B1(n246), .B2(n219), .A(n220), .ZN(n214) );
  INV_X1 U394 ( .A(n134), .ZN(n132) );
  INV_X1 U395 ( .A(n240), .ZN(n234) );
  INV_X1 U396 ( .A(n152), .ZN(n150) );
  INV_X1 U397 ( .A(n247), .ZN(n246) );
  AOI21_X1 U398 ( .B1(n267), .B2(n258), .A(n259), .ZN(n257) );
  AOI21_X1 U399 ( .B1(n122), .B2(n150), .A(n123), .ZN(n121) );
  NOR2_X1 U400 ( .A1(n437), .A2(n124), .ZN(n122) );
  INV_X1 U401 ( .A(n203), .ZN(n201) );
  INV_X1 U402 ( .A(n220), .ZN(n218) );
  INV_X1 U403 ( .A(n422), .ZN(n134) );
  OAI21_X1 U404 ( .B1(n246), .B2(n188), .A(n189), .ZN(n187) );
  AOI21_X1 U405 ( .B1(n190), .B2(n218), .A(n191), .ZN(n189) );
  NAND2_X1 U406 ( .A1(n190), .A2(n217), .ZN(n188) );
  NOR2_X1 U407 ( .A1(n201), .A2(n194), .ZN(n190) );
  INV_X1 U408 ( .A(n268), .ZN(n267) );
  NAND2_X1 U409 ( .A1(n239), .A2(n221), .ZN(n219) );
  INV_X1 U410 ( .A(n204), .ZN(n202) );
  INV_X1 U411 ( .A(n277), .ZN(n276) );
  INV_X1 U412 ( .A(n170), .ZN(n168) );
  INV_X1 U413 ( .A(n172), .ZN(n170) );
  INV_X1 U414 ( .A(n239), .ZN(n237) );
  NAND2_X1 U415 ( .A1(n239), .A2(n228), .ZN(n226) );
  INV_X1 U416 ( .A(n60), .ZN(n58) );
  INV_X1 U417 ( .A(n5), .ZN(n76) );
  NOR2_X1 U418 ( .A1(n244), .A2(n241), .ZN(n239) );
  OAI21_X1 U419 ( .B1(n241), .B2(n245), .A(n242), .ZN(n240) );
  AOI21_X1 U420 ( .B1(n221), .B2(n240), .A(n222), .ZN(n220) );
  OAI21_X1 U421 ( .B1(n223), .B2(n231), .A(n224), .ZN(n222) );
  OAI21_X1 U422 ( .B1(n173), .B2(n177), .A(n174), .ZN(n172) );
  OAI21_X1 U423 ( .B1(n205), .B2(n213), .A(n206), .ZN(n204) );
  NAND2_X1 U424 ( .A1(n171), .A2(n160), .ZN(n158) );
  AOI21_X1 U425 ( .B1(n168), .B2(n160), .A(n161), .ZN(n159) );
  INV_X1 U426 ( .A(n162), .ZN(n160) );
  AOI21_X1 U427 ( .B1(n269), .B2(n277), .A(n270), .ZN(n268) );
  NOR2_X1 U428 ( .A1(n274), .A2(n271), .ZN(n269) );
  OAI21_X1 U429 ( .B1(n271), .B2(n275), .A(n272), .ZN(n270) );
  OAI21_X1 U430 ( .B1(n260), .B2(n266), .A(n261), .ZN(n259) );
  OAI21_X1 U431 ( .B1(n278), .B2(n281), .A(n279), .ZN(n277) );
  NOR2_X1 U432 ( .A1(n265), .A2(n260), .ZN(n258) );
  OAI21_X1 U433 ( .B1(n433), .B2(n145), .A(n138), .ZN(n136) );
  INV_X1 U434 ( .A(n51), .ZN(n49) );
  BUF_X1 U435 ( .A(n112), .Z(n3) );
  INV_X1 U436 ( .A(n106), .ZN(n104) );
  AOI21_X1 U437 ( .B1(n150), .B2(n142), .A(n143), .ZN(n141) );
  INV_X1 U438 ( .A(n144), .ZN(n142) );
  AOI21_X1 U439 ( .B1(n240), .B2(n228), .A(n229), .ZN(n227) );
  INV_X1 U440 ( .A(n231), .ZN(n229) );
  OAI21_X1 U441 ( .B1(n268), .B2(n248), .A(n249), .ZN(n247) );
  AOI21_X1 U442 ( .B1(n250), .B2(n259), .A(n251), .ZN(n249) );
  NAND2_X1 U443 ( .A1(n258), .A2(n250), .ZN(n248) );
  NOR2_X1 U444 ( .A1(n255), .A2(n252), .ZN(n250) );
  NOR2_X1 U445 ( .A1(n230), .A2(n223), .ZN(n221) );
  OAI21_X1 U446 ( .B1(n252), .B2(n256), .A(n253), .ZN(n251) );
  AOI21_X1 U447 ( .B1(n267), .B2(n309), .A(n264), .ZN(n262) );
  INV_X1 U448 ( .A(n266), .ZN(n264) );
  OAI21_X1 U449 ( .B1(n134), .B2(n124), .A(n127), .ZN(n123) );
  OAI21_X1 U450 ( .B1(n202), .B2(n194), .A(n195), .ZN(n191) );
  OAI21_X1 U451 ( .B1(n276), .B2(n274), .A(n275), .ZN(n273) );
  OAI21_X1 U452 ( .B1(n257), .B2(n255), .A(n256), .ZN(n254) );
  OAI21_X1 U453 ( .B1(n246), .B2(n244), .A(n245), .ZN(n243) );
  OAI21_X1 U454 ( .B1(n246), .B2(n208), .A(n209), .ZN(n207) );
  AOI21_X1 U455 ( .B1(n218), .B2(n210), .A(n211), .ZN(n209) );
  NAND2_X1 U456 ( .A1(n217), .A2(n210), .ZN(n208) );
  INV_X1 U457 ( .A(n213), .ZN(n211) );
  INV_X1 U458 ( .A(n230), .ZN(n228) );
  INV_X1 U459 ( .A(n205), .ZN(n300) );
  INV_X1 U460 ( .A(n212), .ZN(n210) );
  INV_X1 U461 ( .A(n427), .ZN(n284) );
  INV_X1 U462 ( .A(n176), .ZN(n297) );
  INV_X1 U463 ( .A(n425), .ZN(n290) );
  INV_X1 U464 ( .A(n418), .ZN(n286) );
  INV_X1 U465 ( .A(n145), .ZN(n143) );
  INV_X1 U466 ( .A(n125), .ZN(n124) );
  INV_X1 U467 ( .A(n423), .ZN(n125) );
  INV_X1 U468 ( .A(n137), .ZN(n292) );
  INV_X1 U469 ( .A(n194), .ZN(n193) );
  INV_X1 U470 ( .A(n255), .ZN(n307) );
  INV_X1 U471 ( .A(n274), .ZN(n311) );
  INV_X1 U472 ( .A(n260), .ZN(n308) );
  INV_X1 U473 ( .A(n271), .ZN(n310) );
  INV_X1 U474 ( .A(n252), .ZN(n306) );
  INV_X1 U475 ( .A(n265), .ZN(n309) );
  NAND2_X1 U476 ( .A1(n228), .A2(n231), .ZN(n28) );
  NAND2_X1 U477 ( .A1(n302), .A2(n224), .ZN(n27) );
  INV_X1 U478 ( .A(n223), .ZN(n302) );
  INV_X1 U479 ( .A(n244), .ZN(n305) );
  INV_X1 U480 ( .A(n173), .ZN(n296) );
  INV_X1 U481 ( .A(n241), .ZN(n304) );
  INV_X1 U482 ( .A(n278), .ZN(n312) );
  INV_X1 U483 ( .A(n426), .ZN(n294) );
  INV_X1 U484 ( .A(n185), .ZN(n298) );
  INV_X1 U485 ( .A(n163), .ZN(n161) );
  INV_X1 U486 ( .A(n107), .ZN(n105) );
  INV_X1 U487 ( .A(n429), .ZN(n86) );
  INV_X1 U488 ( .A(n69), .ZN(n68) );
  INV_X1 U489 ( .A(n70), .ZN(n69) );
  NOR2_X1 U490 ( .A1(B[22]), .A2(A[22]), .ZN(n126) );
  NOR2_X1 U491 ( .A1(A[26]), .A2(B[26]), .ZN(n88) );
  NOR2_X1 U492 ( .A1(A[24]), .A2(B[24]), .ZN(n106) );
  NOR2_X1 U493 ( .A1(A[17]), .A2(B[17]), .ZN(n173) );
  NOR2_X1 U494 ( .A1(B[21]), .A2(A[21]), .ZN(n137) );
  NOR2_X1 U495 ( .A1(A[9]), .A2(B[9]), .ZN(n241) );
  NAND2_X1 U496 ( .A1(A[24]), .A2(B[24]), .ZN(n107) );
  NAND2_X1 U497 ( .A1(n297), .A2(n177), .ZN(n22) );
  NOR2_X1 U498 ( .A1(A[18]), .A2(B[18]), .ZN(n162) );
  NOR2_X1 U499 ( .A1(A[14]), .A2(B[14]), .ZN(n194) );
  NOR2_X1 U500 ( .A1(A[28]), .A2(B[28]), .ZN(n70) );
  NOR2_X1 U501 ( .A1(A[19]), .A2(B[19]), .ZN(n155) );
  NOR2_X1 U502 ( .A1(A[15]), .A2(B[15]), .ZN(n185) );
  AND2_X1 U503 ( .A1(n440), .A2(n281), .ZN(SUM[0]) );
  NAND2_X1 U504 ( .A1(A[4]), .A2(B[4]), .ZN(n266) );
  NAND2_X1 U505 ( .A1(A[2]), .A2(B[2]), .ZN(n275) );
  NAND2_X1 U506 ( .A1(A[6]), .A2(B[6]), .ZN(n256) );
  NAND2_X1 U507 ( .A1(A[8]), .A2(B[8]), .ZN(n245) );
  XOR2_X1 U508 ( .A(n257), .B(n32), .Z(SUM[6]) );
  NAND2_X1 U509 ( .A1(n307), .A2(n256), .ZN(n32) );
  NAND2_X1 U510 ( .A1(A[10]), .A2(B[10]), .ZN(n231) );
  NAND2_X1 U511 ( .A1(n284), .A2(n62), .ZN(n9) );
  NAND2_X1 U512 ( .A1(n417), .A2(n51), .ZN(n8) );
  NAND2_X1 U513 ( .A1(n441), .A2(n40), .ZN(n7) );
  NAND2_X1 U514 ( .A1(n286), .A2(n80), .ZN(n11) );
  NAND2_X1 U515 ( .A1(n431), .A2(n100), .ZN(n13) );
  NAND2_X1 U516 ( .A1(n429), .A2(n89), .ZN(n12) );
  NAND2_X1 U517 ( .A1(n69), .A2(n71), .ZN(n10) );
  NAND2_X1 U518 ( .A1(n290), .A2(n118), .ZN(n15) );
  XNOR2_X1 U519 ( .A(n146), .B(n18), .ZN(SUM[20]) );
  NAND2_X1 U520 ( .A1(n292), .A2(n138), .ZN(n17) );
  NAND2_X1 U521 ( .A1(n125), .A2(n127), .ZN(n16) );
  XOR2_X1 U522 ( .A(n37), .B(n281), .Z(SUM[1]) );
  NAND2_X1 U523 ( .A1(n312), .A2(n279), .ZN(n37) );
  XOR2_X1 U524 ( .A(n276), .B(n36), .Z(SUM[2]) );
  NAND2_X1 U525 ( .A1(n311), .A2(n275), .ZN(n36) );
  XNOR2_X1 U526 ( .A(n273), .B(n35), .ZN(SUM[3]) );
  NAND2_X1 U527 ( .A1(n310), .A2(n272), .ZN(n35) );
  XOR2_X1 U528 ( .A(n262), .B(n33), .Z(SUM[5]) );
  NAND2_X1 U529 ( .A1(n308), .A2(n261), .ZN(n33) );
  XNOR2_X1 U530 ( .A(n187), .B(n23), .ZN(SUM[15]) );
  NAND2_X1 U531 ( .A1(n298), .A2(n186), .ZN(n23) );
  XNOR2_X1 U532 ( .A(n157), .B(n19), .ZN(SUM[19]) );
  NAND2_X1 U533 ( .A1(n294), .A2(n156), .ZN(n19) );
  XNOR2_X1 U534 ( .A(n207), .B(n25), .ZN(SUM[13]) );
  NAND2_X1 U535 ( .A1(n300), .A2(n206), .ZN(n25) );
  XNOR2_X1 U536 ( .A(n196), .B(n24), .ZN(SUM[14]) );
  NAND2_X1 U537 ( .A1(n193), .A2(n195), .ZN(n24) );
  XNOR2_X1 U538 ( .A(n214), .B(n26), .ZN(SUM[12]) );
  NAND2_X1 U539 ( .A1(n210), .A2(n213), .ZN(n26) );
  XNOR2_X1 U540 ( .A(n225), .B(n27), .ZN(SUM[11]) );
  OAI21_X1 U541 ( .B1(n246), .B2(n226), .A(n227), .ZN(n225) );
  XNOR2_X1 U542 ( .A(n232), .B(n28), .ZN(SUM[10]) );
  OAI21_X1 U543 ( .B1(n246), .B2(n237), .A(n234), .ZN(n232) );
  XNOR2_X1 U544 ( .A(n254), .B(n31), .ZN(SUM[7]) );
  NAND2_X1 U545 ( .A1(n306), .A2(n253), .ZN(n31) );
  XOR2_X1 U546 ( .A(n246), .B(n30), .Z(SUM[8]) );
  NAND2_X1 U547 ( .A1(n305), .A2(n245), .ZN(n30) );
  XNOR2_X1 U548 ( .A(n108), .B(n14), .ZN(SUM[24]) );
  NAND2_X1 U549 ( .A1(n104), .A2(n419), .ZN(n14) );
  NAND2_X1 U550 ( .A1(A[11]), .A2(B[11]), .ZN(n224) );
  NAND2_X1 U551 ( .A1(A[12]), .A2(B[12]), .ZN(n213) );
  NAND2_X1 U552 ( .A1(A[0]), .A2(B[0]), .ZN(n281) );
  NAND2_X1 U553 ( .A1(A[5]), .A2(B[5]), .ZN(n261) );
  NAND2_X1 U554 ( .A1(A[7]), .A2(B[7]), .ZN(n253) );
  NAND2_X1 U555 ( .A1(A[3]), .A2(B[3]), .ZN(n272) );
  XNOR2_X1 U556 ( .A(n175), .B(n21), .ZN(SUM[17]) );
  NAND2_X1 U557 ( .A1(n296), .A2(n174), .ZN(n21) );
  NAND2_X1 U558 ( .A1(A[18]), .A2(B[18]), .ZN(n163) );
  NAND2_X1 U559 ( .A1(A[14]), .A2(B[14]), .ZN(n195) );
  NAND2_X1 U560 ( .A1(A[9]), .A2(B[9]), .ZN(n242) );
  XNOR2_X1 U561 ( .A(n243), .B(n29), .ZN(SUM[9]) );
  NAND2_X1 U562 ( .A1(n304), .A2(n242), .ZN(n29) );
  XNOR2_X1 U563 ( .A(n164), .B(n20), .ZN(SUM[18]) );
  NAND2_X1 U564 ( .A1(n160), .A2(n163), .ZN(n20) );
  NAND2_X1 U565 ( .A1(A[15]), .A2(B[15]), .ZN(n186) );
  NAND2_X1 U566 ( .A1(A[19]), .A2(B[19]), .ZN(n156) );
  NAND2_X1 U567 ( .A1(A[1]), .A2(B[1]), .ZN(n279) );
  NAND2_X1 U568 ( .A1(A[28]), .A2(B[28]), .ZN(n71) );
  NAND2_X1 U569 ( .A1(A[31]), .A2(B[31]), .ZN(n40) );
  XNOR2_X1 U570 ( .A(n267), .B(n34), .ZN(SUM[4]) );
  NAND2_X1 U571 ( .A1(n309), .A2(n266), .ZN(n34) );
  OR2_X1 U572 ( .A1(A[0]), .A2(B[0]), .ZN(n440) );
  OR2_X1 U573 ( .A1(A[31]), .A2(B[31]), .ZN(n441) );
  NOR2_X1 U574 ( .A1(n106), .A2(n416), .ZN(n97) );
  NOR2_X1 U575 ( .A1(B[25]), .A2(A[25]), .ZN(n99) );
  NOR2_X1 U576 ( .A1(n117), .A2(n126), .ZN(n115) );
  NAND2_X1 U577 ( .A1(A[29]), .A2(B[29]), .ZN(n62) );
  NOR2_X1 U578 ( .A1(B[29]), .A2(A[29]), .ZN(n61) );
  NOR2_X1 U579 ( .A1(n95), .A2(n86), .ZN(n84) );
  INV_X1 U580 ( .A(n95), .ZN(n93) );
  INV_X1 U581 ( .A(n97), .ZN(n95) );
  AOI21_X1 U582 ( .B1(n247), .B2(n179), .A(n180), .ZN(n178) );
  NOR2_X1 U583 ( .A1(B[23]), .A2(A[23]), .ZN(n117) );
  NAND2_X1 U584 ( .A1(n122), .A2(n149), .ZN(n120) );
  NAND2_X1 U585 ( .A1(n149), .A2(n131), .ZN(n129) );
  NAND2_X1 U586 ( .A1(n149), .A2(n142), .ZN(n140) );
  INV_X1 U587 ( .A(n149), .ZN(n147) );
  INV_X1 U588 ( .A(n151), .ZN(n149) );
  OAI21_X1 U589 ( .B1(n96), .B2(n86), .A(n89), .ZN(n85) );
  XNOR2_X1 U590 ( .A(n72), .B(n10), .ZN(SUM[28]) );
  XNOR2_X1 U591 ( .A(n101), .B(n13), .ZN(SUM[25]) );
  XNOR2_X1 U592 ( .A(n52), .B(n8), .ZN(SUM[30]) );
  XNOR2_X1 U593 ( .A(n63), .B(n9), .ZN(SUM[29]) );
  NAND2_X1 U594 ( .A1(A[17]), .A2(B[17]), .ZN(n174) );
  NAND2_X1 U595 ( .A1(A[13]), .A2(B[13]), .ZN(n206) );
  NOR2_X1 U596 ( .A1(A[13]), .A2(B[13]), .ZN(n205) );
  NOR2_X1 U597 ( .A1(n88), .A2(n79), .ZN(n77) );
  INV_X1 U598 ( .A(n171), .ZN(n169) );
  NOR2_X1 U599 ( .A1(n176), .A2(n173), .ZN(n171) );
  INV_X1 U600 ( .A(n420), .ZN(n96) );
  NAND2_X1 U601 ( .A1(A[30]), .A2(B[30]), .ZN(n51) );
  XNOR2_X1 U602 ( .A(n128), .B(n16), .ZN(SUM[22]) );
  NAND2_X1 U603 ( .A1(A[16]), .A2(B[16]), .ZN(n177) );
  NOR2_X1 U604 ( .A1(A[16]), .A2(B[16]), .ZN(n176) );
  XNOR2_X1 U605 ( .A(n139), .B(n17), .ZN(SUM[21]) );
  INV_X1 U606 ( .A(n59), .ZN(n57) );
  NOR2_X1 U607 ( .A1(n6), .A2(n57), .ZN(n55) );
  NAND2_X1 U608 ( .A1(A[26]), .A2(B[26]), .ZN(n89) );
  OAI21_X1 U609 ( .B1(n2), .B2(n109), .A(n110), .ZN(n108) );
  NOR2_X1 U610 ( .A1(B[20]), .A2(A[20]), .ZN(n144) );
  NAND2_X1 U611 ( .A1(B[20]), .A2(A[20]), .ZN(n145) );
  OAI21_X1 U612 ( .B1(n99), .B2(n107), .A(n100), .ZN(n98) );
  NAND2_X1 U613 ( .A1(B[22]), .A2(A[22]), .ZN(n127) );
  XNOR2_X1 U614 ( .A(n119), .B(n15), .ZN(SUM[23]) );
  XNOR2_X1 U615 ( .A(n90), .B(n12), .ZN(SUM[26]) );
  INV_X1 U616 ( .A(n3), .ZN(n110) );
  AOI21_X1 U617 ( .B1(n60), .B2(n417), .A(n49), .ZN(n47) );
  NAND2_X1 U618 ( .A1(B[23]), .A2(A[23]), .ZN(n118) );
  NOR2_X1 U619 ( .A1(n219), .A2(n181), .ZN(n179) );
  OAI21_X1 U620 ( .B1(n220), .B2(n181), .A(n182), .ZN(n180) );
  XNOR2_X1 U621 ( .A(n81), .B(n11), .ZN(SUM[27]) );
  INV_X1 U622 ( .A(n111), .ZN(n109) );
  AOI21_X1 U623 ( .B1(n153), .B2(n172), .A(n154), .ZN(n152) );
  NAND2_X1 U624 ( .A1(n171), .A2(n153), .ZN(n151) );
  NOR2_X1 U625 ( .A1(n162), .A2(n426), .ZN(n153) );
  AOI21_X1 U626 ( .B1(n183), .B2(n204), .A(n184), .ZN(n182) );
  NAND2_X1 U627 ( .A1(n203), .A2(n183), .ZN(n181) );
  AOI21_X1 U628 ( .B1(n136), .B2(n430), .A(n116), .ZN(n114) );
  XOR2_X1 U629 ( .A(n1), .B(n22), .Z(SUM[16]) );
  OAI21_X1 U630 ( .B1(n1), .B2(n120), .A(n121), .ZN(n119) );
  OAI21_X1 U631 ( .B1(n1), .B2(n129), .A(n130), .ZN(n128) );
  OAI21_X1 U632 ( .B1(n1), .B2(n140), .A(n141), .ZN(n139) );
  OAI21_X1 U633 ( .B1(n1), .B2(n147), .A(n148), .ZN(n146) );
  OAI21_X1 U634 ( .B1(n1), .B2(n158), .A(n159), .ZN(n157) );
  OAI21_X1 U635 ( .B1(n1), .B2(n169), .A(n170), .ZN(n164) );
  OAI21_X1 U636 ( .B1(n1), .B2(n176), .A(n177), .ZN(n175) );
  NOR2_X1 U637 ( .A1(n212), .A2(n205), .ZN(n203) );
  NAND2_X1 U638 ( .A1(n142), .A2(n145), .ZN(n18) );
  OAI21_X1 U639 ( .B1(n2), .B2(n91), .A(n92), .ZN(n90) );
  OAI21_X1 U640 ( .B1(n2), .B2(n102), .A(n103), .ZN(n101) );
  OAI21_X1 U641 ( .B1(n155), .B2(n163), .A(n156), .ZN(n154) );
  OAI21_X1 U642 ( .B1(n2), .B2(n53), .A(n54), .ZN(n52) );
  OAI21_X1 U643 ( .B1(n2), .B2(n73), .A(n74), .ZN(n72) );
  NAND2_X1 U644 ( .A1(B[25]), .A2(A[25]), .ZN(n100) );
  NAND2_X1 U645 ( .A1(n421), .A2(n44), .ZN(n42) );
  NAND2_X1 U646 ( .A1(n111), .A2(n66), .ZN(n64) );
  NAND2_X1 U647 ( .A1(n421), .A2(n84), .ZN(n82) );
  NAND2_X1 U648 ( .A1(n421), .A2(n104), .ZN(n102) );
  NAND2_X1 U649 ( .A1(n111), .A2(n55), .ZN(n53) );
  NAND2_X1 U650 ( .A1(n421), .A2(n75), .ZN(n73) );
  NAND2_X1 U651 ( .A1(n111), .A2(n93), .ZN(n91) );
  NAND2_X1 U652 ( .A1(n59), .A2(n417), .ZN(n46) );
  NOR2_X1 U653 ( .A1(n70), .A2(n61), .ZN(n59) );
  OAI21_X1 U654 ( .B1(n2), .B2(n82), .A(n83), .ZN(n81) );
  INV_X1 U655 ( .A(n6), .ZN(n75) );
  NOR2_X1 U656 ( .A1(n6), .A2(n68), .ZN(n66) );
  NOR2_X1 U657 ( .A1(n6), .A2(n46), .ZN(n44) );
  NAND2_X1 U658 ( .A1(n77), .A2(n97), .ZN(n6) );
  XNOR2_X1 U659 ( .A(n41), .B(n7), .ZN(SUM[31]) );
  OAI21_X1 U660 ( .B1(n61), .B2(n71), .A(n62), .ZN(n60) );
  NOR2_X1 U661 ( .A1(n194), .A2(n185), .ZN(n183) );
  OAI21_X1 U662 ( .B1(n185), .B2(n195), .A(n186), .ZN(n184) );
  OAI21_X1 U663 ( .B1(n2), .B2(n42), .A(n43), .ZN(n41) );
  NOR2_X1 U664 ( .A1(n151), .A2(n113), .ZN(n111) );
  OAI21_X1 U665 ( .B1(n113), .B2(n152), .A(n114), .ZN(n112) );
  NAND2_X1 U666 ( .A1(n135), .A2(n115), .ZN(n113) );
  OAI21_X1 U667 ( .B1(n2), .B2(n64), .A(n65), .ZN(n63) );
  AOI21_X1 U668 ( .B1(n3), .B2(n104), .A(n105), .ZN(n103) );
  AOI21_X1 U669 ( .B1(n438), .B2(n93), .A(n420), .ZN(n92) );
  AOI21_X1 U670 ( .B1(n3), .B2(n75), .A(n76), .ZN(n74) );
  AOI21_X1 U671 ( .B1(n438), .B2(n84), .A(n85), .ZN(n83) );
  AOI21_X1 U672 ( .B1(n438), .B2(n44), .A(n45), .ZN(n43) );
  AOI21_X1 U673 ( .B1(n3), .B2(n55), .A(n56), .ZN(n54) );
  AOI21_X1 U674 ( .B1(n438), .B2(n66), .A(n67), .ZN(n65) );
  OAI21_X1 U675 ( .B1(n5), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U676 ( .B1(n5), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U677 ( .B1(n5), .B2(n68), .A(n71), .ZN(n67) );
  OAI21_X1 U678 ( .B1(n436), .B2(n89), .A(n80), .ZN(n78) );
  NAND2_X1 U679 ( .A1(A[27]), .A2(B[27]), .ZN(n80) );
  NOR2_X1 U680 ( .A1(A[27]), .A2(B[27]), .ZN(n79) );
  NOR2_X1 U681 ( .A1(n137), .A2(n144), .ZN(n135) );
  NAND2_X1 U682 ( .A1(B[21]), .A2(A[21]), .ZN(n138) );
  OAI21_X1 U683 ( .B1(n432), .B2(n127), .A(n118), .ZN(n116) );
endmodule


module datapath_DW01_add_9 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n40, n41, n42, n43, n44, n45, n46,
         n47, n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n134, n135, n137, n138, n139, n140, n141,
         n143, n144, n145, n146, n147, n149, n150, n151, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n193, n194, n195, n196, n197, n198, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n234, n237, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n281, n284, n286, n287, n288, n290, n292, n293, n294, n296,
         n297, n298, n300, n302, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n416, n417, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444;

  CLKBUF_X1 U349 ( .A(n61), .Z(n416) );
  BUF_X1 U350 ( .A(n432), .Z(n427) );
  NOR2_X2 U351 ( .A1(B[19]), .A2(A[19]), .ZN(n155) );
  OR2_X1 U352 ( .A1(A[30]), .A2(B[30]), .ZN(n417) );
  AND2_X1 U353 ( .A1(n420), .A2(n281), .ZN(SUM[0]) );
  NOR2_X1 U354 ( .A1(A[26]), .A2(n436), .ZN(n419) );
  BUF_X1 U355 ( .A(n435), .Z(n437) );
  OR2_X1 U356 ( .A1(A[0]), .A2(B[0]), .ZN(n420) );
  AOI21_X1 U357 ( .B1(n77), .B2(n98), .A(n78), .ZN(n421) );
  AOI21_X1 U358 ( .B1(n77), .B2(n98), .A(n78), .ZN(n5) );
  BUF_X1 U359 ( .A(n112), .Z(n422) );
  CLKBUF_X1 U360 ( .A(n112), .Z(n3) );
  BUF_X1 U361 ( .A(n428), .Z(n423) );
  CLKBUF_X1 U362 ( .A(n430), .Z(n424) );
  BUF_X1 U363 ( .A(n178), .Z(n425) );
  BUF_X1 U364 ( .A(n178), .Z(n426) );
  AOI21_X2 U365 ( .B1(n247), .B2(n179), .A(n180), .ZN(n178) );
  NOR2_X1 U366 ( .A1(n151), .A2(n113), .ZN(n428) );
  NOR2_X1 U367 ( .A1(n88), .A2(n430), .ZN(n429) );
  NOR2_X1 U368 ( .A1(B[27]), .A2(A[27]), .ZN(n430) );
  NOR2_X1 U369 ( .A1(B[27]), .A2(A[27]), .ZN(n79) );
  BUF_X1 U370 ( .A(n112), .Z(n431) );
  AOI21_X1 U371 ( .B1(n153), .B2(n172), .A(n154), .ZN(n432) );
  INV_X1 U372 ( .A(n143), .ZN(n433) );
  CLKBUF_X1 U373 ( .A(n137), .Z(n434) );
  OAI21_X1 U374 ( .B1(n443), .B2(n145), .A(n138), .ZN(n435) );
  CLKBUF_X1 U375 ( .A(B[26]), .Z(n436) );
  CLKBUF_X1 U376 ( .A(n117), .Z(n438) );
  NOR2_X1 U377 ( .A1(B[22]), .A2(A[22]), .ZN(n126) );
  NOR2_X1 U378 ( .A1(B[26]), .A2(A[26]), .ZN(n88) );
  NOR2_X1 U379 ( .A1(B[25]), .A2(A[25]), .ZN(n439) );
  NOR2_X1 U380 ( .A1(n117), .A2(n126), .ZN(n440) );
  OR2_X1 U381 ( .A1(n144), .A2(n434), .ZN(n441) );
  NOR2_X1 U382 ( .A1(B[23]), .A2(A[23]), .ZN(n442) );
  NOR2_X1 U383 ( .A1(A[25]), .A2(B[25]), .ZN(n99) );
  NOR2_X1 U384 ( .A1(A[21]), .A2(B[21]), .ZN(n443) );
  NOR2_X1 U385 ( .A1(A[10]), .A2(B[10]), .ZN(n230) );
  NOR2_X1 U386 ( .A1(A[12]), .A2(B[12]), .ZN(n212) );
  NOR2_X1 U387 ( .A1(A[4]), .A2(B[4]), .ZN(n265) );
  NOR2_X1 U388 ( .A1(A[3]), .A2(B[3]), .ZN(n271) );
  NOR2_X1 U389 ( .A1(A[5]), .A2(B[5]), .ZN(n260) );
  NOR2_X1 U390 ( .A1(A[9]), .A2(B[9]), .ZN(n241) );
  NOR2_X1 U391 ( .A1(A[7]), .A2(B[7]), .ZN(n252) );
  NOR2_X1 U392 ( .A1(A[8]), .A2(B[8]), .ZN(n244) );
  NOR2_X1 U393 ( .A1(A[6]), .A2(B[6]), .ZN(n255) );
  NOR2_X1 U394 ( .A1(A[2]), .A2(B[2]), .ZN(n274) );
  NOR2_X1 U395 ( .A1(A[1]), .A2(B[1]), .ZN(n278) );
  NAND2_X1 U396 ( .A1(A[24]), .A2(B[24]), .ZN(n107) );
  OR2_X1 U397 ( .A1(A[31]), .A2(B[31]), .ZN(n444) );
  INV_X1 U398 ( .A(n151), .ZN(n149) );
  INV_X1 U399 ( .A(n149), .ZN(n147) );
  NAND2_X1 U400 ( .A1(n149), .A2(n131), .ZN(n129) );
  AOI21_X1 U401 ( .B1(n150), .B2(n131), .A(n437), .ZN(n130) );
  INV_X1 U402 ( .A(n441), .ZN(n131) );
  INV_X1 U403 ( .A(n219), .ZN(n217) );
  OAI21_X1 U404 ( .B1(n246), .B2(n237), .A(n234), .ZN(n232) );
  INV_X1 U405 ( .A(n240), .ZN(n234) );
  OAI21_X1 U406 ( .B1(n246), .B2(n219), .A(n220), .ZN(n214) );
  BUF_X1 U407 ( .A(n178), .Z(n2) );
  BUF_X1 U408 ( .A(n428), .Z(n4) );
  BUF_X1 U409 ( .A(n178), .Z(n1) );
  OAI21_X1 U410 ( .B1(n246), .B2(n197), .A(n198), .ZN(n196) );
  AOI21_X1 U411 ( .B1(n218), .B2(n203), .A(n204), .ZN(n198) );
  NAND2_X1 U412 ( .A1(n217), .A2(n203), .ZN(n197) );
  INV_X1 U413 ( .A(n96), .ZN(n94) );
  INV_X1 U414 ( .A(n427), .ZN(n150) );
  INV_X1 U415 ( .A(n247), .ZN(n246) );
  NAND2_X1 U416 ( .A1(n122), .A2(n149), .ZN(n120) );
  AOI21_X1 U417 ( .B1(n122), .B2(n150), .A(n123), .ZN(n121) );
  NOR2_X1 U418 ( .A1(n441), .A2(n124), .ZN(n122) );
  AOI21_X1 U419 ( .B1(n267), .B2(n258), .A(n259), .ZN(n257) );
  NOR2_X1 U420 ( .A1(n201), .A2(n194), .ZN(n190) );
  INV_X1 U421 ( .A(n6), .ZN(n75) );
  INV_X1 U422 ( .A(n220), .ZN(n218) );
  NAND2_X1 U423 ( .A1(n97), .A2(n429), .ZN(n6) );
  INV_X1 U424 ( .A(n268), .ZN(n267) );
  INV_X1 U425 ( .A(n203), .ZN(n201) );
  NAND2_X1 U426 ( .A1(n239), .A2(n221), .ZN(n219) );
  INV_X1 U427 ( .A(n204), .ZN(n202) );
  INV_X1 U428 ( .A(n170), .ZN(n168) );
  INV_X1 U429 ( .A(n172), .ZN(n170) );
  OAI21_X1 U430 ( .B1(n2), .B2(n109), .A(n110), .ZN(n108) );
  INV_X1 U431 ( .A(n111), .ZN(n109) );
  INV_X1 U432 ( .A(n277), .ZN(n276) );
  INV_X1 U433 ( .A(n171), .ZN(n169) );
  INV_X1 U434 ( .A(n239), .ZN(n237) );
  INV_X1 U435 ( .A(n59), .ZN(n57) );
  INV_X1 U436 ( .A(n421), .ZN(n76) );
  NOR2_X1 U437 ( .A1(n230), .A2(n223), .ZN(n221) );
  OAI21_X1 U438 ( .B1(n205), .B2(n213), .A(n206), .ZN(n204) );
  AOI21_X1 U439 ( .B1(n168), .B2(n160), .A(n161), .ZN(n159) );
  NAND2_X1 U440 ( .A1(n171), .A2(n160), .ZN(n158) );
  NAND2_X1 U441 ( .A1(n149), .A2(n293), .ZN(n140) );
  AOI21_X1 U442 ( .B1(n150), .B2(n293), .A(n143), .ZN(n141) );
  AOI21_X1 U443 ( .B1(n269), .B2(n277), .A(n270), .ZN(n268) );
  OAI21_X1 U444 ( .B1(n271), .B2(n275), .A(n272), .ZN(n270) );
  NOR2_X1 U445 ( .A1(n274), .A2(n271), .ZN(n269) );
  NOR2_X1 U446 ( .A1(n176), .A2(n173), .ZN(n171) );
  OAI21_X1 U447 ( .B1(n241), .B2(n245), .A(n242), .ZN(n240) );
  OAI21_X1 U448 ( .B1(n260), .B2(n266), .A(n261), .ZN(n259) );
  OAI21_X1 U449 ( .B1(n278), .B2(n281), .A(n279), .ZN(n277) );
  OAI21_X1 U450 ( .B1(n268), .B2(n248), .A(n249), .ZN(n247) );
  AOI21_X1 U451 ( .B1(n250), .B2(n259), .A(n251), .ZN(n249) );
  NAND2_X1 U452 ( .A1(n258), .A2(n250), .ZN(n248) );
  OAI21_X1 U453 ( .B1(n252), .B2(n256), .A(n253), .ZN(n251) );
  NOR2_X1 U454 ( .A1(n88), .A2(n430), .ZN(n77) );
  NOR2_X1 U455 ( .A1(n265), .A2(n260), .ZN(n258) );
  NOR2_X1 U456 ( .A1(n255), .A2(n252), .ZN(n250) );
  AOI21_X1 U457 ( .B1(n221), .B2(n240), .A(n222), .ZN(n220) );
  NOR2_X1 U458 ( .A1(n244), .A2(n241), .ZN(n239) );
  INV_X1 U459 ( .A(n51), .ZN(n49) );
  AOI21_X1 U460 ( .B1(n267), .B2(n309), .A(n264), .ZN(n262) );
  INV_X1 U461 ( .A(n266), .ZN(n264) );
  OAI21_X1 U462 ( .B1(n134), .B2(n124), .A(n127), .ZN(n123) );
  INV_X1 U463 ( .A(n125), .ZN(n124) );
  OAI21_X1 U464 ( .B1(n246), .B2(n244), .A(n245), .ZN(n243) );
  OAI21_X1 U465 ( .B1(n257), .B2(n255), .A(n256), .ZN(n254) );
  OAI21_X1 U466 ( .B1(n276), .B2(n274), .A(n275), .ZN(n273) );
  OAI21_X1 U467 ( .B1(n246), .B2(n188), .A(n189), .ZN(n187) );
  AOI21_X1 U468 ( .B1(n190), .B2(n218), .A(n191), .ZN(n189) );
  NAND2_X1 U469 ( .A1(n190), .A2(n217), .ZN(n188) );
  OAI21_X1 U470 ( .B1(n202), .B2(n194), .A(n195), .ZN(n191) );
  OAI21_X1 U471 ( .B1(n246), .B2(n208), .A(n209), .ZN(n207) );
  NAND2_X1 U472 ( .A1(n217), .A2(n210), .ZN(n208) );
  AOI21_X1 U473 ( .B1(n218), .B2(n210), .A(n211), .ZN(n209) );
  INV_X1 U474 ( .A(n212), .ZN(n210) );
  OAI21_X1 U475 ( .B1(n246), .B2(n226), .A(n227), .ZN(n225) );
  NAND2_X1 U476 ( .A1(n239), .A2(n228), .ZN(n226) );
  AOI21_X1 U477 ( .B1(n240), .B2(n228), .A(n229), .ZN(n227) );
  INV_X1 U478 ( .A(n230), .ZN(n228) );
  INV_X1 U479 ( .A(n434), .ZN(n292) );
  INV_X1 U480 ( .A(n163), .ZN(n161) );
  INV_X1 U481 ( .A(n194), .ZN(n193) );
  NAND2_X1 U482 ( .A1(n417), .A2(n51), .ZN(n8) );
  NAND2_X1 U483 ( .A1(n309), .A2(n266), .ZN(n34) );
  INV_X1 U484 ( .A(n265), .ZN(n309) );
  NAND2_X1 U485 ( .A1(n310), .A2(n272), .ZN(n35) );
  INV_X1 U486 ( .A(n271), .ZN(n310) );
  NAND2_X1 U487 ( .A1(n307), .A2(n256), .ZN(n32) );
  INV_X1 U488 ( .A(n255), .ZN(n307) );
  NAND2_X1 U489 ( .A1(n305), .A2(n245), .ZN(n30) );
  INV_X1 U490 ( .A(n244), .ZN(n305) );
  INV_X1 U491 ( .A(n88), .ZN(n287) );
  NAND2_X1 U492 ( .A1(n306), .A2(n253), .ZN(n31) );
  INV_X1 U493 ( .A(n252), .ZN(n306) );
  NAND2_X1 U494 ( .A1(n304), .A2(n242), .ZN(n29) );
  INV_X1 U495 ( .A(n241), .ZN(n304) );
  NAND2_X1 U496 ( .A1(n210), .A2(n213), .ZN(n26) );
  NAND2_X1 U497 ( .A1(n308), .A2(n261), .ZN(n33) );
  INV_X1 U498 ( .A(n260), .ZN(n308) );
  NAND2_X1 U499 ( .A1(n311), .A2(n275), .ZN(n36) );
  INV_X1 U500 ( .A(n274), .ZN(n311) );
  NAND2_X1 U501 ( .A1(n228), .A2(n231), .ZN(n28) );
  NAND2_X1 U502 ( .A1(n193), .A2(n195), .ZN(n24) );
  INV_X1 U503 ( .A(n424), .ZN(n286) );
  NAND2_X1 U504 ( .A1(n300), .A2(n206), .ZN(n25) );
  INV_X1 U505 ( .A(n205), .ZN(n300) );
  NAND2_X1 U506 ( .A1(n298), .A2(n186), .ZN(n23) );
  INV_X1 U507 ( .A(n185), .ZN(n298) );
  NAND2_X1 U508 ( .A1(n312), .A2(n279), .ZN(n37) );
  INV_X1 U509 ( .A(n278), .ZN(n312) );
  INV_X1 U510 ( .A(n145), .ZN(n143) );
  INV_X1 U511 ( .A(n155), .ZN(n294) );
  NAND2_X1 U512 ( .A1(n302), .A2(n224), .ZN(n27) );
  INV_X1 U513 ( .A(n213), .ZN(n211) );
  INV_X1 U514 ( .A(n231), .ZN(n229) );
  INV_X1 U515 ( .A(n439), .ZN(n288) );
  NAND2_X1 U516 ( .A1(n104), .A2(n107), .ZN(n14) );
  NAND2_X1 U517 ( .A1(n69), .A2(n71), .ZN(n10) );
  NAND2_X1 U518 ( .A1(n297), .A2(n177), .ZN(n22) );
  INV_X1 U519 ( .A(n69), .ZN(n68) );
  INV_X1 U520 ( .A(n70), .ZN(n69) );
  INV_X1 U521 ( .A(n107), .ZN(n105) );
  NAND2_X1 U522 ( .A1(n444), .A2(n40), .ZN(n7) );
  NAND2_X1 U523 ( .A1(A[31]), .A2(B[31]), .ZN(n40) );
  NOR2_X1 U524 ( .A1(A[28]), .A2(B[28]), .ZN(n70) );
  NOR2_X1 U525 ( .A1(A[17]), .A2(B[17]), .ZN(n173) );
  NAND2_X1 U526 ( .A1(A[20]), .A2(B[20]), .ZN(n145) );
  NAND2_X1 U527 ( .A1(A[22]), .A2(B[22]), .ZN(n127) );
  NOR2_X1 U528 ( .A1(A[18]), .A2(B[18]), .ZN(n162) );
  NOR2_X1 U529 ( .A1(B[23]), .A2(A[23]), .ZN(n117) );
  NOR2_X1 U530 ( .A1(A[14]), .A2(B[14]), .ZN(n194) );
  NOR2_X1 U531 ( .A1(A[13]), .A2(B[13]), .ZN(n205) );
  NOR2_X1 U532 ( .A1(A[15]), .A2(B[15]), .ZN(n185) );
  NAND2_X1 U533 ( .A1(A[4]), .A2(B[4]), .ZN(n266) );
  NAND2_X1 U534 ( .A1(A[6]), .A2(B[6]), .ZN(n256) );
  NAND2_X1 U535 ( .A1(A[8]), .A2(B[8]), .ZN(n245) );
  NAND2_X1 U536 ( .A1(B[26]), .A2(A[26]), .ZN(n89) );
  NAND2_X1 U537 ( .A1(A[2]), .A2(B[2]), .ZN(n275) );
  NAND2_X1 U538 ( .A1(A[5]), .A2(B[5]), .ZN(n261) );
  NAND2_X1 U539 ( .A1(A[9]), .A2(B[9]), .ZN(n242) );
  NAND2_X1 U540 ( .A1(A[7]), .A2(B[7]), .ZN(n253) );
  NAND2_X1 U541 ( .A1(A[12]), .A2(B[12]), .ZN(n213) );
  NAND2_X1 U542 ( .A1(A[0]), .A2(B[0]), .ZN(n281) );
  NAND2_X1 U543 ( .A1(A[19]), .A2(B[19]), .ZN(n156) );
  NAND2_X1 U544 ( .A1(A[10]), .A2(B[10]), .ZN(n231) );
  NAND2_X1 U545 ( .A1(A[14]), .A2(B[14]), .ZN(n195) );
  NAND2_X1 U546 ( .A1(A[1]), .A2(B[1]), .ZN(n279) );
  NAND2_X1 U547 ( .A1(A[3]), .A2(B[3]), .ZN(n272) );
  NAND2_X1 U548 ( .A1(A[13]), .A2(B[13]), .ZN(n206) );
  NAND2_X1 U549 ( .A1(A[15]), .A2(B[15]), .ZN(n186) );
  NAND2_X1 U550 ( .A1(A[28]), .A2(B[28]), .ZN(n71) );
  NAND2_X1 U551 ( .A1(A[16]), .A2(B[16]), .ZN(n177) );
  NAND2_X1 U552 ( .A1(A[11]), .A2(B[11]), .ZN(n224) );
  XNOR2_X1 U553 ( .A(n119), .B(n15), .ZN(SUM[23]) );
  NAND2_X1 U554 ( .A1(n290), .A2(n118), .ZN(n15) );
  XNOR2_X1 U555 ( .A(n175), .B(n21), .ZN(SUM[17]) );
  NAND2_X1 U556 ( .A1(n296), .A2(n174), .ZN(n21) );
  XNOR2_X1 U557 ( .A(n157), .B(n19), .ZN(SUM[19]) );
  NAND2_X1 U558 ( .A1(n294), .A2(n156), .ZN(n19) );
  XNOR2_X1 U559 ( .A(n146), .B(n18), .ZN(SUM[20]) );
  NAND2_X1 U560 ( .A1(n293), .A2(n433), .ZN(n18) );
  XNOR2_X1 U561 ( .A(n139), .B(n17), .ZN(SUM[21]) );
  NAND2_X1 U562 ( .A1(n292), .A2(n138), .ZN(n17) );
  XNOR2_X1 U563 ( .A(n164), .B(n20), .ZN(SUM[18]) );
  NAND2_X1 U564 ( .A1(n160), .A2(n163), .ZN(n20) );
  XNOR2_X1 U565 ( .A(n128), .B(n16), .ZN(SUM[22]) );
  NAND2_X1 U566 ( .A1(n125), .A2(n127), .ZN(n16) );
  NAND2_X1 U567 ( .A1(n287), .A2(n89), .ZN(n12) );
  NAND2_X1 U568 ( .A1(n286), .A2(n80), .ZN(n11) );
  XNOR2_X1 U569 ( .A(n273), .B(n35), .ZN(SUM[3]) );
  XNOR2_X1 U570 ( .A(n267), .B(n34), .ZN(SUM[4]) );
  XOR2_X1 U571 ( .A(n262), .B(n33), .Z(SUM[5]) );
  XNOR2_X1 U572 ( .A(n187), .B(n23), .ZN(SUM[15]) );
  XNOR2_X1 U573 ( .A(n196), .B(n24), .ZN(SUM[14]) );
  XNOR2_X1 U574 ( .A(n207), .B(n25), .ZN(SUM[13]) );
  XNOR2_X1 U575 ( .A(n243), .B(n29), .ZN(SUM[9]) );
  XNOR2_X1 U576 ( .A(n232), .B(n28), .ZN(SUM[10]) );
  XNOR2_X1 U577 ( .A(n225), .B(n27), .ZN(SUM[11]) );
  XNOR2_X1 U578 ( .A(n214), .B(n26), .ZN(SUM[12]) );
  XOR2_X1 U579 ( .A(n257), .B(n32), .Z(SUM[6]) );
  XNOR2_X1 U580 ( .A(n254), .B(n31), .ZN(SUM[7]) );
  XOR2_X1 U581 ( .A(n37), .B(n281), .Z(SUM[1]) );
  XOR2_X1 U582 ( .A(n276), .B(n36), .Z(SUM[2]) );
  XOR2_X1 U583 ( .A(n246), .B(n30), .Z(SUM[8]) );
  INV_X1 U584 ( .A(n106), .ZN(n104) );
  NOR2_X1 U585 ( .A1(n106), .A2(n439), .ZN(n97) );
  NOR2_X1 U586 ( .A1(A[24]), .A2(B[24]), .ZN(n106) );
  INV_X1 U587 ( .A(n126), .ZN(n125) );
  INV_X1 U588 ( .A(n176), .ZN(n297) );
  NOR2_X1 U589 ( .A1(A[16]), .A2(B[16]), .ZN(n176) );
  INV_X1 U590 ( .A(n173), .ZN(n296) );
  INV_X1 U591 ( .A(n223), .ZN(n302) );
  OAI21_X1 U592 ( .B1(n223), .B2(n231), .A(n224), .ZN(n222) );
  NOR2_X1 U593 ( .A1(A[11]), .A2(B[11]), .ZN(n223) );
  INV_X1 U594 ( .A(n162), .ZN(n160) );
  NOR2_X1 U595 ( .A1(n162), .A2(n155), .ZN(n153) );
  INV_X1 U596 ( .A(n438), .ZN(n290) );
  NOR2_X1 U597 ( .A1(A[29]), .A2(B[29]), .ZN(n61) );
  NAND2_X1 U598 ( .A1(A[29]), .A2(B[29]), .ZN(n62) );
  NAND2_X1 U599 ( .A1(n284), .A2(n62), .ZN(n9) );
  INV_X1 U600 ( .A(n416), .ZN(n284) );
  NAND2_X1 U601 ( .A1(A[30]), .A2(B[30]), .ZN(n51) );
  INV_X1 U602 ( .A(n437), .ZN(n134) );
  INV_X1 U603 ( .A(n431), .ZN(n110) );
  INV_X1 U604 ( .A(n144), .ZN(n293) );
  OAI21_X1 U605 ( .B1(n173), .B2(n177), .A(n174), .ZN(n172) );
  INV_X1 U606 ( .A(n95), .ZN(n93) );
  NOR2_X1 U607 ( .A1(n95), .A2(n419), .ZN(n84) );
  INV_X1 U608 ( .A(n97), .ZN(n95) );
  NAND2_X1 U609 ( .A1(A[18]), .A2(B[18]), .ZN(n163) );
  OAI21_X1 U610 ( .B1(n96), .B2(n419), .A(n89), .ZN(n85) );
  XNOR2_X1 U611 ( .A(n72), .B(n10), .ZN(SUM[28]) );
  NAND2_X1 U612 ( .A1(n288), .A2(n100), .ZN(n13) );
  NAND2_X1 U613 ( .A1(A[17]), .A2(B[17]), .ZN(n174) );
  NOR2_X1 U614 ( .A1(B[20]), .A2(A[20]), .ZN(n144) );
  XNOR2_X1 U615 ( .A(n90), .B(n12), .ZN(SUM[26]) );
  XNOR2_X1 U616 ( .A(n101), .B(n13), .ZN(SUM[25]) );
  XNOR2_X1 U617 ( .A(n81), .B(n11), .ZN(SUM[27]) );
  NOR2_X1 U618 ( .A1(n219), .A2(n181), .ZN(n179) );
  OAI21_X1 U619 ( .B1(n220), .B2(n181), .A(n182), .ZN(n180) );
  AOI21_X1 U620 ( .B1(n60), .B2(n417), .A(n49), .ZN(n47) );
  INV_X1 U621 ( .A(n60), .ZN(n58) );
  OAI21_X1 U622 ( .B1(n53), .B2(n2), .A(n54), .ZN(n52) );
  OAI21_X1 U623 ( .B1(n2), .B2(n64), .A(n65), .ZN(n63) );
  NAND2_X1 U624 ( .A1(n171), .A2(n153), .ZN(n151) );
  XNOR2_X1 U625 ( .A(n108), .B(n14), .ZN(SUM[24]) );
  NOR2_X1 U626 ( .A1(n6), .A2(n46), .ZN(n44) );
  NAND2_X1 U627 ( .A1(B[25]), .A2(A[25]), .ZN(n100) );
  AOI21_X1 U628 ( .B1(n183), .B2(n204), .A(n184), .ZN(n182) );
  NAND2_X1 U629 ( .A1(n203), .A2(n183), .ZN(n181) );
  OAI21_X1 U630 ( .B1(n2), .B2(n102), .A(n103), .ZN(n101) );
  XOR2_X1 U631 ( .A(n1), .B(n22), .Z(SUM[16]) );
  OAI21_X1 U632 ( .B1(n425), .B2(n120), .A(n121), .ZN(n119) );
  OAI21_X1 U633 ( .B1(n426), .B2(n129), .A(n130), .ZN(n128) );
  OAI21_X1 U634 ( .B1(n425), .B2(n140), .A(n141), .ZN(n139) );
  OAI21_X1 U635 ( .B1(n426), .B2(n147), .A(n427), .ZN(n146) );
  OAI21_X1 U636 ( .B1(n1), .B2(n158), .A(n159), .ZN(n157) );
  OAI21_X1 U637 ( .B1(n425), .B2(n169), .A(n170), .ZN(n164) );
  OAI21_X1 U638 ( .B1(n426), .B2(n176), .A(n177), .ZN(n175) );
  NOR2_X1 U639 ( .A1(n212), .A2(n205), .ZN(n203) );
  NAND2_X1 U640 ( .A1(B[27]), .A2(A[27]), .ZN(n80) );
  XNOR2_X1 U641 ( .A(n41), .B(n7), .ZN(SUM[31]) );
  INV_X1 U642 ( .A(n98), .ZN(n96) );
  NAND2_X1 U643 ( .A1(n59), .A2(n417), .ZN(n46) );
  NOR2_X1 U644 ( .A1(n70), .A2(n61), .ZN(n59) );
  XNOR2_X1 U645 ( .A(n52), .B(n8), .ZN(SUM[30]) );
  XNOR2_X1 U646 ( .A(n63), .B(n9), .ZN(SUM[29]) );
  OAI21_X1 U647 ( .B1(n99), .B2(n107), .A(n100), .ZN(n98) );
  OAI21_X1 U648 ( .B1(n1), .B2(n73), .A(n74), .ZN(n72) );
  OAI21_X1 U649 ( .B1(n426), .B2(n91), .A(n92), .ZN(n90) );
  OAI21_X1 U650 ( .B1(n155), .B2(n163), .A(n156), .ZN(n154) );
  OAI21_X1 U651 ( .B1(n425), .B2(n82), .A(n83), .ZN(n81) );
  OAI21_X1 U652 ( .B1(n1), .B2(n42), .A(n43), .ZN(n41) );
  OAI21_X1 U653 ( .B1(n61), .B2(n71), .A(n62), .ZN(n60) );
  NOR2_X1 U654 ( .A1(n6), .A2(n57), .ZN(n55) );
  NOR2_X1 U655 ( .A1(n6), .A2(n68), .ZN(n66) );
  NOR2_X1 U656 ( .A1(n194), .A2(n185), .ZN(n183) );
  OAI21_X1 U657 ( .B1(n185), .B2(n195), .A(n186), .ZN(n184) );
  NAND2_X1 U658 ( .A1(n423), .A2(n75), .ZN(n73) );
  NAND2_X1 U659 ( .A1(n4), .A2(n44), .ZN(n42) );
  NAND2_X1 U660 ( .A1(n55), .A2(n423), .ZN(n53) );
  NAND2_X1 U661 ( .A1(n111), .A2(n66), .ZN(n64) );
  NAND2_X1 U662 ( .A1(n111), .A2(n84), .ZN(n82) );
  NAND2_X1 U663 ( .A1(n4), .A2(n93), .ZN(n91) );
  NAND2_X1 U664 ( .A1(n111), .A2(n104), .ZN(n102) );
  OAI21_X1 U665 ( .B1(n113), .B2(n432), .A(n114), .ZN(n112) );
  NOR2_X1 U666 ( .A1(n151), .A2(n113), .ZN(n111) );
  AOI21_X1 U667 ( .B1(n422), .B2(n93), .A(n94), .ZN(n92) );
  AOI21_X1 U668 ( .B1(n422), .B2(n104), .A(n105), .ZN(n103) );
  AOI21_X1 U669 ( .B1(n431), .B2(n75), .A(n76), .ZN(n74) );
  AOI21_X1 U670 ( .B1(n422), .B2(n84), .A(n85), .ZN(n83) );
  AOI21_X1 U671 ( .B1(n3), .B2(n44), .A(n45), .ZN(n43) );
  AOI21_X1 U672 ( .B1(n3), .B2(n55), .A(n56), .ZN(n54) );
  AOI21_X1 U673 ( .B1(n431), .B2(n66), .A(n67), .ZN(n65) );
  NAND2_X1 U674 ( .A1(n440), .A2(n135), .ZN(n113) );
  NOR2_X1 U675 ( .A1(n144), .A2(n137), .ZN(n135) );
  OAI21_X1 U676 ( .B1(n5), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U677 ( .B1(n5), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U678 ( .B1(n421), .B2(n68), .A(n71), .ZN(n67) );
  OAI21_X1 U679 ( .B1(n79), .B2(n89), .A(n80), .ZN(n78) );
  OAI21_X1 U680 ( .B1(n442), .B2(n127), .A(n118), .ZN(n116) );
  NAND2_X1 U681 ( .A1(B[23]), .A2(A[23]), .ZN(n118) );
  NOR2_X1 U682 ( .A1(n117), .A2(n126), .ZN(n115) );
  AOI21_X1 U683 ( .B1(n115), .B2(n435), .A(n116), .ZN(n114) );
  NAND2_X1 U684 ( .A1(B[21]), .A2(A[21]), .ZN(n138) );
  NOR2_X1 U685 ( .A1(B[21]), .A2(A[21]), .ZN(n137) );
endmodule


module datapath_DW01_add_10 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n40, n41, n42, n43, n44, n45, n46,
         n47, n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n193, n194, n195, n196, n197, n198,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n234, n237, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n281, n284, n286, n288, n290,
         n292, n294, n296, n297, n298, n300, n302, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n438, n439, n440;

  CLKBUF_X1 U349 ( .A(n427), .Z(n418) );
  BUF_X2 U350 ( .A(n111), .Z(n4) );
  OR2_X1 U351 ( .A1(A[30]), .A2(B[30]), .ZN(n416) );
  OR2_X1 U352 ( .A1(n144), .A2(n418), .ZN(n417) );
  CLKBUF_X3 U353 ( .A(n178), .Z(n1) );
  CLKBUF_X3 U354 ( .A(n178), .Z(n2) );
  CLKBUF_X1 U355 ( .A(n425), .Z(n419) );
  CLKBUF_X1 U356 ( .A(n127), .Z(n420) );
  OR2_X1 U357 ( .A1(n106), .A2(n99), .ZN(n421) );
  CLKBUF_X1 U358 ( .A(n79), .Z(n422) );
  CLKBUF_X1 U359 ( .A(n61), .Z(n423) );
  CLKBUF_X1 U360 ( .A(n136), .Z(n424) );
  NOR2_X1 U361 ( .A1(A[19]), .A2(B[19]), .ZN(n425) );
  CLKBUF_X1 U362 ( .A(n144), .Z(n426) );
  NOR2_X1 U363 ( .A1(B[21]), .A2(A[21]), .ZN(n427) );
  NOR2_X1 U364 ( .A1(A[27]), .A2(B[27]), .ZN(n428) );
  NOR2_X1 U365 ( .A1(B[25]), .A2(A[25]), .ZN(n429) );
  NOR2_X1 U366 ( .A1(B[25]), .A2(A[25]), .ZN(n99) );
  NOR2_X1 U367 ( .A1(n431), .A2(n126), .ZN(n430) );
  NOR2_X1 U368 ( .A1(B[23]), .A2(A[23]), .ZN(n431) );
  CLKBUF_X1 U369 ( .A(n118), .Z(n432) );
  CLKBUF_X1 U370 ( .A(n112), .Z(n433) );
  BUF_X1 U371 ( .A(n112), .Z(n434) );
  CLKBUF_X1 U372 ( .A(n431), .Z(n435) );
  BUF_X1 U373 ( .A(n111), .Z(n436) );
  NOR2_X1 U374 ( .A1(A[10]), .A2(B[10]), .ZN(n230) );
  NOR2_X1 U375 ( .A1(A[4]), .A2(B[4]), .ZN(n265) );
  NOR2_X1 U376 ( .A1(A[12]), .A2(B[12]), .ZN(n212) );
  NOR2_X1 U377 ( .A1(A[3]), .A2(B[3]), .ZN(n271) );
  NOR2_X1 U378 ( .A1(A[5]), .A2(B[5]), .ZN(n260) );
  NOR2_X1 U379 ( .A1(A[7]), .A2(B[7]), .ZN(n252) );
  NOR2_X1 U380 ( .A1(A[8]), .A2(B[8]), .ZN(n244) );
  NOR2_X1 U381 ( .A1(A[2]), .A2(B[2]), .ZN(n274) );
  NOR2_X1 U382 ( .A1(A[6]), .A2(B[6]), .ZN(n255) );
  NOR2_X1 U383 ( .A1(A[1]), .A2(B[1]), .ZN(n278) );
  NAND2_X1 U384 ( .A1(n149), .A2(n131), .ZN(n129) );
  AOI21_X1 U385 ( .B1(n150), .B2(n131), .A(n424), .ZN(n130) );
  INV_X1 U386 ( .A(n417), .ZN(n131) );
  INV_X1 U387 ( .A(n150), .ZN(n148) );
  INV_X1 U388 ( .A(n149), .ZN(n147) );
  INV_X1 U389 ( .A(n151), .ZN(n149) );
  INV_X1 U390 ( .A(n219), .ZN(n217) );
  OAI21_X1 U391 ( .B1(n246), .B2(n197), .A(n198), .ZN(n196) );
  NAND2_X1 U392 ( .A1(n217), .A2(n203), .ZN(n197) );
  AOI21_X1 U393 ( .B1(n218), .B2(n203), .A(n204), .ZN(n198) );
  OAI21_X1 U394 ( .B1(n246), .B2(n219), .A(n220), .ZN(n214) );
  OAI21_X1 U395 ( .B1(n246), .B2(n237), .A(n234), .ZN(n232) );
  INV_X1 U396 ( .A(n240), .ZN(n234) );
  INV_X1 U397 ( .A(n96), .ZN(n94) );
  INV_X1 U398 ( .A(n152), .ZN(n150) );
  INV_X1 U399 ( .A(n247), .ZN(n246) );
  AOI21_X1 U400 ( .B1(n247), .B2(n179), .A(n180), .ZN(n178) );
  NOR2_X1 U401 ( .A1(n219), .A2(n181), .ZN(n179) );
  AOI21_X1 U402 ( .B1(n267), .B2(n258), .A(n259), .ZN(n257) );
  NOR2_X1 U403 ( .A1(n421), .A2(n86), .ZN(n84) );
  INV_X1 U404 ( .A(n421), .ZN(n93) );
  NAND2_X1 U405 ( .A1(n122), .A2(n149), .ZN(n120) );
  AOI21_X1 U406 ( .B1(n122), .B2(n150), .A(n123), .ZN(n121) );
  NOR2_X1 U407 ( .A1(n417), .A2(n124), .ZN(n122) );
  INV_X1 U408 ( .A(n436), .ZN(n109) );
  INV_X1 U409 ( .A(n434), .ZN(n110) );
  INV_X1 U410 ( .A(n60), .ZN(n58) );
  INV_X1 U411 ( .A(n220), .ZN(n218) );
  INV_X1 U412 ( .A(n424), .ZN(n134) );
  INV_X1 U413 ( .A(n170), .ZN(n168) );
  OAI21_X1 U414 ( .B1(n246), .B2(n188), .A(n189), .ZN(n187) );
  NAND2_X1 U415 ( .A1(n190), .A2(n217), .ZN(n188) );
  AOI21_X1 U416 ( .B1(n190), .B2(n218), .A(n191), .ZN(n189) );
  NOR2_X1 U417 ( .A1(n201), .A2(n194), .ZN(n190) );
  NAND2_X1 U418 ( .A1(n239), .A2(n221), .ZN(n219) );
  INV_X1 U419 ( .A(n204), .ZN(n202) );
  INV_X1 U420 ( .A(n268), .ZN(n267) );
  INV_X1 U421 ( .A(n203), .ZN(n201) );
  INV_X1 U422 ( .A(n277), .ZN(n276) );
  INV_X1 U423 ( .A(n169), .ZN(n167) );
  INV_X1 U424 ( .A(n171), .ZN(n169) );
  INV_X1 U425 ( .A(n239), .ZN(n237) );
  INV_X1 U426 ( .A(n59), .ZN(n57) );
  OAI21_X1 U427 ( .B1(n241), .B2(n245), .A(n242), .ZN(n240) );
  NOR2_X1 U428 ( .A1(n230), .A2(n223), .ZN(n221) );
  NOR2_X1 U429 ( .A1(n244), .A2(n241), .ZN(n239) );
  NAND2_X1 U430 ( .A1(n167), .A2(n160), .ZN(n158) );
  AOI21_X1 U431 ( .B1(n168), .B2(n160), .A(n161), .ZN(n159) );
  INV_X1 U432 ( .A(n162), .ZN(n160) );
  AOI21_X1 U433 ( .B1(n269), .B2(n277), .A(n270), .ZN(n268) );
  OAI21_X1 U434 ( .B1(n271), .B2(n275), .A(n272), .ZN(n270) );
  NOR2_X1 U435 ( .A1(n274), .A2(n271), .ZN(n269) );
  NOR2_X1 U436 ( .A1(n212), .A2(n205), .ZN(n203) );
  AOI21_X1 U437 ( .B1(n153), .B2(n172), .A(n154), .ZN(n152) );
  OAI21_X1 U438 ( .B1(n260), .B2(n266), .A(n261), .ZN(n259) );
  OAI21_X1 U439 ( .B1(n278), .B2(n281), .A(n279), .ZN(n277) );
  BUF_X1 U440 ( .A(n112), .Z(n3) );
  NOR2_X1 U441 ( .A1(n265), .A2(n260), .ZN(n258) );
  NOR2_X1 U442 ( .A1(n255), .A2(n252), .ZN(n250) );
  AOI21_X1 U443 ( .B1(n221), .B2(n240), .A(n222), .ZN(n220) );
  INV_X1 U444 ( .A(n106), .ZN(n104) );
  AOI21_X1 U445 ( .B1(n150), .B2(n142), .A(n143), .ZN(n141) );
  NAND2_X1 U446 ( .A1(n149), .A2(n142), .ZN(n140) );
  OAI21_X1 U447 ( .B1(n268), .B2(n248), .A(n249), .ZN(n247) );
  AOI21_X1 U448 ( .B1(n250), .B2(n259), .A(n251), .ZN(n249) );
  NAND2_X1 U449 ( .A1(n258), .A2(n250), .ZN(n248) );
  OAI21_X1 U450 ( .B1(n252), .B2(n256), .A(n253), .ZN(n251) );
  NOR2_X1 U451 ( .A1(n162), .A2(n425), .ZN(n153) );
  INV_X1 U452 ( .A(n51), .ZN(n49) );
  AOI21_X1 U453 ( .B1(n267), .B2(n309), .A(n264), .ZN(n262) );
  INV_X1 U454 ( .A(n266), .ZN(n264) );
  OAI21_X1 U455 ( .B1(n134), .B2(n124), .A(n420), .ZN(n123) );
  OAI21_X1 U456 ( .B1(n202), .B2(n194), .A(n195), .ZN(n191) );
  INV_X1 U457 ( .A(n125), .ZN(n124) );
  OAI21_X1 U458 ( .B1(n246), .B2(n244), .A(n245), .ZN(n243) );
  OAI21_X1 U459 ( .B1(n276), .B2(n274), .A(n275), .ZN(n273) );
  OAI21_X1 U460 ( .B1(n246), .B2(n208), .A(n209), .ZN(n207) );
  AOI21_X1 U461 ( .B1(n218), .B2(n210), .A(n211), .ZN(n209) );
  NAND2_X1 U462 ( .A1(n217), .A2(n210), .ZN(n208) );
  INV_X1 U463 ( .A(n213), .ZN(n211) );
  OAI21_X1 U464 ( .B1(n246), .B2(n226), .A(n227), .ZN(n225) );
  NAND2_X1 U465 ( .A1(n239), .A2(n228), .ZN(n226) );
  AOI21_X1 U466 ( .B1(n240), .B2(n228), .A(n229), .ZN(n227) );
  INV_X1 U467 ( .A(n230), .ZN(n228) );
  INV_X1 U468 ( .A(n212), .ZN(n210) );
  INV_X1 U469 ( .A(n194), .ZN(n193) );
  NAND2_X1 U470 ( .A1(n296), .A2(n174), .ZN(n21) );
  INV_X1 U471 ( .A(n173), .ZN(n296) );
  INV_X1 U472 ( .A(n255), .ZN(n307) );
  INV_X1 U473 ( .A(n274), .ZN(n311) );
  INV_X1 U474 ( .A(n265), .ZN(n309) );
  NAND2_X1 U475 ( .A1(n294), .A2(n156), .ZN(n19) );
  NAND2_X1 U476 ( .A1(n298), .A2(n186), .ZN(n23) );
  INV_X1 U477 ( .A(n185), .ZN(n298) );
  INV_X1 U478 ( .A(n260), .ZN(n308) );
  INV_X1 U479 ( .A(n271), .ZN(n310) );
  NAND2_X1 U480 ( .A1(n160), .A2(n163), .ZN(n20) );
  NAND2_X1 U481 ( .A1(n306), .A2(n253), .ZN(n31) );
  INV_X1 U482 ( .A(n252), .ZN(n306) );
  INV_X1 U483 ( .A(n244), .ZN(n305) );
  NAND2_X1 U484 ( .A1(n297), .A2(n177), .ZN(n22) );
  NAND2_X1 U485 ( .A1(n210), .A2(n213), .ZN(n26) );
  NAND2_X1 U486 ( .A1(n228), .A2(n231), .ZN(n28) );
  NAND2_X1 U487 ( .A1(n193), .A2(n195), .ZN(n24) );
  XOR2_X1 U488 ( .A(n37), .B(n281), .Z(SUM[1]) );
  NAND2_X1 U489 ( .A1(n312), .A2(n279), .ZN(n37) );
  XOR2_X1 U490 ( .A(n276), .B(n36), .Z(SUM[2]) );
  NAND2_X1 U491 ( .A1(n311), .A2(n275), .ZN(n36) );
  XNOR2_X1 U492 ( .A(n273), .B(n35), .ZN(SUM[3]) );
  NAND2_X1 U493 ( .A1(n310), .A2(n272), .ZN(n35) );
  XNOR2_X1 U494 ( .A(n267), .B(n34), .ZN(SUM[4]) );
  NAND2_X1 U495 ( .A1(n309), .A2(n266), .ZN(n34) );
  XOR2_X1 U496 ( .A(n262), .B(n33), .Z(SUM[5]) );
  NAND2_X1 U497 ( .A1(n308), .A2(n261), .ZN(n33) );
  XOR2_X1 U498 ( .A(n246), .B(n30), .Z(SUM[8]) );
  NAND2_X1 U499 ( .A1(n305), .A2(n245), .ZN(n30) );
  XOR2_X1 U500 ( .A(n257), .B(n32), .Z(SUM[6]) );
  NAND2_X1 U501 ( .A1(n307), .A2(n256), .ZN(n32) );
  XNOR2_X1 U502 ( .A(n254), .B(n31), .ZN(SUM[7]) );
  OAI21_X1 U503 ( .B1(n257), .B2(n255), .A(n256), .ZN(n254) );
  NAND2_X1 U504 ( .A1(n304), .A2(n242), .ZN(n29) );
  NAND2_X1 U505 ( .A1(n300), .A2(n206), .ZN(n25) );
  INV_X1 U506 ( .A(n205), .ZN(n300) );
  NAND2_X1 U507 ( .A1(n292), .A2(n138), .ZN(n17) );
  INV_X1 U508 ( .A(n278), .ZN(n312) );
  NAND2_X1 U509 ( .A1(n302), .A2(n224), .ZN(n27) );
  INV_X1 U510 ( .A(n163), .ZN(n161) );
  INV_X1 U511 ( .A(n87), .ZN(n86) );
  INV_X1 U512 ( .A(n88), .ZN(n87) );
  INV_X1 U513 ( .A(n107), .ZN(n105) );
  INV_X1 U514 ( .A(n423), .ZN(n284) );
  INV_X1 U515 ( .A(n231), .ZN(n229) );
  INV_X1 U516 ( .A(n69), .ZN(n68) );
  INV_X1 U517 ( .A(n70), .ZN(n69) );
  AND2_X1 U518 ( .A1(n438), .A2(n281), .ZN(SUM[0]) );
  NOR2_X1 U519 ( .A1(A[18]), .A2(B[18]), .ZN(n162) );
  OR2_X1 U520 ( .A1(A[0]), .A2(B[0]), .ZN(n438) );
  NOR2_X1 U521 ( .A1(A[13]), .A2(B[13]), .ZN(n205) );
  NOR2_X1 U522 ( .A1(B[26]), .A2(A[26]), .ZN(n88) );
  NOR2_X1 U523 ( .A1(A[24]), .A2(B[24]), .ZN(n106) );
  NOR2_X1 U524 ( .A1(B[29]), .A2(A[29]), .ZN(n61) );
  NOR2_X1 U525 ( .A1(A[15]), .A2(B[15]), .ZN(n185) );
  NOR2_X1 U526 ( .A1(A[9]), .A2(B[9]), .ZN(n241) );
  NOR2_X1 U527 ( .A1(B[19]), .A2(A[19]), .ZN(n155) );
  NOR2_X1 U528 ( .A1(A[11]), .A2(B[11]), .ZN(n223) );
  NOR2_X1 U529 ( .A1(A[17]), .A2(B[17]), .ZN(n173) );
  NAND2_X1 U530 ( .A1(A[18]), .A2(B[18]), .ZN(n163) );
  NOR2_X1 U531 ( .A1(A[14]), .A2(B[14]), .ZN(n194) );
  NAND2_X1 U532 ( .A1(A[4]), .A2(B[4]), .ZN(n266) );
  NAND2_X1 U533 ( .A1(A[6]), .A2(B[6]), .ZN(n256) );
  NAND2_X1 U534 ( .A1(A[8]), .A2(B[8]), .ZN(n245) );
  NAND2_X1 U535 ( .A1(A[2]), .A2(B[2]), .ZN(n275) );
  NAND2_X1 U536 ( .A1(A[7]), .A2(B[7]), .ZN(n253) );
  NAND2_X1 U537 ( .A1(A[0]), .A2(B[0]), .ZN(n281) );
  XNOR2_X1 U538 ( .A(n243), .B(n29), .ZN(SUM[9]) );
  NAND2_X1 U539 ( .A1(A[14]), .A2(B[14]), .ZN(n195) );
  NAND2_X1 U540 ( .A1(A[12]), .A2(B[12]), .ZN(n213) );
  NAND2_X1 U541 ( .A1(A[10]), .A2(B[10]), .ZN(n231) );
  NAND2_X1 U542 ( .A1(A[5]), .A2(B[5]), .ZN(n261) );
  NAND2_X1 U543 ( .A1(A[1]), .A2(B[1]), .ZN(n279) );
  NAND2_X1 U544 ( .A1(A[3]), .A2(B[3]), .ZN(n272) );
  NAND2_X1 U545 ( .A1(A[9]), .A2(B[9]), .ZN(n242) );
  NAND2_X1 U546 ( .A1(A[13]), .A2(B[13]), .ZN(n206) );
  NAND2_X1 U547 ( .A1(A[31]), .A2(B[31]), .ZN(n40) );
  NAND2_X1 U548 ( .A1(A[11]), .A2(B[11]), .ZN(n224) );
  NAND2_X1 U549 ( .A1(n284), .A2(n62), .ZN(n9) );
  NAND2_X1 U550 ( .A1(n416), .A2(n51), .ZN(n8) );
  NAND2_X1 U551 ( .A1(n286), .A2(n80), .ZN(n11) );
  NAND2_X1 U552 ( .A1(n288), .A2(n100), .ZN(n13) );
  NAND2_X1 U553 ( .A1(n87), .A2(n89), .ZN(n12) );
  NAND2_X1 U554 ( .A1(n69), .A2(n71), .ZN(n10) );
  NAND2_X1 U555 ( .A1(n439), .A2(n40), .ZN(n7) );
  NAND2_X1 U556 ( .A1(n104), .A2(n107), .ZN(n14) );
  XNOR2_X1 U557 ( .A(n232), .B(n28), .ZN(SUM[10]) );
  XNOR2_X1 U558 ( .A(n225), .B(n27), .ZN(SUM[11]) );
  XNOR2_X1 U559 ( .A(n128), .B(n16), .ZN(SUM[22]) );
  NAND2_X1 U560 ( .A1(n125), .A2(n420), .ZN(n16) );
  NAND2_X1 U561 ( .A1(n290), .A2(n432), .ZN(n15) );
  XNOR2_X1 U562 ( .A(n175), .B(n21), .ZN(SUM[17]) );
  XNOR2_X1 U563 ( .A(n157), .B(n19), .ZN(SUM[19]) );
  XNOR2_X1 U564 ( .A(n146), .B(n18), .ZN(SUM[20]) );
  XNOR2_X1 U565 ( .A(n164), .B(n20), .ZN(SUM[18]) );
  XNOR2_X1 U566 ( .A(n196), .B(n24), .ZN(SUM[14]) );
  XNOR2_X1 U567 ( .A(n187), .B(n23), .ZN(SUM[15]) );
  XNOR2_X1 U568 ( .A(n207), .B(n25), .ZN(SUM[13]) );
  XNOR2_X1 U569 ( .A(n214), .B(n26), .ZN(SUM[12]) );
  OR2_X1 U570 ( .A1(A[31]), .A2(B[31]), .ZN(n439) );
  NAND2_X1 U571 ( .A1(A[30]), .A2(B[30]), .ZN(n51) );
  INV_X1 U572 ( .A(n176), .ZN(n297) );
  NOR2_X1 U573 ( .A1(A[16]), .A2(B[16]), .ZN(n176) );
  NAND2_X1 U574 ( .A1(A[15]), .A2(B[15]), .ZN(n186) );
  INV_X1 U575 ( .A(n435), .ZN(n290) );
  INV_X1 U576 ( .A(n223), .ZN(n302) );
  OAI21_X1 U577 ( .B1(n223), .B2(n231), .A(n224), .ZN(n222) );
  NAND2_X1 U578 ( .A1(A[28]), .A2(B[28]), .ZN(n71) );
  NOR2_X1 U579 ( .A1(A[28]), .A2(B[28]), .ZN(n70) );
  NAND2_X1 U580 ( .A1(B[29]), .A2(A[29]), .ZN(n62) );
  INV_X1 U581 ( .A(n426), .ZN(n142) );
  NOR2_X1 U582 ( .A1(A[20]), .A2(B[20]), .ZN(n144) );
  INV_X1 U583 ( .A(n422), .ZN(n286) );
  NOR2_X1 U584 ( .A1(n88), .A2(n428), .ZN(n77) );
  NAND2_X1 U585 ( .A1(B[26]), .A2(A[26]), .ZN(n89) );
  INV_X1 U586 ( .A(n172), .ZN(n170) );
  OAI21_X1 U587 ( .B1(n173), .B2(n177), .A(n174), .ZN(n172) );
  NAND2_X1 U588 ( .A1(n142), .A2(n145), .ZN(n18) );
  INV_X1 U589 ( .A(n145), .ZN(n143) );
  NAND2_X1 U590 ( .A1(B[21]), .A2(A[21]), .ZN(n138) );
  NOR2_X1 U591 ( .A1(B[21]), .A2(A[21]), .ZN(n137) );
  INV_X1 U592 ( .A(n429), .ZN(n288) );
  NOR2_X1 U593 ( .A1(n106), .A2(n99), .ZN(n97) );
  NAND2_X1 U594 ( .A1(B[25]), .A2(A[25]), .ZN(n100) );
  INV_X1 U595 ( .A(n126), .ZN(n125) );
  XNOR2_X1 U596 ( .A(n41), .B(n7), .ZN(SUM[31]) );
  INV_X1 U597 ( .A(n418), .ZN(n292) );
  OAI21_X1 U598 ( .B1(n96), .B2(n86), .A(n89), .ZN(n85) );
  INV_X1 U599 ( .A(n98), .ZN(n96) );
  NAND2_X1 U600 ( .A1(B[23]), .A2(A[23]), .ZN(n118) );
  NOR2_X1 U601 ( .A1(B[23]), .A2(A[23]), .ZN(n117) );
  NOR2_X1 U602 ( .A1(n176), .A2(n173), .ZN(n171) );
  INV_X1 U603 ( .A(n241), .ZN(n304) );
  INV_X1 U604 ( .A(n6), .ZN(n75) );
  AOI21_X1 U605 ( .B1(n98), .B2(n77), .A(n78), .ZN(n440) );
  AOI21_X1 U606 ( .B1(n98), .B2(n77), .A(n78), .ZN(n5) );
  XNOR2_X1 U607 ( .A(n72), .B(n10), .ZN(SUM[28]) );
  NAND2_X1 U608 ( .A1(A[17]), .A2(B[17]), .ZN(n174) );
  AOI21_X1 U609 ( .B1(n60), .B2(n416), .A(n49), .ZN(n47) );
  NAND2_X1 U610 ( .A1(n97), .A2(n77), .ZN(n6) );
  XNOR2_X1 U611 ( .A(n101), .B(n13), .ZN(SUM[25]) );
  NAND2_X1 U612 ( .A1(B[22]), .A2(A[22]), .ZN(n127) );
  NOR2_X1 U613 ( .A1(B[22]), .A2(A[22]), .ZN(n126) );
  XNOR2_X1 U614 ( .A(n90), .B(n12), .ZN(SUM[26]) );
  NAND2_X1 U615 ( .A1(A[24]), .A2(B[24]), .ZN(n107) );
  XNOR2_X1 U616 ( .A(n139), .B(n17), .ZN(SUM[21]) );
  OAI21_X1 U617 ( .B1(n155), .B2(n163), .A(n156), .ZN(n154) );
  INV_X1 U618 ( .A(n419), .ZN(n294) );
  OAI21_X1 U619 ( .B1(n429), .B2(n107), .A(n100), .ZN(n98) );
  NAND2_X1 U620 ( .A1(n171), .A2(n153), .ZN(n151) );
  NAND2_X1 U621 ( .A1(A[16]), .A2(B[16]), .ZN(n177) );
  XNOR2_X1 U622 ( .A(n52), .B(n8), .ZN(SUM[30]) );
  XNOR2_X1 U623 ( .A(n108), .B(n14), .ZN(SUM[24]) );
  XNOR2_X1 U624 ( .A(n81), .B(n11), .ZN(SUM[27]) );
  XNOR2_X1 U625 ( .A(n119), .B(n15), .ZN(SUM[23]) );
  OAI21_X1 U626 ( .B1(n2), .B2(n64), .A(n65), .ZN(n63) );
  OAI21_X1 U627 ( .B1(n2), .B2(n109), .A(n110), .ZN(n108) );
  OAI21_X1 U628 ( .B1(n102), .B2(n2), .A(n103), .ZN(n101) );
  OAI21_X1 U629 ( .B1(n73), .B2(n2), .A(n74), .ZN(n72) );
  OAI21_X1 U630 ( .B1(n1), .B2(n91), .A(n92), .ZN(n90) );
  OAI21_X1 U631 ( .B1(n220), .B2(n181), .A(n182), .ZN(n180) );
  OAI21_X1 U632 ( .B1(n205), .B2(n213), .A(n206), .ZN(n204) );
  OAI21_X1 U633 ( .B1(n2), .B2(n82), .A(n83), .ZN(n81) );
  XOR2_X1 U634 ( .A(n2), .B(n22), .Z(SUM[16]) );
  OAI21_X1 U635 ( .B1(n1), .B2(n120), .A(n121), .ZN(n119) );
  OAI21_X1 U636 ( .B1(n1), .B2(n129), .A(n130), .ZN(n128) );
  OAI21_X1 U637 ( .B1(n1), .B2(n140), .A(n141), .ZN(n139) );
  OAI21_X1 U638 ( .B1(n1), .B2(n169), .A(n170), .ZN(n164) );
  OAI21_X1 U639 ( .B1(n1), .B2(n158), .A(n159), .ZN(n157) );
  OAI21_X1 U640 ( .B1(n1), .B2(n147), .A(n148), .ZN(n146) );
  OAI21_X1 U641 ( .B1(n1), .B2(n176), .A(n177), .ZN(n175) );
  AOI21_X1 U642 ( .B1(n183), .B2(n204), .A(n184), .ZN(n182) );
  NAND2_X1 U643 ( .A1(n203), .A2(n183), .ZN(n181) );
  OAI21_X1 U644 ( .B1(n42), .B2(n2), .A(n43), .ZN(n41) );
  NOR2_X1 U645 ( .A1(n6), .A2(n57), .ZN(n55) );
  NOR2_X1 U646 ( .A1(n6), .A2(n68), .ZN(n66) );
  NOR2_X1 U647 ( .A1(n6), .A2(n46), .ZN(n44) );
  OAI21_X1 U648 ( .B1(n2), .B2(n53), .A(n54), .ZN(n52) );
  INV_X1 U649 ( .A(n5), .ZN(n76) );
  NAND2_X1 U650 ( .A1(n4), .A2(n66), .ZN(n64) );
  NAND2_X1 U651 ( .A1(n4), .A2(n84), .ZN(n82) );
  NAND2_X1 U652 ( .A1(n4), .A2(n93), .ZN(n91) );
  NAND2_X1 U653 ( .A1(n436), .A2(n75), .ZN(n73) );
  NAND2_X1 U654 ( .A1(n436), .A2(n44), .ZN(n42) );
  NAND2_X1 U655 ( .A1(n4), .A2(n55), .ZN(n53) );
  NAND2_X1 U656 ( .A1(n436), .A2(n104), .ZN(n102) );
  NAND2_X1 U657 ( .A1(A[19]), .A2(B[19]), .ZN(n156) );
  NAND2_X1 U658 ( .A1(n59), .A2(n416), .ZN(n46) );
  NOR2_X1 U659 ( .A1(n70), .A2(n61), .ZN(n59) );
  OAI21_X1 U660 ( .B1(n152), .B2(n113), .A(n114), .ZN(n112) );
  NOR2_X1 U661 ( .A1(n113), .A2(n151), .ZN(n111) );
  OAI21_X1 U662 ( .B1(n61), .B2(n71), .A(n62), .ZN(n60) );
  NAND2_X1 U663 ( .A1(n430), .A2(n135), .ZN(n113) );
  NOR2_X1 U664 ( .A1(n144), .A2(n427), .ZN(n135) );
  XNOR2_X1 U665 ( .A(n63), .B(n9), .ZN(SUM[29]) );
  NOR2_X1 U666 ( .A1(n194), .A2(n185), .ZN(n183) );
  OAI21_X1 U667 ( .B1(n185), .B2(n195), .A(n186), .ZN(n184) );
  AOI21_X1 U668 ( .B1(n433), .B2(n93), .A(n94), .ZN(n92) );
  AOI21_X1 U669 ( .B1(n3), .B2(n104), .A(n105), .ZN(n103) );
  AOI21_X1 U670 ( .B1(n434), .B2(n75), .A(n76), .ZN(n74) );
  AOI21_X1 U671 ( .B1(n433), .B2(n84), .A(n85), .ZN(n83) );
  AOI21_X1 U672 ( .B1(n3), .B2(n44), .A(n45), .ZN(n43) );
  AOI21_X1 U673 ( .B1(n3), .B2(n55), .A(n56), .ZN(n54) );
  AOI21_X1 U674 ( .B1(n434), .B2(n66), .A(n67), .ZN(n65) );
  AOI21_X1 U675 ( .B1(n430), .B2(n136), .A(n116), .ZN(n114) );
  NAND2_X1 U676 ( .A1(B[20]), .A2(A[20]), .ZN(n145) );
  OAI21_X1 U677 ( .B1(n440), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U678 ( .B1(n440), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U679 ( .B1(n5), .B2(n68), .A(n71), .ZN(n67) );
  OAI21_X1 U680 ( .B1(n79), .B2(n89), .A(n80), .ZN(n78) );
  NAND2_X1 U681 ( .A1(A[27]), .A2(B[27]), .ZN(n80) );
  NOR2_X1 U682 ( .A1(B[27]), .A2(A[27]), .ZN(n79) );
  OAI21_X1 U683 ( .B1(n117), .B2(n127), .A(n118), .ZN(n116) );
  OAI21_X1 U684 ( .B1(n137), .B2(n145), .A(n138), .ZN(n136) );
endmodule


module datapath_DW01_add_12 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n39, n41, n42, n43, n44, n45, n46,
         n47, n49, n51, n52, n53, n54, n55, n56, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n193, n194, n195, n196, n197, n198, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n234, n237, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n281, n284, n286, n288, n290,
         n292, n294, n296, n297, n298, n300, n302, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n416, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440;

  NOR2_X2 U349 ( .A1(A[14]), .A2(B[14]), .ZN(n194) );
  OR2_X1 U350 ( .A1(A[30]), .A2(B[30]), .ZN(n416) );
  AND2_X1 U351 ( .A1(n418), .A2(n281), .ZN(SUM[0]) );
  OR2_X1 U352 ( .A1(A[0]), .A2(B[0]), .ZN(n418) );
  NAND2_X1 U353 ( .A1(n97), .A2(n77), .ZN(n419) );
  INV_X1 U354 ( .A(n143), .ZN(n420) );
  CLKBUF_X1 U355 ( .A(n127), .Z(n421) );
  NOR2_X1 U356 ( .A1(B[25]), .A2(A[25]), .ZN(n422) );
  NOR2_X1 U357 ( .A1(B[25]), .A2(A[25]), .ZN(n99) );
  NOR2_X2 U358 ( .A1(n79), .A2(n88), .ZN(n77) );
  CLKBUF_X1 U359 ( .A(n118), .Z(n423) );
  CLKBUF_X1 U360 ( .A(n88), .Z(n424) );
  OR2_X1 U361 ( .A1(n70), .A2(n61), .ZN(n425) );
  NOR2_X1 U362 ( .A1(A[29]), .A2(B[29]), .ZN(n426) );
  NOR2_X1 U363 ( .A1(B[27]), .A2(A[27]), .ZN(n427) );
  NOR2_X1 U364 ( .A1(A[19]), .A2(B[19]), .ZN(n428) );
  OR2_X1 U365 ( .A1(n144), .A2(n137), .ZN(n429) );
  CLKBUF_X1 U366 ( .A(n136), .Z(n430) );
  NOR2_X1 U367 ( .A1(A[21]), .A2(B[21]), .ZN(n431) );
  CLKBUF_X1 U368 ( .A(n144), .Z(n432) );
  CLKBUF_X1 U369 ( .A(n427), .Z(n433) );
  NOR2_X1 U370 ( .A1(B[23]), .A2(A[23]), .ZN(n434) );
  CLKBUF_X1 U371 ( .A(n137), .Z(n435) );
  CLKBUF_X1 U372 ( .A(n117), .Z(n436) );
  BUF_X1 U373 ( .A(n112), .Z(n437) );
  BUF_X1 U374 ( .A(n111), .Z(n438) );
  NOR2_X1 U375 ( .A1(A[10]), .A2(B[10]), .ZN(n230) );
  NOR2_X1 U376 ( .A1(A[4]), .A2(B[4]), .ZN(n265) );
  NOR2_X1 U377 ( .A1(A[12]), .A2(B[12]), .ZN(n212) );
  NOR2_X1 U378 ( .A1(A[3]), .A2(B[3]), .ZN(n271) );
  NOR2_X1 U379 ( .A1(A[5]), .A2(B[5]), .ZN(n260) );
  NOR2_X1 U380 ( .A1(A[9]), .A2(B[9]), .ZN(n241) );
  NOR2_X1 U381 ( .A1(A[7]), .A2(B[7]), .ZN(n252) );
  NOR2_X1 U382 ( .A1(A[8]), .A2(B[8]), .ZN(n244) );
  NOR2_X1 U383 ( .A1(A[6]), .A2(B[6]), .ZN(n255) );
  NOR2_X1 U384 ( .A1(A[2]), .A2(B[2]), .ZN(n274) );
  NOR2_X1 U385 ( .A1(A[1]), .A2(B[1]), .ZN(n278) );
  INV_X1 U386 ( .A(n150), .ZN(n148) );
  INV_X1 U387 ( .A(n151), .ZN(n149) );
  BUF_X1 U388 ( .A(n178), .Z(n1) );
  INV_X1 U389 ( .A(n219), .ZN(n217) );
  OAI21_X1 U390 ( .B1(n246), .B2(n197), .A(n198), .ZN(n196) );
  AOI21_X1 U391 ( .B1(n218), .B2(n203), .A(n200), .ZN(n198) );
  NAND2_X1 U392 ( .A1(n217), .A2(n203), .ZN(n197) );
  INV_X1 U393 ( .A(n202), .ZN(n200) );
  OAI21_X1 U394 ( .B1(n246), .B2(n219), .A(n220), .ZN(n214) );
  OAI21_X1 U395 ( .B1(n246), .B2(n237), .A(n234), .ZN(n232) );
  INV_X1 U396 ( .A(n240), .ZN(n234) );
  BUF_X1 U397 ( .A(n178), .Z(n2) );
  BUF_X1 U398 ( .A(n111), .Z(n4) );
  NAND2_X1 U399 ( .A1(n149), .A2(n131), .ZN(n129) );
  AOI21_X1 U400 ( .B1(n150), .B2(n131), .A(n430), .ZN(n130) );
  INV_X1 U401 ( .A(n429), .ZN(n131) );
  INV_X1 U402 ( .A(n152), .ZN(n150) );
  INV_X1 U403 ( .A(n247), .ZN(n246) );
  NAND2_X1 U404 ( .A1(n122), .A2(n149), .ZN(n120) );
  AOI21_X1 U405 ( .B1(n122), .B2(n150), .A(n123), .ZN(n121) );
  NOR2_X1 U406 ( .A1(n429), .A2(n124), .ZN(n122) );
  AOI21_X1 U407 ( .B1(n267), .B2(n258), .A(n259), .ZN(n257) );
  AOI21_X1 U408 ( .B1(n247), .B2(n179), .A(n180), .ZN(n178) );
  NOR2_X1 U409 ( .A1(n201), .A2(n194), .ZN(n190) );
  INV_X1 U410 ( .A(n60), .ZN(n58) );
  INV_X1 U411 ( .A(n220), .ZN(n218) );
  INV_X1 U412 ( .A(n430), .ZN(n134) );
  INV_X1 U413 ( .A(n204), .ZN(n202) );
  NAND2_X1 U414 ( .A1(n203), .A2(n183), .ZN(n181) );
  OAI21_X1 U415 ( .B1(n2), .B2(n109), .A(n110), .ZN(n108) );
  INV_X1 U416 ( .A(n3), .ZN(n110) );
  INV_X1 U417 ( .A(n438), .ZN(n109) );
  NAND2_X1 U418 ( .A1(n239), .A2(n221), .ZN(n219) );
  INV_X1 U419 ( .A(n203), .ZN(n201) );
  INV_X1 U420 ( .A(n268), .ZN(n267) );
  INV_X1 U421 ( .A(n170), .ZN(n168) );
  INV_X1 U422 ( .A(n172), .ZN(n170) );
  INV_X1 U423 ( .A(n277), .ZN(n276) );
  INV_X1 U424 ( .A(n169), .ZN(n167) );
  INV_X1 U425 ( .A(n171), .ZN(n169) );
  INV_X1 U426 ( .A(n239), .ZN(n237) );
  OAI21_X1 U427 ( .B1(n426), .B2(n71), .A(n62), .ZN(n60) );
  AOI21_X1 U428 ( .B1(n150), .B2(n142), .A(n143), .ZN(n141) );
  NAND2_X1 U429 ( .A1(n149), .A2(n142), .ZN(n140) );
  INV_X1 U430 ( .A(n145), .ZN(n143) );
  NAND2_X1 U431 ( .A1(n167), .A2(n160), .ZN(n158) );
  AOI21_X1 U432 ( .B1(n168), .B2(n160), .A(n161), .ZN(n159) );
  INV_X1 U433 ( .A(n162), .ZN(n160) );
  AOI21_X1 U434 ( .B1(n269), .B2(n277), .A(n270), .ZN(n268) );
  OAI21_X1 U435 ( .B1(n271), .B2(n275), .A(n272), .ZN(n270) );
  NOR2_X1 U436 ( .A1(n274), .A2(n271), .ZN(n269) );
  OAI21_X1 U437 ( .B1(n241), .B2(n245), .A(n242), .ZN(n240) );
  AOI21_X1 U438 ( .B1(n153), .B2(n172), .A(n154), .ZN(n152) );
  OAI21_X1 U439 ( .B1(n260), .B2(n266), .A(n261), .ZN(n259) );
  OAI21_X1 U440 ( .B1(n278), .B2(n281), .A(n279), .ZN(n277) );
  BUF_X1 U441 ( .A(n112), .Z(n3) );
  NOR2_X1 U442 ( .A1(n255), .A2(n252), .ZN(n250) );
  AOI21_X1 U443 ( .B1(n221), .B2(n240), .A(n222), .ZN(n220) );
  NOR2_X1 U444 ( .A1(n244), .A2(n241), .ZN(n239) );
  NOR2_X1 U445 ( .A1(n265), .A2(n260), .ZN(n258) );
  INV_X1 U446 ( .A(n106), .ZN(n104) );
  OAI21_X1 U447 ( .B1(n268), .B2(n248), .A(n249), .ZN(n247) );
  AOI21_X1 U448 ( .B1(n250), .B2(n259), .A(n251), .ZN(n249) );
  NAND2_X1 U449 ( .A1(n258), .A2(n250), .ZN(n248) );
  OAI21_X1 U450 ( .B1(n252), .B2(n256), .A(n253), .ZN(n251) );
  NOR2_X1 U451 ( .A1(n162), .A2(n428), .ZN(n153) );
  AOI21_X1 U452 ( .B1(n267), .B2(n309), .A(n264), .ZN(n262) );
  INV_X1 U453 ( .A(n266), .ZN(n264) );
  INV_X1 U454 ( .A(n432), .ZN(n142) );
  OAI21_X1 U455 ( .B1(n134), .B2(n124), .A(n421), .ZN(n123) );
  OAI21_X1 U456 ( .B1(n246), .B2(n244), .A(n245), .ZN(n243) );
  OAI21_X1 U457 ( .B1(n257), .B2(n255), .A(n256), .ZN(n254) );
  OAI21_X1 U458 ( .B1(n276), .B2(n274), .A(n275), .ZN(n273) );
  OAI21_X1 U459 ( .B1(n246), .B2(n188), .A(n189), .ZN(n187) );
  AOI21_X1 U460 ( .B1(n190), .B2(n218), .A(n191), .ZN(n189) );
  NAND2_X1 U461 ( .A1(n190), .A2(n217), .ZN(n188) );
  OAI21_X1 U462 ( .B1(n202), .B2(n194), .A(n195), .ZN(n191) );
  OAI21_X1 U463 ( .B1(n246), .B2(n208), .A(n209), .ZN(n207) );
  AOI21_X1 U464 ( .B1(n218), .B2(n210), .A(n211), .ZN(n209) );
  NAND2_X1 U465 ( .A1(n217), .A2(n210), .ZN(n208) );
  INV_X1 U466 ( .A(n213), .ZN(n211) );
  OAI21_X1 U467 ( .B1(n246), .B2(n226), .A(n227), .ZN(n225) );
  NAND2_X1 U468 ( .A1(n239), .A2(n228), .ZN(n226) );
  AOI21_X1 U469 ( .B1(n240), .B2(n228), .A(n229), .ZN(n227) );
  INV_X1 U470 ( .A(n230), .ZN(n228) );
  INV_X1 U471 ( .A(n212), .ZN(n210) );
  INV_X1 U472 ( .A(n194), .ZN(n193) );
  INV_X1 U473 ( .A(n125), .ZN(n124) );
  INV_X1 U474 ( .A(n126), .ZN(n125) );
  NAND2_X1 U475 ( .A1(n69), .A2(n71), .ZN(n10) );
  NAND2_X1 U476 ( .A1(n310), .A2(n272), .ZN(n35) );
  INV_X1 U477 ( .A(n271), .ZN(n310) );
  NAND2_X1 U478 ( .A1(n305), .A2(n245), .ZN(n30) );
  INV_X1 U479 ( .A(n244), .ZN(n305) );
  NAND2_X1 U480 ( .A1(n307), .A2(n256), .ZN(n32) );
  INV_X1 U481 ( .A(n255), .ZN(n307) );
  NAND2_X1 U482 ( .A1(n292), .A2(n138), .ZN(n17) );
  INV_X1 U483 ( .A(n435), .ZN(n292) );
  NAND2_X1 U484 ( .A1(n290), .A2(n423), .ZN(n15) );
  NAND2_X1 U485 ( .A1(n302), .A2(n224), .ZN(n27) );
  INV_X1 U486 ( .A(n223), .ZN(n302) );
  NAND2_X1 U487 ( .A1(n296), .A2(n174), .ZN(n21) );
  INV_X1 U488 ( .A(n173), .ZN(n296) );
  NAND2_X1 U489 ( .A1(n104), .A2(n107), .ZN(n14) );
  NAND2_X1 U490 ( .A1(n300), .A2(n206), .ZN(n25) );
  NAND2_X1 U491 ( .A1(n142), .A2(n420), .ZN(n18) );
  NAND2_X1 U492 ( .A1(n193), .A2(n195), .ZN(n24) );
  NAND2_X1 U493 ( .A1(n306), .A2(n253), .ZN(n31) );
  INV_X1 U494 ( .A(n252), .ZN(n306) );
  NAND2_X1 U495 ( .A1(n304), .A2(n242), .ZN(n29) );
  INV_X1 U496 ( .A(n241), .ZN(n304) );
  NAND2_X1 U497 ( .A1(n309), .A2(n266), .ZN(n34) );
  INV_X1 U498 ( .A(n265), .ZN(n309) );
  NAND2_X1 U499 ( .A1(n284), .A2(n62), .ZN(n9) );
  NAND2_X1 U500 ( .A1(n297), .A2(n177), .ZN(n22) );
  INV_X1 U501 ( .A(n176), .ZN(n297) );
  NAND2_X1 U502 ( .A1(n294), .A2(n156), .ZN(n19) );
  INV_X1 U503 ( .A(n428), .ZN(n294) );
  NAND2_X1 U504 ( .A1(n298), .A2(n186), .ZN(n23) );
  INV_X1 U505 ( .A(n185), .ZN(n298) );
  NAND2_X1 U506 ( .A1(n311), .A2(n275), .ZN(n36) );
  INV_X1 U507 ( .A(n274), .ZN(n311) );
  NAND2_X1 U508 ( .A1(n160), .A2(n163), .ZN(n20) );
  NAND2_X1 U509 ( .A1(n228), .A2(n231), .ZN(n28) );
  NAND2_X1 U510 ( .A1(n210), .A2(n213), .ZN(n26) );
  NAND2_X1 U511 ( .A1(n286), .A2(n80), .ZN(n11) );
  INV_X1 U512 ( .A(n433), .ZN(n286) );
  NAND2_X1 U513 ( .A1(n288), .A2(n100), .ZN(n13) );
  NAND2_X1 U514 ( .A1(n308), .A2(n261), .ZN(n33) );
  INV_X1 U515 ( .A(n260), .ZN(n308) );
  NAND2_X1 U516 ( .A1(n312), .A2(n279), .ZN(n37) );
  INV_X1 U517 ( .A(n278), .ZN(n312) );
  INV_X1 U518 ( .A(n231), .ZN(n229) );
  INV_X1 U519 ( .A(n163), .ZN(n161) );
  INV_X1 U520 ( .A(n69), .ZN(n68) );
  INV_X1 U521 ( .A(n107), .ZN(n105) );
  NOR2_X1 U522 ( .A1(A[20]), .A2(B[20]), .ZN(n144) );
  NOR2_X1 U523 ( .A1(B[22]), .A2(A[22]), .ZN(n126) );
  NOR2_X1 U524 ( .A1(A[11]), .A2(B[11]), .ZN(n223) );
  NOR2_X1 U525 ( .A1(B[27]), .A2(A[27]), .ZN(n79) );
  NOR2_X1 U526 ( .A1(B[26]), .A2(A[26]), .ZN(n88) );
  NOR2_X1 U527 ( .A1(A[17]), .A2(B[17]), .ZN(n173) );
  NOR2_X1 U528 ( .A1(A[18]), .A2(B[18]), .ZN(n162) );
  NOR2_X1 U529 ( .A1(A[19]), .A2(B[19]), .ZN(n155) );
  NAND2_X1 U530 ( .A1(A[24]), .A2(B[24]), .ZN(n107) );
  NAND2_X1 U531 ( .A1(B[20]), .A2(A[20]), .ZN(n145) );
  NAND2_X1 U532 ( .A1(B[22]), .A2(A[22]), .ZN(n127) );
  NAND2_X1 U533 ( .A1(A[14]), .A2(B[14]), .ZN(n195) );
  NOR2_X1 U534 ( .A1(A[13]), .A2(B[13]), .ZN(n205) );
  NOR2_X1 U535 ( .A1(A[24]), .A2(B[24]), .ZN(n106) );
  NOR2_X1 U536 ( .A1(A[15]), .A2(B[15]), .ZN(n185) );
  NAND2_X1 U537 ( .A1(A[6]), .A2(B[6]), .ZN(n256) );
  NAND2_X1 U538 ( .A1(A[8]), .A2(B[8]), .ZN(n245) );
  NAND2_X1 U539 ( .A1(A[4]), .A2(B[4]), .ZN(n266) );
  NAND2_X1 U540 ( .A1(A[2]), .A2(B[2]), .ZN(n275) );
  NAND2_X1 U541 ( .A1(A[9]), .A2(B[9]), .ZN(n242) );
  NAND2_X1 U542 ( .A1(A[7]), .A2(B[7]), .ZN(n253) );
  NAND2_X1 U543 ( .A1(A[0]), .A2(B[0]), .ZN(n281) );
  XNOR2_X1 U544 ( .A(n157), .B(n19), .ZN(SUM[19]) );
  XNOR2_X1 U545 ( .A(n108), .B(n14), .ZN(SUM[24]) );
  NAND2_X1 U546 ( .A1(A[19]), .A2(B[19]), .ZN(n156) );
  NAND2_X1 U547 ( .A1(A[15]), .A2(B[15]), .ZN(n186) );
  NAND2_X1 U548 ( .A1(A[18]), .A2(B[18]), .ZN(n163) );
  NAND2_X1 U549 ( .A1(A[12]), .A2(B[12]), .ZN(n213) );
  NAND2_X1 U550 ( .A1(A[10]), .A2(B[10]), .ZN(n231) );
  NAND2_X1 U551 ( .A1(A[5]), .A2(B[5]), .ZN(n261) );
  NAND2_X1 U552 ( .A1(A[1]), .A2(B[1]), .ZN(n279) );
  NAND2_X1 U553 ( .A1(A[3]), .A2(B[3]), .ZN(n272) );
  OR2_X1 U554 ( .A1(n39), .A2(n439), .ZN(n7) );
  AND2_X1 U555 ( .A1(A[31]), .A2(B[31]), .ZN(n439) );
  XNOR2_X1 U556 ( .A(n119), .B(n15), .ZN(SUM[23]) );
  XOR2_X1 U557 ( .A(n37), .B(n281), .Z(SUM[1]) );
  XOR2_X1 U558 ( .A(n276), .B(n36), .Z(SUM[2]) );
  XNOR2_X1 U559 ( .A(n273), .B(n35), .ZN(SUM[3]) );
  XNOR2_X1 U560 ( .A(n267), .B(n34), .ZN(SUM[4]) );
  XOR2_X1 U561 ( .A(n262), .B(n33), .Z(SUM[5]) );
  XNOR2_X1 U562 ( .A(n128), .B(n16), .ZN(SUM[22]) );
  NAND2_X1 U563 ( .A1(n125), .A2(n421), .ZN(n16) );
  XNOR2_X1 U564 ( .A(n90), .B(n12), .ZN(SUM[26]) );
  NAND2_X1 U565 ( .A1(n87), .A2(n89), .ZN(n12) );
  XNOR2_X1 U566 ( .A(n139), .B(n17), .ZN(SUM[21]) );
  XNOR2_X1 U567 ( .A(n146), .B(n18), .ZN(SUM[20]) );
  XNOR2_X1 U568 ( .A(n175), .B(n21), .ZN(SUM[17]) );
  XNOR2_X1 U569 ( .A(n164), .B(n20), .ZN(SUM[18]) );
  XNOR2_X1 U570 ( .A(n187), .B(n23), .ZN(SUM[15]) );
  XNOR2_X1 U571 ( .A(n196), .B(n24), .ZN(SUM[14]) );
  XNOR2_X1 U572 ( .A(n207), .B(n25), .ZN(SUM[13]) );
  XNOR2_X1 U573 ( .A(n214), .B(n26), .ZN(SUM[12]) );
  XNOR2_X1 U574 ( .A(n243), .B(n29), .ZN(SUM[9]) );
  XNOR2_X1 U575 ( .A(n232), .B(n28), .ZN(SUM[10]) );
  XNOR2_X1 U576 ( .A(n225), .B(n27), .ZN(SUM[11]) );
  XOR2_X1 U577 ( .A(n246), .B(n30), .Z(SUM[8]) );
  XOR2_X1 U578 ( .A(n257), .B(n32), .Z(SUM[6]) );
  XNOR2_X1 U579 ( .A(n254), .B(n31), .ZN(SUM[7]) );
  INV_X1 U580 ( .A(n205), .ZN(n300) );
  NOR2_X1 U581 ( .A1(n212), .A2(n205), .ZN(n203) );
  INV_X1 U582 ( .A(n436), .ZN(n290) );
  NOR2_X1 U583 ( .A1(n230), .A2(n223), .ZN(n221) );
  OAI21_X1 U584 ( .B1(n223), .B2(n231), .A(n224), .ZN(n222) );
  NAND2_X1 U585 ( .A1(A[11]), .A2(B[11]), .ZN(n224) );
  OAI21_X1 U586 ( .B1(n173), .B2(n177), .A(n174), .ZN(n172) );
  NAND2_X1 U587 ( .A1(A[29]), .A2(B[29]), .ZN(n62) );
  NOR2_X1 U588 ( .A1(A[29]), .A2(B[29]), .ZN(n61) );
  NOR2_X1 U589 ( .A1(A[31]), .A2(B[31]), .ZN(n39) );
  AOI21_X1 U590 ( .B1(n77), .B2(n98), .A(n78), .ZN(n440) );
  AOI21_X1 U591 ( .B1(n77), .B2(n98), .A(n78), .ZN(n5) );
  OAI21_X1 U592 ( .B1(n2), .B2(n102), .A(n103), .ZN(n101) );
  AOI21_X1 U593 ( .B1(n60), .B2(n416), .A(n49), .ZN(n47) );
  NOR2_X1 U594 ( .A1(n219), .A2(n181), .ZN(n179) );
  OAI21_X1 U595 ( .B1(n220), .B2(n181), .A(n182), .ZN(n180) );
  NAND2_X1 U596 ( .A1(A[13]), .A2(B[13]), .ZN(n206) );
  NAND2_X1 U597 ( .A1(B[23]), .A2(A[23]), .ZN(n118) );
  NOR2_X1 U598 ( .A1(B[23]), .A2(A[23]), .ZN(n117) );
  NAND2_X1 U599 ( .A1(A[17]), .A2(B[17]), .ZN(n174) );
  INV_X1 U600 ( .A(n51), .ZN(n49) );
  NAND2_X1 U601 ( .A1(n416), .A2(n51), .ZN(n8) );
  INV_X1 U602 ( .A(n5), .ZN(n76) );
  XNOR2_X1 U603 ( .A(n72), .B(n10), .ZN(SUM[28]) );
  NAND2_X1 U604 ( .A1(n171), .A2(n153), .ZN(n151) );
  NOR2_X1 U605 ( .A1(n176), .A2(n173), .ZN(n171) );
  NAND2_X1 U606 ( .A1(A[16]), .A2(B[16]), .ZN(n177) );
  NOR2_X1 U607 ( .A1(A[16]), .A2(B[16]), .ZN(n176) );
  XNOR2_X1 U608 ( .A(n81), .B(n11), .ZN(SUM[27]) );
  OAI21_X1 U609 ( .B1(n2), .B2(n82), .A(n83), .ZN(n81) );
  NOR2_X1 U610 ( .A1(n95), .A2(n424), .ZN(n84) );
  INV_X1 U611 ( .A(n95), .ZN(n93) );
  INV_X1 U612 ( .A(n97), .ZN(n95) );
  NAND2_X1 U613 ( .A1(A[30]), .A2(B[30]), .ZN(n51) );
  NAND2_X1 U614 ( .A1(A[28]), .A2(B[28]), .ZN(n71) );
  XNOR2_X1 U615 ( .A(n101), .B(n13), .ZN(SUM[25]) );
  OAI21_X1 U616 ( .B1(n205), .B2(n213), .A(n206), .ZN(n204) );
  INV_X1 U617 ( .A(n96), .ZN(n94) );
  INV_X1 U618 ( .A(n98), .ZN(n96) );
  INV_X1 U619 ( .A(n422), .ZN(n288) );
  NOR2_X1 U620 ( .A1(n106), .A2(n422), .ZN(n97) );
  NAND2_X1 U621 ( .A1(B[26]), .A2(A[26]), .ZN(n89) );
  NAND2_X1 U622 ( .A1(B[25]), .A2(A[25]), .ZN(n100) );
  INV_X1 U623 ( .A(n419), .ZN(n75) );
  NOR2_X1 U624 ( .A1(n6), .A2(n68), .ZN(n66) );
  NOR2_X1 U625 ( .A1(n6), .A2(n425), .ZN(n55) );
  NOR2_X1 U626 ( .A1(n419), .A2(n46), .ZN(n44) );
  NAND2_X1 U627 ( .A1(n97), .A2(n77), .ZN(n6) );
  XOR2_X1 U628 ( .A(n1), .B(n22), .Z(SUM[16]) );
  OAI21_X1 U629 ( .B1(n1), .B2(n120), .A(n121), .ZN(n119) );
  OAI21_X1 U630 ( .B1(n1), .B2(n129), .A(n130), .ZN(n128) );
  OAI21_X1 U631 ( .B1(n1), .B2(n140), .A(n141), .ZN(n139) );
  OAI21_X1 U632 ( .B1(n1), .B2(n151), .A(n148), .ZN(n146) );
  OAI21_X1 U633 ( .B1(n1), .B2(n158), .A(n159), .ZN(n157) );
  OAI21_X1 U634 ( .B1(n1), .B2(n169), .A(n170), .ZN(n164) );
  OAI21_X1 U635 ( .B1(n1), .B2(n176), .A(n177), .ZN(n175) );
  AOI21_X1 U636 ( .B1(n183), .B2(n204), .A(n184), .ZN(n182) );
  OAI21_X1 U637 ( .B1(n155), .B2(n163), .A(n156), .ZN(n154) );
  XNOR2_X1 U638 ( .A(n52), .B(n8), .ZN(SUM[30]) );
  NAND2_X1 U639 ( .A1(B[27]), .A2(A[27]), .ZN(n80) );
  XNOR2_X1 U640 ( .A(n63), .B(n9), .ZN(SUM[29]) );
  INV_X1 U641 ( .A(n424), .ZN(n87) );
  OAI21_X1 U642 ( .B1(n2), .B2(n91), .A(n92), .ZN(n90) );
  OAI21_X1 U643 ( .B1(n2), .B2(n42), .A(n43), .ZN(n41) );
  NAND2_X1 U644 ( .A1(n59), .A2(n416), .ZN(n46) );
  INV_X1 U645 ( .A(n426), .ZN(n284) );
  OAI21_X1 U646 ( .B1(n96), .B2(n424), .A(n89), .ZN(n85) );
  NAND2_X1 U647 ( .A1(n4), .A2(n75), .ZN(n73) );
  NAND2_X1 U648 ( .A1(n438), .A2(n55), .ZN(n53) );
  NAND2_X1 U649 ( .A1(n4), .A2(n66), .ZN(n64) );
  NAND2_X1 U650 ( .A1(n4), .A2(n44), .ZN(n42) );
  NAND2_X1 U651 ( .A1(n438), .A2(n93), .ZN(n91) );
  NAND2_X1 U652 ( .A1(n4), .A2(n84), .ZN(n82) );
  NAND2_X1 U653 ( .A1(n438), .A2(n104), .ZN(n102) );
  OAI21_X1 U654 ( .B1(n2), .B2(n73), .A(n74), .ZN(n72) );
  OAI21_X1 U655 ( .B1(n2), .B2(n53), .A(n54), .ZN(n52) );
  NOR2_X1 U656 ( .A1(n70), .A2(n61), .ZN(n59) );
  INV_X1 U657 ( .A(n70), .ZN(n69) );
  NOR2_X1 U658 ( .A1(A[28]), .A2(B[28]), .ZN(n70) );
  XNOR2_X1 U659 ( .A(n41), .B(n7), .ZN(SUM[31]) );
  OAI21_X1 U660 ( .B1(n2), .B2(n64), .A(n65), .ZN(n63) );
  OAI21_X1 U661 ( .B1(n99), .B2(n107), .A(n100), .ZN(n98) );
  NOR2_X1 U662 ( .A1(n194), .A2(n185), .ZN(n183) );
  OAI21_X1 U663 ( .B1(n185), .B2(n195), .A(n186), .ZN(n184) );
  OAI21_X1 U664 ( .B1(n152), .B2(n113), .A(n114), .ZN(n112) );
  NOR2_X1 U665 ( .A1(n113), .A2(n151), .ZN(n111) );
  AOI21_X1 U666 ( .B1(n437), .B2(n93), .A(n94), .ZN(n92) );
  AOI21_X1 U667 ( .B1(n3), .B2(n104), .A(n105), .ZN(n103) );
  AOI21_X1 U668 ( .B1(n437), .B2(n75), .A(n76), .ZN(n74) );
  AOI21_X1 U669 ( .B1(n3), .B2(n84), .A(n85), .ZN(n83) );
  AOI21_X1 U670 ( .B1(n437), .B2(n44), .A(n45), .ZN(n43) );
  AOI21_X1 U671 ( .B1(n3), .B2(n55), .A(n56), .ZN(n54) );
  AOI21_X1 U672 ( .B1(n437), .B2(n66), .A(n67), .ZN(n65) );
  NAND2_X1 U673 ( .A1(n115), .A2(n135), .ZN(n113) );
  NOR2_X1 U674 ( .A1(n144), .A2(n137), .ZN(n135) );
  OAI21_X1 U675 ( .B1(n440), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U676 ( .B1(n5), .B2(n425), .A(n58), .ZN(n56) );
  OAI21_X1 U677 ( .B1(n440), .B2(n68), .A(n71), .ZN(n67) );
  OAI21_X1 U678 ( .B1(n427), .B2(n89), .A(n80), .ZN(n78) );
  OAI21_X1 U679 ( .B1(n434), .B2(n127), .A(n118), .ZN(n116) );
  NOR2_X1 U680 ( .A1(n117), .A2(n126), .ZN(n115) );
  AOI21_X1 U681 ( .B1(n136), .B2(n115), .A(n116), .ZN(n114) );
  OAI21_X1 U682 ( .B1(n431), .B2(n145), .A(n138), .ZN(n136) );
  NAND2_X1 U683 ( .A1(A[21]), .A2(B[21]), .ZN(n138) );
  NOR2_X1 U684 ( .A1(B[21]), .A2(A[21]), .ZN(n137) );
endmodule


module datapath_DW01_add_13 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n40, n41, n42, n43, n44, n45, n46,
         n47, n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n88, n89, n90, n91, n92,
         n93, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n126, n127, n128, n129,
         n130, n131, n133, n134, n135, n136, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n193, n194, n195, n196, n197, n198, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n234, n237, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n281, n284, n286, n287, n290, n291,
         n292, n294, n296, n297, n298, n300, n302, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n416, n417, n418, n419, n420, n421,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446;

  CLKBUF_X1 U349 ( .A(n420), .Z(n416) );
  CLKBUF_X1 U350 ( .A(n88), .Z(n417) );
  CLKBUF_X1 U351 ( .A(n126), .Z(n418) );
  CLKBUF_X1 U352 ( .A(n135), .Z(n419) );
  NOR2_X1 U353 ( .A1(B[21]), .A2(A[21]), .ZN(n420) );
  OR2_X1 U354 ( .A1(A[30]), .A2(B[30]), .ZN(n421) );
  AND2_X1 U355 ( .A1(n425), .A2(n281), .ZN(SUM[0]) );
  NOR2_X1 U356 ( .A1(A[26]), .A2(n431), .ZN(n423) );
  NOR2_X1 U357 ( .A1(A[22]), .A2(n436), .ZN(n424) );
  OR2_X1 U358 ( .A1(A[0]), .A2(B[0]), .ZN(n425) );
  CLKBUF_X1 U359 ( .A(n112), .Z(n443) );
  CLKBUF_X1 U360 ( .A(n61), .Z(n426) );
  BUF_X1 U361 ( .A(n112), .Z(n444) );
  CLKBUF_X1 U362 ( .A(B[25]), .Z(n427) );
  CLKBUF_X1 U363 ( .A(n144), .Z(n428) );
  NOR2_X1 U364 ( .A1(B[27]), .A2(A[27]), .ZN(n429) );
  OR2_X1 U365 ( .A1(n427), .A2(A[25]), .ZN(n430) );
  NOR2_X1 U366 ( .A1(B[25]), .A2(A[25]), .ZN(n99) );
  CLKBUF_X1 U367 ( .A(B[26]), .Z(n431) );
  CLKBUF_X1 U368 ( .A(n98), .Z(n432) );
  NOR2_X1 U369 ( .A1(n126), .A2(n435), .ZN(n433) );
  NOR2_X1 U370 ( .A1(A[19]), .A2(B[19]), .ZN(n434) );
  NOR2_X1 U371 ( .A1(B[23]), .A2(A[23]), .ZN(n435) );
  CLKBUF_X1 U372 ( .A(B[22]), .Z(n436) );
  NAND2_X1 U373 ( .A1(A[24]), .A2(B[24]), .ZN(n107) );
  NAND2_X1 U374 ( .A1(n98), .A2(n77), .ZN(n437) );
  INV_X1 U375 ( .A(n78), .ZN(n438) );
  AND2_X2 U376 ( .A1(n437), .A2(n438), .ZN(n5) );
  CLKBUF_X1 U377 ( .A(n429), .Z(n439) );
  CLKBUF_X1 U378 ( .A(n136), .Z(n440) );
  NOR2_X1 U379 ( .A1(B[21]), .A2(A[21]), .ZN(n441) );
  CLKBUF_X1 U380 ( .A(n435), .Z(n442) );
  BUF_X1 U381 ( .A(n111), .Z(n445) );
  NOR2_X1 U382 ( .A1(A[10]), .A2(B[10]), .ZN(n230) );
  NOR2_X1 U383 ( .A1(A[4]), .A2(B[4]), .ZN(n265) );
  NOR2_X1 U384 ( .A1(A[12]), .A2(B[12]), .ZN(n212) );
  NOR2_X1 U385 ( .A1(A[3]), .A2(B[3]), .ZN(n271) );
  NOR2_X1 U386 ( .A1(A[5]), .A2(B[5]), .ZN(n260) );
  NOR2_X1 U387 ( .A1(A[7]), .A2(B[7]), .ZN(n252) );
  NOR2_X1 U388 ( .A1(A[8]), .A2(B[8]), .ZN(n244) );
  NOR2_X1 U389 ( .A1(A[6]), .A2(B[6]), .ZN(n255) );
  NOR2_X1 U390 ( .A1(A[2]), .A2(B[2]), .ZN(n274) );
  NOR2_X1 U391 ( .A1(A[1]), .A2(B[1]), .ZN(n278) );
  INV_X1 U392 ( .A(n150), .ZN(n148) );
  INV_X1 U393 ( .A(n149), .ZN(n147) );
  INV_X1 U394 ( .A(n219), .ZN(n217) );
  OAI21_X1 U395 ( .B1(n246), .B2(n197), .A(n198), .ZN(n196) );
  AOI21_X1 U396 ( .B1(n218), .B2(n203), .A(n200), .ZN(n198) );
  NAND2_X1 U397 ( .A1(n217), .A2(n203), .ZN(n197) );
  OAI21_X1 U398 ( .B1(n246), .B2(n219), .A(n220), .ZN(n214) );
  OAI21_X1 U399 ( .B1(n246), .B2(n237), .A(n234), .ZN(n232) );
  INV_X1 U400 ( .A(n240), .ZN(n234) );
  INV_X1 U401 ( .A(n151), .ZN(n149) );
  BUF_X1 U402 ( .A(n178), .Z(n1) );
  BUF_X1 U403 ( .A(n178), .Z(n2) );
  BUF_X1 U404 ( .A(n111), .Z(n4) );
  INV_X1 U405 ( .A(n202), .ZN(n200) );
  INV_X1 U406 ( .A(n247), .ZN(n246) );
  AOI21_X1 U407 ( .B1(n247), .B2(n179), .A(n180), .ZN(n178) );
  NOR2_X1 U408 ( .A1(n219), .A2(n181), .ZN(n179) );
  AOI21_X1 U409 ( .B1(n267), .B2(n258), .A(n259), .ZN(n257) );
  NOR2_X1 U410 ( .A1(n201), .A2(n194), .ZN(n190) );
  NOR2_X1 U411 ( .A1(n95), .A2(n423), .ZN(n84) );
  INV_X1 U412 ( .A(n95), .ZN(n93) );
  INV_X1 U413 ( .A(n6), .ZN(n75) );
  INV_X1 U414 ( .A(n203), .ZN(n201) );
  INV_X1 U415 ( .A(n220), .ZN(n218) );
  NAND2_X1 U416 ( .A1(n239), .A2(n221), .ZN(n219) );
  INV_X1 U417 ( .A(n268), .ZN(n267) );
  INV_X1 U418 ( .A(n204), .ZN(n202) );
  INV_X1 U419 ( .A(n170), .ZN(n168) );
  INV_X1 U420 ( .A(n172), .ZN(n170) );
  INV_X1 U421 ( .A(n277), .ZN(n276) );
  INV_X1 U422 ( .A(n169), .ZN(n167) );
  INV_X1 U423 ( .A(n239), .ZN(n237) );
  INV_X1 U424 ( .A(n419), .ZN(n133) );
  INV_X1 U425 ( .A(n59), .ZN(n57) );
  OAI21_X1 U426 ( .B1(n241), .B2(n245), .A(n242), .ZN(n240) );
  NOR2_X1 U427 ( .A1(n230), .A2(n223), .ZN(n221) );
  NOR2_X1 U428 ( .A1(n244), .A2(n241), .ZN(n239) );
  OAI21_X1 U429 ( .B1(n205), .B2(n213), .A(n206), .ZN(n204) );
  NAND2_X1 U430 ( .A1(n167), .A2(n160), .ZN(n158) );
  AOI21_X1 U431 ( .B1(n168), .B2(n160), .A(n161), .ZN(n159) );
  INV_X1 U432 ( .A(n162), .ZN(n160) );
  AOI21_X1 U433 ( .B1(n150), .B2(n142), .A(n143), .ZN(n141) );
  NAND2_X1 U434 ( .A1(n149), .A2(n142), .ZN(n140) );
  AOI21_X1 U435 ( .B1(n269), .B2(n277), .A(n270), .ZN(n268) );
  OAI21_X1 U436 ( .B1(n271), .B2(n275), .A(n272), .ZN(n270) );
  NOR2_X1 U437 ( .A1(n274), .A2(n271), .ZN(n269) );
  OAI21_X1 U438 ( .B1(n260), .B2(n266), .A(n261), .ZN(n259) );
  OAI21_X1 U439 ( .B1(n278), .B2(n281), .A(n279), .ZN(n277) );
  NOR2_X1 U440 ( .A1(n265), .A2(n260), .ZN(n258) );
  AOI21_X1 U441 ( .B1(n221), .B2(n240), .A(n222), .ZN(n220) );
  INV_X1 U442 ( .A(n51), .ZN(n49) );
  OAI21_X1 U443 ( .B1(n268), .B2(n248), .A(n249), .ZN(n247) );
  AOI21_X1 U444 ( .B1(n250), .B2(n259), .A(n251), .ZN(n249) );
  NAND2_X1 U445 ( .A1(n258), .A2(n250), .ZN(n248) );
  NOR2_X1 U446 ( .A1(n255), .A2(n252), .ZN(n250) );
  NOR2_X1 U447 ( .A1(n70), .A2(n61), .ZN(n59) );
  OAI21_X1 U448 ( .B1(n252), .B2(n256), .A(n253), .ZN(n251) );
  AOI21_X1 U449 ( .B1(n267), .B2(n309), .A(n264), .ZN(n262) );
  INV_X1 U450 ( .A(n266), .ZN(n264) );
  INV_X1 U451 ( .A(n428), .ZN(n142) );
  BUF_X1 U452 ( .A(n112), .Z(n3) );
  OAI21_X1 U453 ( .B1(n257), .B2(n255), .A(n256), .ZN(n254) );
  OAI21_X1 U454 ( .B1(n246), .B2(n244), .A(n245), .ZN(n243) );
  OAI21_X1 U455 ( .B1(n276), .B2(n274), .A(n275), .ZN(n273) );
  OAI21_X1 U456 ( .B1(n246), .B2(n188), .A(n189), .ZN(n187) );
  AOI21_X1 U457 ( .B1(n190), .B2(n218), .A(n191), .ZN(n189) );
  NAND2_X1 U458 ( .A1(n190), .A2(n217), .ZN(n188) );
  OAI21_X1 U459 ( .B1(n202), .B2(n194), .A(n195), .ZN(n191) );
  OAI21_X1 U460 ( .B1(n246), .B2(n208), .A(n209), .ZN(n207) );
  AOI21_X1 U461 ( .B1(n218), .B2(n210), .A(n211), .ZN(n209) );
  NAND2_X1 U462 ( .A1(n217), .A2(n210), .ZN(n208) );
  INV_X1 U463 ( .A(n213), .ZN(n211) );
  OAI21_X1 U464 ( .B1(n246), .B2(n226), .A(n227), .ZN(n225) );
  AOI21_X1 U465 ( .B1(n240), .B2(n228), .A(n229), .ZN(n227) );
  NAND2_X1 U466 ( .A1(n239), .A2(n228), .ZN(n226) );
  INV_X1 U467 ( .A(n231), .ZN(n229) );
  INV_X1 U468 ( .A(n212), .ZN(n210) );
  OAI21_X1 U469 ( .B1(n96), .B2(n423), .A(n89), .ZN(n85) );
  INV_X1 U470 ( .A(n230), .ZN(n228) );
  INV_X1 U471 ( .A(n442), .ZN(n290) );
  NAND2_X1 U472 ( .A1(n160), .A2(n163), .ZN(n20) );
  INV_X1 U473 ( .A(n69), .ZN(n68) );
  INV_X1 U474 ( .A(n70), .ZN(n69) );
  INV_X1 U475 ( .A(n163), .ZN(n161) );
  INV_X1 U476 ( .A(n194), .ZN(n193) );
  INV_X1 U477 ( .A(n417), .ZN(n287) );
  NAND2_X1 U478 ( .A1(n300), .A2(n206), .ZN(n25) );
  INV_X1 U479 ( .A(n205), .ZN(n300) );
  NAND2_X1 U480 ( .A1(n309), .A2(n266), .ZN(n34) );
  INV_X1 U481 ( .A(n265), .ZN(n309) );
  NAND2_X1 U482 ( .A1(n307), .A2(n256), .ZN(n32) );
  INV_X1 U483 ( .A(n255), .ZN(n307) );
  NAND2_X1 U484 ( .A1(n210), .A2(n213), .ZN(n26) );
  NAND2_X1 U485 ( .A1(n302), .A2(n224), .ZN(n27) );
  INV_X1 U486 ( .A(n223), .ZN(n302) );
  NAND2_X1 U487 ( .A1(n296), .A2(n174), .ZN(n21) );
  INV_X1 U488 ( .A(n173), .ZN(n296) );
  NAND2_X1 U489 ( .A1(n305), .A2(n245), .ZN(n30) );
  INV_X1 U490 ( .A(n244), .ZN(n305) );
  NAND2_X1 U491 ( .A1(n306), .A2(n253), .ZN(n31) );
  INV_X1 U492 ( .A(n252), .ZN(n306) );
  NAND2_X1 U493 ( .A1(n308), .A2(n261), .ZN(n33) );
  INV_X1 U494 ( .A(n260), .ZN(n308) );
  NAND2_X1 U495 ( .A1(n298), .A2(n186), .ZN(n23) );
  INV_X1 U496 ( .A(n185), .ZN(n298) );
  NAND2_X1 U497 ( .A1(n311), .A2(n275), .ZN(n36) );
  INV_X1 U498 ( .A(n274), .ZN(n311) );
  NAND2_X1 U499 ( .A1(n228), .A2(n231), .ZN(n28) );
  NAND2_X1 U500 ( .A1(n193), .A2(n195), .ZN(n24) );
  INV_X1 U501 ( .A(n426), .ZN(n284) );
  INV_X1 U502 ( .A(n418), .ZN(n291) );
  NAND2_X1 U503 ( .A1(n310), .A2(n272), .ZN(n35) );
  INV_X1 U504 ( .A(n271), .ZN(n310) );
  NAND2_X1 U505 ( .A1(n104), .A2(n107), .ZN(n14) );
  XNOR2_X1 U506 ( .A(n128), .B(n16), .ZN(SUM[22]) );
  NAND2_X1 U507 ( .A1(n291), .A2(n127), .ZN(n16) );
  XNOR2_X1 U508 ( .A(n119), .B(n15), .ZN(SUM[23]) );
  NAND2_X1 U509 ( .A1(n290), .A2(n118), .ZN(n15) );
  XNOR2_X1 U510 ( .A(n139), .B(n17), .ZN(SUM[21]) );
  NAND2_X1 U511 ( .A1(n292), .A2(n138), .ZN(n17) );
  XNOR2_X1 U512 ( .A(n146), .B(n18), .ZN(SUM[20]) );
  NAND2_X1 U513 ( .A1(n304), .A2(n242), .ZN(n29) );
  NAND2_X1 U514 ( .A1(n312), .A2(n279), .ZN(n37) );
  INV_X1 U515 ( .A(n278), .ZN(n312) );
  NAND2_X1 U516 ( .A1(n294), .A2(n156), .ZN(n19) );
  INV_X1 U517 ( .A(n434), .ZN(n294) );
  INV_X1 U518 ( .A(n439), .ZN(n286) );
  NAND2_X1 U519 ( .A1(n297), .A2(n177), .ZN(n22) );
  INV_X1 U520 ( .A(n107), .ZN(n105) );
  NOR2_X1 U521 ( .A1(A[28]), .A2(B[28]), .ZN(n70) );
  NOR2_X1 U522 ( .A1(A[29]), .A2(B[29]), .ZN(n61) );
  NOR2_X1 U523 ( .A1(A[11]), .A2(B[11]), .ZN(n223) );
  NOR2_X1 U524 ( .A1(A[18]), .A2(B[18]), .ZN(n162) );
  NOR2_X1 U525 ( .A1(B[22]), .A2(A[22]), .ZN(n126) );
  NOR2_X1 U526 ( .A1(B[20]), .A2(A[20]), .ZN(n144) );
  NOR2_X1 U527 ( .A1(A[13]), .A2(B[13]), .ZN(n205) );
  NOR2_X1 U528 ( .A1(A[19]), .A2(B[19]), .ZN(n155) );
  NOR2_X1 U529 ( .A1(B[27]), .A2(A[27]), .ZN(n79) );
  NOR2_X1 U530 ( .A1(A[9]), .A2(B[9]), .ZN(n241) );
  NOR2_X1 U531 ( .A1(B[26]), .A2(A[26]), .ZN(n88) );
  NAND2_X1 U532 ( .A1(B[26]), .A2(A[26]), .ZN(n89) );
  NOR2_X1 U533 ( .A1(A[24]), .A2(B[24]), .ZN(n106) );
  NOR2_X1 U534 ( .A1(A[14]), .A2(B[14]), .ZN(n194) );
  NOR2_X1 U535 ( .A1(A[15]), .A2(B[15]), .ZN(n185) );
  NAND2_X1 U536 ( .A1(A[4]), .A2(B[4]), .ZN(n266) );
  NAND2_X1 U537 ( .A1(A[6]), .A2(B[6]), .ZN(n256) );
  NAND2_X1 U538 ( .A1(A[12]), .A2(B[12]), .ZN(n213) );
  NAND2_X1 U539 ( .A1(A[8]), .A2(B[8]), .ZN(n245) );
  XOR2_X1 U540 ( .A(n257), .B(n32), .Z(SUM[6]) );
  NAND2_X1 U541 ( .A1(A[2]), .A2(B[2]), .ZN(n275) );
  NAND2_X1 U542 ( .A1(A[5]), .A2(B[5]), .ZN(n261) );
  NAND2_X1 U543 ( .A1(A[7]), .A2(B[7]), .ZN(n253) );
  NAND2_X1 U544 ( .A1(A[0]), .A2(B[0]), .ZN(n281) );
  NAND2_X1 U545 ( .A1(A[30]), .A2(B[30]), .ZN(n51) );
  XNOR2_X1 U546 ( .A(n243), .B(n29), .ZN(SUM[9]) );
  NAND2_X1 U547 ( .A1(A[15]), .A2(B[15]), .ZN(n186) );
  NAND2_X1 U548 ( .A1(A[14]), .A2(B[14]), .ZN(n195) );
  NAND2_X1 U549 ( .A1(A[10]), .A2(B[10]), .ZN(n231) );
  NAND2_X1 U550 ( .A1(A[1]), .A2(B[1]), .ZN(n279) );
  NAND2_X1 U551 ( .A1(A[3]), .A2(B[3]), .ZN(n272) );
  NAND2_X1 U552 ( .A1(A[9]), .A2(B[9]), .ZN(n242) );
  NAND2_X1 U553 ( .A1(A[31]), .A2(B[31]), .ZN(n40) );
  NAND2_X1 U554 ( .A1(A[29]), .A2(B[29]), .ZN(n62) );
  NAND2_X1 U555 ( .A1(A[16]), .A2(B[16]), .ZN(n177) );
  NAND2_X1 U556 ( .A1(n446), .A2(n40), .ZN(n7) );
  NAND2_X1 U557 ( .A1(n421), .A2(n51), .ZN(n8) );
  NAND2_X1 U558 ( .A1(n284), .A2(n62), .ZN(n9) );
  NAND2_X1 U559 ( .A1(n286), .A2(n80), .ZN(n11) );
  XOR2_X1 U560 ( .A(n37), .B(n281), .Z(SUM[1]) );
  XOR2_X1 U561 ( .A(n276), .B(n36), .Z(SUM[2]) );
  XNOR2_X1 U562 ( .A(n273), .B(n35), .ZN(SUM[3]) );
  XNOR2_X1 U563 ( .A(n267), .B(n34), .ZN(SUM[4]) );
  XOR2_X1 U564 ( .A(n262), .B(n33), .Z(SUM[5]) );
  NAND2_X1 U565 ( .A1(n287), .A2(n89), .ZN(n12) );
  NAND2_X1 U566 ( .A1(n69), .A2(n71), .ZN(n10) );
  NAND2_X1 U567 ( .A1(n430), .A2(n100), .ZN(n13) );
  XNOR2_X1 U568 ( .A(n175), .B(n21), .ZN(SUM[17]) );
  XNOR2_X1 U569 ( .A(n157), .B(n19), .ZN(SUM[19]) );
  XNOR2_X1 U570 ( .A(n164), .B(n20), .ZN(SUM[18]) );
  XNOR2_X1 U571 ( .A(n187), .B(n23), .ZN(SUM[15]) );
  XNOR2_X1 U572 ( .A(n207), .B(n25), .ZN(SUM[13]) );
  XNOR2_X1 U573 ( .A(n196), .B(n24), .ZN(SUM[14]) );
  XNOR2_X1 U574 ( .A(n214), .B(n26), .ZN(SUM[12]) );
  XNOR2_X1 U575 ( .A(n225), .B(n27), .ZN(SUM[11]) );
  XNOR2_X1 U576 ( .A(n232), .B(n28), .ZN(SUM[10]) );
  XOR2_X1 U577 ( .A(n246), .B(n30), .Z(SUM[8]) );
  XNOR2_X1 U578 ( .A(n254), .B(n31), .ZN(SUM[7]) );
  OR2_X1 U579 ( .A1(A[31]), .A2(B[31]), .ZN(n446) );
  NAND2_X1 U580 ( .A1(B[22]), .A2(A[22]), .ZN(n127) );
  INV_X1 U581 ( .A(n416), .ZN(n292) );
  NOR2_X1 U582 ( .A1(n144), .A2(n441), .ZN(n135) );
  INV_X1 U583 ( .A(n5), .ZN(n76) );
  NAND2_X1 U584 ( .A1(A[19]), .A2(B[19]), .ZN(n156) );
  INV_X1 U585 ( .A(n432), .ZN(n96) );
  NAND2_X1 U586 ( .A1(A[28]), .A2(B[28]), .ZN(n71) );
  NAND2_X1 U587 ( .A1(n149), .A2(n131), .ZN(n129) );
  XNOR2_X1 U588 ( .A(n108), .B(n14), .ZN(SUM[24]) );
  NOR2_X1 U589 ( .A1(n88), .A2(n79), .ZN(n77) );
  XNOR2_X1 U590 ( .A(n90), .B(n12), .ZN(SUM[26]) );
  XNOR2_X1 U591 ( .A(n101), .B(n13), .ZN(SUM[25]) );
  XNOR2_X1 U592 ( .A(n72), .B(n10), .ZN(SUM[28]) );
  XNOR2_X1 U593 ( .A(n63), .B(n9), .ZN(SUM[29]) );
  NAND2_X1 U594 ( .A1(n97), .A2(n77), .ZN(n6) );
  XOR2_X1 U595 ( .A(n1), .B(n22), .Z(SUM[16]) );
  OAI21_X1 U596 ( .B1(n1), .B2(n140), .A(n141), .ZN(n139) );
  OAI21_X1 U597 ( .B1(n1), .B2(n158), .A(n159), .ZN(n157) );
  OAI21_X1 U598 ( .B1(n1), .B2(n169), .A(n170), .ZN(n164) );
  OAI21_X1 U599 ( .B1(n1), .B2(n129), .A(n130), .ZN(n128) );
  OAI21_X1 U600 ( .B1(n1), .B2(n120), .A(n121), .ZN(n119) );
  OAI21_X1 U601 ( .B1(n1), .B2(n147), .A(n148), .ZN(n146) );
  NAND2_X1 U602 ( .A1(n122), .A2(n149), .ZN(n120) );
  AOI21_X1 U603 ( .B1(n122), .B2(n150), .A(n123), .ZN(n121) );
  NOR2_X1 U604 ( .A1(n133), .A2(n424), .ZN(n122) );
  XNOR2_X1 U605 ( .A(n52), .B(n8), .ZN(SUM[30]) );
  AOI21_X1 U606 ( .B1(n150), .B2(n131), .A(n440), .ZN(n130) );
  INV_X1 U607 ( .A(n133), .ZN(n131) );
  INV_X1 U608 ( .A(n241), .ZN(n304) );
  OAI21_X1 U609 ( .B1(n2), .B2(n109), .A(n110), .ZN(n108) );
  INV_X1 U610 ( .A(n4), .ZN(n109) );
  INV_X1 U611 ( .A(n3), .ZN(n110) );
  NAND2_X1 U612 ( .A1(n203), .A2(n183), .ZN(n181) );
  NAND2_X1 U613 ( .A1(A[13]), .A2(B[13]), .ZN(n206) );
  AOI21_X1 U614 ( .B1(n60), .B2(n421), .A(n49), .ZN(n47) );
  INV_X1 U615 ( .A(n60), .ZN(n58) );
  NOR2_X1 U616 ( .A1(n113), .A2(n151), .ZN(n111) );
  OAI21_X1 U617 ( .B1(n134), .B2(n424), .A(n127), .ZN(n123) );
  INV_X1 U618 ( .A(n145), .ZN(n143) );
  NAND2_X1 U619 ( .A1(n142), .A2(n145), .ZN(n18) );
  NOR2_X1 U620 ( .A1(A[23]), .A2(B[23]), .ZN(n117) );
  NAND2_X1 U621 ( .A1(B[23]), .A2(A[23]), .ZN(n118) );
  NOR2_X1 U622 ( .A1(n6), .A2(n46), .ZN(n44) );
  NOR2_X1 U623 ( .A1(n6), .A2(n68), .ZN(n66) );
  NOR2_X1 U624 ( .A1(n6), .A2(n57), .ZN(n55) );
  OAI21_X1 U625 ( .B1(n2), .B2(n82), .A(n83), .ZN(n81) );
  OAI21_X1 U626 ( .B1(n223), .B2(n231), .A(n224), .ZN(n222) );
  NAND2_X1 U627 ( .A1(A[11]), .A2(B[11]), .ZN(n224) );
  NAND2_X1 U628 ( .A1(n59), .A2(n421), .ZN(n46) );
  OAI21_X1 U629 ( .B1(n2), .B2(n91), .A(n92), .ZN(n90) );
  INV_X1 U630 ( .A(n106), .ZN(n104) );
  NAND2_X1 U631 ( .A1(n171), .A2(n153), .ZN(n151) );
  INV_X1 U632 ( .A(n171), .ZN(n169) );
  NOR2_X1 U633 ( .A1(n176), .A2(n173), .ZN(n171) );
  INV_X1 U634 ( .A(n176), .ZN(n297) );
  OAI21_X1 U635 ( .B1(n1), .B2(n176), .A(n177), .ZN(n175) );
  NOR2_X1 U636 ( .A1(A[16]), .A2(B[16]), .ZN(n176) );
  OAI21_X1 U637 ( .B1(n2), .B2(n102), .A(n103), .ZN(n101) );
  OAI21_X1 U638 ( .B1(n220), .B2(n181), .A(n182), .ZN(n180) );
  NAND2_X1 U639 ( .A1(A[18]), .A2(B[18]), .ZN(n163) );
  OAI21_X1 U640 ( .B1(n2), .B2(n42), .A(n43), .ZN(n41) );
  NAND2_X1 U641 ( .A1(A[27]), .A2(B[27]), .ZN(n80) );
  OAI21_X1 U642 ( .B1(n2), .B2(n73), .A(n74), .ZN(n72) );
  INV_X1 U643 ( .A(n97), .ZN(n95) );
  NAND2_X1 U644 ( .A1(B[25]), .A2(A[25]), .ZN(n100) );
  AOI21_X1 U645 ( .B1(n3), .B2(n84), .A(n85), .ZN(n83) );
  NAND2_X1 U646 ( .A1(B[20]), .A2(A[20]), .ZN(n145) );
  INV_X1 U647 ( .A(n440), .ZN(n134) );
  AOI21_X1 U648 ( .B1(n183), .B2(n204), .A(n184), .ZN(n182) );
  NOR2_X1 U649 ( .A1(n212), .A2(n205), .ZN(n203) );
  OAI21_X1 U650 ( .B1(n2), .B2(n64), .A(n65), .ZN(n63) );
  INV_X1 U651 ( .A(n152), .ZN(n150) );
  NOR2_X1 U652 ( .A1(n162), .A2(n434), .ZN(n153) );
  OAI21_X1 U653 ( .B1(n155), .B2(n163), .A(n156), .ZN(n154) );
  NAND2_X1 U654 ( .A1(n4), .A2(n55), .ZN(n53) );
  NAND2_X1 U655 ( .A1(n445), .A2(n84), .ZN(n82) );
  NAND2_X1 U656 ( .A1(n4), .A2(n44), .ZN(n42) );
  NAND2_X1 U657 ( .A1(n445), .A2(n93), .ZN(n91) );
  NAND2_X1 U658 ( .A1(n445), .A2(n75), .ZN(n73) );
  NAND2_X1 U659 ( .A1(n445), .A2(n66), .ZN(n64) );
  NAND2_X1 U660 ( .A1(n4), .A2(n104), .ZN(n102) );
  OAI21_X1 U661 ( .B1(n152), .B2(n113), .A(n114), .ZN(n112) );
  AOI21_X1 U662 ( .B1(n153), .B2(n172), .A(n154), .ZN(n152) );
  OAI21_X1 U663 ( .B1(n173), .B2(n177), .A(n174), .ZN(n172) );
  NAND2_X1 U664 ( .A1(A[17]), .A2(B[17]), .ZN(n174) );
  NOR2_X1 U665 ( .A1(A[17]), .A2(B[17]), .ZN(n173) );
  OAI21_X1 U666 ( .B1(n2), .B2(n53), .A(n54), .ZN(n52) );
  OAI21_X1 U667 ( .B1(n61), .B2(n71), .A(n62), .ZN(n60) );
  XNOR2_X1 U668 ( .A(n41), .B(n7), .ZN(SUM[31]) );
  OAI21_X1 U669 ( .B1(n99), .B2(n107), .A(n100), .ZN(n98) );
  NOR2_X1 U670 ( .A1(n106), .A2(n99), .ZN(n97) );
  NOR2_X1 U671 ( .A1(n194), .A2(n185), .ZN(n183) );
  OAI21_X1 U672 ( .B1(n185), .B2(n195), .A(n186), .ZN(n184) );
  AOI21_X1 U673 ( .B1(n3), .B2(n66), .A(n67), .ZN(n65) );
  AOI21_X1 U674 ( .B1(n443), .B2(n55), .A(n56), .ZN(n54) );
  AOI21_X1 U675 ( .B1(n443), .B2(n75), .A(n76), .ZN(n74) );
  AOI21_X1 U676 ( .B1(n444), .B2(n44), .A(n45), .ZN(n43) );
  AOI21_X1 U677 ( .B1(n444), .B2(n104), .A(n105), .ZN(n103) );
  AOI21_X1 U678 ( .B1(n444), .B2(n93), .A(n432), .ZN(n92) );
  OAI21_X1 U679 ( .B1(n5), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U680 ( .B1(n5), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U681 ( .B1(n5), .B2(n68), .A(n71), .ZN(n67) );
  OAI21_X1 U682 ( .B1(n429), .B2(n89), .A(n80), .ZN(n78) );
  OAI21_X1 U683 ( .B1(n117), .B2(n127), .A(n118), .ZN(n116) );
  NOR2_X1 U684 ( .A1(n435), .A2(n126), .ZN(n115) );
  XNOR2_X1 U685 ( .A(n81), .B(n11), .ZN(SUM[27]) );
  NAND2_X1 U686 ( .A1(n135), .A2(n433), .ZN(n113) );
  AOI21_X1 U687 ( .B1(n136), .B2(n115), .A(n116), .ZN(n114) );
  OAI21_X1 U688 ( .B1(n145), .B2(n420), .A(n138), .ZN(n136) );
  NAND2_X1 U689 ( .A1(B[21]), .A2(A[21]), .ZN(n138) );
endmodule


module datapath_DW01_add_14 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n40, n41, n42, n43, n45, n46, n47,
         n49, n51, n52, n53, n54, n55, n56, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n88, n89, n90, n91, n92, n93,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n193, n194, n195, n196, n197, n198, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n234, n237, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n281, n284, n286, n288, n290,
         n292, n294, n296, n297, n300, n302, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n444, n445;

  BUF_X1 U349 ( .A(n112), .Z(n416) );
  CLKBUF_X1 U350 ( .A(n112), .Z(n3) );
  CLKBUF_X1 U351 ( .A(n71), .Z(n417) );
  CLKBUF_X1 U352 ( .A(n89), .Z(n418) );
  NOR2_X1 U353 ( .A1(n6), .A2(n46), .ZN(n419) );
  OR2_X1 U354 ( .A1(A[30]), .A2(B[30]), .ZN(n420) );
  OR2_X1 U355 ( .A1(A[15]), .A2(B[15]), .ZN(n421) );
  CLKBUF_X1 U356 ( .A(B[26]), .Z(n422) );
  CLKBUF_X1 U357 ( .A(n127), .Z(n423) );
  NOR2_X1 U358 ( .A1(A[17]), .A2(B[17]), .ZN(n173) );
  NOR2_X1 U359 ( .A1(n176), .A2(n173), .ZN(n171) );
  OR2_X1 U360 ( .A1(n422), .A2(A[26]), .ZN(n424) );
  NOR2_X1 U361 ( .A1(A[15]), .A2(B[15]), .ZN(n425) );
  CLKBUF_X1 U362 ( .A(n441), .Z(n426) );
  NOR2_X1 U363 ( .A1(B[25]), .A2(A[25]), .ZN(n427) );
  NOR2_X1 U364 ( .A1(B[25]), .A2(A[25]), .ZN(n99) );
  OAI21_X1 U365 ( .B1(n427), .B2(n107), .A(n100), .ZN(n428) );
  CLKBUF_X1 U366 ( .A(n438), .Z(n429) );
  NOR2_X1 U367 ( .A1(A[19]), .A2(B[19]), .ZN(n430) );
  OR2_X1 U368 ( .A1(n61), .A2(n70), .ZN(n431) );
  NOR2_X2 U369 ( .A1(A[29]), .A2(B[29]), .ZN(n61) );
  NOR2_X1 U370 ( .A1(A[22]), .A2(B[22]), .ZN(n432) );
  NOR2_X1 U371 ( .A1(B[19]), .A2(A[19]), .ZN(n155) );
  BUF_X1 U372 ( .A(n178), .Z(n433) );
  BUF_X1 U373 ( .A(n178), .Z(n434) );
  AOI21_X2 U374 ( .B1(n247), .B2(n179), .A(n180), .ZN(n178) );
  BUF_X1 U375 ( .A(n112), .Z(n435) );
  OR2_X1 U376 ( .A1(n137), .A2(n144), .ZN(n436) );
  NOR2_X1 U377 ( .A1(n440), .A2(n126), .ZN(n437) );
  NOR2_X1 U378 ( .A1(B[27]), .A2(A[27]), .ZN(n438) );
  NOR2_X1 U379 ( .A1(B[21]), .A2(A[21]), .ZN(n439) );
  NOR2_X1 U380 ( .A1(A[23]), .A2(B[23]), .ZN(n440) );
  AOI21_X1 U381 ( .B1(n153), .B2(n172), .A(n154), .ZN(n441) );
  AOI21_X2 U382 ( .B1(n98), .B2(n77), .A(n78), .ZN(n5) );
  CLKBUF_X1 U383 ( .A(n117), .Z(n442) );
  NOR2_X1 U384 ( .A1(A[4]), .A2(B[4]), .ZN(n265) );
  NOR2_X1 U385 ( .A1(A[12]), .A2(B[12]), .ZN(n212) );
  NOR2_X1 U386 ( .A1(A[10]), .A2(B[10]), .ZN(n230) );
  NOR2_X1 U387 ( .A1(A[5]), .A2(B[5]), .ZN(n260) );
  NOR2_X1 U388 ( .A1(A[7]), .A2(B[7]), .ZN(n252) );
  NOR2_X1 U389 ( .A1(A[8]), .A2(B[8]), .ZN(n244) );
  NOR2_X1 U390 ( .A1(A[3]), .A2(B[3]), .ZN(n271) );
  NOR2_X1 U391 ( .A1(A[6]), .A2(B[6]), .ZN(n255) );
  NOR2_X1 U392 ( .A1(A[2]), .A2(B[2]), .ZN(n274) );
  NOR2_X1 U393 ( .A1(A[1]), .A2(B[1]), .ZN(n278) );
  INV_X1 U394 ( .A(n151), .ZN(n149) );
  NAND2_X1 U395 ( .A1(n149), .A2(n131), .ZN(n129) );
  INV_X1 U396 ( .A(n134), .ZN(n132) );
  INV_X1 U397 ( .A(n149), .ZN(n147) );
  BUF_X1 U398 ( .A(n178), .Z(n1) );
  INV_X1 U399 ( .A(n219), .ZN(n217) );
  BUF_X1 U400 ( .A(n178), .Z(n2) );
  OAI21_X1 U401 ( .B1(n246), .B2(n197), .A(n198), .ZN(n196) );
  AOI21_X1 U402 ( .B1(n218), .B2(n203), .A(n200), .ZN(n198) );
  NAND2_X1 U403 ( .A1(n217), .A2(n203), .ZN(n197) );
  INV_X1 U404 ( .A(n202), .ZN(n200) );
  OAI21_X1 U405 ( .B1(n246), .B2(n219), .A(n220), .ZN(n214) );
  OAI21_X1 U406 ( .B1(n246), .B2(n237), .A(n234), .ZN(n232) );
  INV_X1 U407 ( .A(n240), .ZN(n234) );
  CLKBUF_X3 U408 ( .A(n111), .Z(n4) );
  INV_X1 U409 ( .A(n436), .ZN(n131) );
  INV_X1 U410 ( .A(n6), .ZN(n75) );
  INV_X1 U411 ( .A(n95), .ZN(n93) );
  INV_X1 U412 ( .A(n247), .ZN(n246) );
  AOI21_X1 U413 ( .B1(n267), .B2(n258), .A(n259), .ZN(n257) );
  NOR2_X1 U414 ( .A1(n201), .A2(n194), .ZN(n190) );
  NOR2_X1 U415 ( .A1(n95), .A2(n86), .ZN(n84) );
  INV_X1 U416 ( .A(n428), .ZN(n96) );
  INV_X1 U417 ( .A(n220), .ZN(n218) );
  INV_X1 U418 ( .A(n136), .ZN(n134) );
  NOR2_X1 U419 ( .A1(n436), .A2(n124), .ZN(n122) );
  NAND2_X1 U420 ( .A1(n97), .A2(n77), .ZN(n6) );
  NAND2_X1 U421 ( .A1(n239), .A2(n221), .ZN(n219) );
  INV_X1 U422 ( .A(n204), .ZN(n202) );
  INV_X1 U423 ( .A(n268), .ZN(n267) );
  INV_X1 U424 ( .A(n203), .ZN(n201) );
  INV_X1 U425 ( .A(n277), .ZN(n276) );
  INV_X1 U426 ( .A(n170), .ZN(n168) );
  INV_X1 U427 ( .A(n172), .ZN(n170) );
  INV_X1 U428 ( .A(n169), .ZN(n167) );
  INV_X1 U429 ( .A(n171), .ZN(n169) );
  INV_X1 U430 ( .A(n60), .ZN(n58) );
  INV_X1 U431 ( .A(n239), .ZN(n237) );
  OAI21_X1 U432 ( .B1(n241), .B2(n245), .A(n242), .ZN(n240) );
  NOR2_X1 U433 ( .A1(n244), .A2(n241), .ZN(n239) );
  OAI21_X1 U434 ( .B1(n173), .B2(n177), .A(n174), .ZN(n172) );
  NAND2_X1 U435 ( .A1(n149), .A2(n142), .ZN(n140) );
  AOI21_X1 U436 ( .B1(n168), .B2(n160), .A(n161), .ZN(n159) );
  NAND2_X1 U437 ( .A1(n167), .A2(n160), .ZN(n158) );
  INV_X1 U438 ( .A(n163), .ZN(n161) );
  AOI21_X1 U439 ( .B1(n269), .B2(n277), .A(n270), .ZN(n268) );
  OAI21_X1 U440 ( .B1(n271), .B2(n275), .A(n272), .ZN(n270) );
  NOR2_X1 U441 ( .A1(n274), .A2(n271), .ZN(n269) );
  OAI21_X1 U442 ( .B1(n260), .B2(n266), .A(n261), .ZN(n259) );
  OAI21_X1 U443 ( .B1(n278), .B2(n281), .A(n279), .ZN(n277) );
  AOI21_X1 U444 ( .B1(n221), .B2(n240), .A(n222), .ZN(n220) );
  NOR2_X1 U445 ( .A1(n265), .A2(n260), .ZN(n258) );
  INV_X1 U446 ( .A(n107), .ZN(n105) );
  NAND2_X1 U447 ( .A1(n122), .A2(n149), .ZN(n120) );
  OAI21_X1 U448 ( .B1(n134), .B2(n124), .A(n423), .ZN(n123) );
  OAI21_X1 U449 ( .B1(n268), .B2(n248), .A(n249), .ZN(n247) );
  AOI21_X1 U450 ( .B1(n250), .B2(n259), .A(n251), .ZN(n249) );
  NAND2_X1 U451 ( .A1(n258), .A2(n250), .ZN(n248) );
  NOR2_X1 U452 ( .A1(n255), .A2(n252), .ZN(n250) );
  OAI21_X1 U453 ( .B1(n252), .B2(n256), .A(n253), .ZN(n251) );
  AOI21_X1 U454 ( .B1(n267), .B2(n309), .A(n264), .ZN(n262) );
  INV_X1 U455 ( .A(n266), .ZN(n264) );
  INV_X1 U456 ( .A(n424), .ZN(n86) );
  XOR2_X1 U457 ( .A(n257), .B(n32), .Z(SUM[6]) );
  NAND2_X1 U458 ( .A1(n307), .A2(n256), .ZN(n32) );
  AOI21_X1 U459 ( .B1(n60), .B2(n420), .A(n49), .ZN(n47) );
  INV_X1 U460 ( .A(n51), .ZN(n49) );
  OAI21_X1 U461 ( .B1(n276), .B2(n274), .A(n275), .ZN(n273) );
  OAI21_X1 U462 ( .B1(n257), .B2(n255), .A(n256), .ZN(n254) );
  OAI21_X1 U463 ( .B1(n246), .B2(n244), .A(n245), .ZN(n243) );
  OAI21_X1 U464 ( .B1(n246), .B2(n208), .A(n209), .ZN(n207) );
  AOI21_X1 U465 ( .B1(n218), .B2(n210), .A(n211), .ZN(n209) );
  NAND2_X1 U466 ( .A1(n217), .A2(n210), .ZN(n208) );
  INV_X1 U467 ( .A(n213), .ZN(n211) );
  INV_X1 U468 ( .A(n106), .ZN(n104) );
  OAI21_X1 U469 ( .B1(n246), .B2(n188), .A(n189), .ZN(n187) );
  AOI21_X1 U470 ( .B1(n190), .B2(n218), .A(n191), .ZN(n189) );
  NAND2_X1 U471 ( .A1(n190), .A2(n217), .ZN(n188) );
  OAI21_X1 U472 ( .B1(n202), .B2(n194), .A(n195), .ZN(n191) );
  OAI21_X1 U473 ( .B1(n96), .B2(n86), .A(n418), .ZN(n85) );
  INV_X1 U474 ( .A(n230), .ZN(n228) );
  INV_X1 U475 ( .A(n212), .ZN(n210) );
  INV_X1 U476 ( .A(n125), .ZN(n124) );
  INV_X1 U477 ( .A(n427), .ZN(n288) );
  INV_X1 U478 ( .A(n442), .ZN(n290) );
  INV_X1 U479 ( .A(n255), .ZN(n307) );
  INV_X1 U480 ( .A(n274), .ZN(n311) );
  INV_X1 U481 ( .A(n260), .ZN(n308) );
  INV_X1 U482 ( .A(n252), .ZN(n306) );
  INV_X1 U483 ( .A(n265), .ZN(n309) );
  INV_X1 U484 ( .A(n271), .ZN(n310) );
  NAND2_X1 U485 ( .A1(n297), .A2(n177), .ZN(n22) );
  INV_X1 U486 ( .A(n176), .ZN(n297) );
  OAI21_X1 U487 ( .B1(n246), .B2(n226), .A(n227), .ZN(n225) );
  AOI21_X1 U488 ( .B1(n240), .B2(n228), .A(n229), .ZN(n227) );
  NAND2_X1 U489 ( .A1(n239), .A2(n228), .ZN(n226) );
  INV_X1 U490 ( .A(n231), .ZN(n229) );
  NAND2_X1 U491 ( .A1(n302), .A2(n224), .ZN(n27) );
  INV_X1 U492 ( .A(n223), .ZN(n302) );
  INV_X1 U493 ( .A(n244), .ZN(n305) );
  NAND2_X1 U494 ( .A1(n210), .A2(n213), .ZN(n26) );
  NAND2_X1 U495 ( .A1(n228), .A2(n231), .ZN(n28) );
  NAND2_X1 U496 ( .A1(n284), .A2(n62), .ZN(n9) );
  NAND2_X1 U497 ( .A1(n445), .A2(n40), .ZN(n7) );
  NAND2_X1 U498 ( .A1(n288), .A2(n100), .ZN(n13) );
  NAND2_X1 U499 ( .A1(n424), .A2(n418), .ZN(n12) );
  NAND2_X1 U500 ( .A1(n286), .A2(n80), .ZN(n11) );
  NAND2_X1 U501 ( .A1(n69), .A2(n417), .ZN(n10) );
  XOR2_X1 U502 ( .A(n276), .B(n36), .Z(SUM[2]) );
  NAND2_X1 U503 ( .A1(n311), .A2(n275), .ZN(n36) );
  XNOR2_X1 U504 ( .A(n273), .B(n35), .ZN(SUM[3]) );
  NAND2_X1 U505 ( .A1(n310), .A2(n272), .ZN(n35) );
  XOR2_X1 U506 ( .A(n246), .B(n30), .Z(SUM[8]) );
  NAND2_X1 U507 ( .A1(n305), .A2(n245), .ZN(n30) );
  XNOR2_X1 U508 ( .A(n254), .B(n31), .ZN(SUM[7]) );
  NAND2_X1 U509 ( .A1(n306), .A2(n253), .ZN(n31) );
  XOR2_X1 U510 ( .A(n262), .B(n33), .Z(SUM[5]) );
  NAND2_X1 U511 ( .A1(n308), .A2(n261), .ZN(n33) );
  XNOR2_X1 U512 ( .A(n267), .B(n34), .ZN(SUM[4]) );
  NAND2_X1 U513 ( .A1(n309), .A2(n266), .ZN(n34) );
  XOR2_X1 U514 ( .A(n37), .B(n281), .Z(SUM[1]) );
  NAND2_X1 U515 ( .A1(n312), .A2(n279), .ZN(n37) );
  AND2_X1 U516 ( .A1(n444), .A2(n281), .ZN(SUM[0]) );
  NAND2_X1 U517 ( .A1(n420), .A2(n51), .ZN(n8) );
  NAND2_X1 U518 ( .A1(n300), .A2(n206), .ZN(n25) );
  INV_X1 U519 ( .A(n205), .ZN(n300) );
  NAND2_X1 U520 ( .A1(n193), .A2(n195), .ZN(n24) );
  NAND2_X1 U521 ( .A1(n304), .A2(n242), .ZN(n29) );
  NAND2_X1 U522 ( .A1(n421), .A2(n186), .ZN(n23) );
  NAND2_X1 U523 ( .A1(n296), .A2(n174), .ZN(n21) );
  INV_X1 U524 ( .A(n173), .ZN(n296) );
  INV_X1 U525 ( .A(n278), .ZN(n312) );
  INV_X1 U526 ( .A(n145), .ZN(n143) );
  INV_X1 U527 ( .A(n439), .ZN(n292) );
  INV_X1 U528 ( .A(n155), .ZN(n294) );
  INV_X1 U529 ( .A(n69), .ZN(n68) );
  OR2_X1 U530 ( .A1(A[0]), .A2(B[0]), .ZN(n444) );
  NOR2_X1 U531 ( .A1(A[13]), .A2(B[13]), .ZN(n205) );
  NOR2_X1 U532 ( .A1(A[11]), .A2(B[11]), .ZN(n223) );
  NOR2_X1 U533 ( .A1(B[21]), .A2(A[21]), .ZN(n137) );
  NOR2_X1 U534 ( .A1(B[28]), .A2(A[28]), .ZN(n70) );
  NAND2_X1 U535 ( .A1(A[8]), .A2(B[8]), .ZN(n245) );
  NOR2_X1 U536 ( .A1(B[23]), .A2(A[23]), .ZN(n117) );
  NOR2_X1 U537 ( .A1(A[14]), .A2(B[14]), .ZN(n194) );
  NAND2_X1 U538 ( .A1(A[30]), .A2(B[30]), .ZN(n51) );
  NAND2_X1 U539 ( .A1(A[4]), .A2(B[4]), .ZN(n266) );
  NAND2_X1 U540 ( .A1(A[6]), .A2(B[6]), .ZN(n256) );
  NAND2_X1 U541 ( .A1(A[2]), .A2(B[2]), .ZN(n275) );
  NAND2_X1 U542 ( .A1(A[5]), .A2(B[5]), .ZN(n261) );
  NAND2_X1 U543 ( .A1(A[7]), .A2(B[7]), .ZN(n253) );
  NAND2_X1 U544 ( .A1(A[0]), .A2(B[0]), .ZN(n281) );
  XNOR2_X1 U545 ( .A(n243), .B(n29), .ZN(SUM[9]) );
  NAND2_X1 U546 ( .A1(B[26]), .A2(A[26]), .ZN(n89) );
  NAND2_X1 U547 ( .A1(A[12]), .A2(B[12]), .ZN(n213) );
  NAND2_X1 U548 ( .A1(A[10]), .A2(B[10]), .ZN(n231) );
  NAND2_X1 U549 ( .A1(A[14]), .A2(B[14]), .ZN(n195) );
  NAND2_X1 U550 ( .A1(A[3]), .A2(B[3]), .ZN(n272) );
  NAND2_X1 U551 ( .A1(A[1]), .A2(B[1]), .ZN(n279) );
  NAND2_X1 U552 ( .A1(A[13]), .A2(B[13]), .ZN(n206) );
  NAND2_X1 U553 ( .A1(A[9]), .A2(B[9]), .ZN(n242) );
  NAND2_X1 U554 ( .A1(A[17]), .A2(B[17]), .ZN(n174) );
  NAND2_X1 U555 ( .A1(A[31]), .A2(B[31]), .ZN(n40) );
  NAND2_X1 U556 ( .A1(A[29]), .A2(B[29]), .ZN(n62) );
  NAND2_X1 U557 ( .A1(n104), .A2(n107), .ZN(n14) );
  XNOR2_X1 U558 ( .A(n128), .B(n16), .ZN(SUM[22]) );
  NAND2_X1 U559 ( .A1(n125), .A2(n423), .ZN(n16) );
  XNOR2_X1 U560 ( .A(n139), .B(n17), .ZN(SUM[21]) );
  NAND2_X1 U561 ( .A1(n292), .A2(n138), .ZN(n17) );
  XNOR2_X1 U562 ( .A(n146), .B(n18), .ZN(SUM[20]) );
  NAND2_X1 U563 ( .A1(n142), .A2(n145), .ZN(n18) );
  NAND2_X1 U564 ( .A1(n290), .A2(n118), .ZN(n15) );
  XNOR2_X1 U565 ( .A(n157), .B(n19), .ZN(SUM[19]) );
  NAND2_X1 U566 ( .A1(n294), .A2(n156), .ZN(n19) );
  XNOR2_X1 U567 ( .A(n164), .B(n20), .ZN(SUM[18]) );
  XNOR2_X1 U568 ( .A(n207), .B(n25), .ZN(SUM[13]) );
  XNOR2_X1 U569 ( .A(n196), .B(n24), .ZN(SUM[14]) );
  XNOR2_X1 U570 ( .A(n214), .B(n26), .ZN(SUM[12]) );
  XNOR2_X1 U571 ( .A(n175), .B(n21), .ZN(SUM[17]) );
  XNOR2_X1 U572 ( .A(n225), .B(n27), .ZN(SUM[11]) );
  XNOR2_X1 U573 ( .A(n232), .B(n28), .ZN(SUM[10]) );
  OR2_X1 U574 ( .A1(A[31]), .A2(B[31]), .ZN(n445) );
  NOR2_X1 U575 ( .A1(n438), .A2(n88), .ZN(n77) );
  NOR2_X1 U576 ( .A1(B[24]), .A2(A[24]), .ZN(n106) );
  NAND2_X1 U577 ( .A1(B[24]), .A2(A[24]), .ZN(n107) );
  XNOR2_X1 U578 ( .A(n187), .B(n23), .ZN(SUM[15]) );
  AOI21_X1 U579 ( .B1(n122), .B2(n150), .A(n123), .ZN(n121) );
  AOI21_X1 U580 ( .B1(n150), .B2(n131), .A(n132), .ZN(n130) );
  AOI21_X1 U581 ( .B1(n150), .B2(n142), .A(n143), .ZN(n141) );
  INV_X1 U582 ( .A(n150), .ZN(n148) );
  XNOR2_X1 U583 ( .A(n108), .B(n14), .ZN(SUM[24]) );
  NAND2_X1 U584 ( .A1(n160), .A2(n163), .ZN(n20) );
  INV_X1 U585 ( .A(n426), .ZN(n150) );
  NAND2_X1 U586 ( .A1(B[22]), .A2(A[22]), .ZN(n127) );
  NOR2_X1 U587 ( .A1(A[22]), .A2(B[22]), .ZN(n126) );
  XNOR2_X1 U588 ( .A(n81), .B(n11), .ZN(SUM[27]) );
  XNOR2_X1 U589 ( .A(n72), .B(n10), .ZN(SUM[28]) );
  NOR2_X1 U590 ( .A1(A[16]), .A2(B[16]), .ZN(n176) );
  NAND2_X1 U591 ( .A1(A[16]), .A2(B[16]), .ZN(n177) );
  INV_X1 U592 ( .A(n144), .ZN(n142) );
  NAND2_X1 U593 ( .A1(A[20]), .A2(B[20]), .ZN(n145) );
  INV_X1 U594 ( .A(n61), .ZN(n284) );
  NOR2_X1 U595 ( .A1(n70), .A2(n61), .ZN(n59) );
  NAND2_X1 U596 ( .A1(A[18]), .A2(B[18]), .ZN(n163) );
  XNOR2_X1 U597 ( .A(n90), .B(n12), .ZN(SUM[26]) );
  INV_X1 U598 ( .A(n4), .ZN(n109) );
  INV_X1 U599 ( .A(n435), .ZN(n110) );
  XNOR2_X1 U600 ( .A(n119), .B(n15), .ZN(SUM[23]) );
  INV_X1 U601 ( .A(n432), .ZN(n125) );
  NOR2_X1 U602 ( .A1(n106), .A2(n99), .ZN(n97) );
  INV_X1 U603 ( .A(n97), .ZN(n95) );
  XNOR2_X1 U604 ( .A(n63), .B(n9), .ZN(SUM[29]) );
  INV_X1 U605 ( .A(n429), .ZN(n286) );
  NOR2_X1 U606 ( .A1(n6), .A2(n431), .ZN(n55) );
  NOR2_X1 U607 ( .A1(n6), .A2(n68), .ZN(n66) );
  OAI21_X1 U608 ( .B1(n433), .B2(n102), .A(n103), .ZN(n101) );
  OAI21_X1 U609 ( .B1(n434), .B2(n42), .A(n43), .ZN(n41) );
  OAI21_X1 U610 ( .B1(n2), .B2(n109), .A(n110), .ZN(n108) );
  NAND2_X1 U611 ( .A1(A[15]), .A2(B[15]), .ZN(n186) );
  NOR2_X1 U612 ( .A1(A[15]), .A2(B[15]), .ZN(n185) );
  NOR2_X1 U613 ( .A1(n144), .A2(n137), .ZN(n135) );
  NOR2_X1 U614 ( .A1(A[20]), .A2(B[20]), .ZN(n144) );
  INV_X1 U615 ( .A(n241), .ZN(n304) );
  NOR2_X1 U616 ( .A1(A[9]), .A2(B[9]), .ZN(n241) );
  INV_X1 U617 ( .A(n70), .ZN(n69) );
  NAND2_X1 U618 ( .A1(B[28]), .A2(A[28]), .ZN(n71) );
  INV_X1 U619 ( .A(n162), .ZN(n160) );
  NOR2_X1 U620 ( .A1(A[18]), .A2(B[18]), .ZN(n162) );
  NOR2_X1 U621 ( .A1(n230), .A2(n223), .ZN(n221) );
  OAI21_X1 U622 ( .B1(n223), .B2(n231), .A(n224), .ZN(n222) );
  NAND2_X1 U623 ( .A1(A[11]), .A2(B[11]), .ZN(n224) );
  OAI21_X1 U624 ( .B1(n61), .B2(n71), .A(n62), .ZN(n60) );
  NOR2_X1 U625 ( .A1(B[26]), .A2(A[26]), .ZN(n88) );
  OAI21_X1 U626 ( .B1(n220), .B2(n181), .A(n182), .ZN(n180) );
  NOR2_X1 U627 ( .A1(n219), .A2(n181), .ZN(n179) );
  OAI21_X1 U628 ( .B1(n205), .B2(n213), .A(n206), .ZN(n204) );
  NAND2_X1 U629 ( .A1(n203), .A2(n183), .ZN(n181) );
  AOI21_X1 U630 ( .B1(n183), .B2(n204), .A(n184), .ZN(n182) );
  NOR2_X1 U631 ( .A1(n194), .A2(n425), .ZN(n183) );
  INV_X1 U632 ( .A(n194), .ZN(n193) );
  NAND2_X1 U633 ( .A1(n171), .A2(n153), .ZN(n151) );
  XNOR2_X1 U634 ( .A(n52), .B(n8), .ZN(SUM[30]) );
  NAND2_X1 U635 ( .A1(n59), .A2(n420), .ZN(n46) );
  XNOR2_X1 U636 ( .A(n41), .B(n7), .ZN(SUM[31]) );
  OAI21_X1 U637 ( .B1(n2), .B2(n91), .A(n92), .ZN(n90) );
  INV_X1 U638 ( .A(n5), .ZN(n76) );
  XNOR2_X1 U639 ( .A(n101), .B(n13), .ZN(SUM[25]) );
  OAI21_X1 U640 ( .B1(n434), .B2(n82), .A(n83), .ZN(n81) );
  NAND2_X1 U641 ( .A1(A[25]), .A2(B[25]), .ZN(n100) );
  XOR2_X1 U642 ( .A(n2), .B(n22), .Z(SUM[16]) );
  OAI21_X1 U643 ( .B1(n433), .B2(n120), .A(n121), .ZN(n119) );
  OAI21_X1 U644 ( .B1(n434), .B2(n129), .A(n130), .ZN(n128) );
  OAI21_X1 U645 ( .B1(n2), .B2(n140), .A(n141), .ZN(n139) );
  OAI21_X1 U646 ( .B1(n1), .B2(n147), .A(n148), .ZN(n146) );
  OAI21_X1 U647 ( .B1(n1), .B2(n158), .A(n159), .ZN(n157) );
  OAI21_X1 U648 ( .B1(n1), .B2(n169), .A(n170), .ZN(n164) );
  OAI21_X1 U649 ( .B1(n1), .B2(n176), .A(n177), .ZN(n175) );
  NOR2_X1 U650 ( .A1(n212), .A2(n205), .ZN(n203) );
  OAI21_X1 U651 ( .B1(n433), .B2(n73), .A(n74), .ZN(n72) );
  NOR2_X1 U652 ( .A1(n151), .A2(n113), .ZN(n111) );
  OAI21_X1 U653 ( .B1(n441), .B2(n113), .A(n114), .ZN(n112) );
  OAI21_X1 U654 ( .B1(n53), .B2(n434), .A(n54), .ZN(n52) );
  NOR2_X1 U655 ( .A1(n162), .A2(n155), .ZN(n153) );
  OAI21_X1 U656 ( .B1(n430), .B2(n163), .A(n156), .ZN(n154) );
  NAND2_X1 U657 ( .A1(B[19]), .A2(A[19]), .ZN(n156) );
  OAI21_X1 U658 ( .B1(n64), .B2(n433), .A(n65), .ZN(n63) );
  NAND2_X1 U659 ( .A1(n419), .A2(n4), .ZN(n42) );
  NAND2_X1 U660 ( .A1(n55), .A2(n4), .ZN(n53) );
  NAND2_X1 U661 ( .A1(n66), .A2(n4), .ZN(n64) );
  NAND2_X1 U662 ( .A1(n4), .A2(n75), .ZN(n73) );
  NAND2_X1 U663 ( .A1(n4), .A2(n84), .ZN(n82) );
  NAND2_X1 U664 ( .A1(n4), .A2(n93), .ZN(n91) );
  NAND2_X1 U665 ( .A1(n4), .A2(n104), .ZN(n102) );
  NAND2_X1 U666 ( .A1(n135), .A2(n437), .ZN(n113) );
  NAND2_X1 U667 ( .A1(B[21]), .A2(A[21]), .ZN(n138) );
  AOI21_X1 U668 ( .B1(n416), .B2(n93), .A(n428), .ZN(n92) );
  AOI21_X1 U669 ( .B1(n416), .B2(n104), .A(n105), .ZN(n103) );
  AOI21_X1 U670 ( .B1(n416), .B2(n75), .A(n76), .ZN(n74) );
  AOI21_X1 U671 ( .B1(n435), .B2(n84), .A(n85), .ZN(n83) );
  AOI21_X1 U672 ( .B1(n435), .B2(n419), .A(n45), .ZN(n43) );
  AOI21_X1 U673 ( .B1(n3), .B2(n55), .A(n56), .ZN(n54) );
  AOI21_X1 U674 ( .B1(n3), .B2(n66), .A(n67), .ZN(n65) );
  OAI21_X1 U675 ( .B1(n99), .B2(n107), .A(n100), .ZN(n98) );
  OAI21_X1 U676 ( .B1(n185), .B2(n195), .A(n186), .ZN(n184) );
  AOI21_X1 U677 ( .B1(n136), .B2(n115), .A(n116), .ZN(n114) );
  NOR2_X1 U678 ( .A1(n432), .A2(n440), .ZN(n115) );
  OAI21_X1 U679 ( .B1(n5), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U680 ( .B1(n5), .B2(n431), .A(n58), .ZN(n56) );
  OAI21_X1 U681 ( .B1(n5), .B2(n68), .A(n417), .ZN(n67) );
  OAI21_X1 U682 ( .B1(n79), .B2(n89), .A(n80), .ZN(n78) );
  NAND2_X1 U683 ( .A1(B[27]), .A2(A[27]), .ZN(n80) );
  NOR2_X1 U684 ( .A1(B[27]), .A2(A[27]), .ZN(n79) );
  OAI21_X1 U685 ( .B1(n117), .B2(n127), .A(n118), .ZN(n116) );
  NAND2_X1 U686 ( .A1(B[23]), .A2(A[23]), .ZN(n118) );
  OAI21_X1 U687 ( .B1(n439), .B2(n145), .A(n138), .ZN(n136) );
endmodule


module datapath_DW01_add_15 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n40, n41, n42, n43, n44, n45, n46,
         n47, n49, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n125, n126, n127, n128,
         n129, n130, n131, n132, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n166, n167, n169, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n193, n194, n195, n196, n197, n198, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n234, n237, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n281, n284, n286, n287, n288, n290, n292,
         n294, n296, n297, n298, n300, n302, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n444, n445;

  BUF_X1 U349 ( .A(n112), .Z(n416) );
  AOI21_X2 U350 ( .B1(n247), .B2(n179), .A(n180), .ZN(n178) );
  BUF_X1 U351 ( .A(n424), .Z(n439) );
  BUF_X1 U352 ( .A(n152), .Z(n432) );
  OR2_X1 U353 ( .A1(A[30]), .A2(B[30]), .ZN(n417) );
  CLKBUF_X1 U354 ( .A(n172), .Z(n430) );
  INV_X1 U355 ( .A(n143), .ZN(n418) );
  NAND2_X1 U356 ( .A1(n98), .A2(n77), .ZN(n419) );
  INV_X1 U357 ( .A(n78), .ZN(n420) );
  AND2_X2 U358 ( .A1(n419), .A2(n420), .ZN(n5) );
  NOR2_X1 U359 ( .A1(n79), .A2(n88), .ZN(n77) );
  NOR2_X1 U360 ( .A1(A[15]), .A2(B[15]), .ZN(n421) );
  NOR2_X1 U361 ( .A1(A[15]), .A2(B[15]), .ZN(n185) );
  OR2_X1 U362 ( .A1(n439), .A2(n144), .ZN(n422) );
  NOR2_X1 U363 ( .A1(B[27]), .A2(A[27]), .ZN(n423) );
  NOR2_X1 U364 ( .A1(A[21]), .A2(B[21]), .ZN(n424) );
  CLKBUF_X1 U365 ( .A(n61), .Z(n425) );
  CLKBUF_X1 U366 ( .A(n88), .Z(n426) );
  INV_X1 U367 ( .A(n297), .ZN(n427) );
  NAND2_X1 U368 ( .A1(A[24]), .A2(B[24]), .ZN(n107) );
  NOR2_X1 U369 ( .A1(B[25]), .A2(A[25]), .ZN(n428) );
  NOR2_X1 U370 ( .A1(n126), .A2(n117), .ZN(n429) );
  CLKBUF_X1 U371 ( .A(n136), .Z(n431) );
  BUF_X1 U372 ( .A(n178), .Z(n433) );
  BUF_X1 U373 ( .A(n178), .Z(n434) );
  NOR2_X1 U374 ( .A1(B[23]), .A2(A[23]), .ZN(n435) );
  NOR2_X1 U375 ( .A1(B[25]), .A2(A[25]), .ZN(n99) );
  CLKBUF_X1 U376 ( .A(n423), .Z(n436) );
  CLKBUF_X1 U377 ( .A(n126), .Z(n437) );
  CLKBUF_X1 U378 ( .A(n144), .Z(n438) );
  CLKBUF_X1 U379 ( .A(n435), .Z(n440) );
  BUF_X1 U380 ( .A(n112), .Z(n441) );
  BUF_X1 U381 ( .A(n111), .Z(n442) );
  NOR2_X1 U382 ( .A1(A[12]), .A2(B[12]), .ZN(n212) );
  NOR2_X1 U383 ( .A1(A[4]), .A2(B[4]), .ZN(n265) );
  NOR2_X1 U384 ( .A1(A[3]), .A2(B[3]), .ZN(n271) );
  NOR2_X1 U385 ( .A1(A[5]), .A2(B[5]), .ZN(n260) );
  NOR2_X1 U386 ( .A1(A[9]), .A2(B[9]), .ZN(n241) );
  NOR2_X1 U387 ( .A1(A[7]), .A2(B[7]), .ZN(n252) );
  NOR2_X1 U388 ( .A1(A[8]), .A2(B[8]), .ZN(n244) );
  NOR2_X1 U389 ( .A1(A[2]), .A2(B[2]), .ZN(n274) );
  NOR2_X1 U390 ( .A1(A[6]), .A2(B[6]), .ZN(n255) );
  NOR2_X1 U391 ( .A1(A[1]), .A2(B[1]), .ZN(n278) );
  AOI21_X1 U392 ( .B1(n150), .B2(n131), .A(n132), .ZN(n130) );
  INV_X1 U393 ( .A(n422), .ZN(n131) );
  BUF_X1 U394 ( .A(n178), .Z(n2) );
  BUF_X1 U395 ( .A(n178), .Z(n1) );
  INV_X1 U396 ( .A(n219), .ZN(n217) );
  BUF_X1 U397 ( .A(n111), .Z(n4) );
  OAI21_X1 U398 ( .B1(n246), .B2(n197), .A(n198), .ZN(n196) );
  NAND2_X1 U399 ( .A1(n217), .A2(n203), .ZN(n197) );
  AOI21_X1 U400 ( .B1(n218), .B2(n203), .A(n204), .ZN(n198) );
  OAI21_X1 U401 ( .B1(n246), .B2(n219), .A(n220), .ZN(n214) );
  OAI21_X1 U402 ( .B1(n246), .B2(n237), .A(n234), .ZN(n232) );
  INV_X1 U403 ( .A(n240), .ZN(n234) );
  OAI21_X1 U404 ( .B1(n1), .B2(n147), .A(n432), .ZN(n146) );
  INV_X1 U405 ( .A(n149), .ZN(n147) );
  OAI21_X1 U406 ( .B1(n1), .B2(n169), .A(n166), .ZN(n164) );
  INV_X1 U407 ( .A(n430), .ZN(n166) );
  INV_X1 U408 ( .A(n151), .ZN(n149) );
  INV_X1 U409 ( .A(n134), .ZN(n132) );
  INV_X1 U410 ( .A(n96), .ZN(n94) );
  INV_X1 U411 ( .A(n220), .ZN(n218) );
  INV_X1 U412 ( .A(n247), .ZN(n246) );
  AOI21_X1 U413 ( .B1(n122), .B2(n150), .A(n123), .ZN(n121) );
  NOR2_X1 U414 ( .A1(n422), .A2(n437), .ZN(n122) );
  INV_X1 U415 ( .A(n432), .ZN(n150) );
  AOI21_X1 U416 ( .B1(n267), .B2(n258), .A(n259), .ZN(n257) );
  NOR2_X1 U417 ( .A1(n201), .A2(n194), .ZN(n190) );
  INV_X1 U418 ( .A(n95), .ZN(n93) );
  NOR2_X1 U419 ( .A1(n95), .A2(n426), .ZN(n84) );
  INV_X1 U420 ( .A(n6), .ZN(n75) );
  INV_X1 U421 ( .A(n441), .ZN(n110) );
  INV_X1 U422 ( .A(n60), .ZN(n58) );
  INV_X1 U423 ( .A(n97), .ZN(n95) );
  INV_X1 U424 ( .A(n203), .ZN(n201) );
  INV_X1 U425 ( .A(n431), .ZN(n134) );
  INV_X1 U426 ( .A(n204), .ZN(n202) );
  INV_X1 U427 ( .A(n268), .ZN(n267) );
  NAND2_X1 U428 ( .A1(n239), .A2(n221), .ZN(n219) );
  INV_X1 U429 ( .A(n277), .ZN(n276) );
  INV_X1 U430 ( .A(n169), .ZN(n167) );
  INV_X1 U431 ( .A(n239), .ZN(n237) );
  INV_X1 U432 ( .A(n59), .ZN(n57) );
  AOI21_X1 U433 ( .B1(n269), .B2(n277), .A(n270), .ZN(n268) );
  OAI21_X1 U434 ( .B1(n271), .B2(n275), .A(n272), .ZN(n270) );
  NOR2_X1 U435 ( .A1(n274), .A2(n271), .ZN(n269) );
  AOI21_X1 U436 ( .B1(n221), .B2(n240), .A(n222), .ZN(n220) );
  OAI21_X1 U437 ( .B1(n260), .B2(n266), .A(n261), .ZN(n259) );
  OAI21_X1 U438 ( .B1(n278), .B2(n281), .A(n279), .ZN(n277) );
  NOR2_X1 U439 ( .A1(n255), .A2(n252), .ZN(n250) );
  NOR2_X1 U440 ( .A1(n244), .A2(n241), .ZN(n239) );
  NOR2_X1 U441 ( .A1(n265), .A2(n260), .ZN(n258) );
  INV_X1 U442 ( .A(n106), .ZN(n104) );
  OAI21_X1 U443 ( .B1(n241), .B2(n245), .A(n242), .ZN(n240) );
  NOR2_X1 U444 ( .A1(n137), .A2(n144), .ZN(n135) );
  OAI21_X1 U445 ( .B1(n268), .B2(n248), .A(n249), .ZN(n247) );
  AOI21_X1 U446 ( .B1(n250), .B2(n259), .A(n251), .ZN(n249) );
  NAND2_X1 U447 ( .A1(n258), .A2(n250), .ZN(n248) );
  OAI21_X1 U448 ( .B1(n252), .B2(n256), .A(n253), .ZN(n251) );
  INV_X1 U449 ( .A(n51), .ZN(n49) );
  AOI21_X1 U450 ( .B1(n267), .B2(n309), .A(n264), .ZN(n262) );
  INV_X1 U451 ( .A(n266), .ZN(n264) );
  INV_X1 U452 ( .A(n230), .ZN(n228) );
  BUF_X1 U453 ( .A(n112), .Z(n3) );
  OAI21_X1 U454 ( .B1(n134), .B2(n437), .A(n127), .ZN(n123) );
  OAI21_X1 U455 ( .B1(n246), .B2(n244), .A(n245), .ZN(n243) );
  OAI21_X1 U456 ( .B1(n257), .B2(n255), .A(n256), .ZN(n254) );
  OAI21_X1 U457 ( .B1(n276), .B2(n274), .A(n275), .ZN(n273) );
  OAI21_X1 U458 ( .B1(n246), .B2(n188), .A(n189), .ZN(n187) );
  AOI21_X1 U459 ( .B1(n190), .B2(n218), .A(n191), .ZN(n189) );
  NAND2_X1 U460 ( .A1(n190), .A2(n217), .ZN(n188) );
  OAI21_X1 U461 ( .B1(n202), .B2(n194), .A(n195), .ZN(n191) );
  OAI21_X1 U462 ( .B1(n246), .B2(n208), .A(n209), .ZN(n207) );
  AOI21_X1 U463 ( .B1(n218), .B2(n210), .A(n211), .ZN(n209) );
  NAND2_X1 U464 ( .A1(n217), .A2(n210), .ZN(n208) );
  INV_X1 U465 ( .A(n213), .ZN(n211) );
  OAI21_X1 U466 ( .B1(n246), .B2(n226), .A(n227), .ZN(n225) );
  AOI21_X1 U467 ( .B1(n240), .B2(n228), .A(n229), .ZN(n227) );
  NAND2_X1 U468 ( .A1(n239), .A2(n228), .ZN(n226) );
  INV_X1 U469 ( .A(n231), .ZN(n229) );
  OAI21_X1 U470 ( .B1(n1), .B2(n158), .A(n159), .ZN(n157) );
  NAND2_X1 U471 ( .A1(n167), .A2(n160), .ZN(n158) );
  AOI21_X1 U472 ( .B1(n430), .B2(n160), .A(n161), .ZN(n159) );
  INV_X1 U473 ( .A(n162), .ZN(n160) );
  INV_X1 U474 ( .A(n212), .ZN(n210) );
  INV_X1 U475 ( .A(n425), .ZN(n284) );
  INV_X1 U476 ( .A(n176), .ZN(n297) );
  INV_X1 U477 ( .A(n426), .ZN(n287) );
  INV_X1 U478 ( .A(n436), .ZN(n286) );
  INV_X1 U479 ( .A(n194), .ZN(n193) );
  INV_X1 U480 ( .A(n440), .ZN(n290) );
  INV_X1 U481 ( .A(n428), .ZN(n288) );
  INV_X1 U482 ( .A(n173), .ZN(n296) );
  INV_X1 U483 ( .A(n244), .ZN(n305) );
  INV_X1 U484 ( .A(n255), .ZN(n307) );
  INV_X1 U485 ( .A(n274), .ZN(n311) );
  INV_X1 U486 ( .A(n252), .ZN(n306) );
  INV_X1 U487 ( .A(n241), .ZN(n304) );
  INV_X1 U488 ( .A(n260), .ZN(n308) );
  INV_X1 U489 ( .A(n271), .ZN(n310) );
  INV_X1 U490 ( .A(n265), .ZN(n309) );
  INV_X1 U491 ( .A(n163), .ZN(n161) );
  INV_X1 U492 ( .A(n278), .ZN(n312) );
  INV_X1 U493 ( .A(n155), .ZN(n294) );
  INV_X1 U494 ( .A(n205), .ZN(n300) );
  INV_X1 U495 ( .A(n107), .ZN(n105) );
  INV_X1 U496 ( .A(n69), .ZN(n68) );
  INV_X1 U497 ( .A(n70), .ZN(n69) );
  NOR2_X1 U498 ( .A1(B[18]), .A2(A[18]), .ZN(n162) );
  NOR2_X1 U499 ( .A1(B[19]), .A2(A[19]), .ZN(n155) );
  NOR2_X1 U500 ( .A1(A[13]), .A2(B[13]), .ZN(n205) );
  NOR2_X1 U501 ( .A1(A[21]), .A2(B[21]), .ZN(n137) );
  NOR2_X1 U502 ( .A1(B[22]), .A2(A[22]), .ZN(n126) );
  NOR2_X1 U503 ( .A1(B[17]), .A2(A[17]), .ZN(n173) );
  NOR2_X1 U504 ( .A1(B[23]), .A2(A[23]), .ZN(n117) );
  NAND2_X1 U505 ( .A1(B[22]), .A2(A[22]), .ZN(n127) );
  NAND2_X1 U506 ( .A1(B[18]), .A2(A[18]), .ZN(n163) );
  NOR2_X1 U507 ( .A1(A[14]), .A2(B[14]), .ZN(n194) );
  NOR2_X1 U508 ( .A1(A[10]), .A2(B[10]), .ZN(n230) );
  NOR2_X1 U509 ( .A1(A[28]), .A2(B[28]), .ZN(n70) );
  NOR2_X1 U510 ( .A1(A[11]), .A2(B[11]), .ZN(n223) );
  AND2_X1 U511 ( .A1(n445), .A2(n281), .ZN(SUM[0]) );
  NAND2_X1 U512 ( .A1(A[6]), .A2(B[6]), .ZN(n256) );
  NAND2_X1 U513 ( .A1(A[8]), .A2(B[8]), .ZN(n245) );
  XOR2_X1 U514 ( .A(n2), .B(n22), .Z(SUM[16]) );
  NAND2_X1 U515 ( .A1(n297), .A2(n177), .ZN(n22) );
  NAND2_X1 U516 ( .A1(A[12]), .A2(B[12]), .ZN(n213) );
  NAND2_X1 U517 ( .A1(A[4]), .A2(B[4]), .ZN(n266) );
  NAND2_X1 U518 ( .A1(A[2]), .A2(B[2]), .ZN(n275) );
  XNOR2_X1 U519 ( .A(n119), .B(n15), .ZN(SUM[23]) );
  NAND2_X1 U520 ( .A1(n290), .A2(n118), .ZN(n15) );
  XNOR2_X1 U521 ( .A(n146), .B(n18), .ZN(SUM[20]) );
  XNOR2_X1 U522 ( .A(n128), .B(n16), .ZN(SUM[22]) );
  NAND2_X1 U523 ( .A1(n125), .A2(n127), .ZN(n16) );
  NAND2_X1 U524 ( .A1(n69), .A2(n71), .ZN(n10) );
  NAND2_X1 U525 ( .A1(n284), .A2(n62), .ZN(n9) );
  NAND2_X1 U526 ( .A1(n417), .A2(n51), .ZN(n8) );
  NAND2_X1 U527 ( .A1(n444), .A2(n40), .ZN(n7) );
  NAND2_X1 U528 ( .A1(n288), .A2(n100), .ZN(n13) );
  NAND2_X1 U529 ( .A1(n287), .A2(n89), .ZN(n12) );
  NAND2_X1 U530 ( .A1(n286), .A2(n80), .ZN(n11) );
  XOR2_X1 U531 ( .A(n37), .B(n281), .Z(SUM[1]) );
  NAND2_X1 U532 ( .A1(n312), .A2(n279), .ZN(n37) );
  XNOR2_X1 U533 ( .A(n273), .B(n35), .ZN(SUM[3]) );
  NAND2_X1 U534 ( .A1(n310), .A2(n272), .ZN(n35) );
  XNOR2_X1 U535 ( .A(n267), .B(n34), .ZN(SUM[4]) );
  NAND2_X1 U536 ( .A1(n309), .A2(n266), .ZN(n34) );
  XOR2_X1 U537 ( .A(n262), .B(n33), .Z(SUM[5]) );
  NAND2_X1 U538 ( .A1(n308), .A2(n261), .ZN(n33) );
  NAND2_X1 U539 ( .A1(n104), .A2(n107), .ZN(n14) );
  XNOR2_X1 U540 ( .A(n139), .B(n17), .ZN(SUM[21]) );
  NAND2_X1 U541 ( .A1(n292), .A2(n138), .ZN(n17) );
  XNOR2_X1 U542 ( .A(n175), .B(n21), .ZN(SUM[17]) );
  NAND2_X1 U543 ( .A1(n296), .A2(n174), .ZN(n21) );
  XNOR2_X1 U544 ( .A(n187), .B(n23), .ZN(SUM[15]) );
  NAND2_X1 U545 ( .A1(n298), .A2(n186), .ZN(n23) );
  XNOR2_X1 U546 ( .A(n196), .B(n24), .ZN(SUM[14]) );
  NAND2_X1 U547 ( .A1(n193), .A2(n195), .ZN(n24) );
  XNOR2_X1 U548 ( .A(n207), .B(n25), .ZN(SUM[13]) );
  NAND2_X1 U549 ( .A1(n300), .A2(n206), .ZN(n25) );
  XNOR2_X1 U550 ( .A(n214), .B(n26), .ZN(SUM[12]) );
  NAND2_X1 U551 ( .A1(n210), .A2(n213), .ZN(n26) );
  XNOR2_X1 U552 ( .A(n243), .B(n29), .ZN(SUM[9]) );
  NAND2_X1 U553 ( .A1(n304), .A2(n242), .ZN(n29) );
  XNOR2_X1 U554 ( .A(n232), .B(n28), .ZN(SUM[10]) );
  NAND2_X1 U555 ( .A1(n228), .A2(n231), .ZN(n28) );
  XNOR2_X1 U556 ( .A(n225), .B(n27), .ZN(SUM[11]) );
  NAND2_X1 U557 ( .A1(n302), .A2(n224), .ZN(n27) );
  XOR2_X1 U558 ( .A(n246), .B(n30), .Z(SUM[8]) );
  NAND2_X1 U559 ( .A1(n305), .A2(n245), .ZN(n30) );
  XOR2_X1 U560 ( .A(n257), .B(n32), .Z(SUM[6]) );
  NAND2_X1 U561 ( .A1(n307), .A2(n256), .ZN(n32) );
  XNOR2_X1 U562 ( .A(n254), .B(n31), .ZN(SUM[7]) );
  NAND2_X1 U563 ( .A1(n306), .A2(n253), .ZN(n31) );
  NAND2_X1 U564 ( .A1(A[0]), .A2(B[0]), .ZN(n281) );
  NAND2_X1 U565 ( .A1(A[9]), .A2(B[9]), .ZN(n242) );
  NAND2_X1 U566 ( .A1(A[7]), .A2(B[7]), .ZN(n253) );
  NAND2_X1 U567 ( .A1(A[10]), .A2(B[10]), .ZN(n231) );
  NAND2_X1 U568 ( .A1(A[14]), .A2(B[14]), .ZN(n195) );
  XNOR2_X1 U569 ( .A(n157), .B(n19), .ZN(SUM[19]) );
  NAND2_X1 U570 ( .A1(n294), .A2(n156), .ZN(n19) );
  XNOR2_X1 U571 ( .A(n164), .B(n20), .ZN(SUM[18]) );
  NAND2_X1 U572 ( .A1(n160), .A2(n163), .ZN(n20) );
  NAND2_X1 U573 ( .A1(A[30]), .A2(B[30]), .ZN(n51) );
  NAND2_X1 U574 ( .A1(A[5]), .A2(B[5]), .ZN(n261) );
  NAND2_X1 U575 ( .A1(A[1]), .A2(B[1]), .ZN(n279) );
  NAND2_X1 U576 ( .A1(A[3]), .A2(B[3]), .ZN(n272) );
  NAND2_X1 U577 ( .A1(A[19]), .A2(B[19]), .ZN(n156) );
  NAND2_X1 U578 ( .A1(A[29]), .A2(B[29]), .ZN(n62) );
  NAND2_X1 U579 ( .A1(A[31]), .A2(B[31]), .ZN(n40) );
  NAND2_X1 U580 ( .A1(A[15]), .A2(B[15]), .ZN(n186) );
  NAND2_X1 U581 ( .A1(A[11]), .A2(B[11]), .ZN(n224) );
  XOR2_X1 U582 ( .A(n276), .B(n36), .Z(SUM[2]) );
  NAND2_X1 U583 ( .A1(n311), .A2(n275), .ZN(n36) );
  OR2_X1 U584 ( .A1(A[31]), .A2(B[31]), .ZN(n444) );
  OR2_X1 U585 ( .A1(A[0]), .A2(B[0]), .ZN(n445) );
  XNOR2_X1 U586 ( .A(n81), .B(n11), .ZN(SUM[27]) );
  NAND2_X1 U587 ( .A1(n142), .A2(n418), .ZN(n18) );
  INV_X1 U588 ( .A(n145), .ZN(n143) );
  INV_X1 U589 ( .A(n223), .ZN(n302) );
  OAI21_X1 U590 ( .B1(n223), .B2(n231), .A(n224), .ZN(n222) );
  NOR2_X1 U591 ( .A1(n230), .A2(n223), .ZN(n221) );
  NAND2_X1 U592 ( .A1(B[20]), .A2(A[20]), .ZN(n145) );
  XNOR2_X1 U593 ( .A(n90), .B(n12), .ZN(SUM[26]) );
  NOR2_X1 U594 ( .A1(A[29]), .A2(B[29]), .ZN(n61) );
  XNOR2_X1 U595 ( .A(n101), .B(n13), .ZN(SUM[25]) );
  AOI21_X1 U596 ( .B1(n153), .B2(n172), .A(n154), .ZN(n152) );
  INV_X1 U597 ( .A(n98), .ZN(n96) );
  OAI21_X1 U598 ( .B1(n96), .B2(n426), .A(n89), .ZN(n85) );
  OAI21_X1 U599 ( .B1(n173), .B2(n177), .A(n174), .ZN(n172) );
  NAND2_X1 U600 ( .A1(A[13]), .A2(B[13]), .ZN(n206) );
  OAI21_X1 U601 ( .B1(n2), .B2(n140), .A(n141), .ZN(n139) );
  XNOR2_X1 U602 ( .A(n72), .B(n10), .ZN(SUM[28]) );
  XNOR2_X1 U603 ( .A(n108), .B(n14), .ZN(SUM[24]) );
  NOR2_X1 U604 ( .A1(A[16]), .A2(B[16]), .ZN(n176) );
  NAND2_X1 U605 ( .A1(A[16]), .A2(B[16]), .ZN(n177) );
  NOR2_X1 U606 ( .A1(A[24]), .A2(B[24]), .ZN(n106) );
  XNOR2_X1 U607 ( .A(n52), .B(n8), .ZN(SUM[30]) );
  NOR2_X1 U608 ( .A1(n106), .A2(n428), .ZN(n97) );
  NAND2_X1 U609 ( .A1(B[17]), .A2(A[17]), .ZN(n174) );
  XNOR2_X1 U610 ( .A(n63), .B(n9), .ZN(SUM[29]) );
  NAND2_X1 U611 ( .A1(A[21]), .A2(B[21]), .ZN(n138) );
  OAI21_X1 U612 ( .B1(n1), .B2(n129), .A(n130), .ZN(n128) );
  NAND2_X1 U613 ( .A1(n122), .A2(n149), .ZN(n120) );
  NAND2_X1 U614 ( .A1(n149), .A2(n142), .ZN(n140) );
  NAND2_X1 U615 ( .A1(n149), .A2(n131), .ZN(n129) );
  NOR2_X1 U616 ( .A1(n219), .A2(n181), .ZN(n179) );
  INV_X1 U617 ( .A(n5), .ZN(n76) );
  INV_X1 U618 ( .A(n439), .ZN(n292) );
  AOI21_X1 U619 ( .B1(n150), .B2(n142), .A(n143), .ZN(n141) );
  XNOR2_X1 U620 ( .A(n41), .B(n7), .ZN(SUM[31]) );
  INV_X1 U621 ( .A(n171), .ZN(n169) );
  NAND2_X1 U622 ( .A1(B[26]), .A2(A[26]), .ZN(n89) );
  NOR2_X1 U623 ( .A1(A[26]), .A2(B[26]), .ZN(n88) );
  OAI21_X1 U624 ( .B1(n109), .B2(n433), .A(n110), .ZN(n108) );
  NAND2_X1 U625 ( .A1(B[23]), .A2(A[23]), .ZN(n118) );
  NAND2_X1 U626 ( .A1(n203), .A2(n183), .ZN(n181) );
  OAI21_X1 U627 ( .B1(n433), .B2(n120), .A(n121), .ZN(n119) );
  NOR2_X1 U628 ( .A1(n117), .A2(n126), .ZN(n115) );
  INV_X1 U629 ( .A(n437), .ZN(n125) );
  NOR2_X1 U630 ( .A1(n162), .A2(n155), .ZN(n153) );
  INV_X1 U631 ( .A(n438), .ZN(n142) );
  OAI21_X1 U632 ( .B1(n220), .B2(n181), .A(n182), .ZN(n180) );
  NOR2_X1 U633 ( .A1(n212), .A2(n205), .ZN(n203) );
  OAI21_X1 U634 ( .B1(n205), .B2(n213), .A(n206), .ZN(n204) );
  OAI21_X1 U635 ( .B1(n434), .B2(n73), .A(n74), .ZN(n72) );
  OAI21_X1 U636 ( .B1(n2), .B2(n91), .A(n92), .ZN(n90) );
  INV_X1 U637 ( .A(n4), .ZN(n109) );
  NOR2_X1 U638 ( .A1(n194), .A2(n185), .ZN(n183) );
  AOI21_X1 U639 ( .B1(n183), .B2(n204), .A(n184), .ZN(n182) );
  OAI21_X1 U640 ( .B1(n433), .B2(n102), .A(n103), .ZN(n101) );
  OAI21_X1 U641 ( .B1(n434), .B2(n82), .A(n83), .ZN(n81) );
  OAI21_X1 U642 ( .B1(n2), .B2(n53), .A(n54), .ZN(n52) );
  AOI21_X1 U643 ( .B1(n60), .B2(n417), .A(n49), .ZN(n47) );
  NAND2_X1 U644 ( .A1(A[28]), .A2(B[28]), .ZN(n71) );
  OAI21_X1 U645 ( .B1(n434), .B2(n427), .A(n177), .ZN(n175) );
  NAND2_X1 U646 ( .A1(n153), .A2(n171), .ZN(n151) );
  NAND2_X1 U647 ( .A1(n97), .A2(n77), .ZN(n6) );
  NAND2_X1 U648 ( .A1(B[25]), .A2(A[25]), .ZN(n100) );
  NOR2_X1 U649 ( .A1(n113), .A2(n151), .ZN(n111) );
  OAI21_X1 U650 ( .B1(n152), .B2(n113), .A(n114), .ZN(n112) );
  NOR2_X1 U651 ( .A1(B[20]), .A2(A[20]), .ZN(n144) );
  NOR2_X1 U652 ( .A1(n6), .A2(n46), .ZN(n44) );
  NOR2_X1 U653 ( .A1(n6), .A2(n68), .ZN(n66) );
  NOR2_X1 U654 ( .A1(n6), .A2(n57), .ZN(n55) );
  OAI21_X1 U655 ( .B1(n155), .B2(n163), .A(n156), .ZN(n154) );
  NOR2_X1 U656 ( .A1(n176), .A2(n173), .ZN(n171) );
  NAND2_X1 U657 ( .A1(n59), .A2(n417), .ZN(n46) );
  OAI21_X1 U658 ( .B1(n61), .B2(n71), .A(n62), .ZN(n60) );
  NOR2_X1 U659 ( .A1(n70), .A2(n61), .ZN(n59) );
  NAND2_X1 U660 ( .A1(n115), .A2(n135), .ZN(n113) );
  OAI21_X1 U661 ( .B1(n433), .B2(n64), .A(n65), .ZN(n63) );
  OAI21_X1 U662 ( .B1(n107), .B2(n99), .A(n100), .ZN(n98) );
  OAI21_X1 U663 ( .B1(n421), .B2(n195), .A(n186), .ZN(n184) );
  INV_X1 U664 ( .A(n185), .ZN(n298) );
  NAND2_X1 U665 ( .A1(n4), .A2(n44), .ZN(n42) );
  NAND2_X1 U666 ( .A1(n442), .A2(n104), .ZN(n102) );
  NAND2_X1 U667 ( .A1(n4), .A2(n55), .ZN(n53) );
  NAND2_X1 U668 ( .A1(n4), .A2(n66), .ZN(n64) );
  NAND2_X1 U669 ( .A1(n442), .A2(n75), .ZN(n73) );
  NAND2_X1 U670 ( .A1(n442), .A2(n84), .ZN(n82) );
  NAND2_X1 U671 ( .A1(n442), .A2(n93), .ZN(n91) );
  AOI21_X1 U672 ( .B1(n3), .B2(n44), .A(n45), .ZN(n43) );
  AOI21_X1 U673 ( .B1(n441), .B2(n93), .A(n94), .ZN(n92) );
  AOI21_X1 U674 ( .B1(n416), .B2(n104), .A(n105), .ZN(n103) );
  AOI21_X1 U675 ( .B1(n416), .B2(n75), .A(n76), .ZN(n74) );
  AOI21_X1 U676 ( .B1(n441), .B2(n84), .A(n85), .ZN(n83) );
  AOI21_X1 U677 ( .B1(n3), .B2(n55), .A(n56), .ZN(n54) );
  AOI21_X1 U678 ( .B1(n416), .B2(n66), .A(n67), .ZN(n65) );
  AOI21_X1 U679 ( .B1(n136), .B2(n429), .A(n116), .ZN(n114) );
  OAI21_X1 U680 ( .B1(n5), .B2(n46), .A(n47), .ZN(n45) );
  OAI21_X1 U681 ( .B1(n5), .B2(n57), .A(n58), .ZN(n56) );
  OAI21_X1 U682 ( .B1(n5), .B2(n68), .A(n71), .ZN(n67) );
  OAI21_X1 U683 ( .B1(n423), .B2(n89), .A(n80), .ZN(n78) );
  NAND2_X1 U684 ( .A1(B[27]), .A2(A[27]), .ZN(n80) );
  NOR2_X1 U685 ( .A1(A[27]), .A2(B[27]), .ZN(n79) );
  OAI21_X1 U686 ( .B1(n434), .B2(n42), .A(n43), .ZN(n41) );
  OAI21_X1 U687 ( .B1(n424), .B2(n145), .A(n138), .ZN(n136) );
  OAI21_X1 U688 ( .B1(n435), .B2(n127), .A(n118), .ZN(n116) );
endmodule


module datapath_DW01_add_16 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n8, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n35, n36, n37, n38, n40, n42,
         n43, n44, n45, n46, n47, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n94, n95, n96, n97, n98, n100, n101, n102, n103,
         n104, n105, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n122, n123, n124, n127, n129, n130, n131, n132,
         n133, n135, n137, n138, n139, n140, n141, n142, n143, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n162, n164, n165, n167, n169, n170, n171, n173,
         n175, n176, n177, n178, n180, n182, n183, n184, n185, n186, n187,
         n188, n190, n191, n192, n193, n194, n196, n198, n199, n200, n201,
         n203, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n217, n219, n220, n222, n224, n225, n226, n227, n228, n230,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n246, n247, n248, n249, n254, n255, n258, n261, n365, n366, n367,
         n368, n369, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411;

  CLKBUF_X1 U298 ( .A(n149), .Z(n365) );
  CLKBUF_X1 U299 ( .A(n391), .Z(n366) );
  XNOR2_X1 U300 ( .A(n45), .B(n367), .ZN(SUM[30]) );
  AND2_X1 U301 ( .A1(n232), .A2(n44), .ZN(n367) );
  OR2_X1 U302 ( .A1(n390), .A2(n108), .ZN(n368) );
  NOR2_X1 U303 ( .A1(n59), .A2(n66), .ZN(n369) );
  AND2_X1 U304 ( .A1(B[19]), .A2(A[19]), .ZN(n374) );
  INV_X1 U305 ( .A(n374), .ZN(n122) );
  AND2_X1 U306 ( .A1(n372), .A2(n230), .ZN(SUM[0]) );
  OR2_X1 U307 ( .A1(n43), .A2(n50), .ZN(n371) );
  OR2_X1 U308 ( .A1(B[0]), .A2(A[0]), .ZN(n372) );
  AOI21_X1 U309 ( .B1(n85), .B2(n102), .A(n86), .ZN(n373) );
  NOR2_X1 U310 ( .A1(B[16]), .A2(A[16]), .ZN(n375) );
  NOR2_X1 U311 ( .A1(B[16]), .A2(A[16]), .ZN(n141) );
  XNOR2_X1 U312 ( .A(n61), .B(n376), .ZN(SUM[28]) );
  AND2_X1 U313 ( .A1(n234), .A2(n60), .ZN(n376) );
  XNOR2_X1 U314 ( .A(n96), .B(n377), .ZN(SUM[23]) );
  AND2_X1 U315 ( .A1(n239), .A2(n95), .ZN(n377) );
  XNOR2_X1 U316 ( .A(n105), .B(n378), .ZN(SUM[22]) );
  AND2_X1 U317 ( .A1(n240), .A2(n104), .ZN(n378) );
  XNOR2_X1 U318 ( .A(n89), .B(n379), .ZN(SUM[24]) );
  AND2_X1 U319 ( .A1(n238), .A2(n88), .ZN(n379) );
  NOR2_X1 U320 ( .A1(B[26]), .A2(A[26]), .ZN(n380) );
  NOR2_X1 U321 ( .A1(B[26]), .A2(A[26]), .ZN(n75) );
  AOI21_X1 U322 ( .B1(n403), .B2(n127), .A(n374), .ZN(n381) );
  XNOR2_X1 U323 ( .A(n77), .B(n382), .ZN(SUM[26]) );
  AND2_X1 U324 ( .A1(n236), .A2(n76), .ZN(n382) );
  OAI21_X1 U325 ( .B1(n75), .B2(n81), .A(n76), .ZN(n383) );
  NOR2_X1 U326 ( .A1(A[28]), .A2(B[28]), .ZN(n384) );
  CLKBUF_X1 U327 ( .A(n114), .Z(n385) );
  CLKBUF_X1 U328 ( .A(n140), .Z(n386) );
  CLKBUF_X1 U329 ( .A(n392), .Z(n387) );
  NOR2_X1 U330 ( .A1(n94), .A2(n391), .ZN(n388) );
  AOI21_X1 U331 ( .B1(n57), .B2(n74), .A(n58), .ZN(n389) );
  NOR2_X1 U332 ( .A1(B[22]), .A2(A[22]), .ZN(n390) );
  NOR2_X1 U333 ( .A1(B[24]), .A2(A[24]), .ZN(n391) );
  NOR2_X1 U334 ( .A1(B[20]), .A2(A[20]), .ZN(n114) );
  OAI21_X1 U335 ( .B1(n132), .B2(n149), .A(n133), .ZN(n392) );
  AOI21_X1 U336 ( .B1(n392), .B2(n112), .A(n113), .ZN(n393) );
  XNOR2_X1 U337 ( .A(n36), .B(n394), .ZN(SUM[31]) );
  AND2_X1 U338 ( .A1(n411), .A2(n35), .ZN(n394) );
  CLKBUF_X1 U339 ( .A(n139), .Z(n395) );
  XNOR2_X1 U340 ( .A(n68), .B(n396), .ZN(SUM[27]) );
  AND2_X1 U341 ( .A1(n235), .A2(n67), .ZN(n396) );
  XNOR2_X1 U342 ( .A(n52), .B(n397), .ZN(SUM[29]) );
  AND2_X1 U343 ( .A1(n233), .A2(n51), .ZN(n397) );
  AOI21_X1 U344 ( .B1(n112), .B2(n131), .A(n113), .ZN(n111) );
  OAI21_X1 U345 ( .B1(n393), .B2(n83), .A(n373), .ZN(n398) );
  OAI21_X1 U346 ( .B1(n111), .B2(n83), .A(n84), .ZN(n399) );
  OAI21_X1 U347 ( .B1(n83), .B2(n111), .A(n373), .ZN(n82) );
  NOR2_X1 U348 ( .A1(B[28]), .A2(A[28]), .ZN(n59) );
  OR2_X1 U349 ( .A1(B[9]), .A2(A[9]), .ZN(n400) );
  OR2_X1 U350 ( .A1(B[10]), .A2(A[10]), .ZN(n401) );
  OR2_X1 U351 ( .A1(B[17]), .A2(A[17]), .ZN(n402) );
  OR2_X1 U352 ( .A1(B[19]), .A2(A[19]), .ZN(n403) );
  OR2_X1 U353 ( .A1(B[2]), .A2(A[2]), .ZN(n404) );
  OR2_X1 U354 ( .A1(B[12]), .A2(A[12]), .ZN(n405) );
  OR2_X1 U355 ( .A1(A[18]), .A2(B[18]), .ZN(n406) );
  OR2_X1 U356 ( .A1(B[11]), .A2(A[11]), .ZN(n407) );
  OR2_X1 U357 ( .A1(B[3]), .A2(A[3]), .ZN(n408) );
  OR2_X1 U358 ( .A1(B[5]), .A2(A[5]), .ZN(n409) );
  OR2_X1 U359 ( .A1(B[6]), .A2(A[6]), .ZN(n410) );
  OR2_X1 U360 ( .A1(B[31]), .A2(A[31]), .ZN(n411) );
  NAND2_X1 U361 ( .A1(B[0]), .A2(A[0]), .ZN(n230) );
  NAND2_X1 U362 ( .A1(n258), .A2(n212), .ZN(n29) );
  NAND2_X1 U363 ( .A1(n404), .A2(n224), .ZN(n31) );
  INV_X1 U364 ( .A(n210), .ZN(n208) );
  NAND2_X1 U365 ( .A1(B[31]), .A2(A[31]), .ZN(n35) );
  NAND2_X1 U366 ( .A1(B[4]), .A2(A[4]), .ZN(n212) );
  NAND2_X1 U367 ( .A1(n408), .A2(n404), .ZN(n214) );
  NAND2_X1 U368 ( .A1(B[2]), .A2(A[2]), .ZN(n224) );
  INV_X1 U369 ( .A(n209), .ZN(n207) );
  NOR2_X1 U370 ( .A1(n211), .A2(n214), .ZN(n209) );
  INV_X1 U371 ( .A(n224), .ZN(n222) );
  AOI21_X1 U372 ( .B1(n408), .B2(n222), .A(n217), .ZN(n215) );
  OAI21_X1 U373 ( .B1(n211), .B2(n215), .A(n212), .ZN(n210) );
  NAND2_X1 U374 ( .A1(n408), .A2(n219), .ZN(n30) );
  INV_X1 U375 ( .A(n219), .ZN(n217) );
  NAND2_X1 U376 ( .A1(B[3]), .A2(A[3]), .ZN(n219) );
  INV_X1 U377 ( .A(n211), .ZN(n258) );
  NOR2_X1 U378 ( .A1(B[4]), .A2(A[4]), .ZN(n211) );
  NAND2_X1 U379 ( .A1(B[5]), .A2(A[5]), .ZN(n205) );
  NAND2_X1 U380 ( .A1(n255), .A2(n192), .ZN(n26) );
  INV_X1 U381 ( .A(n192), .ZN(n190) );
  NAND2_X1 U382 ( .A1(B[7]), .A2(A[7]), .ZN(n192) );
  NAND2_X1 U383 ( .A1(n254), .A2(n187), .ZN(n25) );
  INV_X1 U384 ( .A(n191), .ZN(n255) );
  NOR2_X1 U385 ( .A1(B[7]), .A2(A[7]), .ZN(n191) );
  INV_X1 U386 ( .A(n205), .ZN(n203) );
  INV_X1 U387 ( .A(n235), .ZN(n64) );
  INV_X1 U388 ( .A(n239), .ZN(n92) );
  INV_X1 U389 ( .A(n368), .ZN(n97) );
  NAND2_X1 U390 ( .A1(B[8]), .A2(A[8]), .ZN(n187) );
  NAND2_X1 U391 ( .A1(B[30]), .A2(A[30]), .ZN(n44) );
  NAND2_X1 U392 ( .A1(B[29]), .A2(A[29]), .ZN(n51) );
  INV_X1 U393 ( .A(n100), .ZN(n98) );
  NAND2_X1 U394 ( .A1(n400), .A2(n182), .ZN(n24) );
  NAND2_X1 U395 ( .A1(B[9]), .A2(A[9]), .ZN(n182) );
  NAND2_X1 U396 ( .A1(n242), .A2(n115), .ZN(n13) );
  INV_X1 U397 ( .A(n226), .ZN(n225) );
  OAI21_X1 U398 ( .B1(n43), .B2(n51), .A(n44), .ZN(n42) );
  INV_X1 U399 ( .A(n71), .ZN(n69) );
  NOR2_X1 U400 ( .A1(n71), .A2(n64), .ZN(n62) );
  NAND2_X1 U401 ( .A1(B[1]), .A2(A[1]), .ZN(n228) );
  NAND2_X1 U402 ( .A1(n237), .A2(n81), .ZN(n8) );
  INV_X1 U403 ( .A(n81), .ZN(n79) );
  NAND2_X1 U404 ( .A1(B[25]), .A2(A[25]), .ZN(n81) );
  NOR2_X1 U405 ( .A1(n59), .A2(n66), .ZN(n57) );
  NOR2_X1 U406 ( .A1(n380), .A2(n80), .ZN(n73) );
  NAND2_X1 U407 ( .A1(n247), .A2(n147), .ZN(n18) );
  INV_X1 U408 ( .A(n147), .ZN(n145) );
  NAND2_X1 U409 ( .A1(B[15]), .A2(A[15]), .ZN(n147) );
  NOR2_X1 U410 ( .A1(n368), .A2(n92), .ZN(n90) );
  NAND2_X1 U411 ( .A1(n402), .A2(n137), .ZN(n16) );
  NAND2_X1 U412 ( .A1(B[28]), .A2(A[28]), .ZN(n60) );
  OAI21_X1 U413 ( .B1(n100), .B2(n92), .A(n95), .ZN(n91) );
  NAND2_X1 U414 ( .A1(n248), .A2(n153), .ZN(n19) );
  NAND2_X1 U415 ( .A1(B[14]), .A2(A[14]), .ZN(n153) );
  INV_X1 U416 ( .A(n406), .ZN(n124) );
  NAND2_X1 U417 ( .A1(B[22]), .A2(A[22]), .ZN(n104) );
  NAND2_X1 U418 ( .A1(n405), .A2(n164), .ZN(n21) );
  NAND2_X1 U419 ( .A1(n409), .A2(n209), .ZN(n200) );
  AOI21_X1 U420 ( .B1(n409), .B2(n210), .A(n203), .ZN(n201) );
  NAND2_X1 U421 ( .A1(n246), .A2(n142), .ZN(n17) );
  NAND2_X1 U422 ( .A1(B[26]), .A2(A[26]), .ZN(n76) );
  NAND2_X1 U423 ( .A1(B[27]), .A2(A[27]), .ZN(n67) );
  INV_X1 U424 ( .A(n182), .ZN(n180) );
  NAND2_X1 U425 ( .A1(B[24]), .A2(A[24]), .ZN(n88) );
  NAND2_X1 U426 ( .A1(n406), .A2(n129), .ZN(n15) );
  NAND2_X1 U427 ( .A1(B[23]), .A2(A[23]), .ZN(n95) );
  INV_X1 U428 ( .A(n175), .ZN(n173) );
  NAND2_X1 U429 ( .A1(B[10]), .A2(A[10]), .ZN(n175) );
  INV_X1 U430 ( .A(n42), .ZN(n40) );
  NAND2_X1 U431 ( .A1(B[20]), .A2(A[20]), .ZN(n115) );
  INV_X1 U432 ( .A(n186), .ZN(n254) );
  OAI21_X1 U433 ( .B1(n186), .B2(n192), .A(n187), .ZN(n185) );
  NOR2_X1 U434 ( .A1(B[8]), .A2(A[8]), .ZN(n186) );
  NAND2_X1 U435 ( .A1(B[13]), .A2(A[13]), .ZN(n156) );
  INV_X1 U436 ( .A(n72), .ZN(n70) );
  OAI21_X1 U437 ( .B1(n72), .B2(n64), .A(n67), .ZN(n63) );
  NAND2_X1 U438 ( .A1(B[17]), .A2(A[17]), .ZN(n137) );
  INV_X1 U439 ( .A(n146), .ZN(n247) );
  NOR2_X1 U440 ( .A1(B[15]), .A2(A[15]), .ZN(n146) );
  NAND2_X1 U441 ( .A1(B[12]), .A2(A[12]), .ZN(n164) );
  NAND2_X1 U442 ( .A1(n403), .A2(n122), .ZN(n14) );
  INV_X1 U443 ( .A(n55), .ZN(n53) );
  NOR2_X1 U444 ( .A1(n55), .A2(n50), .ZN(n46) );
  NOR2_X1 U445 ( .A1(n55), .A2(n371), .ZN(n37) );
  NAND2_X1 U446 ( .A1(n73), .A2(n369), .ZN(n55) );
  NAND2_X1 U447 ( .A1(B[11]), .A2(A[11]), .ZN(n169) );
  NOR2_X1 U448 ( .A1(n186), .A2(n191), .ZN(n184) );
  INV_X1 U449 ( .A(n383), .ZN(n72) );
  OAI21_X1 U450 ( .B1(n75), .B2(n81), .A(n76), .ZN(n74) );
  NAND2_X1 U451 ( .A1(B[16]), .A2(A[16]), .ZN(n142) );
  INV_X1 U452 ( .A(n155), .ZN(n249) );
  NOR2_X1 U453 ( .A1(B[13]), .A2(A[13]), .ZN(n155) );
  INV_X1 U454 ( .A(n129), .ZN(n127) );
  NAND2_X1 U455 ( .A1(B[18]), .A2(A[18]), .ZN(n129) );
  INV_X1 U456 ( .A(n137), .ZN(n135) );
  AOI21_X1 U457 ( .B1(n410), .B2(n199), .A(n196), .ZN(n194) );
  OAI21_X1 U458 ( .B1(n225), .B2(n200), .A(n201), .ZN(n199) );
  INV_X1 U459 ( .A(n73), .ZN(n71) );
  INV_X1 U460 ( .A(n164), .ZN(n162) );
  INV_X1 U461 ( .A(n169), .ZN(n167) );
  INV_X1 U462 ( .A(n108), .ZN(n241) );
  NOR2_X1 U463 ( .A1(B[21]), .A2(A[21]), .ZN(n108) );
  INV_X1 U464 ( .A(n80), .ZN(n237) );
  NOR2_X1 U465 ( .A1(B[25]), .A2(A[25]), .ZN(n80) );
  NOR2_X1 U466 ( .A1(n390), .A2(n108), .ZN(n101) );
  NAND2_X1 U467 ( .A1(n184), .A2(n400), .ZN(n177) );
  INV_X1 U468 ( .A(n385), .ZN(n242) );
  INV_X1 U469 ( .A(n152), .ZN(n248) );
  OAI21_X1 U470 ( .B1(n152), .B2(n156), .A(n153), .ZN(n151) );
  NOR2_X1 U471 ( .A1(n155), .A2(n152), .ZN(n150) );
  NOR2_X1 U472 ( .A1(B[14]), .A2(A[14]), .ZN(n152) );
  INV_X1 U473 ( .A(n198), .ZN(n196) );
  NAND2_X1 U474 ( .A1(B[6]), .A2(A[6]), .ZN(n198) );
  INV_X1 U475 ( .A(n103), .ZN(n240) );
  NOR2_X1 U476 ( .A1(B[22]), .A2(A[22]), .ZN(n103) );
  INV_X1 U477 ( .A(n94), .ZN(n239) );
  NOR2_X1 U478 ( .A1(n94), .A2(n391), .ZN(n85) );
  NOR2_X1 U479 ( .A1(B[23]), .A2(A[23]), .ZN(n94) );
  INV_X1 U480 ( .A(n102), .ZN(n100) );
  AOI21_X1 U481 ( .B1(n85), .B2(n102), .A(n86), .ZN(n84) );
  OAI21_X1 U482 ( .B1(n103), .B2(n109), .A(n104), .ZN(n102) );
  INV_X1 U483 ( .A(n375), .ZN(n246) );
  INV_X1 U484 ( .A(n389), .ZN(n54) );
  OAI21_X1 U485 ( .B1(n56), .B2(n50), .A(n51), .ZN(n47) );
  OAI21_X1 U486 ( .B1(n389), .B2(n371), .A(n40), .ZN(n38) );
  AOI21_X1 U487 ( .B1(n57), .B2(n383), .A(n58), .ZN(n56) );
  INV_X1 U488 ( .A(n43), .ZN(n232) );
  NOR2_X1 U489 ( .A1(B[30]), .A2(A[30]), .ZN(n43) );
  AOI21_X1 U490 ( .B1(n405), .B2(n167), .A(n162), .ZN(n160) );
  INV_X1 U491 ( .A(n366), .ZN(n238) );
  OAI21_X1 U492 ( .B1(n87), .B2(n95), .A(n88), .ZN(n86) );
  NOR2_X1 U493 ( .A1(A[24]), .A2(B[24]), .ZN(n87) );
  OAI21_X1 U494 ( .B1(n141), .B2(n147), .A(n142), .ZN(n140) );
  NAND2_X1 U495 ( .A1(n406), .A2(n403), .ZN(n117) );
  NAND2_X1 U496 ( .A1(n241), .A2(n109), .ZN(n12) );
  INV_X1 U497 ( .A(n109), .ZN(n107) );
  NAND2_X1 U498 ( .A1(B[21]), .A2(A[21]), .ZN(n109) );
  NOR2_X1 U499 ( .A1(n375), .A2(n146), .ZN(n139) );
  OAI21_X1 U500 ( .B1(n159), .B2(n171), .A(n160), .ZN(n158) );
  NAND2_X1 U501 ( .A1(n407), .A2(n405), .ZN(n159) );
  INV_X1 U502 ( .A(n50), .ZN(n233) );
  NOR2_X1 U503 ( .A1(B[29]), .A2(A[29]), .ZN(n50) );
  OAI21_X1 U504 ( .B1(n194), .B2(n177), .A(n178), .ZN(n176) );
  AOI21_X1 U505 ( .B1(n185), .B2(n400), .A(n180), .ZN(n178) );
  INV_X1 U506 ( .A(n59), .ZN(n234) );
  OAI21_X1 U507 ( .B1(n384), .B2(n67), .A(n60), .ZN(n58) );
  INV_X1 U508 ( .A(n66), .ZN(n235) );
  NOR2_X1 U509 ( .A1(B[27]), .A2(A[27]), .ZN(n66) );
  INV_X1 U510 ( .A(n380), .ZN(n236) );
  NAND2_X1 U511 ( .A1(n388), .A2(n101), .ZN(n83) );
  NOR2_X1 U512 ( .A1(n117), .A2(n114), .ZN(n112) );
  AOI21_X1 U513 ( .B1(n403), .B2(n127), .A(n374), .ZN(n118) );
  NAND2_X1 U514 ( .A1(n139), .A2(n402), .ZN(n132) );
  AOI21_X1 U515 ( .B1(n140), .B2(n402), .A(n135), .ZN(n133) );
  AOI21_X1 U516 ( .B1(n150), .B2(n158), .A(n151), .ZN(n149) );
  INV_X1 U517 ( .A(n227), .ZN(n261) );
  OAI21_X1 U518 ( .B1(n227), .B2(n230), .A(n228), .ZN(n226) );
  NOR2_X1 U519 ( .A1(B[1]), .A2(A[1]), .ZN(n227) );
  OAI21_X1 U520 ( .B1(n118), .B2(n114), .A(n115), .ZN(n113) );
  OAI21_X1 U521 ( .B1(n132), .B2(n149), .A(n133), .ZN(n131) );
  AOI21_X1 U522 ( .B1(n176), .B2(n401), .A(n173), .ZN(n171) );
  XOR2_X1 U523 ( .A(n220), .B(n30), .Z(SUM[3]) );
  AOI21_X1 U524 ( .B1(n226), .B2(n404), .A(n222), .ZN(n220) );
  XOR2_X1 U525 ( .A(n225), .B(n31), .Z(SUM[2]) );
  NAND2_X1 U526 ( .A1(n409), .A2(n205), .ZN(n28) );
  XNOR2_X1 U527 ( .A(n206), .B(n28), .ZN(SUM[5]) );
  OAI21_X1 U528 ( .B1(n225), .B2(n207), .A(n208), .ZN(n206) );
  XNOR2_X1 U529 ( .A(n213), .B(n29), .ZN(SUM[4]) );
  OAI21_X1 U530 ( .B1(n225), .B2(n214), .A(n215), .ZN(n213) );
  XOR2_X1 U531 ( .A(n32), .B(n230), .Z(SUM[1]) );
  NAND2_X1 U532 ( .A1(n261), .A2(n228), .ZN(n32) );
  XNOR2_X1 U533 ( .A(n193), .B(n26), .ZN(SUM[7]) );
  INV_X1 U534 ( .A(n194), .ZN(n193) );
  XNOR2_X1 U535 ( .A(n27), .B(n199), .ZN(SUM[6]) );
  NAND2_X1 U536 ( .A1(n410), .A2(n198), .ZN(n27) );
  XNOR2_X1 U537 ( .A(n176), .B(n23), .ZN(SUM[10]) );
  NAND2_X1 U538 ( .A1(n401), .A2(n175), .ZN(n23) );
  XOR2_X1 U539 ( .A(n188), .B(n25), .Z(SUM[8]) );
  AOI21_X1 U540 ( .B1(n193), .B2(n255), .A(n190), .ZN(n188) );
  XOR2_X1 U541 ( .A(n183), .B(n24), .Z(SUM[9]) );
  AOI21_X1 U542 ( .B1(n193), .B2(n184), .A(n185), .ZN(n183) );
  NAND2_X1 U543 ( .A1(n407), .A2(n169), .ZN(n22) );
  XNOR2_X1 U544 ( .A(n22), .B(n170), .ZN(SUM[11]) );
  INV_X1 U545 ( .A(n171), .ZN(n170) );
  NAND2_X1 U546 ( .A1(n249), .A2(n156), .ZN(n20) );
  XOR2_X1 U547 ( .A(n165), .B(n21), .Z(SUM[12]) );
  AOI21_X1 U548 ( .B1(n170), .B2(n407), .A(n167), .ZN(n165) );
  XOR2_X1 U549 ( .A(n157), .B(n20), .Z(SUM[13]) );
  INV_X1 U550 ( .A(n158), .ZN(n157) );
  XNOR2_X1 U551 ( .A(n154), .B(n19), .ZN(SUM[14]) );
  OAI21_X1 U552 ( .B1(n157), .B2(n155), .A(n156), .ZN(n154) );
  XNOR2_X1 U553 ( .A(n148), .B(n18), .ZN(SUM[15]) );
  INV_X1 U554 ( .A(n365), .ZN(n148) );
  XOR2_X1 U555 ( .A(n143), .B(n17), .Z(SUM[16]) );
  AOI21_X1 U556 ( .B1(n148), .B2(n247), .A(n145), .ZN(n143) );
  XOR2_X1 U557 ( .A(n138), .B(n16), .Z(SUM[17]) );
  AOI21_X1 U558 ( .B1(n148), .B2(n395), .A(n386), .ZN(n138) );
  XOR2_X1 U559 ( .A(n130), .B(n15), .Z(SUM[18]) );
  INV_X1 U560 ( .A(n387), .ZN(n130) );
  XNOR2_X1 U561 ( .A(n123), .B(n14), .ZN(SUM[19]) );
  OAI21_X1 U562 ( .B1(n130), .B2(n124), .A(n129), .ZN(n123) );
  XNOR2_X1 U563 ( .A(n116), .B(n13), .ZN(SUM[20]) );
  OAI21_X1 U564 ( .B1(n130), .B2(n117), .A(n381), .ZN(n116) );
  XNOR2_X1 U565 ( .A(n110), .B(n12), .ZN(SUM[21]) );
  INV_X1 U566 ( .A(n393), .ZN(n110) );
  AOI21_X1 U567 ( .B1(n110), .B2(n97), .A(n98), .ZN(n96) );
  AOI21_X1 U568 ( .B1(n110), .B2(n241), .A(n107), .ZN(n105) );
  AOI21_X1 U569 ( .B1(n110), .B2(n90), .A(n91), .ZN(n89) );
  XNOR2_X1 U570 ( .A(n398), .B(n8), .ZN(SUM[25]) );
  AOI21_X1 U571 ( .B1(n399), .B2(n69), .A(n70), .ZN(n68) );
  AOI21_X1 U572 ( .B1(n399), .B2(n53), .A(n54), .ZN(n52) );
  AOI21_X1 U573 ( .B1(n398), .B2(n237), .A(n79), .ZN(n77) );
  AOI21_X1 U574 ( .B1(n399), .B2(n62), .A(n63), .ZN(n61) );
  AOI21_X1 U575 ( .B1(n82), .B2(n46), .A(n47), .ZN(n45) );
  AOI21_X1 U576 ( .B1(n82), .B2(n37), .A(n38), .ZN(n36) );
endmodule


module datapath ( clk, data_in, addr_x, wr_en_x, addr_a1, addr_a2, addr_a3, 
        addr_a4, addr_a5, addr_a6, addr_a7, addr_a8, wr_en_a1, wr_en_a2, 
        wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6, wr_en_a7, wr_en_a8, addr_y, 
        wr_en_y, clear_acc, clc, clc1, data_out );
  input [15:0] data_in;
  input [2:0] addr_x;
  input [2:0] addr_a1;
  input [2:0] addr_a2;
  input [2:0] addr_a3;
  input [2:0] addr_a4;
  input [2:0] addr_a5;
  input [2:0] addr_a6;
  input [2:0] addr_a7;
  input [2:0] addr_a8;
  input [2:0] addr_y;
  output [31:0] data_out;
  input clk, wr_en_x, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5,
         wr_en_a6, wr_en_a7, wr_en_a8, wr_en_y, clear_acc, clc, clc1;
  wire   n16, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n274, n275, n276, n277, n280, n281, n285,
         n286, n287, n288, n291, n292, n295, n296, n299, n300, n303, n304,
         n307, n308, n311, n312, n315, n316, n319, n320, n323, n324, n327,
         n328, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n410, n411, n412, n413, n414, n415, n416, n417, n419, n420,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, \mul_out1[9] , \mul_out1[8] , \mul_out1[7] ,
         \mul_out1[6] , \mul_out1[5] , \mul_out1[4] , \mul_out1[3] ,
         \mul_out1[31] , \mul_out1[30] , \mul_out1[2] , \mul_out1[29] ,
         \mul_out1[28] , \mul_out1[27] , \mul_out1[26] , \mul_out1[25] ,
         \mul_out1[24] , \mul_out1[23] , \mul_out1[22] , \mul_out1[21] ,
         \mul_out1[20] , \mul_out1[1] , \mul_out1[19] , \mul_out1[18] ,
         \mul_out1[17] , \mul_out1[16] , \mul_out1[15] , \mul_out1[14] ,
         \mul_out1[13] , \mul_out1[12] , \mul_out1[11] , \mul_out1[10] ,
         \mul_out1[0] , \mul_out2[9] , \mul_out2[8] , \mul_out2[7] ,
         \mul_out2[6] , \mul_out2[5] , \mul_out2[4] , \mul_out2[3] ,
         \mul_out2[31] , \mul_out2[30] , \mul_out2[2] , \mul_out2[29] ,
         \mul_out2[28] , \mul_out2[27] , \mul_out2[26] , \mul_out2[25] ,
         \mul_out2[24] , \mul_out2[23] , \mul_out2[22] , \mul_out2[21] ,
         \mul_out2[20] , \mul_out2[1] , \mul_out2[19] , \mul_out2[18] ,
         \mul_out2[17] , \mul_out2[16] , \mul_out2[15] , \mul_out2[14] ,
         \mul_out2[13] , \mul_out2[12] , \mul_out2[11] , \mul_out2[10] ,
         \mul_out2[0] , \mul_out3[9] , \mul_out3[8] , \mul_out3[7] ,
         \mul_out3[6] , \mul_out3[5] , \mul_out3[4] , \mul_out3[3] ,
         \mul_out3[31] , \mul_out3[30] , \mul_out3[2] , \mul_out3[29] ,
         \mul_out3[28] , \mul_out3[27] , \mul_out3[26] , \mul_out3[25] ,
         \mul_out3[24] , \mul_out3[23] , \mul_out3[22] , \mul_out3[21] ,
         \mul_out3[20] , \mul_out3[1] , \mul_out3[19] , \mul_out3[18] ,
         \mul_out3[17] , \mul_out3[16] , \mul_out3[15] , \mul_out3[14] ,
         \mul_out3[13] , \mul_out3[12] , \mul_out3[11] , \mul_out3[10] ,
         \mul_out3[0] , \mul_out4[9] , \mul_out4[8] , \mul_out4[7] ,
         \mul_out4[6] , \mul_out4[5] , \mul_out4[4] , \mul_out4[3] ,
         \mul_out4[31] , \mul_out4[30] , \mul_out4[2] , \mul_out4[29] ,
         \mul_out4[28] , \mul_out4[27] , \mul_out4[26] , \mul_out4[25] ,
         \mul_out4[24] , \mul_out4[23] , \mul_out4[22] , \mul_out4[21] ,
         \mul_out4[20] , \mul_out4[1] , \mul_out4[19] , \mul_out4[18] ,
         \mul_out4[17] , \mul_out4[16] , \mul_out4[15] , \mul_out4[14] ,
         \mul_out4[13] , \mul_out4[12] , \mul_out4[11] , \mul_out4[10] ,
         \mul_out4[0] , \mul_out5[9] , \mul_out5[8] , \mul_out5[7] ,
         \mul_out5[6] , \mul_out5[5] , \mul_out5[4] , \mul_out5[3] ,
         \mul_out5[31] , \mul_out5[30] , \mul_out5[2] , \mul_out5[29] ,
         \mul_out5[28] , \mul_out5[27] , \mul_out5[26] , \mul_out5[25] ,
         \mul_out5[24] , \mul_out5[23] , \mul_out5[22] , \mul_out5[21] ,
         \mul_out5[20] , \mul_out5[1] , \mul_out5[19] , \mul_out5[18] ,
         \mul_out5[17] , \mul_out5[16] , \mul_out5[15] , \mul_out5[14] ,
         \mul_out5[13] , \mul_out5[12] , \mul_out5[11] , \mul_out5[10] ,
         \mul_out5[0] , \mul_out6[9] , \mul_out6[8] , \mul_out6[7] ,
         \mul_out6[6] , \mul_out6[5] , \mul_out6[4] , \mul_out6[3] ,
         \mul_out6[31] , \mul_out6[30] , \mul_out6[2] , \mul_out6[29] ,
         \mul_out6[28] , \mul_out6[27] , \mul_out6[26] , \mul_out6[25] ,
         \mul_out6[24] , \mul_out6[23] , \mul_out6[22] , \mul_out6[21] ,
         \mul_out6[20] , \mul_out6[1] , \mul_out6[19] , \mul_out6[18] ,
         \mul_out6[17] , \mul_out6[16] , \mul_out6[15] , \mul_out6[14] ,
         \mul_out6[13] , \mul_out6[12] , \mul_out6[11] , \mul_out6[10] ,
         \mul_out6[0] , \mul_out7[9] , \mul_out7[8] , \mul_out7[7] ,
         \mul_out7[6] , \mul_out7[5] , \mul_out7[4] , \mul_out7[3] ,
         \mul_out7[31] , \mul_out7[30] , \mul_out7[2] , \mul_out7[29] ,
         \mul_out7[28] , \mul_out7[27] , \mul_out7[26] , \mul_out7[25] ,
         \mul_out7[24] , \mul_out7[23] , \mul_out7[22] , \mul_out7[21] ,
         \mul_out7[20] , \mul_out7[1] , \mul_out7[19] , \mul_out7[18] ,
         \mul_out7[17] , \mul_out7[16] , \mul_out7[15] , \mul_out7[14] ,
         \mul_out7[13] , \mul_out7[12] , \mul_out7[11] , \mul_out7[10] ,
         \mul_out7[0] , \mul_out8[9] , \mul_out8[8] , \mul_out8[7] ,
         \mul_out8[6] , \mul_out8[5] , \mul_out8[4] , \mul_out8[3] ,
         \mul_out8[31] , \mul_out8[30] , \mul_out8[2] , \mul_out8[29] ,
         \mul_out8[28] , \mul_out8[27] , \mul_out8[26] , \mul_out8[25] ,
         \mul_out8[24] , \mul_out8[23] , \mul_out8[22] , \mul_out8[21] ,
         \mul_out8[20] , \mul_out8[1] , \mul_out8[19] , \mul_out8[18] ,
         \mul_out8[17] , \mul_out8[16] , \mul_out8[15] , \mul_out8[14] ,
         \mul_out8[13] , \mul_out8[12] , \mul_out8[11] , \mul_out8[10] ,
         \mul_out8[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n17, n18, n19, n20, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n96, n97, n98, n99, n100, n101, n102, n103, n104, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n278, n279, n282, n283,
         n284, n289, n290, n293, n294, n297, n298, n301, n302, n305, n306,
         n309, n310, n313, n314, n317, n318, n321, n322, n325, n326, n329,
         n330, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n418, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071;
  wire   [15:0] data_out_x;
  wire   [15:0] data_out_a1;
  wire   [15:0] data_out_a2;
  wire   [15:0] data_out_a3;
  wire   [15:0] data_out_a4;
  wire   [15:0] data_out_a5;
  wire   [15:0] data_out_a6;
  wire   [15:0] data_out_a7;
  wire   [15:0] data_out_a8;
  wire   [31:0] f;
  wire   [31:0] f1;
  wire   [31:0] f2;
  wire   [31:0] f3;
  wire   [31:0] f4;
  wire   [31:0] f5;
  wire   [31:0] f6;
  wire   [31:0] f7;
  wire   [31:0] f8;
  wire   [31:0] add_r1;
  wire   [31:0] add_r2;
  wire   [31:0] add_r3;
  wire   [31:0] add_r4;
  wire   [31:0] add_r5;
  wire   [31:0] add_r6;
  wire   [31:0] add_r7;
  wire   [31:0] add_r8;

  DFF_X1 \f1_reg[31]  ( .D(n966), .CK(clk), .Q(f1[31]), .QN(n1058) );
  DFF_X1 \f1_reg[29]  ( .D(n964), .CK(clk), .Q(f1[29]), .QN(n1050) );
  DFF_X1 \f1_reg[23]  ( .D(n958), .CK(clk), .Q(f1[23]), .QN(n1027) );
  DFF_X1 \f1_reg[22]  ( .D(n957), .CK(clk), .Q(f1[22]), .QN(n1023) );
  DFF_X1 \f1_reg[21]  ( .D(n956), .CK(clk), .Q(f1[21]), .QN(n1019) );
  DFF_X1 \f1_reg[20]  ( .D(n955), .CK(clk), .Q(f1[20]), .QN(n1015) );
  DFF_X1 \f1_reg[19]  ( .D(n954), .CK(clk), .Q(f1[19]), .QN(n21) );
  DFF_X1 \f1_reg[18]  ( .D(n953), .CK(clk), .Q(f1[18]), .QN(n22) );
  DFF_X1 \f1_reg[17]  ( .D(n952), .CK(clk), .Q(f1[17]), .QN(n23) );
  DFF_X1 \f2_reg[24]  ( .D(n927), .CK(clk), .Q(f2[24]), .QN(n48) );
  DFF_X1 \f2_reg[23]  ( .D(n926), .CK(clk), .Q(n650), .QN(n49) );
  DFF_X1 \f2_reg[22]  ( .D(n925), .CK(clk), .Q(n652), .QN(n50) );
  DFF_X1 \f2_reg[21]  ( .D(n924), .CK(clk), .Q(n654), .QN(n51) );
  DFF_X1 \f2_reg[20]  ( .D(n923), .CK(clk), .Q(n656), .QN(n52) );
  DFF_X1 \f2_reg[19]  ( .D(n922), .CK(clk), .Q(n658), .QN(n53) );
  DFF_X1 \f2_reg[18]  ( .D(n921), .CK(clk), .Q(n660), .QN(n54) );
  DFF_X1 \f2_reg[17]  ( .D(n920), .CK(clk), .Q(n662), .QN(n55) );
  DFF_X1 \f3_reg[24]  ( .D(n895), .CK(clk), .Q(n577), .QN(n80) );
  DFF_X1 \f3_reg[23]  ( .D(n894), .CK(clk), .Q(n579), .QN(n81) );
  DFF_X1 \f3_reg[22]  ( .D(n893), .CK(clk), .Q(n581), .QN(n82) );
  DFF_X1 \f3_reg[21]  ( .D(n892), .CK(clk), .Q(f3[21]), .QN(n83) );
  DFF_X1 \f3_reg[20]  ( .D(n891), .CK(clk), .Q(f3[20]), .QN(n84) );
  DFF_X1 \f3_reg[19]  ( .D(n890), .CK(clk), .Q(f3[19]), .QN(n85) );
  DFF_X1 \f3_reg[18]  ( .D(n889), .CK(clk), .Q(f3[18]), .QN(n86) );
  DFF_X1 \f3_reg[17]  ( .D(n888), .CK(clk), .Q(f3[17]), .QN(n87) );
  DFF_X1 \f4_reg[31]  ( .D(n870), .CK(clk), .Q(f4[31]), .QN(n105) );
  DFF_X1 \f4_reg[30]  ( .D(n869), .CK(clk), .Q(f4[30]), .QN(n106) );
  DFF_X1 \f4_reg[29]  ( .D(n868), .CK(clk), .Q(f4[29]), .QN(n107) );
  DFF_X1 \f4_reg[26]  ( .D(n865), .CK(clk), .Q(f4[26]), .QN(n110) );
  DFF_X1 \f4_reg[24]  ( .D(n863), .CK(clk), .Q(f4[24]), .QN(n112) );
  DFF_X1 \f4_reg[23]  ( .D(n862), .CK(clk), .Q(f4[23]), .QN(n113) );
  DFF_X1 \f4_reg[22]  ( .D(n861), .CK(clk), .Q(f4[22]), .QN(n114) );
  DFF_X1 \f4_reg[20]  ( .D(n859), .CK(clk), .Q(f4[20]), .QN(n116) );
  DFF_X1 \f4_reg[19]  ( .D(n858), .CK(clk), .Q(f4[19]), .QN(n117) );
  DFF_X1 \f5_reg[24]  ( .D(n831), .CK(clk), .Q(f5[24]), .QN(n144) );
  DFF_X1 \f5_reg[23]  ( .D(n830), .CK(clk), .Q(f5[23]), .QN(n145) );
  DFF_X1 \f5_reg[22]  ( .D(n829), .CK(clk), .Q(n615), .QN(n146) );
  DFF_X1 \f5_reg[21]  ( .D(n828), .CK(clk), .Q(f5[21]), .QN(n147) );
  DFF_X1 \f5_reg[20]  ( .D(n827), .CK(clk), .Q(f5[20]), .QN(n148) );
  DFF_X1 \f5_reg[19]  ( .D(n826), .CK(clk), .Q(f5[19]), .QN(n149) );
  DFF_X1 \f5_reg[18]  ( .D(n825), .CK(clk), .Q(f5[18]), .QN(n150) );
  DFF_X1 \f5_reg[17]  ( .D(n824), .CK(clk), .Q(f5[17]), .QN(n151) );
  DFF_X1 \f6_reg[25]  ( .D(n800), .CK(clk), .Q(n1036) );
  DFF_X1 \f6_reg[24]  ( .D(n799), .CK(clk), .Q(f6[24]) );
  DFF_X1 \f6_reg[23]  ( .D(n798), .CK(clk), .Q(f6[23]) );
  DFF_X1 \f6_reg[22]  ( .D(n797), .CK(clk), .Q(f6[22]) );
  DFF_X1 \f6_reg[21]  ( .D(n796), .CK(clk), .Q(f6[21]) );
  DFF_X1 \f6_reg[20]  ( .D(n795), .CK(clk), .Q(f6[20]) );
  DFF_X1 \f6_reg[19]  ( .D(n794), .CK(clk), .Q(f6[19]), .QN(n181) );
  DFF_X1 \f6_reg[18]  ( .D(n793), .CK(clk), .Q(f6[18]), .QN(n182) );
  DFF_X1 \f6_reg[17]  ( .D(n792), .CK(clk), .Q(f6[17]), .QN(n183) );
  DFF_X1 \f7_reg[24]  ( .D(n767), .CK(clk), .Q(n1032) );
  DFF_X1 \f7_reg[23]  ( .D(n766), .CK(clk), .Q(n1029) );
  DFF_X1 \f7_reg[22]  ( .D(n765), .CK(clk), .Q(n1025) );
  DFF_X1 \f7_reg[21]  ( .D(n764), .CK(clk), .Q(n1021) );
  DFF_X1 \f7_reg[20]  ( .D(n763), .CK(clk), .Q(n1017) );
  DFF_X1 \f7_reg[19]  ( .D(n762), .CK(clk), .Q(n477), .QN(n213) );
  DFF_X1 \f7_reg[18]  ( .D(n761), .CK(clk), .Q(n479), .QN(n214) );
  DFF_X1 \f_reg[31]  ( .D(n679), .CK(clk), .Q(f[31]), .QN(n37) );
  DFF_X1 \f_reg[30]  ( .D(n680), .CK(clk), .Q(f[30]), .QN(n36) );
  DFF_X1 \f_reg[29]  ( .D(n681), .CK(clk), .Q(f[29]), .QN(n35) );
  DFF_X1 \f8_reg[28]  ( .D(n739), .CK(clk), .Q(f8[28]), .QN(n236) );
  DFF_X1 \f_reg[28]  ( .D(n682), .CK(clk), .Q(f[28]), .QN(n34) );
  DFF_X1 \f_reg[27]  ( .D(n683), .CK(clk), .Q(f[27]), .QN(n33) );
  DFF_X1 \f_reg[26]  ( .D(n684), .CK(clk), .Q(f[26]), .QN(n32) );
  DFF_X1 \f8_reg[25]  ( .D(n736), .CK(clk), .Q(f8[25]), .QN(n239) );
  DFF_X1 \f_reg[25]  ( .D(n685), .CK(clk), .Q(f[25]), .QN(n20) );
  DFF_X1 \f_reg[24]  ( .D(n686), .CK(clk), .Q(f[24]), .QN(n19) );
  DFF_X1 \f8_reg[23]  ( .D(n734), .CK(clk), .Q(f8[23]), .QN(n241) );
  DFF_X1 \f_reg[23]  ( .D(n687), .CK(clk), .Q(f[23]), .QN(n18) );
  DFF_X1 \f8_reg[22]  ( .D(n733), .CK(clk), .Q(f8[22]), .QN(n242) );
  DFF_X1 \f_reg[22]  ( .D(n688), .CK(clk), .Q(f[22]), .QN(n17) );
  DFF_X1 \f8_reg[21]  ( .D(n732), .CK(clk), .Q(f8[21]), .QN(n243) );
  DFF_X1 \f_reg[21]  ( .D(n689), .CK(clk), .Q(f[21]), .QN(n15) );
  DFF_X1 \f8_reg[20]  ( .D(n731), .CK(clk), .Q(f8[20]), .QN(n244) );
  DFF_X1 \f_reg[20]  ( .D(n690), .CK(clk), .Q(f[20]), .QN(n14) );
  DFF_X1 \f8_reg[19]  ( .D(n730), .CK(clk), .Q(f8[19]), .QN(n245) );
  DFF_X1 \f_reg[19]  ( .D(n691), .CK(clk), .Q(f[19]) );
  DFF_X1 \f8_reg[18]  ( .D(n729), .CK(clk), .Q(f8[18]), .QN(n246) );
  DFF_X1 \f_reg[18]  ( .D(n692), .CK(clk), .Q(f[18]) );
  DFF_X1 \f8_reg[17]  ( .D(n728), .CK(clk), .Q(f8[17]), .QN(n247) );
  DFF_X1 \f_reg[17]  ( .D(n693), .CK(clk), .Q(f[17]) );
  DFF_X1 \f8_reg[16]  ( .D(n727), .CK(clk), .Q(f8[16]), .QN(n248) );
  DFF_X1 \f_reg[16]  ( .D(n694), .CK(clk), .Q(f[16]) );
  DFF_X1 \f_reg[15]  ( .D(n695), .CK(clk), .Q(f[15]) );
  DFF_X1 \f_reg[14]  ( .D(n696), .CK(clk), .Q(f[14]) );
  DFF_X1 \f_reg[13]  ( .D(n697), .CK(clk), .Q(f[13]) );
  DFF_X1 \f_reg[12]  ( .D(n698), .CK(clk), .Q(f[12]) );
  DFF_X1 \f_reg[11]  ( .D(n699), .CK(clk), .Q(f[11]) );
  DFF_X1 \f_reg[10]  ( .D(n700), .CK(clk), .Q(f[10]) );
  DFF_X1 \f_reg[9]  ( .D(n701), .CK(clk), .Q(f[9]) );
  DFF_X1 \f_reg[8]  ( .D(n702), .CK(clk), .Q(f[8]), .QN(n38) );
  DFF_X1 \f_reg[7]  ( .D(n703), .CK(clk), .Q(f[7]), .QN(n39) );
  DFF_X1 \f_reg[6]  ( .D(n704), .CK(clk), .Q(f[6]), .QN(n40) );
  DFF_X1 \f_reg[5]  ( .D(n705), .CK(clk), .Q(f[5]), .QN(n96) );
  DFF_X1 \f_reg[4]  ( .D(n706), .CK(clk), .Q(f[4]), .QN(n97) );
  DFF_X1 \f_reg[3]  ( .D(n707), .CK(clk), .Q(f[3]), .QN(n98) );
  DFF_X1 \f_reg[2]  ( .D(n708), .CK(clk), .Q(f[2]), .QN(n99) );
  DFF_X1 \f_reg[1]  ( .D(n709), .CK(clk), .Q(f[1]), .QN(n100) );
  DFF_X1 \f_reg[0]  ( .D(n710), .CK(clk), .Q(f[0]), .QN(n101) );
  memory_WIDTH16_SIZE8_LOGSIZE3_0 mem_x ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_x), .addr(addr_x), .wr_en(wr_en_x) );
  memory_WIDTH16_SIZE8_LOGSIZE3_8 mem_a1 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a1), .addr(addr_a1), .wr_en(wr_en_a1) );
  memory_WIDTH16_SIZE8_LOGSIZE3_7 mem_a2 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a2), .addr(addr_a2), .wr_en(wr_en_a2) );
  memory_WIDTH16_SIZE8_LOGSIZE3_6 mem_a3 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a3), .addr(addr_a3), .wr_en(wr_en_a3) );
  memory_WIDTH16_SIZE8_LOGSIZE3_5 mem_a4 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a4), .addr(addr_a4), .wr_en(wr_en_a4) );
  memory_WIDTH16_SIZE8_LOGSIZE3_4 mem_a5 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a5), .addr(addr_a5), .wr_en(wr_en_a5) );
  memory_WIDTH16_SIZE8_LOGSIZE3_3 mem_a6 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a6), .addr(addr_a6), .wr_en(wr_en_a6) );
  memory_WIDTH16_SIZE8_LOGSIZE3_2 mem_a7 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a7), .addr(addr_a7), .wr_en(wr_en_a7) );
  memory_WIDTH16_SIZE8_LOGSIZE3_1 mem_a8 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a8), .addr(addr_a8), .wr_en(wr_en_a8) );
  memory_WIDTH32_SIZE8_LOGSIZE3 mem_y ( .clk(clk), .data_in(f), .data_out(
        data_out), .addr(addr_y), .wr_en(wr_en_y) );
  datapath_DW_mult_tc_8 mult_84 ( .a(data_out_a1), .b({data_out_x[15], n203, 
        data_out_x[13], n2, data_out_x[11], n202, n171, n169, data_out_x[7], 
        n201, n204, data_out_x[4:0]}), .product({\mul_out1[31] , 
        \mul_out1[30] , \mul_out1[29] , \mul_out1[28] , \mul_out1[27] , 
        \mul_out1[26] , \mul_out1[25] , \mul_out1[24] , \mul_out1[23] , 
        \mul_out1[22] , \mul_out1[21] , \mul_out1[20] , \mul_out1[19] , 
        \mul_out1[18] , \mul_out1[17] , \mul_out1[16] , \mul_out1[15] , 
        \mul_out1[14] , \mul_out1[13] , \mul_out1[12] , \mul_out1[11] , 
        \mul_out1[10] , \mul_out1[9] , \mul_out1[8] , \mul_out1[7] , 
        \mul_out1[6] , \mul_out1[5] , \mul_out1[4] , \mul_out1[3] , 
        \mul_out1[2] , \mul_out1[1] , \mul_out1[0] }) );
  datapath_DW_mult_tc_9 mult_86 ( .a(data_out_a2), .b({data_out_x[15], n203, 
        data_out_x[13:11], n202, data_out_x[9:7], n179, data_out_x[5:0]}), 
        .product({\mul_out2[31] , \mul_out2[30] , \mul_out2[29] , 
        \mul_out2[28] , \mul_out2[27] , \mul_out2[26] , \mul_out2[25] , 
        \mul_out2[24] , \mul_out2[23] , \mul_out2[22] , \mul_out2[21] , 
        \mul_out2[20] , \mul_out2[19] , \mul_out2[18] , \mul_out2[17] , 
        \mul_out2[16] , \mul_out2[15] , \mul_out2[14] , \mul_out2[13] , 
        \mul_out2[12] , \mul_out2[11] , \mul_out2[10] , \mul_out2[9] , 
        \mul_out2[8] , \mul_out2[7] , \mul_out2[6] , \mul_out2[5] , 
        \mul_out2[4] , \mul_out2[3] , \mul_out2[2] , \mul_out2[1] , 
        \mul_out2[0] }) );
  datapath_DW_mult_tc_10 mult_88 ( .a(data_out_a3), .b({data_out_x[15], n203, 
        data_out_x[13], n3, data_out_x[11], n202, n172, n170, data_out_x[7], 
        n179, n204, data_out_x[4:0]}), .product({\mul_out3[31] , 
        \mul_out3[30] , \mul_out3[29] , \mul_out3[28] , \mul_out3[27] , 
        \mul_out3[26] , \mul_out3[25] , \mul_out3[24] , \mul_out3[23] , 
        \mul_out3[22] , \mul_out3[21] , \mul_out3[20] , \mul_out3[19] , 
        \mul_out3[18] , \mul_out3[17] , \mul_out3[16] , \mul_out3[15] , 
        \mul_out3[14] , \mul_out3[13] , \mul_out3[12] , \mul_out3[11] , 
        \mul_out3[10] , \mul_out3[9] , \mul_out3[8] , \mul_out3[7] , 
        \mul_out3[6] , \mul_out3[5] , \mul_out3[4] , \mul_out3[3] , 
        \mul_out3[2] , \mul_out3[1] , \mul_out3[0] }) );
  datapath_DW_mult_tc_11 mult_90 ( .a(data_out_a4), .b({data_out_x[15], n203, 
        data_out_x[13], n2, data_out_x[11], n202, n172, n169, data_out_x[7], 
        n180, n204, data_out_x[4:0]}), .product({\mul_out4[31] , 
        \mul_out4[30] , \mul_out4[29] , \mul_out4[28] , \mul_out4[27] , 
        \mul_out4[26] , \mul_out4[25] , \mul_out4[24] , \mul_out4[23] , 
        \mul_out4[22] , \mul_out4[21] , \mul_out4[20] , \mul_out4[19] , 
        \mul_out4[18] , \mul_out4[17] , \mul_out4[16] , \mul_out4[15] , 
        \mul_out4[14] , \mul_out4[13] , \mul_out4[12] , \mul_out4[11] , 
        \mul_out4[10] , \mul_out4[9] , \mul_out4[8] , \mul_out4[7] , 
        \mul_out4[6] , \mul_out4[5] , \mul_out4[4] , \mul_out4[3] , 
        \mul_out4[2] , \mul_out4[1] , \mul_out4[0] }) );
  datapath_DW_mult_tc_12 mult_92 ( .a(data_out_a5), .b({data_out_x[15:11], 
        n202, data_out_x[9:7], n201, n204, data_out_x[4:0]}), .product({
        \mul_out5[31] , \mul_out5[30] , \mul_out5[29] , \mul_out5[28] , 
        \mul_out5[27] , \mul_out5[26] , \mul_out5[25] , \mul_out5[24] , 
        \mul_out5[23] , \mul_out5[22] , \mul_out5[21] , \mul_out5[20] , 
        \mul_out5[19] , \mul_out5[18] , \mul_out5[17] , \mul_out5[16] , 
        \mul_out5[15] , \mul_out5[14] , \mul_out5[13] , \mul_out5[12] , 
        \mul_out5[11] , \mul_out5[10] , \mul_out5[9] , \mul_out5[8] , 
        \mul_out5[7] , \mul_out5[6] , \mul_out5[5] , \mul_out5[4] , 
        \mul_out5[3] , \mul_out5[2] , \mul_out5[1] , \mul_out5[0] }) );
  datapath_DW_mult_tc_13 mult_94 ( .a(data_out_a6), .b({data_out_x[15], n203, 
        data_out_x[13], n2, data_out_x[11], n202, n205, data_out_x[8:7], n201, 
        n204, data_out_x[4:0]}), .product({\mul_out6[31] , \mul_out6[30] , 
        \mul_out6[29] , \mul_out6[28] , \mul_out6[27] , \mul_out6[26] , 
        \mul_out6[25] , \mul_out6[24] , \mul_out6[23] , \mul_out6[22] , 
        \mul_out6[21] , \mul_out6[20] , \mul_out6[19] , \mul_out6[18] , 
        \mul_out6[17] , \mul_out6[16] , \mul_out6[15] , \mul_out6[14] , 
        \mul_out6[13] , \mul_out6[12] , \mul_out6[11] , \mul_out6[10] , 
        \mul_out6[9] , \mul_out6[8] , \mul_out6[7] , \mul_out6[6] , 
        \mul_out6[5] , \mul_out6[4] , \mul_out6[3] , \mul_out6[2] , 
        \mul_out6[1] , \mul_out6[0] }) );
  datapath_DW_mult_tc_14 mult_96 ( .a(data_out_a7), .b({data_out_x[15], n203, 
        data_out_x[13], n3, data_out_x[11], n202, n205, n170, data_out_x[7], 
        n179, n204, data_out_x[4:0]}), .product({\mul_out7[31] , 
        \mul_out7[30] , \mul_out7[29] , \mul_out7[28] , \mul_out7[27] , 
        \mul_out7[26] , \mul_out7[25] , \mul_out7[24] , \mul_out7[23] , 
        \mul_out7[22] , \mul_out7[21] , \mul_out7[20] , \mul_out7[19] , 
        \mul_out7[18] , \mul_out7[17] , \mul_out7[16] , \mul_out7[15] , 
        \mul_out7[14] , \mul_out7[13] , \mul_out7[12] , \mul_out7[11] , 
        \mul_out7[10] , \mul_out7[9] , \mul_out7[8] , \mul_out7[7] , 
        \mul_out7[6] , \mul_out7[5] , \mul_out7[4] , \mul_out7[3] , 
        \mul_out7[2] , \mul_out7[1] , \mul_out7[0] }) );
  datapath_DW_mult_tc_15 mult_98 ( .a(data_out_a8), .b({data_out_x[15], n203, 
        data_out_x[13], n3, data_out_x[11], n202, n171, n169, data_out_x[7], 
        n180, n204, data_out_x[4:0]}), .product({\mul_out8[31] , 
        \mul_out8[30] , \mul_out8[29] , \mul_out8[28] , \mul_out8[27] , 
        \mul_out8[26] , \mul_out8[25] , \mul_out8[24] , \mul_out8[23] , 
        \mul_out8[22] , \mul_out8[21] , \mul_out8[20] , \mul_out8[19] , 
        \mul_out8[18] , \mul_out8[17] , \mul_out8[16] , \mul_out8[15] , 
        \mul_out8[14] , \mul_out8[13] , \mul_out8[12] , \mul_out8[11] , 
        \mul_out8[10] , \mul_out8[9] , \mul_out8[8] , \mul_out8[7] , 
        \mul_out8[6] , \mul_out8[5] , \mul_out8[4] , \mul_out8[3] , 
        \mul_out8[2] , \mul_out8[1] , \mul_out8[0] }) );
  datapath_DW01_add_8 add_85 ( .A(f1), .B({\mul_out1[31] , \mul_out1[30] , 
        \mul_out1[29] , \mul_out1[28] , \mul_out1[27] , \mul_out1[26] , 
        \mul_out1[25] , \mul_out1[24] , \mul_out1[23] , \mul_out1[22] , 
        \mul_out1[21] , \mul_out1[20] , \mul_out1[19] , \mul_out1[18] , 
        \mul_out1[17] , \mul_out1[16] , \mul_out1[15] , \mul_out1[14] , 
        \mul_out1[13] , \mul_out1[12] , \mul_out1[11] , \mul_out1[10] , 
        \mul_out1[9] , \mul_out1[8] , \mul_out1[7] , \mul_out1[6] , 
        \mul_out1[5] , \mul_out1[4] , \mul_out1[3] , \mul_out1[2] , 
        \mul_out1[1] , \mul_out1[0] }), .CI(1'b0), .SUM(add_r1) );
  datapath_DW01_add_9 add_87 ( .A({f2[31:28], n643, n645, n647, f2[24], n650, 
        n652, n654, n656, n658, n660, n662, f2[16:0]}), .B({\mul_out2[31] , 
        \mul_out2[30] , \mul_out2[29] , \mul_out2[28] , \mul_out2[27] , 
        \mul_out2[26] , \mul_out2[25] , \mul_out2[24] , \mul_out2[23] , 
        \mul_out2[22] , \mul_out2[21] , \mul_out2[20] , \mul_out2[19] , 
        \mul_out2[18] , \mul_out2[17] , \mul_out2[16] , \mul_out2[15] , 
        \mul_out2[14] , \mul_out2[13] , \mul_out2[12] , \mul_out2[11] , 
        \mul_out2[10] , \mul_out2[9] , \mul_out2[8] , \mul_out2[7] , 
        \mul_out2[6] , \mul_out2[5] , \mul_out2[4] , \mul_out2[3] , 
        \mul_out2[2] , \mul_out2[1] , \mul_out2[0] }), .CI(1'b0), .SUM(add_r2)
         );
  datapath_DW01_add_10 add_89 ( .A({n563, n565, n567, n569, n571, n573, n575, 
        n577, n579, n581, f3[21:0]}), .B({\mul_out3[31] , \mul_out3[30] , 
        \mul_out3[29] , \mul_out3[28] , \mul_out3[27] , \mul_out3[26] , 
        \mul_out3[25] , \mul_out3[24] , \mul_out3[23] , \mul_out3[22] , 
        \mul_out3[21] , \mul_out3[20] , \mul_out3[19] , \mul_out3[18] , 
        \mul_out3[17] , \mul_out3[16] , \mul_out3[15] , \mul_out3[14] , 
        \mul_out3[13] , \mul_out3[12] , \mul_out3[11] , \mul_out3[10] , 
        \mul_out3[9] , \mul_out3[8] , \mul_out3[7] , \mul_out3[6] , 
        \mul_out3[5] , \mul_out3[4] , \mul_out3[3] , \mul_out3[2] , 
        \mul_out3[1] , \mul_out3[0] }), .CI(1'b0), .SUM(add_r3) );
  datapath_DW01_add_12 add_93 ( .A({f5[31:27], n610, f5[25:23], n615, f5[21:0]}), .B({\mul_out5[31] , \mul_out5[30] , \mul_out5[29] , \mul_out5[28] , 
        \mul_out5[27] , \mul_out5[26] , \mul_out5[25] , \mul_out5[24] , 
        \mul_out5[23] , \mul_out5[22] , \mul_out5[21] , \mul_out5[20] , 
        \mul_out5[19] , \mul_out5[18] , \mul_out5[17] , \mul_out5[16] , 
        \mul_out5[15] , \mul_out5[14] , \mul_out5[13] , \mul_out5[12] , 
        \mul_out5[11] , \mul_out5[10] , \mul_out5[9] , \mul_out5[8] , 
        \mul_out5[7] , \mul_out5[6] , \mul_out5[5] , \mul_out5[4] , 
        \mul_out5[3] , \mul_out5[2] , \mul_out5[1] , \mul_out5[0] }), .CI(1'b0), .SUM(add_r5) );
  datapath_DW01_add_13 add_95 ( .A({n1064, n1056, n1052, n1048, n1044, n1040, 
        n1036, f6[24:0]}), .B({\mul_out6[31] , \mul_out6[30] , \mul_out6[29] , 
        \mul_out6[28] , \mul_out6[27] , \mul_out6[26] , \mul_out6[25] , 
        \mul_out6[24] , \mul_out6[23] , \mul_out6[22] , \mul_out6[21] , 
        \mul_out6[20] , \mul_out6[19] , \mul_out6[18] , \mul_out6[17] , 
        \mul_out6[16] , \mul_out6[15] , \mul_out6[14] , \mul_out6[13] , 
        \mul_out6[12] , \mul_out6[11] , \mul_out6[10] , \mul_out6[9] , 
        \mul_out6[8] , \mul_out6[7] , \mul_out6[6] , \mul_out6[5] , 
        \mul_out6[4] , \mul_out6[3] , \mul_out6[2] , \mul_out6[1] , 
        \mul_out6[0] }), .CI(1'b0), .SUM(add_r6) );
  datapath_DW01_add_14 add_97 ( .A({f7[31:25], n1032, n1029, n1025, n1021, 
        n1017, n477, n479, f7[17:0]}), .B({\mul_out7[31] , \mul_out7[30] , 
        \mul_out7[29] , \mul_out7[28] , \mul_out7[27] , \mul_out7[26] , 
        \mul_out7[25] , \mul_out7[24] , \mul_out7[23] , \mul_out7[22] , 
        \mul_out7[21] , \mul_out7[20] , \mul_out7[19] , \mul_out7[18] , 
        \mul_out7[17] , \mul_out7[16] , \mul_out7[15] , \mul_out7[14] , 
        \mul_out7[13] , \mul_out7[12] , \mul_out7[11] , \mul_out7[10] , 
        \mul_out7[9] , \mul_out7[8] , \mul_out7[7] , \mul_out7[6] , 
        \mul_out7[5] , \mul_out7[4] , \mul_out7[3] , \mul_out7[2] , 
        \mul_out7[1] , \mul_out7[0] }), .CI(1'b0), .SUM(add_r7) );
  datapath_DW01_add_15 add_99 ( .A(f8), .B({\mul_out8[31] , \mul_out8[30] , 
        \mul_out8[29] , \mul_out8[28] , \mul_out8[27] , \mul_out8[26] , 
        \mul_out8[25] , \mul_out8[24] , \mul_out8[23] , \mul_out8[22] , 
        \mul_out8[21] , \mul_out8[20] , \mul_out8[19] , \mul_out8[18] , 
        \mul_out8[17] , \mul_out8[16] , \mul_out8[15] , \mul_out8[14] , 
        \mul_out8[13] , \mul_out8[12] , \mul_out8[11] , \mul_out8[10] , 
        \mul_out8[9] , \mul_out8[8] , \mul_out8[7] , \mul_out8[6] , 
        \mul_out8[5] , \mul_out8[4] , \mul_out8[3] , \mul_out8[2] , 
        \mul_out8[1] , \mul_out8[0] }), .CI(1'b0), .SUM(add_r8) );
  datapath_DW01_add_16 add_91 ( .A(f4), .B({\mul_out4[31] , \mul_out4[30] , 
        \mul_out4[29] , \mul_out4[28] , \mul_out4[27] , \mul_out4[26] , 
        \mul_out4[25] , \mul_out4[24] , \mul_out4[23] , \mul_out4[22] , 
        \mul_out4[21] , \mul_out4[20] , \mul_out4[19] , \mul_out4[18] , 
        \mul_out4[17] , \mul_out4[16] , \mul_out4[15] , \mul_out4[14] , 
        \mul_out4[13] , \mul_out4[12] , \mul_out4[11] , \mul_out4[10] , 
        \mul_out4[9] , \mul_out4[8] , \mul_out4[7] , \mul_out4[6] , 
        \mul_out4[5] , \mul_out4[4] , \mul_out4[3] , \mul_out4[2] , 
        \mul_out4[1] , \mul_out4[0] }), .CI(1'b0), .SUM(add_r4) );
  DFF_X1 \f1_reg[24]  ( .D(n959), .CK(clk), .Q(f1[24]), .QN(n16) );
  DFF_X1 \f4_reg[28]  ( .D(n867), .CK(clk), .Q(f4[28]), .QN(n108) );
  DFF_X1 \f6_reg[3]  ( .D(n778), .CK(clk), .Q(f6[3]), .QN(n197) );
  DFF_X1 \f6_reg[2]  ( .D(n777), .CK(clk), .Q(f6[2]), .QN(n198) );
  DFF_X1 \f6_reg[1]  ( .D(n776), .CK(clk), .Q(f6[1]), .QN(n199) );
  DFF_X1 \f6_reg[0]  ( .D(n775), .CK(clk), .Q(f6[0]), .QN(n200) );
  DFF_X1 \f4_reg[3]  ( .D(n842), .CK(clk), .Q(f4[3]), .QN(n133) );
  DFF_X1 \f4_reg[2]  ( .D(n841), .CK(clk), .Q(f4[2]), .QN(n134) );
  DFF_X1 \f4_reg[1]  ( .D(n840), .CK(clk), .Q(f4[1]), .QN(n135) );
  DFF_X1 \f4_reg[0]  ( .D(n839), .CK(clk), .Q(f4[0]), .QN(n136) );
  DFF_X1 \f8_reg[0]  ( .D(n711), .CK(clk), .Q(f8[0]), .QN(n264) );
  DFF_X1 \f8_reg[3]  ( .D(n714), .CK(clk), .Q(f8[3]), .QN(n261) );
  DFF_X1 \f8_reg[2]  ( .D(n713), .CK(clk), .Q(f8[2]), .QN(n262) );
  DFF_X1 \f8_reg[1]  ( .D(n712), .CK(clk), .Q(f8[1]), .QN(n263) );
  DFF_X1 \f1_reg[3]  ( .D(n938), .CK(clk), .Q(f1[3]), .QN(n995) );
  DFF_X1 \f1_reg[2]  ( .D(n937), .CK(clk), .Q(f1[2]), .QN(n1000) );
  DFF_X1 \f1_reg[1]  ( .D(n936), .CK(clk), .Q(f1[1]), .QN(n1005) );
  DFF_X1 \f1_reg[0]  ( .D(n935), .CK(clk), .Q(f1[0]), .QN(n1010) );
  DFF_X1 \f2_reg[2]  ( .D(n905), .CK(clk), .Q(f2[2]), .QN(n70) );
  DFF_X1 \f2_reg[1]  ( .D(n904), .CK(clk), .Q(f2[1]), .QN(n71) );
  DFF_X1 \f2_reg[0]  ( .D(n903), .CK(clk), .Q(f2[0]), .QN(n72) );
  DFF_X1 \f7_reg[3]  ( .D(n746), .CK(clk), .Q(f7[3]) );
  DFF_X1 \f7_reg[2]  ( .D(n745), .CK(clk), .Q(f7[2]) );
  DFF_X1 \f7_reg[1]  ( .D(n744), .CK(clk), .Q(f7[1]) );
  DFF_X1 \f7_reg[0]  ( .D(n743), .CK(clk), .Q(f7[0]) );
  DFF_X1 \f5_reg[3]  ( .D(n810), .CK(clk), .Q(f5[3]), .QN(n165) );
  DFF_X1 \f5_reg[2]  ( .D(n809), .CK(clk), .Q(f5[2]), .QN(n166) );
  DFF_X1 \f5_reg[1]  ( .D(n808), .CK(clk), .Q(f5[1]), .QN(n167) );
  DFF_X1 \f5_reg[0]  ( .D(n807), .CK(clk), .Q(f5[0]), .QN(n168) );
  DFF_X1 \f3_reg[3]  ( .D(n874), .CK(clk), .Q(f3[3]) );
  DFF_X1 \f3_reg[2]  ( .D(n873), .CK(clk), .Q(f3[2]) );
  DFF_X1 \f3_reg[1]  ( .D(n872), .CK(clk), .Q(f3[1]) );
  DFF_X1 \f3_reg[0]  ( .D(n871), .CK(clk), .Q(f3[0]) );
  DFF_X1 \f2_reg[3]  ( .D(n906), .CK(clk), .Q(f2[3]), .QN(n69) );
  DFF_X1 \f4_reg[4]  ( .D(n843), .CK(clk), .Q(f4[4]), .QN(n132) );
  DFF_X1 \f8_reg[4]  ( .D(n715), .CK(clk), .Q(f8[4]), .QN(n260) );
  DFF_X1 \f1_reg[4]  ( .D(n939), .CK(clk), .Q(f1[4]), .QN(n990) );
  DFF_X1 \f3_reg[4]  ( .D(n875), .CK(clk), .Q(f3[4]) );
  DFF_X1 \f6_reg[4]  ( .D(n779), .CK(clk), .Q(f6[4]), .QN(n196) );
  DFF_X1 \f5_reg[4]  ( .D(n811), .CK(clk), .Q(f5[4]), .QN(n164) );
  DFF_X1 \f7_reg[4]  ( .D(n747), .CK(clk), .Q(f7[4]) );
  DFF_X1 \f2_reg[4]  ( .D(n907), .CK(clk), .Q(f2[4]), .QN(n68) );
  DFF_X1 \f4_reg[5]  ( .D(n844), .CK(clk), .Q(f4[5]), .QN(n131) );
  DFF_X1 \f8_reg[5]  ( .D(n716), .CK(clk), .Q(f8[5]), .QN(n259) );
  DFF_X1 \f6_reg[5]  ( .D(n780), .CK(clk), .Q(f6[5]), .QN(n195) );
  DFF_X1 \f3_reg[5]  ( .D(n876), .CK(clk), .Q(f3[5]) );
  DFF_X1 \f5_reg[5]  ( .D(n812), .CK(clk), .Q(f5[5]), .QN(n163) );
  DFF_X1 \f1_reg[5]  ( .D(n940), .CK(clk), .Q(f1[5]), .QN(n985) );
  DFF_X1 \f2_reg[5]  ( .D(n908), .CK(clk), .Q(f2[5]), .QN(n67) );
  DFF_X1 \f7_reg[5]  ( .D(n748), .CK(clk), .Q(f7[5]) );
  DFF_X1 \f4_reg[6]  ( .D(n845), .CK(clk), .Q(f4[6]), .QN(n130) );
  DFF_X1 \f8_reg[6]  ( .D(n717), .CK(clk), .Q(f8[6]), .QN(n258) );
  DFF_X1 \f8_reg[7]  ( .D(n718), .CK(clk), .Q(f8[7]), .QN(n257) );
  DFF_X1 \f1_reg[6]  ( .D(n941), .CK(clk), .Q(f1[6]), .QN(n980) );
  DFF_X1 \f6_reg[6]  ( .D(n781), .CK(clk), .Q(f6[6]), .QN(n194) );
  DFF_X1 \f5_reg[6]  ( .D(n813), .CK(clk), .Q(f5[6]), .QN(n162) );
  DFF_X1 \f6_reg[7]  ( .D(n782), .CK(clk), .Q(f6[7]), .QN(n193) );
  DFF_X1 \f3_reg[6]  ( .D(n877), .CK(clk), .Q(f3[6]) );
  DFF_X1 \f5_reg[7]  ( .D(n814), .CK(clk), .Q(f5[7]), .QN(n161) );
  DFF_X1 \f3_reg[7]  ( .D(n878), .CK(clk), .Q(f3[7]) );
  DFF_X1 \f2_reg[6]  ( .D(n909), .CK(clk), .Q(f2[6]), .QN(n66) );
  DFF_X1 \f2_reg[7]  ( .D(n910), .CK(clk), .Q(f2[7]), .QN(n65) );
  DFF_X1 \f7_reg[6]  ( .D(n749), .CK(clk), .Q(f7[6]) );
  DFF_X1 \f1_reg[7]  ( .D(n942), .CK(clk), .Q(f1[7]), .QN(n975) );
  DFF_X1 \f7_reg[7]  ( .D(n750), .CK(clk), .Q(f7[7]) );
  DFF_X1 \f4_reg[7]  ( .D(n846), .CK(clk), .Q(f4[7]), .QN(n129) );
  DFF_X1 \f4_reg[8]  ( .D(n847), .CK(clk), .Q(f4[8]), .QN(n128) );
  DFF_X1 \f4_reg[9]  ( .D(n848), .CK(clk), .Q(f4[9]), .QN(n127) );
  DFF_X1 \f6_reg[8]  ( .D(n783), .CK(clk), .Q(f6[8]), .QN(n192) );
  DFF_X1 \f4_reg[10]  ( .D(n849), .CK(clk), .Q(f4[10]), .QN(n126) );
  DFF_X1 \f8_reg[8]  ( .D(n719), .CK(clk), .Q(f8[8]), .QN(n256) );
  DFF_X1 \f5_reg[8]  ( .D(n815), .CK(clk), .Q(f5[8]), .QN(n160) );
  DFF_X1 \f3_reg[8]  ( .D(n879), .CK(clk), .Q(f3[8]) );
  DFF_X1 \f2_reg[8]  ( .D(n911), .CK(clk), .Q(f2[8]), .QN(n64) );
  DFF_X1 \f7_reg[8]  ( .D(n751), .CK(clk), .Q(f7[8]) );
  DFF_X1 \f8_reg[9]  ( .D(n720), .CK(clk), .Q(f8[9]), .QN(n255) );
  DFF_X1 \f6_reg[9]  ( .D(n784), .CK(clk), .Q(f6[9]), .QN(n191) );
  DFF_X1 \f8_reg[10]  ( .D(n721), .CK(clk), .Q(f8[10]), .QN(n254) );
  DFF_X1 \f1_reg[8]  ( .D(n943), .CK(clk), .Q(f1[8]), .QN(n970) );
  DFF_X1 \f5_reg[9]  ( .D(n816), .CK(clk), .Q(f5[9]), .QN(n159) );
  DFF_X1 \f3_reg[9]  ( .D(n880), .CK(clk), .Q(f3[9]), .QN(n95) );
  DFF_X1 \f2_reg[10]  ( .D(n913), .CK(clk), .Q(f2[10]), .QN(n62) );
  DFF_X1 \f2_reg[9]  ( .D(n912), .CK(clk), .Q(f2[9]), .QN(n63) );
  DFF_X1 \f7_reg[9]  ( .D(n752), .CK(clk), .Q(f7[9]), .QN(n223) );
  DFF_X1 \f1_reg[10]  ( .D(n945), .CK(clk), .Q(f1[10]), .QN(n30) );
  DFF_X1 \f1_reg[9]  ( .D(n944), .CK(clk), .Q(f1[9]), .QN(n31) );
  DFF_X1 \f8_reg[11]  ( .D(n722), .CK(clk), .Q(f8[11]), .QN(n253) );
  DFF_X1 \f6_reg[10]  ( .D(n785), .CK(clk), .Q(f6[10]), .QN(n190) );
  DFF_X1 \f4_reg[11]  ( .D(n850), .CK(clk), .Q(f4[11]), .QN(n125) );
  DFF_X1 \f1_reg[11]  ( .D(n946), .CK(clk), .Q(f1[11]), .QN(n29) );
  DFF_X1 \f7_reg[10]  ( .D(n753), .CK(clk), .Q(f7[10]), .QN(n222) );
  DFF_X1 \f6_reg[11]  ( .D(n786), .CK(clk), .Q(f6[11]), .QN(n189) );
  DFF_X1 \f2_reg[11]  ( .D(n914), .CK(clk), .Q(f2[11]), .QN(n61) );
  DFF_X1 \f5_reg[10]  ( .D(n817), .CK(clk), .Q(f5[10]), .QN(n158) );
  DFF_X1 \f3_reg[10]  ( .D(n881), .CK(clk), .Q(f3[10]), .QN(n94) );
  DFF_X1 \f7_reg[11]  ( .D(n754), .CK(clk), .Q(f7[11]), .QN(n221) );
  DFF_X1 \f5_reg[11]  ( .D(n818), .CK(clk), .Q(f5[11]), .QN(n157) );
  DFF_X1 \f3_reg[11]  ( .D(n882), .CK(clk), .Q(f3[11]), .QN(n93) );
  DFF_X1 \f4_reg[12]  ( .D(n851), .CK(clk), .Q(f4[12]), .QN(n124) );
  DFF_X1 \f4_reg[13]  ( .D(n852), .CK(clk), .Q(f4[13]), .QN(n123) );
  DFF_X1 \f4_reg[14]  ( .D(n853), .CK(clk), .Q(f4[14]), .QN(n122) );
  DFF_X1 \f6_reg[12]  ( .D(n787), .CK(clk), .Q(f6[12]), .QN(n188) );
  DFF_X1 \f8_reg[12]  ( .D(n723), .CK(clk), .Q(f8[12]), .QN(n252) );
  DFF_X1 \f8_reg[13]  ( .D(n724), .CK(clk), .Q(f8[13]), .QN(n251) );
  DFF_X1 \f2_reg[12]  ( .D(n915), .CK(clk), .Q(f2[12]), .QN(n60) );
  DFF_X1 \f1_reg[12]  ( .D(n947), .CK(clk), .Q(f1[12]), .QN(n28) );
  DFF_X1 \f6_reg[13]  ( .D(n788), .CK(clk), .Q(f6[13]), .QN(n187) );
  DFF_X1 \f1_reg[13]  ( .D(n948), .CK(clk), .Q(f1[13]), .QN(n27) );
  DFF_X1 \f5_reg[12]  ( .D(n819), .CK(clk), .Q(f5[12]), .QN(n156) );
  DFF_X1 \f2_reg[13]  ( .D(n916), .CK(clk), .Q(f2[13]), .QN(n59) );
  DFF_X1 \f7_reg[12]  ( .D(n755), .CK(clk), .Q(f7[12]), .QN(n220) );
  DFF_X1 \f3_reg[12]  ( .D(n883), .CK(clk), .Q(f3[12]), .QN(n92) );
  DFF_X1 \f8_reg[14]  ( .D(n725), .CK(clk), .Q(f8[14]), .QN(n250) );
  DFF_X1 \f4_reg[15]  ( .D(n854), .CK(clk), .Q(f4[15]), .QN(n121) );
  DFF_X1 \f5_reg[13]  ( .D(n820), .CK(clk), .Q(f5[13]), .QN(n155) );
  DFF_X1 \f8_reg[15]  ( .D(n726), .CK(clk), .Q(f8[15]), .QN(n249) );
  DFF_X1 \f7_reg[13]  ( .D(n756), .CK(clk), .Q(f7[13]), .QN(n219) );
  DFF_X1 \f6_reg[14]  ( .D(n789), .CK(clk), .Q(f6[14]), .QN(n186) );
  DFF_X1 \f3_reg[13]  ( .D(n884), .CK(clk), .Q(f3[13]), .QN(n91) );
  DFF_X1 \f2_reg[14]  ( .D(n917), .CK(clk), .Q(f2[14]), .QN(n58) );
  DFF_X1 \f6_reg[15]  ( .D(n790), .CK(clk), .Q(f6[15]), .QN(n185) );
  DFF_X1 \f1_reg[14]  ( .D(n949), .CK(clk), .Q(f1[14]), .QN(n26) );
  DFF_X1 \f2_reg[15]  ( .D(n918), .CK(clk), .Q(f2[15]), .QN(n57) );
  DFF_X1 \f5_reg[14]  ( .D(n821), .CK(clk), .Q(f5[14]), .QN(n154) );
  DFF_X1 \f3_reg[14]  ( .D(n885), .CK(clk), .Q(f3[14]), .QN(n90) );
  DFF_X1 \f1_reg[15]  ( .D(n950), .CK(clk), .Q(f1[15]), .QN(n25) );
  DFF_X1 \f7_reg[14]  ( .D(n757), .CK(clk), .Q(f7[14]), .QN(n218) );
  DFF_X1 \f5_reg[15]  ( .D(n822), .CK(clk), .Q(f5[15]), .QN(n153) );
  DFF_X1 \f3_reg[15]  ( .D(n886), .CK(clk), .Q(f3[15]), .QN(n89) );
  DFF_X1 \f7_reg[15]  ( .D(n758), .CK(clk), .Q(f7[15]), .QN(n217) );
  DFF_X1 \f4_reg[17]  ( .D(n856), .CK(clk), .Q(f4[17]), .QN(n119) );
  DFF_X1 \f4_reg[16]  ( .D(n855), .CK(clk), .Q(f4[16]), .QN(n120) );
  DFF_X1 \f4_reg[18]  ( .D(n857), .CK(clk), .Q(f4[18]), .QN(n118) );
  DFF_X1 \f2_reg[16]  ( .D(n919), .CK(clk), .Q(f2[16]), .QN(n56) );
  DFF_X1 \f4_reg[21]  ( .D(n860), .CK(clk), .Q(f4[21]), .QN(n115) );
  DFF_X1 \f6_reg[16]  ( .D(n791), .CK(clk), .Q(f6[16]), .QN(n184) );
  DFF_X1 \f4_reg[25]  ( .D(n864), .CK(clk), .Q(f4[25]), .QN(n111) );
  DFF_X1 \f7_reg[16]  ( .D(n759), .CK(clk), .Q(f7[16]), .QN(n216) );
  DFF_X1 \f3_reg[16]  ( .D(n887), .CK(clk), .Q(f3[16]), .QN(n88) );
  DFF_X1 \f5_reg[16]  ( .D(n823), .CK(clk), .Q(f5[16]), .QN(n152) );
  DFF_X1 \f1_reg[16]  ( .D(n951), .CK(clk), .Q(f1[16]), .QN(n24) );
  DFF_X1 \f7_reg[17]  ( .D(n760), .CK(clk), .Q(f7[17]), .QN(n215) );
  DFF_X1 \f7_reg[25]  ( .D(n768), .CK(clk), .Q(f7[25]) );
  DFF_X1 \f7_reg[28]  ( .D(n771), .CK(clk), .Q(f7[28]) );
  DFF_X1 \f7_reg[26]  ( .D(n769), .CK(clk), .Q(f7[26]) );
  DFF_X1 \f7_reg[30]  ( .D(n773), .CK(clk), .Q(f7[30]) );
  DFF_X1 \f5_reg[28]  ( .D(n835), .CK(clk), .Q(f5[28]), .QN(n140) );
  DFF_X1 \f5_reg[27]  ( .D(n834), .CK(clk), .Q(f5[27]), .QN(n141) );
  DFF_X1 \f7_reg[27]  ( .D(n770), .CK(clk), .Q(f7[27]) );
  DFF_X1 \f3_reg[31]  ( .D(n902), .CK(clk), .Q(n563), .QN(n73) );
  DFF_X1 \f3_reg[30]  ( .D(n901), .CK(clk), .Q(n565), .QN(n74) );
  DFF_X1 \f3_reg[29]  ( .D(n900), .CK(clk), .Q(n567), .QN(n75) );
  DFF_X1 \f3_reg[26]  ( .D(n897), .CK(clk), .Q(n573), .QN(n78) );
  DFF_X1 \f2_reg[31]  ( .D(n934), .CK(clk), .Q(f2[31]), .QN(n41) );
  DFF_X1 \f2_reg[30]  ( .D(n933), .CK(clk), .Q(f2[30]), .QN(n42) );
  DFF_X1 \f2_reg[29]  ( .D(n932), .CK(clk), .Q(f2[29]), .QN(n43) );
  DFF_X1 \f2_reg[27]  ( .D(n930), .CK(clk), .Q(n643), .QN(n45) );
  DFF_X1 \f5_reg[29]  ( .D(n836), .CK(clk), .Q(f5[29]), .QN(n139) );
  DFF_X1 \f2_reg[28]  ( .D(n931), .CK(clk), .Q(f2[28]), .QN(n44) );
  DFF_X1 \f2_reg[26]  ( .D(n929), .CK(clk), .Q(n645), .QN(n46) );
  DFF_X1 \f2_reg[25]  ( .D(n928), .CK(clk), .Q(n647), .QN(n47) );
  DFF_X1 \f5_reg[30]  ( .D(n837), .CK(clk), .Q(f5[30]), .QN(n138) );
  DFF_X1 \f5_reg[26]  ( .D(n833), .CK(clk), .Q(n610), .QN(n142) );
  DFF_X1 \f5_reg[25]  ( .D(n832), .CK(clk), .Q(f5[25]), .QN(n143) );
  DFF_X1 \f3_reg[28]  ( .D(n899), .CK(clk), .Q(n569), .QN(n76) );
  DFF_X1 \f3_reg[27]  ( .D(n898), .CK(clk), .Q(n571), .QN(n77) );
  DFF_X1 \f3_reg[25]  ( .D(n896), .CK(clk), .Q(n575), .QN(n79) );
  DFF_X1 \f5_reg[31]  ( .D(n838), .CK(clk), .Q(f5[31]), .QN(n137) );
  DFF_X1 \f7_reg[31]  ( .D(n774), .CK(clk), .Q(f7[31]) );
  DFF_X1 \f7_reg[29]  ( .D(n772), .CK(clk), .Q(f7[29]) );
  DFF_X1 \f6_reg[27]  ( .D(n802), .CK(clk), .Q(n1044) );
  DFF_X1 \f6_reg[29]  ( .D(n804), .CK(clk), .Q(n1052) );
  DFF_X1 \f6_reg[26]  ( .D(n801), .CK(clk), .Q(n1040) );
  DFF_X1 \f6_reg[31]  ( .D(n806), .CK(clk), .Q(n1064) );
  DFF_X1 \f6_reg[28]  ( .D(n803), .CK(clk), .Q(n1048) );
  DFF_X1 \f6_reg[30]  ( .D(n805), .CK(clk), .Q(n1056) );
  DFF_X2 \f8_reg[31]  ( .D(n742), .CK(clk), .Q(f8[31]), .QN(n233) );
  DFF_X1 \f8_reg[26]  ( .D(n737), .CK(clk), .Q(f8[26]), .QN(n238) );
  DFF_X1 \f8_reg[27]  ( .D(n738), .CK(clk), .Q(f8[27]), .QN(n237) );
  DFF_X1 \f4_reg[27]  ( .D(n866), .CK(clk), .Q(f4[27]), .QN(n109) );
  DFF_X1 \f1_reg[27]  ( .D(n962), .CK(clk), .Q(f1[27]), .QN(n1042) );
  DFF_X1 \f1_reg[25]  ( .D(n960), .CK(clk), .Q(f1[25]), .QN(n1034) );
  DFF_X1 \f1_reg[26]  ( .D(n961), .CK(clk), .Q(f1[26]), .QN(n1038) );
  DFF_X1 \f1_reg[28]  ( .D(n963), .CK(clk), .Q(f1[28]), .QN(n1046) );
  DFF_X1 \f1_reg[30]  ( .D(n965), .CK(clk), .Q(f1[30]), .QN(n1054) );
  DFF_X2 \f8_reg[24]  ( .D(n735), .CK(clk), .Q(f8[24]), .QN(n240) );
  DFF_X1 \f8_reg[30]  ( .D(n741), .CK(clk), .Q(f8[30]), .QN(n234) );
  DFF_X1 \f8_reg[29]  ( .D(n740), .CK(clk), .Q(f8[29]), .QN(n235) );
  BUF_X1 U3 ( .A(data_out_x[12]), .Z(n3) );
  OR2_X1 U4 ( .A1(n110), .A2(n330), .ZN(n1) );
  NAND2_X1 U5 ( .A1(n1), .A2(n536), .ZN(n865) );
  CLKBUF_X1 U6 ( .A(data_out_x[9]), .Z(n172) );
  CLKBUF_X1 U7 ( .A(data_out_x[9]), .Z(n171) );
  BUF_X1 U8 ( .A(data_out_x[12]), .Z(n2) );
  BUF_X1 U9 ( .A(data_out_x[9]), .Z(n205) );
  BUF_X1 U10 ( .A(data_out_x[8]), .Z(n170) );
  BUF_X1 U11 ( .A(data_out_x[6]), .Z(n179) );
  OR2_X1 U12 ( .A1(n237), .A2(n322), .ZN(n4) );
  NAND2_X1 U13 ( .A1(n503), .A2(n4), .ZN(n738) );
  OR2_X1 U14 ( .A1(n238), .A2(n322), .ZN(n5) );
  NAND2_X1 U15 ( .A1(n504), .A2(n5), .ZN(n737) );
  OR2_X1 U16 ( .A1(n1054), .A2(n376), .ZN(n6) );
  NAND2_X1 U17 ( .A1(n392), .A2(n6), .ZN(n965) );
  OR2_X1 U18 ( .A1(n1046), .A2(n376), .ZN(n7) );
  NAND2_X1 U19 ( .A1(n394), .A2(n7), .ZN(n963) );
  OR2_X1 U20 ( .A1(n1038), .A2(n376), .ZN(n8) );
  NAND2_X1 U21 ( .A1(n396), .A2(n8), .ZN(n961) );
  OR2_X1 U22 ( .A1(n1034), .A2(n314), .ZN(n9) );
  NAND2_X1 U23 ( .A1(n397), .A2(n9), .ZN(n960) );
  OR2_X1 U24 ( .A1(n1042), .A2(n376), .ZN(n10) );
  NAND2_X1 U25 ( .A1(n395), .A2(n10), .ZN(n962) );
  OR2_X1 U26 ( .A1(n235), .A2(n322), .ZN(n11) );
  NAND2_X1 U27 ( .A1(n501), .A2(n11), .ZN(n740) );
  OR2_X1 U28 ( .A1(n234), .A2(n321), .ZN(n12) );
  NAND2_X1 U29 ( .A1(n500), .A2(n12), .ZN(n741) );
  OR2_X1 U30 ( .A1(n233), .A2(n321), .ZN(n13) );
  NAND2_X1 U31 ( .A1(n499), .A2(n13), .ZN(n742) );
  BUF_X1 U32 ( .A(data_out_x[6]), .Z(n201) );
  OR2_X1 U33 ( .A1(n107), .A2(n329), .ZN(n102) );
  NAND2_X1 U34 ( .A1(n102), .A2(n533), .ZN(n868) );
  OR2_X1 U35 ( .A1(n106), .A2(n329), .ZN(n103) );
  NAND2_X1 U36 ( .A1(n103), .A2(n532), .ZN(n869) );
  AOI22_X1 U37 ( .A1(n968), .A2(n1056), .B1(add_r6[30]), .B2(n177), .ZN(n434)
         );
  OR2_X1 U38 ( .A1(n1058), .A2(n376), .ZN(n104) );
  NAND2_X1 U39 ( .A1(n391), .A2(n104), .ZN(n966) );
  BUF_X1 U40 ( .A(data_out_x[8]), .Z(n169) );
  BUF_X2 U41 ( .A(data_out_x[10]), .Z(n202) );
  OR2_X1 U42 ( .A1(n108), .A2(n329), .ZN(n173) );
  NAND2_X1 U43 ( .A1(n173), .A2(n534), .ZN(n867) );
  BUF_X1 U44 ( .A(data_out_x[6]), .Z(n180) );
  OR2_X1 U45 ( .A1(n239), .A2(n322), .ZN(n174) );
  NAND2_X1 U46 ( .A1(n505), .A2(n174), .ZN(n736) );
  OR2_X1 U47 ( .A1(n236), .A2(n322), .ZN(n175) );
  NAND2_X1 U48 ( .A1(n502), .A2(n175), .ZN(n739) );
  OR2_X1 U49 ( .A1(n1050), .A2(n376), .ZN(n176) );
  NAND2_X1 U50 ( .A1(n393), .A2(n176), .ZN(n964) );
  BUF_X2 U51 ( .A(data_out_x[5]), .Z(n204) );
  AND2_X1 U52 ( .A1(n380), .A2(n1067), .ZN(n177) );
  BUF_X1 U53 ( .A(n207), .Z(n227) );
  BUF_X1 U54 ( .A(n207), .Z(n228) );
  BUF_X1 U55 ( .A(n207), .Z(n225) );
  BUF_X1 U56 ( .A(n207), .Z(n226) );
  BUF_X1 U57 ( .A(n208), .Z(n231) );
  BUF_X1 U58 ( .A(n207), .Z(n229) );
  BUF_X1 U59 ( .A(n208), .Z(n230) );
  BUF_X1 U60 ( .A(n207), .Z(n224) );
  INV_X1 U61 ( .A(n313), .ZN(n297) );
  INV_X1 U62 ( .A(n310), .ZN(n309) );
  BUF_X1 U63 ( .A(n209), .Z(n273) );
  BUF_X1 U64 ( .A(n210), .Z(n278) );
  BUF_X1 U65 ( .A(n210), .Z(n279) );
  BUF_X1 U66 ( .A(n210), .Z(n282) );
  BUF_X1 U67 ( .A(n209), .Z(n269) );
  BUF_X1 U68 ( .A(n208), .Z(n232) );
  BUF_X1 U69 ( .A(n209), .Z(n271) );
  BUF_X1 U70 ( .A(n209), .Z(n272) );
  BUF_X1 U71 ( .A(n208), .Z(n265) );
  BUF_X1 U72 ( .A(n209), .Z(n270) );
  BUF_X1 U73 ( .A(n208), .Z(n266) );
  BUF_X1 U74 ( .A(n208), .Z(n267) );
  BUF_X1 U75 ( .A(n209), .Z(n268) );
  INV_X1 U76 ( .A(n178), .ZN(n384) );
  BUF_X1 U77 ( .A(n277), .Z(n385) );
  BUF_X1 U78 ( .A(n281), .Z(n382) );
  BUF_X1 U79 ( .A(n280), .Z(n383) );
  BUF_X1 U80 ( .A(n276), .Z(n386) );
  BUF_X1 U81 ( .A(n379), .Z(n313) );
  BUF_X1 U82 ( .A(n379), .Z(n310) );
  BUF_X1 U83 ( .A(n377), .Z(n326) );
  BUF_X1 U84 ( .A(n377), .Z(n325) );
  BUF_X1 U85 ( .A(n378), .Z(n322) );
  BUF_X1 U86 ( .A(n377), .Z(n375) );
  BUF_X1 U87 ( .A(n377), .Z(n330) );
  BUF_X1 U88 ( .A(n377), .Z(n329) );
  BUF_X1 U89 ( .A(n378), .Z(n321) );
  BUF_X1 U90 ( .A(n376), .Z(n318) );
  BUF_X1 U91 ( .A(n376), .Z(n317) );
  BUF_X1 U92 ( .A(n377), .Z(n314) );
  BUF_X1 U93 ( .A(n211), .Z(n209) );
  BUF_X1 U94 ( .A(n212), .Z(n208) );
  BUF_X1 U95 ( .A(n212), .Z(n207) );
  INV_X1 U96 ( .A(n414), .ZN(n1069) );
  BUF_X1 U97 ( .A(n211), .Z(n210) );
  NAND2_X1 U98 ( .A1(n1059), .A2(n420), .ZN(n1060) );
  NAND2_X1 U99 ( .A1(n419), .A2(n1071), .ZN(n286) );
  NAND2_X1 U100 ( .A1(n416), .A2(n415), .ZN(n206) );
  NOR3_X1 U101 ( .A1(n412), .A2(n413), .A3(n414), .ZN(n410) );
  NAND2_X1 U102 ( .A1(n416), .A2(n415), .ZN(n285) );
  NAND2_X1 U103 ( .A1(n415), .A2(n1070), .ZN(n414) );
  INV_X1 U104 ( .A(n416), .ZN(n1070) );
  AND2_X1 U105 ( .A1(n410), .A2(n411), .ZN(n178) );
  NAND2_X1 U106 ( .A1(n410), .A2(n1068), .ZN(n281) );
  INV_X1 U107 ( .A(n411), .ZN(n1068) );
  AND2_X1 U108 ( .A1(n417), .A2(n1071), .ZN(n276) );
  NAND2_X1 U109 ( .A1(n1069), .A2(n412), .ZN(n280) );
  AND2_X1 U110 ( .A1(n413), .A2(n1069), .ZN(n277) );
  BUF_X1 U111 ( .A(n177), .Z(n211) );
  BUF_X1 U112 ( .A(n177), .Z(n212) );
  BUF_X1 U113 ( .A(n378), .Z(n379) );
  BUF_X1 U114 ( .A(n380), .Z(n377) );
  BUF_X1 U115 ( .A(n380), .Z(n378) );
  BUF_X1 U116 ( .A(n380), .Z(n376) );
  NOR3_X1 U117 ( .A1(n417), .A2(n419), .A3(n420), .ZN(n415) );
  NOR3_X1 U118 ( .A1(n387), .A2(addr_y[2]), .A3(n388), .ZN(n412) );
  NOR3_X1 U119 ( .A1(n387), .A2(addr_y[1]), .A3(n389), .ZN(n419) );
  NOR3_X1 U120 ( .A1(n389), .A2(addr_y[0]), .A3(n388), .ZN(n417) );
  NOR2_X1 U121 ( .A1(n389), .A2(addr_y[0]), .ZN(n416) );
  NOR2_X1 U122 ( .A1(n387), .A2(addr_y[1]), .ZN(n411) );
  NOR2_X1 U123 ( .A1(n388), .A2(addr_y[0]), .ZN(n413) );
  INV_X1 U124 ( .A(n420), .ZN(n1071) );
  INV_X1 U125 ( .A(n968), .ZN(n380) );
  NAND2_X1 U126 ( .A1(n311), .A2(n312), .ZN(n686) );
  NAND2_X1 U127 ( .A1(n295), .A2(n296), .ZN(n682) );
  NAND2_X1 U128 ( .A1(n291), .A2(n292), .ZN(n681) );
  NAND2_X1 U129 ( .A1(n287), .A2(n288), .ZN(n680) );
  NAND2_X1 U130 ( .A1(n274), .A2(n275), .ZN(n679) );
  OAI222_X1 U131 ( .A1(n384), .A2(n95), .B1(n280), .B2(n159), .C1(n281), .C2(
        n63), .ZN(n373) );
  OAI222_X1 U132 ( .A1(n384), .A2(n94), .B1(n280), .B2(n158), .C1(n281), .C2(
        n62), .ZN(n369) );
  OAI222_X1 U133 ( .A1(n384), .A2(n93), .B1(n280), .B2(n157), .C1(n281), .C2(
        n61), .ZN(n365) );
  OAI222_X1 U134 ( .A1(n384), .A2(n92), .B1(n280), .B2(n156), .C1(n281), .C2(
        n60), .ZN(n361) );
  OAI222_X1 U135 ( .A1(n384), .A2(n91), .B1(n280), .B2(n155), .C1(n281), .C2(
        n59), .ZN(n357) );
  OAI222_X1 U136 ( .A1(n384), .A2(n90), .B1(n280), .B2(n154), .C1(n281), .C2(
        n58), .ZN(n353) );
  OAI222_X1 U137 ( .A1(n384), .A2(n89), .B1(n280), .B2(n153), .C1(n281), .C2(
        n57), .ZN(n349) );
  OAI222_X1 U138 ( .A1(n384), .A2(n88), .B1(n280), .B2(n152), .C1(n281), .C2(
        n56), .ZN(n345) );
  OAI222_X1 U139 ( .A1(n384), .A2(n87), .B1(n280), .B2(n151), .C1(n281), .C2(
        n55), .ZN(n341) );
  OAI222_X1 U140 ( .A1(n384), .A2(n86), .B1(n280), .B2(n150), .C1(n281), .C2(
        n54), .ZN(n337) );
  OAI222_X1 U141 ( .A1(n384), .A2(n85), .B1(n280), .B2(n149), .C1(n281), .C2(
        n53), .ZN(n333) );
  NAND2_X1 U142 ( .A1(clc1), .A2(n1067), .ZN(n420) );
  NAND2_X1 U143 ( .A1(n327), .A2(n328), .ZN(n690) );
  NAND2_X1 U144 ( .A1(n323), .A2(n324), .ZN(n689) );
  NAND2_X1 U145 ( .A1(n319), .A2(n320), .ZN(n688) );
  NAND2_X1 U146 ( .A1(n315), .A2(n316), .ZN(n687) );
  NAND2_X1 U147 ( .A1(n307), .A2(n308), .ZN(n685) );
  NAND2_X1 U148 ( .A1(n303), .A2(n304), .ZN(n684) );
  NAND2_X1 U149 ( .A1(n299), .A2(n300), .ZN(n683) );
  NAND2_X1 U150 ( .A1(n371), .A2(n372), .ZN(n701) );
  AOI221_X1 U151 ( .B1(f1[9]), .B2(n381), .C1(f[9]), .C2(n1066), .A(n374), 
        .ZN(n371) );
  AOI221_X1 U152 ( .B1(f8[9]), .B2(n386), .C1(f4[9]), .C2(n385), .A(n373), 
        .ZN(n372) );
  OAI22_X1 U153 ( .A1(n206), .A2(n191), .B1(n286), .B2(n223), .ZN(n374) );
  NAND2_X1 U154 ( .A1(n367), .A2(n368), .ZN(n700) );
  AOI221_X1 U155 ( .B1(f1[10]), .B2(n381), .C1(f[10]), .C2(n1066), .A(n370), 
        .ZN(n367) );
  AOI221_X1 U156 ( .B1(f8[10]), .B2(n386), .C1(f4[10]), .C2(n385), .A(n369), 
        .ZN(n368) );
  OAI22_X1 U157 ( .A1(n285), .A2(n190), .B1(n286), .B2(n222), .ZN(n370) );
  NAND2_X1 U158 ( .A1(n363), .A2(n364), .ZN(n699) );
  AOI221_X1 U159 ( .B1(f1[11]), .B2(n381), .C1(f[11]), .C2(n1066), .A(n366), 
        .ZN(n363) );
  AOI221_X1 U160 ( .B1(f8[11]), .B2(n386), .C1(f4[11]), .C2(n385), .A(n365), 
        .ZN(n364) );
  OAI22_X1 U161 ( .A1(n206), .A2(n189), .B1(n286), .B2(n221), .ZN(n366) );
  NAND2_X1 U162 ( .A1(n359), .A2(n360), .ZN(n698) );
  AOI221_X1 U163 ( .B1(f1[12]), .B2(n381), .C1(f[12]), .C2(n1066), .A(n362), 
        .ZN(n359) );
  AOI221_X1 U164 ( .B1(f8[12]), .B2(n386), .C1(f4[12]), .C2(n385), .A(n361), 
        .ZN(n360) );
  OAI22_X1 U165 ( .A1(n285), .A2(n188), .B1(n286), .B2(n220), .ZN(n362) );
  NAND2_X1 U166 ( .A1(n355), .A2(n356), .ZN(n697) );
  AOI221_X1 U167 ( .B1(f1[13]), .B2(n381), .C1(f[13]), .C2(n1066), .A(n358), 
        .ZN(n355) );
  AOI221_X1 U168 ( .B1(f8[13]), .B2(n386), .C1(f4[13]), .C2(n385), .A(n357), 
        .ZN(n356) );
  OAI22_X1 U169 ( .A1(n206), .A2(n187), .B1(n286), .B2(n219), .ZN(n358) );
  NAND2_X1 U170 ( .A1(n351), .A2(n352), .ZN(n696) );
  AOI221_X1 U171 ( .B1(f1[14]), .B2(n381), .C1(f[14]), .C2(n1066), .A(n354), 
        .ZN(n351) );
  AOI221_X1 U172 ( .B1(f8[14]), .B2(n386), .C1(f4[14]), .C2(n385), .A(n353), 
        .ZN(n352) );
  OAI22_X1 U173 ( .A1(n285), .A2(n186), .B1(n286), .B2(n218), .ZN(n354) );
  NAND2_X1 U174 ( .A1(n347), .A2(n348), .ZN(n695) );
  AOI221_X1 U175 ( .B1(f1[15]), .B2(n381), .C1(f[15]), .C2(n1066), .A(n350), 
        .ZN(n347) );
  AOI221_X1 U176 ( .B1(f8[15]), .B2(n386), .C1(f4[15]), .C2(n385), .A(n349), 
        .ZN(n348) );
  OAI22_X1 U177 ( .A1(n206), .A2(n185), .B1(n286), .B2(n217), .ZN(n350) );
  NAND2_X1 U178 ( .A1(n343), .A2(n344), .ZN(n694) );
  AOI221_X1 U179 ( .B1(f1[16]), .B2(n381), .C1(f[16]), .C2(n1066), .A(n346), 
        .ZN(n343) );
  AOI221_X1 U180 ( .B1(f8[16]), .B2(n386), .C1(f4[16]), .C2(n385), .A(n345), 
        .ZN(n344) );
  OAI22_X1 U181 ( .A1(n285), .A2(n184), .B1(n286), .B2(n216), .ZN(n346) );
  NAND2_X1 U182 ( .A1(n339), .A2(n340), .ZN(n693) );
  AOI221_X1 U183 ( .B1(f1[17]), .B2(n381), .C1(f[17]), .C2(n1066), .A(n342), 
        .ZN(n339) );
  AOI221_X1 U184 ( .B1(f8[17]), .B2(n386), .C1(f4[17]), .C2(n385), .A(n341), 
        .ZN(n340) );
  OAI22_X1 U185 ( .A1(n206), .A2(n183), .B1(n286), .B2(n215), .ZN(n342) );
  NAND2_X1 U186 ( .A1(n335), .A2(n336), .ZN(n692) );
  AOI221_X1 U187 ( .B1(f1[18]), .B2(n381), .C1(f[18]), .C2(n1066), .A(n338), 
        .ZN(n335) );
  AOI221_X1 U188 ( .B1(f8[18]), .B2(n386), .C1(f4[18]), .C2(n385), .A(n337), 
        .ZN(n336) );
  OAI22_X1 U189 ( .A1(n285), .A2(n182), .B1(n286), .B2(n214), .ZN(n338) );
  NAND2_X1 U190 ( .A1(n331), .A2(n332), .ZN(n691) );
  AOI221_X1 U191 ( .B1(f1[19]), .B2(n381), .C1(f[19]), .C2(n1066), .A(n334), 
        .ZN(n331) );
  AOI221_X1 U192 ( .B1(f8[19]), .B2(n386), .C1(f4[19]), .C2(n385), .A(n333), 
        .ZN(n332) );
  OAI22_X1 U193 ( .A1(n206), .A2(n181), .B1(n286), .B2(n213), .ZN(n334) );
  BUF_X2 U194 ( .A(data_out_x[14]), .Z(n203) );
  CLKBUF_X1 U195 ( .A(n210), .Z(n283) );
  INV_X1 U196 ( .A(n313), .ZN(n284) );
  INV_X1 U197 ( .A(n313), .ZN(n289) );
  INV_X1 U198 ( .A(n313), .ZN(n290) );
  INV_X1 U199 ( .A(n313), .ZN(n293) );
  INV_X1 U200 ( .A(n313), .ZN(n294) );
  INV_X1 U201 ( .A(n310), .ZN(n298) );
  INV_X1 U202 ( .A(n310), .ZN(n301) );
  INV_X1 U203 ( .A(n310), .ZN(n302) );
  INV_X1 U204 ( .A(n310), .ZN(n305) );
  INV_X1 U205 ( .A(n310), .ZN(n306) );
  INV_X1 U206 ( .A(n1059), .ZN(n381) );
  INV_X1 U207 ( .A(addr_y[0]), .ZN(n387) );
  INV_X1 U208 ( .A(addr_y[1]), .ZN(n388) );
  INV_X1 U209 ( .A(addr_y[2]), .ZN(n389) );
  INV_X1 U210 ( .A(clc1), .ZN(n390) );
  INV_X1 U211 ( .A(clear_acc), .ZN(n1067) );
  NAND3_X1 U212 ( .A1(clc), .A2(n1067), .A3(n390), .ZN(n1059) );
  OAI21_X1 U213 ( .B1(clear_acc), .B2(n390), .A(n1059), .ZN(n968) );
  NAND2_X1 U214 ( .A1(add_r1[31]), .A2(n224), .ZN(n391) );
  NAND2_X1 U215 ( .A1(add_r1[30]), .A2(n230), .ZN(n392) );
  NAND2_X1 U216 ( .A1(add_r1[29]), .A2(n230), .ZN(n393) );
  NAND2_X1 U217 ( .A1(add_r1[28]), .A2(n229), .ZN(n394) );
  NAND2_X1 U218 ( .A1(add_r1[27]), .A2(n230), .ZN(n395) );
  NAND2_X1 U219 ( .A1(add_r1[26]), .A2(n229), .ZN(n396) );
  NAND2_X1 U220 ( .A1(add_r1[25]), .A2(n229), .ZN(n397) );
  NAND2_X1 U221 ( .A1(add_r1[24]), .A2(n230), .ZN(n398) );
  OAI21_X1 U222 ( .B1(n16), .B2(n314), .A(n398), .ZN(n959) );
  NAND2_X1 U223 ( .A1(add_r1[23]), .A2(n229), .ZN(n399) );
  OAI21_X1 U224 ( .B1(n1027), .B2(n314), .A(n399), .ZN(n958) );
  NAND2_X1 U225 ( .A1(add_r1[22]), .A2(n230), .ZN(n400) );
  OAI21_X1 U226 ( .B1(n1023), .B2(n314), .A(n400), .ZN(n957) );
  NAND2_X1 U227 ( .A1(add_r1[21]), .A2(n230), .ZN(n401) );
  OAI21_X1 U228 ( .B1(n1019), .B2(n314), .A(n401), .ZN(n956) );
  NAND2_X1 U229 ( .A1(add_r1[20]), .A2(n229), .ZN(n402) );
  OAI21_X1 U230 ( .B1(n1015), .B2(n314), .A(n402), .ZN(n955) );
  NAND2_X1 U231 ( .A1(add_r1[19]), .A2(n231), .ZN(n403) );
  OAI21_X1 U232 ( .B1(n21), .B2(n314), .A(n403), .ZN(n954) );
  NAND2_X1 U233 ( .A1(add_r1[18]), .A2(n231), .ZN(n404) );
  OAI21_X1 U234 ( .B1(n22), .B2(n317), .A(n404), .ZN(n953) );
  NAND2_X1 U235 ( .A1(add_r1[17]), .A2(n230), .ZN(n405) );
  OAI21_X1 U236 ( .B1(n23), .B2(n317), .A(n405), .ZN(n952) );
  NAND2_X1 U237 ( .A1(add_r1[16]), .A2(n229), .ZN(n406) );
  OAI21_X1 U238 ( .B1(n24), .B2(n317), .A(n406), .ZN(n951) );
  NAND2_X1 U239 ( .A1(add_r1[15]), .A2(n230), .ZN(n407) );
  OAI21_X1 U240 ( .B1(n25), .B2(n317), .A(n407), .ZN(n950) );
  NAND2_X1 U241 ( .A1(add_r1[14]), .A2(n231), .ZN(n408) );
  OAI21_X1 U242 ( .B1(n26), .B2(n317), .A(n408), .ZN(n949) );
  NAND2_X1 U243 ( .A1(add_r1[13]), .A2(n229), .ZN(n409) );
  OAI21_X1 U244 ( .B1(n27), .B2(n317), .A(n409), .ZN(n948) );
  NAND2_X1 U245 ( .A1(add_r1[12]), .A2(n231), .ZN(n418) );
  OAI21_X1 U246 ( .B1(n28), .B2(n317), .A(n418), .ZN(n947) );
  NAND2_X1 U247 ( .A1(add_r1[11]), .A2(n230), .ZN(n421) );
  OAI21_X1 U248 ( .B1(n29), .B2(n318), .A(n421), .ZN(n946) );
  NAND2_X1 U249 ( .A1(add_r1[10]), .A2(n231), .ZN(n422) );
  OAI21_X1 U250 ( .B1(n30), .B2(n318), .A(n422), .ZN(n945) );
  NAND2_X1 U251 ( .A1(add_r1[9]), .A2(n230), .ZN(n423) );
  OAI21_X1 U252 ( .B1(n31), .B2(n318), .A(n423), .ZN(n944) );
  NAND2_X1 U253 ( .A1(add_r1[7]), .A2(n231), .ZN(n424) );
  OAI21_X1 U254 ( .B1(n975), .B2(n318), .A(n424), .ZN(n942) );
  NAND2_X1 U255 ( .A1(add_r1[6]), .A2(n231), .ZN(n425) );
  OAI21_X1 U256 ( .B1(n980), .B2(n318), .A(n425), .ZN(n941) );
  NAND2_X1 U257 ( .A1(add_r1[5]), .A2(n230), .ZN(n426) );
  OAI21_X1 U258 ( .B1(n985), .B2(n318), .A(n426), .ZN(n940) );
  NAND2_X1 U259 ( .A1(add_r1[4]), .A2(n231), .ZN(n427) );
  OAI21_X1 U260 ( .B1(n990), .B2(n318), .A(n427), .ZN(n939) );
  NAND2_X1 U261 ( .A1(add_r1[3]), .A2(n231), .ZN(n428) );
  OAI21_X1 U262 ( .B1(n995), .B2(n321), .A(n428), .ZN(n938) );
  NAND2_X1 U263 ( .A1(add_r1[2]), .A2(n231), .ZN(n429) );
  OAI21_X1 U264 ( .B1(n1000), .B2(n321), .A(n429), .ZN(n937) );
  NAND2_X1 U265 ( .A1(add_r1[1]), .A2(n230), .ZN(n430) );
  OAI21_X1 U266 ( .B1(n1005), .B2(n321), .A(n430), .ZN(n936) );
  NAND2_X1 U267 ( .A1(add_r1[0]), .A2(n231), .ZN(n431) );
  OAI21_X1 U268 ( .B1(n1010), .B2(n321), .A(n431), .ZN(n935) );
  NAND2_X1 U269 ( .A1(add_r1[8]), .A2(n231), .ZN(n432) );
  OAI21_X1 U270 ( .B1(n970), .B2(n321), .A(n432), .ZN(n943) );
  AOI22_X1 U271 ( .A1(n294), .A2(n1064), .B1(add_r6[31]), .B2(n265), .ZN(n433)
         );
  INV_X1 U272 ( .A(n433), .ZN(n806) );
  INV_X1 U273 ( .A(n434), .ZN(n805) );
  AOI22_X1 U274 ( .A1(n297), .A2(n1052), .B1(add_r6[29]), .B2(n283), .ZN(n435)
         );
  INV_X1 U275 ( .A(n435), .ZN(n804) );
  AOI22_X1 U276 ( .A1(n306), .A2(n1048), .B1(add_r6[28]), .B2(n283), .ZN(n436)
         );
  INV_X1 U277 ( .A(n436), .ZN(n803) );
  AOI22_X1 U278 ( .A1(n305), .A2(n1044), .B1(add_r6[27]), .B2(n283), .ZN(n437)
         );
  INV_X1 U279 ( .A(n437), .ZN(n802) );
  AOI22_X1 U280 ( .A1(n293), .A2(n1040), .B1(add_r6[26]), .B2(n282), .ZN(n438)
         );
  INV_X1 U281 ( .A(n438), .ZN(n801) );
  AOI22_X1 U282 ( .A1(n290), .A2(n1036), .B1(add_r6[25]), .B2(n282), .ZN(n439)
         );
  INV_X1 U283 ( .A(n439), .ZN(n800) );
  AOI22_X1 U284 ( .A1(n289), .A2(f6[24]), .B1(add_r6[24]), .B2(n282), .ZN(n440) );
  INV_X1 U285 ( .A(n440), .ZN(n799) );
  AOI22_X1 U286 ( .A1(n284), .A2(f6[23]), .B1(add_r6[23]), .B2(n282), .ZN(n441) );
  INV_X1 U287 ( .A(n441), .ZN(n798) );
  AOI22_X1 U288 ( .A1(n297), .A2(f6[22]), .B1(add_r6[22]), .B2(n282), .ZN(n442) );
  INV_X1 U289 ( .A(n442), .ZN(n797) );
  AOI22_X1 U290 ( .A1(n306), .A2(f6[21]), .B1(add_r6[21]), .B2(n282), .ZN(n443) );
  INV_X1 U291 ( .A(n443), .ZN(n796) );
  AOI22_X1 U292 ( .A1(n305), .A2(f6[20]), .B1(add_r6[20]), .B2(n282), .ZN(n444) );
  INV_X1 U293 ( .A(n444), .ZN(n795) );
  AOI22_X1 U294 ( .A1(n284), .A2(f6[19]), .B1(add_r6[19]), .B2(n282), .ZN(n445) );
  INV_X1 U295 ( .A(n445), .ZN(n794) );
  AOI22_X1 U296 ( .A1(n284), .A2(f6[18]), .B1(add_r6[18]), .B2(n282), .ZN(n446) );
  INV_X1 U297 ( .A(n446), .ZN(n793) );
  AOI22_X1 U298 ( .A1(n284), .A2(f6[17]), .B1(add_r6[17]), .B2(n282), .ZN(n447) );
  INV_X1 U299 ( .A(n447), .ZN(n792) );
  AOI22_X1 U300 ( .A1(n284), .A2(f6[16]), .B1(add_r6[16]), .B2(n282), .ZN(n448) );
  INV_X1 U301 ( .A(n448), .ZN(n791) );
  AOI22_X1 U302 ( .A1(n284), .A2(f6[15]), .B1(add_r6[15]), .B2(n282), .ZN(n449) );
  INV_X1 U303 ( .A(n449), .ZN(n790) );
  AOI22_X1 U304 ( .A1(n284), .A2(f6[14]), .B1(add_r6[14]), .B2(n279), .ZN(n450) );
  INV_X1 U305 ( .A(n450), .ZN(n789) );
  AOI22_X1 U306 ( .A1(n284), .A2(f6[13]), .B1(add_r6[13]), .B2(n279), .ZN(n451) );
  INV_X1 U307 ( .A(n451), .ZN(n788) );
  AOI22_X1 U308 ( .A1(n284), .A2(f6[12]), .B1(add_r6[12]), .B2(n279), .ZN(n452) );
  INV_X1 U309 ( .A(n452), .ZN(n787) );
  AOI22_X1 U310 ( .A1(n284), .A2(f6[11]), .B1(add_r6[11]), .B2(n279), .ZN(n453) );
  INV_X1 U311 ( .A(n453), .ZN(n786) );
  AOI22_X1 U312 ( .A1(n284), .A2(f6[10]), .B1(add_r6[10]), .B2(n279), .ZN(n454) );
  INV_X1 U313 ( .A(n454), .ZN(n785) );
  AOI22_X1 U314 ( .A1(n284), .A2(f6[9]), .B1(add_r6[9]), .B2(n279), .ZN(n455)
         );
  INV_X1 U315 ( .A(n455), .ZN(n784) );
  AOI22_X1 U316 ( .A1(n284), .A2(f6[7]), .B1(add_r6[7]), .B2(n279), .ZN(n456)
         );
  INV_X1 U317 ( .A(n456), .ZN(n782) );
  AOI22_X1 U318 ( .A1(n289), .A2(f6[6]), .B1(add_r6[6]), .B2(n279), .ZN(n457)
         );
  INV_X1 U319 ( .A(n457), .ZN(n781) );
  AOI22_X1 U320 ( .A1(n289), .A2(f6[5]), .B1(add_r6[5]), .B2(n279), .ZN(n458)
         );
  INV_X1 U321 ( .A(n458), .ZN(n780) );
  AOI22_X1 U322 ( .A1(n289), .A2(f6[4]), .B1(add_r6[4]), .B2(n279), .ZN(n459)
         );
  INV_X1 U323 ( .A(n459), .ZN(n779) );
  AOI22_X1 U324 ( .A1(n289), .A2(f6[3]), .B1(add_r6[3]), .B2(n279), .ZN(n460)
         );
  INV_X1 U325 ( .A(n460), .ZN(n778) );
  AOI22_X1 U326 ( .A1(n289), .A2(f6[2]), .B1(add_r6[2]), .B2(n279), .ZN(n461)
         );
  INV_X1 U327 ( .A(n461), .ZN(n777) );
  AOI22_X1 U328 ( .A1(n289), .A2(f6[1]), .B1(add_r6[1]), .B2(n278), .ZN(n462)
         );
  INV_X1 U329 ( .A(n462), .ZN(n776) );
  AOI22_X1 U330 ( .A1(n289), .A2(f6[0]), .B1(add_r6[0]), .B2(n278), .ZN(n463)
         );
  INV_X1 U331 ( .A(n463), .ZN(n775) );
  AOI22_X1 U332 ( .A1(n289), .A2(f6[8]), .B1(add_r6[8]), .B2(n278), .ZN(n464)
         );
  INV_X1 U333 ( .A(n464), .ZN(n783) );
  AOI22_X1 U334 ( .A1(n289), .A2(f7[31]), .B1(add_r7[31]), .B2(n278), .ZN(n465) );
  INV_X1 U335 ( .A(n465), .ZN(n774) );
  AOI22_X1 U336 ( .A1(n289), .A2(f7[30]), .B1(add_r7[30]), .B2(n278), .ZN(n466) );
  INV_X1 U337 ( .A(n466), .ZN(n773) );
  AOI22_X1 U338 ( .A1(n289), .A2(f7[29]), .B1(add_r7[29]), .B2(n278), .ZN(n467) );
  INV_X1 U339 ( .A(n467), .ZN(n772) );
  AOI22_X1 U340 ( .A1(n289), .A2(f7[28]), .B1(add_r7[28]), .B2(n278), .ZN(n468) );
  INV_X1 U341 ( .A(n468), .ZN(n771) );
  AOI22_X1 U342 ( .A1(n290), .A2(f7[27]), .B1(add_r7[27]), .B2(n278), .ZN(n469) );
  INV_X1 U343 ( .A(n469), .ZN(n770) );
  AOI22_X1 U344 ( .A1(n290), .A2(f7[26]), .B1(add_r7[26]), .B2(n278), .ZN(n470) );
  INV_X1 U345 ( .A(n470), .ZN(n769) );
  AOI22_X1 U346 ( .A1(n290), .A2(f7[25]), .B1(add_r7[25]), .B2(n278), .ZN(n471) );
  INV_X1 U347 ( .A(n471), .ZN(n768) );
  AOI22_X1 U348 ( .A1(n290), .A2(n1032), .B1(add_r7[24]), .B2(n278), .ZN(n472)
         );
  INV_X1 U349 ( .A(n472), .ZN(n767) );
  AOI22_X1 U350 ( .A1(n290), .A2(n1029), .B1(add_r7[23]), .B2(n278), .ZN(n473)
         );
  INV_X1 U351 ( .A(n473), .ZN(n766) );
  AOI22_X1 U352 ( .A1(n290), .A2(n1025), .B1(add_r7[22]), .B2(n273), .ZN(n474)
         );
  INV_X1 U353 ( .A(n474), .ZN(n765) );
  AOI22_X1 U354 ( .A1(n290), .A2(n1021), .B1(add_r7[21]), .B2(n273), .ZN(n475)
         );
  INV_X1 U355 ( .A(n475), .ZN(n764) );
  AOI22_X1 U356 ( .A1(n290), .A2(n1017), .B1(add_r7[20]), .B2(n273), .ZN(n476)
         );
  INV_X1 U357 ( .A(n476), .ZN(n763) );
  AOI22_X1 U358 ( .A1(n290), .A2(n477), .B1(add_r7[19]), .B2(n273), .ZN(n478)
         );
  INV_X1 U359 ( .A(n478), .ZN(n762) );
  AOI22_X1 U360 ( .A1(n290), .A2(n479), .B1(add_r7[18]), .B2(n273), .ZN(n480)
         );
  INV_X1 U361 ( .A(n480), .ZN(n761) );
  AOI22_X1 U362 ( .A1(n290), .A2(f7[17]), .B1(add_r7[17]), .B2(n273), .ZN(n481) );
  INV_X1 U363 ( .A(n481), .ZN(n760) );
  AOI22_X1 U364 ( .A1(n290), .A2(f7[16]), .B1(add_r7[16]), .B2(n273), .ZN(n482) );
  INV_X1 U365 ( .A(n482), .ZN(n759) );
  AOI22_X1 U366 ( .A1(n293), .A2(f7[15]), .B1(add_r7[15]), .B2(n273), .ZN(n483) );
  INV_X1 U367 ( .A(n483), .ZN(n758) );
  AOI22_X1 U368 ( .A1(n293), .A2(f7[14]), .B1(add_r7[14]), .B2(n273), .ZN(n484) );
  INV_X1 U369 ( .A(n484), .ZN(n757) );
  AOI22_X1 U370 ( .A1(n293), .A2(f7[13]), .B1(add_r7[13]), .B2(n273), .ZN(n485) );
  INV_X1 U371 ( .A(n485), .ZN(n756) );
  AOI22_X1 U372 ( .A1(n293), .A2(f7[12]), .B1(add_r7[12]), .B2(n273), .ZN(n486) );
  INV_X1 U373 ( .A(n486), .ZN(n755) );
  AOI22_X1 U374 ( .A1(n293), .A2(f7[11]), .B1(add_r7[11]), .B2(n273), .ZN(n487) );
  INV_X1 U375 ( .A(n487), .ZN(n754) );
  AOI22_X1 U376 ( .A1(n293), .A2(f7[10]), .B1(add_r7[10]), .B2(n272), .ZN(n488) );
  INV_X1 U377 ( .A(n488), .ZN(n753) );
  AOI22_X1 U378 ( .A1(n293), .A2(f7[9]), .B1(add_r7[9]), .B2(n272), .ZN(n489)
         );
  INV_X1 U379 ( .A(n489), .ZN(n752) );
  AOI22_X1 U380 ( .A1(n293), .A2(f7[7]), .B1(add_r7[7]), .B2(n272), .ZN(n490)
         );
  INV_X1 U381 ( .A(n490), .ZN(n750) );
  AOI22_X1 U382 ( .A1(n293), .A2(f7[6]), .B1(add_r7[6]), .B2(n272), .ZN(n491)
         );
  INV_X1 U383 ( .A(n491), .ZN(n749) );
  AOI22_X1 U384 ( .A1(n293), .A2(f7[5]), .B1(add_r7[5]), .B2(n272), .ZN(n492)
         );
  INV_X1 U385 ( .A(n492), .ZN(n748) );
  AOI22_X1 U386 ( .A1(n293), .A2(f7[4]), .B1(add_r7[4]), .B2(n272), .ZN(n493)
         );
  INV_X1 U387 ( .A(n493), .ZN(n747) );
  AOI22_X1 U388 ( .A1(n293), .A2(f7[3]), .B1(add_r7[3]), .B2(n272), .ZN(n494)
         );
  INV_X1 U389 ( .A(n494), .ZN(n746) );
  AOI22_X1 U390 ( .A1(n294), .A2(f7[2]), .B1(add_r7[2]), .B2(n272), .ZN(n495)
         );
  INV_X1 U391 ( .A(n495), .ZN(n745) );
  AOI22_X1 U392 ( .A1(n294), .A2(f7[1]), .B1(add_r7[1]), .B2(n272), .ZN(n496)
         );
  INV_X1 U393 ( .A(n496), .ZN(n744) );
  AOI22_X1 U394 ( .A1(n294), .A2(f7[0]), .B1(add_r7[0]), .B2(n272), .ZN(n497)
         );
  INV_X1 U395 ( .A(n497), .ZN(n743) );
  AOI22_X1 U396 ( .A1(n294), .A2(f7[8]), .B1(add_r7[8]), .B2(n272), .ZN(n498)
         );
  INV_X1 U397 ( .A(n498), .ZN(n751) );
  NAND2_X1 U398 ( .A1(add_r8[31]), .A2(n229), .ZN(n499) );
  NAND2_X1 U399 ( .A1(add_r8[30]), .A2(n229), .ZN(n500) );
  NAND2_X1 U400 ( .A1(add_r8[29]), .A2(n229), .ZN(n501) );
  NAND2_X1 U401 ( .A1(add_r8[28]), .A2(n229), .ZN(n502) );
  NAND2_X1 U402 ( .A1(add_r8[27]), .A2(n228), .ZN(n503) );
  NAND2_X1 U403 ( .A1(add_r8[26]), .A2(n228), .ZN(n504) );
  NAND2_X1 U404 ( .A1(add_r8[25]), .A2(n228), .ZN(n505) );
  NAND2_X1 U405 ( .A1(add_r8[24]), .A2(n228), .ZN(n506) );
  OAI21_X1 U406 ( .B1(n240), .B2(n322), .A(n506), .ZN(n735) );
  NAND2_X1 U407 ( .A1(add_r8[23]), .A2(n228), .ZN(n507) );
  OAI21_X1 U408 ( .B1(n241), .B2(n322), .A(n507), .ZN(n734) );
  NAND2_X1 U409 ( .A1(add_r8[22]), .A2(n228), .ZN(n508) );
  OAI21_X1 U410 ( .B1(n242), .B2(n325), .A(n508), .ZN(n733) );
  NAND2_X1 U411 ( .A1(add_r8[21]), .A2(n228), .ZN(n509) );
  OAI21_X1 U412 ( .B1(n243), .B2(n325), .A(n509), .ZN(n732) );
  NAND2_X1 U413 ( .A1(add_r8[20]), .A2(n228), .ZN(n510) );
  OAI21_X1 U414 ( .B1(n244), .B2(n325), .A(n510), .ZN(n731) );
  NAND2_X1 U415 ( .A1(add_r8[19]), .A2(n228), .ZN(n511) );
  OAI21_X1 U416 ( .B1(n245), .B2(n325), .A(n511), .ZN(n730) );
  NAND2_X1 U417 ( .A1(add_r8[18]), .A2(n228), .ZN(n512) );
  OAI21_X1 U418 ( .B1(n246), .B2(n325), .A(n512), .ZN(n729) );
  NAND2_X1 U419 ( .A1(add_r8[17]), .A2(n228), .ZN(n513) );
  OAI21_X1 U420 ( .B1(n247), .B2(n325), .A(n513), .ZN(n728) );
  NAND2_X1 U421 ( .A1(add_r8[16]), .A2(n228), .ZN(n514) );
  OAI21_X1 U422 ( .B1(n248), .B2(n325), .A(n514), .ZN(n727) );
  NAND2_X1 U423 ( .A1(add_r8[15]), .A2(n227), .ZN(n515) );
  OAI21_X1 U424 ( .B1(n249), .B2(n326), .A(n515), .ZN(n726) );
  NAND2_X1 U425 ( .A1(add_r8[14]), .A2(n227), .ZN(n516) );
  OAI21_X1 U426 ( .B1(n250), .B2(n326), .A(n516), .ZN(n725) );
  NAND2_X1 U427 ( .A1(add_r8[13]), .A2(n227), .ZN(n517) );
  OAI21_X1 U428 ( .B1(n251), .B2(n326), .A(n517), .ZN(n724) );
  NAND2_X1 U429 ( .A1(add_r8[12]), .A2(n227), .ZN(n518) );
  OAI21_X1 U430 ( .B1(n252), .B2(n326), .A(n518), .ZN(n723) );
  NAND2_X1 U431 ( .A1(add_r8[11]), .A2(n227), .ZN(n519) );
  OAI21_X1 U432 ( .B1(n253), .B2(n326), .A(n519), .ZN(n722) );
  NAND2_X1 U433 ( .A1(add_r8[10]), .A2(n227), .ZN(n520) );
  OAI21_X1 U434 ( .B1(n254), .B2(n326), .A(n520), .ZN(n721) );
  NAND2_X1 U435 ( .A1(add_r8[9]), .A2(n227), .ZN(n521) );
  OAI21_X1 U436 ( .B1(n255), .B2(n326), .A(n521), .ZN(n720) );
  NAND2_X1 U437 ( .A1(add_r8[7]), .A2(n227), .ZN(n522) );
  OAI21_X1 U438 ( .B1(n257), .B2(n326), .A(n522), .ZN(n718) );
  NAND2_X1 U439 ( .A1(add_r8[6]), .A2(n227), .ZN(n523) );
  OAI21_X1 U440 ( .B1(n258), .B2(n375), .A(n523), .ZN(n717) );
  NAND2_X1 U441 ( .A1(add_r8[5]), .A2(n227), .ZN(n524) );
  OAI21_X1 U442 ( .B1(n259), .B2(n325), .A(n524), .ZN(n716) );
  NAND2_X1 U443 ( .A1(add_r8[4]), .A2(n227), .ZN(n525) );
  OAI21_X1 U444 ( .B1(n260), .B2(n330), .A(n525), .ZN(n715) );
  NAND2_X1 U445 ( .A1(add_r8[3]), .A2(n227), .ZN(n526) );
  OAI21_X1 U446 ( .B1(n261), .B2(n326), .A(n526), .ZN(n714) );
  NAND2_X1 U447 ( .A1(add_r8[2]), .A2(n226), .ZN(n527) );
  OAI21_X1 U448 ( .B1(n262), .B2(n375), .A(n527), .ZN(n713) );
  NAND2_X1 U449 ( .A1(add_r8[1]), .A2(n226), .ZN(n528) );
  OAI21_X1 U450 ( .B1(n263), .B2(n325), .A(n528), .ZN(n712) );
  NAND2_X1 U451 ( .A1(add_r8[0]), .A2(n226), .ZN(n529) );
  OAI21_X1 U452 ( .B1(n264), .B2(n329), .A(n529), .ZN(n711) );
  NAND2_X1 U453 ( .A1(add_r8[8]), .A2(n226), .ZN(n530) );
  OAI21_X1 U454 ( .B1(n256), .B2(n329), .A(n530), .ZN(n719) );
  NAND2_X1 U455 ( .A1(add_r4[31]), .A2(n226), .ZN(n531) );
  OAI21_X1 U456 ( .B1(n105), .B2(n329), .A(n531), .ZN(n870) );
  NAND2_X1 U457 ( .A1(add_r4[30]), .A2(n226), .ZN(n532) );
  NAND2_X1 U458 ( .A1(add_r4[29]), .A2(n226), .ZN(n533) );
  NAND2_X1 U459 ( .A1(add_r4[28]), .A2(n229), .ZN(n534) );
  NAND2_X1 U460 ( .A1(add_r4[27]), .A2(n226), .ZN(n535) );
  OAI21_X1 U461 ( .B1(n109), .B2(n329), .A(n535), .ZN(n866) );
  NAND2_X1 U462 ( .A1(add_r4[26]), .A2(n226), .ZN(n536) );
  NAND2_X1 U463 ( .A1(add_r4[25]), .A2(n226), .ZN(n537) );
  OAI21_X1 U464 ( .B1(n111), .B2(n330), .A(n537), .ZN(n864) );
  NAND2_X1 U465 ( .A1(add_r4[24]), .A2(n226), .ZN(n538) );
  OAI21_X1 U466 ( .B1(n112), .B2(n330), .A(n538), .ZN(n863) );
  NAND2_X1 U467 ( .A1(add_r4[23]), .A2(n226), .ZN(n539) );
  OAI21_X1 U468 ( .B1(n113), .B2(n330), .A(n539), .ZN(n862) );
  NAND2_X1 U469 ( .A1(add_r4[22]), .A2(n225), .ZN(n540) );
  OAI21_X1 U470 ( .B1(n114), .B2(n330), .A(n540), .ZN(n861) );
  NAND2_X1 U471 ( .A1(add_r4[21]), .A2(n225), .ZN(n541) );
  OAI21_X1 U472 ( .B1(n115), .B2(n330), .A(n541), .ZN(n860) );
  NAND2_X1 U473 ( .A1(add_r4[20]), .A2(n225), .ZN(n542) );
  OAI21_X1 U474 ( .B1(n116), .B2(n330), .A(n542), .ZN(n859) );
  NAND2_X1 U475 ( .A1(add_r4[19]), .A2(n225), .ZN(n543) );
  OAI21_X1 U476 ( .B1(n117), .B2(n375), .A(n543), .ZN(n858) );
  NAND2_X1 U477 ( .A1(add_r4[18]), .A2(n225), .ZN(n544) );
  OAI21_X1 U478 ( .B1(n118), .B2(n375), .A(n544), .ZN(n857) );
  NAND2_X1 U479 ( .A1(add_r4[17]), .A2(n225), .ZN(n545) );
  OAI21_X1 U480 ( .B1(n119), .B2(n375), .A(n545), .ZN(n856) );
  NAND2_X1 U481 ( .A1(add_r4[16]), .A2(n225), .ZN(n546) );
  OAI21_X1 U482 ( .B1(n120), .B2(n375), .A(n546), .ZN(n855) );
  NAND2_X1 U483 ( .A1(add_r4[15]), .A2(n225), .ZN(n547) );
  OAI21_X1 U484 ( .B1(n121), .B2(n375), .A(n547), .ZN(n854) );
  NAND2_X1 U485 ( .A1(add_r4[14]), .A2(n225), .ZN(n548) );
  OAI21_X1 U486 ( .B1(n122), .B2(n375), .A(n548), .ZN(n853) );
  NAND2_X1 U487 ( .A1(add_r4[13]), .A2(n225), .ZN(n549) );
  OAI21_X1 U488 ( .B1(n123), .B2(n375), .A(n549), .ZN(n852) );
  NAND2_X1 U489 ( .A1(add_r4[12]), .A2(n225), .ZN(n550) );
  OAI21_X1 U490 ( .B1(n124), .B2(n376), .A(n550), .ZN(n851) );
  NAND2_X1 U491 ( .A1(add_r4[11]), .A2(n225), .ZN(n551) );
  OAI21_X1 U492 ( .B1(n125), .B2(n376), .A(n551), .ZN(n850) );
  NAND2_X1 U493 ( .A1(add_r4[10]), .A2(n224), .ZN(n552) );
  OAI21_X1 U494 ( .B1(n126), .B2(n376), .A(n552), .ZN(n849) );
  NAND2_X1 U495 ( .A1(add_r4[9]), .A2(n224), .ZN(n553) );
  OAI21_X1 U496 ( .B1(n127), .B2(n376), .A(n553), .ZN(n848) );
  NAND2_X1 U497 ( .A1(add_r4[7]), .A2(n224), .ZN(n554) );
  OAI21_X1 U498 ( .B1(n129), .B2(n376), .A(n554), .ZN(n846) );
  NAND2_X1 U499 ( .A1(add_r4[6]), .A2(n224), .ZN(n555) );
  OAI21_X1 U500 ( .B1(n130), .B2(n376), .A(n555), .ZN(n845) );
  NAND2_X1 U501 ( .A1(add_r4[5]), .A2(n224), .ZN(n556) );
  OAI21_X1 U502 ( .B1(n131), .B2(n376), .A(n556), .ZN(n844) );
  NAND2_X1 U503 ( .A1(add_r4[4]), .A2(n224), .ZN(n557) );
  OAI21_X1 U504 ( .B1(n132), .B2(n330), .A(n557), .ZN(n843) );
  NAND2_X1 U505 ( .A1(add_r4[3]), .A2(n224), .ZN(n558) );
  OAI21_X1 U506 ( .B1(n133), .B2(n376), .A(n558), .ZN(n842) );
  NAND2_X1 U507 ( .A1(add_r4[2]), .A2(n224), .ZN(n559) );
  OAI21_X1 U508 ( .B1(n134), .B2(n376), .A(n559), .ZN(n841) );
  NAND2_X1 U509 ( .A1(add_r4[1]), .A2(n224), .ZN(n560) );
  OAI21_X1 U510 ( .B1(n135), .B2(n326), .A(n560), .ZN(n840) );
  NAND2_X1 U511 ( .A1(add_r4[0]), .A2(n224), .ZN(n561) );
  OAI21_X1 U512 ( .B1(n136), .B2(n376), .A(n561), .ZN(n839) );
  NAND2_X1 U513 ( .A1(add_r4[8]), .A2(n224), .ZN(n562) );
  OAI21_X1 U514 ( .B1(n128), .B2(n376), .A(n562), .ZN(n847) );
  AOI22_X1 U515 ( .A1(n294), .A2(n563), .B1(add_r3[31]), .B2(n272), .ZN(n564)
         );
  INV_X1 U516 ( .A(n564), .ZN(n902) );
  AOI22_X1 U517 ( .A1(n294), .A2(n565), .B1(add_r3[30]), .B2(n271), .ZN(n566)
         );
  INV_X1 U518 ( .A(n566), .ZN(n901) );
  AOI22_X1 U519 ( .A1(n294), .A2(n567), .B1(add_r3[29]), .B2(n271), .ZN(n568)
         );
  INV_X1 U520 ( .A(n568), .ZN(n900) );
  AOI22_X1 U521 ( .A1(n294), .A2(n569), .B1(add_r3[28]), .B2(n271), .ZN(n570)
         );
  INV_X1 U522 ( .A(n570), .ZN(n899) );
  AOI22_X1 U523 ( .A1(n294), .A2(n571), .B1(add_r3[27]), .B2(n271), .ZN(n572)
         );
  INV_X1 U524 ( .A(n572), .ZN(n898) );
  AOI22_X1 U525 ( .A1(n294), .A2(n573), .B1(add_r3[26]), .B2(n271), .ZN(n574)
         );
  INV_X1 U526 ( .A(n574), .ZN(n897) );
  AOI22_X1 U527 ( .A1(n294), .A2(n575), .B1(add_r3[25]), .B2(n271), .ZN(n576)
         );
  INV_X1 U528 ( .A(n576), .ZN(n896) );
  AOI22_X1 U529 ( .A1(n294), .A2(n577), .B1(add_r3[24]), .B2(n271), .ZN(n578)
         );
  INV_X1 U530 ( .A(n578), .ZN(n895) );
  AOI22_X1 U531 ( .A1(n297), .A2(n579), .B1(add_r3[23]), .B2(n271), .ZN(n580)
         );
  INV_X1 U532 ( .A(n580), .ZN(n894) );
  AOI22_X1 U533 ( .A1(n297), .A2(n581), .B1(add_r3[22]), .B2(n271), .ZN(n582)
         );
  INV_X1 U534 ( .A(n582), .ZN(n893) );
  AOI22_X1 U535 ( .A1(n297), .A2(f3[21]), .B1(add_r3[21]), .B2(n271), .ZN(n583) );
  INV_X1 U536 ( .A(n583), .ZN(n892) );
  AOI22_X1 U537 ( .A1(n297), .A2(f3[20]), .B1(add_r3[20]), .B2(n271), .ZN(n584) );
  INV_X1 U538 ( .A(n584), .ZN(n891) );
  AOI22_X1 U539 ( .A1(n297), .A2(f3[19]), .B1(add_r3[19]), .B2(n271), .ZN(n585) );
  INV_X1 U540 ( .A(n585), .ZN(n890) );
  AOI22_X1 U541 ( .A1(n297), .A2(f3[18]), .B1(add_r3[18]), .B2(n270), .ZN(n586) );
  INV_X1 U542 ( .A(n586), .ZN(n889) );
  AOI22_X1 U543 ( .A1(n297), .A2(f3[17]), .B1(add_r3[17]), .B2(n270), .ZN(n587) );
  INV_X1 U544 ( .A(n587), .ZN(n888) );
  AOI22_X1 U545 ( .A1(n297), .A2(f3[16]), .B1(add_r3[16]), .B2(n270), .ZN(n588) );
  INV_X1 U546 ( .A(n588), .ZN(n887) );
  AOI22_X1 U547 ( .A1(n297), .A2(f3[15]), .B1(add_r3[15]), .B2(n265), .ZN(n589) );
  INV_X1 U548 ( .A(n589), .ZN(n886) );
  AOI22_X1 U549 ( .A1(n297), .A2(f3[14]), .B1(add_r3[14]), .B2(n232), .ZN(n590) );
  INV_X1 U550 ( .A(n590), .ZN(n885) );
  AOI22_X1 U551 ( .A1(n297), .A2(f3[13]), .B1(add_r3[13]), .B2(n232), .ZN(n591) );
  INV_X1 U552 ( .A(n591), .ZN(n884) );
  AOI22_X1 U553 ( .A1(n297), .A2(f3[12]), .B1(add_r3[12]), .B2(n232), .ZN(n592) );
  INV_X1 U554 ( .A(n592), .ZN(n883) );
  AOI22_X1 U555 ( .A1(n298), .A2(f3[11]), .B1(add_r3[11]), .B2(n232), .ZN(n593) );
  INV_X1 U556 ( .A(n593), .ZN(n882) );
  AOI22_X1 U557 ( .A1(n298), .A2(f3[10]), .B1(add_r3[10]), .B2(n232), .ZN(n594) );
  INV_X1 U558 ( .A(n594), .ZN(n881) );
  AOI22_X1 U559 ( .A1(n298), .A2(f3[9]), .B1(add_r3[9]), .B2(n232), .ZN(n595)
         );
  INV_X1 U560 ( .A(n595), .ZN(n880) );
  AOI22_X1 U561 ( .A1(n298), .A2(f3[7]), .B1(add_r3[7]), .B2(n232), .ZN(n596)
         );
  INV_X1 U562 ( .A(n596), .ZN(n878) );
  AOI22_X1 U563 ( .A1(n298), .A2(f3[6]), .B1(add_r3[6]), .B2(n232), .ZN(n597)
         );
  INV_X1 U564 ( .A(n597), .ZN(n877) );
  AOI22_X1 U565 ( .A1(n298), .A2(f3[5]), .B1(add_r3[5]), .B2(n232), .ZN(n598)
         );
  INV_X1 U566 ( .A(n598), .ZN(n876) );
  AOI22_X1 U567 ( .A1(n298), .A2(f3[4]), .B1(add_r3[4]), .B2(n232), .ZN(n599)
         );
  INV_X1 U568 ( .A(n599), .ZN(n875) );
  AOI22_X1 U569 ( .A1(n298), .A2(f3[3]), .B1(add_r3[3]), .B2(n265), .ZN(n600)
         );
  INV_X1 U570 ( .A(n600), .ZN(n874) );
  AOI22_X1 U571 ( .A1(n298), .A2(f3[2]), .B1(add_r3[2]), .B2(n232), .ZN(n601)
         );
  INV_X1 U572 ( .A(n601), .ZN(n873) );
  AOI22_X1 U573 ( .A1(n298), .A2(f3[1]), .B1(add_r3[1]), .B2(n265), .ZN(n602)
         );
  INV_X1 U574 ( .A(n602), .ZN(n872) );
  AOI22_X1 U575 ( .A1(n298), .A2(f3[0]), .B1(add_r3[0]), .B2(n232), .ZN(n603)
         );
  INV_X1 U576 ( .A(n603), .ZN(n871) );
  AOI22_X1 U577 ( .A1(n298), .A2(f3[8]), .B1(add_r3[8]), .B2(n265), .ZN(n604)
         );
  INV_X1 U578 ( .A(n604), .ZN(n879) );
  AOI22_X1 U579 ( .A1(n301), .A2(f5[31]), .B1(add_r5[31]), .B2(n268), .ZN(n605) );
  INV_X1 U580 ( .A(n605), .ZN(n838) );
  AOI22_X1 U581 ( .A1(n301), .A2(f5[30]), .B1(add_r5[30]), .B2(n268), .ZN(n606) );
  INV_X1 U582 ( .A(n606), .ZN(n837) );
  AOI22_X1 U583 ( .A1(n301), .A2(f5[29]), .B1(add_r5[29]), .B2(n268), .ZN(n607) );
  INV_X1 U584 ( .A(n607), .ZN(n836) );
  AOI22_X1 U585 ( .A1(n301), .A2(f5[28]), .B1(add_r5[28]), .B2(n266), .ZN(n608) );
  INV_X1 U586 ( .A(n608), .ZN(n835) );
  AOI22_X1 U587 ( .A1(n301), .A2(f5[27]), .B1(add_r5[27]), .B2(n268), .ZN(n609) );
  INV_X1 U588 ( .A(n609), .ZN(n834) );
  AOI22_X1 U589 ( .A1(n301), .A2(n610), .B1(add_r5[26]), .B2(n268), .ZN(n611)
         );
  INV_X1 U590 ( .A(n611), .ZN(n833) );
  AOI22_X1 U591 ( .A1(n301), .A2(f5[25]), .B1(add_r5[25]), .B2(n268), .ZN(n612) );
  INV_X1 U592 ( .A(n612), .ZN(n832) );
  AOI22_X1 U593 ( .A1(n301), .A2(f5[24]), .B1(add_r5[24]), .B2(n268), .ZN(n613) );
  INV_X1 U594 ( .A(n613), .ZN(n831) );
  AOI22_X1 U595 ( .A1(n301), .A2(f5[23]), .B1(add_r5[23]), .B2(n268), .ZN(n614) );
  INV_X1 U596 ( .A(n614), .ZN(n830) );
  AOI22_X1 U597 ( .A1(n301), .A2(n615), .B1(add_r5[22]), .B2(n268), .ZN(n616)
         );
  INV_X1 U598 ( .A(n616), .ZN(n829) );
  AOI22_X1 U599 ( .A1(n301), .A2(f5[21]), .B1(add_r5[21]), .B2(n269), .ZN(n617) );
  INV_X1 U600 ( .A(n617), .ZN(n828) );
  AOI22_X1 U601 ( .A1(n301), .A2(f5[20]), .B1(add_r5[20]), .B2(n269), .ZN(n618) );
  INV_X1 U602 ( .A(n618), .ZN(n827) );
  AOI22_X1 U603 ( .A1(n302), .A2(f5[19]), .B1(add_r5[19]), .B2(n269), .ZN(n619) );
  INV_X1 U604 ( .A(n619), .ZN(n826) );
  AOI22_X1 U605 ( .A1(n302), .A2(f5[18]), .B1(add_r5[18]), .B2(n269), .ZN(n620) );
  INV_X1 U606 ( .A(n620), .ZN(n825) );
  AOI22_X1 U607 ( .A1(n302), .A2(f5[17]), .B1(add_r5[17]), .B2(n269), .ZN(n621) );
  INV_X1 U608 ( .A(n621), .ZN(n824) );
  AOI22_X1 U609 ( .A1(n302), .A2(f5[16]), .B1(add_r5[16]), .B2(n269), .ZN(n622) );
  INV_X1 U610 ( .A(n622), .ZN(n823) );
  AOI22_X1 U611 ( .A1(n302), .A2(f5[15]), .B1(add_r5[15]), .B2(n269), .ZN(n623) );
  INV_X1 U612 ( .A(n623), .ZN(n822) );
  AOI22_X1 U613 ( .A1(n302), .A2(f5[14]), .B1(add_r5[14]), .B2(n269), .ZN(n624) );
  INV_X1 U614 ( .A(n624), .ZN(n821) );
  AOI22_X1 U615 ( .A1(n302), .A2(f5[13]), .B1(add_r5[13]), .B2(n269), .ZN(n625) );
  INV_X1 U616 ( .A(n625), .ZN(n820) );
  AOI22_X1 U617 ( .A1(n302), .A2(f5[12]), .B1(add_r5[12]), .B2(n269), .ZN(n626) );
  INV_X1 U618 ( .A(n626), .ZN(n819) );
  AOI22_X1 U619 ( .A1(n302), .A2(f5[11]), .B1(add_r5[11]), .B2(n269), .ZN(n627) );
  INV_X1 U620 ( .A(n627), .ZN(n818) );
  AOI22_X1 U621 ( .A1(n302), .A2(f5[10]), .B1(add_r5[10]), .B2(n269), .ZN(n628) );
  INV_X1 U622 ( .A(n628), .ZN(n817) );
  AOI22_X1 U623 ( .A1(n302), .A2(f5[9]), .B1(add_r5[9]), .B2(n270), .ZN(n629)
         );
  INV_X1 U624 ( .A(n629), .ZN(n816) );
  AOI22_X1 U625 ( .A1(n302), .A2(f5[7]), .B1(add_r5[7]), .B2(n270), .ZN(n630)
         );
  INV_X1 U626 ( .A(n630), .ZN(n814) );
  AOI22_X1 U627 ( .A1(n305), .A2(f5[6]), .B1(add_r5[6]), .B2(n270), .ZN(n631)
         );
  INV_X1 U628 ( .A(n631), .ZN(n813) );
  AOI22_X1 U629 ( .A1(n305), .A2(f5[5]), .B1(add_r5[5]), .B2(n270), .ZN(n632)
         );
  INV_X1 U630 ( .A(n632), .ZN(n812) );
  AOI22_X1 U631 ( .A1(n305), .A2(f5[4]), .B1(add_r5[4]), .B2(n270), .ZN(n633)
         );
  INV_X1 U632 ( .A(n633), .ZN(n811) );
  AOI22_X1 U633 ( .A1(n305), .A2(f5[3]), .B1(add_r5[3]), .B2(n270), .ZN(n634)
         );
  INV_X1 U634 ( .A(n634), .ZN(n810) );
  AOI22_X1 U635 ( .A1(n305), .A2(f5[2]), .B1(add_r5[2]), .B2(n270), .ZN(n635)
         );
  INV_X1 U636 ( .A(n635), .ZN(n809) );
  AOI22_X1 U637 ( .A1(n305), .A2(f5[1]), .B1(add_r5[1]), .B2(n270), .ZN(n636)
         );
  INV_X1 U638 ( .A(n636), .ZN(n808) );
  AOI22_X1 U639 ( .A1(n305), .A2(f5[0]), .B1(add_r5[0]), .B2(n265), .ZN(n637)
         );
  INV_X1 U640 ( .A(n637), .ZN(n807) );
  AOI22_X1 U641 ( .A1(n305), .A2(f5[8]), .B1(add_r5[8]), .B2(n268), .ZN(n638)
         );
  INV_X1 U642 ( .A(n638), .ZN(n815) );
  AOI22_X1 U643 ( .A1(n305), .A2(f2[31]), .B1(add_r2[31]), .B2(n268), .ZN(n639) );
  INV_X1 U644 ( .A(n639), .ZN(n934) );
  AOI22_X1 U645 ( .A1(n305), .A2(f2[30]), .B1(add_r2[30]), .B2(n268), .ZN(n640) );
  INV_X1 U646 ( .A(n640), .ZN(n933) );
  AOI22_X1 U647 ( .A1(n305), .A2(f2[29]), .B1(add_r2[29]), .B2(n267), .ZN(n641) );
  INV_X1 U648 ( .A(n641), .ZN(n932) );
  AOI22_X1 U649 ( .A1(n305), .A2(f2[28]), .B1(add_r2[28]), .B2(n267), .ZN(n642) );
  INV_X1 U650 ( .A(n642), .ZN(n931) );
  AOI22_X1 U651 ( .A1(n306), .A2(n643), .B1(add_r2[27]), .B2(n267), .ZN(n644)
         );
  INV_X1 U652 ( .A(n644), .ZN(n930) );
  AOI22_X1 U653 ( .A1(n306), .A2(n645), .B1(add_r2[26]), .B2(n267), .ZN(n646)
         );
  INV_X1 U654 ( .A(n646), .ZN(n929) );
  AOI22_X1 U655 ( .A1(n306), .A2(n647), .B1(add_r2[25]), .B2(n267), .ZN(n648)
         );
  INV_X1 U656 ( .A(n648), .ZN(n928) );
  AOI22_X1 U657 ( .A1(n306), .A2(f2[24]), .B1(add_r2[24]), .B2(n267), .ZN(n649) );
  INV_X1 U658 ( .A(n649), .ZN(n927) );
  AOI22_X1 U659 ( .A1(n306), .A2(n650), .B1(add_r2[23]), .B2(n267), .ZN(n651)
         );
  INV_X1 U660 ( .A(n651), .ZN(n926) );
  AOI22_X1 U661 ( .A1(n306), .A2(n652), .B1(add_r2[22]), .B2(n267), .ZN(n653)
         );
  INV_X1 U662 ( .A(n653), .ZN(n925) );
  AOI22_X1 U663 ( .A1(n306), .A2(n654), .B1(add_r2[21]), .B2(n267), .ZN(n655)
         );
  INV_X1 U664 ( .A(n655), .ZN(n924) );
  AOI22_X1 U665 ( .A1(n306), .A2(n656), .B1(add_r2[20]), .B2(n267), .ZN(n657)
         );
  INV_X1 U666 ( .A(n657), .ZN(n923) );
  AOI22_X1 U667 ( .A1(n306), .A2(n658), .B1(add_r2[19]), .B2(n267), .ZN(n659)
         );
  INV_X1 U668 ( .A(n659), .ZN(n922) );
  AOI22_X1 U669 ( .A1(n306), .A2(n660), .B1(add_r2[18]), .B2(n267), .ZN(n661)
         );
  INV_X1 U670 ( .A(n661), .ZN(n921) );
  AOI22_X1 U671 ( .A1(n306), .A2(n662), .B1(add_r2[17]), .B2(n266), .ZN(n663)
         );
  INV_X1 U672 ( .A(n663), .ZN(n920) );
  AOI22_X1 U673 ( .A1(n306), .A2(f2[16]), .B1(add_r2[16]), .B2(n266), .ZN(n664) );
  INV_X1 U674 ( .A(n664), .ZN(n919) );
  AOI22_X1 U675 ( .A1(n309), .A2(f2[15]), .B1(add_r2[15]), .B2(n266), .ZN(n665) );
  INV_X1 U676 ( .A(n665), .ZN(n918) );
  AOI22_X1 U677 ( .A1(n309), .A2(f2[14]), .B1(add_r2[14]), .B2(n266), .ZN(n666) );
  INV_X1 U678 ( .A(n666), .ZN(n917) );
  AOI22_X1 U679 ( .A1(n309), .A2(f2[13]), .B1(add_r2[13]), .B2(n266), .ZN(n667) );
  INV_X1 U680 ( .A(n667), .ZN(n916) );
  AOI22_X1 U681 ( .A1(n309), .A2(f2[12]), .B1(add_r2[12]), .B2(n266), .ZN(n668) );
  INV_X1 U682 ( .A(n668), .ZN(n915) );
  AOI22_X1 U683 ( .A1(n309), .A2(f2[11]), .B1(add_r2[11]), .B2(n266), .ZN(n669) );
  INV_X1 U684 ( .A(n669), .ZN(n914) );
  AOI22_X1 U685 ( .A1(n309), .A2(f2[10]), .B1(add_r2[10]), .B2(n266), .ZN(n670) );
  INV_X1 U686 ( .A(n670), .ZN(n913) );
  AOI22_X1 U687 ( .A1(n309), .A2(f2[9]), .B1(add_r2[9]), .B2(n266), .ZN(n671)
         );
  INV_X1 U688 ( .A(n671), .ZN(n912) );
  AOI22_X1 U689 ( .A1(n309), .A2(f2[7]), .B1(add_r2[7]), .B2(n266), .ZN(n672)
         );
  INV_X1 U690 ( .A(n672), .ZN(n910) );
  AOI22_X1 U691 ( .A1(n309), .A2(f2[6]), .B1(add_r2[6]), .B2(n266), .ZN(n673)
         );
  INV_X1 U692 ( .A(n673), .ZN(n909) );
  AOI22_X1 U693 ( .A1(n309), .A2(f2[5]), .B1(add_r2[5]), .B2(n265), .ZN(n674)
         );
  INV_X1 U694 ( .A(n674), .ZN(n908) );
  AOI22_X1 U695 ( .A1(n309), .A2(f2[4]), .B1(add_r2[4]), .B2(n265), .ZN(n675)
         );
  INV_X1 U696 ( .A(n675), .ZN(n907) );
  AOI22_X1 U697 ( .A1(n309), .A2(f2[3]), .B1(add_r2[3]), .B2(n265), .ZN(n676)
         );
  INV_X1 U698 ( .A(n676), .ZN(n906) );
  AOI22_X1 U699 ( .A1(n302), .A2(f2[2]), .B1(add_r2[2]), .B2(n265), .ZN(n677)
         );
  INV_X1 U700 ( .A(n677), .ZN(n905) );
  AOI22_X1 U701 ( .A1(n301), .A2(f2[1]), .B1(add_r2[1]), .B2(n265), .ZN(n678)
         );
  INV_X1 U702 ( .A(n678), .ZN(n904) );
  AOI22_X1 U703 ( .A1(n298), .A2(f2[0]), .B1(add_r2[0]), .B2(n265), .ZN(n967)
         );
  INV_X1 U704 ( .A(n967), .ZN(n903) );
  AOI22_X1 U705 ( .A1(n309), .A2(f2[8]), .B1(add_r2[8]), .B2(n270), .ZN(n969)
         );
  INV_X1 U706 ( .A(n969), .ZN(n911) );
  INV_X1 U707 ( .A(n286), .ZN(n1062) );
  OAI222_X1 U708 ( .A1(n1060), .A2(n38), .B1(n1059), .B2(n970), .C1(n206), 
        .C2(n192), .ZN(n971) );
  AOI221_X1 U709 ( .B1(f7[8]), .B2(n1062), .C1(f8[8]), .C2(n386), .A(n971), 
        .ZN(n974) );
  OAI22_X1 U710 ( .A1(n382), .A2(n64), .B1(n383), .B2(n160), .ZN(n972) );
  AOI221_X1 U711 ( .B1(f4[8]), .B2(n277), .C1(f3[8]), .C2(n178), .A(n972), 
        .ZN(n973) );
  NAND2_X1 U712 ( .A1(n974), .A2(n973), .ZN(n702) );
  OAI222_X1 U713 ( .A1(n1060), .A2(n39), .B1(n1059), .B2(n975), .C1(n206), 
        .C2(n193), .ZN(n976) );
  AOI221_X1 U714 ( .B1(f7[7]), .B2(n1062), .C1(f8[7]), .C2(n386), .A(n976), 
        .ZN(n979) );
  OAI22_X1 U715 ( .A1(n281), .A2(n65), .B1(n280), .B2(n161), .ZN(n977) );
  AOI221_X1 U716 ( .B1(f4[7]), .B2(n277), .C1(f3[7]), .C2(n178), .A(n977), 
        .ZN(n978) );
  NAND2_X1 U717 ( .A1(n979), .A2(n978), .ZN(n703) );
  OAI222_X1 U718 ( .A1(n1060), .A2(n40), .B1(n1059), .B2(n980), .C1(n285), 
        .C2(n194), .ZN(n981) );
  AOI221_X1 U719 ( .B1(f7[6]), .B2(n1062), .C1(f8[6]), .C2(n276), .A(n981), 
        .ZN(n984) );
  OAI22_X1 U720 ( .A1(n382), .A2(n66), .B1(n383), .B2(n162), .ZN(n982) );
  AOI221_X1 U721 ( .B1(f4[6]), .B2(n277), .C1(f3[6]), .C2(n178), .A(n982), 
        .ZN(n983) );
  NAND2_X1 U722 ( .A1(n984), .A2(n983), .ZN(n704) );
  OAI222_X1 U723 ( .A1(n1060), .A2(n96), .B1(n1059), .B2(n985), .C1(n206), 
        .C2(n195), .ZN(n986) );
  AOI221_X1 U724 ( .B1(f7[5]), .B2(n1062), .C1(f8[5]), .C2(n276), .A(n986), 
        .ZN(n989) );
  OAI22_X1 U725 ( .A1(n382), .A2(n67), .B1(n383), .B2(n163), .ZN(n987) );
  AOI221_X1 U726 ( .B1(f4[5]), .B2(n277), .C1(f3[5]), .C2(n178), .A(n987), 
        .ZN(n988) );
  NAND2_X1 U727 ( .A1(n989), .A2(n988), .ZN(n705) );
  OAI222_X1 U728 ( .A1(n1060), .A2(n97), .B1(n1059), .B2(n990), .C1(n285), 
        .C2(n196), .ZN(n991) );
  AOI221_X1 U729 ( .B1(f7[4]), .B2(n1062), .C1(f8[4]), .C2(n276), .A(n991), 
        .ZN(n994) );
  OAI22_X1 U730 ( .A1(n382), .A2(n68), .B1(n383), .B2(n164), .ZN(n992) );
  AOI221_X1 U731 ( .B1(f4[4]), .B2(n277), .C1(f3[4]), .C2(n178), .A(n992), 
        .ZN(n993) );
  NAND2_X1 U732 ( .A1(n994), .A2(n993), .ZN(n706) );
  OAI222_X1 U733 ( .A1(n1060), .A2(n98), .B1(n1059), .B2(n995), .C1(n206), 
        .C2(n197), .ZN(n996) );
  AOI221_X1 U734 ( .B1(f7[3]), .B2(n1062), .C1(f8[3]), .C2(n276), .A(n996), 
        .ZN(n999) );
  OAI22_X1 U735 ( .A1(n382), .A2(n69), .B1(n383), .B2(n165), .ZN(n997) );
  AOI221_X1 U736 ( .B1(f4[3]), .B2(n277), .C1(f3[3]), .C2(n178), .A(n997), 
        .ZN(n998) );
  NAND2_X1 U737 ( .A1(n999), .A2(n998), .ZN(n707) );
  OAI222_X1 U738 ( .A1(n1060), .A2(n99), .B1(n1059), .B2(n1000), .C1(n285), 
        .C2(n198), .ZN(n1001) );
  AOI221_X1 U739 ( .B1(f7[2]), .B2(n1062), .C1(f8[2]), .C2(n276), .A(n1001), 
        .ZN(n1004) );
  OAI22_X1 U740 ( .A1(n382), .A2(n70), .B1(n383), .B2(n166), .ZN(n1002) );
  AOI221_X1 U741 ( .B1(f4[2]), .B2(n277), .C1(f3[2]), .C2(n178), .A(n1002), 
        .ZN(n1003) );
  NAND2_X1 U742 ( .A1(n1004), .A2(n1003), .ZN(n708) );
  OAI222_X1 U743 ( .A1(n1060), .A2(n100), .B1(n1059), .B2(n1005), .C1(n206), 
        .C2(n199), .ZN(n1006) );
  AOI221_X1 U744 ( .B1(f7[1]), .B2(n1062), .C1(f8[1]), .C2(n276), .A(n1006), 
        .ZN(n1009) );
  OAI22_X1 U745 ( .A1(n382), .A2(n71), .B1(n383), .B2(n167), .ZN(n1007) );
  AOI221_X1 U746 ( .B1(f4[1]), .B2(n277), .C1(f3[1]), .C2(n178), .A(n1007), 
        .ZN(n1008) );
  NAND2_X1 U747 ( .A1(n1009), .A2(n1008), .ZN(n709) );
  OAI222_X1 U748 ( .A1(n1060), .A2(n101), .B1(n1059), .B2(n1010), .C1(n285), 
        .C2(n200), .ZN(n1011) );
  AOI221_X1 U749 ( .B1(f7[0]), .B2(n1062), .C1(f8[0]), .C2(n276), .A(n1011), 
        .ZN(n1014) );
  OAI22_X1 U750 ( .A1(n382), .A2(n72), .B1(n383), .B2(n168), .ZN(n1012) );
  AOI221_X1 U751 ( .B1(f4[0]), .B2(n277), .C1(f3[0]), .C2(n178), .A(n1012), 
        .ZN(n1013) );
  NAND2_X1 U752 ( .A1(n1014), .A2(n1013), .ZN(n710) );
  INV_X1 U753 ( .A(n1060), .ZN(n1066) );
  INV_X1 U754 ( .A(n285), .ZN(n1063) );
  OAI22_X1 U755 ( .A1(n1060), .A2(n14), .B1(n1059), .B2(n1015), .ZN(n1016) );
  AOI221_X1 U756 ( .B1(f6[20]), .B2(n1063), .C1(n1017), .C2(n1062), .A(n1016), 
        .ZN(n327) );
  OAI222_X1 U757 ( .A1(n383), .A2(n148), .B1(n384), .B2(n84), .C1(n382), .C2(
        n52), .ZN(n1018) );
  AOI221_X1 U758 ( .B1(f4[20]), .B2(n277), .C1(f8[20]), .C2(n276), .A(n1018), 
        .ZN(n328) );
  OAI22_X1 U759 ( .A1(n1060), .A2(n15), .B1(n1059), .B2(n1019), .ZN(n1020) );
  AOI221_X1 U760 ( .B1(f6[21]), .B2(n1063), .C1(n1021), .C2(n1062), .A(n1020), 
        .ZN(n323) );
  OAI222_X1 U761 ( .A1(n383), .A2(n147), .B1(n384), .B2(n83), .C1(n382), .C2(
        n51), .ZN(n1022) );
  AOI221_X1 U762 ( .B1(f4[21]), .B2(n277), .C1(f8[21]), .C2(n276), .A(n1022), 
        .ZN(n324) );
  OAI22_X1 U763 ( .A1(n1060), .A2(n17), .B1(n1059), .B2(n1023), .ZN(n1024) );
  AOI221_X1 U764 ( .B1(f6[22]), .B2(n1063), .C1(n1025), .C2(n1062), .A(n1024), 
        .ZN(n319) );
  OAI222_X1 U765 ( .A1(n383), .A2(n146), .B1(n384), .B2(n82), .C1(n382), .C2(
        n50), .ZN(n1026) );
  AOI221_X1 U766 ( .B1(f4[22]), .B2(n277), .C1(f8[22]), .C2(n276), .A(n1026), 
        .ZN(n320) );
  OAI22_X1 U767 ( .A1(n1060), .A2(n18), .B1(n1059), .B2(n1027), .ZN(n1028) );
  AOI221_X1 U768 ( .B1(f6[23]), .B2(n1063), .C1(n1029), .C2(n1062), .A(n1028), 
        .ZN(n315) );
  OAI222_X1 U769 ( .A1(n383), .A2(n145), .B1(n384), .B2(n81), .C1(n382), .C2(
        n49), .ZN(n1030) );
  AOI221_X1 U770 ( .B1(f4[23]), .B2(n277), .C1(f8[23]), .C2(n276), .A(n1030), 
        .ZN(n316) );
  OAI22_X1 U771 ( .A1(n1060), .A2(n19), .B1(n1059), .B2(n16), .ZN(n1031) );
  AOI221_X1 U772 ( .B1(f6[24]), .B2(n1063), .C1(n1032), .C2(n1062), .A(n1031), 
        .ZN(n311) );
  OAI222_X1 U773 ( .A1(n383), .A2(n144), .B1(n384), .B2(n80), .C1(n382), .C2(
        n48), .ZN(n1033) );
  AOI221_X1 U774 ( .B1(f4[24]), .B2(n277), .C1(f8[24]), .C2(n276), .A(n1033), 
        .ZN(n312) );
  OAI22_X1 U775 ( .A1(n1060), .A2(n20), .B1(n1059), .B2(n1034), .ZN(n1035) );
  AOI221_X1 U776 ( .B1(n1036), .B2(n1063), .C1(f7[25]), .C2(n1062), .A(n1035), 
        .ZN(n307) );
  OAI222_X1 U777 ( .A1(n383), .A2(n143), .B1(n384), .B2(n79), .C1(n382), .C2(
        n47), .ZN(n1037) );
  AOI221_X1 U778 ( .B1(f4[25]), .B2(n277), .C1(f8[25]), .C2(n276), .A(n1037), 
        .ZN(n308) );
  OAI22_X1 U779 ( .A1(n1060), .A2(n32), .B1(n1059), .B2(n1038), .ZN(n1039) );
  AOI221_X1 U780 ( .B1(n1040), .B2(n1063), .C1(f7[26]), .C2(n1062), .A(n1039), 
        .ZN(n303) );
  OAI222_X1 U781 ( .A1(n383), .A2(n142), .B1(n384), .B2(n78), .C1(n382), .C2(
        n46), .ZN(n1041) );
  AOI221_X1 U782 ( .B1(f4[26]), .B2(n277), .C1(f8[26]), .C2(n276), .A(n1041), 
        .ZN(n304) );
  OAI22_X1 U783 ( .A1(n1060), .A2(n33), .B1(n1059), .B2(n1042), .ZN(n1043) );
  AOI221_X1 U784 ( .B1(n1044), .B2(n1063), .C1(f7[27]), .C2(n1062), .A(n1043), 
        .ZN(n299) );
  OAI222_X1 U785 ( .A1(n383), .A2(n141), .B1(n384), .B2(n77), .C1(n382), .C2(
        n45), .ZN(n1045) );
  AOI221_X1 U786 ( .B1(f4[27]), .B2(n277), .C1(f8[27]), .C2(n276), .A(n1045), 
        .ZN(n300) );
  OAI22_X1 U787 ( .A1(n1060), .A2(n34), .B1(n1059), .B2(n1046), .ZN(n1047) );
  AOI221_X1 U788 ( .B1(n1048), .B2(n1063), .C1(f7[28]), .C2(n1062), .A(n1047), 
        .ZN(n295) );
  OAI222_X1 U789 ( .A1(n383), .A2(n140), .B1(n384), .B2(n76), .C1(n382), .C2(
        n44), .ZN(n1049) );
  AOI221_X1 U790 ( .B1(f4[28]), .B2(n277), .C1(f8[28]), .C2(n276), .A(n1049), 
        .ZN(n296) );
  OAI22_X1 U791 ( .A1(n1060), .A2(n35), .B1(n1059), .B2(n1050), .ZN(n1051) );
  AOI221_X1 U792 ( .B1(n1052), .B2(n1063), .C1(f7[29]), .C2(n1062), .A(n1051), 
        .ZN(n291) );
  OAI222_X1 U793 ( .A1(n383), .A2(n139), .B1(n384), .B2(n75), .C1(n382), .C2(
        n43), .ZN(n1053) );
  AOI221_X1 U794 ( .B1(f4[29]), .B2(n277), .C1(f8[29]), .C2(n276), .A(n1053), 
        .ZN(n292) );
  OAI22_X1 U795 ( .A1(n1060), .A2(n36), .B1(n1059), .B2(n1054), .ZN(n1055) );
  AOI221_X1 U796 ( .B1(n1056), .B2(n1063), .C1(f7[30]), .C2(n1062), .A(n1055), 
        .ZN(n287) );
  OAI222_X1 U797 ( .A1(n383), .A2(n138), .B1(n384), .B2(n74), .C1(n382), .C2(
        n42), .ZN(n1057) );
  AOI221_X1 U798 ( .B1(f4[30]), .B2(n277), .C1(f8[30]), .C2(n276), .A(n1057), 
        .ZN(n288) );
  OAI22_X1 U799 ( .A1(n1060), .A2(n37), .B1(n1059), .B2(n1058), .ZN(n1061) );
  AOI221_X1 U800 ( .B1(n1064), .B2(n1063), .C1(f7[31]), .C2(n1062), .A(n1061), 
        .ZN(n274) );
  OAI222_X1 U801 ( .A1(n383), .A2(n137), .B1(n384), .B2(n73), .C1(n382), .C2(
        n41), .ZN(n1065) );
  AOI221_X1 U802 ( .B1(f4[31]), .B2(n385), .C1(f8[31]), .C2(n386), .A(n1065), 
        .ZN(n275) );
endmodule


module ctrlpath ( clk, reset, start, addr_x, wr_en_x, addr_a1, addr_a2, 
        addr_a3, addr_a4, addr_a5, addr_a6, addr_a7, addr_a8, wr_en_a1, 
        wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6, wr_en_a7, wr_en_a8, 
        clear_acc, clc, clc1, addr_y, wr_en_y, done, loadMatrix, loadVector );
  output [2:0] addr_x;
  output [2:0] addr_a1;
  output [2:0] addr_a2;
  output [2:0] addr_a3;
  output [2:0] addr_a4;
  output [2:0] addr_a5;
  output [2:0] addr_a6;
  output [2:0] addr_a7;
  output [2:0] addr_a8;
  output [2:0] addr_y;
  input clk, reset, start, loadMatrix, loadVector;
  output wr_en_x, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6,
         wr_en_a7, wr_en_a8, clear_acc, clc, clc1, wr_en_y, done;
  wire   N32, N33, N34, N35, N37, N45, N46, N56, N57, N67, N68, N78, N79, N89,
         N90, N100, N101, N111, N112, N122, N123, N131, N132, N133, N141, N142,
         N143, N146, N147, N148, n76, n79, n80, n81, n83, n84, n85, n86, n87,
         n88, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n111, n112, n113, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39;
  wire   [4:0] state;

  DFF_X1 \state_reg[3]  ( .D(N35), .CK(clk), .Q(state[3]) );
  DFF_X1 done_reg ( .D(N37), .CK(clk), .Q(done) );
  DFF_X1 \addr_x_reg[0]  ( .D(N131), .CK(clk), .Q(addr_x[0]) );
  DFF_X1 \addr_x_reg[1]  ( .D(N132), .CK(clk), .Q(addr_x[1]) );
  DFF_X1 clear_acc_reg ( .D(N146), .CK(clk), .Q(clear_acc) );
  DFF_X1 clc_reg ( .D(N147), .CK(clk), .Q(clc) );
  DFF_X1 clc1_reg ( .D(N148), .CK(clk), .Q(clc1) );
  NAND3_X1 U201 ( .A1(n127), .A2(n97), .A3(addr_a5[0]), .ZN(n129) );
  NAND3_X1 U202 ( .A1(n133), .A2(n121), .A3(n134), .ZN(n132) );
  NAND3_X1 U203 ( .A1(n137), .A2(n94), .A3(addr_a4[0]), .ZN(n139) );
  NAND3_X1 U204 ( .A1(n120), .A2(n119), .A3(n142), .ZN(n141) );
  NAND3_X1 U205 ( .A1(n145), .A2(n91), .A3(addr_a3[0]), .ZN(n147) );
  NAND3_X1 U206 ( .A1(n142), .A2(n120), .A3(n27), .ZN(n149) );
  NAND3_X1 U207 ( .A1(n153), .A2(n87), .A3(addr_a2[0]), .ZN(n155) );
  NAND3_X1 U208 ( .A1(n119), .A2(n118), .A3(n142), .ZN(n157) );
  NAND3_X1 U209 ( .A1(n162), .A2(n84), .A3(addr_a1[0]), .ZN(n164) );
  NAND3_X1 U210 ( .A1(n133), .A2(n167), .A3(n134), .ZN(n166) );
  NAND3_X1 U211 ( .A1(n178), .A2(n179), .A3(n31), .ZN(n175) );
  NAND3_X1 U212 ( .A1(addr_a8[1]), .A2(addr_a8[0]), .A3(addr_a8[2]), .ZN(n170)
         );
  NAND3_X1 U213 ( .A1(addr_a7[1]), .A2(addr_a7[0]), .A3(addr_a7[2]), .ZN(n195)
         );
  NAND3_X1 U214 ( .A1(addr_y[0]), .A2(n112), .A3(n216), .ZN(n218) );
  NAND3_X1 U215 ( .A1(n219), .A2(n30), .A3(addr_y[0]), .ZN(n220) );
  NAND3_X1 U216 ( .A1(addr_x[0]), .A2(n224), .A3(addr_x[1]), .ZN(n223) );
  NAND3_X1 U217 ( .A1(n228), .A2(n106), .A3(addr_a8[0]), .ZN(n230) );
  NAND3_X1 U218 ( .A1(n233), .A2(n172), .A3(n134), .ZN(n232) );
  NAND3_X1 U219 ( .A1(n236), .A2(n103), .A3(addr_a7[0]), .ZN(n238) );
  NAND3_X1 U220 ( .A1(n233), .A2(n173), .A3(n134), .ZN(n240) );
  NAND3_X1 U221 ( .A1(n123), .A2(n100), .A3(addr_a6[0]), .ZN(n244) );
  NAND3_X1 U222 ( .A1(n22), .A2(n158), .A3(n28), .ZN(n245) );
  NAND3_X1 U223 ( .A1(n119), .A2(n118), .A3(n120), .ZN(n246) );
  NAND3_X1 U224 ( .A1(addr_x[1]), .A2(addr_x[0]), .A3(addr_x[2]), .ZN(n205) );
  DFF_X1 \state_reg[4]  ( .D(n21), .CK(clk), .Q(state[4]), .QN(n76) );
  DFF_X1 \state_reg[2]  ( .D(N34), .CK(clk), .Q(state[2]), .QN(n79) );
  DFF_X1 \addr_y_reg[0]  ( .D(N141), .CK(clk), .Q(addr_y[0]), .QN(n113) );
  DFF_X1 \addr_y_reg[1]  ( .D(N142), .CK(clk), .Q(addr_y[1]), .QN(n112) );
  DFF_X1 \state_reg[1]  ( .D(N33), .CK(clk), .Q(state[1]), .QN(n80) );
  DFF_X1 \addr_y_reg[2]  ( .D(N143), .CK(clk), .Q(addr_y[2]), .QN(n111) );
  DFF_X1 \state_reg[0]  ( .D(N32), .CK(clk), .Q(state[0]), .QN(n81) );
  DFF_X1 \addr_x_reg[2]  ( .D(N133), .CK(clk), .Q(addr_x[2]), .QN(n108) );
  DFF_X1 \addr_a8_reg[0]  ( .D(n8), .CK(clk), .Q(addr_a8[0]), .QN(n107) );
  DFF_X1 \addr_a7_reg[0]  ( .D(n6), .CK(clk), .Q(addr_a7[0]), .QN(n104) );
  DFF_X1 \addr_a6_reg[0]  ( .D(n5), .CK(clk), .Q(addr_a6[0]), .QN(n101) );
  DFF_X1 \addr_a5_reg[0]  ( .D(n19), .CK(clk), .Q(addr_a5[0]), .QN(n98) );
  DFF_X1 \addr_a4_reg[0]  ( .D(n17), .CK(clk), .Q(addr_a4[0]), .QN(n95) );
  DFF_X1 \addr_a3_reg[0]  ( .D(n15), .CK(clk), .Q(addr_a3[0]), .QN(n92) );
  DFF_X1 \addr_a2_reg[0]  ( .D(n13), .CK(clk), .Q(addr_a2[0]), .QN(n88) );
  DFF_X1 \addr_a1_reg[0]  ( .D(n11), .CK(clk), .Q(addr_a1[0]), .QN(n85) );
  DFF_X1 \addr_a8_reg[1]  ( .D(N122), .CK(clk), .Q(addr_a8[1]), .QN(n106) );
  DFF_X1 \addr_a7_reg[1]  ( .D(N111), .CK(clk), .Q(addr_a7[1]), .QN(n103) );
  DFF_X1 \addr_a6_reg[1]  ( .D(N100), .CK(clk), .Q(addr_a6[1]), .QN(n100) );
  DFF_X1 \addr_a5_reg[1]  ( .D(N89), .CK(clk), .Q(addr_a5[1]), .QN(n97) );
  DFF_X1 \addr_a4_reg[1]  ( .D(N78), .CK(clk), .Q(addr_a4[1]), .QN(n94) );
  DFF_X1 \addr_a3_reg[1]  ( .D(N67), .CK(clk), .Q(addr_a3[1]), .QN(n91) );
  DFF_X1 \addr_a2_reg[1]  ( .D(N56), .CK(clk), .Q(addr_a2[1]), .QN(n87) );
  DFF_X1 \addr_a1_reg[1]  ( .D(N45), .CK(clk), .Q(addr_a1[1]), .QN(n84) );
  DFF_X1 \addr_a8_reg[2]  ( .D(N123), .CK(clk), .Q(addr_a8[2]), .QN(n105) );
  DFF_X1 \addr_a7_reg[2]  ( .D(N112), .CK(clk), .Q(addr_a7[2]), .QN(n102) );
  DFF_X1 \addr_a6_reg[2]  ( .D(N101), .CK(clk), .Q(addr_a6[2]), .QN(n99) );
  DFF_X1 \addr_a5_reg[2]  ( .D(N90), .CK(clk), .Q(addr_a5[2]), .QN(n96) );
  DFF_X1 \addr_a4_reg[2]  ( .D(N79), .CK(clk), .Q(addr_a4[2]), .QN(n93) );
  DFF_X1 \addr_a3_reg[2]  ( .D(N68), .CK(clk), .Q(addr_a3[2]), .QN(n90) );
  DFF_X1 \addr_a2_reg[2]  ( .D(N57), .CK(clk), .Q(addr_a2[2]), .QN(n86) );
  DFF_X1 \addr_a1_reg[2]  ( .D(N46), .CK(clk), .Q(addr_a1[2]), .QN(n83) );
  INV_X1 U3 ( .A(n248), .ZN(n22) );
  INV_X1 U4 ( .A(n224), .ZN(n10) );
  INV_X1 U5 ( .A(n246), .ZN(n28) );
  NAND2_X1 U6 ( .A1(n233), .A2(n133), .ZN(n248) );
  NAND2_X1 U7 ( .A1(n131), .A2(n245), .ZN(n123) );
  NAND2_X1 U8 ( .A1(n131), .A2(n149), .ZN(n145) );
  INV_X1 U9 ( .A(n150), .ZN(n27) );
  NAND2_X1 U10 ( .A1(n131), .A2(n157), .ZN(n153) );
  NAND2_X1 U11 ( .A1(n131), .A2(n141), .ZN(n137) );
  NAND2_X1 U12 ( .A1(n131), .A2(n132), .ZN(n127) );
  NAND2_X1 U13 ( .A1(n131), .A2(n166), .ZN(n162) );
  NOR2_X1 U14 ( .A1(n32), .A2(n23), .ZN(n133) );
  OAI21_X1 U15 ( .B1(n37), .B2(n117), .A(n131), .ZN(n224) );
  NAND2_X1 U16 ( .A1(n202), .A2(n116), .ZN(N148) );
  AND2_X1 U17 ( .A1(n207), .A2(n180), .ZN(n191) );
  NAND2_X1 U18 ( .A1(n117), .A2(n180), .ZN(N146) );
  INV_X1 U19 ( .A(n210), .ZN(n29) );
  AND2_X1 U20 ( .A1(n121), .A2(n167), .ZN(n233) );
  AND4_X1 U21 ( .A1(n247), .A2(n178), .A3(n210), .A4(n26), .ZN(n158) );
  INV_X1 U22 ( .A(N148), .ZN(n26) );
  OR2_X1 U23 ( .A1(n189), .A2(N37), .ZN(n188) );
  OAI211_X2 U24 ( .C1(n205), .C2(n210), .A(n116), .B(n178), .ZN(n124) );
  OAI221_X1 U25 ( .B1(n169), .B2(n167), .C1(n121), .C2(n35), .A(n28), .ZN(n177) );
  INV_X1 U26 ( .A(n184), .ZN(n35) );
  AOI21_X1 U27 ( .B1(n251), .B2(n33), .A(n189), .ZN(n178) );
  OAI22_X1 U28 ( .A1(n117), .A2(n205), .B1(n173), .B2(n170), .ZN(n176) );
  NAND4_X1 U29 ( .A1(n202), .A2(n159), .A3(n247), .A4(n249), .ZN(n131) );
  NOR3_X1 U30 ( .A1(n124), .A2(n248), .A3(n246), .ZN(n249) );
  OAI22_X1 U31 ( .A1(n37), .A2(n117), .B1(n172), .B2(n195), .ZN(n192) );
  NAND2_X1 U32 ( .A1(n222), .A2(n252), .ZN(n116) );
  NAND2_X1 U33 ( .A1(n254), .A2(n251), .ZN(n117) );
  OAI21_X1 U34 ( .B1(n119), .B2(n36), .A(n118), .ZN(n150) );
  INV_X1 U35 ( .A(n194), .ZN(n36) );
  OAI21_X1 U36 ( .B1(n190), .B2(n208), .A(n209), .ZN(n183) );
  NAND2_X1 U37 ( .A1(n254), .A2(n252), .ZN(n121) );
  NAND2_X1 U38 ( .A1(n131), .A2(n232), .ZN(n228) );
  NAND2_X1 U39 ( .A1(n131), .A2(n240), .ZN(n236) );
  NAND2_X1 U40 ( .A1(n250), .A2(n252), .ZN(n119) );
  NAND2_X1 U41 ( .A1(n255), .A2(n254), .ZN(n210) );
  NAND2_X1 U42 ( .A1(n255), .A2(n250), .ZN(n167) );
  NAND2_X1 U43 ( .A1(n250), .A2(n251), .ZN(n118) );
  INV_X1 U44 ( .A(n205), .ZN(n37) );
  NAND2_X1 U45 ( .A1(n251), .A2(n222), .ZN(n209) );
  NAND2_X1 U46 ( .A1(n221), .A2(n250), .ZN(n120) );
  INV_X1 U47 ( .A(n216), .ZN(n30) );
  NAND2_X1 U48 ( .A1(n33), .A2(n221), .ZN(n202) );
  INV_X1 U49 ( .A(n212), .ZN(n33) );
  NAND2_X1 U50 ( .A1(n33), .A2(n252), .ZN(n180) );
  NAND2_X1 U51 ( .A1(n255), .A2(n222), .ZN(n208) );
  NOR2_X1 U52 ( .A1(n2), .A2(n116), .ZN(N37) );
  INV_X1 U53 ( .A(n190), .ZN(n2) );
  INV_X1 U54 ( .A(n172), .ZN(n32) );
  NAND2_X1 U55 ( .A1(n221), .A2(n254), .ZN(n207) );
  AND3_X1 U56 ( .A1(n158), .A2(n159), .A3(n28), .ZN(n134) );
  INV_X1 U57 ( .A(n222), .ZN(n34) );
  AND4_X1 U58 ( .A1(n207), .A2(n25), .A3(n209), .A4(n256), .ZN(n247) );
  AND2_X1 U59 ( .A1(n208), .A2(n31), .ZN(n256) );
  INV_X1 U60 ( .A(N146), .ZN(n25) );
  AND3_X1 U61 ( .A1(n158), .A2(n159), .A3(n22), .ZN(n142) );
  INV_X1 U62 ( .A(n193), .ZN(n3) );
  AND2_X1 U63 ( .A1(n221), .A2(n222), .ZN(n189) );
  INV_X1 U64 ( .A(n173), .ZN(n23) );
  INV_X1 U65 ( .A(n168), .ZN(n21) );
  AOI221_X1 U66 ( .B1(n169), .B2(wr_en_a5), .C1(n170), .C2(wr_en_a8), .A(n171), 
        .ZN(n168) );
  OR2_X1 U67 ( .A1(wr_en_a7), .A2(wr_en_a6), .ZN(n171) );
  OAI22_X1 U68 ( .A1(n190), .A2(n116), .B1(n184), .B2(n121), .ZN(n204) );
  AOI211_X1 U69 ( .C1(n80), .C2(n81), .A(state[4]), .B(n34), .ZN(n216) );
  NOR3_X1 U70 ( .A1(state[0]), .A2(state[4]), .A3(n80), .ZN(n251) );
  NOR2_X1 U71 ( .A1(state[3]), .A2(state[2]), .ZN(n254) );
  NOR3_X1 U72 ( .A1(n97), .A2(n98), .A3(n96), .ZN(n169) );
  NOR3_X1 U73 ( .A1(n112), .A2(n113), .A3(n111), .ZN(n190) );
  NOR3_X1 U74 ( .A1(n81), .A2(state[4]), .A3(n80), .ZN(n255) );
  AOI211_X1 U75 ( .C1(n205), .C2(n29), .A(n183), .B(n206), .ZN(n193) );
  OAI22_X1 U76 ( .A1(n39), .A2(n191), .B1(n167), .B2(n169), .ZN(n206) );
  INV_X1 U77 ( .A(start), .ZN(n39) );
  NOR2_X1 U78 ( .A1(n79), .A2(state[3]), .ZN(n222) );
  NOR2_X1 U79 ( .A1(n211), .A2(state[0]), .ZN(n221) );
  NOR2_X1 U80 ( .A1(n81), .A2(n211), .ZN(n252) );
  NOR3_X1 U81 ( .A1(n91), .A2(n92), .A3(n90), .ZN(n194) );
  OAI221_X1 U82 ( .B1(n191), .B2(n38), .C1(n194), .C2(n119), .A(n202), .ZN(
        n198) );
  INV_X1 U83 ( .A(loadMatrix), .ZN(n38) );
  NAND4_X1 U84 ( .A1(state[4]), .A2(n254), .A3(state[0]), .A4(n80), .ZN(n172)
         );
  AOI22_X1 U85 ( .A1(n113), .A2(n216), .B1(n30), .B2(n219), .ZN(n217) );
  AOI21_X1 U86 ( .B1(n101), .B2(n123), .A(n124), .ZN(n243) );
  AOI21_X1 U87 ( .B1(n92), .B2(n145), .A(n124), .ZN(n146) );
  AOI21_X1 U88 ( .B1(n88), .B2(n153), .A(n124), .ZN(n154) );
  AOI21_X1 U89 ( .B1(n95), .B2(n137), .A(n124), .ZN(n138) );
  AOI21_X1 U90 ( .B1(n98), .B2(n127), .A(n124), .ZN(n128) );
  AOI21_X1 U91 ( .B1(n85), .B2(n162), .A(n124), .ZN(n163) );
  AOI21_X1 U92 ( .B1(n107), .B2(n228), .A(n124), .ZN(n229) );
  AOI21_X1 U93 ( .B1(n104), .B2(n236), .A(n124), .ZN(n237) );
  NOR2_X1 U94 ( .A1(n173), .A2(reset), .ZN(wr_en_a8) );
  NOR2_X1 U95 ( .A1(n167), .A2(reset), .ZN(wr_en_a5) );
  NOR2_X1 U96 ( .A1(n172), .A2(reset), .ZN(wr_en_a7) );
  NAND2_X1 U97 ( .A1(n253), .A2(n80), .ZN(n159) );
  NOR2_X1 U98 ( .A1(n159), .A2(reset), .ZN(wr_en_a6) );
  INV_X1 U99 ( .A(n257), .ZN(n31) );
  OAI21_X1 U100 ( .B1(n254), .B2(n76), .A(n258), .ZN(n257) );
  OAI211_X1 U101 ( .C1(n33), .C2(state[4]), .A(state[0]), .B(state[1]), .ZN(
        n258) );
  NOR2_X1 U102 ( .A1(reset), .A2(n117), .ZN(wr_en_x) );
  NOR2_X1 U103 ( .A1(reset), .A2(n116), .ZN(wr_en_y) );
  NOR2_X1 U104 ( .A1(reset), .A2(n121), .ZN(wr_en_a1) );
  OAI211_X1 U105 ( .C1(loadVector), .C2(n180), .A(n24), .B(n193), .ZN(n203) );
  INV_X1 U106 ( .A(n176), .ZN(n24) );
  NOR2_X1 U107 ( .A1(reset), .A2(n118), .ZN(wr_en_a4) );
  NOR2_X1 U108 ( .A1(reset), .A2(n120), .ZN(wr_en_a2) );
  NOR2_X1 U109 ( .A1(reset), .A2(n119), .ZN(wr_en_a3) );
  AND2_X1 U110 ( .A1(state[3]), .A2(state[2]), .ZN(n250) );
  NAND2_X1 U111 ( .A1(n76), .A2(n80), .ZN(n211) );
  NAND2_X1 U112 ( .A1(n253), .A2(state[1]), .ZN(n173) );
  AOI21_X1 U113 ( .B1(n181), .B2(n182), .A(reset), .ZN(N34) );
  AOI21_X1 U114 ( .B1(n29), .B2(n37), .A(N148), .ZN(n182) );
  NOR2_X1 U115 ( .A1(n177), .A2(n183), .ZN(n181) );
  AOI21_X1 U116 ( .B1(n185), .B2(n186), .A(reset), .ZN(N33) );
  AOI221_X1 U117 ( .B1(n187), .B2(loadVector), .C1(n23), .C2(n170), .A(n188), 
        .ZN(n186) );
  NOR3_X1 U118 ( .A1(n192), .A2(n150), .A3(n3), .ZN(n185) );
  NOR2_X1 U119 ( .A1(loadMatrix), .A2(n191), .ZN(n187) );
  AOI21_X1 U120 ( .B1(n196), .B2(n197), .A(reset), .ZN(N32) );
  NOR4_X1 U121 ( .A1(n198), .A2(n199), .A3(n200), .A4(n201), .ZN(n197) );
  AOI211_X1 U122 ( .C1(n32), .C2(n195), .A(n203), .B(n204), .ZN(n196) );
  NOR4_X1 U123 ( .A1(n118), .A2(n95), .A3(n94), .A4(n93), .ZN(n201) );
  NAND2_X1 U124 ( .A1(n221), .A2(n79), .ZN(n219) );
  OAI21_X1 U125 ( .B1(n243), .B2(n100), .A(n244), .ZN(N100) );
  OAI21_X1 U126 ( .B1(n237), .B2(n103), .A(n238), .ZN(N111) );
  OAI21_X1 U127 ( .B1(n229), .B2(n106), .A(n230), .ZN(N122) );
  OAI21_X1 U128 ( .B1(n146), .B2(n91), .A(n147), .ZN(N67) );
  OAI21_X1 U129 ( .B1(n154), .B2(n87), .A(n155), .ZN(N56) );
  OAI21_X1 U130 ( .B1(n138), .B2(n94), .A(n139), .ZN(N78) );
  OAI21_X1 U131 ( .B1(n163), .B2(n84), .A(n164), .ZN(N45) );
  OAI21_X1 U132 ( .B1(n128), .B2(n97), .A(n129), .ZN(N89) );
  OAI21_X1 U133 ( .B1(n217), .B2(n112), .A(n218), .ZN(N142) );
  OAI21_X1 U134 ( .B1(n214), .B2(n111), .A(n215), .ZN(N143) );
  NAND4_X1 U135 ( .A1(n216), .A2(addr_y[1]), .A3(addr_y[0]), .A4(n111), .ZN(
        n215) );
  AOI21_X1 U136 ( .B1(n216), .B2(n112), .A(n1), .ZN(n214) );
  INV_X1 U137 ( .A(n217), .ZN(n1) );
  AND3_X1 U138 ( .A1(n254), .A2(n81), .A3(state[4]), .ZN(n253) );
  NAND2_X1 U139 ( .A1(state[3]), .A2(n79), .ZN(n212) );
  OAI21_X1 U140 ( .B1(n241), .B2(n99), .A(n242), .ZN(N101) );
  NAND4_X1 U141 ( .A1(addr_a6[1]), .A2(addr_a6[0]), .A3(n123), .A4(n99), .ZN(
        n242) );
  AOI21_X1 U142 ( .B1(n123), .B2(n100), .A(n4), .ZN(n241) );
  INV_X1 U143 ( .A(n243), .ZN(n4) );
  OAI21_X1 U144 ( .B1(n151), .B2(n86), .A(n152), .ZN(N57) );
  NAND4_X1 U145 ( .A1(addr_a2[1]), .A2(addr_a2[0]), .A3(n153), .A4(n86), .ZN(
        n152) );
  AOI21_X1 U146 ( .B1(n153), .B2(n87), .A(n14), .ZN(n151) );
  INV_X1 U147 ( .A(n154), .ZN(n14) );
  OAI21_X1 U148 ( .B1(n135), .B2(n93), .A(n136), .ZN(N79) );
  NAND4_X1 U149 ( .A1(addr_a4[1]), .A2(addr_a4[0]), .A3(n137), .A4(n93), .ZN(
        n136) );
  AOI21_X1 U150 ( .B1(n137), .B2(n94), .A(n18), .ZN(n135) );
  INV_X1 U151 ( .A(n138), .ZN(n18) );
  OAI21_X1 U152 ( .B1(n143), .B2(n90), .A(n144), .ZN(N68) );
  NAND4_X1 U153 ( .A1(addr_a3[1]), .A2(addr_a3[0]), .A3(n145), .A4(n90), .ZN(
        n144) );
  AOI21_X1 U154 ( .B1(n145), .B2(n91), .A(n16), .ZN(n143) );
  INV_X1 U155 ( .A(n146), .ZN(n16) );
  OAI21_X1 U156 ( .B1(n125), .B2(n96), .A(n126), .ZN(N90) );
  NAND4_X1 U157 ( .A1(addr_a5[1]), .A2(addr_a5[0]), .A3(n127), .A4(n96), .ZN(
        n126) );
  AOI21_X1 U158 ( .B1(n127), .B2(n97), .A(n20), .ZN(n125) );
  INV_X1 U159 ( .A(n128), .ZN(n20) );
  OAI21_X1 U160 ( .B1(n160), .B2(n83), .A(n161), .ZN(N46) );
  NAND4_X1 U161 ( .A1(addr_a1[1]), .A2(addr_a1[0]), .A3(n162), .A4(n83), .ZN(
        n161) );
  AOI21_X1 U162 ( .B1(n162), .B2(n84), .A(n12), .ZN(n160) );
  INV_X1 U163 ( .A(n163), .ZN(n12) );
  OAI21_X1 U164 ( .B1(addr_y[0]), .B2(n30), .A(n220), .ZN(N141) );
  OAI21_X1 U165 ( .B1(n226), .B2(n105), .A(n227), .ZN(N123) );
  NAND4_X1 U166 ( .A1(addr_a8[1]), .A2(addr_a8[0]), .A3(n228), .A4(n105), .ZN(
        n227) );
  AOI21_X1 U167 ( .B1(n228), .B2(n106), .A(n9), .ZN(n226) );
  INV_X1 U168 ( .A(n229), .ZN(n9) );
  OAI21_X1 U169 ( .B1(n234), .B2(n102), .A(n235), .ZN(N112) );
  NAND4_X1 U170 ( .A1(addr_a7[1]), .A2(addr_a7[0]), .A3(n236), .A4(n102), .ZN(
        n235) );
  AOI21_X1 U171 ( .B1(n236), .B2(n103), .A(n7), .ZN(n234) );
  INV_X1 U172 ( .A(n237), .ZN(n7) );
  OAI21_X1 U173 ( .B1(n10), .B2(n108), .A(n223), .ZN(N133) );
  NOR2_X1 U174 ( .A1(addr_x[0]), .A2(n10), .ZN(N131) );
  NOR2_X1 U175 ( .A1(n10), .A2(n225), .ZN(N132) );
  XNOR2_X1 U176 ( .A(addr_x[1]), .B(addr_x[0]), .ZN(n225) );
  NOR2_X1 U177 ( .A1(reset), .A2(n174), .ZN(N35) );
  NOR3_X1 U178 ( .A1(n175), .A2(n176), .A3(n177), .ZN(n174) );
  OR4_X1 U179 ( .A1(n180), .A2(loadMatrix), .A3(loadVector), .A4(start), .ZN(
        n179) );
  INV_X1 U180 ( .A(n122), .ZN(n5) );
  AOI22_X1 U181 ( .A1(n101), .A2(n123), .B1(n124), .B2(addr_a6[0]), .ZN(n122)
         );
  INV_X1 U182 ( .A(n148), .ZN(n15) );
  AOI22_X1 U183 ( .A1(n92), .A2(n145), .B1(n124), .B2(addr_a3[0]), .ZN(n148)
         );
  INV_X1 U184 ( .A(n156), .ZN(n13) );
  AOI22_X1 U185 ( .A1(n88), .A2(n153), .B1(n124), .B2(addr_a2[0]), .ZN(n156)
         );
  INV_X1 U186 ( .A(n140), .ZN(n17) );
  AOI22_X1 U187 ( .A1(n95), .A2(n137), .B1(n124), .B2(addr_a4[0]), .ZN(n140)
         );
  INV_X1 U188 ( .A(n130), .ZN(n19) );
  AOI22_X1 U189 ( .A1(n98), .A2(n127), .B1(n124), .B2(addr_a5[0]), .ZN(n130)
         );
  INV_X1 U190 ( .A(n165), .ZN(n11) );
  AOI22_X1 U191 ( .A1(n85), .A2(n162), .B1(n124), .B2(addr_a1[0]), .ZN(n165)
         );
  INV_X1 U192 ( .A(n231), .ZN(n8) );
  AOI22_X1 U193 ( .A1(n107), .A2(n228), .B1(n124), .B2(addr_a8[0]), .ZN(n231)
         );
  INV_X1 U194 ( .A(n239), .ZN(n6) );
  AOI22_X1 U195 ( .A1(n104), .A2(n236), .B1(n124), .B2(addr_a7[0]), .ZN(n239)
         );
  NOR4_X1 U196 ( .A1(n159), .A2(n101), .A3(n100), .A4(n99), .ZN(n200) );
  NOR4_X1 U197 ( .A1(n120), .A2(n88), .A3(n87), .A4(n86), .ZN(n199) );
  NOR3_X1 U198 ( .A1(n84), .A2(n85), .A3(n83), .ZN(n184) );
  OAI22_X1 U199 ( .A1(n211), .A2(n34), .B1(n212), .B2(n213), .ZN(N147) );
  NAND2_X1 U200 ( .A1(n81), .A2(n76), .ZN(n213) );
endmodule


module mvm_8_8_16_1 ( clk, reset, loadMatrix, loadVector, start, done, data_in, 
        data_out );
  input [15:0] data_in;
  output [31:0] data_out;
  input clk, reset, loadMatrix, loadVector, start;
  output done;
  wire   wr_en_x, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6,
         wr_en_a7, wr_en_a8, wr_en_y, clear_acc, clc, clc1;
  wire   [2:0] addr_x;
  wire   [2:0] addr_a1;
  wire   [2:0] addr_a2;
  wire   [2:0] addr_a3;
  wire   [2:0] addr_a4;
  wire   [2:0] addr_a5;
  wire   [2:0] addr_a6;
  wire   [2:0] addr_a7;
  wire   [2:0] addr_a8;
  wire   [2:0] addr_y;

  datapath d ( .clk(clk), .data_in(data_in), .addr_x(addr_x), .wr_en_x(wr_en_x), .addr_a1(addr_a1), .addr_a2(addr_a2), .addr_a3(addr_a3), .addr_a4(addr_a4), 
        .addr_a5(addr_a5), .addr_a6(addr_a6), .addr_a7(addr_a7), .addr_a8(
        addr_a8), .wr_en_a1(wr_en_a1), .wr_en_a2(wr_en_a2), .wr_en_a3(wr_en_a3), .wr_en_a4(wr_en_a4), .wr_en_a5(wr_en_a5), .wr_en_a6(wr_en_a6), .wr_en_a7(
        wr_en_a7), .wr_en_a8(wr_en_a8), .addr_y(addr_y), .wr_en_y(wr_en_y), 
        .clear_acc(clear_acc), .clc(clc), .clc1(clc1), .data_out(data_out) );
  ctrlpath c ( .clk(clk), .reset(reset), .start(start), .addr_x(addr_x), 
        .wr_en_x(wr_en_x), .addr_a1(addr_a1), .addr_a2(addr_a2), .addr_a3(
        addr_a3), .addr_a4(addr_a4), .addr_a5(addr_a5), .addr_a6(addr_a6), 
        .addr_a7(addr_a7), .addr_a8(addr_a8), .wr_en_a1(wr_en_a1), .wr_en_a2(
        wr_en_a2), .wr_en_a3(wr_en_a3), .wr_en_a4(wr_en_a4), .wr_en_a5(
        wr_en_a5), .wr_en_a6(wr_en_a6), .wr_en_a7(wr_en_a7), .wr_en_a8(
        wr_en_a8), .clear_acc(clear_acc), .clc(clc), .clc1(clc1), .addr_y(
        addr_y), .wr_en_y(wr_en_y), .done(done), .loadMatrix(loadMatrix), 
        .loadVector(loadVector) );
endmodule

