include "s_thakkar_mvm_8_8_8_1.sv";
// Testbench, with parameters k=8, p=8, b=8, g=1

//This Test bench shows values on normal computation and in the next cycle only the vector is updated keeping the matrix same
 module tb1();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_8_8_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

// Set input values.
initial begin  
start=0; reset=1; data_in=8'bx;
@(posedge clk);
#1; reset=0; loadMatrix=1;
@(posedge clk);
#1; loadMatrix=0; data_in = 1;
@(posedge clk);
#1;data_in = 2;
@(posedge clk);
#1;data_in = 3;
@(posedge clk);
#1;data_in = 4;
@(posedge clk);
#1;data_in = 5;
@(posedge clk);
#1;data_in = 6;
@(posedge clk);
#1;data_in = 7;
@(posedge clk);
#1;data_in = 8;
@(posedge clk);
#1;data_in = 9;
@(posedge clk);
#1;data_in = 10;
@(posedge clk);
#1;data_in = 11;
@(posedge clk);
#1;data_in = 12;
@(posedge clk);
#1;data_in = 13;
@(posedge clk);
#1;data_in = 14;
@(posedge clk);
#1;data_in = 15;
@(posedge clk);
#1;data_in = 16;
@(posedge clk);
#1;data_in = 17;
@(posedge clk);
#1;data_in = 18;
@(posedge clk);
#1;data_in = 19;
@(posedge clk);
#1;data_in = 20;
@(posedge clk);
#1;data_in = 21;
@(posedge clk);
#1;data_in = 22;
@(posedge clk);
#1;data_in = 23;
@(posedge clk);
#1;data_in = 24;
@(posedge clk);
#1;data_in = 25;
@(posedge clk);
#1;data_in = 26;
@(posedge clk);
#1;data_in = 27;
@(posedge clk);
#1;data_in = 28;
@(posedge clk);
#1;data_in = 29;
@(posedge clk);
#1;data_in = 30;
@(posedge clk);
#1;data_in = 31;
@(posedge clk);
#1;data_in = 32;
@(posedge clk);
#1;data_in = 33;
@(posedge clk);
#1;data_in = 34;
@(posedge clk);
#1;data_in = 35;
@(posedge clk);
#1;data_in = 36;
@(posedge clk);
#1;data_in = 37;
@(posedge clk);
#1;data_in = 38;
@(posedge clk);
#1;data_in = 39;
@(posedge clk);
#1;data_in = 40;
@(posedge clk);
#1;data_in = 41;
@(posedge clk);
#1;data_in = 42;
@(posedge clk);
#1;data_in = 43;
@(posedge clk);
#1;data_in = 44;
@(posedge clk);
#1;data_in = 45;
@(posedge clk);
#1;data_in = 46;
@(posedge clk);
#1;data_in = 47;
@(posedge clk);
#1;data_in = 48;
@(posedge clk);
#1;data_in = 49;
@(posedge clk);
#1;data_in = 50;
@(posedge clk);
#1;data_in = 51;
@(posedge clk);
#1;data_in = 52;
@(posedge clk);
#1;data_in = 53;
@(posedge clk);
#1;data_in = 54;
@(posedge clk);
#1;data_in = 55;
@(posedge clk);
#1;data_in = 56;
@(posedge clk);
#1;data_in = 57;
@(posedge clk);
#1;data_in = 58;
@(posedge clk);
#1;data_in = 59;
@(posedge clk);
#1;data_in = 60;
@(posedge clk);
#1;data_in = 61;
@(posedge clk);
#1;data_in = 62;
@(posedge clk);
#1;data_in = 63;
@(posedge clk);
#1;data_in = 64;
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=1; 
@(posedge clk);
#1;data_in = 2;
@(posedge clk);
#1;data_in = 3;
@(posedge clk);
#1;data_in = 4;
@(posedge clk);
#1;data_in = 5;
@(posedge clk);
#1;data_in = 6;
@(posedge clk);
#1;data_in = 7;
@(posedge clk);
#1;data_in = 8;
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 end

integer filehandle=$fopen("proj3_outValuestb1");
// wait for done signal and output  
initial begin
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; loadVector=1;
@(posedge clk);
#1; loadVector=0;
data_in = 1;
@(posedge clk);
#1;data_in = -3;
@(posedge clk);
#1;data_in = -4;
@(posedge clk);
#1;data_in = -5;
@(posedge clk);
#1;data_in = -6;
@(posedge clk);
#1;data_in = -7;
@(posedge clk);
#1;data_in = -8;
@(posedge clk);
#1;data_in = -9;
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
//This testbench incorporates two iterations in the first iteration the values are computed according to the values and in the next iteration only the Matrix is updated keeping vector
module tb2();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_8_8_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

// Set input values.
initial begin  
start = 0; reset = 1;data_in=8'bx;
@(posedge clk);
#1; reset=0;
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
@(posedge clk);
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
start=0; reset=1; data_in=8'bx;
@(posedge clk);
#1; reset=0; loadMatrix=1;
@(posedge clk);
#1; loadMatrix=0; data_in = 1;
@(posedge clk);
#1;data_in = 2;
@(posedge clk);
#1;data_in = 3;
@(posedge clk);
#1;data_in = 4;
@(posedge clk);
#1;data_in = 5;
@(posedge clk);
#1;data_in = 6;
@(posedge clk);
#1;data_in = 7;
@(posedge clk);
#1;data_in = 8;
@(posedge clk);
#1;data_in = 9;
@(posedge clk);
#1;data_in = 10;
@(posedge clk);
#1;data_in = 11;
@(posedge clk);
#1;data_in = 12;
@(posedge clk);
#1;data_in = 13;
@(posedge clk);
#1;data_in = 14;
@(posedge clk);
#1;data_in = 15;
@(posedge clk);
#1;data_in = 16;
@(posedge clk);
#1;data_in = 17;
@(posedge clk);
#1;data_in = 18;
@(posedge clk);
#1;data_in = 19;
@(posedge clk);
#1;data_in = 20;
@(posedge clk);
#1;data_in = 21;
@(posedge clk);
#1;data_in = 22;
@(posedge clk);
#1;data_in = 23;
@(posedge clk);
#1;data_in = 24;
@(posedge clk);
#1;data_in = 25;
@(posedge clk);
#1;data_in = 26;
@(posedge clk);
#1;data_in = 27;
@(posedge clk);
#1;data_in = 28;
@(posedge clk);
#1;data_in = 29;
@(posedge clk);
#1;data_in = 30;
@(posedge clk);
#1;data_in = 31;
@(posedge clk);
#1;data_in = 32;
@(posedge clk);
#1;data_in = 33;
@(posedge clk);
#1;data_in = 34;
@(posedge clk);
#1;data_in = 35;
@(posedge clk);
#1;data_in = 36;
@(posedge clk);
#1;data_in = 37;
@(posedge clk);
#1;data_in = 38;
@(posedge clk);
#1;data_in = 39;
@(posedge clk);
#1;data_in = 40;
@(posedge clk);
#1;data_in = 41;
@(posedge clk);
#1;data_in = 42;
@(posedge clk);
#1;data_in = 43;
@(posedge clk);
#1;data_in = 44;
@(posedge clk);
#1;data_in = 45;
@(posedge clk);
#1;data_in = 46;
@(posedge clk);
#1;data_in = 47;
@(posedge clk);
#1;data_in = 48;
@(posedge clk);
#1;data_in = 49;
@(posedge clk);
#1;data_in = 50;
@(posedge clk);
#1;data_in = 51;
@(posedge clk);
#1;data_in = 52;
@(posedge clk);
#1;data_in = 53;
@(posedge clk);
#1;data_in = 54;
@(posedge clk);
#1;data_in = 55;
@(posedge clk);
#1;data_in = 56;
@(posedge clk);
#1;data_in = 57;
@(posedge clk);
#1;data_in = 58;
@(posedge clk);
#1;data_in = 59;
@(posedge clk);
#1;data_in = 60;
@(posedge clk);
#1;data_in = 61;
@(posedge clk);
#1;data_in = 62;
@(posedge clk);
#1;data_in = 63;
@(posedge clk);
#1;data_in = 64;
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=1; 
@(posedge clk);
#1;data_in = 2;
@(posedge clk);
#1;data_in = 3;
@(posedge clk);
#1;data_in = 4;
@(posedge clk);
#1;data_in = 5;
@(posedge clk);
#1;data_in = 6;
@(posedge clk);
#1;data_in = 7;
@(posedge clk);
#1;data_in = 8;
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 end

integer filehandle=$fopen("proj3_outValuestb2");
// wait for done signal and output  
initial begin
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; loadMatrix=1;
@(posedge clk);
#1; loadMatrix=0;
data_in = 1;
@(posedge clk);
#1;data_in = -5;
@(posedge clk);
#1;data_in = -6;
@(posedge clk);
#1;data_in = -7;
@(posedge clk);
#1;data_in = -8;
@(posedge clk);
#1;data_in = -9;
@(posedge clk);
#1;data_in = -10;
@(posedge clk);
#1;data_in = -11;
@(posedge clk);
#1;data_in = -12;
@(posedge clk);
#1;data_in = -13;
@(posedge clk);
#1;data_in = -14;
@(posedge clk);
#1;data_in = -15;
@(posedge clk);
#1;data_in = -16;
@(posedge clk);
#1;data_in = -17;
@(posedge clk);
#1;data_in = -18;
@(posedge clk);
#1;data_in = -19;
@(posedge clk);
#1;data_in = -20;
@(posedge clk);
#1;data_in = -21;
@(posedge clk);
#1;data_in = -22;
@(posedge clk);
#1;data_in = -23;
@(posedge clk);
#1;data_in = -24;
@(posedge clk);
#1;data_in = -25;
@(posedge clk);
#1;data_in = -26;
@(posedge clk);
#1;data_in = -27;
@(posedge clk);
#1;data_in = -28;
@(posedge clk);
#1;data_in = -29;
@(posedge clk);
#1;data_in = -30;
@(posedge clk);
#1;data_in = -31;
@(posedge clk);
#1;data_in = -32;
@(posedge clk);
#1;data_in = -33;
@(posedge clk);
#1;data_in = -34;
@(posedge clk);
#1;data_in = -35;
@(posedge clk);
#1;data_in = -36;
@(posedge clk);
#1;data_in = -37;
@(posedge clk);
#1;data_in = -38;
@(posedge clk);
#1;data_in = -39;
@(posedge clk);
#1;data_in = -40;
@(posedge clk);
#1;data_in = -41;
@(posedge clk);
#1;data_in = -42;
@(posedge clk);
#1;data_in = -43;
@(posedge clk);
#1;data_in = -44;
@(posedge clk);
#1;data_in = -45;
@(posedge clk);
#1;data_in = -46;
@(posedge clk);
#1;data_in = -47;
@(posedge clk);
#1;data_in = -48;
@(posedge clk);
#1;data_in = -49;
@(posedge clk);
#1;data_in = -50;
@(posedge clk);
#1;data_in = -51;
@(posedge clk);
#1;data_in = -52;
@(posedge clk);
#1;data_in = -53;
@(posedge clk);
#1;data_in = -54;
@(posedge clk);
#1;data_in = -55;
@(posedge clk);
#1;data_in = -56;
@(posedge clk);
#1;data_in = -57;
@(posedge clk);
#1;data_in = -58;
@(posedge clk);
#1;data_in = -59;
@(posedge clk);
#1;data_in = -60;
@(posedge clk);
#1;data_in = -61;
@(posedge clk);
#1;data_in = -62;
@(posedge clk);
#1;data_in = -63;
@(posedge clk);
#1;data_in = -64;
@(posedge clk);
#1;data_in = -65;
@(posedge clk);
#1;data_in = -66;
@(posedge clk);
#1;data_in = -67;
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
// Testbench, with parameters k=8, p=8, b=8, g=1

module tb3();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_8_8_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

logic [7:0] testData3[71:0];
   //read input from C file inputDatapart2     
 initial $readmemh("proj3_inputDatatb3", testData3);
 integer i;
 integer filehandle=$fopen("proj3_outValuestb3");
  initial begin 
  $monitor("Data in : %x",data_in);       
start  = 0; reset  = 1; data_in = 8'bx;
 @(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData3[0];
@(posedge clk);
#1;data_in = testData3[1];
@(posedge clk);
#1;data_in = testData3[2];
@(posedge clk);
#1;data_in = testData3[3];
@(posedge clk);
#1;data_in = testData3[4];
@(posedge clk);
#1;data_in = testData3[5];
@(posedge clk);
#1;data_in = testData3[6];
@(posedge clk);
#1;data_in = testData3[7];
@(posedge clk);
#1;data_in = testData3[8];
@(posedge clk);
#1;data_in = testData3[9];
@(posedge clk);
#1;data_in = testData3[10];
@(posedge clk);
#1;data_in = testData3[11];
@(posedge clk);
#1;data_in = testData3[12];
@(posedge clk);
#1;data_in = testData3[13];
@(posedge clk);
#1;data_in = testData3[14];
@(posedge clk);
#1;data_in = testData3[15];
@(posedge clk);
#1;data_in = testData3[16];
@(posedge clk);
#1;data_in = testData3[17];
@(posedge clk);
#1;data_in = testData3[18];
@(posedge clk);
#1;data_in = testData3[19];
@(posedge clk);
#1;data_in = testData3[20];
@(posedge clk);
#1;data_in = testData3[21];
@(posedge clk);
#1;data_in = testData3[22];
@(posedge clk);
#1;data_in = testData3[23];
@(posedge clk);
#1;data_in = testData3[24];
@(posedge clk);
#1;data_in = testData3[25];
@(posedge clk);
#1;data_in = testData3[26];
@(posedge clk);
#1;data_in = testData3[27];
@(posedge clk);
#1;data_in = testData3[28];
@(posedge clk);
#1;data_in = testData3[29];
@(posedge clk);
#1;data_in = testData3[30];
@(posedge clk);
#1;data_in = testData3[31];
@(posedge clk);
#1;data_in = testData3[32];
@(posedge clk);
#1;data_in = testData3[33];
@(posedge clk);
#1;data_in = testData3[34];
@(posedge clk);
#1;data_in = testData3[35];
@(posedge clk);
#1;data_in = testData3[36];
@(posedge clk);
#1;data_in = testData3[37];
@(posedge clk);
#1;data_in = testData3[38];
@(posedge clk);
#1;data_in = testData3[39];
@(posedge clk);
#1;data_in = testData3[40];
@(posedge clk);
#1;data_in = testData3[41];
@(posedge clk);
#1;data_in = testData3[42];
@(posedge clk);
#1;data_in = testData3[43];
@(posedge clk);
#1;data_in = testData3[44];
@(posedge clk);
#1;data_in = testData3[45];
@(posedge clk);
#1;data_in = testData3[46];
@(posedge clk);
#1;data_in = testData3[47];
@(posedge clk);
#1;data_in = testData3[48];
@(posedge clk);
#1;data_in = testData3[49];
@(posedge clk);
#1;data_in = testData3[50];
@(posedge clk);
#1;data_in = testData3[51];
@(posedge clk);
#1;data_in = testData3[52];
@(posedge clk);
#1;data_in = testData3[53];
@(posedge clk);
#1;data_in = testData3[54];
@(posedge clk);
#1;data_in = testData3[55];
@(posedge clk);
#1;data_in = testData3[56];
@(posedge clk);
#1;data_in = testData3[57];
@(posedge clk);
#1;data_in = testData3[58];
@(posedge clk);
#1;data_in = testData3[59];
@(posedge clk);
#1;data_in = testData3[60];
@(posedge clk);
#1;data_in = testData3[61];
@(posedge clk);
#1;data_in = testData3[62];
@(posedge clk);
#1;data_in = testData3[63];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData3[64]; 
@(posedge clk);
#1;data_in = testData3[65];
@(posedge clk);
#1;data_in = testData3[66];
@(posedge clk);
#1;data_in = testData3[67];
@(posedge clk);
#1;data_in = testData3[68];
@(posedge clk);
#1;data_in = testData3[69];
@(posedge clk);
#1;data_in = testData3[70];
@(posedge clk);
#1;data_in = testData3[71];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 end

// wait for done signal and output  
initial begin
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
// Testbench, with parameters k=8, p=8, b=8, g=1

module tb4();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_8_8_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

logic [7:0] testData4[471:0];
   //read input from C file inputDatapart1     
 initial $readmemh("proj3_inputDatatb4", testData4);
 integer i;
 integer filehandle=$fopen("proj3_outValuestb4");
  initial begin 
start  = 0; reset  = 1; data_in = 8'bx;
 @(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData4[0];
@(posedge clk);
#1;data_in = testData4[1];
@(posedge clk);
#1;data_in = testData4[2];
@(posedge clk);
#1;data_in = testData4[3];
@(posedge clk);
#1;data_in = testData4[4];
@(posedge clk);
#1;data_in = testData4[5];
@(posedge clk);
#1;data_in = testData4[6];
@(posedge clk);
#1;data_in = testData4[7];
@(posedge clk);
#1;data_in = testData4[8];
@(posedge clk);
#1;data_in = testData4[9];
@(posedge clk);
#1;data_in = testData4[10];
@(posedge clk);
#1;data_in = testData4[11];
@(posedge clk);
#1;data_in = testData4[12];
@(posedge clk);
#1;data_in = testData4[13];
@(posedge clk);
#1;data_in = testData4[14];
@(posedge clk);
#1;data_in = testData4[15];
@(posedge clk);
#1;data_in = testData4[16];
@(posedge clk);
#1;data_in = testData4[17];
@(posedge clk);
#1;data_in = testData4[18];
@(posedge clk);
#1;data_in = testData4[19];
@(posedge clk);
#1;data_in = testData4[20];
@(posedge clk);
#1;data_in = testData4[21];
@(posedge clk);
#1;data_in = testData4[22];
@(posedge clk);
#1;data_in = testData4[23];
@(posedge clk);
#1;data_in = testData4[24];
@(posedge clk);
#1;data_in = testData4[25];
@(posedge clk);
#1;data_in = testData4[26];
@(posedge clk);
#1;data_in = testData4[27];
@(posedge clk);
#1;data_in = testData4[28];
@(posedge clk);
#1;data_in = testData4[29];
@(posedge clk);
#1;data_in = testData4[30];
@(posedge clk);
#1;data_in = testData4[31];
@(posedge clk);
#1;data_in = testData4[32];
@(posedge clk);
#1;data_in = testData4[33];
@(posedge clk);
#1;data_in = testData4[34];
@(posedge clk);
#1;data_in = testData4[35];
@(posedge clk);
#1;data_in = testData4[36];
@(posedge clk);
#1;data_in = testData4[37];
@(posedge clk);
#1;data_in = testData4[38];
@(posedge clk);
#1;data_in = testData4[39];
@(posedge clk);
#1;data_in = testData4[40];
@(posedge clk);
#1;data_in = testData4[41];
@(posedge clk);
#1;data_in = testData4[42];
@(posedge clk);
#1;data_in = testData4[43];
@(posedge clk);
#1;data_in = testData4[44];
@(posedge clk);
#1;data_in = testData4[45];
@(posedge clk);
#1;data_in = testData4[46];
@(posedge clk);
#1;data_in = testData4[47];
@(posedge clk);
#1;data_in = testData4[48];
@(posedge clk);
#1;data_in = testData4[49];
@(posedge clk);
#1;data_in = testData4[50];
@(posedge clk);
#1;data_in = testData4[51];
@(posedge clk);
#1;data_in = testData4[52];
@(posedge clk);
#1;data_in = testData4[53];
@(posedge clk);
#1;data_in = testData4[54];
@(posedge clk);
#1;data_in = testData4[55];
@(posedge clk);
#1;data_in = testData4[56];
@(posedge clk);
#1;data_in = testData4[57];
@(posedge clk);
#1;data_in = testData4[58];
@(posedge clk);
#1;data_in = testData4[59];
@(posedge clk);
#1;data_in = testData4[60];
@(posedge clk);
#1;data_in = testData4[61];
@(posedge clk);
#1;data_in = testData4[62];
@(posedge clk);
#1;data_in = testData4[63];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData4[64]; 
@(posedge clk);
#1;data_in = testData4[65];
@(posedge clk);
#1;data_in = testData4[66];
@(posedge clk);
#1;data_in = testData4[67];
@(posedge clk);
#1;data_in = testData4[68];
@(posedge clk);
#1;data_in = testData4[69];
@(posedge clk);
#1;data_in = testData4[70];
@(posedge clk);
#1;data_in = testData4[71];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 end

// wait for done signal and output  
initial begin
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[72]; 
@(posedge clk);
#1;data_in = testData4[73];
@(posedge clk);
#1;data_in = testData4[74];
@(posedge clk);
#1;data_in = testData4[75];
@(posedge clk);
#1;data_in = testData4[76];
@(posedge clk);
#1;data_in = testData4[77];
@(posedge clk);
#1;data_in = testData4[78];
@(posedge clk);
#1;data_in = testData4[79];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[80]; 
@(posedge clk);
#1;data_in = testData4[81];
@(posedge clk);
#1;data_in = testData4[82];
@(posedge clk);
#1;data_in = testData4[83];
@(posedge clk);
#1;data_in = testData4[84];
@(posedge clk);
#1;data_in = testData4[85];
@(posedge clk);
#1;data_in = testData4[86];
@(posedge clk);
#1;data_in = testData4[87];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[88]; 
@(posedge clk);
#1;data_in = testData4[89];
@(posedge clk);
#1;data_in = testData4[90];
@(posedge clk);
#1;data_in = testData4[91];
@(posedge clk);
#1;data_in = testData4[92];
@(posedge clk);
#1;data_in = testData4[93];
@(posedge clk);
#1;data_in = testData4[94];
@(posedge clk);
#1;data_in = testData4[95];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[96]; 
@(posedge clk);
#1;data_in = testData4[97];
@(posedge clk);
#1;data_in = testData4[98];
@(posedge clk);
#1;data_in = testData4[99];
@(posedge clk);
#1;data_in = testData4[100];
@(posedge clk);
#1;data_in = testData4[101];
@(posedge clk);
#1;data_in = testData4[102];
@(posedge clk);
#1;data_in = testData4[103];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[104]; 
@(posedge clk);
#1;data_in = testData4[105];
@(posedge clk);
#1;data_in = testData4[106];
@(posedge clk);
#1;data_in = testData4[107];
@(posedge clk);
#1;data_in = testData4[108];
@(posedge clk);
#1;data_in = testData4[109];
@(posedge clk);
#1;data_in = testData4[110];
@(posedge clk);
#1;data_in = testData4[111];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[112]; 
@(posedge clk);
#1;data_in = testData4[113];
@(posedge clk);
#1;data_in = testData4[114];
@(posedge clk);
#1;data_in = testData4[115];
@(posedge clk);
#1;data_in = testData4[116];
@(posedge clk);
#1;data_in = testData4[117];
@(posedge clk);
#1;data_in = testData4[118];
@(posedge clk);
#1;data_in = testData4[119];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[120]; 
@(posedge clk);
#1;data_in = testData4[121];
@(posedge clk);
#1;data_in = testData4[122];
@(posedge clk);
#1;data_in = testData4[123];
@(posedge clk);
#1;data_in = testData4[124];
@(posedge clk);
#1;data_in = testData4[125];
@(posedge clk);
#1;data_in = testData4[126];
@(posedge clk);
#1;data_in = testData4[127];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[128]; 
@(posedge clk);
#1;data_in = testData4[129];
@(posedge clk);
#1;data_in = testData4[130];
@(posedge clk);
#1;data_in = testData4[131];
@(posedge clk);
#1;data_in = testData4[132];
@(posedge clk);
#1;data_in = testData4[133];
@(posedge clk);
#1;data_in = testData4[134];
@(posedge clk);
#1;data_in = testData4[135];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[136]; 
@(posedge clk);
#1;data_in = testData4[137];
@(posedge clk);
#1;data_in = testData4[138];
@(posedge clk);
#1;data_in = testData4[139];
@(posedge clk);
#1;data_in = testData4[140];
@(posedge clk);
#1;data_in = testData4[141];
@(posedge clk);
#1;data_in = testData4[142];
@(posedge clk);
#1;data_in = testData4[143];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[144]; 
@(posedge clk);
#1;data_in = testData4[145];
@(posedge clk);
#1;data_in = testData4[146];
@(posedge clk);
#1;data_in = testData4[147];
@(posedge clk);
#1;data_in = testData4[148];
@(posedge clk);
#1;data_in = testData4[149];
@(posedge clk);
#1;data_in = testData4[150];
@(posedge clk);
#1;data_in = testData4[151];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[152]; 
@(posedge clk);
#1;data_in = testData4[153];
@(posedge clk);
#1;data_in = testData4[154];
@(posedge clk);
#1;data_in = testData4[155];
@(posedge clk);
#1;data_in = testData4[156];
@(posedge clk);
#1;data_in = testData4[157];
@(posedge clk);
#1;data_in = testData4[158];
@(posedge clk);
#1;data_in = testData4[159];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[160]; 
@(posedge clk);
#1;data_in = testData4[161];
@(posedge clk);
#1;data_in = testData4[162];
@(posedge clk);
#1;data_in = testData4[163];
@(posedge clk);
#1;data_in = testData4[164];
@(posedge clk);
#1;data_in = testData4[165];
@(posedge clk);
#1;data_in = testData4[166];
@(posedge clk);
#1;data_in = testData4[167];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[168]; 
@(posedge clk);
#1;data_in = testData4[169];
@(posedge clk);
#1;data_in = testData4[170];
@(posedge clk);
#1;data_in = testData4[171];
@(posedge clk);
#1;data_in = testData4[172];
@(posedge clk);
#1;data_in = testData4[173];
@(posedge clk);
#1;data_in = testData4[174];
@(posedge clk);
#1;data_in = testData4[175];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[176]; 
@(posedge clk);
#1;data_in = testData4[177];
@(posedge clk);
#1;data_in = testData4[178];
@(posedge clk);
#1;data_in = testData4[179];
@(posedge clk);
#1;data_in = testData4[180];
@(posedge clk);
#1;data_in = testData4[181];
@(posedge clk);
#1;data_in = testData4[182];
@(posedge clk);
#1;data_in = testData4[183];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[184]; 
@(posedge clk);
#1;data_in = testData4[185];
@(posedge clk);
#1;data_in = testData4[186];
@(posedge clk);
#1;data_in = testData4[187];
@(posedge clk);
#1;data_in = testData4[188];
@(posedge clk);
#1;data_in = testData4[189];
@(posedge clk);
#1;data_in = testData4[190];
@(posedge clk);
#1;data_in = testData4[191];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[192]; 
@(posedge clk);
#1;data_in = testData4[193];
@(posedge clk);
#1;data_in = testData4[194];
@(posedge clk);
#1;data_in = testData4[195];
@(posedge clk);
#1;data_in = testData4[196];
@(posedge clk);
#1;data_in = testData4[197];
@(posedge clk);
#1;data_in = testData4[198];
@(posedge clk);
#1;data_in = testData4[199];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[200]; 
@(posedge clk);
#1;data_in = testData4[201];
@(posedge clk);
#1;data_in = testData4[202];
@(posedge clk);
#1;data_in = testData4[203];
@(posedge clk);
#1;data_in = testData4[204];
@(posedge clk);
#1;data_in = testData4[205];
@(posedge clk);
#1;data_in = testData4[206];
@(posedge clk);
#1;data_in = testData4[207];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[208]; 
@(posedge clk);
#1;data_in = testData4[209];
@(posedge clk);
#1;data_in = testData4[210];
@(posedge clk);
#1;data_in = testData4[211];
@(posedge clk);
#1;data_in = testData4[212];
@(posedge clk);
#1;data_in = testData4[213];
@(posedge clk);
#1;data_in = testData4[214];
@(posedge clk);
#1;data_in = testData4[215];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[216]; 
@(posedge clk);
#1;data_in = testData4[217];
@(posedge clk);
#1;data_in = testData4[218];
@(posedge clk);
#1;data_in = testData4[219];
@(posedge clk);
#1;data_in = testData4[220];
@(posedge clk);
#1;data_in = testData4[221];
@(posedge clk);
#1;data_in = testData4[222];
@(posedge clk);
#1;data_in = testData4[223];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[224]; 
@(posedge clk);
#1;data_in = testData4[225];
@(posedge clk);
#1;data_in = testData4[226];
@(posedge clk);
#1;data_in = testData4[227];
@(posedge clk);
#1;data_in = testData4[228];
@(posedge clk);
#1;data_in = testData4[229];
@(posedge clk);
#1;data_in = testData4[230];
@(posedge clk);
#1;data_in = testData4[231];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[232]; 
@(posedge clk);
#1;data_in = testData4[233];
@(posedge clk);
#1;data_in = testData4[234];
@(posedge clk);
#1;data_in = testData4[235];
@(posedge clk);
#1;data_in = testData4[236];
@(posedge clk);
#1;data_in = testData4[237];
@(posedge clk);
#1;data_in = testData4[238];
@(posedge clk);
#1;data_in = testData4[239];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[240]; 
@(posedge clk);
#1;data_in = testData4[241];
@(posedge clk);
#1;data_in = testData4[242];
@(posedge clk);
#1;data_in = testData4[243];
@(posedge clk);
#1;data_in = testData4[244];
@(posedge clk);
#1;data_in = testData4[245];
@(posedge clk);
#1;data_in = testData4[246];
@(posedge clk);
#1;data_in = testData4[247];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[248]; 
@(posedge clk);
#1;data_in = testData4[249];
@(posedge clk);
#1;data_in = testData4[250];
@(posedge clk);
#1;data_in = testData4[251];
@(posedge clk);
#1;data_in = testData4[252];
@(posedge clk);
#1;data_in = testData4[253];
@(posedge clk);
#1;data_in = testData4[254];
@(posedge clk);
#1;data_in = testData4[255];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[256]; 
@(posedge clk);
#1;data_in = testData4[257];
@(posedge clk);
#1;data_in = testData4[258];
@(posedge clk);
#1;data_in = testData4[259];
@(posedge clk);
#1;data_in = testData4[260];
@(posedge clk);
#1;data_in = testData4[261];
@(posedge clk);
#1;data_in = testData4[262];
@(posedge clk);
#1;data_in = testData4[263];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[264]; 
@(posedge clk);
#1;data_in = testData4[265];
@(posedge clk);
#1;data_in = testData4[266];
@(posedge clk);
#1;data_in = testData4[267];
@(posedge clk);
#1;data_in = testData4[268];
@(posedge clk);
#1;data_in = testData4[269];
@(posedge clk);
#1;data_in = testData4[270];
@(posedge clk);
#1;data_in = testData4[271];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[272]; 
@(posedge clk);
#1;data_in = testData4[273];
@(posedge clk);
#1;data_in = testData4[274];
@(posedge clk);
#1;data_in = testData4[275];
@(posedge clk);
#1;data_in = testData4[276];
@(posedge clk);
#1;data_in = testData4[277];
@(posedge clk);
#1;data_in = testData4[278];
@(posedge clk);
#1;data_in = testData4[279];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[280]; 
@(posedge clk);
#1;data_in = testData4[281];
@(posedge clk);
#1;data_in = testData4[282];
@(posedge clk);
#1;data_in = testData4[283];
@(posedge clk);
#1;data_in = testData4[284];
@(posedge clk);
#1;data_in = testData4[285];
@(posedge clk);
#1;data_in = testData4[286];
@(posedge clk);
#1;data_in = testData4[287];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[288]; 
@(posedge clk);
#1;data_in = testData4[289];
@(posedge clk);
#1;data_in = testData4[290];
@(posedge clk);
#1;data_in = testData4[291];
@(posedge clk);
#1;data_in = testData4[292];
@(posedge clk);
#1;data_in = testData4[293];
@(posedge clk);
#1;data_in = testData4[294];
@(posedge clk);
#1;data_in = testData4[295];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[296]; 
@(posedge clk);
#1;data_in = testData4[297];
@(posedge clk);
#1;data_in = testData4[298];
@(posedge clk);
#1;data_in = testData4[299];
@(posedge clk);
#1;data_in = testData4[300];
@(posedge clk);
#1;data_in = testData4[301];
@(posedge clk);
#1;data_in = testData4[302];
@(posedge clk);
#1;data_in = testData4[303];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[304]; 
@(posedge clk);
#1;data_in = testData4[305];
@(posedge clk);
#1;data_in = testData4[306];
@(posedge clk);
#1;data_in = testData4[307];
@(posedge clk);
#1;data_in = testData4[308];
@(posedge clk);
#1;data_in = testData4[309];
@(posedge clk);
#1;data_in = testData4[310];
@(posedge clk);
#1;data_in = testData4[311];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[312]; 
@(posedge clk);
#1;data_in = testData4[313];
@(posedge clk);
#1;data_in = testData4[314];
@(posedge clk);
#1;data_in = testData4[315];
@(posedge clk);
#1;data_in = testData4[316];
@(posedge clk);
#1;data_in = testData4[317];
@(posedge clk);
#1;data_in = testData4[318];
@(posedge clk);
#1;data_in = testData4[319];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[320]; 
@(posedge clk);
#1;data_in = testData4[321];
@(posedge clk);
#1;data_in = testData4[322];
@(posedge clk);
#1;data_in = testData4[323];
@(posedge clk);
#1;data_in = testData4[324];
@(posedge clk);
#1;data_in = testData4[325];
@(posedge clk);
#1;data_in = testData4[326];
@(posedge clk);
#1;data_in = testData4[327];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[328]; 
@(posedge clk);
#1;data_in = testData4[329];
@(posedge clk);
#1;data_in = testData4[330];
@(posedge clk);
#1;data_in = testData4[331];
@(posedge clk);
#1;data_in = testData4[332];
@(posedge clk);
#1;data_in = testData4[333];
@(posedge clk);
#1;data_in = testData4[334];
@(posedge clk);
#1;data_in = testData4[335];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[336]; 
@(posedge clk);
#1;data_in = testData4[337];
@(posedge clk);
#1;data_in = testData4[338];
@(posedge clk);
#1;data_in = testData4[339];
@(posedge clk);
#1;data_in = testData4[340];
@(posedge clk);
#1;data_in = testData4[341];
@(posedge clk);
#1;data_in = testData4[342];
@(posedge clk);
#1;data_in = testData4[343];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[344]; 
@(posedge clk);
#1;data_in = testData4[345];
@(posedge clk);
#1;data_in = testData4[346];
@(posedge clk);
#1;data_in = testData4[347];
@(posedge clk);
#1;data_in = testData4[348];
@(posedge clk);
#1;data_in = testData4[349];
@(posedge clk);
#1;data_in = testData4[350];
@(posedge clk);
#1;data_in = testData4[351];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[352]; 
@(posedge clk);
#1;data_in = testData4[353];
@(posedge clk);
#1;data_in = testData4[354];
@(posedge clk);
#1;data_in = testData4[355];
@(posedge clk);
#1;data_in = testData4[356];
@(posedge clk);
#1;data_in = testData4[357];
@(posedge clk);
#1;data_in = testData4[358];
@(posedge clk);
#1;data_in = testData4[359];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[360]; 
@(posedge clk);
#1;data_in = testData4[361];
@(posedge clk);
#1;data_in = testData4[362];
@(posedge clk);
#1;data_in = testData4[363];
@(posedge clk);
#1;data_in = testData4[364];
@(posedge clk);
#1;data_in = testData4[365];
@(posedge clk);
#1;data_in = testData4[366];
@(posedge clk);
#1;data_in = testData4[367];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[368]; 
@(posedge clk);
#1;data_in = testData4[369];
@(posedge clk);
#1;data_in = testData4[370];
@(posedge clk);
#1;data_in = testData4[371];
@(posedge clk);
#1;data_in = testData4[372];
@(posedge clk);
#1;data_in = testData4[373];
@(posedge clk);
#1;data_in = testData4[374];
@(posedge clk);
#1;data_in = testData4[375];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[376]; 
@(posedge clk);
#1;data_in = testData4[377];
@(posedge clk);
#1;data_in = testData4[378];
@(posedge clk);
#1;data_in = testData4[379];
@(posedge clk);
#1;data_in = testData4[380];
@(posedge clk);
#1;data_in = testData4[381];
@(posedge clk);
#1;data_in = testData4[382];
@(posedge clk);
#1;data_in = testData4[383];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[384]; 
@(posedge clk);
#1;data_in = testData4[385];
@(posedge clk);
#1;data_in = testData4[386];
@(posedge clk);
#1;data_in = testData4[387];
@(posedge clk);
#1;data_in = testData4[388];
@(posedge clk);
#1;data_in = testData4[389];
@(posedge clk);
#1;data_in = testData4[390];
@(posedge clk);
#1;data_in = testData4[391];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[392]; 
@(posedge clk);
#1;data_in = testData4[393];
@(posedge clk);
#1;data_in = testData4[394];
@(posedge clk);
#1;data_in = testData4[395];
@(posedge clk);
#1;data_in = testData4[396];
@(posedge clk);
#1;data_in = testData4[397];
@(posedge clk);
#1;data_in = testData4[398];
@(posedge clk);
#1;data_in = testData4[399];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[400]; 
@(posedge clk);
#1;data_in = testData4[401];
@(posedge clk);
#1;data_in = testData4[402];
@(posedge clk);
#1;data_in = testData4[403];
@(posedge clk);
#1;data_in = testData4[404];
@(posedge clk);
#1;data_in = testData4[405];
@(posedge clk);
#1;data_in = testData4[406];
@(posedge clk);
#1;data_in = testData4[407];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[408]; 
@(posedge clk);
#1;data_in = testData4[409];
@(posedge clk);
#1;data_in = testData4[410];
@(posedge clk);
#1;data_in = testData4[411];
@(posedge clk);
#1;data_in = testData4[412];
@(posedge clk);
#1;data_in = testData4[413];
@(posedge clk);
#1;data_in = testData4[414];
@(posedge clk);
#1;data_in = testData4[415];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[416]; 
@(posedge clk);
#1;data_in = testData4[417];
@(posedge clk);
#1;data_in = testData4[418];
@(posedge clk);
#1;data_in = testData4[419];
@(posedge clk);
#1;data_in = testData4[420];
@(posedge clk);
#1;data_in = testData4[421];
@(posedge clk);
#1;data_in = testData4[422];
@(posedge clk);
#1;data_in = testData4[423];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[424]; 
@(posedge clk);
#1;data_in = testData4[425];
@(posedge clk);
#1;data_in = testData4[426];
@(posedge clk);
#1;data_in = testData4[427];
@(posedge clk);
#1;data_in = testData4[428];
@(posedge clk);
#1;data_in = testData4[429];
@(posedge clk);
#1;data_in = testData4[430];
@(posedge clk);
#1;data_in = testData4[431];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[432]; 
@(posedge clk);
#1;data_in = testData4[433];
@(posedge clk);
#1;data_in = testData4[434];
@(posedge clk);
#1;data_in = testData4[435];
@(posedge clk);
#1;data_in = testData4[436];
@(posedge clk);
#1;data_in = testData4[437];
@(posedge clk);
#1;data_in = testData4[438];
@(posedge clk);
#1;data_in = testData4[439];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[440]; 
@(posedge clk);
#1;data_in = testData4[441];
@(posedge clk);
#1;data_in = testData4[442];
@(posedge clk);
#1;data_in = testData4[443];
@(posedge clk);
#1;data_in = testData4[444];
@(posedge clk);
#1;data_in = testData4[445];
@(posedge clk);
#1;data_in = testData4[446];
@(posedge clk);
#1;data_in = testData4[447];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[448]; 
@(posedge clk);
#1;data_in = testData4[449];
@(posedge clk);
#1;data_in = testData4[450];
@(posedge clk);
#1;data_in = testData4[451];
@(posedge clk);
#1;data_in = testData4[452];
@(posedge clk);
#1;data_in = testData4[453];
@(posedge clk);
#1;data_in = testData4[454];
@(posedge clk);
#1;data_in = testData4[455];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[456]; 
@(posedge clk);
#1;data_in = testData4[457];
@(posedge clk);
#1;data_in = testData4[458];
@(posedge clk);
#1;data_in = testData4[459];
@(posedge clk);
#1;data_in = testData4[460];
@(posedge clk);
#1;data_in = testData4[461];
@(posedge clk);
#1;data_in = testData4[462];
@(posedge clk);
#1;data_in = testData4[463];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[464]; 
@(posedge clk);
#1;data_in = testData4[465];
@(posedge clk);
#1;data_in = testData4[466];
@(posedge clk);
#1;data_in = testData4[467];
@(posedge clk);
#1;data_in = testData4[468];
@(posedge clk);
#1;data_in = testData4[469];
@(posedge clk);
#1;data_in = testData4[470];
@(posedge clk);
#1;data_in = testData4[471];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
module tb6();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_8_8_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

logic [7:0] testData6[3671:0];
   //read input from C file inputDatapart2     
 initial $readmemh("proj3_inputDatatb6", testData6);
 integer i;
 integer filehandle=$fopen("proj3_outValuestb6");
  initial begin 
  $monitor("Data in : %x",data_in);       
start  = 0; reset  = 1; data_in = 8'bx;
 @(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[0];
@(posedge clk);
#1;data_in = testData6[1];
@(posedge clk);
#1;data_in = testData6[2];
@(posedge clk);
#1;data_in = testData6[3];
@(posedge clk);
#1;data_in = testData6[4];
@(posedge clk);
#1;data_in = testData6[5];
@(posedge clk);
#1;data_in = testData6[6];
@(posedge clk);
#1;data_in = testData6[7];
@(posedge clk);
#1;data_in = testData6[8];
@(posedge clk);
#1;data_in = testData6[9];
@(posedge clk);
#1;data_in = testData6[10];
@(posedge clk);
#1;data_in = testData6[11];
@(posedge clk);
#1;data_in = testData6[12];
@(posedge clk);
#1;data_in = testData6[13];
@(posedge clk);
#1;data_in = testData6[14];
@(posedge clk);
#1;data_in = testData6[15];
@(posedge clk);
#1;data_in = testData6[16];
@(posedge clk);
#1;data_in = testData6[17];
@(posedge clk);
#1;data_in = testData6[18];
@(posedge clk);
#1;data_in = testData6[19];
@(posedge clk);
#1;data_in = testData6[20];
@(posedge clk);
#1;data_in = testData6[21];
@(posedge clk);
#1;data_in = testData6[22];
@(posedge clk);
#1;data_in = testData6[23];
@(posedge clk);
#1;data_in = testData6[24];
@(posedge clk);
#1;data_in = testData6[25];
@(posedge clk);
#1;data_in = testData6[26];
@(posedge clk);
#1;data_in = testData6[27];
@(posedge clk);
#1;data_in = testData6[28];
@(posedge clk);
#1;data_in = testData6[29];
@(posedge clk);
#1;data_in = testData6[30];
@(posedge clk);
#1;data_in = testData6[31];
@(posedge clk);
#1;data_in = testData6[32];
@(posedge clk);
#1;data_in = testData6[33];
@(posedge clk);
#1;data_in = testData6[34];
@(posedge clk);
#1;data_in = testData6[35];
@(posedge clk);
#1;data_in = testData6[36];
@(posedge clk);
#1;data_in = testData6[37];
@(posedge clk);
#1;data_in = testData6[38];
@(posedge clk);
#1;data_in = testData6[39];
@(posedge clk);
#1;data_in = testData6[40];
@(posedge clk);
#1;data_in = testData6[41];
@(posedge clk);
#1;data_in = testData6[42];
@(posedge clk);
#1;data_in = testData6[43];
@(posedge clk);
#1;data_in = testData6[44];
@(posedge clk);
#1;data_in = testData6[45];
@(posedge clk);
#1;data_in = testData6[46];
@(posedge clk);
#1;data_in = testData6[47];
@(posedge clk);
#1;data_in = testData6[48];
@(posedge clk);
#1;data_in = testData6[49];
@(posedge clk);
#1;data_in = testData6[50];
@(posedge clk);
#1;data_in = testData6[51];
@(posedge clk);
#1;data_in = testData6[52];
@(posedge clk);
#1;data_in = testData6[53];
@(posedge clk);
#1;data_in = testData6[54];
@(posedge clk);
#1;data_in = testData6[55];
@(posedge clk);
#1;data_in = testData6[56];
@(posedge clk);
#1;data_in = testData6[57];
@(posedge clk);
#1;data_in = testData6[58];
@(posedge clk);
#1;data_in = testData6[59];
@(posedge clk);
#1;data_in = testData6[60];
@(posedge clk);
#1;data_in = testData6[61];
@(posedge clk);
#1;data_in = testData6[62];
@(posedge clk);
#1;data_in = testData6[63];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[64]; 
@(posedge clk);
#1;data_in = testData6[65];
@(posedge clk);
#1;data_in = testData6[66];
@(posedge clk);
#1;data_in = testData6[67];
@(posedge clk);
#1;data_in = testData6[68];
@(posedge clk);
#1;data_in = testData6[69];
@(posedge clk);
#1;data_in = testData6[70];
@(posedge clk);
#1;data_in = testData6[71];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[72];
@(posedge clk);
#1;data_in = testData6[73];
@(posedge clk);
#1;data_in = testData6[74];
@(posedge clk);
#1;data_in = testData6[75];
@(posedge clk);
#1;data_in = testData6[76];
@(posedge clk);
#1;data_in = testData6[77];
@(posedge clk);
#1;data_in = testData6[78];
@(posedge clk);
#1;data_in = testData6[79];
@(posedge clk);
#1;data_in = testData6[80];
@(posedge clk);
#1;data_in = testData6[81];
@(posedge clk);
#1;data_in = testData6[82];
@(posedge clk);
#1;data_in = testData6[83];
@(posedge clk);
#1;data_in = testData6[84];
@(posedge clk);
#1;data_in = testData6[85];
@(posedge clk);
#1;data_in = testData6[86];
@(posedge clk);
#1;data_in = testData6[87];
@(posedge clk);
#1;data_in = testData6[88];
@(posedge clk);
#1;data_in = testData6[89];
@(posedge clk);
#1;data_in = testData6[90];
@(posedge clk);
#1;data_in = testData6[91];
@(posedge clk);
#1;data_in = testData6[92];
@(posedge clk);
#1;data_in = testData6[93];
@(posedge clk);
#1;data_in = testData6[94];
@(posedge clk);
#1;data_in = testData6[95];
@(posedge clk);
#1;data_in = testData6[96];
@(posedge clk);
#1;data_in = testData6[97];
@(posedge clk);
#1;data_in = testData6[98];
@(posedge clk);
#1;data_in = testData6[99];
@(posedge clk);
#1;data_in = testData6[100];
@(posedge clk);
#1;data_in = testData6[101];
@(posedge clk);
#1;data_in = testData6[102];
@(posedge clk);
#1;data_in = testData6[103];
@(posedge clk);
#1;data_in = testData6[104];
@(posedge clk);
#1;data_in = testData6[105];
@(posedge clk);
#1;data_in = testData6[106];
@(posedge clk);
#1;data_in = testData6[107];
@(posedge clk);
#1;data_in = testData6[108];
@(posedge clk);
#1;data_in = testData6[109];
@(posedge clk);
#1;data_in = testData6[110];
@(posedge clk);
#1;data_in = testData6[111];
@(posedge clk);
#1;data_in = testData6[112];
@(posedge clk);
#1;data_in = testData6[113];
@(posedge clk);
#1;data_in = testData6[114];
@(posedge clk);
#1;data_in = testData6[115];
@(posedge clk);
#1;data_in = testData6[116];
@(posedge clk);
#1;data_in = testData6[117];
@(posedge clk);
#1;data_in = testData6[118];
@(posedge clk);
#1;data_in = testData6[119];
@(posedge clk);
#1;data_in = testData6[120];
@(posedge clk);
#1;data_in = testData6[121];
@(posedge clk);
#1;data_in = testData6[122];
@(posedge clk);
#1;data_in = testData6[123];
@(posedge clk);
#1;data_in = testData6[124];
@(posedge clk);
#1;data_in = testData6[125];
@(posedge clk);
#1;data_in = testData6[126];
@(posedge clk);
#1;data_in = testData6[127];
@(posedge clk);
#1;data_in = testData6[128];
@(posedge clk);
#1;data_in = testData6[129];
@(posedge clk);
#1;data_in = testData6[130];
@(posedge clk);
#1;data_in = testData6[131];
@(posedge clk);
#1;data_in = testData6[132];
@(posedge clk);
#1;data_in = testData6[133];
@(posedge clk);
#1;data_in = testData6[134];
@(posedge clk);
#1;data_in = testData6[135];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[136]; 
@(posedge clk);
#1;data_in = testData6[137];
@(posedge clk);
#1;data_in = testData6[138];
@(posedge clk);
#1;data_in = testData6[139];
@(posedge clk);
#1;data_in = testData6[140];
@(posedge clk);
#1;data_in = testData6[141];
@(posedge clk);
#1;data_in = testData6[142];
@(posedge clk);
#1;data_in = testData6[143];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[144];
@(posedge clk);
#1;data_in = testData6[145];
@(posedge clk);
#1;data_in = testData6[146];
@(posedge clk);
#1;data_in = testData6[147];
@(posedge clk);
#1;data_in = testData6[148];
@(posedge clk);
#1;data_in = testData6[149];
@(posedge clk);
#1;data_in = testData6[150];
@(posedge clk);
#1;data_in = testData6[151];
@(posedge clk);
#1;data_in = testData6[152];
@(posedge clk);
#1;data_in = testData6[153];
@(posedge clk);
#1;data_in = testData6[154];
@(posedge clk);
#1;data_in = testData6[155];
@(posedge clk);
#1;data_in = testData6[156];
@(posedge clk);
#1;data_in = testData6[157];
@(posedge clk);
#1;data_in = testData6[158];
@(posedge clk);
#1;data_in = testData6[159];
@(posedge clk);
#1;data_in = testData6[160];
@(posedge clk);
#1;data_in = testData6[161];
@(posedge clk);
#1;data_in = testData6[162];
@(posedge clk);
#1;data_in = testData6[163];
@(posedge clk);
#1;data_in = testData6[164];
@(posedge clk);
#1;data_in = testData6[165];
@(posedge clk);
#1;data_in = testData6[166];
@(posedge clk);
#1;data_in = testData6[167];
@(posedge clk);
#1;data_in = testData6[168];
@(posedge clk);
#1;data_in = testData6[169];
@(posedge clk);
#1;data_in = testData6[170];
@(posedge clk);
#1;data_in = testData6[171];
@(posedge clk);
#1;data_in = testData6[172];
@(posedge clk);
#1;data_in = testData6[173];
@(posedge clk);
#1;data_in = testData6[174];
@(posedge clk);
#1;data_in = testData6[175];
@(posedge clk);
#1;data_in = testData6[176];
@(posedge clk);
#1;data_in = testData6[177];
@(posedge clk);
#1;data_in = testData6[178];
@(posedge clk);
#1;data_in = testData6[179];
@(posedge clk);
#1;data_in = testData6[180];
@(posedge clk);
#1;data_in = testData6[181];
@(posedge clk);
#1;data_in = testData6[182];
@(posedge clk);
#1;data_in = testData6[183];
@(posedge clk);
#1;data_in = testData6[184];
@(posedge clk);
#1;data_in = testData6[185];
@(posedge clk);
#1;data_in = testData6[186];
@(posedge clk);
#1;data_in = testData6[187];
@(posedge clk);
#1;data_in = testData6[188];
@(posedge clk);
#1;data_in = testData6[189];
@(posedge clk);
#1;data_in = testData6[190];
@(posedge clk);
#1;data_in = testData6[191];
@(posedge clk);
#1;data_in = testData6[192];
@(posedge clk);
#1;data_in = testData6[193];
@(posedge clk);
#1;data_in = testData6[194];
@(posedge clk);
#1;data_in = testData6[195];
@(posedge clk);
#1;data_in = testData6[196];
@(posedge clk);
#1;data_in = testData6[197];
@(posedge clk);
#1;data_in = testData6[198];
@(posedge clk);
#1;data_in = testData6[199];
@(posedge clk);
#1;data_in = testData6[200];
@(posedge clk);
#1;data_in = testData6[201];
@(posedge clk);
#1;data_in = testData6[202];
@(posedge clk);
#1;data_in = testData6[203];
@(posedge clk);
#1;data_in = testData6[204];
@(posedge clk);
#1;data_in = testData6[205];
@(posedge clk);
#1;data_in = testData6[206];
@(posedge clk);
#1;data_in = testData6[207];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[208]; 
@(posedge clk);
#1;data_in = testData6[209];
@(posedge clk);
#1;data_in = testData6[210];
@(posedge clk);
#1;data_in = testData6[211];
@(posedge clk);
#1;data_in = testData6[212];
@(posedge clk);
#1;data_in = testData6[213];
@(posedge clk);
#1;data_in = testData6[214];
@(posedge clk);
#1;data_in = testData6[215];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[216];
@(posedge clk);
#1;data_in = testData6[217];
@(posedge clk);
#1;data_in = testData6[218];
@(posedge clk);
#1;data_in = testData6[219];
@(posedge clk);
#1;data_in = testData6[220];
@(posedge clk);
#1;data_in = testData6[221];
@(posedge clk);
#1;data_in = testData6[222];
@(posedge clk);
#1;data_in = testData6[223];
@(posedge clk);
#1;data_in = testData6[224];
@(posedge clk);
#1;data_in = testData6[225];
@(posedge clk);
#1;data_in = testData6[226];
@(posedge clk);
#1;data_in = testData6[227];
@(posedge clk);
#1;data_in = testData6[228];
@(posedge clk);
#1;data_in = testData6[229];
@(posedge clk);
#1;data_in = testData6[230];
@(posedge clk);
#1;data_in = testData6[231];
@(posedge clk);
#1;data_in = testData6[232];
@(posedge clk);
#1;data_in = testData6[233];
@(posedge clk);
#1;data_in = testData6[234];
@(posedge clk);
#1;data_in = testData6[235];
@(posedge clk);
#1;data_in = testData6[236];
@(posedge clk);
#1;data_in = testData6[237];
@(posedge clk);
#1;data_in = testData6[238];
@(posedge clk);
#1;data_in = testData6[239];
@(posedge clk);
#1;data_in = testData6[240];
@(posedge clk);
#1;data_in = testData6[241];
@(posedge clk);
#1;data_in = testData6[242];
@(posedge clk);
#1;data_in = testData6[243];
@(posedge clk);
#1;data_in = testData6[244];
@(posedge clk);
#1;data_in = testData6[245];
@(posedge clk);
#1;data_in = testData6[246];
@(posedge clk);
#1;data_in = testData6[247];
@(posedge clk);
#1;data_in = testData6[248];
@(posedge clk);
#1;data_in = testData6[249];
@(posedge clk);
#1;data_in = testData6[250];
@(posedge clk);
#1;data_in = testData6[251];
@(posedge clk);
#1;data_in = testData6[252];
@(posedge clk);
#1;data_in = testData6[253];
@(posedge clk);
#1;data_in = testData6[254];
@(posedge clk);
#1;data_in = testData6[255];
@(posedge clk);
#1;data_in = testData6[256];
@(posedge clk);
#1;data_in = testData6[257];
@(posedge clk);
#1;data_in = testData6[258];
@(posedge clk);
#1;data_in = testData6[259];
@(posedge clk);
#1;data_in = testData6[260];
@(posedge clk);
#1;data_in = testData6[261];
@(posedge clk);
#1;data_in = testData6[262];
@(posedge clk);
#1;data_in = testData6[263];
@(posedge clk);
#1;data_in = testData6[264];
@(posedge clk);
#1;data_in = testData6[265];
@(posedge clk);
#1;data_in = testData6[266];
@(posedge clk);
#1;data_in = testData6[267];
@(posedge clk);
#1;data_in = testData6[268];
@(posedge clk);
#1;data_in = testData6[269];
@(posedge clk);
#1;data_in = testData6[270];
@(posedge clk);
#1;data_in = testData6[271];
@(posedge clk);
#1;data_in = testData6[272];
@(posedge clk);
#1;data_in = testData6[273];
@(posedge clk);
#1;data_in = testData6[274];
@(posedge clk);
#1;data_in = testData6[275];
@(posedge clk);
#1;data_in = testData6[276];
@(posedge clk);
#1;data_in = testData6[277];
@(posedge clk);
#1;data_in = testData6[278];
@(posedge clk);
#1;data_in = testData6[279];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[280]; 
@(posedge clk);
#1;data_in = testData6[281];
@(posedge clk);
#1;data_in = testData6[282];
@(posedge clk);
#1;data_in = testData6[283];
@(posedge clk);
#1;data_in = testData6[284];
@(posedge clk);
#1;data_in = testData6[285];
@(posedge clk);
#1;data_in = testData6[286];
@(posedge clk);
#1;data_in = testData6[287];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[288];
@(posedge clk);
#1;data_in = testData6[289];
@(posedge clk);
#1;data_in = testData6[290];
@(posedge clk);
#1;data_in = testData6[291];
@(posedge clk);
#1;data_in = testData6[292];
@(posedge clk);
#1;data_in = testData6[293];
@(posedge clk);
#1;data_in = testData6[294];
@(posedge clk);
#1;data_in = testData6[295];
@(posedge clk);
#1;data_in = testData6[296];
@(posedge clk);
#1;data_in = testData6[297];
@(posedge clk);
#1;data_in = testData6[298];
@(posedge clk);
#1;data_in = testData6[299];
@(posedge clk);
#1;data_in = testData6[300];
@(posedge clk);
#1;data_in = testData6[301];
@(posedge clk);
#1;data_in = testData6[302];
@(posedge clk);
#1;data_in = testData6[303];
@(posedge clk);
#1;data_in = testData6[304];
@(posedge clk);
#1;data_in = testData6[305];
@(posedge clk);
#1;data_in = testData6[306];
@(posedge clk);
#1;data_in = testData6[307];
@(posedge clk);
#1;data_in = testData6[308];
@(posedge clk);
#1;data_in = testData6[309];
@(posedge clk);
#1;data_in = testData6[310];
@(posedge clk);
#1;data_in = testData6[311];
@(posedge clk);
#1;data_in = testData6[312];
@(posedge clk);
#1;data_in = testData6[313];
@(posedge clk);
#1;data_in = testData6[314];
@(posedge clk);
#1;data_in = testData6[315];
@(posedge clk);
#1;data_in = testData6[316];
@(posedge clk);
#1;data_in = testData6[317];
@(posedge clk);
#1;data_in = testData6[318];
@(posedge clk);
#1;data_in = testData6[319];
@(posedge clk);
#1;data_in = testData6[320];
@(posedge clk);
#1;data_in = testData6[321];
@(posedge clk);
#1;data_in = testData6[322];
@(posedge clk);
#1;data_in = testData6[323];
@(posedge clk);
#1;data_in = testData6[324];
@(posedge clk);
#1;data_in = testData6[325];
@(posedge clk);
#1;data_in = testData6[326];
@(posedge clk);
#1;data_in = testData6[327];
@(posedge clk);
#1;data_in = testData6[328];
@(posedge clk);
#1;data_in = testData6[329];
@(posedge clk);
#1;data_in = testData6[330];
@(posedge clk);
#1;data_in = testData6[331];
@(posedge clk);
#1;data_in = testData6[332];
@(posedge clk);
#1;data_in = testData6[333];
@(posedge clk);
#1;data_in = testData6[334];
@(posedge clk);
#1;data_in = testData6[335];
@(posedge clk);
#1;data_in = testData6[336];
@(posedge clk);
#1;data_in = testData6[337];
@(posedge clk);
#1;data_in = testData6[338];
@(posedge clk);
#1;data_in = testData6[339];
@(posedge clk);
#1;data_in = testData6[340];
@(posedge clk);
#1;data_in = testData6[341];
@(posedge clk);
#1;data_in = testData6[342];
@(posedge clk);
#1;data_in = testData6[343];
@(posedge clk);
#1;data_in = testData6[344];
@(posedge clk);
#1;data_in = testData6[345];
@(posedge clk);
#1;data_in = testData6[346];
@(posedge clk);
#1;data_in = testData6[347];
@(posedge clk);
#1;data_in = testData6[348];
@(posedge clk);
#1;data_in = testData6[349];
@(posedge clk);
#1;data_in = testData6[350];
@(posedge clk);
#1;data_in = testData6[351];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[352]; 
@(posedge clk);
#1;data_in = testData6[353];
@(posedge clk);
#1;data_in = testData6[354];
@(posedge clk);
#1;data_in = testData6[355];
@(posedge clk);
#1;data_in = testData6[356];
@(posedge clk);
#1;data_in = testData6[357];
@(posedge clk);
#1;data_in = testData6[358];
@(posedge clk);
#1;data_in = testData6[359];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[360];
@(posedge clk);
#1;data_in = testData6[361];
@(posedge clk);
#1;data_in = testData6[362];
@(posedge clk);
#1;data_in = testData6[363];
@(posedge clk);
#1;data_in = testData6[364];
@(posedge clk);
#1;data_in = testData6[365];
@(posedge clk);
#1;data_in = testData6[366];
@(posedge clk);
#1;data_in = testData6[367];
@(posedge clk);
#1;data_in = testData6[368];
@(posedge clk);
#1;data_in = testData6[369];
@(posedge clk);
#1;data_in = testData6[370];
@(posedge clk);
#1;data_in = testData6[371];
@(posedge clk);
#1;data_in = testData6[372];
@(posedge clk);
#1;data_in = testData6[373];
@(posedge clk);
#1;data_in = testData6[374];
@(posedge clk);
#1;data_in = testData6[375];
@(posedge clk);
#1;data_in = testData6[376];
@(posedge clk);
#1;data_in = testData6[377];
@(posedge clk);
#1;data_in = testData6[378];
@(posedge clk);
#1;data_in = testData6[379];
@(posedge clk);
#1;data_in = testData6[380];
@(posedge clk);
#1;data_in = testData6[381];
@(posedge clk);
#1;data_in = testData6[382];
@(posedge clk);
#1;data_in = testData6[383];
@(posedge clk);
#1;data_in = testData6[384];
@(posedge clk);
#1;data_in = testData6[385];
@(posedge clk);
#1;data_in = testData6[386];
@(posedge clk);
#1;data_in = testData6[387];
@(posedge clk);
#1;data_in = testData6[388];
@(posedge clk);
#1;data_in = testData6[389];
@(posedge clk);
#1;data_in = testData6[390];
@(posedge clk);
#1;data_in = testData6[391];
@(posedge clk);
#1;data_in = testData6[392];
@(posedge clk);
#1;data_in = testData6[393];
@(posedge clk);
#1;data_in = testData6[394];
@(posedge clk);
#1;data_in = testData6[395];
@(posedge clk);
#1;data_in = testData6[396];
@(posedge clk);
#1;data_in = testData6[397];
@(posedge clk);
#1;data_in = testData6[398];
@(posedge clk);
#1;data_in = testData6[399];
@(posedge clk);
#1;data_in = testData6[400];
@(posedge clk);
#1;data_in = testData6[401];
@(posedge clk);
#1;data_in = testData6[402];
@(posedge clk);
#1;data_in = testData6[403];
@(posedge clk);
#1;data_in = testData6[404];
@(posedge clk);
#1;data_in = testData6[405];
@(posedge clk);
#1;data_in = testData6[406];
@(posedge clk);
#1;data_in = testData6[407];
@(posedge clk);
#1;data_in = testData6[408];
@(posedge clk);
#1;data_in = testData6[409];
@(posedge clk);
#1;data_in = testData6[410];
@(posedge clk);
#1;data_in = testData6[411];
@(posedge clk);
#1;data_in = testData6[412];
@(posedge clk);
#1;data_in = testData6[413];
@(posedge clk);
#1;data_in = testData6[414];
@(posedge clk);
#1;data_in = testData6[415];
@(posedge clk);
#1;data_in = testData6[416];
@(posedge clk);
#1;data_in = testData6[417];
@(posedge clk);
#1;data_in = testData6[418];
@(posedge clk);
#1;data_in = testData6[419];
@(posedge clk);
#1;data_in = testData6[420];
@(posedge clk);
#1;data_in = testData6[421];
@(posedge clk);
#1;data_in = testData6[422];
@(posedge clk);
#1;data_in = testData6[423];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[424]; 
@(posedge clk);
#1;data_in = testData6[425];
@(posedge clk);
#1;data_in = testData6[426];
@(posedge clk);
#1;data_in = testData6[427];
@(posedge clk);
#1;data_in = testData6[428];
@(posedge clk);
#1;data_in = testData6[429];
@(posedge clk);
#1;data_in = testData6[430];
@(posedge clk);
#1;data_in = testData6[431];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[432];
@(posedge clk);
#1;data_in = testData6[433];
@(posedge clk);
#1;data_in = testData6[434];
@(posedge clk);
#1;data_in = testData6[435];
@(posedge clk);
#1;data_in = testData6[436];
@(posedge clk);
#1;data_in = testData6[437];
@(posedge clk);
#1;data_in = testData6[438];
@(posedge clk);
#1;data_in = testData6[439];
@(posedge clk);
#1;data_in = testData6[440];
@(posedge clk);
#1;data_in = testData6[441];
@(posedge clk);
#1;data_in = testData6[442];
@(posedge clk);
#1;data_in = testData6[443];
@(posedge clk);
#1;data_in = testData6[444];
@(posedge clk);
#1;data_in = testData6[445];
@(posedge clk);
#1;data_in = testData6[446];
@(posedge clk);
#1;data_in = testData6[447];
@(posedge clk);
#1;data_in = testData6[448];
@(posedge clk);
#1;data_in = testData6[449];
@(posedge clk);
#1;data_in = testData6[450];
@(posedge clk);
#1;data_in = testData6[451];
@(posedge clk);
#1;data_in = testData6[452];
@(posedge clk);
#1;data_in = testData6[453];
@(posedge clk);
#1;data_in = testData6[454];
@(posedge clk);
#1;data_in = testData6[455];
@(posedge clk);
#1;data_in = testData6[456];
@(posedge clk);
#1;data_in = testData6[457];
@(posedge clk);
#1;data_in = testData6[458];
@(posedge clk);
#1;data_in = testData6[459];
@(posedge clk);
#1;data_in = testData6[460];
@(posedge clk);
#1;data_in = testData6[461];
@(posedge clk);
#1;data_in = testData6[462];
@(posedge clk);
#1;data_in = testData6[463];
@(posedge clk);
#1;data_in = testData6[464];
@(posedge clk);
#1;data_in = testData6[465];
@(posedge clk);
#1;data_in = testData6[466];
@(posedge clk);
#1;data_in = testData6[467];
@(posedge clk);
#1;data_in = testData6[468];
@(posedge clk);
#1;data_in = testData6[469];
@(posedge clk);
#1;data_in = testData6[470];
@(posedge clk);
#1;data_in = testData6[471];
@(posedge clk);
#1;data_in = testData6[472];
@(posedge clk);
#1;data_in = testData6[473];
@(posedge clk);
#1;data_in = testData6[474];
@(posedge clk);
#1;data_in = testData6[475];
@(posedge clk);
#1;data_in = testData6[476];
@(posedge clk);
#1;data_in = testData6[477];
@(posedge clk);
#1;data_in = testData6[478];
@(posedge clk);
#1;data_in = testData6[479];
@(posedge clk);
#1;data_in = testData6[480];
@(posedge clk);
#1;data_in = testData6[481];
@(posedge clk);
#1;data_in = testData6[482];
@(posedge clk);
#1;data_in = testData6[483];
@(posedge clk);
#1;data_in = testData6[484];
@(posedge clk);
#1;data_in = testData6[485];
@(posedge clk);
#1;data_in = testData6[486];
@(posedge clk);
#1;data_in = testData6[487];
@(posedge clk);
#1;data_in = testData6[488];
@(posedge clk);
#1;data_in = testData6[489];
@(posedge clk);
#1;data_in = testData6[490];
@(posedge clk);
#1;data_in = testData6[491];
@(posedge clk);
#1;data_in = testData6[492];
@(posedge clk);
#1;data_in = testData6[493];
@(posedge clk);
#1;data_in = testData6[494];
@(posedge clk);
#1;data_in = testData6[495];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[496]; 
@(posedge clk);
#1;data_in = testData6[497];
@(posedge clk);
#1;data_in = testData6[498];
@(posedge clk);
#1;data_in = testData6[499];
@(posedge clk);
#1;data_in = testData6[500];
@(posedge clk);
#1;data_in = testData6[501];
@(posedge clk);
#1;data_in = testData6[502];
@(posedge clk);
#1;data_in = testData6[503];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[504];
@(posedge clk);
#1;data_in = testData6[505];
@(posedge clk);
#1;data_in = testData6[506];
@(posedge clk);
#1;data_in = testData6[507];
@(posedge clk);
#1;data_in = testData6[508];
@(posedge clk);
#1;data_in = testData6[509];
@(posedge clk);
#1;data_in = testData6[510];
@(posedge clk);
#1;data_in = testData6[511];
@(posedge clk);
#1;data_in = testData6[512];
@(posedge clk);
#1;data_in = testData6[513];
@(posedge clk);
#1;data_in = testData6[514];
@(posedge clk);
#1;data_in = testData6[515];
@(posedge clk);
#1;data_in = testData6[516];
@(posedge clk);
#1;data_in = testData6[517];
@(posedge clk);
#1;data_in = testData6[518];
@(posedge clk);
#1;data_in = testData6[519];
@(posedge clk);
#1;data_in = testData6[520];
@(posedge clk);
#1;data_in = testData6[521];
@(posedge clk);
#1;data_in = testData6[522];
@(posedge clk);
#1;data_in = testData6[523];
@(posedge clk);
#1;data_in = testData6[524];
@(posedge clk);
#1;data_in = testData6[525];
@(posedge clk);
#1;data_in = testData6[526];
@(posedge clk);
#1;data_in = testData6[527];
@(posedge clk);
#1;data_in = testData6[528];
@(posedge clk);
#1;data_in = testData6[529];
@(posedge clk);
#1;data_in = testData6[530];
@(posedge clk);
#1;data_in = testData6[531];
@(posedge clk);
#1;data_in = testData6[532];
@(posedge clk);
#1;data_in = testData6[533];
@(posedge clk);
#1;data_in = testData6[534];
@(posedge clk);
#1;data_in = testData6[535];
@(posedge clk);
#1;data_in = testData6[536];
@(posedge clk);
#1;data_in = testData6[537];
@(posedge clk);
#1;data_in = testData6[538];
@(posedge clk);
#1;data_in = testData6[539];
@(posedge clk);
#1;data_in = testData6[540];
@(posedge clk);
#1;data_in = testData6[541];
@(posedge clk);
#1;data_in = testData6[542];
@(posedge clk);
#1;data_in = testData6[543];
@(posedge clk);
#1;data_in = testData6[544];
@(posedge clk);
#1;data_in = testData6[545];
@(posedge clk);
#1;data_in = testData6[546];
@(posedge clk);
#1;data_in = testData6[547];
@(posedge clk);
#1;data_in = testData6[548];
@(posedge clk);
#1;data_in = testData6[549];
@(posedge clk);
#1;data_in = testData6[550];
@(posedge clk);
#1;data_in = testData6[551];
@(posedge clk);
#1;data_in = testData6[552];
@(posedge clk);
#1;data_in = testData6[553];
@(posedge clk);
#1;data_in = testData6[554];
@(posedge clk);
#1;data_in = testData6[555];
@(posedge clk);
#1;data_in = testData6[556];
@(posedge clk);
#1;data_in = testData6[557];
@(posedge clk);
#1;data_in = testData6[558];
@(posedge clk);
#1;data_in = testData6[559];
@(posedge clk);
#1;data_in = testData6[560];
@(posedge clk);
#1;data_in = testData6[561];
@(posedge clk);
#1;data_in = testData6[562];
@(posedge clk);
#1;data_in = testData6[563];
@(posedge clk);
#1;data_in = testData6[564];
@(posedge clk);
#1;data_in = testData6[565];
@(posedge clk);
#1;data_in = testData6[566];
@(posedge clk);
#1;data_in = testData6[567];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[568]; 
@(posedge clk);
#1;data_in = testData6[569];
@(posedge clk);
#1;data_in = testData6[570];
@(posedge clk);
#1;data_in = testData6[571];
@(posedge clk);
#1;data_in = testData6[572];
@(posedge clk);
#1;data_in = testData6[573];
@(posedge clk);
#1;data_in = testData6[574];
@(posedge clk);
#1;data_in = testData6[575];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[576];
@(posedge clk);
#1;data_in = testData6[577];
@(posedge clk);
#1;data_in = testData6[578];
@(posedge clk);
#1;data_in = testData6[579];
@(posedge clk);
#1;data_in = testData6[580];
@(posedge clk);
#1;data_in = testData6[581];
@(posedge clk);
#1;data_in = testData6[582];
@(posedge clk);
#1;data_in = testData6[583];
@(posedge clk);
#1;data_in = testData6[584];
@(posedge clk);
#1;data_in = testData6[585];
@(posedge clk);
#1;data_in = testData6[586];
@(posedge clk);
#1;data_in = testData6[587];
@(posedge clk);
#1;data_in = testData6[588];
@(posedge clk);
#1;data_in = testData6[589];
@(posedge clk);
#1;data_in = testData6[590];
@(posedge clk);
#1;data_in = testData6[591];
@(posedge clk);
#1;data_in = testData6[592];
@(posedge clk);
#1;data_in = testData6[593];
@(posedge clk);
#1;data_in = testData6[594];
@(posedge clk);
#1;data_in = testData6[595];
@(posedge clk);
#1;data_in = testData6[596];
@(posedge clk);
#1;data_in = testData6[597];
@(posedge clk);
#1;data_in = testData6[598];
@(posedge clk);
#1;data_in = testData6[599];
@(posedge clk);
#1;data_in = testData6[600];
@(posedge clk);
#1;data_in = testData6[601];
@(posedge clk);
#1;data_in = testData6[602];
@(posedge clk);
#1;data_in = testData6[603];
@(posedge clk);
#1;data_in = testData6[604];
@(posedge clk);
#1;data_in = testData6[605];
@(posedge clk);
#1;data_in = testData6[606];
@(posedge clk);
#1;data_in = testData6[607];
@(posedge clk);
#1;data_in = testData6[608];
@(posedge clk);
#1;data_in = testData6[609];
@(posedge clk);
#1;data_in = testData6[610];
@(posedge clk);
#1;data_in = testData6[611];
@(posedge clk);
#1;data_in = testData6[612];
@(posedge clk);
#1;data_in = testData6[613];
@(posedge clk);
#1;data_in = testData6[614];
@(posedge clk);
#1;data_in = testData6[615];
@(posedge clk);
#1;data_in = testData6[616];
@(posedge clk);
#1;data_in = testData6[617];
@(posedge clk);
#1;data_in = testData6[618];
@(posedge clk);
#1;data_in = testData6[619];
@(posedge clk);
#1;data_in = testData6[620];
@(posedge clk);
#1;data_in = testData6[621];
@(posedge clk);
#1;data_in = testData6[622];
@(posedge clk);
#1;data_in = testData6[623];
@(posedge clk);
#1;data_in = testData6[624];
@(posedge clk);
#1;data_in = testData6[625];
@(posedge clk);
#1;data_in = testData6[626];
@(posedge clk);
#1;data_in = testData6[627];
@(posedge clk);
#1;data_in = testData6[628];
@(posedge clk);
#1;data_in = testData6[629];
@(posedge clk);
#1;data_in = testData6[630];
@(posedge clk);
#1;data_in = testData6[631];
@(posedge clk);
#1;data_in = testData6[632];
@(posedge clk);
#1;data_in = testData6[633];
@(posedge clk);
#1;data_in = testData6[634];
@(posedge clk);
#1;data_in = testData6[635];
@(posedge clk);
#1;data_in = testData6[636];
@(posedge clk);
#1;data_in = testData6[637];
@(posedge clk);
#1;data_in = testData6[638];
@(posedge clk);
#1;data_in = testData6[639];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[640]; 
@(posedge clk);
#1;data_in = testData6[641];
@(posedge clk);
#1;data_in = testData6[642];
@(posedge clk);
#1;data_in = testData6[643];
@(posedge clk);
#1;data_in = testData6[644];
@(posedge clk);
#1;data_in = testData6[645];
@(posedge clk);
#1;data_in = testData6[646];
@(posedge clk);
#1;data_in = testData6[647];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[648];
@(posedge clk);
#1;data_in = testData6[649];
@(posedge clk);
#1;data_in = testData6[650];
@(posedge clk);
#1;data_in = testData6[651];
@(posedge clk);
#1;data_in = testData6[652];
@(posedge clk);
#1;data_in = testData6[653];
@(posedge clk);
#1;data_in = testData6[654];
@(posedge clk);
#1;data_in = testData6[655];
@(posedge clk);
#1;data_in = testData6[656];
@(posedge clk);
#1;data_in = testData6[657];
@(posedge clk);
#1;data_in = testData6[658];
@(posedge clk);
#1;data_in = testData6[659];
@(posedge clk);
#1;data_in = testData6[660];
@(posedge clk);
#1;data_in = testData6[661];
@(posedge clk);
#1;data_in = testData6[662];
@(posedge clk);
#1;data_in = testData6[663];
@(posedge clk);
#1;data_in = testData6[664];
@(posedge clk);
#1;data_in = testData6[665];
@(posedge clk);
#1;data_in = testData6[666];
@(posedge clk);
#1;data_in = testData6[667];
@(posedge clk);
#1;data_in = testData6[668];
@(posedge clk);
#1;data_in = testData6[669];
@(posedge clk);
#1;data_in = testData6[670];
@(posedge clk);
#1;data_in = testData6[671];
@(posedge clk);
#1;data_in = testData6[672];
@(posedge clk);
#1;data_in = testData6[673];
@(posedge clk);
#1;data_in = testData6[674];
@(posedge clk);
#1;data_in = testData6[675];
@(posedge clk);
#1;data_in = testData6[676];
@(posedge clk);
#1;data_in = testData6[677];
@(posedge clk);
#1;data_in = testData6[678];
@(posedge clk);
#1;data_in = testData6[679];
@(posedge clk);
#1;data_in = testData6[680];
@(posedge clk);
#1;data_in = testData6[681];
@(posedge clk);
#1;data_in = testData6[682];
@(posedge clk);
#1;data_in = testData6[683];
@(posedge clk);
#1;data_in = testData6[684];
@(posedge clk);
#1;data_in = testData6[685];
@(posedge clk);
#1;data_in = testData6[686];
@(posedge clk);
#1;data_in = testData6[687];
@(posedge clk);
#1;data_in = testData6[688];
@(posedge clk);
#1;data_in = testData6[689];
@(posedge clk);
#1;data_in = testData6[690];
@(posedge clk);
#1;data_in = testData6[691];
@(posedge clk);
#1;data_in = testData6[692];
@(posedge clk);
#1;data_in = testData6[693];
@(posedge clk);
#1;data_in = testData6[694];
@(posedge clk);
#1;data_in = testData6[695];
@(posedge clk);
#1;data_in = testData6[696];
@(posedge clk);
#1;data_in = testData6[697];
@(posedge clk);
#1;data_in = testData6[698];
@(posedge clk);
#1;data_in = testData6[699];
@(posedge clk);
#1;data_in = testData6[700];
@(posedge clk);
#1;data_in = testData6[701];
@(posedge clk);
#1;data_in = testData6[702];
@(posedge clk);
#1;data_in = testData6[703];
@(posedge clk);
#1;data_in = testData6[704];
@(posedge clk);
#1;data_in = testData6[705];
@(posedge clk);
#1;data_in = testData6[706];
@(posedge clk);
#1;data_in = testData6[707];
@(posedge clk);
#1;data_in = testData6[708];
@(posedge clk);
#1;data_in = testData6[709];
@(posedge clk);
#1;data_in = testData6[710];
@(posedge clk);
#1;data_in = testData6[711];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[712]; 
@(posedge clk);
#1;data_in = testData6[713];
@(posedge clk);
#1;data_in = testData6[714];
@(posedge clk);
#1;data_in = testData6[715];
@(posedge clk);
#1;data_in = testData6[716];
@(posedge clk);
#1;data_in = testData6[717];
@(posedge clk);
#1;data_in = testData6[718];
@(posedge clk);
#1;data_in = testData6[719];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[720];
@(posedge clk);
#1;data_in = testData6[721];
@(posedge clk);
#1;data_in = testData6[722];
@(posedge clk);
#1;data_in = testData6[723];
@(posedge clk);
#1;data_in = testData6[724];
@(posedge clk);
#1;data_in = testData6[725];
@(posedge clk);
#1;data_in = testData6[726];
@(posedge clk);
#1;data_in = testData6[727];
@(posedge clk);
#1;data_in = testData6[728];
@(posedge clk);
#1;data_in = testData6[729];
@(posedge clk);
#1;data_in = testData6[730];
@(posedge clk);
#1;data_in = testData6[731];
@(posedge clk);
#1;data_in = testData6[732];
@(posedge clk);
#1;data_in = testData6[733];
@(posedge clk);
#1;data_in = testData6[734];
@(posedge clk);
#1;data_in = testData6[735];
@(posedge clk);
#1;data_in = testData6[736];
@(posedge clk);
#1;data_in = testData6[737];
@(posedge clk);
#1;data_in = testData6[738];
@(posedge clk);
#1;data_in = testData6[739];
@(posedge clk);
#1;data_in = testData6[740];
@(posedge clk);
#1;data_in = testData6[741];
@(posedge clk);
#1;data_in = testData6[742];
@(posedge clk);
#1;data_in = testData6[743];
@(posedge clk);
#1;data_in = testData6[744];
@(posedge clk);
#1;data_in = testData6[745];
@(posedge clk);
#1;data_in = testData6[746];
@(posedge clk);
#1;data_in = testData6[747];
@(posedge clk);
#1;data_in = testData6[748];
@(posedge clk);
#1;data_in = testData6[749];
@(posedge clk);
#1;data_in = testData6[750];
@(posedge clk);
#1;data_in = testData6[751];
@(posedge clk);
#1;data_in = testData6[752];
@(posedge clk);
#1;data_in = testData6[753];
@(posedge clk);
#1;data_in = testData6[754];
@(posedge clk);
#1;data_in = testData6[755];
@(posedge clk);
#1;data_in = testData6[756];
@(posedge clk);
#1;data_in = testData6[757];
@(posedge clk);
#1;data_in = testData6[758];
@(posedge clk);
#1;data_in = testData6[759];
@(posedge clk);
#1;data_in = testData6[760];
@(posedge clk);
#1;data_in = testData6[761];
@(posedge clk);
#1;data_in = testData6[762];
@(posedge clk);
#1;data_in = testData6[763];
@(posedge clk);
#1;data_in = testData6[764];
@(posedge clk);
#1;data_in = testData6[765];
@(posedge clk);
#1;data_in = testData6[766];
@(posedge clk);
#1;data_in = testData6[767];
@(posedge clk);
#1;data_in = testData6[768];
@(posedge clk);
#1;data_in = testData6[769];
@(posedge clk);
#1;data_in = testData6[770];
@(posedge clk);
#1;data_in = testData6[771];
@(posedge clk);
#1;data_in = testData6[772];
@(posedge clk);
#1;data_in = testData6[773];
@(posedge clk);
#1;data_in = testData6[774];
@(posedge clk);
#1;data_in = testData6[775];
@(posedge clk);
#1;data_in = testData6[776];
@(posedge clk);
#1;data_in = testData6[777];
@(posedge clk);
#1;data_in = testData6[778];
@(posedge clk);
#1;data_in = testData6[779];
@(posedge clk);
#1;data_in = testData6[780];
@(posedge clk);
#1;data_in = testData6[781];
@(posedge clk);
#1;data_in = testData6[782];
@(posedge clk);
#1;data_in = testData6[783];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[784]; 
@(posedge clk);
#1;data_in = testData6[785];
@(posedge clk);
#1;data_in = testData6[786];
@(posedge clk);
#1;data_in = testData6[787];
@(posedge clk);
#1;data_in = testData6[788];
@(posedge clk);
#1;data_in = testData6[789];
@(posedge clk);
#1;data_in = testData6[790];
@(posedge clk);
#1;data_in = testData6[791];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[792];
@(posedge clk);
#1;data_in = testData6[793];
@(posedge clk);
#1;data_in = testData6[794];
@(posedge clk);
#1;data_in = testData6[795];
@(posedge clk);
#1;data_in = testData6[796];
@(posedge clk);
#1;data_in = testData6[797];
@(posedge clk);
#1;data_in = testData6[798];
@(posedge clk);
#1;data_in = testData6[799];
@(posedge clk);
#1;data_in = testData6[800];
@(posedge clk);
#1;data_in = testData6[801];
@(posedge clk);
#1;data_in = testData6[802];
@(posedge clk);
#1;data_in = testData6[803];
@(posedge clk);
#1;data_in = testData6[804];
@(posedge clk);
#1;data_in = testData6[805];
@(posedge clk);
#1;data_in = testData6[806];
@(posedge clk);
#1;data_in = testData6[807];
@(posedge clk);
#1;data_in = testData6[808];
@(posedge clk);
#1;data_in = testData6[809];
@(posedge clk);
#1;data_in = testData6[810];
@(posedge clk);
#1;data_in = testData6[811];
@(posedge clk);
#1;data_in = testData6[812];
@(posedge clk);
#1;data_in = testData6[813];
@(posedge clk);
#1;data_in = testData6[814];
@(posedge clk);
#1;data_in = testData6[815];
@(posedge clk);
#1;data_in = testData6[816];
@(posedge clk);
#1;data_in = testData6[817];
@(posedge clk);
#1;data_in = testData6[818];
@(posedge clk);
#1;data_in = testData6[819];
@(posedge clk);
#1;data_in = testData6[820];
@(posedge clk);
#1;data_in = testData6[821];
@(posedge clk);
#1;data_in = testData6[822];
@(posedge clk);
#1;data_in = testData6[823];
@(posedge clk);
#1;data_in = testData6[824];
@(posedge clk);
#1;data_in = testData6[825];
@(posedge clk);
#1;data_in = testData6[826];
@(posedge clk);
#1;data_in = testData6[827];
@(posedge clk);
#1;data_in = testData6[828];
@(posedge clk);
#1;data_in = testData6[829];
@(posedge clk);
#1;data_in = testData6[830];
@(posedge clk);
#1;data_in = testData6[831];
@(posedge clk);
#1;data_in = testData6[832];
@(posedge clk);
#1;data_in = testData6[833];
@(posedge clk);
#1;data_in = testData6[834];
@(posedge clk);
#1;data_in = testData6[835];
@(posedge clk);
#1;data_in = testData6[836];
@(posedge clk);
#1;data_in = testData6[837];
@(posedge clk);
#1;data_in = testData6[838];
@(posedge clk);
#1;data_in = testData6[839];
@(posedge clk);
#1;data_in = testData6[840];
@(posedge clk);
#1;data_in = testData6[841];
@(posedge clk);
#1;data_in = testData6[842];
@(posedge clk);
#1;data_in = testData6[843];
@(posedge clk);
#1;data_in = testData6[844];
@(posedge clk);
#1;data_in = testData6[845];
@(posedge clk);
#1;data_in = testData6[846];
@(posedge clk);
#1;data_in = testData6[847];
@(posedge clk);
#1;data_in = testData6[848];
@(posedge clk);
#1;data_in = testData6[849];
@(posedge clk);
#1;data_in = testData6[850];
@(posedge clk);
#1;data_in = testData6[851];
@(posedge clk);
#1;data_in = testData6[852];
@(posedge clk);
#1;data_in = testData6[853];
@(posedge clk);
#1;data_in = testData6[854];
@(posedge clk);
#1;data_in = testData6[855];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[856]; 
@(posedge clk);
#1;data_in = testData6[857];
@(posedge clk);
#1;data_in = testData6[858];
@(posedge clk);
#1;data_in = testData6[859];
@(posedge clk);
#1;data_in = testData6[860];
@(posedge clk);
#1;data_in = testData6[861];
@(posedge clk);
#1;data_in = testData6[862];
@(posedge clk);
#1;data_in = testData6[863];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[864];
@(posedge clk);
#1;data_in = testData6[865];
@(posedge clk);
#1;data_in = testData6[866];
@(posedge clk);
#1;data_in = testData6[867];
@(posedge clk);
#1;data_in = testData6[868];
@(posedge clk);
#1;data_in = testData6[869];
@(posedge clk);
#1;data_in = testData6[870];
@(posedge clk);
#1;data_in = testData6[871];
@(posedge clk);
#1;data_in = testData6[872];
@(posedge clk);
#1;data_in = testData6[873];
@(posedge clk);
#1;data_in = testData6[874];
@(posedge clk);
#1;data_in = testData6[875];
@(posedge clk);
#1;data_in = testData6[876];
@(posedge clk);
#1;data_in = testData6[877];
@(posedge clk);
#1;data_in = testData6[878];
@(posedge clk);
#1;data_in = testData6[879];
@(posedge clk);
#1;data_in = testData6[880];
@(posedge clk);
#1;data_in = testData6[881];
@(posedge clk);
#1;data_in = testData6[882];
@(posedge clk);
#1;data_in = testData6[883];
@(posedge clk);
#1;data_in = testData6[884];
@(posedge clk);
#1;data_in = testData6[885];
@(posedge clk);
#1;data_in = testData6[886];
@(posedge clk);
#1;data_in = testData6[887];
@(posedge clk);
#1;data_in = testData6[888];
@(posedge clk);
#1;data_in = testData6[889];
@(posedge clk);
#1;data_in = testData6[890];
@(posedge clk);
#1;data_in = testData6[891];
@(posedge clk);
#1;data_in = testData6[892];
@(posedge clk);
#1;data_in = testData6[893];
@(posedge clk);
#1;data_in = testData6[894];
@(posedge clk);
#1;data_in = testData6[895];
@(posedge clk);
#1;data_in = testData6[896];
@(posedge clk);
#1;data_in = testData6[897];
@(posedge clk);
#1;data_in = testData6[898];
@(posedge clk);
#1;data_in = testData6[899];
@(posedge clk);
#1;data_in = testData6[900];
@(posedge clk);
#1;data_in = testData6[901];
@(posedge clk);
#1;data_in = testData6[902];
@(posedge clk);
#1;data_in = testData6[903];
@(posedge clk);
#1;data_in = testData6[904];
@(posedge clk);
#1;data_in = testData6[905];
@(posedge clk);
#1;data_in = testData6[906];
@(posedge clk);
#1;data_in = testData6[907];
@(posedge clk);
#1;data_in = testData6[908];
@(posedge clk);
#1;data_in = testData6[909];
@(posedge clk);
#1;data_in = testData6[910];
@(posedge clk);
#1;data_in = testData6[911];
@(posedge clk);
#1;data_in = testData6[912];
@(posedge clk);
#1;data_in = testData6[913];
@(posedge clk);
#1;data_in = testData6[914];
@(posedge clk);
#1;data_in = testData6[915];
@(posedge clk);
#1;data_in = testData6[916];
@(posedge clk);
#1;data_in = testData6[917];
@(posedge clk);
#1;data_in = testData6[918];
@(posedge clk);
#1;data_in = testData6[919];
@(posedge clk);
#1;data_in = testData6[920];
@(posedge clk);
#1;data_in = testData6[921];
@(posedge clk);
#1;data_in = testData6[922];
@(posedge clk);
#1;data_in = testData6[923];
@(posedge clk);
#1;data_in = testData6[924];
@(posedge clk);
#1;data_in = testData6[925];
@(posedge clk);
#1;data_in = testData6[926];
@(posedge clk);
#1;data_in = testData6[927];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[928]; 
@(posedge clk);
#1;data_in = testData6[929];
@(posedge clk);
#1;data_in = testData6[930];
@(posedge clk);
#1;data_in = testData6[931];
@(posedge clk);
#1;data_in = testData6[932];
@(posedge clk);
#1;data_in = testData6[933];
@(posedge clk);
#1;data_in = testData6[934];
@(posedge clk);
#1;data_in = testData6[935];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[936];
@(posedge clk);
#1;data_in = testData6[937];
@(posedge clk);
#1;data_in = testData6[938];
@(posedge clk);
#1;data_in = testData6[939];
@(posedge clk);
#1;data_in = testData6[940];
@(posedge clk);
#1;data_in = testData6[941];
@(posedge clk);
#1;data_in = testData6[942];
@(posedge clk);
#1;data_in = testData6[943];
@(posedge clk);
#1;data_in = testData6[944];
@(posedge clk);
#1;data_in = testData6[945];
@(posedge clk);
#1;data_in = testData6[946];
@(posedge clk);
#1;data_in = testData6[947];
@(posedge clk);
#1;data_in = testData6[948];
@(posedge clk);
#1;data_in = testData6[949];
@(posedge clk);
#1;data_in = testData6[950];
@(posedge clk);
#1;data_in = testData6[951];
@(posedge clk);
#1;data_in = testData6[952];
@(posedge clk);
#1;data_in = testData6[953];
@(posedge clk);
#1;data_in = testData6[954];
@(posedge clk);
#1;data_in = testData6[955];
@(posedge clk);
#1;data_in = testData6[956];
@(posedge clk);
#1;data_in = testData6[957];
@(posedge clk);
#1;data_in = testData6[958];
@(posedge clk);
#1;data_in = testData6[959];
@(posedge clk);
#1;data_in = testData6[960];
@(posedge clk);
#1;data_in = testData6[961];
@(posedge clk);
#1;data_in = testData6[962];
@(posedge clk);
#1;data_in = testData6[963];
@(posedge clk);
#1;data_in = testData6[964];
@(posedge clk);
#1;data_in = testData6[965];
@(posedge clk);
#1;data_in = testData6[966];
@(posedge clk);
#1;data_in = testData6[967];
@(posedge clk);
#1;data_in = testData6[968];
@(posedge clk);
#1;data_in = testData6[969];
@(posedge clk);
#1;data_in = testData6[970];
@(posedge clk);
#1;data_in = testData6[971];
@(posedge clk);
#1;data_in = testData6[972];
@(posedge clk);
#1;data_in = testData6[973];
@(posedge clk);
#1;data_in = testData6[974];
@(posedge clk);
#1;data_in = testData6[975];
@(posedge clk);
#1;data_in = testData6[976];
@(posedge clk);
#1;data_in = testData6[977];
@(posedge clk);
#1;data_in = testData6[978];
@(posedge clk);
#1;data_in = testData6[979];
@(posedge clk);
#1;data_in = testData6[980];
@(posedge clk);
#1;data_in = testData6[981];
@(posedge clk);
#1;data_in = testData6[982];
@(posedge clk);
#1;data_in = testData6[983];
@(posedge clk);
#1;data_in = testData6[984];
@(posedge clk);
#1;data_in = testData6[985];
@(posedge clk);
#1;data_in = testData6[986];
@(posedge clk);
#1;data_in = testData6[987];
@(posedge clk);
#1;data_in = testData6[988];
@(posedge clk);
#1;data_in = testData6[989];
@(posedge clk);
#1;data_in = testData6[990];
@(posedge clk);
#1;data_in = testData6[991];
@(posedge clk);
#1;data_in = testData6[992];
@(posedge clk);
#1;data_in = testData6[993];
@(posedge clk);
#1;data_in = testData6[994];
@(posedge clk);
#1;data_in = testData6[995];
@(posedge clk);
#1;data_in = testData6[996];
@(posedge clk);
#1;data_in = testData6[997];
@(posedge clk);
#1;data_in = testData6[998];
@(posedge clk);
#1;data_in = testData6[999];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1000]; 
@(posedge clk);
#1;data_in = testData6[1001];
@(posedge clk);
#1;data_in = testData6[1002];
@(posedge clk);
#1;data_in = testData6[1003];
@(posedge clk);
#1;data_in = testData6[1004];
@(posedge clk);
#1;data_in = testData6[1005];
@(posedge clk);
#1;data_in = testData6[1006];
@(posedge clk);
#1;data_in = testData6[1007];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1008];
@(posedge clk);
#1;data_in = testData6[1009];
@(posedge clk);
#1;data_in = testData6[1010];
@(posedge clk);
#1;data_in = testData6[1011];
@(posedge clk);
#1;data_in = testData6[1012];
@(posedge clk);
#1;data_in = testData6[1013];
@(posedge clk);
#1;data_in = testData6[1014];
@(posedge clk);
#1;data_in = testData6[1015];
@(posedge clk);
#1;data_in = testData6[1016];
@(posedge clk);
#1;data_in = testData6[1017];
@(posedge clk);
#1;data_in = testData6[1018];
@(posedge clk);
#1;data_in = testData6[1019];
@(posedge clk);
#1;data_in = testData6[1020];
@(posedge clk);
#1;data_in = testData6[1021];
@(posedge clk);
#1;data_in = testData6[1022];
@(posedge clk);
#1;data_in = testData6[1023];
@(posedge clk);
#1;data_in = testData6[1024];
@(posedge clk);
#1;data_in = testData6[1025];
@(posedge clk);
#1;data_in = testData6[1026];
@(posedge clk);
#1;data_in = testData6[1027];
@(posedge clk);
#1;data_in = testData6[1028];
@(posedge clk);
#1;data_in = testData6[1029];
@(posedge clk);
#1;data_in = testData6[1030];
@(posedge clk);
#1;data_in = testData6[1031];
@(posedge clk);
#1;data_in = testData6[1032];
@(posedge clk);
#1;data_in = testData6[1033];
@(posedge clk);
#1;data_in = testData6[1034];
@(posedge clk);
#1;data_in = testData6[1035];
@(posedge clk);
#1;data_in = testData6[1036];
@(posedge clk);
#1;data_in = testData6[1037];
@(posedge clk);
#1;data_in = testData6[1038];
@(posedge clk);
#1;data_in = testData6[1039];
@(posedge clk);
#1;data_in = testData6[1040];
@(posedge clk);
#1;data_in = testData6[1041];
@(posedge clk);
#1;data_in = testData6[1042];
@(posedge clk);
#1;data_in = testData6[1043];
@(posedge clk);
#1;data_in = testData6[1044];
@(posedge clk);
#1;data_in = testData6[1045];
@(posedge clk);
#1;data_in = testData6[1046];
@(posedge clk);
#1;data_in = testData6[1047];
@(posedge clk);
#1;data_in = testData6[1048];
@(posedge clk);
#1;data_in = testData6[1049];
@(posedge clk);
#1;data_in = testData6[1050];
@(posedge clk);
#1;data_in = testData6[1051];
@(posedge clk);
#1;data_in = testData6[1052];
@(posedge clk);
#1;data_in = testData6[1053];
@(posedge clk);
#1;data_in = testData6[1054];
@(posedge clk);
#1;data_in = testData6[1055];
@(posedge clk);
#1;data_in = testData6[1056];
@(posedge clk);
#1;data_in = testData6[1057];
@(posedge clk);
#1;data_in = testData6[1058];
@(posedge clk);
#1;data_in = testData6[1059];
@(posedge clk);
#1;data_in = testData6[1060];
@(posedge clk);
#1;data_in = testData6[1061];
@(posedge clk);
#1;data_in = testData6[1062];
@(posedge clk);
#1;data_in = testData6[1063];
@(posedge clk);
#1;data_in = testData6[1064];
@(posedge clk);
#1;data_in = testData6[1065];
@(posedge clk);
#1;data_in = testData6[1066];
@(posedge clk);
#1;data_in = testData6[1067];
@(posedge clk);
#1;data_in = testData6[1068];
@(posedge clk);
#1;data_in = testData6[1069];
@(posedge clk);
#1;data_in = testData6[1070];
@(posedge clk);
#1;data_in = testData6[1071];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1072]; 
@(posedge clk);
#1;data_in = testData6[1073];
@(posedge clk);
#1;data_in = testData6[1074];
@(posedge clk);
#1;data_in = testData6[1075];
@(posedge clk);
#1;data_in = testData6[1076];
@(posedge clk);
#1;data_in = testData6[1077];
@(posedge clk);
#1;data_in = testData6[1078];
@(posedge clk);
#1;data_in = testData6[1079];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1080];
@(posedge clk);
#1;data_in = testData6[1081];
@(posedge clk);
#1;data_in = testData6[1082];
@(posedge clk);
#1;data_in = testData6[1083];
@(posedge clk);
#1;data_in = testData6[1084];
@(posedge clk);
#1;data_in = testData6[1085];
@(posedge clk);
#1;data_in = testData6[1086];
@(posedge clk);
#1;data_in = testData6[1087];
@(posedge clk);
#1;data_in = testData6[1088];
@(posedge clk);
#1;data_in = testData6[1089];
@(posedge clk);
#1;data_in = testData6[1090];
@(posedge clk);
#1;data_in = testData6[1091];
@(posedge clk);
#1;data_in = testData6[1092];
@(posedge clk);
#1;data_in = testData6[1093];
@(posedge clk);
#1;data_in = testData6[1094];
@(posedge clk);
#1;data_in = testData6[1095];
@(posedge clk);
#1;data_in = testData6[1096];
@(posedge clk);
#1;data_in = testData6[1097];
@(posedge clk);
#1;data_in = testData6[1098];
@(posedge clk);
#1;data_in = testData6[1099];
@(posedge clk);
#1;data_in = testData6[1100];
@(posedge clk);
#1;data_in = testData6[1101];
@(posedge clk);
#1;data_in = testData6[1102];
@(posedge clk);
#1;data_in = testData6[1103];
@(posedge clk);
#1;data_in = testData6[1104];
@(posedge clk);
#1;data_in = testData6[1105];
@(posedge clk);
#1;data_in = testData6[1106];
@(posedge clk);
#1;data_in = testData6[1107];
@(posedge clk);
#1;data_in = testData6[1108];
@(posedge clk);
#1;data_in = testData6[1109];
@(posedge clk);
#1;data_in = testData6[1110];
@(posedge clk);
#1;data_in = testData6[1111];
@(posedge clk);
#1;data_in = testData6[1112];
@(posedge clk);
#1;data_in = testData6[1113];
@(posedge clk);
#1;data_in = testData6[1114];
@(posedge clk);
#1;data_in = testData6[1115];
@(posedge clk);
#1;data_in = testData6[1116];
@(posedge clk);
#1;data_in = testData6[1117];
@(posedge clk);
#1;data_in = testData6[1118];
@(posedge clk);
#1;data_in = testData6[1119];
@(posedge clk);
#1;data_in = testData6[1120];
@(posedge clk);
#1;data_in = testData6[1121];
@(posedge clk);
#1;data_in = testData6[1122];
@(posedge clk);
#1;data_in = testData6[1123];
@(posedge clk);
#1;data_in = testData6[1124];
@(posedge clk);
#1;data_in = testData6[1125];
@(posedge clk);
#1;data_in = testData6[1126];
@(posedge clk);
#1;data_in = testData6[1127];
@(posedge clk);
#1;data_in = testData6[1128];
@(posedge clk);
#1;data_in = testData6[1129];
@(posedge clk);
#1;data_in = testData6[1130];
@(posedge clk);
#1;data_in = testData6[1131];
@(posedge clk);
#1;data_in = testData6[1132];
@(posedge clk);
#1;data_in = testData6[1133];
@(posedge clk);
#1;data_in = testData6[1134];
@(posedge clk);
#1;data_in = testData6[1135];
@(posedge clk);
#1;data_in = testData6[1136];
@(posedge clk);
#1;data_in = testData6[1137];
@(posedge clk);
#1;data_in = testData6[1138];
@(posedge clk);
#1;data_in = testData6[1139];
@(posedge clk);
#1;data_in = testData6[1140];
@(posedge clk);
#1;data_in = testData6[1141];
@(posedge clk);
#1;data_in = testData6[1142];
@(posedge clk);
#1;data_in = testData6[1143];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1144]; 
@(posedge clk);
#1;data_in = testData6[1145];
@(posedge clk);
#1;data_in = testData6[1146];
@(posedge clk);
#1;data_in = testData6[1147];
@(posedge clk);
#1;data_in = testData6[1148];
@(posedge clk);
#1;data_in = testData6[1149];
@(posedge clk);
#1;data_in = testData6[1150];
@(posedge clk);
#1;data_in = testData6[1151];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1152];
@(posedge clk);
#1;data_in = testData6[1153];
@(posedge clk);
#1;data_in = testData6[1154];
@(posedge clk);
#1;data_in = testData6[1155];
@(posedge clk);
#1;data_in = testData6[1156];
@(posedge clk);
#1;data_in = testData6[1157];
@(posedge clk);
#1;data_in = testData6[1158];
@(posedge clk);
#1;data_in = testData6[1159];
@(posedge clk);
#1;data_in = testData6[1160];
@(posedge clk);
#1;data_in = testData6[1161];
@(posedge clk);
#1;data_in = testData6[1162];
@(posedge clk);
#1;data_in = testData6[1163];
@(posedge clk);
#1;data_in = testData6[1164];
@(posedge clk);
#1;data_in = testData6[1165];
@(posedge clk);
#1;data_in = testData6[1166];
@(posedge clk);
#1;data_in = testData6[1167];
@(posedge clk);
#1;data_in = testData6[1168];
@(posedge clk);
#1;data_in = testData6[1169];
@(posedge clk);
#1;data_in = testData6[1170];
@(posedge clk);
#1;data_in = testData6[1171];
@(posedge clk);
#1;data_in = testData6[1172];
@(posedge clk);
#1;data_in = testData6[1173];
@(posedge clk);
#1;data_in = testData6[1174];
@(posedge clk);
#1;data_in = testData6[1175];
@(posedge clk);
#1;data_in = testData6[1176];
@(posedge clk);
#1;data_in = testData6[1177];
@(posedge clk);
#1;data_in = testData6[1178];
@(posedge clk);
#1;data_in = testData6[1179];
@(posedge clk);
#1;data_in = testData6[1180];
@(posedge clk);
#1;data_in = testData6[1181];
@(posedge clk);
#1;data_in = testData6[1182];
@(posedge clk);
#1;data_in = testData6[1183];
@(posedge clk);
#1;data_in = testData6[1184];
@(posedge clk);
#1;data_in = testData6[1185];
@(posedge clk);
#1;data_in = testData6[1186];
@(posedge clk);
#1;data_in = testData6[1187];
@(posedge clk);
#1;data_in = testData6[1188];
@(posedge clk);
#1;data_in = testData6[1189];
@(posedge clk);
#1;data_in = testData6[1190];
@(posedge clk);
#1;data_in = testData6[1191];
@(posedge clk);
#1;data_in = testData6[1192];
@(posedge clk);
#1;data_in = testData6[1193];
@(posedge clk);
#1;data_in = testData6[1194];
@(posedge clk);
#1;data_in = testData6[1195];
@(posedge clk);
#1;data_in = testData6[1196];
@(posedge clk);
#1;data_in = testData6[1197];
@(posedge clk);
#1;data_in = testData6[1198];
@(posedge clk);
#1;data_in = testData6[1199];
@(posedge clk);
#1;data_in = testData6[1200];
@(posedge clk);
#1;data_in = testData6[1201];
@(posedge clk);
#1;data_in = testData6[1202];
@(posedge clk);
#1;data_in = testData6[1203];
@(posedge clk);
#1;data_in = testData6[1204];
@(posedge clk);
#1;data_in = testData6[1205];
@(posedge clk);
#1;data_in = testData6[1206];
@(posedge clk);
#1;data_in = testData6[1207];
@(posedge clk);
#1;data_in = testData6[1208];
@(posedge clk);
#1;data_in = testData6[1209];
@(posedge clk);
#1;data_in = testData6[1210];
@(posedge clk);
#1;data_in = testData6[1211];
@(posedge clk);
#1;data_in = testData6[1212];
@(posedge clk);
#1;data_in = testData6[1213];
@(posedge clk);
#1;data_in = testData6[1214];
@(posedge clk);
#1;data_in = testData6[1215];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1216]; 
@(posedge clk);
#1;data_in = testData6[1217];
@(posedge clk);
#1;data_in = testData6[1218];
@(posedge clk);
#1;data_in = testData6[1219];
@(posedge clk);
#1;data_in = testData6[1220];
@(posedge clk);
#1;data_in = testData6[1221];
@(posedge clk);
#1;data_in = testData6[1222];
@(posedge clk);
#1;data_in = testData6[1223];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1224];
@(posedge clk);
#1;data_in = testData6[1225];
@(posedge clk);
#1;data_in = testData6[1226];
@(posedge clk);
#1;data_in = testData6[1227];
@(posedge clk);
#1;data_in = testData6[1228];
@(posedge clk);
#1;data_in = testData6[1229];
@(posedge clk);
#1;data_in = testData6[1230];
@(posedge clk);
#1;data_in = testData6[1231];
@(posedge clk);
#1;data_in = testData6[1232];
@(posedge clk);
#1;data_in = testData6[1233];
@(posedge clk);
#1;data_in = testData6[1234];
@(posedge clk);
#1;data_in = testData6[1235];
@(posedge clk);
#1;data_in = testData6[1236];
@(posedge clk);
#1;data_in = testData6[1237];
@(posedge clk);
#1;data_in = testData6[1238];
@(posedge clk);
#1;data_in = testData6[1239];
@(posedge clk);
#1;data_in = testData6[1240];
@(posedge clk);
#1;data_in = testData6[1241];
@(posedge clk);
#1;data_in = testData6[1242];
@(posedge clk);
#1;data_in = testData6[1243];
@(posedge clk);
#1;data_in = testData6[1244];
@(posedge clk);
#1;data_in = testData6[1245];
@(posedge clk);
#1;data_in = testData6[1246];
@(posedge clk);
#1;data_in = testData6[1247];
@(posedge clk);
#1;data_in = testData6[1248];
@(posedge clk);
#1;data_in = testData6[1249];
@(posedge clk);
#1;data_in = testData6[1250];
@(posedge clk);
#1;data_in = testData6[1251];
@(posedge clk);
#1;data_in = testData6[1252];
@(posedge clk);
#1;data_in = testData6[1253];
@(posedge clk);
#1;data_in = testData6[1254];
@(posedge clk);
#1;data_in = testData6[1255];
@(posedge clk);
#1;data_in = testData6[1256];
@(posedge clk);
#1;data_in = testData6[1257];
@(posedge clk);
#1;data_in = testData6[1258];
@(posedge clk);
#1;data_in = testData6[1259];
@(posedge clk);
#1;data_in = testData6[1260];
@(posedge clk);
#1;data_in = testData6[1261];
@(posedge clk);
#1;data_in = testData6[1262];
@(posedge clk);
#1;data_in = testData6[1263];
@(posedge clk);
#1;data_in = testData6[1264];
@(posedge clk);
#1;data_in = testData6[1265];
@(posedge clk);
#1;data_in = testData6[1266];
@(posedge clk);
#1;data_in = testData6[1267];
@(posedge clk);
#1;data_in = testData6[1268];
@(posedge clk);
#1;data_in = testData6[1269];
@(posedge clk);
#1;data_in = testData6[1270];
@(posedge clk);
#1;data_in = testData6[1271];
@(posedge clk);
#1;data_in = testData6[1272];
@(posedge clk);
#1;data_in = testData6[1273];
@(posedge clk);
#1;data_in = testData6[1274];
@(posedge clk);
#1;data_in = testData6[1275];
@(posedge clk);
#1;data_in = testData6[1276];
@(posedge clk);
#1;data_in = testData6[1277];
@(posedge clk);
#1;data_in = testData6[1278];
@(posedge clk);
#1;data_in = testData6[1279];
@(posedge clk);
#1;data_in = testData6[1280];
@(posedge clk);
#1;data_in = testData6[1281];
@(posedge clk);
#1;data_in = testData6[1282];
@(posedge clk);
#1;data_in = testData6[1283];
@(posedge clk);
#1;data_in = testData6[1284];
@(posedge clk);
#1;data_in = testData6[1285];
@(posedge clk);
#1;data_in = testData6[1286];
@(posedge clk);
#1;data_in = testData6[1287];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1288]; 
@(posedge clk);
#1;data_in = testData6[1289];
@(posedge clk);
#1;data_in = testData6[1290];
@(posedge clk);
#1;data_in = testData6[1291];
@(posedge clk);
#1;data_in = testData6[1292];
@(posedge clk);
#1;data_in = testData6[1293];
@(posedge clk);
#1;data_in = testData6[1294];
@(posedge clk);
#1;data_in = testData6[1295];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1296];
@(posedge clk);
#1;data_in = testData6[1297];
@(posedge clk);
#1;data_in = testData6[1298];
@(posedge clk);
#1;data_in = testData6[1299];
@(posedge clk);
#1;data_in = testData6[1300];
@(posedge clk);
#1;data_in = testData6[1301];
@(posedge clk);
#1;data_in = testData6[1302];
@(posedge clk);
#1;data_in = testData6[1303];
@(posedge clk);
#1;data_in = testData6[1304];
@(posedge clk);
#1;data_in = testData6[1305];
@(posedge clk);
#1;data_in = testData6[1306];
@(posedge clk);
#1;data_in = testData6[1307];
@(posedge clk);
#1;data_in = testData6[1308];
@(posedge clk);
#1;data_in = testData6[1309];
@(posedge clk);
#1;data_in = testData6[1310];
@(posedge clk);
#1;data_in = testData6[1311];
@(posedge clk);
#1;data_in = testData6[1312];
@(posedge clk);
#1;data_in = testData6[1313];
@(posedge clk);
#1;data_in = testData6[1314];
@(posedge clk);
#1;data_in = testData6[1315];
@(posedge clk);
#1;data_in = testData6[1316];
@(posedge clk);
#1;data_in = testData6[1317];
@(posedge clk);
#1;data_in = testData6[1318];
@(posedge clk);
#1;data_in = testData6[1319];
@(posedge clk);
#1;data_in = testData6[1320];
@(posedge clk);
#1;data_in = testData6[1321];
@(posedge clk);
#1;data_in = testData6[1322];
@(posedge clk);
#1;data_in = testData6[1323];
@(posedge clk);
#1;data_in = testData6[1324];
@(posedge clk);
#1;data_in = testData6[1325];
@(posedge clk);
#1;data_in = testData6[1326];
@(posedge clk);
#1;data_in = testData6[1327];
@(posedge clk);
#1;data_in = testData6[1328];
@(posedge clk);
#1;data_in = testData6[1329];
@(posedge clk);
#1;data_in = testData6[1330];
@(posedge clk);
#1;data_in = testData6[1331];
@(posedge clk);
#1;data_in = testData6[1332];
@(posedge clk);
#1;data_in = testData6[1333];
@(posedge clk);
#1;data_in = testData6[1334];
@(posedge clk);
#1;data_in = testData6[1335];
@(posedge clk);
#1;data_in = testData6[1336];
@(posedge clk);
#1;data_in = testData6[1337];
@(posedge clk);
#1;data_in = testData6[1338];
@(posedge clk);
#1;data_in = testData6[1339];
@(posedge clk);
#1;data_in = testData6[1340];
@(posedge clk);
#1;data_in = testData6[1341];
@(posedge clk);
#1;data_in = testData6[1342];
@(posedge clk);
#1;data_in = testData6[1343];
@(posedge clk);
#1;data_in = testData6[1344];
@(posedge clk);
#1;data_in = testData6[1345];
@(posedge clk);
#1;data_in = testData6[1346];
@(posedge clk);
#1;data_in = testData6[1347];
@(posedge clk);
#1;data_in = testData6[1348];
@(posedge clk);
#1;data_in = testData6[1349];
@(posedge clk);
#1;data_in = testData6[1350];
@(posedge clk);
#1;data_in = testData6[1351];
@(posedge clk);
#1;data_in = testData6[1352];
@(posedge clk);
#1;data_in = testData6[1353];
@(posedge clk);
#1;data_in = testData6[1354];
@(posedge clk);
#1;data_in = testData6[1355];
@(posedge clk);
#1;data_in = testData6[1356];
@(posedge clk);
#1;data_in = testData6[1357];
@(posedge clk);
#1;data_in = testData6[1358];
@(posedge clk);
#1;data_in = testData6[1359];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1360]; 
@(posedge clk);
#1;data_in = testData6[1361];
@(posedge clk);
#1;data_in = testData6[1362];
@(posedge clk);
#1;data_in = testData6[1363];
@(posedge clk);
#1;data_in = testData6[1364];
@(posedge clk);
#1;data_in = testData6[1365];
@(posedge clk);
#1;data_in = testData6[1366];
@(posedge clk);
#1;data_in = testData6[1367];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1368];
@(posedge clk);
#1;data_in = testData6[1369];
@(posedge clk);
#1;data_in = testData6[1370];
@(posedge clk);
#1;data_in = testData6[1371];
@(posedge clk);
#1;data_in = testData6[1372];
@(posedge clk);
#1;data_in = testData6[1373];
@(posedge clk);
#1;data_in = testData6[1374];
@(posedge clk);
#1;data_in = testData6[1375];
@(posedge clk);
#1;data_in = testData6[1376];
@(posedge clk);
#1;data_in = testData6[1377];
@(posedge clk);
#1;data_in = testData6[1378];
@(posedge clk);
#1;data_in = testData6[1379];
@(posedge clk);
#1;data_in = testData6[1380];
@(posedge clk);
#1;data_in = testData6[1381];
@(posedge clk);
#1;data_in = testData6[1382];
@(posedge clk);
#1;data_in = testData6[1383];
@(posedge clk);
#1;data_in = testData6[1384];
@(posedge clk);
#1;data_in = testData6[1385];
@(posedge clk);
#1;data_in = testData6[1386];
@(posedge clk);
#1;data_in = testData6[1387];
@(posedge clk);
#1;data_in = testData6[1388];
@(posedge clk);
#1;data_in = testData6[1389];
@(posedge clk);
#1;data_in = testData6[1390];
@(posedge clk);
#1;data_in = testData6[1391];
@(posedge clk);
#1;data_in = testData6[1392];
@(posedge clk);
#1;data_in = testData6[1393];
@(posedge clk);
#1;data_in = testData6[1394];
@(posedge clk);
#1;data_in = testData6[1395];
@(posedge clk);
#1;data_in = testData6[1396];
@(posedge clk);
#1;data_in = testData6[1397];
@(posedge clk);
#1;data_in = testData6[1398];
@(posedge clk);
#1;data_in = testData6[1399];
@(posedge clk);
#1;data_in = testData6[1400];
@(posedge clk);
#1;data_in = testData6[1401];
@(posedge clk);
#1;data_in = testData6[1402];
@(posedge clk);
#1;data_in = testData6[1403];
@(posedge clk);
#1;data_in = testData6[1404];
@(posedge clk);
#1;data_in = testData6[1405];
@(posedge clk);
#1;data_in = testData6[1406];
@(posedge clk);
#1;data_in = testData6[1407];
@(posedge clk);
#1;data_in = testData6[1408];
@(posedge clk);
#1;data_in = testData6[1409];
@(posedge clk);
#1;data_in = testData6[1410];
@(posedge clk);
#1;data_in = testData6[1411];
@(posedge clk);
#1;data_in = testData6[1412];
@(posedge clk);
#1;data_in = testData6[1413];
@(posedge clk);
#1;data_in = testData6[1414];
@(posedge clk);
#1;data_in = testData6[1415];
@(posedge clk);
#1;data_in = testData6[1416];
@(posedge clk);
#1;data_in = testData6[1417];
@(posedge clk);
#1;data_in = testData6[1418];
@(posedge clk);
#1;data_in = testData6[1419];
@(posedge clk);
#1;data_in = testData6[1420];
@(posedge clk);
#1;data_in = testData6[1421];
@(posedge clk);
#1;data_in = testData6[1422];
@(posedge clk);
#1;data_in = testData6[1423];
@(posedge clk);
#1;data_in = testData6[1424];
@(posedge clk);
#1;data_in = testData6[1425];
@(posedge clk);
#1;data_in = testData6[1426];
@(posedge clk);
#1;data_in = testData6[1427];
@(posedge clk);
#1;data_in = testData6[1428];
@(posedge clk);
#1;data_in = testData6[1429];
@(posedge clk);
#1;data_in = testData6[1430];
@(posedge clk);
#1;data_in = testData6[1431];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1432]; 
@(posedge clk);
#1;data_in = testData6[1433];
@(posedge clk);
#1;data_in = testData6[1434];
@(posedge clk);
#1;data_in = testData6[1435];
@(posedge clk);
#1;data_in = testData6[1436];
@(posedge clk);
#1;data_in = testData6[1437];
@(posedge clk);
#1;data_in = testData6[1438];
@(posedge clk);
#1;data_in = testData6[1439];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1440];
@(posedge clk);
#1;data_in = testData6[1441];
@(posedge clk);
#1;data_in = testData6[1442];
@(posedge clk);
#1;data_in = testData6[1443];
@(posedge clk);
#1;data_in = testData6[1444];
@(posedge clk);
#1;data_in = testData6[1445];
@(posedge clk);
#1;data_in = testData6[1446];
@(posedge clk);
#1;data_in = testData6[1447];
@(posedge clk);
#1;data_in = testData6[1448];
@(posedge clk);
#1;data_in = testData6[1449];
@(posedge clk);
#1;data_in = testData6[1450];
@(posedge clk);
#1;data_in = testData6[1451];
@(posedge clk);
#1;data_in = testData6[1452];
@(posedge clk);
#1;data_in = testData6[1453];
@(posedge clk);
#1;data_in = testData6[1454];
@(posedge clk);
#1;data_in = testData6[1455];
@(posedge clk);
#1;data_in = testData6[1456];
@(posedge clk);
#1;data_in = testData6[1457];
@(posedge clk);
#1;data_in = testData6[1458];
@(posedge clk);
#1;data_in = testData6[1459];
@(posedge clk);
#1;data_in = testData6[1460];
@(posedge clk);
#1;data_in = testData6[1461];
@(posedge clk);
#1;data_in = testData6[1462];
@(posedge clk);
#1;data_in = testData6[1463];
@(posedge clk);
#1;data_in = testData6[1464];
@(posedge clk);
#1;data_in = testData6[1465];
@(posedge clk);
#1;data_in = testData6[1466];
@(posedge clk);
#1;data_in = testData6[1467];
@(posedge clk);
#1;data_in = testData6[1468];
@(posedge clk);
#1;data_in = testData6[1469];
@(posedge clk);
#1;data_in = testData6[1470];
@(posedge clk);
#1;data_in = testData6[1471];
@(posedge clk);
#1;data_in = testData6[1472];
@(posedge clk);
#1;data_in = testData6[1473];
@(posedge clk);
#1;data_in = testData6[1474];
@(posedge clk);
#1;data_in = testData6[1475];
@(posedge clk);
#1;data_in = testData6[1476];
@(posedge clk);
#1;data_in = testData6[1477];
@(posedge clk);
#1;data_in = testData6[1478];
@(posedge clk);
#1;data_in = testData6[1479];
@(posedge clk);
#1;data_in = testData6[1480];
@(posedge clk);
#1;data_in = testData6[1481];
@(posedge clk);
#1;data_in = testData6[1482];
@(posedge clk);
#1;data_in = testData6[1483];
@(posedge clk);
#1;data_in = testData6[1484];
@(posedge clk);
#1;data_in = testData6[1485];
@(posedge clk);
#1;data_in = testData6[1486];
@(posedge clk);
#1;data_in = testData6[1487];
@(posedge clk);
#1;data_in = testData6[1488];
@(posedge clk);
#1;data_in = testData6[1489];
@(posedge clk);
#1;data_in = testData6[1490];
@(posedge clk);
#1;data_in = testData6[1491];
@(posedge clk);
#1;data_in = testData6[1492];
@(posedge clk);
#1;data_in = testData6[1493];
@(posedge clk);
#1;data_in = testData6[1494];
@(posedge clk);
#1;data_in = testData6[1495];
@(posedge clk);
#1;data_in = testData6[1496];
@(posedge clk);
#1;data_in = testData6[1497];
@(posedge clk);
#1;data_in = testData6[1498];
@(posedge clk);
#1;data_in = testData6[1499];
@(posedge clk);
#1;data_in = testData6[1500];
@(posedge clk);
#1;data_in = testData6[1501];
@(posedge clk);
#1;data_in = testData6[1502];
@(posedge clk);
#1;data_in = testData6[1503];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1504]; 
@(posedge clk);
#1;data_in = testData6[1505];
@(posedge clk);
#1;data_in = testData6[1506];
@(posedge clk);
#1;data_in = testData6[1507];
@(posedge clk);
#1;data_in = testData6[1508];
@(posedge clk);
#1;data_in = testData6[1509];
@(posedge clk);
#1;data_in = testData6[1510];
@(posedge clk);
#1;data_in = testData6[1511];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1512];
@(posedge clk);
#1;data_in = testData6[1513];
@(posedge clk);
#1;data_in = testData6[1514];
@(posedge clk);
#1;data_in = testData6[1515];
@(posedge clk);
#1;data_in = testData6[1516];
@(posedge clk);
#1;data_in = testData6[1517];
@(posedge clk);
#1;data_in = testData6[1518];
@(posedge clk);
#1;data_in = testData6[1519];
@(posedge clk);
#1;data_in = testData6[1520];
@(posedge clk);
#1;data_in = testData6[1521];
@(posedge clk);
#1;data_in = testData6[1522];
@(posedge clk);
#1;data_in = testData6[1523];
@(posedge clk);
#1;data_in = testData6[1524];
@(posedge clk);
#1;data_in = testData6[1525];
@(posedge clk);
#1;data_in = testData6[1526];
@(posedge clk);
#1;data_in = testData6[1527];
@(posedge clk);
#1;data_in = testData6[1528];
@(posedge clk);
#1;data_in = testData6[1529];
@(posedge clk);
#1;data_in = testData6[1530];
@(posedge clk);
#1;data_in = testData6[1531];
@(posedge clk);
#1;data_in = testData6[1532];
@(posedge clk);
#1;data_in = testData6[1533];
@(posedge clk);
#1;data_in = testData6[1534];
@(posedge clk);
#1;data_in = testData6[1535];
@(posedge clk);
#1;data_in = testData6[1536];
@(posedge clk);
#1;data_in = testData6[1537];
@(posedge clk);
#1;data_in = testData6[1538];
@(posedge clk);
#1;data_in = testData6[1539];
@(posedge clk);
#1;data_in = testData6[1540];
@(posedge clk);
#1;data_in = testData6[1541];
@(posedge clk);
#1;data_in = testData6[1542];
@(posedge clk);
#1;data_in = testData6[1543];
@(posedge clk);
#1;data_in = testData6[1544];
@(posedge clk);
#1;data_in = testData6[1545];
@(posedge clk);
#1;data_in = testData6[1546];
@(posedge clk);
#1;data_in = testData6[1547];
@(posedge clk);
#1;data_in = testData6[1548];
@(posedge clk);
#1;data_in = testData6[1549];
@(posedge clk);
#1;data_in = testData6[1550];
@(posedge clk);
#1;data_in = testData6[1551];
@(posedge clk);
#1;data_in = testData6[1552];
@(posedge clk);
#1;data_in = testData6[1553];
@(posedge clk);
#1;data_in = testData6[1554];
@(posedge clk);
#1;data_in = testData6[1555];
@(posedge clk);
#1;data_in = testData6[1556];
@(posedge clk);
#1;data_in = testData6[1557];
@(posedge clk);
#1;data_in = testData6[1558];
@(posedge clk);
#1;data_in = testData6[1559];
@(posedge clk);
#1;data_in = testData6[1560];
@(posedge clk);
#1;data_in = testData6[1561];
@(posedge clk);
#1;data_in = testData6[1562];
@(posedge clk);
#1;data_in = testData6[1563];
@(posedge clk);
#1;data_in = testData6[1564];
@(posedge clk);
#1;data_in = testData6[1565];
@(posedge clk);
#1;data_in = testData6[1566];
@(posedge clk);
#1;data_in = testData6[1567];
@(posedge clk);
#1;data_in = testData6[1568];
@(posedge clk);
#1;data_in = testData6[1569];
@(posedge clk);
#1;data_in = testData6[1570];
@(posedge clk);
#1;data_in = testData6[1571];
@(posedge clk);
#1;data_in = testData6[1572];
@(posedge clk);
#1;data_in = testData6[1573];
@(posedge clk);
#1;data_in = testData6[1574];
@(posedge clk);
#1;data_in = testData6[1575];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1576]; 
@(posedge clk);
#1;data_in = testData6[1577];
@(posedge clk);
#1;data_in = testData6[1578];
@(posedge clk);
#1;data_in = testData6[1579];
@(posedge clk);
#1;data_in = testData6[1580];
@(posedge clk);
#1;data_in = testData6[1581];
@(posedge clk);
#1;data_in = testData6[1582];
@(posedge clk);
#1;data_in = testData6[1583];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1584];
@(posedge clk);
#1;data_in = testData6[1585];
@(posedge clk);
#1;data_in = testData6[1586];
@(posedge clk);
#1;data_in = testData6[1587];
@(posedge clk);
#1;data_in = testData6[1588];
@(posedge clk);
#1;data_in = testData6[1589];
@(posedge clk);
#1;data_in = testData6[1590];
@(posedge clk);
#1;data_in = testData6[1591];
@(posedge clk);
#1;data_in = testData6[1592];
@(posedge clk);
#1;data_in = testData6[1593];
@(posedge clk);
#1;data_in = testData6[1594];
@(posedge clk);
#1;data_in = testData6[1595];
@(posedge clk);
#1;data_in = testData6[1596];
@(posedge clk);
#1;data_in = testData6[1597];
@(posedge clk);
#1;data_in = testData6[1598];
@(posedge clk);
#1;data_in = testData6[1599];
@(posedge clk);
#1;data_in = testData6[1600];
@(posedge clk);
#1;data_in = testData6[1601];
@(posedge clk);
#1;data_in = testData6[1602];
@(posedge clk);
#1;data_in = testData6[1603];
@(posedge clk);
#1;data_in = testData6[1604];
@(posedge clk);
#1;data_in = testData6[1605];
@(posedge clk);
#1;data_in = testData6[1606];
@(posedge clk);
#1;data_in = testData6[1607];
@(posedge clk);
#1;data_in = testData6[1608];
@(posedge clk);
#1;data_in = testData6[1609];
@(posedge clk);
#1;data_in = testData6[1610];
@(posedge clk);
#1;data_in = testData6[1611];
@(posedge clk);
#1;data_in = testData6[1612];
@(posedge clk);
#1;data_in = testData6[1613];
@(posedge clk);
#1;data_in = testData6[1614];
@(posedge clk);
#1;data_in = testData6[1615];
@(posedge clk);
#1;data_in = testData6[1616];
@(posedge clk);
#1;data_in = testData6[1617];
@(posedge clk);
#1;data_in = testData6[1618];
@(posedge clk);
#1;data_in = testData6[1619];
@(posedge clk);
#1;data_in = testData6[1620];
@(posedge clk);
#1;data_in = testData6[1621];
@(posedge clk);
#1;data_in = testData6[1622];
@(posedge clk);
#1;data_in = testData6[1623];
@(posedge clk);
#1;data_in = testData6[1624];
@(posedge clk);
#1;data_in = testData6[1625];
@(posedge clk);
#1;data_in = testData6[1626];
@(posedge clk);
#1;data_in = testData6[1627];
@(posedge clk);
#1;data_in = testData6[1628];
@(posedge clk);
#1;data_in = testData6[1629];
@(posedge clk);
#1;data_in = testData6[1630];
@(posedge clk);
#1;data_in = testData6[1631];
@(posedge clk);
#1;data_in = testData6[1632];
@(posedge clk);
#1;data_in = testData6[1633];
@(posedge clk);
#1;data_in = testData6[1634];
@(posedge clk);
#1;data_in = testData6[1635];
@(posedge clk);
#1;data_in = testData6[1636];
@(posedge clk);
#1;data_in = testData6[1637];
@(posedge clk);
#1;data_in = testData6[1638];
@(posedge clk);
#1;data_in = testData6[1639];
@(posedge clk);
#1;data_in = testData6[1640];
@(posedge clk);
#1;data_in = testData6[1641];
@(posedge clk);
#1;data_in = testData6[1642];
@(posedge clk);
#1;data_in = testData6[1643];
@(posedge clk);
#1;data_in = testData6[1644];
@(posedge clk);
#1;data_in = testData6[1645];
@(posedge clk);
#1;data_in = testData6[1646];
@(posedge clk);
#1;data_in = testData6[1647];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1648]; 
@(posedge clk);
#1;data_in = testData6[1649];
@(posedge clk);
#1;data_in = testData6[1650];
@(posedge clk);
#1;data_in = testData6[1651];
@(posedge clk);
#1;data_in = testData6[1652];
@(posedge clk);
#1;data_in = testData6[1653];
@(posedge clk);
#1;data_in = testData6[1654];
@(posedge clk);
#1;data_in = testData6[1655];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1656];
@(posedge clk);
#1;data_in = testData6[1657];
@(posedge clk);
#1;data_in = testData6[1658];
@(posedge clk);
#1;data_in = testData6[1659];
@(posedge clk);
#1;data_in = testData6[1660];
@(posedge clk);
#1;data_in = testData6[1661];
@(posedge clk);
#1;data_in = testData6[1662];
@(posedge clk);
#1;data_in = testData6[1663];
@(posedge clk);
#1;data_in = testData6[1664];
@(posedge clk);
#1;data_in = testData6[1665];
@(posedge clk);
#1;data_in = testData6[1666];
@(posedge clk);
#1;data_in = testData6[1667];
@(posedge clk);
#1;data_in = testData6[1668];
@(posedge clk);
#1;data_in = testData6[1669];
@(posedge clk);
#1;data_in = testData6[1670];
@(posedge clk);
#1;data_in = testData6[1671];
@(posedge clk);
#1;data_in = testData6[1672];
@(posedge clk);
#1;data_in = testData6[1673];
@(posedge clk);
#1;data_in = testData6[1674];
@(posedge clk);
#1;data_in = testData6[1675];
@(posedge clk);
#1;data_in = testData6[1676];
@(posedge clk);
#1;data_in = testData6[1677];
@(posedge clk);
#1;data_in = testData6[1678];
@(posedge clk);
#1;data_in = testData6[1679];
@(posedge clk);
#1;data_in = testData6[1680];
@(posedge clk);
#1;data_in = testData6[1681];
@(posedge clk);
#1;data_in = testData6[1682];
@(posedge clk);
#1;data_in = testData6[1683];
@(posedge clk);
#1;data_in = testData6[1684];
@(posedge clk);
#1;data_in = testData6[1685];
@(posedge clk);
#1;data_in = testData6[1686];
@(posedge clk);
#1;data_in = testData6[1687];
@(posedge clk);
#1;data_in = testData6[1688];
@(posedge clk);
#1;data_in = testData6[1689];
@(posedge clk);
#1;data_in = testData6[1690];
@(posedge clk);
#1;data_in = testData6[1691];
@(posedge clk);
#1;data_in = testData6[1692];
@(posedge clk);
#1;data_in = testData6[1693];
@(posedge clk);
#1;data_in = testData6[1694];
@(posedge clk);
#1;data_in = testData6[1695];
@(posedge clk);
#1;data_in = testData6[1696];
@(posedge clk);
#1;data_in = testData6[1697];
@(posedge clk);
#1;data_in = testData6[1698];
@(posedge clk);
#1;data_in = testData6[1699];
@(posedge clk);
#1;data_in = testData6[1700];
@(posedge clk);
#1;data_in = testData6[1701];
@(posedge clk);
#1;data_in = testData6[1702];
@(posedge clk);
#1;data_in = testData6[1703];
@(posedge clk);
#1;data_in = testData6[1704];
@(posedge clk);
#1;data_in = testData6[1705];
@(posedge clk);
#1;data_in = testData6[1706];
@(posedge clk);
#1;data_in = testData6[1707];
@(posedge clk);
#1;data_in = testData6[1708];
@(posedge clk);
#1;data_in = testData6[1709];
@(posedge clk);
#1;data_in = testData6[1710];
@(posedge clk);
#1;data_in = testData6[1711];
@(posedge clk);
#1;data_in = testData6[1712];
@(posedge clk);
#1;data_in = testData6[1713];
@(posedge clk);
#1;data_in = testData6[1714];
@(posedge clk);
#1;data_in = testData6[1715];
@(posedge clk);
#1;data_in = testData6[1716];
@(posedge clk);
#1;data_in = testData6[1717];
@(posedge clk);
#1;data_in = testData6[1718];
@(posedge clk);
#1;data_in = testData6[1719];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1720]; 
@(posedge clk);
#1;data_in = testData6[1721];
@(posedge clk);
#1;data_in = testData6[1722];
@(posedge clk);
#1;data_in = testData6[1723];
@(posedge clk);
#1;data_in = testData6[1724];
@(posedge clk);
#1;data_in = testData6[1725];
@(posedge clk);
#1;data_in = testData6[1726];
@(posedge clk);
#1;data_in = testData6[1727];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1728];
@(posedge clk);
#1;data_in = testData6[1729];
@(posedge clk);
#1;data_in = testData6[1730];
@(posedge clk);
#1;data_in = testData6[1731];
@(posedge clk);
#1;data_in = testData6[1732];
@(posedge clk);
#1;data_in = testData6[1733];
@(posedge clk);
#1;data_in = testData6[1734];
@(posedge clk);
#1;data_in = testData6[1735];
@(posedge clk);
#1;data_in = testData6[1736];
@(posedge clk);
#1;data_in = testData6[1737];
@(posedge clk);
#1;data_in = testData6[1738];
@(posedge clk);
#1;data_in = testData6[1739];
@(posedge clk);
#1;data_in = testData6[1740];
@(posedge clk);
#1;data_in = testData6[1741];
@(posedge clk);
#1;data_in = testData6[1742];
@(posedge clk);
#1;data_in = testData6[1743];
@(posedge clk);
#1;data_in = testData6[1744];
@(posedge clk);
#1;data_in = testData6[1745];
@(posedge clk);
#1;data_in = testData6[1746];
@(posedge clk);
#1;data_in = testData6[1747];
@(posedge clk);
#1;data_in = testData6[1748];
@(posedge clk);
#1;data_in = testData6[1749];
@(posedge clk);
#1;data_in = testData6[1750];
@(posedge clk);
#1;data_in = testData6[1751];
@(posedge clk);
#1;data_in = testData6[1752];
@(posedge clk);
#1;data_in = testData6[1753];
@(posedge clk);
#1;data_in = testData6[1754];
@(posedge clk);
#1;data_in = testData6[1755];
@(posedge clk);
#1;data_in = testData6[1756];
@(posedge clk);
#1;data_in = testData6[1757];
@(posedge clk);
#1;data_in = testData6[1758];
@(posedge clk);
#1;data_in = testData6[1759];
@(posedge clk);
#1;data_in = testData6[1760];
@(posedge clk);
#1;data_in = testData6[1761];
@(posedge clk);
#1;data_in = testData6[1762];
@(posedge clk);
#1;data_in = testData6[1763];
@(posedge clk);
#1;data_in = testData6[1764];
@(posedge clk);
#1;data_in = testData6[1765];
@(posedge clk);
#1;data_in = testData6[1766];
@(posedge clk);
#1;data_in = testData6[1767];
@(posedge clk);
#1;data_in = testData6[1768];
@(posedge clk);
#1;data_in = testData6[1769];
@(posedge clk);
#1;data_in = testData6[1770];
@(posedge clk);
#1;data_in = testData6[1771];
@(posedge clk);
#1;data_in = testData6[1772];
@(posedge clk);
#1;data_in = testData6[1773];
@(posedge clk);
#1;data_in = testData6[1774];
@(posedge clk);
#1;data_in = testData6[1775];
@(posedge clk);
#1;data_in = testData6[1776];
@(posedge clk);
#1;data_in = testData6[1777];
@(posedge clk);
#1;data_in = testData6[1778];
@(posedge clk);
#1;data_in = testData6[1779];
@(posedge clk);
#1;data_in = testData6[1780];
@(posedge clk);
#1;data_in = testData6[1781];
@(posedge clk);
#1;data_in = testData6[1782];
@(posedge clk);
#1;data_in = testData6[1783];
@(posedge clk);
#1;data_in = testData6[1784];
@(posedge clk);
#1;data_in = testData6[1785];
@(posedge clk);
#1;data_in = testData6[1786];
@(posedge clk);
#1;data_in = testData6[1787];
@(posedge clk);
#1;data_in = testData6[1788];
@(posedge clk);
#1;data_in = testData6[1789];
@(posedge clk);
#1;data_in = testData6[1790];
@(posedge clk);
#1;data_in = testData6[1791];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1792]; 
@(posedge clk);
#1;data_in = testData6[1793];
@(posedge clk);
#1;data_in = testData6[1794];
@(posedge clk);
#1;data_in = testData6[1795];
@(posedge clk);
#1;data_in = testData6[1796];
@(posedge clk);
#1;data_in = testData6[1797];
@(posedge clk);
#1;data_in = testData6[1798];
@(posedge clk);
#1;data_in = testData6[1799];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1800];
@(posedge clk);
#1;data_in = testData6[1801];
@(posedge clk);
#1;data_in = testData6[1802];
@(posedge clk);
#1;data_in = testData6[1803];
@(posedge clk);
#1;data_in = testData6[1804];
@(posedge clk);
#1;data_in = testData6[1805];
@(posedge clk);
#1;data_in = testData6[1806];
@(posedge clk);
#1;data_in = testData6[1807];
@(posedge clk);
#1;data_in = testData6[1808];
@(posedge clk);
#1;data_in = testData6[1809];
@(posedge clk);
#1;data_in = testData6[1810];
@(posedge clk);
#1;data_in = testData6[1811];
@(posedge clk);
#1;data_in = testData6[1812];
@(posedge clk);
#1;data_in = testData6[1813];
@(posedge clk);
#1;data_in = testData6[1814];
@(posedge clk);
#1;data_in = testData6[1815];
@(posedge clk);
#1;data_in = testData6[1816];
@(posedge clk);
#1;data_in = testData6[1817];
@(posedge clk);
#1;data_in = testData6[1818];
@(posedge clk);
#1;data_in = testData6[1819];
@(posedge clk);
#1;data_in = testData6[1820];
@(posedge clk);
#1;data_in = testData6[1821];
@(posedge clk);
#1;data_in = testData6[1822];
@(posedge clk);
#1;data_in = testData6[1823];
@(posedge clk);
#1;data_in = testData6[1824];
@(posedge clk);
#1;data_in = testData6[1825];
@(posedge clk);
#1;data_in = testData6[1826];
@(posedge clk);
#1;data_in = testData6[1827];
@(posedge clk);
#1;data_in = testData6[1828];
@(posedge clk);
#1;data_in = testData6[1829];
@(posedge clk);
#1;data_in = testData6[1830];
@(posedge clk);
#1;data_in = testData6[1831];
@(posedge clk);
#1;data_in = testData6[1832];
@(posedge clk);
#1;data_in = testData6[1833];
@(posedge clk);
#1;data_in = testData6[1834];
@(posedge clk);
#1;data_in = testData6[1835];
@(posedge clk);
#1;data_in = testData6[1836];
@(posedge clk);
#1;data_in = testData6[1837];
@(posedge clk);
#1;data_in = testData6[1838];
@(posedge clk);
#1;data_in = testData6[1839];
@(posedge clk);
#1;data_in = testData6[1840];
@(posedge clk);
#1;data_in = testData6[1841];
@(posedge clk);
#1;data_in = testData6[1842];
@(posedge clk);
#1;data_in = testData6[1843];
@(posedge clk);
#1;data_in = testData6[1844];
@(posedge clk);
#1;data_in = testData6[1845];
@(posedge clk);
#1;data_in = testData6[1846];
@(posedge clk);
#1;data_in = testData6[1847];
@(posedge clk);
#1;data_in = testData6[1848];
@(posedge clk);
#1;data_in = testData6[1849];
@(posedge clk);
#1;data_in = testData6[1850];
@(posedge clk);
#1;data_in = testData6[1851];
@(posedge clk);
#1;data_in = testData6[1852];
@(posedge clk);
#1;data_in = testData6[1853];
@(posedge clk);
#1;data_in = testData6[1854];
@(posedge clk);
#1;data_in = testData6[1855];
@(posedge clk);
#1;data_in = testData6[1856];
@(posedge clk);
#1;data_in = testData6[1857];
@(posedge clk);
#1;data_in = testData6[1858];
@(posedge clk);
#1;data_in = testData6[1859];
@(posedge clk);
#1;data_in = testData6[1860];
@(posedge clk);
#1;data_in = testData6[1861];
@(posedge clk);
#1;data_in = testData6[1862];
@(posedge clk);
#1;data_in = testData6[1863];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1864]; 
@(posedge clk);
#1;data_in = testData6[1865];
@(posedge clk);
#1;data_in = testData6[1866];
@(posedge clk);
#1;data_in = testData6[1867];
@(posedge clk);
#1;data_in = testData6[1868];
@(posedge clk);
#1;data_in = testData6[1869];
@(posedge clk);
#1;data_in = testData6[1870];
@(posedge clk);
#1;data_in = testData6[1871];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1872];
@(posedge clk);
#1;data_in = testData6[1873];
@(posedge clk);
#1;data_in = testData6[1874];
@(posedge clk);
#1;data_in = testData6[1875];
@(posedge clk);
#1;data_in = testData6[1876];
@(posedge clk);
#1;data_in = testData6[1877];
@(posedge clk);
#1;data_in = testData6[1878];
@(posedge clk);
#1;data_in = testData6[1879];
@(posedge clk);
#1;data_in = testData6[1880];
@(posedge clk);
#1;data_in = testData6[1881];
@(posedge clk);
#1;data_in = testData6[1882];
@(posedge clk);
#1;data_in = testData6[1883];
@(posedge clk);
#1;data_in = testData6[1884];
@(posedge clk);
#1;data_in = testData6[1885];
@(posedge clk);
#1;data_in = testData6[1886];
@(posedge clk);
#1;data_in = testData6[1887];
@(posedge clk);
#1;data_in = testData6[1888];
@(posedge clk);
#1;data_in = testData6[1889];
@(posedge clk);
#1;data_in = testData6[1890];
@(posedge clk);
#1;data_in = testData6[1891];
@(posedge clk);
#1;data_in = testData6[1892];
@(posedge clk);
#1;data_in = testData6[1893];
@(posedge clk);
#1;data_in = testData6[1894];
@(posedge clk);
#1;data_in = testData6[1895];
@(posedge clk);
#1;data_in = testData6[1896];
@(posedge clk);
#1;data_in = testData6[1897];
@(posedge clk);
#1;data_in = testData6[1898];
@(posedge clk);
#1;data_in = testData6[1899];
@(posedge clk);
#1;data_in = testData6[1900];
@(posedge clk);
#1;data_in = testData6[1901];
@(posedge clk);
#1;data_in = testData6[1902];
@(posedge clk);
#1;data_in = testData6[1903];
@(posedge clk);
#1;data_in = testData6[1904];
@(posedge clk);
#1;data_in = testData6[1905];
@(posedge clk);
#1;data_in = testData6[1906];
@(posedge clk);
#1;data_in = testData6[1907];
@(posedge clk);
#1;data_in = testData6[1908];
@(posedge clk);
#1;data_in = testData6[1909];
@(posedge clk);
#1;data_in = testData6[1910];
@(posedge clk);
#1;data_in = testData6[1911];
@(posedge clk);
#1;data_in = testData6[1912];
@(posedge clk);
#1;data_in = testData6[1913];
@(posedge clk);
#1;data_in = testData6[1914];
@(posedge clk);
#1;data_in = testData6[1915];
@(posedge clk);
#1;data_in = testData6[1916];
@(posedge clk);
#1;data_in = testData6[1917];
@(posedge clk);
#1;data_in = testData6[1918];
@(posedge clk);
#1;data_in = testData6[1919];
@(posedge clk);
#1;data_in = testData6[1920];
@(posedge clk);
#1;data_in = testData6[1921];
@(posedge clk);
#1;data_in = testData6[1922];
@(posedge clk);
#1;data_in = testData6[1923];
@(posedge clk);
#1;data_in = testData6[1924];
@(posedge clk);
#1;data_in = testData6[1925];
@(posedge clk);
#1;data_in = testData6[1926];
@(posedge clk);
#1;data_in = testData6[1927];
@(posedge clk);
#1;data_in = testData6[1928];
@(posedge clk);
#1;data_in = testData6[1929];
@(posedge clk);
#1;data_in = testData6[1930];
@(posedge clk);
#1;data_in = testData6[1931];
@(posedge clk);
#1;data_in = testData6[1932];
@(posedge clk);
#1;data_in = testData6[1933];
@(posedge clk);
#1;data_in = testData6[1934];
@(posedge clk);
#1;data_in = testData6[1935];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1936]; 
@(posedge clk);
#1;data_in = testData6[1937];
@(posedge clk);
#1;data_in = testData6[1938];
@(posedge clk);
#1;data_in = testData6[1939];
@(posedge clk);
#1;data_in = testData6[1940];
@(posedge clk);
#1;data_in = testData6[1941];
@(posedge clk);
#1;data_in = testData6[1942];
@(posedge clk);
#1;data_in = testData6[1943];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1944];
@(posedge clk);
#1;data_in = testData6[1945];
@(posedge clk);
#1;data_in = testData6[1946];
@(posedge clk);
#1;data_in = testData6[1947];
@(posedge clk);
#1;data_in = testData6[1948];
@(posedge clk);
#1;data_in = testData6[1949];
@(posedge clk);
#1;data_in = testData6[1950];
@(posedge clk);
#1;data_in = testData6[1951];
@(posedge clk);
#1;data_in = testData6[1952];
@(posedge clk);
#1;data_in = testData6[1953];
@(posedge clk);
#1;data_in = testData6[1954];
@(posedge clk);
#1;data_in = testData6[1955];
@(posedge clk);
#1;data_in = testData6[1956];
@(posedge clk);
#1;data_in = testData6[1957];
@(posedge clk);
#1;data_in = testData6[1958];
@(posedge clk);
#1;data_in = testData6[1959];
@(posedge clk);
#1;data_in = testData6[1960];
@(posedge clk);
#1;data_in = testData6[1961];
@(posedge clk);
#1;data_in = testData6[1962];
@(posedge clk);
#1;data_in = testData6[1963];
@(posedge clk);
#1;data_in = testData6[1964];
@(posedge clk);
#1;data_in = testData6[1965];
@(posedge clk);
#1;data_in = testData6[1966];
@(posedge clk);
#1;data_in = testData6[1967];
@(posedge clk);
#1;data_in = testData6[1968];
@(posedge clk);
#1;data_in = testData6[1969];
@(posedge clk);
#1;data_in = testData6[1970];
@(posedge clk);
#1;data_in = testData6[1971];
@(posedge clk);
#1;data_in = testData6[1972];
@(posedge clk);
#1;data_in = testData6[1973];
@(posedge clk);
#1;data_in = testData6[1974];
@(posedge clk);
#1;data_in = testData6[1975];
@(posedge clk);
#1;data_in = testData6[1976];
@(posedge clk);
#1;data_in = testData6[1977];
@(posedge clk);
#1;data_in = testData6[1978];
@(posedge clk);
#1;data_in = testData6[1979];
@(posedge clk);
#1;data_in = testData6[1980];
@(posedge clk);
#1;data_in = testData6[1981];
@(posedge clk);
#1;data_in = testData6[1982];
@(posedge clk);
#1;data_in = testData6[1983];
@(posedge clk);
#1;data_in = testData6[1984];
@(posedge clk);
#1;data_in = testData6[1985];
@(posedge clk);
#1;data_in = testData6[1986];
@(posedge clk);
#1;data_in = testData6[1987];
@(posedge clk);
#1;data_in = testData6[1988];
@(posedge clk);
#1;data_in = testData6[1989];
@(posedge clk);
#1;data_in = testData6[1990];
@(posedge clk);
#1;data_in = testData6[1991];
@(posedge clk);
#1;data_in = testData6[1992];
@(posedge clk);
#1;data_in = testData6[1993];
@(posedge clk);
#1;data_in = testData6[1994];
@(posedge clk);
#1;data_in = testData6[1995];
@(posedge clk);
#1;data_in = testData6[1996];
@(posedge clk);
#1;data_in = testData6[1997];
@(posedge clk);
#1;data_in = testData6[1998];
@(posedge clk);
#1;data_in = testData6[1999];
@(posedge clk);
#1;data_in = testData6[2000];
@(posedge clk);
#1;data_in = testData6[2001];
@(posedge clk);
#1;data_in = testData6[2002];
@(posedge clk);
#1;data_in = testData6[2003];
@(posedge clk);
#1;data_in = testData6[2004];
@(posedge clk);
#1;data_in = testData6[2005];
@(posedge clk);
#1;data_in = testData6[2006];
@(posedge clk);
#1;data_in = testData6[2007];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2008]; 
@(posedge clk);
#1;data_in = testData6[2009];
@(posedge clk);
#1;data_in = testData6[2010];
@(posedge clk);
#1;data_in = testData6[2011];
@(posedge clk);
#1;data_in = testData6[2012];
@(posedge clk);
#1;data_in = testData6[2013];
@(posedge clk);
#1;data_in = testData6[2014];
@(posedge clk);
#1;data_in = testData6[2015];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2016];
@(posedge clk);
#1;data_in = testData6[2017];
@(posedge clk);
#1;data_in = testData6[2018];
@(posedge clk);
#1;data_in = testData6[2019];
@(posedge clk);
#1;data_in = testData6[2020];
@(posedge clk);
#1;data_in = testData6[2021];
@(posedge clk);
#1;data_in = testData6[2022];
@(posedge clk);
#1;data_in = testData6[2023];
@(posedge clk);
#1;data_in = testData6[2024];
@(posedge clk);
#1;data_in = testData6[2025];
@(posedge clk);
#1;data_in = testData6[2026];
@(posedge clk);
#1;data_in = testData6[2027];
@(posedge clk);
#1;data_in = testData6[2028];
@(posedge clk);
#1;data_in = testData6[2029];
@(posedge clk);
#1;data_in = testData6[2030];
@(posedge clk);
#1;data_in = testData6[2031];
@(posedge clk);
#1;data_in = testData6[2032];
@(posedge clk);
#1;data_in = testData6[2033];
@(posedge clk);
#1;data_in = testData6[2034];
@(posedge clk);
#1;data_in = testData6[2035];
@(posedge clk);
#1;data_in = testData6[2036];
@(posedge clk);
#1;data_in = testData6[2037];
@(posedge clk);
#1;data_in = testData6[2038];
@(posedge clk);
#1;data_in = testData6[2039];
@(posedge clk);
#1;data_in = testData6[2040];
@(posedge clk);
#1;data_in = testData6[2041];
@(posedge clk);
#1;data_in = testData6[2042];
@(posedge clk);
#1;data_in = testData6[2043];
@(posedge clk);
#1;data_in = testData6[2044];
@(posedge clk);
#1;data_in = testData6[2045];
@(posedge clk);
#1;data_in = testData6[2046];
@(posedge clk);
#1;data_in = testData6[2047];
@(posedge clk);
#1;data_in = testData6[2048];
@(posedge clk);
#1;data_in = testData6[2049];
@(posedge clk);
#1;data_in = testData6[2050];
@(posedge clk);
#1;data_in = testData6[2051];
@(posedge clk);
#1;data_in = testData6[2052];
@(posedge clk);
#1;data_in = testData6[2053];
@(posedge clk);
#1;data_in = testData6[2054];
@(posedge clk);
#1;data_in = testData6[2055];
@(posedge clk);
#1;data_in = testData6[2056];
@(posedge clk);
#1;data_in = testData6[2057];
@(posedge clk);
#1;data_in = testData6[2058];
@(posedge clk);
#1;data_in = testData6[2059];
@(posedge clk);
#1;data_in = testData6[2060];
@(posedge clk);
#1;data_in = testData6[2061];
@(posedge clk);
#1;data_in = testData6[2062];
@(posedge clk);
#1;data_in = testData6[2063];
@(posedge clk);
#1;data_in = testData6[2064];
@(posedge clk);
#1;data_in = testData6[2065];
@(posedge clk);
#1;data_in = testData6[2066];
@(posedge clk);
#1;data_in = testData6[2067];
@(posedge clk);
#1;data_in = testData6[2068];
@(posedge clk);
#1;data_in = testData6[2069];
@(posedge clk);
#1;data_in = testData6[2070];
@(posedge clk);
#1;data_in = testData6[2071];
@(posedge clk);
#1;data_in = testData6[2072];
@(posedge clk);
#1;data_in = testData6[2073];
@(posedge clk);
#1;data_in = testData6[2074];
@(posedge clk);
#1;data_in = testData6[2075];
@(posedge clk);
#1;data_in = testData6[2076];
@(posedge clk);
#1;data_in = testData6[2077];
@(posedge clk);
#1;data_in = testData6[2078];
@(posedge clk);
#1;data_in = testData6[2079];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2080]; 
@(posedge clk);
#1;data_in = testData6[2081];
@(posedge clk);
#1;data_in = testData6[2082];
@(posedge clk);
#1;data_in = testData6[2083];
@(posedge clk);
#1;data_in = testData6[2084];
@(posedge clk);
#1;data_in = testData6[2085];
@(posedge clk);
#1;data_in = testData6[2086];
@(posedge clk);
#1;data_in = testData6[2087];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2088];
@(posedge clk);
#1;data_in = testData6[2089];
@(posedge clk);
#1;data_in = testData6[2090];
@(posedge clk);
#1;data_in = testData6[2091];
@(posedge clk);
#1;data_in = testData6[2092];
@(posedge clk);
#1;data_in = testData6[2093];
@(posedge clk);
#1;data_in = testData6[2094];
@(posedge clk);
#1;data_in = testData6[2095];
@(posedge clk);
#1;data_in = testData6[2096];
@(posedge clk);
#1;data_in = testData6[2097];
@(posedge clk);
#1;data_in = testData6[2098];
@(posedge clk);
#1;data_in = testData6[2099];
@(posedge clk);
#1;data_in = testData6[2100];
@(posedge clk);
#1;data_in = testData6[2101];
@(posedge clk);
#1;data_in = testData6[2102];
@(posedge clk);
#1;data_in = testData6[2103];
@(posedge clk);
#1;data_in = testData6[2104];
@(posedge clk);
#1;data_in = testData6[2105];
@(posedge clk);
#1;data_in = testData6[2106];
@(posedge clk);
#1;data_in = testData6[2107];
@(posedge clk);
#1;data_in = testData6[2108];
@(posedge clk);
#1;data_in = testData6[2109];
@(posedge clk);
#1;data_in = testData6[2110];
@(posedge clk);
#1;data_in = testData6[2111];
@(posedge clk);
#1;data_in = testData6[2112];
@(posedge clk);
#1;data_in = testData6[2113];
@(posedge clk);
#1;data_in = testData6[2114];
@(posedge clk);
#1;data_in = testData6[2115];
@(posedge clk);
#1;data_in = testData6[2116];
@(posedge clk);
#1;data_in = testData6[2117];
@(posedge clk);
#1;data_in = testData6[2118];
@(posedge clk);
#1;data_in = testData6[2119];
@(posedge clk);
#1;data_in = testData6[2120];
@(posedge clk);
#1;data_in = testData6[2121];
@(posedge clk);
#1;data_in = testData6[2122];
@(posedge clk);
#1;data_in = testData6[2123];
@(posedge clk);
#1;data_in = testData6[2124];
@(posedge clk);
#1;data_in = testData6[2125];
@(posedge clk);
#1;data_in = testData6[2126];
@(posedge clk);
#1;data_in = testData6[2127];
@(posedge clk);
#1;data_in = testData6[2128];
@(posedge clk);
#1;data_in = testData6[2129];
@(posedge clk);
#1;data_in = testData6[2130];
@(posedge clk);
#1;data_in = testData6[2131];
@(posedge clk);
#1;data_in = testData6[2132];
@(posedge clk);
#1;data_in = testData6[2133];
@(posedge clk);
#1;data_in = testData6[2134];
@(posedge clk);
#1;data_in = testData6[2135];
@(posedge clk);
#1;data_in = testData6[2136];
@(posedge clk);
#1;data_in = testData6[2137];
@(posedge clk);
#1;data_in = testData6[2138];
@(posedge clk);
#1;data_in = testData6[2139];
@(posedge clk);
#1;data_in = testData6[2140];
@(posedge clk);
#1;data_in = testData6[2141];
@(posedge clk);
#1;data_in = testData6[2142];
@(posedge clk);
#1;data_in = testData6[2143];
@(posedge clk);
#1;data_in = testData6[2144];
@(posedge clk);
#1;data_in = testData6[2145];
@(posedge clk);
#1;data_in = testData6[2146];
@(posedge clk);
#1;data_in = testData6[2147];
@(posedge clk);
#1;data_in = testData6[2148];
@(posedge clk);
#1;data_in = testData6[2149];
@(posedge clk);
#1;data_in = testData6[2150];
@(posedge clk);
#1;data_in = testData6[2151];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2152]; 
@(posedge clk);
#1;data_in = testData6[2153];
@(posedge clk);
#1;data_in = testData6[2154];
@(posedge clk);
#1;data_in = testData6[2155];
@(posedge clk);
#1;data_in = testData6[2156];
@(posedge clk);
#1;data_in = testData6[2157];
@(posedge clk);
#1;data_in = testData6[2158];
@(posedge clk);
#1;data_in = testData6[2159];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2160];
@(posedge clk);
#1;data_in = testData6[2161];
@(posedge clk);
#1;data_in = testData6[2162];
@(posedge clk);
#1;data_in = testData6[2163];
@(posedge clk);
#1;data_in = testData6[2164];
@(posedge clk);
#1;data_in = testData6[2165];
@(posedge clk);
#1;data_in = testData6[2166];
@(posedge clk);
#1;data_in = testData6[2167];
@(posedge clk);
#1;data_in = testData6[2168];
@(posedge clk);
#1;data_in = testData6[2169];
@(posedge clk);
#1;data_in = testData6[2170];
@(posedge clk);
#1;data_in = testData6[2171];
@(posedge clk);
#1;data_in = testData6[2172];
@(posedge clk);
#1;data_in = testData6[2173];
@(posedge clk);
#1;data_in = testData6[2174];
@(posedge clk);
#1;data_in = testData6[2175];
@(posedge clk);
#1;data_in = testData6[2176];
@(posedge clk);
#1;data_in = testData6[2177];
@(posedge clk);
#1;data_in = testData6[2178];
@(posedge clk);
#1;data_in = testData6[2179];
@(posedge clk);
#1;data_in = testData6[2180];
@(posedge clk);
#1;data_in = testData6[2181];
@(posedge clk);
#1;data_in = testData6[2182];
@(posedge clk);
#1;data_in = testData6[2183];
@(posedge clk);
#1;data_in = testData6[2184];
@(posedge clk);
#1;data_in = testData6[2185];
@(posedge clk);
#1;data_in = testData6[2186];
@(posedge clk);
#1;data_in = testData6[2187];
@(posedge clk);
#1;data_in = testData6[2188];
@(posedge clk);
#1;data_in = testData6[2189];
@(posedge clk);
#1;data_in = testData6[2190];
@(posedge clk);
#1;data_in = testData6[2191];
@(posedge clk);
#1;data_in = testData6[2192];
@(posedge clk);
#1;data_in = testData6[2193];
@(posedge clk);
#1;data_in = testData6[2194];
@(posedge clk);
#1;data_in = testData6[2195];
@(posedge clk);
#1;data_in = testData6[2196];
@(posedge clk);
#1;data_in = testData6[2197];
@(posedge clk);
#1;data_in = testData6[2198];
@(posedge clk);
#1;data_in = testData6[2199];
@(posedge clk);
#1;data_in = testData6[2200];
@(posedge clk);
#1;data_in = testData6[2201];
@(posedge clk);
#1;data_in = testData6[2202];
@(posedge clk);
#1;data_in = testData6[2203];
@(posedge clk);
#1;data_in = testData6[2204];
@(posedge clk);
#1;data_in = testData6[2205];
@(posedge clk);
#1;data_in = testData6[2206];
@(posedge clk);
#1;data_in = testData6[2207];
@(posedge clk);
#1;data_in = testData6[2208];
@(posedge clk);
#1;data_in = testData6[2209];
@(posedge clk);
#1;data_in = testData6[2210];
@(posedge clk);
#1;data_in = testData6[2211];
@(posedge clk);
#1;data_in = testData6[2212];
@(posedge clk);
#1;data_in = testData6[2213];
@(posedge clk);
#1;data_in = testData6[2214];
@(posedge clk);
#1;data_in = testData6[2215];
@(posedge clk);
#1;data_in = testData6[2216];
@(posedge clk);
#1;data_in = testData6[2217];
@(posedge clk);
#1;data_in = testData6[2218];
@(posedge clk);
#1;data_in = testData6[2219];
@(posedge clk);
#1;data_in = testData6[2220];
@(posedge clk);
#1;data_in = testData6[2221];
@(posedge clk);
#1;data_in = testData6[2222];
@(posedge clk);
#1;data_in = testData6[2223];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2224]; 
@(posedge clk);
#1;data_in = testData6[2225];
@(posedge clk);
#1;data_in = testData6[2226];
@(posedge clk);
#1;data_in = testData6[2227];
@(posedge clk);
#1;data_in = testData6[2228];
@(posedge clk);
#1;data_in = testData6[2229];
@(posedge clk);
#1;data_in = testData6[2230];
@(posedge clk);
#1;data_in = testData6[2231];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2232];
@(posedge clk);
#1;data_in = testData6[2233];
@(posedge clk);
#1;data_in = testData6[2234];
@(posedge clk);
#1;data_in = testData6[2235];
@(posedge clk);
#1;data_in = testData6[2236];
@(posedge clk);
#1;data_in = testData6[2237];
@(posedge clk);
#1;data_in = testData6[2238];
@(posedge clk);
#1;data_in = testData6[2239];
@(posedge clk);
#1;data_in = testData6[2240];
@(posedge clk);
#1;data_in = testData6[2241];
@(posedge clk);
#1;data_in = testData6[2242];
@(posedge clk);
#1;data_in = testData6[2243];
@(posedge clk);
#1;data_in = testData6[2244];
@(posedge clk);
#1;data_in = testData6[2245];
@(posedge clk);
#1;data_in = testData6[2246];
@(posedge clk);
#1;data_in = testData6[2247];
@(posedge clk);
#1;data_in = testData6[2248];
@(posedge clk);
#1;data_in = testData6[2249];
@(posedge clk);
#1;data_in = testData6[2250];
@(posedge clk);
#1;data_in = testData6[2251];
@(posedge clk);
#1;data_in = testData6[2252];
@(posedge clk);
#1;data_in = testData6[2253];
@(posedge clk);
#1;data_in = testData6[2254];
@(posedge clk);
#1;data_in = testData6[2255];
@(posedge clk);
#1;data_in = testData6[2256];
@(posedge clk);
#1;data_in = testData6[2257];
@(posedge clk);
#1;data_in = testData6[2258];
@(posedge clk);
#1;data_in = testData6[2259];
@(posedge clk);
#1;data_in = testData6[2260];
@(posedge clk);
#1;data_in = testData6[2261];
@(posedge clk);
#1;data_in = testData6[2262];
@(posedge clk);
#1;data_in = testData6[2263];
@(posedge clk);
#1;data_in = testData6[2264];
@(posedge clk);
#1;data_in = testData6[2265];
@(posedge clk);
#1;data_in = testData6[2266];
@(posedge clk);
#1;data_in = testData6[2267];
@(posedge clk);
#1;data_in = testData6[2268];
@(posedge clk);
#1;data_in = testData6[2269];
@(posedge clk);
#1;data_in = testData6[2270];
@(posedge clk);
#1;data_in = testData6[2271];
@(posedge clk);
#1;data_in = testData6[2272];
@(posedge clk);
#1;data_in = testData6[2273];
@(posedge clk);
#1;data_in = testData6[2274];
@(posedge clk);
#1;data_in = testData6[2275];
@(posedge clk);
#1;data_in = testData6[2276];
@(posedge clk);
#1;data_in = testData6[2277];
@(posedge clk);
#1;data_in = testData6[2278];
@(posedge clk);
#1;data_in = testData6[2279];
@(posedge clk);
#1;data_in = testData6[2280];
@(posedge clk);
#1;data_in = testData6[2281];
@(posedge clk);
#1;data_in = testData6[2282];
@(posedge clk);
#1;data_in = testData6[2283];
@(posedge clk);
#1;data_in = testData6[2284];
@(posedge clk);
#1;data_in = testData6[2285];
@(posedge clk);
#1;data_in = testData6[2286];
@(posedge clk);
#1;data_in = testData6[2287];
@(posedge clk);
#1;data_in = testData6[2288];
@(posedge clk);
#1;data_in = testData6[2289];
@(posedge clk);
#1;data_in = testData6[2290];
@(posedge clk);
#1;data_in = testData6[2291];
@(posedge clk);
#1;data_in = testData6[2292];
@(posedge clk);
#1;data_in = testData6[2293];
@(posedge clk);
#1;data_in = testData6[2294];
@(posedge clk);
#1;data_in = testData6[2295];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2296]; 
@(posedge clk);
#1;data_in = testData6[2297];
@(posedge clk);
#1;data_in = testData6[2298];
@(posedge clk);
#1;data_in = testData6[2299];
@(posedge clk);
#1;data_in = testData6[2300];
@(posedge clk);
#1;data_in = testData6[2301];
@(posedge clk);
#1;data_in = testData6[2302];
@(posedge clk);
#1;data_in = testData6[2303];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2304];
@(posedge clk);
#1;data_in = testData6[2305];
@(posedge clk);
#1;data_in = testData6[2306];
@(posedge clk);
#1;data_in = testData6[2307];
@(posedge clk);
#1;data_in = testData6[2308];
@(posedge clk);
#1;data_in = testData6[2309];
@(posedge clk);
#1;data_in = testData6[2310];
@(posedge clk);
#1;data_in = testData6[2311];
@(posedge clk);
#1;data_in = testData6[2312];
@(posedge clk);
#1;data_in = testData6[2313];
@(posedge clk);
#1;data_in = testData6[2314];
@(posedge clk);
#1;data_in = testData6[2315];
@(posedge clk);
#1;data_in = testData6[2316];
@(posedge clk);
#1;data_in = testData6[2317];
@(posedge clk);
#1;data_in = testData6[2318];
@(posedge clk);
#1;data_in = testData6[2319];
@(posedge clk);
#1;data_in = testData6[2320];
@(posedge clk);
#1;data_in = testData6[2321];
@(posedge clk);
#1;data_in = testData6[2322];
@(posedge clk);
#1;data_in = testData6[2323];
@(posedge clk);
#1;data_in = testData6[2324];
@(posedge clk);
#1;data_in = testData6[2325];
@(posedge clk);
#1;data_in = testData6[2326];
@(posedge clk);
#1;data_in = testData6[2327];
@(posedge clk);
#1;data_in = testData6[2328];
@(posedge clk);
#1;data_in = testData6[2329];
@(posedge clk);
#1;data_in = testData6[2330];
@(posedge clk);
#1;data_in = testData6[2331];
@(posedge clk);
#1;data_in = testData6[2332];
@(posedge clk);
#1;data_in = testData6[2333];
@(posedge clk);
#1;data_in = testData6[2334];
@(posedge clk);
#1;data_in = testData6[2335];
@(posedge clk);
#1;data_in = testData6[2336];
@(posedge clk);
#1;data_in = testData6[2337];
@(posedge clk);
#1;data_in = testData6[2338];
@(posedge clk);
#1;data_in = testData6[2339];
@(posedge clk);
#1;data_in = testData6[2340];
@(posedge clk);
#1;data_in = testData6[2341];
@(posedge clk);
#1;data_in = testData6[2342];
@(posedge clk);
#1;data_in = testData6[2343];
@(posedge clk);
#1;data_in = testData6[2344];
@(posedge clk);
#1;data_in = testData6[2345];
@(posedge clk);
#1;data_in = testData6[2346];
@(posedge clk);
#1;data_in = testData6[2347];
@(posedge clk);
#1;data_in = testData6[2348];
@(posedge clk);
#1;data_in = testData6[2349];
@(posedge clk);
#1;data_in = testData6[2350];
@(posedge clk);
#1;data_in = testData6[2351];
@(posedge clk);
#1;data_in = testData6[2352];
@(posedge clk);
#1;data_in = testData6[2353];
@(posedge clk);
#1;data_in = testData6[2354];
@(posedge clk);
#1;data_in = testData6[2355];
@(posedge clk);
#1;data_in = testData6[2356];
@(posedge clk);
#1;data_in = testData6[2357];
@(posedge clk);
#1;data_in = testData6[2358];
@(posedge clk);
#1;data_in = testData6[2359];
@(posedge clk);
#1;data_in = testData6[2360];
@(posedge clk);
#1;data_in = testData6[2361];
@(posedge clk);
#1;data_in = testData6[2362];
@(posedge clk);
#1;data_in = testData6[2363];
@(posedge clk);
#1;data_in = testData6[2364];
@(posedge clk);
#1;data_in = testData6[2365];
@(posedge clk);
#1;data_in = testData6[2366];
@(posedge clk);
#1;data_in = testData6[2367];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2368]; 
@(posedge clk);
#1;data_in = testData6[2369];
@(posedge clk);
#1;data_in = testData6[2370];
@(posedge clk);
#1;data_in = testData6[2371];
@(posedge clk);
#1;data_in = testData6[2372];
@(posedge clk);
#1;data_in = testData6[2373];
@(posedge clk);
#1;data_in = testData6[2374];
@(posedge clk);
#1;data_in = testData6[2375];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2376];
@(posedge clk);
#1;data_in = testData6[2377];
@(posedge clk);
#1;data_in = testData6[2378];
@(posedge clk);
#1;data_in = testData6[2379];
@(posedge clk);
#1;data_in = testData6[2380];
@(posedge clk);
#1;data_in = testData6[2381];
@(posedge clk);
#1;data_in = testData6[2382];
@(posedge clk);
#1;data_in = testData6[2383];
@(posedge clk);
#1;data_in = testData6[2384];
@(posedge clk);
#1;data_in = testData6[2385];
@(posedge clk);
#1;data_in = testData6[2386];
@(posedge clk);
#1;data_in = testData6[2387];
@(posedge clk);
#1;data_in = testData6[2388];
@(posedge clk);
#1;data_in = testData6[2389];
@(posedge clk);
#1;data_in = testData6[2390];
@(posedge clk);
#1;data_in = testData6[2391];
@(posedge clk);
#1;data_in = testData6[2392];
@(posedge clk);
#1;data_in = testData6[2393];
@(posedge clk);
#1;data_in = testData6[2394];
@(posedge clk);
#1;data_in = testData6[2395];
@(posedge clk);
#1;data_in = testData6[2396];
@(posedge clk);
#1;data_in = testData6[2397];
@(posedge clk);
#1;data_in = testData6[2398];
@(posedge clk);
#1;data_in = testData6[2399];
@(posedge clk);
#1;data_in = testData6[2400];
@(posedge clk);
#1;data_in = testData6[2401];
@(posedge clk);
#1;data_in = testData6[2402];
@(posedge clk);
#1;data_in = testData6[2403];
@(posedge clk);
#1;data_in = testData6[2404];
@(posedge clk);
#1;data_in = testData6[2405];
@(posedge clk);
#1;data_in = testData6[2406];
@(posedge clk);
#1;data_in = testData6[2407];
@(posedge clk);
#1;data_in = testData6[2408];
@(posedge clk);
#1;data_in = testData6[2409];
@(posedge clk);
#1;data_in = testData6[2410];
@(posedge clk);
#1;data_in = testData6[2411];
@(posedge clk);
#1;data_in = testData6[2412];
@(posedge clk);
#1;data_in = testData6[2413];
@(posedge clk);
#1;data_in = testData6[2414];
@(posedge clk);
#1;data_in = testData6[2415];
@(posedge clk);
#1;data_in = testData6[2416];
@(posedge clk);
#1;data_in = testData6[2417];
@(posedge clk);
#1;data_in = testData6[2418];
@(posedge clk);
#1;data_in = testData6[2419];
@(posedge clk);
#1;data_in = testData6[2420];
@(posedge clk);
#1;data_in = testData6[2421];
@(posedge clk);
#1;data_in = testData6[2422];
@(posedge clk);
#1;data_in = testData6[2423];
@(posedge clk);
#1;data_in = testData6[2424];
@(posedge clk);
#1;data_in = testData6[2425];
@(posedge clk);
#1;data_in = testData6[2426];
@(posedge clk);
#1;data_in = testData6[2427];
@(posedge clk);
#1;data_in = testData6[2428];
@(posedge clk);
#1;data_in = testData6[2429];
@(posedge clk);
#1;data_in = testData6[2430];
@(posedge clk);
#1;data_in = testData6[2431];
@(posedge clk);
#1;data_in = testData6[2432];
@(posedge clk);
#1;data_in = testData6[2433];
@(posedge clk);
#1;data_in = testData6[2434];
@(posedge clk);
#1;data_in = testData6[2435];
@(posedge clk);
#1;data_in = testData6[2436];
@(posedge clk);
#1;data_in = testData6[2437];
@(posedge clk);
#1;data_in = testData6[2438];
@(posedge clk);
#1;data_in = testData6[2439];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2440]; 
@(posedge clk);
#1;data_in = testData6[2441];
@(posedge clk);
#1;data_in = testData6[2442];
@(posedge clk);
#1;data_in = testData6[2443];
@(posedge clk);
#1;data_in = testData6[2444];
@(posedge clk);
#1;data_in = testData6[2445];
@(posedge clk);
#1;data_in = testData6[2446];
@(posedge clk);
#1;data_in = testData6[2447];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2448];
@(posedge clk);
#1;data_in = testData6[2449];
@(posedge clk);
#1;data_in = testData6[2450];
@(posedge clk);
#1;data_in = testData6[2451];
@(posedge clk);
#1;data_in = testData6[2452];
@(posedge clk);
#1;data_in = testData6[2453];
@(posedge clk);
#1;data_in = testData6[2454];
@(posedge clk);
#1;data_in = testData6[2455];
@(posedge clk);
#1;data_in = testData6[2456];
@(posedge clk);
#1;data_in = testData6[2457];
@(posedge clk);
#1;data_in = testData6[2458];
@(posedge clk);
#1;data_in = testData6[2459];
@(posedge clk);
#1;data_in = testData6[2460];
@(posedge clk);
#1;data_in = testData6[2461];
@(posedge clk);
#1;data_in = testData6[2462];
@(posedge clk);
#1;data_in = testData6[2463];
@(posedge clk);
#1;data_in = testData6[2464];
@(posedge clk);
#1;data_in = testData6[2465];
@(posedge clk);
#1;data_in = testData6[2466];
@(posedge clk);
#1;data_in = testData6[2467];
@(posedge clk);
#1;data_in = testData6[2468];
@(posedge clk);
#1;data_in = testData6[2469];
@(posedge clk);
#1;data_in = testData6[2470];
@(posedge clk);
#1;data_in = testData6[2471];
@(posedge clk);
#1;data_in = testData6[2472];
@(posedge clk);
#1;data_in = testData6[2473];
@(posedge clk);
#1;data_in = testData6[2474];
@(posedge clk);
#1;data_in = testData6[2475];
@(posedge clk);
#1;data_in = testData6[2476];
@(posedge clk);
#1;data_in = testData6[2477];
@(posedge clk);
#1;data_in = testData6[2478];
@(posedge clk);
#1;data_in = testData6[2479];
@(posedge clk);
#1;data_in = testData6[2480];
@(posedge clk);
#1;data_in = testData6[2481];
@(posedge clk);
#1;data_in = testData6[2482];
@(posedge clk);
#1;data_in = testData6[2483];
@(posedge clk);
#1;data_in = testData6[2484];
@(posedge clk);
#1;data_in = testData6[2485];
@(posedge clk);
#1;data_in = testData6[2486];
@(posedge clk);
#1;data_in = testData6[2487];
@(posedge clk);
#1;data_in = testData6[2488];
@(posedge clk);
#1;data_in = testData6[2489];
@(posedge clk);
#1;data_in = testData6[2490];
@(posedge clk);
#1;data_in = testData6[2491];
@(posedge clk);
#1;data_in = testData6[2492];
@(posedge clk);
#1;data_in = testData6[2493];
@(posedge clk);
#1;data_in = testData6[2494];
@(posedge clk);
#1;data_in = testData6[2495];
@(posedge clk);
#1;data_in = testData6[2496];
@(posedge clk);
#1;data_in = testData6[2497];
@(posedge clk);
#1;data_in = testData6[2498];
@(posedge clk);
#1;data_in = testData6[2499];
@(posedge clk);
#1;data_in = testData6[2500];
@(posedge clk);
#1;data_in = testData6[2501];
@(posedge clk);
#1;data_in = testData6[2502];
@(posedge clk);
#1;data_in = testData6[2503];
@(posedge clk);
#1;data_in = testData6[2504];
@(posedge clk);
#1;data_in = testData6[2505];
@(posedge clk);
#1;data_in = testData6[2506];
@(posedge clk);
#1;data_in = testData6[2507];
@(posedge clk);
#1;data_in = testData6[2508];
@(posedge clk);
#1;data_in = testData6[2509];
@(posedge clk);
#1;data_in = testData6[2510];
@(posedge clk);
#1;data_in = testData6[2511];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2512]; 
@(posedge clk);
#1;data_in = testData6[2513];
@(posedge clk);
#1;data_in = testData6[2514];
@(posedge clk);
#1;data_in = testData6[2515];
@(posedge clk);
#1;data_in = testData6[2516];
@(posedge clk);
#1;data_in = testData6[2517];
@(posedge clk);
#1;data_in = testData6[2518];
@(posedge clk);
#1;data_in = testData6[2519];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2520];
@(posedge clk);
#1;data_in = testData6[2521];
@(posedge clk);
#1;data_in = testData6[2522];
@(posedge clk);
#1;data_in = testData6[2523];
@(posedge clk);
#1;data_in = testData6[2524];
@(posedge clk);
#1;data_in = testData6[2525];
@(posedge clk);
#1;data_in = testData6[2526];
@(posedge clk);
#1;data_in = testData6[2527];
@(posedge clk);
#1;data_in = testData6[2528];
@(posedge clk);
#1;data_in = testData6[2529];
@(posedge clk);
#1;data_in = testData6[2530];
@(posedge clk);
#1;data_in = testData6[2531];
@(posedge clk);
#1;data_in = testData6[2532];
@(posedge clk);
#1;data_in = testData6[2533];
@(posedge clk);
#1;data_in = testData6[2534];
@(posedge clk);
#1;data_in = testData6[2535];
@(posedge clk);
#1;data_in = testData6[2536];
@(posedge clk);
#1;data_in = testData6[2537];
@(posedge clk);
#1;data_in = testData6[2538];
@(posedge clk);
#1;data_in = testData6[2539];
@(posedge clk);
#1;data_in = testData6[2540];
@(posedge clk);
#1;data_in = testData6[2541];
@(posedge clk);
#1;data_in = testData6[2542];
@(posedge clk);
#1;data_in = testData6[2543];
@(posedge clk);
#1;data_in = testData6[2544];
@(posedge clk);
#1;data_in = testData6[2545];
@(posedge clk);
#1;data_in = testData6[2546];
@(posedge clk);
#1;data_in = testData6[2547];
@(posedge clk);
#1;data_in = testData6[2548];
@(posedge clk);
#1;data_in = testData6[2549];
@(posedge clk);
#1;data_in = testData6[2550];
@(posedge clk);
#1;data_in = testData6[2551];
@(posedge clk);
#1;data_in = testData6[2552];
@(posedge clk);
#1;data_in = testData6[2553];
@(posedge clk);
#1;data_in = testData6[2554];
@(posedge clk);
#1;data_in = testData6[2555];
@(posedge clk);
#1;data_in = testData6[2556];
@(posedge clk);
#1;data_in = testData6[2557];
@(posedge clk);
#1;data_in = testData6[2558];
@(posedge clk);
#1;data_in = testData6[2559];
@(posedge clk);
#1;data_in = testData6[2560];
@(posedge clk);
#1;data_in = testData6[2561];
@(posedge clk);
#1;data_in = testData6[2562];
@(posedge clk);
#1;data_in = testData6[2563];
@(posedge clk);
#1;data_in = testData6[2564];
@(posedge clk);
#1;data_in = testData6[2565];
@(posedge clk);
#1;data_in = testData6[2566];
@(posedge clk);
#1;data_in = testData6[2567];
@(posedge clk);
#1;data_in = testData6[2568];
@(posedge clk);
#1;data_in = testData6[2569];
@(posedge clk);
#1;data_in = testData6[2570];
@(posedge clk);
#1;data_in = testData6[2571];
@(posedge clk);
#1;data_in = testData6[2572];
@(posedge clk);
#1;data_in = testData6[2573];
@(posedge clk);
#1;data_in = testData6[2574];
@(posedge clk);
#1;data_in = testData6[2575];
@(posedge clk);
#1;data_in = testData6[2576];
@(posedge clk);
#1;data_in = testData6[2577];
@(posedge clk);
#1;data_in = testData6[2578];
@(posedge clk);
#1;data_in = testData6[2579];
@(posedge clk);
#1;data_in = testData6[2580];
@(posedge clk);
#1;data_in = testData6[2581];
@(posedge clk);
#1;data_in = testData6[2582];
@(posedge clk);
#1;data_in = testData6[2583];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2584]; 
@(posedge clk);
#1;data_in = testData6[2585];
@(posedge clk);
#1;data_in = testData6[2586];
@(posedge clk);
#1;data_in = testData6[2587];
@(posedge clk);
#1;data_in = testData6[2588];
@(posedge clk);
#1;data_in = testData6[2589];
@(posedge clk);
#1;data_in = testData6[2590];
@(posedge clk);
#1;data_in = testData6[2591];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2592];
@(posedge clk);
#1;data_in = testData6[2593];
@(posedge clk);
#1;data_in = testData6[2594];
@(posedge clk);
#1;data_in = testData6[2595];
@(posedge clk);
#1;data_in = testData6[2596];
@(posedge clk);
#1;data_in = testData6[2597];
@(posedge clk);
#1;data_in = testData6[2598];
@(posedge clk);
#1;data_in = testData6[2599];
@(posedge clk);
#1;data_in = testData6[2600];
@(posedge clk);
#1;data_in = testData6[2601];
@(posedge clk);
#1;data_in = testData6[2602];
@(posedge clk);
#1;data_in = testData6[2603];
@(posedge clk);
#1;data_in = testData6[2604];
@(posedge clk);
#1;data_in = testData6[2605];
@(posedge clk);
#1;data_in = testData6[2606];
@(posedge clk);
#1;data_in = testData6[2607];
@(posedge clk);
#1;data_in = testData6[2608];
@(posedge clk);
#1;data_in = testData6[2609];
@(posedge clk);
#1;data_in = testData6[2610];
@(posedge clk);
#1;data_in = testData6[2611];
@(posedge clk);
#1;data_in = testData6[2612];
@(posedge clk);
#1;data_in = testData6[2613];
@(posedge clk);
#1;data_in = testData6[2614];
@(posedge clk);
#1;data_in = testData6[2615];
@(posedge clk);
#1;data_in = testData6[2616];
@(posedge clk);
#1;data_in = testData6[2617];
@(posedge clk);
#1;data_in = testData6[2618];
@(posedge clk);
#1;data_in = testData6[2619];
@(posedge clk);
#1;data_in = testData6[2620];
@(posedge clk);
#1;data_in = testData6[2621];
@(posedge clk);
#1;data_in = testData6[2622];
@(posedge clk);
#1;data_in = testData6[2623];
@(posedge clk);
#1;data_in = testData6[2624];
@(posedge clk);
#1;data_in = testData6[2625];
@(posedge clk);
#1;data_in = testData6[2626];
@(posedge clk);
#1;data_in = testData6[2627];
@(posedge clk);
#1;data_in = testData6[2628];
@(posedge clk);
#1;data_in = testData6[2629];
@(posedge clk);
#1;data_in = testData6[2630];
@(posedge clk);
#1;data_in = testData6[2631];
@(posedge clk);
#1;data_in = testData6[2632];
@(posedge clk);
#1;data_in = testData6[2633];
@(posedge clk);
#1;data_in = testData6[2634];
@(posedge clk);
#1;data_in = testData6[2635];
@(posedge clk);
#1;data_in = testData6[2636];
@(posedge clk);
#1;data_in = testData6[2637];
@(posedge clk);
#1;data_in = testData6[2638];
@(posedge clk);
#1;data_in = testData6[2639];
@(posedge clk);
#1;data_in = testData6[2640];
@(posedge clk);
#1;data_in = testData6[2641];
@(posedge clk);
#1;data_in = testData6[2642];
@(posedge clk);
#1;data_in = testData6[2643];
@(posedge clk);
#1;data_in = testData6[2644];
@(posedge clk);
#1;data_in = testData6[2645];
@(posedge clk);
#1;data_in = testData6[2646];
@(posedge clk);
#1;data_in = testData6[2647];
@(posedge clk);
#1;data_in = testData6[2648];
@(posedge clk);
#1;data_in = testData6[2649];
@(posedge clk);
#1;data_in = testData6[2650];
@(posedge clk);
#1;data_in = testData6[2651];
@(posedge clk);
#1;data_in = testData6[2652];
@(posedge clk);
#1;data_in = testData6[2653];
@(posedge clk);
#1;data_in = testData6[2654];
@(posedge clk);
#1;data_in = testData6[2655];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2656]; 
@(posedge clk);
#1;data_in = testData6[2657];
@(posedge clk);
#1;data_in = testData6[2658];
@(posedge clk);
#1;data_in = testData6[2659];
@(posedge clk);
#1;data_in = testData6[2660];
@(posedge clk);
#1;data_in = testData6[2661];
@(posedge clk);
#1;data_in = testData6[2662];
@(posedge clk);
#1;data_in = testData6[2663];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2664];
@(posedge clk);
#1;data_in = testData6[2665];
@(posedge clk);
#1;data_in = testData6[2666];
@(posedge clk);
#1;data_in = testData6[2667];
@(posedge clk);
#1;data_in = testData6[2668];
@(posedge clk);
#1;data_in = testData6[2669];
@(posedge clk);
#1;data_in = testData6[2670];
@(posedge clk);
#1;data_in = testData6[2671];
@(posedge clk);
#1;data_in = testData6[2672];
@(posedge clk);
#1;data_in = testData6[2673];
@(posedge clk);
#1;data_in = testData6[2674];
@(posedge clk);
#1;data_in = testData6[2675];
@(posedge clk);
#1;data_in = testData6[2676];
@(posedge clk);
#1;data_in = testData6[2677];
@(posedge clk);
#1;data_in = testData6[2678];
@(posedge clk);
#1;data_in = testData6[2679];
@(posedge clk);
#1;data_in = testData6[2680];
@(posedge clk);
#1;data_in = testData6[2681];
@(posedge clk);
#1;data_in = testData6[2682];
@(posedge clk);
#1;data_in = testData6[2683];
@(posedge clk);
#1;data_in = testData6[2684];
@(posedge clk);
#1;data_in = testData6[2685];
@(posedge clk);
#1;data_in = testData6[2686];
@(posedge clk);
#1;data_in = testData6[2687];
@(posedge clk);
#1;data_in = testData6[2688];
@(posedge clk);
#1;data_in = testData6[2689];
@(posedge clk);
#1;data_in = testData6[2690];
@(posedge clk);
#1;data_in = testData6[2691];
@(posedge clk);
#1;data_in = testData6[2692];
@(posedge clk);
#1;data_in = testData6[2693];
@(posedge clk);
#1;data_in = testData6[2694];
@(posedge clk);
#1;data_in = testData6[2695];
@(posedge clk);
#1;data_in = testData6[2696];
@(posedge clk);
#1;data_in = testData6[2697];
@(posedge clk);
#1;data_in = testData6[2698];
@(posedge clk);
#1;data_in = testData6[2699];
@(posedge clk);
#1;data_in = testData6[2700];
@(posedge clk);
#1;data_in = testData6[2701];
@(posedge clk);
#1;data_in = testData6[2702];
@(posedge clk);
#1;data_in = testData6[2703];
@(posedge clk);
#1;data_in = testData6[2704];
@(posedge clk);
#1;data_in = testData6[2705];
@(posedge clk);
#1;data_in = testData6[2706];
@(posedge clk);
#1;data_in = testData6[2707];
@(posedge clk);
#1;data_in = testData6[2708];
@(posedge clk);
#1;data_in = testData6[2709];
@(posedge clk);
#1;data_in = testData6[2710];
@(posedge clk);
#1;data_in = testData6[2711];
@(posedge clk);
#1;data_in = testData6[2712];
@(posedge clk);
#1;data_in = testData6[2713];
@(posedge clk);
#1;data_in = testData6[2714];
@(posedge clk);
#1;data_in = testData6[2715];
@(posedge clk);
#1;data_in = testData6[2716];
@(posedge clk);
#1;data_in = testData6[2717];
@(posedge clk);
#1;data_in = testData6[2718];
@(posedge clk);
#1;data_in = testData6[2719];
@(posedge clk);
#1;data_in = testData6[2720];
@(posedge clk);
#1;data_in = testData6[2721];
@(posedge clk);
#1;data_in = testData6[2722];
@(posedge clk);
#1;data_in = testData6[2723];
@(posedge clk);
#1;data_in = testData6[2724];
@(posedge clk);
#1;data_in = testData6[2725];
@(posedge clk);
#1;data_in = testData6[2726];
@(posedge clk);
#1;data_in = testData6[2727];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2728]; 
@(posedge clk);
#1;data_in = testData6[2729];
@(posedge clk);
#1;data_in = testData6[2730];
@(posedge clk);
#1;data_in = testData6[2731];
@(posedge clk);
#1;data_in = testData6[2732];
@(posedge clk);
#1;data_in = testData6[2733];
@(posedge clk);
#1;data_in = testData6[2734];
@(posedge clk);
#1;data_in = testData6[2735];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2736];
@(posedge clk);
#1;data_in = testData6[2737];
@(posedge clk);
#1;data_in = testData6[2738];
@(posedge clk);
#1;data_in = testData6[2739];
@(posedge clk);
#1;data_in = testData6[2740];
@(posedge clk);
#1;data_in = testData6[2741];
@(posedge clk);
#1;data_in = testData6[2742];
@(posedge clk);
#1;data_in = testData6[2743];
@(posedge clk);
#1;data_in = testData6[2744];
@(posedge clk);
#1;data_in = testData6[2745];
@(posedge clk);
#1;data_in = testData6[2746];
@(posedge clk);
#1;data_in = testData6[2747];
@(posedge clk);
#1;data_in = testData6[2748];
@(posedge clk);
#1;data_in = testData6[2749];
@(posedge clk);
#1;data_in = testData6[2750];
@(posedge clk);
#1;data_in = testData6[2751];
@(posedge clk);
#1;data_in = testData6[2752];
@(posedge clk);
#1;data_in = testData6[2753];
@(posedge clk);
#1;data_in = testData6[2754];
@(posedge clk);
#1;data_in = testData6[2755];
@(posedge clk);
#1;data_in = testData6[2756];
@(posedge clk);
#1;data_in = testData6[2757];
@(posedge clk);
#1;data_in = testData6[2758];
@(posedge clk);
#1;data_in = testData6[2759];
@(posedge clk);
#1;data_in = testData6[2760];
@(posedge clk);
#1;data_in = testData6[2761];
@(posedge clk);
#1;data_in = testData6[2762];
@(posedge clk);
#1;data_in = testData6[2763];
@(posedge clk);
#1;data_in = testData6[2764];
@(posedge clk);
#1;data_in = testData6[2765];
@(posedge clk);
#1;data_in = testData6[2766];
@(posedge clk);
#1;data_in = testData6[2767];
@(posedge clk);
#1;data_in = testData6[2768];
@(posedge clk);
#1;data_in = testData6[2769];
@(posedge clk);
#1;data_in = testData6[2770];
@(posedge clk);
#1;data_in = testData6[2771];
@(posedge clk);
#1;data_in = testData6[2772];
@(posedge clk);
#1;data_in = testData6[2773];
@(posedge clk);
#1;data_in = testData6[2774];
@(posedge clk);
#1;data_in = testData6[2775];
@(posedge clk);
#1;data_in = testData6[2776];
@(posedge clk);
#1;data_in = testData6[2777];
@(posedge clk);
#1;data_in = testData6[2778];
@(posedge clk);
#1;data_in = testData6[2779];
@(posedge clk);
#1;data_in = testData6[2780];
@(posedge clk);
#1;data_in = testData6[2781];
@(posedge clk);
#1;data_in = testData6[2782];
@(posedge clk);
#1;data_in = testData6[2783];
@(posedge clk);
#1;data_in = testData6[2784];
@(posedge clk);
#1;data_in = testData6[2785];
@(posedge clk);
#1;data_in = testData6[2786];
@(posedge clk);
#1;data_in = testData6[2787];
@(posedge clk);
#1;data_in = testData6[2788];
@(posedge clk);
#1;data_in = testData6[2789];
@(posedge clk);
#1;data_in = testData6[2790];
@(posedge clk);
#1;data_in = testData6[2791];
@(posedge clk);
#1;data_in = testData6[2792];
@(posedge clk);
#1;data_in = testData6[2793];
@(posedge clk);
#1;data_in = testData6[2794];
@(posedge clk);
#1;data_in = testData6[2795];
@(posedge clk);
#1;data_in = testData6[2796];
@(posedge clk);
#1;data_in = testData6[2797];
@(posedge clk);
#1;data_in = testData6[2798];
@(posedge clk);
#1;data_in = testData6[2799];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2800]; 
@(posedge clk);
#1;data_in = testData6[2801];
@(posedge clk);
#1;data_in = testData6[2802];
@(posedge clk);
#1;data_in = testData6[2803];
@(posedge clk);
#1;data_in = testData6[2804];
@(posedge clk);
#1;data_in = testData6[2805];
@(posedge clk);
#1;data_in = testData6[2806];
@(posedge clk);
#1;data_in = testData6[2807];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2808];
@(posedge clk);
#1;data_in = testData6[2809];
@(posedge clk);
#1;data_in = testData6[2810];
@(posedge clk);
#1;data_in = testData6[2811];
@(posedge clk);
#1;data_in = testData6[2812];
@(posedge clk);
#1;data_in = testData6[2813];
@(posedge clk);
#1;data_in = testData6[2814];
@(posedge clk);
#1;data_in = testData6[2815];
@(posedge clk);
#1;data_in = testData6[2816];
@(posedge clk);
#1;data_in = testData6[2817];
@(posedge clk);
#1;data_in = testData6[2818];
@(posedge clk);
#1;data_in = testData6[2819];
@(posedge clk);
#1;data_in = testData6[2820];
@(posedge clk);
#1;data_in = testData6[2821];
@(posedge clk);
#1;data_in = testData6[2822];
@(posedge clk);
#1;data_in = testData6[2823];
@(posedge clk);
#1;data_in = testData6[2824];
@(posedge clk);
#1;data_in = testData6[2825];
@(posedge clk);
#1;data_in = testData6[2826];
@(posedge clk);
#1;data_in = testData6[2827];
@(posedge clk);
#1;data_in = testData6[2828];
@(posedge clk);
#1;data_in = testData6[2829];
@(posedge clk);
#1;data_in = testData6[2830];
@(posedge clk);
#1;data_in = testData6[2831];
@(posedge clk);
#1;data_in = testData6[2832];
@(posedge clk);
#1;data_in = testData6[2833];
@(posedge clk);
#1;data_in = testData6[2834];
@(posedge clk);
#1;data_in = testData6[2835];
@(posedge clk);
#1;data_in = testData6[2836];
@(posedge clk);
#1;data_in = testData6[2837];
@(posedge clk);
#1;data_in = testData6[2838];
@(posedge clk);
#1;data_in = testData6[2839];
@(posedge clk);
#1;data_in = testData6[2840];
@(posedge clk);
#1;data_in = testData6[2841];
@(posedge clk);
#1;data_in = testData6[2842];
@(posedge clk);
#1;data_in = testData6[2843];
@(posedge clk);
#1;data_in = testData6[2844];
@(posedge clk);
#1;data_in = testData6[2845];
@(posedge clk);
#1;data_in = testData6[2846];
@(posedge clk);
#1;data_in = testData6[2847];
@(posedge clk);
#1;data_in = testData6[2848];
@(posedge clk);
#1;data_in = testData6[2849];
@(posedge clk);
#1;data_in = testData6[2850];
@(posedge clk);
#1;data_in = testData6[2851];
@(posedge clk);
#1;data_in = testData6[2852];
@(posedge clk);
#1;data_in = testData6[2853];
@(posedge clk);
#1;data_in = testData6[2854];
@(posedge clk);
#1;data_in = testData6[2855];
@(posedge clk);
#1;data_in = testData6[2856];
@(posedge clk);
#1;data_in = testData6[2857];
@(posedge clk);
#1;data_in = testData6[2858];
@(posedge clk);
#1;data_in = testData6[2859];
@(posedge clk);
#1;data_in = testData6[2860];
@(posedge clk);
#1;data_in = testData6[2861];
@(posedge clk);
#1;data_in = testData6[2862];
@(posedge clk);
#1;data_in = testData6[2863];
@(posedge clk);
#1;data_in = testData6[2864];
@(posedge clk);
#1;data_in = testData6[2865];
@(posedge clk);
#1;data_in = testData6[2866];
@(posedge clk);
#1;data_in = testData6[2867];
@(posedge clk);
#1;data_in = testData6[2868];
@(posedge clk);
#1;data_in = testData6[2869];
@(posedge clk);
#1;data_in = testData6[2870];
@(posedge clk);
#1;data_in = testData6[2871];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2872]; 
@(posedge clk);
#1;data_in = testData6[2873];
@(posedge clk);
#1;data_in = testData6[2874];
@(posedge clk);
#1;data_in = testData6[2875];
@(posedge clk);
#1;data_in = testData6[2876];
@(posedge clk);
#1;data_in = testData6[2877];
@(posedge clk);
#1;data_in = testData6[2878];
@(posedge clk);
#1;data_in = testData6[2879];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2880];
@(posedge clk);
#1;data_in = testData6[2881];
@(posedge clk);
#1;data_in = testData6[2882];
@(posedge clk);
#1;data_in = testData6[2883];
@(posedge clk);
#1;data_in = testData6[2884];
@(posedge clk);
#1;data_in = testData6[2885];
@(posedge clk);
#1;data_in = testData6[2886];
@(posedge clk);
#1;data_in = testData6[2887];
@(posedge clk);
#1;data_in = testData6[2888];
@(posedge clk);
#1;data_in = testData6[2889];
@(posedge clk);
#1;data_in = testData6[2890];
@(posedge clk);
#1;data_in = testData6[2891];
@(posedge clk);
#1;data_in = testData6[2892];
@(posedge clk);
#1;data_in = testData6[2893];
@(posedge clk);
#1;data_in = testData6[2894];
@(posedge clk);
#1;data_in = testData6[2895];
@(posedge clk);
#1;data_in = testData6[2896];
@(posedge clk);
#1;data_in = testData6[2897];
@(posedge clk);
#1;data_in = testData6[2898];
@(posedge clk);
#1;data_in = testData6[2899];
@(posedge clk);
#1;data_in = testData6[2900];
@(posedge clk);
#1;data_in = testData6[2901];
@(posedge clk);
#1;data_in = testData6[2902];
@(posedge clk);
#1;data_in = testData6[2903];
@(posedge clk);
#1;data_in = testData6[2904];
@(posedge clk);
#1;data_in = testData6[2905];
@(posedge clk);
#1;data_in = testData6[2906];
@(posedge clk);
#1;data_in = testData6[2907];
@(posedge clk);
#1;data_in = testData6[2908];
@(posedge clk);
#1;data_in = testData6[2909];
@(posedge clk);
#1;data_in = testData6[2910];
@(posedge clk);
#1;data_in = testData6[2911];
@(posedge clk);
#1;data_in = testData6[2912];
@(posedge clk);
#1;data_in = testData6[2913];
@(posedge clk);
#1;data_in = testData6[2914];
@(posedge clk);
#1;data_in = testData6[2915];
@(posedge clk);
#1;data_in = testData6[2916];
@(posedge clk);
#1;data_in = testData6[2917];
@(posedge clk);
#1;data_in = testData6[2918];
@(posedge clk);
#1;data_in = testData6[2919];
@(posedge clk);
#1;data_in = testData6[2920];
@(posedge clk);
#1;data_in = testData6[2921];
@(posedge clk);
#1;data_in = testData6[2922];
@(posedge clk);
#1;data_in = testData6[2923];
@(posedge clk);
#1;data_in = testData6[2924];
@(posedge clk);
#1;data_in = testData6[2925];
@(posedge clk);
#1;data_in = testData6[2926];
@(posedge clk);
#1;data_in = testData6[2927];
@(posedge clk);
#1;data_in = testData6[2928];
@(posedge clk);
#1;data_in = testData6[2929];
@(posedge clk);
#1;data_in = testData6[2930];
@(posedge clk);
#1;data_in = testData6[2931];
@(posedge clk);
#1;data_in = testData6[2932];
@(posedge clk);
#1;data_in = testData6[2933];
@(posedge clk);
#1;data_in = testData6[2934];
@(posedge clk);
#1;data_in = testData6[2935];
@(posedge clk);
#1;data_in = testData6[2936];
@(posedge clk);
#1;data_in = testData6[2937];
@(posedge clk);
#1;data_in = testData6[2938];
@(posedge clk);
#1;data_in = testData6[2939];
@(posedge clk);
#1;data_in = testData6[2940];
@(posedge clk);
#1;data_in = testData6[2941];
@(posedge clk);
#1;data_in = testData6[2942];
@(posedge clk);
#1;data_in = testData6[2943];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[2944]; 
@(posedge clk);
#1;data_in = testData6[2945];
@(posedge clk);
#1;data_in = testData6[2946];
@(posedge clk);
#1;data_in = testData6[2947];
@(posedge clk);
#1;data_in = testData6[2948];
@(posedge clk);
#1;data_in = testData6[2949];
@(posedge clk);
#1;data_in = testData6[2950];
@(posedge clk);
#1;data_in = testData6[2951];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[2952];
@(posedge clk);
#1;data_in = testData6[2953];
@(posedge clk);
#1;data_in = testData6[2954];
@(posedge clk);
#1;data_in = testData6[2955];
@(posedge clk);
#1;data_in = testData6[2956];
@(posedge clk);
#1;data_in = testData6[2957];
@(posedge clk);
#1;data_in = testData6[2958];
@(posedge clk);
#1;data_in = testData6[2959];
@(posedge clk);
#1;data_in = testData6[2960];
@(posedge clk);
#1;data_in = testData6[2961];
@(posedge clk);
#1;data_in = testData6[2962];
@(posedge clk);
#1;data_in = testData6[2963];
@(posedge clk);
#1;data_in = testData6[2964];
@(posedge clk);
#1;data_in = testData6[2965];
@(posedge clk);
#1;data_in = testData6[2966];
@(posedge clk);
#1;data_in = testData6[2967];
@(posedge clk);
#1;data_in = testData6[2968];
@(posedge clk);
#1;data_in = testData6[2969];
@(posedge clk);
#1;data_in = testData6[2970];
@(posedge clk);
#1;data_in = testData6[2971];
@(posedge clk);
#1;data_in = testData6[2972];
@(posedge clk);
#1;data_in = testData6[2973];
@(posedge clk);
#1;data_in = testData6[2974];
@(posedge clk);
#1;data_in = testData6[2975];
@(posedge clk);
#1;data_in = testData6[2976];
@(posedge clk);
#1;data_in = testData6[2977];
@(posedge clk);
#1;data_in = testData6[2978];
@(posedge clk);
#1;data_in = testData6[2979];
@(posedge clk);
#1;data_in = testData6[2980];
@(posedge clk);
#1;data_in = testData6[2981];
@(posedge clk);
#1;data_in = testData6[2982];
@(posedge clk);
#1;data_in = testData6[2983];
@(posedge clk);
#1;data_in = testData6[2984];
@(posedge clk);
#1;data_in = testData6[2985];
@(posedge clk);
#1;data_in = testData6[2986];
@(posedge clk);
#1;data_in = testData6[2987];
@(posedge clk);
#1;data_in = testData6[2988];
@(posedge clk);
#1;data_in = testData6[2989];
@(posedge clk);
#1;data_in = testData6[2990];
@(posedge clk);
#1;data_in = testData6[2991];
@(posedge clk);
#1;data_in = testData6[2992];
@(posedge clk);
#1;data_in = testData6[2993];
@(posedge clk);
#1;data_in = testData6[2994];
@(posedge clk);
#1;data_in = testData6[2995];
@(posedge clk);
#1;data_in = testData6[2996];
@(posedge clk);
#1;data_in = testData6[2997];
@(posedge clk);
#1;data_in = testData6[2998];
@(posedge clk);
#1;data_in = testData6[2999];
@(posedge clk);
#1;data_in = testData6[3000];
@(posedge clk);
#1;data_in = testData6[3001];
@(posedge clk);
#1;data_in = testData6[3002];
@(posedge clk);
#1;data_in = testData6[3003];
@(posedge clk);
#1;data_in = testData6[3004];
@(posedge clk);
#1;data_in = testData6[3005];
@(posedge clk);
#1;data_in = testData6[3006];
@(posedge clk);
#1;data_in = testData6[3007];
@(posedge clk);
#1;data_in = testData6[3008];
@(posedge clk);
#1;data_in = testData6[3009];
@(posedge clk);
#1;data_in = testData6[3010];
@(posedge clk);
#1;data_in = testData6[3011];
@(posedge clk);
#1;data_in = testData6[3012];
@(posedge clk);
#1;data_in = testData6[3013];
@(posedge clk);
#1;data_in = testData6[3014];
@(posedge clk);
#1;data_in = testData6[3015];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[3016]; 
@(posedge clk);
#1;data_in = testData6[3017];
@(posedge clk);
#1;data_in = testData6[3018];
@(posedge clk);
#1;data_in = testData6[3019];
@(posedge clk);
#1;data_in = testData6[3020];
@(posedge clk);
#1;data_in = testData6[3021];
@(posedge clk);
#1;data_in = testData6[3022];
@(posedge clk);
#1;data_in = testData6[3023];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[3024];
@(posedge clk);
#1;data_in = testData6[3025];
@(posedge clk);
#1;data_in = testData6[3026];
@(posedge clk);
#1;data_in = testData6[3027];
@(posedge clk);
#1;data_in = testData6[3028];
@(posedge clk);
#1;data_in = testData6[3029];
@(posedge clk);
#1;data_in = testData6[3030];
@(posedge clk);
#1;data_in = testData6[3031];
@(posedge clk);
#1;data_in = testData6[3032];
@(posedge clk);
#1;data_in = testData6[3033];
@(posedge clk);
#1;data_in = testData6[3034];
@(posedge clk);
#1;data_in = testData6[3035];
@(posedge clk);
#1;data_in = testData6[3036];
@(posedge clk);
#1;data_in = testData6[3037];
@(posedge clk);
#1;data_in = testData6[3038];
@(posedge clk);
#1;data_in = testData6[3039];
@(posedge clk);
#1;data_in = testData6[3040];
@(posedge clk);
#1;data_in = testData6[3041];
@(posedge clk);
#1;data_in = testData6[3042];
@(posedge clk);
#1;data_in = testData6[3043];
@(posedge clk);
#1;data_in = testData6[3044];
@(posedge clk);
#1;data_in = testData6[3045];
@(posedge clk);
#1;data_in = testData6[3046];
@(posedge clk);
#1;data_in = testData6[3047];
@(posedge clk);
#1;data_in = testData6[3048];
@(posedge clk);
#1;data_in = testData6[3049];
@(posedge clk);
#1;data_in = testData6[3050];
@(posedge clk);
#1;data_in = testData6[3051];
@(posedge clk);
#1;data_in = testData6[3052];
@(posedge clk);
#1;data_in = testData6[3053];
@(posedge clk);
#1;data_in = testData6[3054];
@(posedge clk);
#1;data_in = testData6[3055];
@(posedge clk);
#1;data_in = testData6[3056];
@(posedge clk);
#1;data_in = testData6[3057];
@(posedge clk);
#1;data_in = testData6[3058];
@(posedge clk);
#1;data_in = testData6[3059];
@(posedge clk);
#1;data_in = testData6[3060];
@(posedge clk);
#1;data_in = testData6[3061];
@(posedge clk);
#1;data_in = testData6[3062];
@(posedge clk);
#1;data_in = testData6[3063];
@(posedge clk);
#1;data_in = testData6[3064];
@(posedge clk);
#1;data_in = testData6[3065];
@(posedge clk);
#1;data_in = testData6[3066];
@(posedge clk);
#1;data_in = testData6[3067];
@(posedge clk);
#1;data_in = testData6[3068];
@(posedge clk);
#1;data_in = testData6[3069];
@(posedge clk);
#1;data_in = testData6[3070];
@(posedge clk);
#1;data_in = testData6[3071];
@(posedge clk);
#1;data_in = testData6[3072];
@(posedge clk);
#1;data_in = testData6[3073];
@(posedge clk);
#1;data_in = testData6[3074];
@(posedge clk);
#1;data_in = testData6[3075];
@(posedge clk);
#1;data_in = testData6[3076];
@(posedge clk);
#1;data_in = testData6[3077];
@(posedge clk);
#1;data_in = testData6[3078];
@(posedge clk);
#1;data_in = testData6[3079];
@(posedge clk);
#1;data_in = testData6[3080];
@(posedge clk);
#1;data_in = testData6[3081];
@(posedge clk);
#1;data_in = testData6[3082];
@(posedge clk);
#1;data_in = testData6[3083];
@(posedge clk);
#1;data_in = testData6[3084];
@(posedge clk);
#1;data_in = testData6[3085];
@(posedge clk);
#1;data_in = testData6[3086];
@(posedge clk);
#1;data_in = testData6[3087];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[3088]; 
@(posedge clk);
#1;data_in = testData6[3089];
@(posedge clk);
#1;data_in = testData6[3090];
@(posedge clk);
#1;data_in = testData6[3091];
@(posedge clk);
#1;data_in = testData6[3092];
@(posedge clk);
#1;data_in = testData6[3093];
@(posedge clk);
#1;data_in = testData6[3094];
@(posedge clk);
#1;data_in = testData6[3095];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[3096];
@(posedge clk);
#1;data_in = testData6[3097];
@(posedge clk);
#1;data_in = testData6[3098];
@(posedge clk);
#1;data_in = testData6[3099];
@(posedge clk);
#1;data_in = testData6[3100];
@(posedge clk);
#1;data_in = testData6[3101];
@(posedge clk);
#1;data_in = testData6[3102];
@(posedge clk);
#1;data_in = testData6[3103];
@(posedge clk);
#1;data_in = testData6[3104];
@(posedge clk);
#1;data_in = testData6[3105];
@(posedge clk);
#1;data_in = testData6[3106];
@(posedge clk);
#1;data_in = testData6[3107];
@(posedge clk);
#1;data_in = testData6[3108];
@(posedge clk);
#1;data_in = testData6[3109];
@(posedge clk);
#1;data_in = testData6[3110];
@(posedge clk);
#1;data_in = testData6[3111];
@(posedge clk);
#1;data_in = testData6[3112];
@(posedge clk);
#1;data_in = testData6[3113];
@(posedge clk);
#1;data_in = testData6[3114];
@(posedge clk);
#1;data_in = testData6[3115];
@(posedge clk);
#1;data_in = testData6[3116];
@(posedge clk);
#1;data_in = testData6[3117];
@(posedge clk);
#1;data_in = testData6[3118];
@(posedge clk);
#1;data_in = testData6[3119];
@(posedge clk);
#1;data_in = testData6[3120];
@(posedge clk);
#1;data_in = testData6[3121];
@(posedge clk);
#1;data_in = testData6[3122];
@(posedge clk);
#1;data_in = testData6[3123];
@(posedge clk);
#1;data_in = testData6[3124];
@(posedge clk);
#1;data_in = testData6[3125];
@(posedge clk);
#1;data_in = testData6[3126];
@(posedge clk);
#1;data_in = testData6[3127];
@(posedge clk);
#1;data_in = testData6[3128];
@(posedge clk);
#1;data_in = testData6[3129];
@(posedge clk);
#1;data_in = testData6[3130];
@(posedge clk);
#1;data_in = testData6[3131];
@(posedge clk);
#1;data_in = testData6[3132];
@(posedge clk);
#1;data_in = testData6[3133];
@(posedge clk);
#1;data_in = testData6[3134];
@(posedge clk);
#1;data_in = testData6[3135];
@(posedge clk);
#1;data_in = testData6[3136];
@(posedge clk);
#1;data_in = testData6[3137];
@(posedge clk);
#1;data_in = testData6[3138];
@(posedge clk);
#1;data_in = testData6[3139];
@(posedge clk);
#1;data_in = testData6[3140];
@(posedge clk);
#1;data_in = testData6[3141];
@(posedge clk);
#1;data_in = testData6[3142];
@(posedge clk);
#1;data_in = testData6[3143];
@(posedge clk);
#1;data_in = testData6[3144];
@(posedge clk);
#1;data_in = testData6[3145];
@(posedge clk);
#1;data_in = testData6[3146];
@(posedge clk);
#1;data_in = testData6[3147];
@(posedge clk);
#1;data_in = testData6[3148];
@(posedge clk);
#1;data_in = testData6[3149];
@(posedge clk);
#1;data_in = testData6[3150];
@(posedge clk);
#1;data_in = testData6[3151];
@(posedge clk);
#1;data_in = testData6[3152];
@(posedge clk);
#1;data_in = testData6[3153];
@(posedge clk);
#1;data_in = testData6[3154];
@(posedge clk);
#1;data_in = testData6[3155];
@(posedge clk);
#1;data_in = testData6[3156];
@(posedge clk);
#1;data_in = testData6[3157];
@(posedge clk);
#1;data_in = testData6[3158];
@(posedge clk);
#1;data_in = testData6[3159];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[3160]; 
@(posedge clk);
#1;data_in = testData6[3161];
@(posedge clk);
#1;data_in = testData6[3162];
@(posedge clk);
#1;data_in = testData6[3163];
@(posedge clk);
#1;data_in = testData6[3164];
@(posedge clk);
#1;data_in = testData6[3165];
@(posedge clk);
#1;data_in = testData6[3166];
@(posedge clk);
#1;data_in = testData6[3167];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[3168];
@(posedge clk);
#1;data_in = testData6[3169];
@(posedge clk);
#1;data_in = testData6[3170];
@(posedge clk);
#1;data_in = testData6[3171];
@(posedge clk);
#1;data_in = testData6[3172];
@(posedge clk);
#1;data_in = testData6[3173];
@(posedge clk);
#1;data_in = testData6[3174];
@(posedge clk);
#1;data_in = testData6[3175];
@(posedge clk);
#1;data_in = testData6[3176];
@(posedge clk);
#1;data_in = testData6[3177];
@(posedge clk);
#1;data_in = testData6[3178];
@(posedge clk);
#1;data_in = testData6[3179];
@(posedge clk);
#1;data_in = testData6[3180];
@(posedge clk);
#1;data_in = testData6[3181];
@(posedge clk);
#1;data_in = testData6[3182];
@(posedge clk);
#1;data_in = testData6[3183];
@(posedge clk);
#1;data_in = testData6[3184];
@(posedge clk);
#1;data_in = testData6[3185];
@(posedge clk);
#1;data_in = testData6[3186];
@(posedge clk);
#1;data_in = testData6[3187];
@(posedge clk);
#1;data_in = testData6[3188];
@(posedge clk);
#1;data_in = testData6[3189];
@(posedge clk);
#1;data_in = testData6[3190];
@(posedge clk);
#1;data_in = testData6[3191];
@(posedge clk);
#1;data_in = testData6[3192];
@(posedge clk);
#1;data_in = testData6[3193];
@(posedge clk);
#1;data_in = testData6[3194];
@(posedge clk);
#1;data_in = testData6[3195];
@(posedge clk);
#1;data_in = testData6[3196];
@(posedge clk);
#1;data_in = testData6[3197];
@(posedge clk);
#1;data_in = testData6[3198];
@(posedge clk);
#1;data_in = testData6[3199];
@(posedge clk);
#1;data_in = testData6[3200];
@(posedge clk);
#1;data_in = testData6[3201];
@(posedge clk);
#1;data_in = testData6[3202];
@(posedge clk);
#1;data_in = testData6[3203];
@(posedge clk);
#1;data_in = testData6[3204];
@(posedge clk);
#1;data_in = testData6[3205];
@(posedge clk);
#1;data_in = testData6[3206];
@(posedge clk);
#1;data_in = testData6[3207];
@(posedge clk);
#1;data_in = testData6[3208];
@(posedge clk);
#1;data_in = testData6[3209];
@(posedge clk);
#1;data_in = testData6[3210];
@(posedge clk);
#1;data_in = testData6[3211];
@(posedge clk);
#1;data_in = testData6[3212];
@(posedge clk);
#1;data_in = testData6[3213];
@(posedge clk);
#1;data_in = testData6[3214];
@(posedge clk);
#1;data_in = testData6[3215];
@(posedge clk);
#1;data_in = testData6[3216];
@(posedge clk);
#1;data_in = testData6[3217];
@(posedge clk);
#1;data_in = testData6[3218];
@(posedge clk);
#1;data_in = testData6[3219];
@(posedge clk);
#1;data_in = testData6[3220];
@(posedge clk);
#1;data_in = testData6[3221];
@(posedge clk);
#1;data_in = testData6[3222];
@(posedge clk);
#1;data_in = testData6[3223];
@(posedge clk);
#1;data_in = testData6[3224];
@(posedge clk);
#1;data_in = testData6[3225];
@(posedge clk);
#1;data_in = testData6[3226];
@(posedge clk);
#1;data_in = testData6[3227];
@(posedge clk);
#1;data_in = testData6[3228];
@(posedge clk);
#1;data_in = testData6[3229];
@(posedge clk);
#1;data_in = testData6[3230];
@(posedge clk);
#1;data_in = testData6[3231];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[3232]; 
@(posedge clk);
#1;data_in = testData6[3233];
@(posedge clk);
#1;data_in = testData6[3234];
@(posedge clk);
#1;data_in = testData6[3235];
@(posedge clk);
#1;data_in = testData6[3236];
@(posedge clk);
#1;data_in = testData6[3237];
@(posedge clk);
#1;data_in = testData6[3238];
@(posedge clk);
#1;data_in = testData6[3239];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[3240];
@(posedge clk);
#1;data_in = testData6[3241];
@(posedge clk);
#1;data_in = testData6[3242];
@(posedge clk);
#1;data_in = testData6[3243];
@(posedge clk);
#1;data_in = testData6[3244];
@(posedge clk);
#1;data_in = testData6[3245];
@(posedge clk);
#1;data_in = testData6[3246];
@(posedge clk);
#1;data_in = testData6[3247];
@(posedge clk);
#1;data_in = testData6[3248];
@(posedge clk);
#1;data_in = testData6[3249];
@(posedge clk);
#1;data_in = testData6[3250];
@(posedge clk);
#1;data_in = testData6[3251];
@(posedge clk);
#1;data_in = testData6[3252];
@(posedge clk);
#1;data_in = testData6[3253];
@(posedge clk);
#1;data_in = testData6[3254];
@(posedge clk);
#1;data_in = testData6[3255];
@(posedge clk);
#1;data_in = testData6[3256];
@(posedge clk);
#1;data_in = testData6[3257];
@(posedge clk);
#1;data_in = testData6[3258];
@(posedge clk);
#1;data_in = testData6[3259];
@(posedge clk);
#1;data_in = testData6[3260];
@(posedge clk);
#1;data_in = testData6[3261];
@(posedge clk);
#1;data_in = testData6[3262];
@(posedge clk);
#1;data_in = testData6[3263];
@(posedge clk);
#1;data_in = testData6[3264];
@(posedge clk);
#1;data_in = testData6[3265];
@(posedge clk);
#1;data_in = testData6[3266];
@(posedge clk);
#1;data_in = testData6[3267];
@(posedge clk);
#1;data_in = testData6[3268];
@(posedge clk);
#1;data_in = testData6[3269];
@(posedge clk);
#1;data_in = testData6[3270];
@(posedge clk);
#1;data_in = testData6[3271];
@(posedge clk);
#1;data_in = testData6[3272];
@(posedge clk);
#1;data_in = testData6[3273];
@(posedge clk);
#1;data_in = testData6[3274];
@(posedge clk);
#1;data_in = testData6[3275];
@(posedge clk);
#1;data_in = testData6[3276];
@(posedge clk);
#1;data_in = testData6[3277];
@(posedge clk);
#1;data_in = testData6[3278];
@(posedge clk);
#1;data_in = testData6[3279];
@(posedge clk);
#1;data_in = testData6[3280];
@(posedge clk);
#1;data_in = testData6[3281];
@(posedge clk);
#1;data_in = testData6[3282];
@(posedge clk);
#1;data_in = testData6[3283];
@(posedge clk);
#1;data_in = testData6[3284];
@(posedge clk);
#1;data_in = testData6[3285];
@(posedge clk);
#1;data_in = testData6[3286];
@(posedge clk);
#1;data_in = testData6[3287];
@(posedge clk);
#1;data_in = testData6[3288];
@(posedge clk);
#1;data_in = testData6[3289];
@(posedge clk);
#1;data_in = testData6[3290];
@(posedge clk);
#1;data_in = testData6[3291];
@(posedge clk);
#1;data_in = testData6[3292];
@(posedge clk);
#1;data_in = testData6[3293];
@(posedge clk);
#1;data_in = testData6[3294];
@(posedge clk);
#1;data_in = testData6[3295];
@(posedge clk);
#1;data_in = testData6[3296];
@(posedge clk);
#1;data_in = testData6[3297];
@(posedge clk);
#1;data_in = testData6[3298];
@(posedge clk);
#1;data_in = testData6[3299];
@(posedge clk);
#1;data_in = testData6[3300];
@(posedge clk);
#1;data_in = testData6[3301];
@(posedge clk);
#1;data_in = testData6[3302];
@(posedge clk);
#1;data_in = testData6[3303];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[3304]; 
@(posedge clk);
#1;data_in = testData6[3305];
@(posedge clk);
#1;data_in = testData6[3306];
@(posedge clk);
#1;data_in = testData6[3307];
@(posedge clk);
#1;data_in = testData6[3308];
@(posedge clk);
#1;data_in = testData6[3309];
@(posedge clk);
#1;data_in = testData6[3310];
@(posedge clk);
#1;data_in = testData6[3311];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[3312];
@(posedge clk);
#1;data_in = testData6[3313];
@(posedge clk);
#1;data_in = testData6[3314];
@(posedge clk);
#1;data_in = testData6[3315];
@(posedge clk);
#1;data_in = testData6[3316];
@(posedge clk);
#1;data_in = testData6[3317];
@(posedge clk);
#1;data_in = testData6[3318];
@(posedge clk);
#1;data_in = testData6[3319];
@(posedge clk);
#1;data_in = testData6[3320];
@(posedge clk);
#1;data_in = testData6[3321];
@(posedge clk);
#1;data_in = testData6[3322];
@(posedge clk);
#1;data_in = testData6[3323];
@(posedge clk);
#1;data_in = testData6[3324];
@(posedge clk);
#1;data_in = testData6[3325];
@(posedge clk);
#1;data_in = testData6[3326];
@(posedge clk);
#1;data_in = testData6[3327];
@(posedge clk);
#1;data_in = testData6[3328];
@(posedge clk);
#1;data_in = testData6[3329];
@(posedge clk);
#1;data_in = testData6[3330];
@(posedge clk);
#1;data_in = testData6[3331];
@(posedge clk);
#1;data_in = testData6[3332];
@(posedge clk);
#1;data_in = testData6[3333];
@(posedge clk);
#1;data_in = testData6[3334];
@(posedge clk);
#1;data_in = testData6[3335];
@(posedge clk);
#1;data_in = testData6[3336];
@(posedge clk);
#1;data_in = testData6[3337];
@(posedge clk);
#1;data_in = testData6[3338];
@(posedge clk);
#1;data_in = testData6[3339];
@(posedge clk);
#1;data_in = testData6[3340];
@(posedge clk);
#1;data_in = testData6[3341];
@(posedge clk);
#1;data_in = testData6[3342];
@(posedge clk);
#1;data_in = testData6[3343];
@(posedge clk);
#1;data_in = testData6[3344];
@(posedge clk);
#1;data_in = testData6[3345];
@(posedge clk);
#1;data_in = testData6[3346];
@(posedge clk);
#1;data_in = testData6[3347];
@(posedge clk);
#1;data_in = testData6[3348];
@(posedge clk);
#1;data_in = testData6[3349];
@(posedge clk);
#1;data_in = testData6[3350];
@(posedge clk);
#1;data_in = testData6[3351];
@(posedge clk);
#1;data_in = testData6[3352];
@(posedge clk);
#1;data_in = testData6[3353];
@(posedge clk);
#1;data_in = testData6[3354];
@(posedge clk);
#1;data_in = testData6[3355];
@(posedge clk);
#1;data_in = testData6[3356];
@(posedge clk);
#1;data_in = testData6[3357];
@(posedge clk);
#1;data_in = testData6[3358];
@(posedge clk);
#1;data_in = testData6[3359];
@(posedge clk);
#1;data_in = testData6[3360];
@(posedge clk);
#1;data_in = testData6[3361];
@(posedge clk);
#1;data_in = testData6[3362];
@(posedge clk);
#1;data_in = testData6[3363];
@(posedge clk);
#1;data_in = testData6[3364];
@(posedge clk);
#1;data_in = testData6[3365];
@(posedge clk);
#1;data_in = testData6[3366];
@(posedge clk);
#1;data_in = testData6[3367];
@(posedge clk);
#1;data_in = testData6[3368];
@(posedge clk);
#1;data_in = testData6[3369];
@(posedge clk);
#1;data_in = testData6[3370];
@(posedge clk);
#1;data_in = testData6[3371];
@(posedge clk);
#1;data_in = testData6[3372];
@(posedge clk);
#1;data_in = testData6[3373];
@(posedge clk);
#1;data_in = testData6[3374];
@(posedge clk);
#1;data_in = testData6[3375];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[3376]; 
@(posedge clk);
#1;data_in = testData6[3377];
@(posedge clk);
#1;data_in = testData6[3378];
@(posedge clk);
#1;data_in = testData6[3379];
@(posedge clk);
#1;data_in = testData6[3380];
@(posedge clk);
#1;data_in = testData6[3381];
@(posedge clk);
#1;data_in = testData6[3382];
@(posedge clk);
#1;data_in = testData6[3383];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[3384];
@(posedge clk);
#1;data_in = testData6[3385];
@(posedge clk);
#1;data_in = testData6[3386];
@(posedge clk);
#1;data_in = testData6[3387];
@(posedge clk);
#1;data_in = testData6[3388];
@(posedge clk);
#1;data_in = testData6[3389];
@(posedge clk);
#1;data_in = testData6[3390];
@(posedge clk);
#1;data_in = testData6[3391];
@(posedge clk);
#1;data_in = testData6[3392];
@(posedge clk);
#1;data_in = testData6[3393];
@(posedge clk);
#1;data_in = testData6[3394];
@(posedge clk);
#1;data_in = testData6[3395];
@(posedge clk);
#1;data_in = testData6[3396];
@(posedge clk);
#1;data_in = testData6[3397];
@(posedge clk);
#1;data_in = testData6[3398];
@(posedge clk);
#1;data_in = testData6[3399];
@(posedge clk);
#1;data_in = testData6[3400];
@(posedge clk);
#1;data_in = testData6[3401];
@(posedge clk);
#1;data_in = testData6[3402];
@(posedge clk);
#1;data_in = testData6[3403];
@(posedge clk);
#1;data_in = testData6[3404];
@(posedge clk);
#1;data_in = testData6[3405];
@(posedge clk);
#1;data_in = testData6[3406];
@(posedge clk);
#1;data_in = testData6[3407];
@(posedge clk);
#1;data_in = testData6[3408];
@(posedge clk);
#1;data_in = testData6[3409];
@(posedge clk);
#1;data_in = testData6[3410];
@(posedge clk);
#1;data_in = testData6[3411];
@(posedge clk);
#1;data_in = testData6[3412];
@(posedge clk);
#1;data_in = testData6[3413];
@(posedge clk);
#1;data_in = testData6[3414];
@(posedge clk);
#1;data_in = testData6[3415];
@(posedge clk);
#1;data_in = testData6[3416];
@(posedge clk);
#1;data_in = testData6[3417];
@(posedge clk);
#1;data_in = testData6[3418];
@(posedge clk);
#1;data_in = testData6[3419];
@(posedge clk);
#1;data_in = testData6[3420];
@(posedge clk);
#1;data_in = testData6[3421];
@(posedge clk);
#1;data_in = testData6[3422];
@(posedge clk);
#1;data_in = testData6[3423];
@(posedge clk);
#1;data_in = testData6[3424];
@(posedge clk);
#1;data_in = testData6[3425];
@(posedge clk);
#1;data_in = testData6[3426];
@(posedge clk);
#1;data_in = testData6[3427];
@(posedge clk);
#1;data_in = testData6[3428];
@(posedge clk);
#1;data_in = testData6[3429];
@(posedge clk);
#1;data_in = testData6[3430];
@(posedge clk);
#1;data_in = testData6[3431];
@(posedge clk);
#1;data_in = testData6[3432];
@(posedge clk);
#1;data_in = testData6[3433];
@(posedge clk);
#1;data_in = testData6[3434];
@(posedge clk);
#1;data_in = testData6[3435];
@(posedge clk);
#1;data_in = testData6[3436];
@(posedge clk);
#1;data_in = testData6[3437];
@(posedge clk);
#1;data_in = testData6[3438];
@(posedge clk);
#1;data_in = testData6[3439];
@(posedge clk);
#1;data_in = testData6[3440];
@(posedge clk);
#1;data_in = testData6[3441];
@(posedge clk);
#1;data_in = testData6[3442];
@(posedge clk);
#1;data_in = testData6[3443];
@(posedge clk);
#1;data_in = testData6[3444];
@(posedge clk);
#1;data_in = testData6[3445];
@(posedge clk);
#1;data_in = testData6[3446];
@(posedge clk);
#1;data_in = testData6[3447];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[3448]; 
@(posedge clk);
#1;data_in = testData6[3449];
@(posedge clk);
#1;data_in = testData6[3450];
@(posedge clk);
#1;data_in = testData6[3451];
@(posedge clk);
#1;data_in = testData6[3452];
@(posedge clk);
#1;data_in = testData6[3453];
@(posedge clk);
#1;data_in = testData6[3454];
@(posedge clk);
#1;data_in = testData6[3455];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[3456];
@(posedge clk);
#1;data_in = testData6[3457];
@(posedge clk);
#1;data_in = testData6[3458];
@(posedge clk);
#1;data_in = testData6[3459];
@(posedge clk);
#1;data_in = testData6[3460];
@(posedge clk);
#1;data_in = testData6[3461];
@(posedge clk);
#1;data_in = testData6[3462];
@(posedge clk);
#1;data_in = testData6[3463];
@(posedge clk);
#1;data_in = testData6[3464];
@(posedge clk);
#1;data_in = testData6[3465];
@(posedge clk);
#1;data_in = testData6[3466];
@(posedge clk);
#1;data_in = testData6[3467];
@(posedge clk);
#1;data_in = testData6[3468];
@(posedge clk);
#1;data_in = testData6[3469];
@(posedge clk);
#1;data_in = testData6[3470];
@(posedge clk);
#1;data_in = testData6[3471];
@(posedge clk);
#1;data_in = testData6[3472];
@(posedge clk);
#1;data_in = testData6[3473];
@(posedge clk);
#1;data_in = testData6[3474];
@(posedge clk);
#1;data_in = testData6[3475];
@(posedge clk);
#1;data_in = testData6[3476];
@(posedge clk);
#1;data_in = testData6[3477];
@(posedge clk);
#1;data_in = testData6[3478];
@(posedge clk);
#1;data_in = testData6[3479];
@(posedge clk);
#1;data_in = testData6[3480];
@(posedge clk);
#1;data_in = testData6[3481];
@(posedge clk);
#1;data_in = testData6[3482];
@(posedge clk);
#1;data_in = testData6[3483];
@(posedge clk);
#1;data_in = testData6[3484];
@(posedge clk);
#1;data_in = testData6[3485];
@(posedge clk);
#1;data_in = testData6[3486];
@(posedge clk);
#1;data_in = testData6[3487];
@(posedge clk);
#1;data_in = testData6[3488];
@(posedge clk);
#1;data_in = testData6[3489];
@(posedge clk);
#1;data_in = testData6[3490];
@(posedge clk);
#1;data_in = testData6[3491];
@(posedge clk);
#1;data_in = testData6[3492];
@(posedge clk);
#1;data_in = testData6[3493];
@(posedge clk);
#1;data_in = testData6[3494];
@(posedge clk);
#1;data_in = testData6[3495];
@(posedge clk);
#1;data_in = testData6[3496];
@(posedge clk);
#1;data_in = testData6[3497];
@(posedge clk);
#1;data_in = testData6[3498];
@(posedge clk);
#1;data_in = testData6[3499];
@(posedge clk);
#1;data_in = testData6[3500];
@(posedge clk);
#1;data_in = testData6[3501];
@(posedge clk);
#1;data_in = testData6[3502];
@(posedge clk);
#1;data_in = testData6[3503];
@(posedge clk);
#1;data_in = testData6[3504];
@(posedge clk);
#1;data_in = testData6[3505];
@(posedge clk);
#1;data_in = testData6[3506];
@(posedge clk);
#1;data_in = testData6[3507];
@(posedge clk);
#1;data_in = testData6[3508];
@(posedge clk);
#1;data_in = testData6[3509];
@(posedge clk);
#1;data_in = testData6[3510];
@(posedge clk);
#1;data_in = testData6[3511];
@(posedge clk);
#1;data_in = testData6[3512];
@(posedge clk);
#1;data_in = testData6[3513];
@(posedge clk);
#1;data_in = testData6[3514];
@(posedge clk);
#1;data_in = testData6[3515];
@(posedge clk);
#1;data_in = testData6[3516];
@(posedge clk);
#1;data_in = testData6[3517];
@(posedge clk);
#1;data_in = testData6[3518];
@(posedge clk);
#1;data_in = testData6[3519];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[3520]; 
@(posedge clk);
#1;data_in = testData6[3521];
@(posedge clk);
#1;data_in = testData6[3522];
@(posedge clk);
#1;data_in = testData6[3523];
@(posedge clk);
#1;data_in = testData6[3524];
@(posedge clk);
#1;data_in = testData6[3525];
@(posedge clk);
#1;data_in = testData6[3526];
@(posedge clk);
#1;data_in = testData6[3527];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[3528];
@(posedge clk);
#1;data_in = testData6[3529];
@(posedge clk);
#1;data_in = testData6[3530];
@(posedge clk);
#1;data_in = testData6[3531];
@(posedge clk);
#1;data_in = testData6[3532];
@(posedge clk);
#1;data_in = testData6[3533];
@(posedge clk);
#1;data_in = testData6[3534];
@(posedge clk);
#1;data_in = testData6[3535];
@(posedge clk);
#1;data_in = testData6[3536];
@(posedge clk);
#1;data_in = testData6[3537];
@(posedge clk);
#1;data_in = testData6[3538];
@(posedge clk);
#1;data_in = testData6[3539];
@(posedge clk);
#1;data_in = testData6[3540];
@(posedge clk);
#1;data_in = testData6[3541];
@(posedge clk);
#1;data_in = testData6[3542];
@(posedge clk);
#1;data_in = testData6[3543];
@(posedge clk);
#1;data_in = testData6[3544];
@(posedge clk);
#1;data_in = testData6[3545];
@(posedge clk);
#1;data_in = testData6[3546];
@(posedge clk);
#1;data_in = testData6[3547];
@(posedge clk);
#1;data_in = testData6[3548];
@(posedge clk);
#1;data_in = testData6[3549];
@(posedge clk);
#1;data_in = testData6[3550];
@(posedge clk);
#1;data_in = testData6[3551];
@(posedge clk);
#1;data_in = testData6[3552];
@(posedge clk);
#1;data_in = testData6[3553];
@(posedge clk);
#1;data_in = testData6[3554];
@(posedge clk);
#1;data_in = testData6[3555];
@(posedge clk);
#1;data_in = testData6[3556];
@(posedge clk);
#1;data_in = testData6[3557];
@(posedge clk);
#1;data_in = testData6[3558];
@(posedge clk);
#1;data_in = testData6[3559];
@(posedge clk);
#1;data_in = testData6[3560];
@(posedge clk);
#1;data_in = testData6[3561];
@(posedge clk);
#1;data_in = testData6[3562];
@(posedge clk);
#1;data_in = testData6[3563];
@(posedge clk);
#1;data_in = testData6[3564];
@(posedge clk);
#1;data_in = testData6[3565];
@(posedge clk);
#1;data_in = testData6[3566];
@(posedge clk);
#1;data_in = testData6[3567];
@(posedge clk);
#1;data_in = testData6[3568];
@(posedge clk);
#1;data_in = testData6[3569];
@(posedge clk);
#1;data_in = testData6[3570];
@(posedge clk);
#1;data_in = testData6[3571];
@(posedge clk);
#1;data_in = testData6[3572];
@(posedge clk);
#1;data_in = testData6[3573];
@(posedge clk);
#1;data_in = testData6[3574];
@(posedge clk);
#1;data_in = testData6[3575];
@(posedge clk);
#1;data_in = testData6[3576];
@(posedge clk);
#1;data_in = testData6[3577];
@(posedge clk);
#1;data_in = testData6[3578];
@(posedge clk);
#1;data_in = testData6[3579];
@(posedge clk);
#1;data_in = testData6[3580];
@(posedge clk);
#1;data_in = testData6[3581];
@(posedge clk);
#1;data_in = testData6[3582];
@(posedge clk);
#1;data_in = testData6[3583];
@(posedge clk);
#1;data_in = testData6[3584];
@(posedge clk);
#1;data_in = testData6[3585];
@(posedge clk);
#1;data_in = testData6[3586];
@(posedge clk);
#1;data_in = testData6[3587];
@(posedge clk);
#1;data_in = testData6[3588];
@(posedge clk);
#1;data_in = testData6[3589];
@(posedge clk);
#1;data_in = testData6[3590];
@(posedge clk);
#1;data_in = testData6[3591];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[3592]; 
@(posedge clk);
#1;data_in = testData6[3593];
@(posedge clk);
#1;data_in = testData6[3594];
@(posedge clk);
#1;data_in = testData6[3595];
@(posedge clk);
#1;data_in = testData6[3596];
@(posedge clk);
#1;data_in = testData6[3597];
@(posedge clk);
#1;data_in = testData6[3598];
@(posedge clk);
#1;data_in = testData6[3599];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[3600];
@(posedge clk);
#1;data_in = testData6[3601];
@(posedge clk);
#1;data_in = testData6[3602];
@(posedge clk);
#1;data_in = testData6[3603];
@(posedge clk);
#1;data_in = testData6[3604];
@(posedge clk);
#1;data_in = testData6[3605];
@(posedge clk);
#1;data_in = testData6[3606];
@(posedge clk);
#1;data_in = testData6[3607];
@(posedge clk);
#1;data_in = testData6[3608];
@(posedge clk);
#1;data_in = testData6[3609];
@(posedge clk);
#1;data_in = testData6[3610];
@(posedge clk);
#1;data_in = testData6[3611];
@(posedge clk);
#1;data_in = testData6[3612];
@(posedge clk);
#1;data_in = testData6[3613];
@(posedge clk);
#1;data_in = testData6[3614];
@(posedge clk);
#1;data_in = testData6[3615];
@(posedge clk);
#1;data_in = testData6[3616];
@(posedge clk);
#1;data_in = testData6[3617];
@(posedge clk);
#1;data_in = testData6[3618];
@(posedge clk);
#1;data_in = testData6[3619];
@(posedge clk);
#1;data_in = testData6[3620];
@(posedge clk);
#1;data_in = testData6[3621];
@(posedge clk);
#1;data_in = testData6[3622];
@(posedge clk);
#1;data_in = testData6[3623];
@(posedge clk);
#1;data_in = testData6[3624];
@(posedge clk);
#1;data_in = testData6[3625];
@(posedge clk);
#1;data_in = testData6[3626];
@(posedge clk);
#1;data_in = testData6[3627];
@(posedge clk);
#1;data_in = testData6[3628];
@(posedge clk);
#1;data_in = testData6[3629];
@(posedge clk);
#1;data_in = testData6[3630];
@(posedge clk);
#1;data_in = testData6[3631];
@(posedge clk);
#1;data_in = testData6[3632];
@(posedge clk);
#1;data_in = testData6[3633];
@(posedge clk);
#1;data_in = testData6[3634];
@(posedge clk);
#1;data_in = testData6[3635];
@(posedge clk);
#1;data_in = testData6[3636];
@(posedge clk);
#1;data_in = testData6[3637];
@(posedge clk);
#1;data_in = testData6[3638];
@(posedge clk);
#1;data_in = testData6[3639];
@(posedge clk);
#1;data_in = testData6[3640];
@(posedge clk);
#1;data_in = testData6[3641];
@(posedge clk);
#1;data_in = testData6[3642];
@(posedge clk);
#1;data_in = testData6[3643];
@(posedge clk);
#1;data_in = testData6[3644];
@(posedge clk);
#1;data_in = testData6[3645];
@(posedge clk);
#1;data_in = testData6[3646];
@(posedge clk);
#1;data_in = testData6[3647];
@(posedge clk);
#1;data_in = testData6[3648];
@(posedge clk);
#1;data_in = testData6[3649];
@(posedge clk);
#1;data_in = testData6[3650];
@(posedge clk);
#1;data_in = testData6[3651];
@(posedge clk);
#1;data_in = testData6[3652];
@(posedge clk);
#1;data_in = testData6[3653];
@(posedge clk);
#1;data_in = testData6[3654];
@(posedge clk);
#1;data_in = testData6[3655];
@(posedge clk);
#1;data_in = testData6[3656];
@(posedge clk);
#1;data_in = testData6[3657];
@(posedge clk);
#1;data_in = testData6[3658];
@(posedge clk);
#1;data_in = testData6[3659];
@(posedge clk);
#1;data_in = testData6[3660];
@(posedge clk);
#1;data_in = testData6[3661];
@(posedge clk);
#1;data_in = testData6[3662];
@(posedge clk);
#1;data_in = testData6[3663];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[3664]; 
@(posedge clk);
#1;data_in = testData6[3665];
@(posedge clk);
#1;data_in = testData6[3666];
@(posedge clk);
#1;data_in = testData6[3667];
@(posedge clk);
#1;data_in = testData6[3668];
@(posedge clk);
#1;data_in = testData6[3669];
@(posedge clk);
#1;data_in = testData6[3670];
@(posedge clk);
#1;data_in = testData6[3671];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
// Testbench, with parameters k=8, p=8, b=8, g=1

module tb5();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_8_8_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

logic [7:0] testData5[3271:0];
   //read input from C file inputDatapart1     
 initial $readmemh("proj3_inputDatatb5", testData5);
 integer i;
 integer filehandle=$fopen("proj3_outValuestb5");
  initial begin 
  $monitor("Data in : %x",data_in);       
start  = 0; reset  = 1; data_in = 8'bx;
 @(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData5[0];
@(posedge clk);
#1;data_in = testData5[1];
@(posedge clk);
#1;data_in = testData5[2];
@(posedge clk);
#1;data_in = testData5[3];
@(posedge clk);
#1;data_in = testData5[4];
@(posedge clk);
#1;data_in = testData5[5];
@(posedge clk);
#1;data_in = testData5[6];
@(posedge clk);
#1;data_in = testData5[7];
@(posedge clk);
#1;data_in = testData5[8];
@(posedge clk);
#1;data_in = testData5[9];
@(posedge clk);
#1;data_in = testData5[10];
@(posedge clk);
#1;data_in = testData5[11];
@(posedge clk);
#1;data_in = testData5[12];
@(posedge clk);
#1;data_in = testData5[13];
@(posedge clk);
#1;data_in = testData5[14];
@(posedge clk);
#1;data_in = testData5[15];
@(posedge clk);
#1;data_in = testData5[16];
@(posedge clk);
#1;data_in = testData5[17];
@(posedge clk);
#1;data_in = testData5[18];
@(posedge clk);
#1;data_in = testData5[19];
@(posedge clk);
#1;data_in = testData5[20];
@(posedge clk);
#1;data_in = testData5[21];
@(posedge clk);
#1;data_in = testData5[22];
@(posedge clk);
#1;data_in = testData5[23];
@(posedge clk);
#1;data_in = testData5[24];
@(posedge clk);
#1;data_in = testData5[25];
@(posedge clk);
#1;data_in = testData5[26];
@(posedge clk);
#1;data_in = testData5[27];
@(posedge clk);
#1;data_in = testData5[28];
@(posedge clk);
#1;data_in = testData5[29];
@(posedge clk);
#1;data_in = testData5[30];
@(posedge clk);
#1;data_in = testData5[31];
@(posedge clk);
#1;data_in = testData5[32];
@(posedge clk);
#1;data_in = testData5[33];
@(posedge clk);
#1;data_in = testData5[34];
@(posedge clk);
#1;data_in = testData5[35];
@(posedge clk);
#1;data_in = testData5[36];
@(posedge clk);
#1;data_in = testData5[37];
@(posedge clk);
#1;data_in = testData5[38];
@(posedge clk);
#1;data_in = testData5[39];
@(posedge clk);
#1;data_in = testData5[40];
@(posedge clk);
#1;data_in = testData5[41];
@(posedge clk);
#1;data_in = testData5[42];
@(posedge clk);
#1;data_in = testData5[43];
@(posedge clk);
#1;data_in = testData5[44];
@(posedge clk);
#1;data_in = testData5[45];
@(posedge clk);
#1;data_in = testData5[46];
@(posedge clk);
#1;data_in = testData5[47];
@(posedge clk);
#1;data_in = testData5[48];
@(posedge clk);
#1;data_in = testData5[49];
@(posedge clk);
#1;data_in = testData5[50];
@(posedge clk);
#1;data_in = testData5[51];
@(posedge clk);
#1;data_in = testData5[52];
@(posedge clk);
#1;data_in = testData5[53];
@(posedge clk);
#1;data_in = testData5[54];
@(posedge clk);
#1;data_in = testData5[55];
@(posedge clk);
#1;data_in = testData5[56];
@(posedge clk);
#1;data_in = testData5[57];
@(posedge clk);
#1;data_in = testData5[58];
@(posedge clk);
#1;data_in = testData5[59];
@(posedge clk);
#1;data_in = testData5[60];
@(posedge clk);
#1;data_in = testData5[61];
@(posedge clk);
#1;data_in = testData5[62];
@(posedge clk);
#1;data_in = testData5[63];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData5[64]; 
@(posedge clk);
#1;data_in = testData5[65];
@(posedge clk);
#1;data_in = testData5[66];
@(posedge clk);
#1;data_in = testData5[67];
@(posedge clk);
#1;data_in = testData5[68];
@(posedge clk);
#1;data_in = testData5[69];
@(posedge clk);
#1;data_in = testData5[70];
@(posedge clk);
#1;data_in = testData5[71];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[72]; 
@(posedge clk);
#1;data_in = testData5[73];
@(posedge clk);
#1;data_in = testData5[74];
@(posedge clk);
#1;data_in = testData5[75];
@(posedge clk);
#1;data_in = testData5[76];
@(posedge clk);
#1;data_in = testData5[77];
@(posedge clk);
#1;data_in = testData5[78];
@(posedge clk);
#1;data_in = testData5[79];
@(posedge clk);
#1;data_in = testData5[80];
@(posedge clk);
#1;data_in = testData5[81];
@(posedge clk);
#1;data_in = testData5[82];
@(posedge clk);
#1;data_in = testData5[83];
@(posedge clk);
#1;data_in = testData5[84];
@(posedge clk);
#1;data_in = testData5[85];
@(posedge clk);
#1;data_in = testData5[86];
@(posedge clk);
#1;data_in = testData5[87];
@(posedge clk);
#1;data_in = testData5[88];
@(posedge clk);
#1;data_in = testData5[89];
@(posedge clk);
#1;data_in = testData5[90];
@(posedge clk);
#1;data_in = testData5[91];
@(posedge clk);
#1;data_in = testData5[92];
@(posedge clk);
#1;data_in = testData5[93];
@(posedge clk);
#1;data_in = testData5[94];
@(posedge clk);
#1;data_in = testData5[95];
@(posedge clk);
#1;data_in = testData5[96];
@(posedge clk);
#1;data_in = testData5[97];
@(posedge clk);
#1;data_in = testData5[98];
@(posedge clk);
#1;data_in = testData5[99];
@(posedge clk);
#1;data_in = testData5[100];
@(posedge clk);
#1;data_in = testData5[101];
@(posedge clk);
#1;data_in = testData5[102];
@(posedge clk);
#1;data_in = testData5[103];
@(posedge clk);
#1;data_in = testData5[104];
@(posedge clk);
#1;data_in = testData5[105];
@(posedge clk);
#1;data_in = testData5[106];
@(posedge clk);
#1;data_in = testData5[107];
@(posedge clk);
#1;data_in = testData5[108];
@(posedge clk);
#1;data_in = testData5[109];
@(posedge clk);
#1;data_in = testData5[110];
@(posedge clk);
#1;data_in = testData5[111];
@(posedge clk);
#1;data_in = testData5[112];
@(posedge clk);
#1;data_in = testData5[113];
@(posedge clk);
#1;data_in = testData5[114];
@(posedge clk);
#1;data_in = testData5[115];
@(posedge clk);
#1;data_in = testData5[116];
@(posedge clk);
#1;data_in = testData5[117];
@(posedge clk);
#1;data_in = testData5[118];
@(posedge clk);
#1;data_in = testData5[119];
@(posedge clk);
#1;data_in = testData5[120];
@(posedge clk);
#1;data_in = testData5[121];
@(posedge clk);
#1;data_in = testData5[122];
@(posedge clk);
#1;data_in = testData5[123];
@(posedge clk);
#1;data_in = testData5[124];
@(posedge clk);
#1;data_in = testData5[125];
@(posedge clk);
#1;data_in = testData5[126];
@(posedge clk);
#1;data_in = testData5[127];
@(posedge clk);
#1;data_in = testData5[128];
@(posedge clk);
#1;data_in = testData5[129];
@(posedge clk);
#1;data_in = testData5[130];
@(posedge clk);
#1;data_in = testData5[131];
@(posedge clk);
#1;data_in = testData5[132];
@(posedge clk);
#1;data_in = testData5[133];
@(posedge clk);
#1;data_in = testData5[134];
@(posedge clk);
#1;data_in = testData5[135];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[136]; 
@(posedge clk);
#1;data_in = testData5[137];
@(posedge clk);
#1;data_in = testData5[138];
@(posedge clk);
#1;data_in = testData5[139];
@(posedge clk);
#1;data_in = testData5[140];
@(posedge clk);
#1;data_in = testData5[141];
@(posedge clk);
#1;data_in = testData5[142];
@(posedge clk);
#1;data_in = testData5[143];
@(posedge clk);
#1;data_in = testData5[144];
@(posedge clk);
#1;data_in = testData5[145];
@(posedge clk);
#1;data_in = testData5[146];
@(posedge clk);
#1;data_in = testData5[147];
@(posedge clk);
#1;data_in = testData5[148];
@(posedge clk);
#1;data_in = testData5[149];
@(posedge clk);
#1;data_in = testData5[150];
@(posedge clk);
#1;data_in = testData5[151];
@(posedge clk);
#1;data_in = testData5[152];
@(posedge clk);
#1;data_in = testData5[153];
@(posedge clk);
#1;data_in = testData5[154];
@(posedge clk);
#1;data_in = testData5[155];
@(posedge clk);
#1;data_in = testData5[156];
@(posedge clk);
#1;data_in = testData5[157];
@(posedge clk);
#1;data_in = testData5[158];
@(posedge clk);
#1;data_in = testData5[159];
@(posedge clk);
#1;data_in = testData5[160];
@(posedge clk);
#1;data_in = testData5[161];
@(posedge clk);
#1;data_in = testData5[162];
@(posedge clk);
#1;data_in = testData5[163];
@(posedge clk);
#1;data_in = testData5[164];
@(posedge clk);
#1;data_in = testData5[165];
@(posedge clk);
#1;data_in = testData5[166];
@(posedge clk);
#1;data_in = testData5[167];
@(posedge clk);
#1;data_in = testData5[168];
@(posedge clk);
#1;data_in = testData5[169];
@(posedge clk);
#1;data_in = testData5[170];
@(posedge clk);
#1;data_in = testData5[171];
@(posedge clk);
#1;data_in = testData5[172];
@(posedge clk);
#1;data_in = testData5[173];
@(posedge clk);
#1;data_in = testData5[174];
@(posedge clk);
#1;data_in = testData5[175];
@(posedge clk);
#1;data_in = testData5[176];
@(posedge clk);
#1;data_in = testData5[177];
@(posedge clk);
#1;data_in = testData5[178];
@(posedge clk);
#1;data_in = testData5[179];
@(posedge clk);
#1;data_in = testData5[180];
@(posedge clk);
#1;data_in = testData5[181];
@(posedge clk);
#1;data_in = testData5[182];
@(posedge clk);
#1;data_in = testData5[183];
@(posedge clk);
#1;data_in = testData5[184];
@(posedge clk);
#1;data_in = testData5[185];
@(posedge clk);
#1;data_in = testData5[186];
@(posedge clk);
#1;data_in = testData5[187];
@(posedge clk);
#1;data_in = testData5[188];
@(posedge clk);
#1;data_in = testData5[189];
@(posedge clk);
#1;data_in = testData5[190];
@(posedge clk);
#1;data_in = testData5[191];
@(posedge clk);
#1;data_in = testData5[192];
@(posedge clk);
#1;data_in = testData5[193];
@(posedge clk);
#1;data_in = testData5[194];
@(posedge clk);
#1;data_in = testData5[195];
@(posedge clk);
#1;data_in = testData5[196];
@(posedge clk);
#1;data_in = testData5[197];
@(posedge clk);
#1;data_in = testData5[198];
@(posedge clk);
#1;data_in = testData5[199];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[200]; 
@(posedge clk);
#1;data_in = testData5[201];
@(posedge clk);
#1;data_in = testData5[202];
@(posedge clk);
#1;data_in = testData5[203];
@(posedge clk);
#1;data_in = testData5[204];
@(posedge clk);
#1;data_in = testData5[205];
@(posedge clk);
#1;data_in = testData5[206];
@(posedge clk);
#1;data_in = testData5[207];
@(posedge clk);
#1;data_in = testData5[208];
@(posedge clk);
#1;data_in = testData5[209];
@(posedge clk);
#1;data_in = testData5[210];
@(posedge clk);
#1;data_in = testData5[211];
@(posedge clk);
#1;data_in = testData5[212];
@(posedge clk);
#1;data_in = testData5[213];
@(posedge clk);
#1;data_in = testData5[214];
@(posedge clk);
#1;data_in = testData5[215];
@(posedge clk);
#1;data_in = testData5[216];
@(posedge clk);
#1;data_in = testData5[217];
@(posedge clk);
#1;data_in = testData5[218];
@(posedge clk);
#1;data_in = testData5[219];
@(posedge clk);
#1;data_in = testData5[220];
@(posedge clk);
#1;data_in = testData5[221];
@(posedge clk);
#1;data_in = testData5[222];
@(posedge clk);
#1;data_in = testData5[223];
@(posedge clk);
#1;data_in = testData5[224];
@(posedge clk);
#1;data_in = testData5[225];
@(posedge clk);
#1;data_in = testData5[226];
@(posedge clk);
#1;data_in = testData5[227];
@(posedge clk);
#1;data_in = testData5[228];
@(posedge clk);
#1;data_in = testData5[229];
@(posedge clk);
#1;data_in = testData5[230];
@(posedge clk);
#1;data_in = testData5[231];
@(posedge clk);
#1;data_in = testData5[232];
@(posedge clk);
#1;data_in = testData5[233];
@(posedge clk);
#1;data_in = testData5[234];
@(posedge clk);
#1;data_in = testData5[235];
@(posedge clk);
#1;data_in = testData5[236];
@(posedge clk);
#1;data_in = testData5[237];
@(posedge clk);
#1;data_in = testData5[238];
@(posedge clk);
#1;data_in = testData5[239];
@(posedge clk);
#1;data_in = testData5[240];
@(posedge clk);
#1;data_in = testData5[241];
@(posedge clk);
#1;data_in = testData5[242];
@(posedge clk);
#1;data_in = testData5[243];
@(posedge clk);
#1;data_in = testData5[244];
@(posedge clk);
#1;data_in = testData5[245];
@(posedge clk);
#1;data_in = testData5[246];
@(posedge clk);
#1;data_in = testData5[247];
@(posedge clk);
#1;data_in = testData5[248];
@(posedge clk);
#1;data_in = testData5[249];
@(posedge clk);
#1;data_in = testData5[250];
@(posedge clk);
#1;data_in = testData5[251];
@(posedge clk);
#1;data_in = testData5[252];
@(posedge clk);
#1;data_in = testData5[253];
@(posedge clk);
#1;data_in = testData5[254];
@(posedge clk);
#1;data_in = testData5[255];
@(posedge clk);
#1;data_in = testData5[256];
@(posedge clk);
#1;data_in = testData5[257];
@(posedge clk);
#1;data_in = testData5[258];
@(posedge clk);
#1;data_in = testData5[259];
@(posedge clk);
#1;data_in = testData5[260];
@(posedge clk);
#1;data_in = testData5[261];
@(posedge clk);
#1;data_in = testData5[262];
@(posedge clk);
#1;data_in = testData5[263];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[264]; 
@(posedge clk);
#1;data_in = testData5[265];
@(posedge clk);
#1;data_in = testData5[266];
@(posedge clk);
#1;data_in = testData5[267];
@(posedge clk);
#1;data_in = testData5[268];
@(posedge clk);
#1;data_in = testData5[269];
@(posedge clk);
#1;data_in = testData5[270];
@(posedge clk);
#1;data_in = testData5[271];
@(posedge clk);
#1;data_in = testData5[272];
@(posedge clk);
#1;data_in = testData5[273];
@(posedge clk);
#1;data_in = testData5[274];
@(posedge clk);
#1;data_in = testData5[275];
@(posedge clk);
#1;data_in = testData5[276];
@(posedge clk);
#1;data_in = testData5[277];
@(posedge clk);
#1;data_in = testData5[278];
@(posedge clk);
#1;data_in = testData5[279];
@(posedge clk);
#1;data_in = testData5[280];
@(posedge clk);
#1;data_in = testData5[281];
@(posedge clk);
#1;data_in = testData5[282];
@(posedge clk);
#1;data_in = testData5[283];
@(posedge clk);
#1;data_in = testData5[284];
@(posedge clk);
#1;data_in = testData5[285];
@(posedge clk);
#1;data_in = testData5[286];
@(posedge clk);
#1;data_in = testData5[287];
@(posedge clk);
#1;data_in = testData5[288];
@(posedge clk);
#1;data_in = testData5[289];
@(posedge clk);
#1;data_in = testData5[290];
@(posedge clk);
#1;data_in = testData5[291];
@(posedge clk);
#1;data_in = testData5[292];
@(posedge clk);
#1;data_in = testData5[293];
@(posedge clk);
#1;data_in = testData5[294];
@(posedge clk);
#1;data_in = testData5[295];
@(posedge clk);
#1;data_in = testData5[296];
@(posedge clk);
#1;data_in = testData5[297];
@(posedge clk);
#1;data_in = testData5[298];
@(posedge clk);
#1;data_in = testData5[299];
@(posedge clk);
#1;data_in = testData5[300];
@(posedge clk);
#1;data_in = testData5[301];
@(posedge clk);
#1;data_in = testData5[302];
@(posedge clk);
#1;data_in = testData5[303];
@(posedge clk);
#1;data_in = testData5[304];
@(posedge clk);
#1;data_in = testData5[305];
@(posedge clk);
#1;data_in = testData5[306];
@(posedge clk);
#1;data_in = testData5[307];
@(posedge clk);
#1;data_in = testData5[308];
@(posedge clk);
#1;data_in = testData5[309];
@(posedge clk);
#1;data_in = testData5[310];
@(posedge clk);
#1;data_in = testData5[311];
@(posedge clk);
#1;data_in = testData5[312];
@(posedge clk);
#1;data_in = testData5[313];
@(posedge clk);
#1;data_in = testData5[314];
@(posedge clk);
#1;data_in = testData5[315];
@(posedge clk);
#1;data_in = testData5[316];
@(posedge clk);
#1;data_in = testData5[317];
@(posedge clk);
#1;data_in = testData5[318];
@(posedge clk);
#1;data_in = testData5[319];
@(posedge clk);
#1;data_in = testData5[320];
@(posedge clk);
#1;data_in = testData5[321];
@(posedge clk);
#1;data_in = testData5[322];
@(posedge clk);
#1;data_in = testData5[323];
@(posedge clk);
#1;data_in = testData5[324];
@(posedge clk);
#1;data_in = testData5[325];
@(posedge clk);
#1;data_in = testData5[326];
@(posedge clk);
#1;data_in = testData5[327];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[328]; 
@(posedge clk);
#1;data_in = testData5[329];
@(posedge clk);
#1;data_in = testData5[330];
@(posedge clk);
#1;data_in = testData5[331];
@(posedge clk);
#1;data_in = testData5[332];
@(posedge clk);
#1;data_in = testData5[333];
@(posedge clk);
#1;data_in = testData5[334];
@(posedge clk);
#1;data_in = testData5[335];
@(posedge clk);
#1;data_in = testData5[336];
@(posedge clk);
#1;data_in = testData5[337];
@(posedge clk);
#1;data_in = testData5[338];
@(posedge clk);
#1;data_in = testData5[339];
@(posedge clk);
#1;data_in = testData5[340];
@(posedge clk);
#1;data_in = testData5[341];
@(posedge clk);
#1;data_in = testData5[342];
@(posedge clk);
#1;data_in = testData5[343];
@(posedge clk);
#1;data_in = testData5[344];
@(posedge clk);
#1;data_in = testData5[345];
@(posedge clk);
#1;data_in = testData5[346];
@(posedge clk);
#1;data_in = testData5[347];
@(posedge clk);
#1;data_in = testData5[348];
@(posedge clk);
#1;data_in = testData5[349];
@(posedge clk);
#1;data_in = testData5[350];
@(posedge clk);
#1;data_in = testData5[351];
@(posedge clk);
#1;data_in = testData5[352];
@(posedge clk);
#1;data_in = testData5[353];
@(posedge clk);
#1;data_in = testData5[354];
@(posedge clk);
#1;data_in = testData5[355];
@(posedge clk);
#1;data_in = testData5[356];
@(posedge clk);
#1;data_in = testData5[357];
@(posedge clk);
#1;data_in = testData5[358];
@(posedge clk);
#1;data_in = testData5[359];
@(posedge clk);
#1;data_in = testData5[360];
@(posedge clk);
#1;data_in = testData5[361];
@(posedge clk);
#1;data_in = testData5[362];
@(posedge clk);
#1;data_in = testData5[363];
@(posedge clk);
#1;data_in = testData5[364];
@(posedge clk);
#1;data_in = testData5[365];
@(posedge clk);
#1;data_in = testData5[366];
@(posedge clk);
#1;data_in = testData5[367];
@(posedge clk);
#1;data_in = testData5[368];
@(posedge clk);
#1;data_in = testData5[369];
@(posedge clk);
#1;data_in = testData5[370];
@(posedge clk);
#1;data_in = testData5[371];
@(posedge clk);
#1;data_in = testData5[372];
@(posedge clk);
#1;data_in = testData5[373];
@(posedge clk);
#1;data_in = testData5[374];
@(posedge clk);
#1;data_in = testData5[375];
@(posedge clk);
#1;data_in = testData5[376];
@(posedge clk);
#1;data_in = testData5[377];
@(posedge clk);
#1;data_in = testData5[378];
@(posedge clk);
#1;data_in = testData5[379];
@(posedge clk);
#1;data_in = testData5[380];
@(posedge clk);
#1;data_in = testData5[381];
@(posedge clk);
#1;data_in = testData5[382];
@(posedge clk);
#1;data_in = testData5[383];
@(posedge clk);
#1;data_in = testData5[384];
@(posedge clk);
#1;data_in = testData5[385];
@(posedge clk);
#1;data_in = testData5[386];
@(posedge clk);
#1;data_in = testData5[387];
@(posedge clk);
#1;data_in = testData5[388];
@(posedge clk);
#1;data_in = testData5[389];
@(posedge clk);
#1;data_in = testData5[390];
@(posedge clk);
#1;data_in = testData5[391];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[392]; 
@(posedge clk);
#1;data_in = testData5[393];
@(posedge clk);
#1;data_in = testData5[394];
@(posedge clk);
#1;data_in = testData5[395];
@(posedge clk);
#1;data_in = testData5[396];
@(posedge clk);
#1;data_in = testData5[397];
@(posedge clk);
#1;data_in = testData5[398];
@(posedge clk);
#1;data_in = testData5[399];
@(posedge clk);
#1;data_in = testData5[400];
@(posedge clk);
#1;data_in = testData5[401];
@(posedge clk);
#1;data_in = testData5[402];
@(posedge clk);
#1;data_in = testData5[403];
@(posedge clk);
#1;data_in = testData5[404];
@(posedge clk);
#1;data_in = testData5[405];
@(posedge clk);
#1;data_in = testData5[406];
@(posedge clk);
#1;data_in = testData5[407];
@(posedge clk);
#1;data_in = testData5[408];
@(posedge clk);
#1;data_in = testData5[409];
@(posedge clk);
#1;data_in = testData5[410];
@(posedge clk);
#1;data_in = testData5[411];
@(posedge clk);
#1;data_in = testData5[412];
@(posedge clk);
#1;data_in = testData5[413];
@(posedge clk);
#1;data_in = testData5[414];
@(posedge clk);
#1;data_in = testData5[415];
@(posedge clk);
#1;data_in = testData5[416];
@(posedge clk);
#1;data_in = testData5[417];
@(posedge clk);
#1;data_in = testData5[418];
@(posedge clk);
#1;data_in = testData5[419];
@(posedge clk);
#1;data_in = testData5[420];
@(posedge clk);
#1;data_in = testData5[421];
@(posedge clk);
#1;data_in = testData5[422];
@(posedge clk);
#1;data_in = testData5[423];
@(posedge clk);
#1;data_in = testData5[424];
@(posedge clk);
#1;data_in = testData5[425];
@(posedge clk);
#1;data_in = testData5[426];
@(posedge clk);
#1;data_in = testData5[427];
@(posedge clk);
#1;data_in = testData5[428];
@(posedge clk);
#1;data_in = testData5[429];
@(posedge clk);
#1;data_in = testData5[430];
@(posedge clk);
#1;data_in = testData5[431];
@(posedge clk);
#1;data_in = testData5[432];
@(posedge clk);
#1;data_in = testData5[433];
@(posedge clk);
#1;data_in = testData5[434];
@(posedge clk);
#1;data_in = testData5[435];
@(posedge clk);
#1;data_in = testData5[436];
@(posedge clk);
#1;data_in = testData5[437];
@(posedge clk);
#1;data_in = testData5[438];
@(posedge clk);
#1;data_in = testData5[439];
@(posedge clk);
#1;data_in = testData5[440];
@(posedge clk);
#1;data_in = testData5[441];
@(posedge clk);
#1;data_in = testData5[442];
@(posedge clk);
#1;data_in = testData5[443];
@(posedge clk);
#1;data_in = testData5[444];
@(posedge clk);
#1;data_in = testData5[445];
@(posedge clk);
#1;data_in = testData5[446];
@(posedge clk);
#1;data_in = testData5[447];
@(posedge clk);
#1;data_in = testData5[448];
@(posedge clk);
#1;data_in = testData5[449];
@(posedge clk);
#1;data_in = testData5[450];
@(posedge clk);
#1;data_in = testData5[451];
@(posedge clk);
#1;data_in = testData5[452];
@(posedge clk);
#1;data_in = testData5[453];
@(posedge clk);
#1;data_in = testData5[454];
@(posedge clk);
#1;data_in = testData5[455];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[456]; 
@(posedge clk);
#1;data_in = testData5[457];
@(posedge clk);
#1;data_in = testData5[458];
@(posedge clk);
#1;data_in = testData5[459];
@(posedge clk);
#1;data_in = testData5[460];
@(posedge clk);
#1;data_in = testData5[461];
@(posedge clk);
#1;data_in = testData5[462];
@(posedge clk);
#1;data_in = testData5[463];
@(posedge clk);
#1;data_in = testData5[464];
@(posedge clk);
#1;data_in = testData5[465];
@(posedge clk);
#1;data_in = testData5[466];
@(posedge clk);
#1;data_in = testData5[467];
@(posedge clk);
#1;data_in = testData5[468];
@(posedge clk);
#1;data_in = testData5[469];
@(posedge clk);
#1;data_in = testData5[470];
@(posedge clk);
#1;data_in = testData5[471];
@(posedge clk);
#1;data_in = testData5[472];
@(posedge clk);
#1;data_in = testData5[473];
@(posedge clk);
#1;data_in = testData5[474];
@(posedge clk);
#1;data_in = testData5[475];
@(posedge clk);
#1;data_in = testData5[476];
@(posedge clk);
#1;data_in = testData5[477];
@(posedge clk);
#1;data_in = testData5[478];
@(posedge clk);
#1;data_in = testData5[479];
@(posedge clk);
#1;data_in = testData5[480];
@(posedge clk);
#1;data_in = testData5[481];
@(posedge clk);
#1;data_in = testData5[482];
@(posedge clk);
#1;data_in = testData5[483];
@(posedge clk);
#1;data_in = testData5[484];
@(posedge clk);
#1;data_in = testData5[485];
@(posedge clk);
#1;data_in = testData5[486];
@(posedge clk);
#1;data_in = testData5[487];
@(posedge clk);
#1;data_in = testData5[488];
@(posedge clk);
#1;data_in = testData5[489];
@(posedge clk);
#1;data_in = testData5[490];
@(posedge clk);
#1;data_in = testData5[491];
@(posedge clk);
#1;data_in = testData5[492];
@(posedge clk);
#1;data_in = testData5[493];
@(posedge clk);
#1;data_in = testData5[494];
@(posedge clk);
#1;data_in = testData5[495];
@(posedge clk);
#1;data_in = testData5[496];
@(posedge clk);
#1;data_in = testData5[497];
@(posedge clk);
#1;data_in = testData5[498];
@(posedge clk);
#1;data_in = testData5[499];
@(posedge clk);
#1;data_in = testData5[500];
@(posedge clk);
#1;data_in = testData5[501];
@(posedge clk);
#1;data_in = testData5[502];
@(posedge clk);
#1;data_in = testData5[503];
@(posedge clk);
#1;data_in = testData5[504];
@(posedge clk);
#1;data_in = testData5[505];
@(posedge clk);
#1;data_in = testData5[506];
@(posedge clk);
#1;data_in = testData5[507];
@(posedge clk);
#1;data_in = testData5[508];
@(posedge clk);
#1;data_in = testData5[509];
@(posedge clk);
#1;data_in = testData5[510];
@(posedge clk);
#1;data_in = testData5[511];
@(posedge clk);
#1;data_in = testData5[512];
@(posedge clk);
#1;data_in = testData5[513];
@(posedge clk);
#1;data_in = testData5[514];
@(posedge clk);
#1;data_in = testData5[515];
@(posedge clk);
#1;data_in = testData5[516];
@(posedge clk);
#1;data_in = testData5[517];
@(posedge clk);
#1;data_in = testData5[518];
@(posedge clk);
#1;data_in = testData5[519];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[520]; 
@(posedge clk);
#1;data_in = testData5[521];
@(posedge clk);
#1;data_in = testData5[522];
@(posedge clk);
#1;data_in = testData5[523];
@(posedge clk);
#1;data_in = testData5[524];
@(posedge clk);
#1;data_in = testData5[525];
@(posedge clk);
#1;data_in = testData5[526];
@(posedge clk);
#1;data_in = testData5[527];
@(posedge clk);
#1;data_in = testData5[528];
@(posedge clk);
#1;data_in = testData5[529];
@(posedge clk);
#1;data_in = testData5[530];
@(posedge clk);
#1;data_in = testData5[531];
@(posedge clk);
#1;data_in = testData5[532];
@(posedge clk);
#1;data_in = testData5[533];
@(posedge clk);
#1;data_in = testData5[534];
@(posedge clk);
#1;data_in = testData5[535];
@(posedge clk);
#1;data_in = testData5[536];
@(posedge clk);
#1;data_in = testData5[537];
@(posedge clk);
#1;data_in = testData5[538];
@(posedge clk);
#1;data_in = testData5[539];
@(posedge clk);
#1;data_in = testData5[540];
@(posedge clk);
#1;data_in = testData5[541];
@(posedge clk);
#1;data_in = testData5[542];
@(posedge clk);
#1;data_in = testData5[543];
@(posedge clk);
#1;data_in = testData5[544];
@(posedge clk);
#1;data_in = testData5[545];
@(posedge clk);
#1;data_in = testData5[546];
@(posedge clk);
#1;data_in = testData5[547];
@(posedge clk);
#1;data_in = testData5[548];
@(posedge clk);
#1;data_in = testData5[549];
@(posedge clk);
#1;data_in = testData5[550];
@(posedge clk);
#1;data_in = testData5[551];
@(posedge clk);
#1;data_in = testData5[552];
@(posedge clk);
#1;data_in = testData5[553];
@(posedge clk);
#1;data_in = testData5[554];
@(posedge clk);
#1;data_in = testData5[555];
@(posedge clk);
#1;data_in = testData5[556];
@(posedge clk);
#1;data_in = testData5[557];
@(posedge clk);
#1;data_in = testData5[558];
@(posedge clk);
#1;data_in = testData5[559];
@(posedge clk);
#1;data_in = testData5[560];
@(posedge clk);
#1;data_in = testData5[561];
@(posedge clk);
#1;data_in = testData5[562];
@(posedge clk);
#1;data_in = testData5[563];
@(posedge clk);
#1;data_in = testData5[564];
@(posedge clk);
#1;data_in = testData5[565];
@(posedge clk);
#1;data_in = testData5[566];
@(posedge clk);
#1;data_in = testData5[567];
@(posedge clk);
#1;data_in = testData5[568];
@(posedge clk);
#1;data_in = testData5[569];
@(posedge clk);
#1;data_in = testData5[570];
@(posedge clk);
#1;data_in = testData5[571];
@(posedge clk);
#1;data_in = testData5[572];
@(posedge clk);
#1;data_in = testData5[573];
@(posedge clk);
#1;data_in = testData5[574];
@(posedge clk);
#1;data_in = testData5[575];
@(posedge clk);
#1;data_in = testData5[576];
@(posedge clk);
#1;data_in = testData5[577];
@(posedge clk);
#1;data_in = testData5[578];
@(posedge clk);
#1;data_in = testData5[579];
@(posedge clk);
#1;data_in = testData5[580];
@(posedge clk);
#1;data_in = testData5[581];
@(posedge clk);
#1;data_in = testData5[582];
@(posedge clk);
#1;data_in = testData5[583];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[584]; 
@(posedge clk);
#1;data_in = testData5[585];
@(posedge clk);
#1;data_in = testData5[586];
@(posedge clk);
#1;data_in = testData5[587];
@(posedge clk);
#1;data_in = testData5[588];
@(posedge clk);
#1;data_in = testData5[589];
@(posedge clk);
#1;data_in = testData5[590];
@(posedge clk);
#1;data_in = testData5[591];
@(posedge clk);
#1;data_in = testData5[592];
@(posedge clk);
#1;data_in = testData5[593];
@(posedge clk);
#1;data_in = testData5[594];
@(posedge clk);
#1;data_in = testData5[595];
@(posedge clk);
#1;data_in = testData5[596];
@(posedge clk);
#1;data_in = testData5[597];
@(posedge clk);
#1;data_in = testData5[598];
@(posedge clk);
#1;data_in = testData5[599];
@(posedge clk);
#1;data_in = testData5[600];
@(posedge clk);
#1;data_in = testData5[601];
@(posedge clk);
#1;data_in = testData5[602];
@(posedge clk);
#1;data_in = testData5[603];
@(posedge clk);
#1;data_in = testData5[604];
@(posedge clk);
#1;data_in = testData5[605];
@(posedge clk);
#1;data_in = testData5[606];
@(posedge clk);
#1;data_in = testData5[607];
@(posedge clk);
#1;data_in = testData5[608];
@(posedge clk);
#1;data_in = testData5[609];
@(posedge clk);
#1;data_in = testData5[610];
@(posedge clk);
#1;data_in = testData5[611];
@(posedge clk);
#1;data_in = testData5[612];
@(posedge clk);
#1;data_in = testData5[613];
@(posedge clk);
#1;data_in = testData5[614];
@(posedge clk);
#1;data_in = testData5[615];
@(posedge clk);
#1;data_in = testData5[616];
@(posedge clk);
#1;data_in = testData5[617];
@(posedge clk);
#1;data_in = testData5[618];
@(posedge clk);
#1;data_in = testData5[619];
@(posedge clk);
#1;data_in = testData5[620];
@(posedge clk);
#1;data_in = testData5[621];
@(posedge clk);
#1;data_in = testData5[622];
@(posedge clk);
#1;data_in = testData5[623];
@(posedge clk);
#1;data_in = testData5[624];
@(posedge clk);
#1;data_in = testData5[625];
@(posedge clk);
#1;data_in = testData5[626];
@(posedge clk);
#1;data_in = testData5[627];
@(posedge clk);
#1;data_in = testData5[628];
@(posedge clk);
#1;data_in = testData5[629];
@(posedge clk);
#1;data_in = testData5[630];
@(posedge clk);
#1;data_in = testData5[631];
@(posedge clk);
#1;data_in = testData5[632];
@(posedge clk);
#1;data_in = testData5[633];
@(posedge clk);
#1;data_in = testData5[634];
@(posedge clk);
#1;data_in = testData5[635];
@(posedge clk);
#1;data_in = testData5[636];
@(posedge clk);
#1;data_in = testData5[637];
@(posedge clk);
#1;data_in = testData5[638];
@(posedge clk);
#1;data_in = testData5[639];
@(posedge clk);
#1;data_in = testData5[640];
@(posedge clk);
#1;data_in = testData5[641];
@(posedge clk);
#1;data_in = testData5[642];
@(posedge clk);
#1;data_in = testData5[643];
@(posedge clk);
#1;data_in = testData5[644];
@(posedge clk);
#1;data_in = testData5[645];
@(posedge clk);
#1;data_in = testData5[646];
@(posedge clk);
#1;data_in = testData5[647];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[648]; 
@(posedge clk);
#1;data_in = testData5[649];
@(posedge clk);
#1;data_in = testData5[650];
@(posedge clk);
#1;data_in = testData5[651];
@(posedge clk);
#1;data_in = testData5[652];
@(posedge clk);
#1;data_in = testData5[653];
@(posedge clk);
#1;data_in = testData5[654];
@(posedge clk);
#1;data_in = testData5[655];
@(posedge clk);
#1;data_in = testData5[656];
@(posedge clk);
#1;data_in = testData5[657];
@(posedge clk);
#1;data_in = testData5[658];
@(posedge clk);
#1;data_in = testData5[659];
@(posedge clk);
#1;data_in = testData5[660];
@(posedge clk);
#1;data_in = testData5[661];
@(posedge clk);
#1;data_in = testData5[662];
@(posedge clk);
#1;data_in = testData5[663];
@(posedge clk);
#1;data_in = testData5[664];
@(posedge clk);
#1;data_in = testData5[665];
@(posedge clk);
#1;data_in = testData5[666];
@(posedge clk);
#1;data_in = testData5[667];
@(posedge clk);
#1;data_in = testData5[668];
@(posedge clk);
#1;data_in = testData5[669];
@(posedge clk);
#1;data_in = testData5[670];
@(posedge clk);
#1;data_in = testData5[671];
@(posedge clk);
#1;data_in = testData5[672];
@(posedge clk);
#1;data_in = testData5[673];
@(posedge clk);
#1;data_in = testData5[674];
@(posedge clk);
#1;data_in = testData5[675];
@(posedge clk);
#1;data_in = testData5[676];
@(posedge clk);
#1;data_in = testData5[677];
@(posedge clk);
#1;data_in = testData5[678];
@(posedge clk);
#1;data_in = testData5[679];
@(posedge clk);
#1;data_in = testData5[680];
@(posedge clk);
#1;data_in = testData5[681];
@(posedge clk);
#1;data_in = testData5[682];
@(posedge clk);
#1;data_in = testData5[683];
@(posedge clk);
#1;data_in = testData5[684];
@(posedge clk);
#1;data_in = testData5[685];
@(posedge clk);
#1;data_in = testData5[686];
@(posedge clk);
#1;data_in = testData5[687];
@(posedge clk);
#1;data_in = testData5[688];
@(posedge clk);
#1;data_in = testData5[689];
@(posedge clk);
#1;data_in = testData5[690];
@(posedge clk);
#1;data_in = testData5[691];
@(posedge clk);
#1;data_in = testData5[692];
@(posedge clk);
#1;data_in = testData5[693];
@(posedge clk);
#1;data_in = testData5[694];
@(posedge clk);
#1;data_in = testData5[695];
@(posedge clk);
#1;data_in = testData5[696];
@(posedge clk);
#1;data_in = testData5[697];
@(posedge clk);
#1;data_in = testData5[698];
@(posedge clk);
#1;data_in = testData5[699];
@(posedge clk);
#1;data_in = testData5[700];
@(posedge clk);
#1;data_in = testData5[701];
@(posedge clk);
#1;data_in = testData5[702];
@(posedge clk);
#1;data_in = testData5[703];
@(posedge clk);
#1;data_in = testData5[704];
@(posedge clk);
#1;data_in = testData5[705];
@(posedge clk);
#1;data_in = testData5[706];
@(posedge clk);
#1;data_in = testData5[707];
@(posedge clk);
#1;data_in = testData5[708];
@(posedge clk);
#1;data_in = testData5[709];
@(posedge clk);
#1;data_in = testData5[710];
@(posedge clk);
#1;data_in = testData5[711];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[712]; 
@(posedge clk);
#1;data_in = testData5[713];
@(posedge clk);
#1;data_in = testData5[714];
@(posedge clk);
#1;data_in = testData5[715];
@(posedge clk);
#1;data_in = testData5[716];
@(posedge clk);
#1;data_in = testData5[717];
@(posedge clk);
#1;data_in = testData5[718];
@(posedge clk);
#1;data_in = testData5[719];
@(posedge clk);
#1;data_in = testData5[720];
@(posedge clk);
#1;data_in = testData5[721];
@(posedge clk);
#1;data_in = testData5[722];
@(posedge clk);
#1;data_in = testData5[723];
@(posedge clk);
#1;data_in = testData5[724];
@(posedge clk);
#1;data_in = testData5[725];
@(posedge clk);
#1;data_in = testData5[726];
@(posedge clk);
#1;data_in = testData5[727];
@(posedge clk);
#1;data_in = testData5[728];
@(posedge clk);
#1;data_in = testData5[729];
@(posedge clk);
#1;data_in = testData5[730];
@(posedge clk);
#1;data_in = testData5[731];
@(posedge clk);
#1;data_in = testData5[732];
@(posedge clk);
#1;data_in = testData5[733];
@(posedge clk);
#1;data_in = testData5[734];
@(posedge clk);
#1;data_in = testData5[735];
@(posedge clk);
#1;data_in = testData5[736];
@(posedge clk);
#1;data_in = testData5[737];
@(posedge clk);
#1;data_in = testData5[738];
@(posedge clk);
#1;data_in = testData5[739];
@(posedge clk);
#1;data_in = testData5[740];
@(posedge clk);
#1;data_in = testData5[741];
@(posedge clk);
#1;data_in = testData5[742];
@(posedge clk);
#1;data_in = testData5[743];
@(posedge clk);
#1;data_in = testData5[744];
@(posedge clk);
#1;data_in = testData5[745];
@(posedge clk);
#1;data_in = testData5[746];
@(posedge clk);
#1;data_in = testData5[747];
@(posedge clk);
#1;data_in = testData5[748];
@(posedge clk);
#1;data_in = testData5[749];
@(posedge clk);
#1;data_in = testData5[750];
@(posedge clk);
#1;data_in = testData5[751];
@(posedge clk);
#1;data_in = testData5[752];
@(posedge clk);
#1;data_in = testData5[753];
@(posedge clk);
#1;data_in = testData5[754];
@(posedge clk);
#1;data_in = testData5[755];
@(posedge clk);
#1;data_in = testData5[756];
@(posedge clk);
#1;data_in = testData5[757];
@(posedge clk);
#1;data_in = testData5[758];
@(posedge clk);
#1;data_in = testData5[759];
@(posedge clk);
#1;data_in = testData5[760];
@(posedge clk);
#1;data_in = testData5[761];
@(posedge clk);
#1;data_in = testData5[762];
@(posedge clk);
#1;data_in = testData5[763];
@(posedge clk);
#1;data_in = testData5[764];
@(posedge clk);
#1;data_in = testData5[765];
@(posedge clk);
#1;data_in = testData5[766];
@(posedge clk);
#1;data_in = testData5[767];
@(posedge clk);
#1;data_in = testData5[768];
@(posedge clk);
#1;data_in = testData5[769];
@(posedge clk);
#1;data_in = testData5[770];
@(posedge clk);
#1;data_in = testData5[771];
@(posedge clk);
#1;data_in = testData5[772];
@(posedge clk);
#1;data_in = testData5[773];
@(posedge clk);
#1;data_in = testData5[774];
@(posedge clk);
#1;data_in = testData5[775];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[776]; 
@(posedge clk);
#1;data_in = testData5[777];
@(posedge clk);
#1;data_in = testData5[778];
@(posedge clk);
#1;data_in = testData5[779];
@(posedge clk);
#1;data_in = testData5[780];
@(posedge clk);
#1;data_in = testData5[781];
@(posedge clk);
#1;data_in = testData5[782];
@(posedge clk);
#1;data_in = testData5[783];
@(posedge clk);
#1;data_in = testData5[784];
@(posedge clk);
#1;data_in = testData5[785];
@(posedge clk);
#1;data_in = testData5[786];
@(posedge clk);
#1;data_in = testData5[787];
@(posedge clk);
#1;data_in = testData5[788];
@(posedge clk);
#1;data_in = testData5[789];
@(posedge clk);
#1;data_in = testData5[790];
@(posedge clk);
#1;data_in = testData5[791];
@(posedge clk);
#1;data_in = testData5[792];
@(posedge clk);
#1;data_in = testData5[793];
@(posedge clk);
#1;data_in = testData5[794];
@(posedge clk);
#1;data_in = testData5[795];
@(posedge clk);
#1;data_in = testData5[796];
@(posedge clk);
#1;data_in = testData5[797];
@(posedge clk);
#1;data_in = testData5[798];
@(posedge clk);
#1;data_in = testData5[799];
@(posedge clk);
#1;data_in = testData5[800];
@(posedge clk);
#1;data_in = testData5[801];
@(posedge clk);
#1;data_in = testData5[802];
@(posedge clk);
#1;data_in = testData5[803];
@(posedge clk);
#1;data_in = testData5[804];
@(posedge clk);
#1;data_in = testData5[805];
@(posedge clk);
#1;data_in = testData5[806];
@(posedge clk);
#1;data_in = testData5[807];
@(posedge clk);
#1;data_in = testData5[808];
@(posedge clk);
#1;data_in = testData5[809];
@(posedge clk);
#1;data_in = testData5[810];
@(posedge clk);
#1;data_in = testData5[811];
@(posedge clk);
#1;data_in = testData5[812];
@(posedge clk);
#1;data_in = testData5[813];
@(posedge clk);
#1;data_in = testData5[814];
@(posedge clk);
#1;data_in = testData5[815];
@(posedge clk);
#1;data_in = testData5[816];
@(posedge clk);
#1;data_in = testData5[817];
@(posedge clk);
#1;data_in = testData5[818];
@(posedge clk);
#1;data_in = testData5[819];
@(posedge clk);
#1;data_in = testData5[820];
@(posedge clk);
#1;data_in = testData5[821];
@(posedge clk);
#1;data_in = testData5[822];
@(posedge clk);
#1;data_in = testData5[823];
@(posedge clk);
#1;data_in = testData5[824];
@(posedge clk);
#1;data_in = testData5[825];
@(posedge clk);
#1;data_in = testData5[826];
@(posedge clk);
#1;data_in = testData5[827];
@(posedge clk);
#1;data_in = testData5[828];
@(posedge clk);
#1;data_in = testData5[829];
@(posedge clk);
#1;data_in = testData5[830];
@(posedge clk);
#1;data_in = testData5[831];
@(posedge clk);
#1;data_in = testData5[832];
@(posedge clk);
#1;data_in = testData5[833];
@(posedge clk);
#1;data_in = testData5[834];
@(posedge clk);
#1;data_in = testData5[835];
@(posedge clk);
#1;data_in = testData5[836];
@(posedge clk);
#1;data_in = testData5[837];
@(posedge clk);
#1;data_in = testData5[838];
@(posedge clk);
#1;data_in = testData5[839];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[840]; 
@(posedge clk);
#1;data_in = testData5[841];
@(posedge clk);
#1;data_in = testData5[842];
@(posedge clk);
#1;data_in = testData5[843];
@(posedge clk);
#1;data_in = testData5[844];
@(posedge clk);
#1;data_in = testData5[845];
@(posedge clk);
#1;data_in = testData5[846];
@(posedge clk);
#1;data_in = testData5[847];
@(posedge clk);
#1;data_in = testData5[848];
@(posedge clk);
#1;data_in = testData5[849];
@(posedge clk);
#1;data_in = testData5[850];
@(posedge clk);
#1;data_in = testData5[851];
@(posedge clk);
#1;data_in = testData5[852];
@(posedge clk);
#1;data_in = testData5[853];
@(posedge clk);
#1;data_in = testData5[854];
@(posedge clk);
#1;data_in = testData5[855];
@(posedge clk);
#1;data_in = testData5[856];
@(posedge clk);
#1;data_in = testData5[857];
@(posedge clk);
#1;data_in = testData5[858];
@(posedge clk);
#1;data_in = testData5[859];
@(posedge clk);
#1;data_in = testData5[860];
@(posedge clk);
#1;data_in = testData5[861];
@(posedge clk);
#1;data_in = testData5[862];
@(posedge clk);
#1;data_in = testData5[863];
@(posedge clk);
#1;data_in = testData5[864];
@(posedge clk);
#1;data_in = testData5[865];
@(posedge clk);
#1;data_in = testData5[866];
@(posedge clk);
#1;data_in = testData5[867];
@(posedge clk);
#1;data_in = testData5[868];
@(posedge clk);
#1;data_in = testData5[869];
@(posedge clk);
#1;data_in = testData5[870];
@(posedge clk);
#1;data_in = testData5[871];
@(posedge clk);
#1;data_in = testData5[872];
@(posedge clk);
#1;data_in = testData5[873];
@(posedge clk);
#1;data_in = testData5[874];
@(posedge clk);
#1;data_in = testData5[875];
@(posedge clk);
#1;data_in = testData5[876];
@(posedge clk);
#1;data_in = testData5[877];
@(posedge clk);
#1;data_in = testData5[878];
@(posedge clk);
#1;data_in = testData5[879];
@(posedge clk);
#1;data_in = testData5[880];
@(posedge clk);
#1;data_in = testData5[881];
@(posedge clk);
#1;data_in = testData5[882];
@(posedge clk);
#1;data_in = testData5[883];
@(posedge clk);
#1;data_in = testData5[884];
@(posedge clk);
#1;data_in = testData5[885];
@(posedge clk);
#1;data_in = testData5[886];
@(posedge clk);
#1;data_in = testData5[887];
@(posedge clk);
#1;data_in = testData5[888];
@(posedge clk);
#1;data_in = testData5[889];
@(posedge clk);
#1;data_in = testData5[890];
@(posedge clk);
#1;data_in = testData5[891];
@(posedge clk);
#1;data_in = testData5[892];
@(posedge clk);
#1;data_in = testData5[893];
@(posedge clk);
#1;data_in = testData5[894];
@(posedge clk);
#1;data_in = testData5[895];
@(posedge clk);
#1;data_in = testData5[896];
@(posedge clk);
#1;data_in = testData5[897];
@(posedge clk);
#1;data_in = testData5[898];
@(posedge clk);
#1;data_in = testData5[899];
@(posedge clk);
#1;data_in = testData5[900];
@(posedge clk);
#1;data_in = testData5[901];
@(posedge clk);
#1;data_in = testData5[902];
@(posedge clk);
#1;data_in = testData5[903];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[904]; 
@(posedge clk);
#1;data_in = testData5[905];
@(posedge clk);
#1;data_in = testData5[906];
@(posedge clk);
#1;data_in = testData5[907];
@(posedge clk);
#1;data_in = testData5[908];
@(posedge clk);
#1;data_in = testData5[909];
@(posedge clk);
#1;data_in = testData5[910];
@(posedge clk);
#1;data_in = testData5[911];
@(posedge clk);
#1;data_in = testData5[912];
@(posedge clk);
#1;data_in = testData5[913];
@(posedge clk);
#1;data_in = testData5[914];
@(posedge clk);
#1;data_in = testData5[915];
@(posedge clk);
#1;data_in = testData5[916];
@(posedge clk);
#1;data_in = testData5[917];
@(posedge clk);
#1;data_in = testData5[918];
@(posedge clk);
#1;data_in = testData5[919];
@(posedge clk);
#1;data_in = testData5[920];
@(posedge clk);
#1;data_in = testData5[921];
@(posedge clk);
#1;data_in = testData5[922];
@(posedge clk);
#1;data_in = testData5[923];
@(posedge clk);
#1;data_in = testData5[924];
@(posedge clk);
#1;data_in = testData5[925];
@(posedge clk);
#1;data_in = testData5[926];
@(posedge clk);
#1;data_in = testData5[927];
@(posedge clk);
#1;data_in = testData5[928];
@(posedge clk);
#1;data_in = testData5[929];
@(posedge clk);
#1;data_in = testData5[930];
@(posedge clk);
#1;data_in = testData5[931];
@(posedge clk);
#1;data_in = testData5[932];
@(posedge clk);
#1;data_in = testData5[933];
@(posedge clk);
#1;data_in = testData5[934];
@(posedge clk);
#1;data_in = testData5[935];
@(posedge clk);
#1;data_in = testData5[936];
@(posedge clk);
#1;data_in = testData5[937];
@(posedge clk);
#1;data_in = testData5[938];
@(posedge clk);
#1;data_in = testData5[939];
@(posedge clk);
#1;data_in = testData5[940];
@(posedge clk);
#1;data_in = testData5[941];
@(posedge clk);
#1;data_in = testData5[942];
@(posedge clk);
#1;data_in = testData5[943];
@(posedge clk);
#1;data_in = testData5[944];
@(posedge clk);
#1;data_in = testData5[945];
@(posedge clk);
#1;data_in = testData5[946];
@(posedge clk);
#1;data_in = testData5[947];
@(posedge clk);
#1;data_in = testData5[948];
@(posedge clk);
#1;data_in = testData5[949];
@(posedge clk);
#1;data_in = testData5[950];
@(posedge clk);
#1;data_in = testData5[951];
@(posedge clk);
#1;data_in = testData5[952];
@(posedge clk);
#1;data_in = testData5[953];
@(posedge clk);
#1;data_in = testData5[954];
@(posedge clk);
#1;data_in = testData5[955];
@(posedge clk);
#1;data_in = testData5[956];
@(posedge clk);
#1;data_in = testData5[957];
@(posedge clk);
#1;data_in = testData5[958];
@(posedge clk);
#1;data_in = testData5[959];
@(posedge clk);
#1;data_in = testData5[960];
@(posedge clk);
#1;data_in = testData5[961];
@(posedge clk);
#1;data_in = testData5[962];
@(posedge clk);
#1;data_in = testData5[963];
@(posedge clk);
#1;data_in = testData5[964];
@(posedge clk);
#1;data_in = testData5[965];
@(posedge clk);
#1;data_in = testData5[966];
@(posedge clk);
#1;data_in = testData5[967];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[968]; 
@(posedge clk);
#1;data_in = testData5[969];
@(posedge clk);
#1;data_in = testData5[970];
@(posedge clk);
#1;data_in = testData5[971];
@(posedge clk);
#1;data_in = testData5[972];
@(posedge clk);
#1;data_in = testData5[973];
@(posedge clk);
#1;data_in = testData5[974];
@(posedge clk);
#1;data_in = testData5[975];
@(posedge clk);
#1;data_in = testData5[976];
@(posedge clk);
#1;data_in = testData5[977];
@(posedge clk);
#1;data_in = testData5[978];
@(posedge clk);
#1;data_in = testData5[979];
@(posedge clk);
#1;data_in = testData5[980];
@(posedge clk);
#1;data_in = testData5[981];
@(posedge clk);
#1;data_in = testData5[982];
@(posedge clk);
#1;data_in = testData5[983];
@(posedge clk);
#1;data_in = testData5[984];
@(posedge clk);
#1;data_in = testData5[985];
@(posedge clk);
#1;data_in = testData5[986];
@(posedge clk);
#1;data_in = testData5[987];
@(posedge clk);
#1;data_in = testData5[988];
@(posedge clk);
#1;data_in = testData5[989];
@(posedge clk);
#1;data_in = testData5[990];
@(posedge clk);
#1;data_in = testData5[991];
@(posedge clk);
#1;data_in = testData5[992];
@(posedge clk);
#1;data_in = testData5[993];
@(posedge clk);
#1;data_in = testData5[994];
@(posedge clk);
#1;data_in = testData5[995];
@(posedge clk);
#1;data_in = testData5[996];
@(posedge clk);
#1;data_in = testData5[997];
@(posedge clk);
#1;data_in = testData5[998];
@(posedge clk);
#1;data_in = testData5[999];
@(posedge clk);
#1;data_in = testData5[1000];
@(posedge clk);
#1;data_in = testData5[1001];
@(posedge clk);
#1;data_in = testData5[1002];
@(posedge clk);
#1;data_in = testData5[1003];
@(posedge clk);
#1;data_in = testData5[1004];
@(posedge clk);
#1;data_in = testData5[1005];
@(posedge clk);
#1;data_in = testData5[1006];
@(posedge clk);
#1;data_in = testData5[1007];
@(posedge clk);
#1;data_in = testData5[1008];
@(posedge clk);
#1;data_in = testData5[1009];
@(posedge clk);
#1;data_in = testData5[1010];
@(posedge clk);
#1;data_in = testData5[1011];
@(posedge clk);
#1;data_in = testData5[1012];
@(posedge clk);
#1;data_in = testData5[1013];
@(posedge clk);
#1;data_in = testData5[1014];
@(posedge clk);
#1;data_in = testData5[1015];
@(posedge clk);
#1;data_in = testData5[1016];
@(posedge clk);
#1;data_in = testData5[1017];
@(posedge clk);
#1;data_in = testData5[1018];
@(posedge clk);
#1;data_in = testData5[1019];
@(posedge clk);
#1;data_in = testData5[1020];
@(posedge clk);
#1;data_in = testData5[1021];
@(posedge clk);
#1;data_in = testData5[1022];
@(posedge clk);
#1;data_in = testData5[1023];
@(posedge clk);
#1;data_in = testData5[1024];
@(posedge clk);
#1;data_in = testData5[1025];
@(posedge clk);
#1;data_in = testData5[1026];
@(posedge clk);
#1;data_in = testData5[1027];
@(posedge clk);
#1;data_in = testData5[1028];
@(posedge clk);
#1;data_in = testData5[1029];
@(posedge clk);
#1;data_in = testData5[1030];
@(posedge clk);
#1;data_in = testData5[1031];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1032]; 
@(posedge clk);
#1;data_in = testData5[1033];
@(posedge clk);
#1;data_in = testData5[1034];
@(posedge clk);
#1;data_in = testData5[1035];
@(posedge clk);
#1;data_in = testData5[1036];
@(posedge clk);
#1;data_in = testData5[1037];
@(posedge clk);
#1;data_in = testData5[1038];
@(posedge clk);
#1;data_in = testData5[1039];
@(posedge clk);
#1;data_in = testData5[1040];
@(posedge clk);
#1;data_in = testData5[1041];
@(posedge clk);
#1;data_in = testData5[1042];
@(posedge clk);
#1;data_in = testData5[1043];
@(posedge clk);
#1;data_in = testData5[1044];
@(posedge clk);
#1;data_in = testData5[1045];
@(posedge clk);
#1;data_in = testData5[1046];
@(posedge clk);
#1;data_in = testData5[1047];
@(posedge clk);
#1;data_in = testData5[1048];
@(posedge clk);
#1;data_in = testData5[1049];
@(posedge clk);
#1;data_in = testData5[1050];
@(posedge clk);
#1;data_in = testData5[1051];
@(posedge clk);
#1;data_in = testData5[1052];
@(posedge clk);
#1;data_in = testData5[1053];
@(posedge clk);
#1;data_in = testData5[1054];
@(posedge clk);
#1;data_in = testData5[1055];
@(posedge clk);
#1;data_in = testData5[1056];
@(posedge clk);
#1;data_in = testData5[1057];
@(posedge clk);
#1;data_in = testData5[1058];
@(posedge clk);
#1;data_in = testData5[1059];
@(posedge clk);
#1;data_in = testData5[1060];
@(posedge clk);
#1;data_in = testData5[1061];
@(posedge clk);
#1;data_in = testData5[1062];
@(posedge clk);
#1;data_in = testData5[1063];
@(posedge clk);
#1;data_in = testData5[1064];
@(posedge clk);
#1;data_in = testData5[1065];
@(posedge clk);
#1;data_in = testData5[1066];
@(posedge clk);
#1;data_in = testData5[1067];
@(posedge clk);
#1;data_in = testData5[1068];
@(posedge clk);
#1;data_in = testData5[1069];
@(posedge clk);
#1;data_in = testData5[1070];
@(posedge clk);
#1;data_in = testData5[1071];
@(posedge clk);
#1;data_in = testData5[1072];
@(posedge clk);
#1;data_in = testData5[1073];
@(posedge clk);
#1;data_in = testData5[1074];
@(posedge clk);
#1;data_in = testData5[1075];
@(posedge clk);
#1;data_in = testData5[1076];
@(posedge clk);
#1;data_in = testData5[1077];
@(posedge clk);
#1;data_in = testData5[1078];
@(posedge clk);
#1;data_in = testData5[1079];
@(posedge clk);
#1;data_in = testData5[1080];
@(posedge clk);
#1;data_in = testData5[1081];
@(posedge clk);
#1;data_in = testData5[1082];
@(posedge clk);
#1;data_in = testData5[1083];
@(posedge clk);
#1;data_in = testData5[1084];
@(posedge clk);
#1;data_in = testData5[1085];
@(posedge clk);
#1;data_in = testData5[1086];
@(posedge clk);
#1;data_in = testData5[1087];
@(posedge clk);
#1;data_in = testData5[1088];
@(posedge clk);
#1;data_in = testData5[1089];
@(posedge clk);
#1;data_in = testData5[1090];
@(posedge clk);
#1;data_in = testData5[1091];
@(posedge clk);
#1;data_in = testData5[1092];
@(posedge clk);
#1;data_in = testData5[1093];
@(posedge clk);
#1;data_in = testData5[1094];
@(posedge clk);
#1;data_in = testData5[1095];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1096]; 
@(posedge clk);
#1;data_in = testData5[1097];
@(posedge clk);
#1;data_in = testData5[1098];
@(posedge clk);
#1;data_in = testData5[1099];
@(posedge clk);
#1;data_in = testData5[1100];
@(posedge clk);
#1;data_in = testData5[1101];
@(posedge clk);
#1;data_in = testData5[1102];
@(posedge clk);
#1;data_in = testData5[1103];
@(posedge clk);
#1;data_in = testData5[1104];
@(posedge clk);
#1;data_in = testData5[1105];
@(posedge clk);
#1;data_in = testData5[1106];
@(posedge clk);
#1;data_in = testData5[1107];
@(posedge clk);
#1;data_in = testData5[1108];
@(posedge clk);
#1;data_in = testData5[1109];
@(posedge clk);
#1;data_in = testData5[1110];
@(posedge clk);
#1;data_in = testData5[1111];
@(posedge clk);
#1;data_in = testData5[1112];
@(posedge clk);
#1;data_in = testData5[1113];
@(posedge clk);
#1;data_in = testData5[1114];
@(posedge clk);
#1;data_in = testData5[1115];
@(posedge clk);
#1;data_in = testData5[1116];
@(posedge clk);
#1;data_in = testData5[1117];
@(posedge clk);
#1;data_in = testData5[1118];
@(posedge clk);
#1;data_in = testData5[1119];
@(posedge clk);
#1;data_in = testData5[1120];
@(posedge clk);
#1;data_in = testData5[1121];
@(posedge clk);
#1;data_in = testData5[1122];
@(posedge clk);
#1;data_in = testData5[1123];
@(posedge clk);
#1;data_in = testData5[1124];
@(posedge clk);
#1;data_in = testData5[1125];
@(posedge clk);
#1;data_in = testData5[1126];
@(posedge clk);
#1;data_in = testData5[1127];
@(posedge clk);
#1;data_in = testData5[1128];
@(posedge clk);
#1;data_in = testData5[1129];
@(posedge clk);
#1;data_in = testData5[1130];
@(posedge clk);
#1;data_in = testData5[1131];
@(posedge clk);
#1;data_in = testData5[1132];
@(posedge clk);
#1;data_in = testData5[1133];
@(posedge clk);
#1;data_in = testData5[1134];
@(posedge clk);
#1;data_in = testData5[1135];
@(posedge clk);
#1;data_in = testData5[1136];
@(posedge clk);
#1;data_in = testData5[1137];
@(posedge clk);
#1;data_in = testData5[1138];
@(posedge clk);
#1;data_in = testData5[1139];
@(posedge clk);
#1;data_in = testData5[1140];
@(posedge clk);
#1;data_in = testData5[1141];
@(posedge clk);
#1;data_in = testData5[1142];
@(posedge clk);
#1;data_in = testData5[1143];
@(posedge clk);
#1;data_in = testData5[1144];
@(posedge clk);
#1;data_in = testData5[1145];
@(posedge clk);
#1;data_in = testData5[1146];
@(posedge clk);
#1;data_in = testData5[1147];
@(posedge clk);
#1;data_in = testData5[1148];
@(posedge clk);
#1;data_in = testData5[1149];
@(posedge clk);
#1;data_in = testData5[1150];
@(posedge clk);
#1;data_in = testData5[1151];
@(posedge clk);
#1;data_in = testData5[1152];
@(posedge clk);
#1;data_in = testData5[1153];
@(posedge clk);
#1;data_in = testData5[1154];
@(posedge clk);
#1;data_in = testData5[1155];
@(posedge clk);
#1;data_in = testData5[1156];
@(posedge clk);
#1;data_in = testData5[1157];
@(posedge clk);
#1;data_in = testData5[1158];
@(posedge clk);
#1;data_in = testData5[1159];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1160]; 
@(posedge clk);
#1;data_in = testData5[1161];
@(posedge clk);
#1;data_in = testData5[1162];
@(posedge clk);
#1;data_in = testData5[1163];
@(posedge clk);
#1;data_in = testData5[1164];
@(posedge clk);
#1;data_in = testData5[1165];
@(posedge clk);
#1;data_in = testData5[1166];
@(posedge clk);
#1;data_in = testData5[1167];
@(posedge clk);
#1;data_in = testData5[1168];
@(posedge clk);
#1;data_in = testData5[1169];
@(posedge clk);
#1;data_in = testData5[1170];
@(posedge clk);
#1;data_in = testData5[1171];
@(posedge clk);
#1;data_in = testData5[1172];
@(posedge clk);
#1;data_in = testData5[1173];
@(posedge clk);
#1;data_in = testData5[1174];
@(posedge clk);
#1;data_in = testData5[1175];
@(posedge clk);
#1;data_in = testData5[1176];
@(posedge clk);
#1;data_in = testData5[1177];
@(posedge clk);
#1;data_in = testData5[1178];
@(posedge clk);
#1;data_in = testData5[1179];
@(posedge clk);
#1;data_in = testData5[1180];
@(posedge clk);
#1;data_in = testData5[1181];
@(posedge clk);
#1;data_in = testData5[1182];
@(posedge clk);
#1;data_in = testData5[1183];
@(posedge clk);
#1;data_in = testData5[1184];
@(posedge clk);
#1;data_in = testData5[1185];
@(posedge clk);
#1;data_in = testData5[1186];
@(posedge clk);
#1;data_in = testData5[1187];
@(posedge clk);
#1;data_in = testData5[1188];
@(posedge clk);
#1;data_in = testData5[1189];
@(posedge clk);
#1;data_in = testData5[1190];
@(posedge clk);
#1;data_in = testData5[1191];
@(posedge clk);
#1;data_in = testData5[1192];
@(posedge clk);
#1;data_in = testData5[1193];
@(posedge clk);
#1;data_in = testData5[1194];
@(posedge clk);
#1;data_in = testData5[1195];
@(posedge clk);
#1;data_in = testData5[1196];
@(posedge clk);
#1;data_in = testData5[1197];
@(posedge clk);
#1;data_in = testData5[1198];
@(posedge clk);
#1;data_in = testData5[1199];
@(posedge clk);
#1;data_in = testData5[1200];
@(posedge clk);
#1;data_in = testData5[1201];
@(posedge clk);
#1;data_in = testData5[1202];
@(posedge clk);
#1;data_in = testData5[1203];
@(posedge clk);
#1;data_in = testData5[1204];
@(posedge clk);
#1;data_in = testData5[1205];
@(posedge clk);
#1;data_in = testData5[1206];
@(posedge clk);
#1;data_in = testData5[1207];
@(posedge clk);
#1;data_in = testData5[1208];
@(posedge clk);
#1;data_in = testData5[1209];
@(posedge clk);
#1;data_in = testData5[1210];
@(posedge clk);
#1;data_in = testData5[1211];
@(posedge clk);
#1;data_in = testData5[1212];
@(posedge clk);
#1;data_in = testData5[1213];
@(posedge clk);
#1;data_in = testData5[1214];
@(posedge clk);
#1;data_in = testData5[1215];
@(posedge clk);
#1;data_in = testData5[1216];
@(posedge clk);
#1;data_in = testData5[1217];
@(posedge clk);
#1;data_in = testData5[1218];
@(posedge clk);
#1;data_in = testData5[1219];
@(posedge clk);
#1;data_in = testData5[1220];
@(posedge clk);
#1;data_in = testData5[1221];
@(posedge clk);
#1;data_in = testData5[1222];
@(posedge clk);
#1;data_in = testData5[1223];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1224]; 
@(posedge clk);
#1;data_in = testData5[1225];
@(posedge clk);
#1;data_in = testData5[1226];
@(posedge clk);
#1;data_in = testData5[1227];
@(posedge clk);
#1;data_in = testData5[1228];
@(posedge clk);
#1;data_in = testData5[1229];
@(posedge clk);
#1;data_in = testData5[1230];
@(posedge clk);
#1;data_in = testData5[1231];
@(posedge clk);
#1;data_in = testData5[1232];
@(posedge clk);
#1;data_in = testData5[1233];
@(posedge clk);
#1;data_in = testData5[1234];
@(posedge clk);
#1;data_in = testData5[1235];
@(posedge clk);
#1;data_in = testData5[1236];
@(posedge clk);
#1;data_in = testData5[1237];
@(posedge clk);
#1;data_in = testData5[1238];
@(posedge clk);
#1;data_in = testData5[1239];
@(posedge clk);
#1;data_in = testData5[1240];
@(posedge clk);
#1;data_in = testData5[1241];
@(posedge clk);
#1;data_in = testData5[1242];
@(posedge clk);
#1;data_in = testData5[1243];
@(posedge clk);
#1;data_in = testData5[1244];
@(posedge clk);
#1;data_in = testData5[1245];
@(posedge clk);
#1;data_in = testData5[1246];
@(posedge clk);
#1;data_in = testData5[1247];
@(posedge clk);
#1;data_in = testData5[1248];
@(posedge clk);
#1;data_in = testData5[1249];
@(posedge clk);
#1;data_in = testData5[1250];
@(posedge clk);
#1;data_in = testData5[1251];
@(posedge clk);
#1;data_in = testData5[1252];
@(posedge clk);
#1;data_in = testData5[1253];
@(posedge clk);
#1;data_in = testData5[1254];
@(posedge clk);
#1;data_in = testData5[1255];
@(posedge clk);
#1;data_in = testData5[1256];
@(posedge clk);
#1;data_in = testData5[1257];
@(posedge clk);
#1;data_in = testData5[1258];
@(posedge clk);
#1;data_in = testData5[1259];
@(posedge clk);
#1;data_in = testData5[1260];
@(posedge clk);
#1;data_in = testData5[1261];
@(posedge clk);
#1;data_in = testData5[1262];
@(posedge clk);
#1;data_in = testData5[1263];
@(posedge clk);
#1;data_in = testData5[1264];
@(posedge clk);
#1;data_in = testData5[1265];
@(posedge clk);
#1;data_in = testData5[1266];
@(posedge clk);
#1;data_in = testData5[1267];
@(posedge clk);
#1;data_in = testData5[1268];
@(posedge clk);
#1;data_in = testData5[1269];
@(posedge clk);
#1;data_in = testData5[1270];
@(posedge clk);
#1;data_in = testData5[1271];
@(posedge clk);
#1;data_in = testData5[1272];
@(posedge clk);
#1;data_in = testData5[1273];
@(posedge clk);
#1;data_in = testData5[1274];
@(posedge clk);
#1;data_in = testData5[1275];
@(posedge clk);
#1;data_in = testData5[1276];
@(posedge clk);
#1;data_in = testData5[1277];
@(posedge clk);
#1;data_in = testData5[1278];
@(posedge clk);
#1;data_in = testData5[1279];
@(posedge clk);
#1;data_in = testData5[1280];
@(posedge clk);
#1;data_in = testData5[1281];
@(posedge clk);
#1;data_in = testData5[1282];
@(posedge clk);
#1;data_in = testData5[1283];
@(posedge clk);
#1;data_in = testData5[1284];
@(posedge clk);
#1;data_in = testData5[1285];
@(posedge clk);
#1;data_in = testData5[1286];
@(posedge clk);
#1;data_in = testData5[1287];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1288]; 
@(posedge clk);
#1;data_in = testData5[1289];
@(posedge clk);
#1;data_in = testData5[1290];
@(posedge clk);
#1;data_in = testData5[1291];
@(posedge clk);
#1;data_in = testData5[1292];
@(posedge clk);
#1;data_in = testData5[1293];
@(posedge clk);
#1;data_in = testData5[1294];
@(posedge clk);
#1;data_in = testData5[1295];
@(posedge clk);
#1;data_in = testData5[1296];
@(posedge clk);
#1;data_in = testData5[1297];
@(posedge clk);
#1;data_in = testData5[1298];
@(posedge clk);
#1;data_in = testData5[1299];
@(posedge clk);
#1;data_in = testData5[1300];
@(posedge clk);
#1;data_in = testData5[1301];
@(posedge clk);
#1;data_in = testData5[1302];
@(posedge clk);
#1;data_in = testData5[1303];
@(posedge clk);
#1;data_in = testData5[1304];
@(posedge clk);
#1;data_in = testData5[1305];
@(posedge clk);
#1;data_in = testData5[1306];
@(posedge clk);
#1;data_in = testData5[1307];
@(posedge clk);
#1;data_in = testData5[1308];
@(posedge clk);
#1;data_in = testData5[1309];
@(posedge clk);
#1;data_in = testData5[1310];
@(posedge clk);
#1;data_in = testData5[1311];
@(posedge clk);
#1;data_in = testData5[1312];
@(posedge clk);
#1;data_in = testData5[1313];
@(posedge clk);
#1;data_in = testData5[1314];
@(posedge clk);
#1;data_in = testData5[1315];
@(posedge clk);
#1;data_in = testData5[1316];
@(posedge clk);
#1;data_in = testData5[1317];
@(posedge clk);
#1;data_in = testData5[1318];
@(posedge clk);
#1;data_in = testData5[1319];
@(posedge clk);
#1;data_in = testData5[1320];
@(posedge clk);
#1;data_in = testData5[1321];
@(posedge clk);
#1;data_in = testData5[1322];
@(posedge clk);
#1;data_in = testData5[1323];
@(posedge clk);
#1;data_in = testData5[1324];
@(posedge clk);
#1;data_in = testData5[1325];
@(posedge clk);
#1;data_in = testData5[1326];
@(posedge clk);
#1;data_in = testData5[1327];
@(posedge clk);
#1;data_in = testData5[1328];
@(posedge clk);
#1;data_in = testData5[1329];
@(posedge clk);
#1;data_in = testData5[1330];
@(posedge clk);
#1;data_in = testData5[1331];
@(posedge clk);
#1;data_in = testData5[1332];
@(posedge clk);
#1;data_in = testData5[1333];
@(posedge clk);
#1;data_in = testData5[1334];
@(posedge clk);
#1;data_in = testData5[1335];
@(posedge clk);
#1;data_in = testData5[1336];
@(posedge clk);
#1;data_in = testData5[1337];
@(posedge clk);
#1;data_in = testData5[1338];
@(posedge clk);
#1;data_in = testData5[1339];
@(posedge clk);
#1;data_in = testData5[1340];
@(posedge clk);
#1;data_in = testData5[1341];
@(posedge clk);
#1;data_in = testData5[1342];
@(posedge clk);
#1;data_in = testData5[1343];
@(posedge clk);
#1;data_in = testData5[1344];
@(posedge clk);
#1;data_in = testData5[1345];
@(posedge clk);
#1;data_in = testData5[1346];
@(posedge clk);
#1;data_in = testData5[1347];
@(posedge clk);
#1;data_in = testData5[1348];
@(posedge clk);
#1;data_in = testData5[1349];
@(posedge clk);
#1;data_in = testData5[1350];
@(posedge clk);
#1;data_in = testData5[1351];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1352]; 
@(posedge clk);
#1;data_in = testData5[1353];
@(posedge clk);
#1;data_in = testData5[1354];
@(posedge clk);
#1;data_in = testData5[1355];
@(posedge clk);
#1;data_in = testData5[1356];
@(posedge clk);
#1;data_in = testData5[1357];
@(posedge clk);
#1;data_in = testData5[1358];
@(posedge clk);
#1;data_in = testData5[1359];
@(posedge clk);
#1;data_in = testData5[1360];
@(posedge clk);
#1;data_in = testData5[1361];
@(posedge clk);
#1;data_in = testData5[1362];
@(posedge clk);
#1;data_in = testData5[1363];
@(posedge clk);
#1;data_in = testData5[1364];
@(posedge clk);
#1;data_in = testData5[1365];
@(posedge clk);
#1;data_in = testData5[1366];
@(posedge clk);
#1;data_in = testData5[1367];
@(posedge clk);
#1;data_in = testData5[1368];
@(posedge clk);
#1;data_in = testData5[1369];
@(posedge clk);
#1;data_in = testData5[1370];
@(posedge clk);
#1;data_in = testData5[1371];
@(posedge clk);
#1;data_in = testData5[1372];
@(posedge clk);
#1;data_in = testData5[1373];
@(posedge clk);
#1;data_in = testData5[1374];
@(posedge clk);
#1;data_in = testData5[1375];
@(posedge clk);
#1;data_in = testData5[1376];
@(posedge clk);
#1;data_in = testData5[1377];
@(posedge clk);
#1;data_in = testData5[1378];
@(posedge clk);
#1;data_in = testData5[1379];
@(posedge clk);
#1;data_in = testData5[1380];
@(posedge clk);
#1;data_in = testData5[1381];
@(posedge clk);
#1;data_in = testData5[1382];
@(posedge clk);
#1;data_in = testData5[1383];
@(posedge clk);
#1;data_in = testData5[1384];
@(posedge clk);
#1;data_in = testData5[1385];
@(posedge clk);
#1;data_in = testData5[1386];
@(posedge clk);
#1;data_in = testData5[1387];
@(posedge clk);
#1;data_in = testData5[1388];
@(posedge clk);
#1;data_in = testData5[1389];
@(posedge clk);
#1;data_in = testData5[1390];
@(posedge clk);
#1;data_in = testData5[1391];
@(posedge clk);
#1;data_in = testData5[1392];
@(posedge clk);
#1;data_in = testData5[1393];
@(posedge clk);
#1;data_in = testData5[1394];
@(posedge clk);
#1;data_in = testData5[1395];
@(posedge clk);
#1;data_in = testData5[1396];
@(posedge clk);
#1;data_in = testData5[1397];
@(posedge clk);
#1;data_in = testData5[1398];
@(posedge clk);
#1;data_in = testData5[1399];
@(posedge clk);
#1;data_in = testData5[1400];
@(posedge clk);
#1;data_in = testData5[1401];
@(posedge clk);
#1;data_in = testData5[1402];
@(posedge clk);
#1;data_in = testData5[1403];
@(posedge clk);
#1;data_in = testData5[1404];
@(posedge clk);
#1;data_in = testData5[1405];
@(posedge clk);
#1;data_in = testData5[1406];
@(posedge clk);
#1;data_in = testData5[1407];
@(posedge clk);
#1;data_in = testData5[1408];
@(posedge clk);
#1;data_in = testData5[1409];
@(posedge clk);
#1;data_in = testData5[1410];
@(posedge clk);
#1;data_in = testData5[1411];
@(posedge clk);
#1;data_in = testData5[1412];
@(posedge clk);
#1;data_in = testData5[1413];
@(posedge clk);
#1;data_in = testData5[1414];
@(posedge clk);
#1;data_in = testData5[1415];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1416]; 
@(posedge clk);
#1;data_in = testData5[1417];
@(posedge clk);
#1;data_in = testData5[1418];
@(posedge clk);
#1;data_in = testData5[1419];
@(posedge clk);
#1;data_in = testData5[1420];
@(posedge clk);
#1;data_in = testData5[1421];
@(posedge clk);
#1;data_in = testData5[1422];
@(posedge clk);
#1;data_in = testData5[1423];
@(posedge clk);
#1;data_in = testData5[1424];
@(posedge clk);
#1;data_in = testData5[1425];
@(posedge clk);
#1;data_in = testData5[1426];
@(posedge clk);
#1;data_in = testData5[1427];
@(posedge clk);
#1;data_in = testData5[1428];
@(posedge clk);
#1;data_in = testData5[1429];
@(posedge clk);
#1;data_in = testData5[1430];
@(posedge clk);
#1;data_in = testData5[1431];
@(posedge clk);
#1;data_in = testData5[1432];
@(posedge clk);
#1;data_in = testData5[1433];
@(posedge clk);
#1;data_in = testData5[1434];
@(posedge clk);
#1;data_in = testData5[1435];
@(posedge clk);
#1;data_in = testData5[1436];
@(posedge clk);
#1;data_in = testData5[1437];
@(posedge clk);
#1;data_in = testData5[1438];
@(posedge clk);
#1;data_in = testData5[1439];
@(posedge clk);
#1;data_in = testData5[1440];
@(posedge clk);
#1;data_in = testData5[1441];
@(posedge clk);
#1;data_in = testData5[1442];
@(posedge clk);
#1;data_in = testData5[1443];
@(posedge clk);
#1;data_in = testData5[1444];
@(posedge clk);
#1;data_in = testData5[1445];
@(posedge clk);
#1;data_in = testData5[1446];
@(posedge clk);
#1;data_in = testData5[1447];
@(posedge clk);
#1;data_in = testData5[1448];
@(posedge clk);
#1;data_in = testData5[1449];
@(posedge clk);
#1;data_in = testData5[1450];
@(posedge clk);
#1;data_in = testData5[1451];
@(posedge clk);
#1;data_in = testData5[1452];
@(posedge clk);
#1;data_in = testData5[1453];
@(posedge clk);
#1;data_in = testData5[1454];
@(posedge clk);
#1;data_in = testData5[1455];
@(posedge clk);
#1;data_in = testData5[1456];
@(posedge clk);
#1;data_in = testData5[1457];
@(posedge clk);
#1;data_in = testData5[1458];
@(posedge clk);
#1;data_in = testData5[1459];
@(posedge clk);
#1;data_in = testData5[1460];
@(posedge clk);
#1;data_in = testData5[1461];
@(posedge clk);
#1;data_in = testData5[1462];
@(posedge clk);
#1;data_in = testData5[1463];
@(posedge clk);
#1;data_in = testData5[1464];
@(posedge clk);
#1;data_in = testData5[1465];
@(posedge clk);
#1;data_in = testData5[1466];
@(posedge clk);
#1;data_in = testData5[1467];
@(posedge clk);
#1;data_in = testData5[1468];
@(posedge clk);
#1;data_in = testData5[1469];
@(posedge clk);
#1;data_in = testData5[1470];
@(posedge clk);
#1;data_in = testData5[1471];
@(posedge clk);
#1;data_in = testData5[1472];
@(posedge clk);
#1;data_in = testData5[1473];
@(posedge clk);
#1;data_in = testData5[1474];
@(posedge clk);
#1;data_in = testData5[1475];
@(posedge clk);
#1;data_in = testData5[1476];
@(posedge clk);
#1;data_in = testData5[1477];
@(posedge clk);
#1;data_in = testData5[1478];
@(posedge clk);
#1;data_in = testData5[1479];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1480]; 
@(posedge clk);
#1;data_in = testData5[1481];
@(posedge clk);
#1;data_in = testData5[1482];
@(posedge clk);
#1;data_in = testData5[1483];
@(posedge clk);
#1;data_in = testData5[1484];
@(posedge clk);
#1;data_in = testData5[1485];
@(posedge clk);
#1;data_in = testData5[1486];
@(posedge clk);
#1;data_in = testData5[1487];
@(posedge clk);
#1;data_in = testData5[1488];
@(posedge clk);
#1;data_in = testData5[1489];
@(posedge clk);
#1;data_in = testData5[1490];
@(posedge clk);
#1;data_in = testData5[1491];
@(posedge clk);
#1;data_in = testData5[1492];
@(posedge clk);
#1;data_in = testData5[1493];
@(posedge clk);
#1;data_in = testData5[1494];
@(posedge clk);
#1;data_in = testData5[1495];
@(posedge clk);
#1;data_in = testData5[1496];
@(posedge clk);
#1;data_in = testData5[1497];
@(posedge clk);
#1;data_in = testData5[1498];
@(posedge clk);
#1;data_in = testData5[1499];
@(posedge clk);
#1;data_in = testData5[1500];
@(posedge clk);
#1;data_in = testData5[1501];
@(posedge clk);
#1;data_in = testData5[1502];
@(posedge clk);
#1;data_in = testData5[1503];
@(posedge clk);
#1;data_in = testData5[1504];
@(posedge clk);
#1;data_in = testData5[1505];
@(posedge clk);
#1;data_in = testData5[1506];
@(posedge clk);
#1;data_in = testData5[1507];
@(posedge clk);
#1;data_in = testData5[1508];
@(posedge clk);
#1;data_in = testData5[1509];
@(posedge clk);
#1;data_in = testData5[1510];
@(posedge clk);
#1;data_in = testData5[1511];
@(posedge clk);
#1;data_in = testData5[1512];
@(posedge clk);
#1;data_in = testData5[1513];
@(posedge clk);
#1;data_in = testData5[1514];
@(posedge clk);
#1;data_in = testData5[1515];
@(posedge clk);
#1;data_in = testData5[1516];
@(posedge clk);
#1;data_in = testData5[1517];
@(posedge clk);
#1;data_in = testData5[1518];
@(posedge clk);
#1;data_in = testData5[1519];
@(posedge clk);
#1;data_in = testData5[1520];
@(posedge clk);
#1;data_in = testData5[1521];
@(posedge clk);
#1;data_in = testData5[1522];
@(posedge clk);
#1;data_in = testData5[1523];
@(posedge clk);
#1;data_in = testData5[1524];
@(posedge clk);
#1;data_in = testData5[1525];
@(posedge clk);
#1;data_in = testData5[1526];
@(posedge clk);
#1;data_in = testData5[1527];
@(posedge clk);
#1;data_in = testData5[1528];
@(posedge clk);
#1;data_in = testData5[1529];
@(posedge clk);
#1;data_in = testData5[1530];
@(posedge clk);
#1;data_in = testData5[1531];
@(posedge clk);
#1;data_in = testData5[1532];
@(posedge clk);
#1;data_in = testData5[1533];
@(posedge clk);
#1;data_in = testData5[1534];
@(posedge clk);
#1;data_in = testData5[1535];
@(posedge clk);
#1;data_in = testData5[1536];
@(posedge clk);
#1;data_in = testData5[1537];
@(posedge clk);
#1;data_in = testData5[1538];
@(posedge clk);
#1;data_in = testData5[1539];
@(posedge clk);
#1;data_in = testData5[1540];
@(posedge clk);
#1;data_in = testData5[1541];
@(posedge clk);
#1;data_in = testData5[1542];
@(posedge clk);
#1;data_in = testData5[1543];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1544]; 
@(posedge clk);
#1;data_in = testData5[1545];
@(posedge clk);
#1;data_in = testData5[1546];
@(posedge clk);
#1;data_in = testData5[1547];
@(posedge clk);
#1;data_in = testData5[1548];
@(posedge clk);
#1;data_in = testData5[1549];
@(posedge clk);
#1;data_in = testData5[1550];
@(posedge clk);
#1;data_in = testData5[1551];
@(posedge clk);
#1;data_in = testData5[1552];
@(posedge clk);
#1;data_in = testData5[1553];
@(posedge clk);
#1;data_in = testData5[1554];
@(posedge clk);
#1;data_in = testData5[1555];
@(posedge clk);
#1;data_in = testData5[1556];
@(posedge clk);
#1;data_in = testData5[1557];
@(posedge clk);
#1;data_in = testData5[1558];
@(posedge clk);
#1;data_in = testData5[1559];
@(posedge clk);
#1;data_in = testData5[1560];
@(posedge clk);
#1;data_in = testData5[1561];
@(posedge clk);
#1;data_in = testData5[1562];
@(posedge clk);
#1;data_in = testData5[1563];
@(posedge clk);
#1;data_in = testData5[1564];
@(posedge clk);
#1;data_in = testData5[1565];
@(posedge clk);
#1;data_in = testData5[1566];
@(posedge clk);
#1;data_in = testData5[1567];
@(posedge clk);
#1;data_in = testData5[1568];
@(posedge clk);
#1;data_in = testData5[1569];
@(posedge clk);
#1;data_in = testData5[1570];
@(posedge clk);
#1;data_in = testData5[1571];
@(posedge clk);
#1;data_in = testData5[1572];
@(posedge clk);
#1;data_in = testData5[1573];
@(posedge clk);
#1;data_in = testData5[1574];
@(posedge clk);
#1;data_in = testData5[1575];
@(posedge clk);
#1;data_in = testData5[1576];
@(posedge clk);
#1;data_in = testData5[1577];
@(posedge clk);
#1;data_in = testData5[1578];
@(posedge clk);
#1;data_in = testData5[1579];
@(posedge clk);
#1;data_in = testData5[1580];
@(posedge clk);
#1;data_in = testData5[1581];
@(posedge clk);
#1;data_in = testData5[1582];
@(posedge clk);
#1;data_in = testData5[1583];
@(posedge clk);
#1;data_in = testData5[1584];
@(posedge clk);
#1;data_in = testData5[1585];
@(posedge clk);
#1;data_in = testData5[1586];
@(posedge clk);
#1;data_in = testData5[1587];
@(posedge clk);
#1;data_in = testData5[1588];
@(posedge clk);
#1;data_in = testData5[1589];
@(posedge clk);
#1;data_in = testData5[1590];
@(posedge clk);
#1;data_in = testData5[1591];
@(posedge clk);
#1;data_in = testData5[1592];
@(posedge clk);
#1;data_in = testData5[1593];
@(posedge clk);
#1;data_in = testData5[1594];
@(posedge clk);
#1;data_in = testData5[1595];
@(posedge clk);
#1;data_in = testData5[1596];
@(posedge clk);
#1;data_in = testData5[1597];
@(posedge clk);
#1;data_in = testData5[1598];
@(posedge clk);
#1;data_in = testData5[1599];
@(posedge clk);
#1;data_in = testData5[1600];
@(posedge clk);
#1;data_in = testData5[1601];
@(posedge clk);
#1;data_in = testData5[1602];
@(posedge clk);
#1;data_in = testData5[1603];
@(posedge clk);
#1;data_in = testData5[1604];
@(posedge clk);
#1;data_in = testData5[1605];
@(posedge clk);
#1;data_in = testData5[1606];
@(posedge clk);
#1;data_in = testData5[1607];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1608]; 
@(posedge clk);
#1;data_in = testData5[1609];
@(posedge clk);
#1;data_in = testData5[1610];
@(posedge clk);
#1;data_in = testData5[1611];
@(posedge clk);
#1;data_in = testData5[1612];
@(posedge clk);
#1;data_in = testData5[1613];
@(posedge clk);
#1;data_in = testData5[1614];
@(posedge clk);
#1;data_in = testData5[1615];
@(posedge clk);
#1;data_in = testData5[1616];
@(posedge clk);
#1;data_in = testData5[1617];
@(posedge clk);
#1;data_in = testData5[1618];
@(posedge clk);
#1;data_in = testData5[1619];
@(posedge clk);
#1;data_in = testData5[1620];
@(posedge clk);
#1;data_in = testData5[1621];
@(posedge clk);
#1;data_in = testData5[1622];
@(posedge clk);
#1;data_in = testData5[1623];
@(posedge clk);
#1;data_in = testData5[1624];
@(posedge clk);
#1;data_in = testData5[1625];
@(posedge clk);
#1;data_in = testData5[1626];
@(posedge clk);
#1;data_in = testData5[1627];
@(posedge clk);
#1;data_in = testData5[1628];
@(posedge clk);
#1;data_in = testData5[1629];
@(posedge clk);
#1;data_in = testData5[1630];
@(posedge clk);
#1;data_in = testData5[1631];
@(posedge clk);
#1;data_in = testData5[1632];
@(posedge clk);
#1;data_in = testData5[1633];
@(posedge clk);
#1;data_in = testData5[1634];
@(posedge clk);
#1;data_in = testData5[1635];
@(posedge clk);
#1;data_in = testData5[1636];
@(posedge clk);
#1;data_in = testData5[1637];
@(posedge clk);
#1;data_in = testData5[1638];
@(posedge clk);
#1;data_in = testData5[1639];
@(posedge clk);
#1;data_in = testData5[1640];
@(posedge clk);
#1;data_in = testData5[1641];
@(posedge clk);
#1;data_in = testData5[1642];
@(posedge clk);
#1;data_in = testData5[1643];
@(posedge clk);
#1;data_in = testData5[1644];
@(posedge clk);
#1;data_in = testData5[1645];
@(posedge clk);
#1;data_in = testData5[1646];
@(posedge clk);
#1;data_in = testData5[1647];
@(posedge clk);
#1;data_in = testData5[1648];
@(posedge clk);
#1;data_in = testData5[1649];
@(posedge clk);
#1;data_in = testData5[1650];
@(posedge clk);
#1;data_in = testData5[1651];
@(posedge clk);
#1;data_in = testData5[1652];
@(posedge clk);
#1;data_in = testData5[1653];
@(posedge clk);
#1;data_in = testData5[1654];
@(posedge clk);
#1;data_in = testData5[1655];
@(posedge clk);
#1;data_in = testData5[1656];
@(posedge clk);
#1;data_in = testData5[1657];
@(posedge clk);
#1;data_in = testData5[1658];
@(posedge clk);
#1;data_in = testData5[1659];
@(posedge clk);
#1;data_in = testData5[1660];
@(posedge clk);
#1;data_in = testData5[1661];
@(posedge clk);
#1;data_in = testData5[1662];
@(posedge clk);
#1;data_in = testData5[1663];
@(posedge clk);
#1;data_in = testData5[1664];
@(posedge clk);
#1;data_in = testData5[1665];
@(posedge clk);
#1;data_in = testData5[1666];
@(posedge clk);
#1;data_in = testData5[1667];
@(posedge clk);
#1;data_in = testData5[1668];
@(posedge clk);
#1;data_in = testData5[1669];
@(posedge clk);
#1;data_in = testData5[1670];
@(posedge clk);
#1;data_in = testData5[1671];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1672]; 
@(posedge clk);
#1;data_in = testData5[1673];
@(posedge clk);
#1;data_in = testData5[1674];
@(posedge clk);
#1;data_in = testData5[1675];
@(posedge clk);
#1;data_in = testData5[1676];
@(posedge clk);
#1;data_in = testData5[1677];
@(posedge clk);
#1;data_in = testData5[1678];
@(posedge clk);
#1;data_in = testData5[1679];
@(posedge clk);
#1;data_in = testData5[1680];
@(posedge clk);
#1;data_in = testData5[1681];
@(posedge clk);
#1;data_in = testData5[1682];
@(posedge clk);
#1;data_in = testData5[1683];
@(posedge clk);
#1;data_in = testData5[1684];
@(posedge clk);
#1;data_in = testData5[1685];
@(posedge clk);
#1;data_in = testData5[1686];
@(posedge clk);
#1;data_in = testData5[1687];
@(posedge clk);
#1;data_in = testData5[1688];
@(posedge clk);
#1;data_in = testData5[1689];
@(posedge clk);
#1;data_in = testData5[1690];
@(posedge clk);
#1;data_in = testData5[1691];
@(posedge clk);
#1;data_in = testData5[1692];
@(posedge clk);
#1;data_in = testData5[1693];
@(posedge clk);
#1;data_in = testData5[1694];
@(posedge clk);
#1;data_in = testData5[1695];
@(posedge clk);
#1;data_in = testData5[1696];
@(posedge clk);
#1;data_in = testData5[1697];
@(posedge clk);
#1;data_in = testData5[1698];
@(posedge clk);
#1;data_in = testData5[1699];
@(posedge clk);
#1;data_in = testData5[1700];
@(posedge clk);
#1;data_in = testData5[1701];
@(posedge clk);
#1;data_in = testData5[1702];
@(posedge clk);
#1;data_in = testData5[1703];
@(posedge clk);
#1;data_in = testData5[1704];
@(posedge clk);
#1;data_in = testData5[1705];
@(posedge clk);
#1;data_in = testData5[1706];
@(posedge clk);
#1;data_in = testData5[1707];
@(posedge clk);
#1;data_in = testData5[1708];
@(posedge clk);
#1;data_in = testData5[1709];
@(posedge clk);
#1;data_in = testData5[1710];
@(posedge clk);
#1;data_in = testData5[1711];
@(posedge clk);
#1;data_in = testData5[1712];
@(posedge clk);
#1;data_in = testData5[1713];
@(posedge clk);
#1;data_in = testData5[1714];
@(posedge clk);
#1;data_in = testData5[1715];
@(posedge clk);
#1;data_in = testData5[1716];
@(posedge clk);
#1;data_in = testData5[1717];
@(posedge clk);
#1;data_in = testData5[1718];
@(posedge clk);
#1;data_in = testData5[1719];
@(posedge clk);
#1;data_in = testData5[1720];
@(posedge clk);
#1;data_in = testData5[1721];
@(posedge clk);
#1;data_in = testData5[1722];
@(posedge clk);
#1;data_in = testData5[1723];
@(posedge clk);
#1;data_in = testData5[1724];
@(posedge clk);
#1;data_in = testData5[1725];
@(posedge clk);
#1;data_in = testData5[1726];
@(posedge clk);
#1;data_in = testData5[1727];
@(posedge clk);
#1;data_in = testData5[1728];
@(posedge clk);
#1;data_in = testData5[1729];
@(posedge clk);
#1;data_in = testData5[1730];
@(posedge clk);
#1;data_in = testData5[1731];
@(posedge clk);
#1;data_in = testData5[1732];
@(posedge clk);
#1;data_in = testData5[1733];
@(posedge clk);
#1;data_in = testData5[1734];
@(posedge clk);
#1;data_in = testData5[1735];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1736]; 
@(posedge clk);
#1;data_in = testData5[1737];
@(posedge clk);
#1;data_in = testData5[1738];
@(posedge clk);
#1;data_in = testData5[1739];
@(posedge clk);
#1;data_in = testData5[1740];
@(posedge clk);
#1;data_in = testData5[1741];
@(posedge clk);
#1;data_in = testData5[1742];
@(posedge clk);
#1;data_in = testData5[1743];
@(posedge clk);
#1;data_in = testData5[1744];
@(posedge clk);
#1;data_in = testData5[1745];
@(posedge clk);
#1;data_in = testData5[1746];
@(posedge clk);
#1;data_in = testData5[1747];
@(posedge clk);
#1;data_in = testData5[1748];
@(posedge clk);
#1;data_in = testData5[1749];
@(posedge clk);
#1;data_in = testData5[1750];
@(posedge clk);
#1;data_in = testData5[1751];
@(posedge clk);
#1;data_in = testData5[1752];
@(posedge clk);
#1;data_in = testData5[1753];
@(posedge clk);
#1;data_in = testData5[1754];
@(posedge clk);
#1;data_in = testData5[1755];
@(posedge clk);
#1;data_in = testData5[1756];
@(posedge clk);
#1;data_in = testData5[1757];
@(posedge clk);
#1;data_in = testData5[1758];
@(posedge clk);
#1;data_in = testData5[1759];
@(posedge clk);
#1;data_in = testData5[1760];
@(posedge clk);
#1;data_in = testData5[1761];
@(posedge clk);
#1;data_in = testData5[1762];
@(posedge clk);
#1;data_in = testData5[1763];
@(posedge clk);
#1;data_in = testData5[1764];
@(posedge clk);
#1;data_in = testData5[1765];
@(posedge clk);
#1;data_in = testData5[1766];
@(posedge clk);
#1;data_in = testData5[1767];
@(posedge clk);
#1;data_in = testData5[1768];
@(posedge clk);
#1;data_in = testData5[1769];
@(posedge clk);
#1;data_in = testData5[1770];
@(posedge clk);
#1;data_in = testData5[1771];
@(posedge clk);
#1;data_in = testData5[1772];
@(posedge clk);
#1;data_in = testData5[1773];
@(posedge clk);
#1;data_in = testData5[1774];
@(posedge clk);
#1;data_in = testData5[1775];
@(posedge clk);
#1;data_in = testData5[1776];
@(posedge clk);
#1;data_in = testData5[1777];
@(posedge clk);
#1;data_in = testData5[1778];
@(posedge clk);
#1;data_in = testData5[1779];
@(posedge clk);
#1;data_in = testData5[1780];
@(posedge clk);
#1;data_in = testData5[1781];
@(posedge clk);
#1;data_in = testData5[1782];
@(posedge clk);
#1;data_in = testData5[1783];
@(posedge clk);
#1;data_in = testData5[1784];
@(posedge clk);
#1;data_in = testData5[1785];
@(posedge clk);
#1;data_in = testData5[1786];
@(posedge clk);
#1;data_in = testData5[1787];
@(posedge clk);
#1;data_in = testData5[1788];
@(posedge clk);
#1;data_in = testData5[1789];
@(posedge clk);
#1;data_in = testData5[1790];
@(posedge clk);
#1;data_in = testData5[1791];
@(posedge clk);
#1;data_in = testData5[1792];
@(posedge clk);
#1;data_in = testData5[1793];
@(posedge clk);
#1;data_in = testData5[1794];
@(posedge clk);
#1;data_in = testData5[1795];
@(posedge clk);
#1;data_in = testData5[1796];
@(posedge clk);
#1;data_in = testData5[1797];
@(posedge clk);
#1;data_in = testData5[1798];
@(posedge clk);
#1;data_in = testData5[1799];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1800]; 
@(posedge clk);
#1;data_in = testData5[1801];
@(posedge clk);
#1;data_in = testData5[1802];
@(posedge clk);
#1;data_in = testData5[1803];
@(posedge clk);
#1;data_in = testData5[1804];
@(posedge clk);
#1;data_in = testData5[1805];
@(posedge clk);
#1;data_in = testData5[1806];
@(posedge clk);
#1;data_in = testData5[1807];
@(posedge clk);
#1;data_in = testData5[1808];
@(posedge clk);
#1;data_in = testData5[1809];
@(posedge clk);
#1;data_in = testData5[1810];
@(posedge clk);
#1;data_in = testData5[1811];
@(posedge clk);
#1;data_in = testData5[1812];
@(posedge clk);
#1;data_in = testData5[1813];
@(posedge clk);
#1;data_in = testData5[1814];
@(posedge clk);
#1;data_in = testData5[1815];
@(posedge clk);
#1;data_in = testData5[1816];
@(posedge clk);
#1;data_in = testData5[1817];
@(posedge clk);
#1;data_in = testData5[1818];
@(posedge clk);
#1;data_in = testData5[1819];
@(posedge clk);
#1;data_in = testData5[1820];
@(posedge clk);
#1;data_in = testData5[1821];
@(posedge clk);
#1;data_in = testData5[1822];
@(posedge clk);
#1;data_in = testData5[1823];
@(posedge clk);
#1;data_in = testData5[1824];
@(posedge clk);
#1;data_in = testData5[1825];
@(posedge clk);
#1;data_in = testData5[1826];
@(posedge clk);
#1;data_in = testData5[1827];
@(posedge clk);
#1;data_in = testData5[1828];
@(posedge clk);
#1;data_in = testData5[1829];
@(posedge clk);
#1;data_in = testData5[1830];
@(posedge clk);
#1;data_in = testData5[1831];
@(posedge clk);
#1;data_in = testData5[1832];
@(posedge clk);
#1;data_in = testData5[1833];
@(posedge clk);
#1;data_in = testData5[1834];
@(posedge clk);
#1;data_in = testData5[1835];
@(posedge clk);
#1;data_in = testData5[1836];
@(posedge clk);
#1;data_in = testData5[1837];
@(posedge clk);
#1;data_in = testData5[1838];
@(posedge clk);
#1;data_in = testData5[1839];
@(posedge clk);
#1;data_in = testData5[1840];
@(posedge clk);
#1;data_in = testData5[1841];
@(posedge clk);
#1;data_in = testData5[1842];
@(posedge clk);
#1;data_in = testData5[1843];
@(posedge clk);
#1;data_in = testData5[1844];
@(posedge clk);
#1;data_in = testData5[1845];
@(posedge clk);
#1;data_in = testData5[1846];
@(posedge clk);
#1;data_in = testData5[1847];
@(posedge clk);
#1;data_in = testData5[1848];
@(posedge clk);
#1;data_in = testData5[1849];
@(posedge clk);
#1;data_in = testData5[1850];
@(posedge clk);
#1;data_in = testData5[1851];
@(posedge clk);
#1;data_in = testData5[1852];
@(posedge clk);
#1;data_in = testData5[1853];
@(posedge clk);
#1;data_in = testData5[1854];
@(posedge clk);
#1;data_in = testData5[1855];
@(posedge clk);
#1;data_in = testData5[1856];
@(posedge clk);
#1;data_in = testData5[1857];
@(posedge clk);
#1;data_in = testData5[1858];
@(posedge clk);
#1;data_in = testData5[1859];
@(posedge clk);
#1;data_in = testData5[1860];
@(posedge clk);
#1;data_in = testData5[1861];
@(posedge clk);
#1;data_in = testData5[1862];
@(posedge clk);
#1;data_in = testData5[1863];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1864]; 
@(posedge clk);
#1;data_in = testData5[1865];
@(posedge clk);
#1;data_in = testData5[1866];
@(posedge clk);
#1;data_in = testData5[1867];
@(posedge clk);
#1;data_in = testData5[1868];
@(posedge clk);
#1;data_in = testData5[1869];
@(posedge clk);
#1;data_in = testData5[1870];
@(posedge clk);
#1;data_in = testData5[1871];
@(posedge clk);
#1;data_in = testData5[1872];
@(posedge clk);
#1;data_in = testData5[1873];
@(posedge clk);
#1;data_in = testData5[1874];
@(posedge clk);
#1;data_in = testData5[1875];
@(posedge clk);
#1;data_in = testData5[1876];
@(posedge clk);
#1;data_in = testData5[1877];
@(posedge clk);
#1;data_in = testData5[1878];
@(posedge clk);
#1;data_in = testData5[1879];
@(posedge clk);
#1;data_in = testData5[1880];
@(posedge clk);
#1;data_in = testData5[1881];
@(posedge clk);
#1;data_in = testData5[1882];
@(posedge clk);
#1;data_in = testData5[1883];
@(posedge clk);
#1;data_in = testData5[1884];
@(posedge clk);
#1;data_in = testData5[1885];
@(posedge clk);
#1;data_in = testData5[1886];
@(posedge clk);
#1;data_in = testData5[1887];
@(posedge clk);
#1;data_in = testData5[1888];
@(posedge clk);
#1;data_in = testData5[1889];
@(posedge clk);
#1;data_in = testData5[1890];
@(posedge clk);
#1;data_in = testData5[1891];
@(posedge clk);
#1;data_in = testData5[1892];
@(posedge clk);
#1;data_in = testData5[1893];
@(posedge clk);
#1;data_in = testData5[1894];
@(posedge clk);
#1;data_in = testData5[1895];
@(posedge clk);
#1;data_in = testData5[1896];
@(posedge clk);
#1;data_in = testData5[1897];
@(posedge clk);
#1;data_in = testData5[1898];
@(posedge clk);
#1;data_in = testData5[1899];
@(posedge clk);
#1;data_in = testData5[1900];
@(posedge clk);
#1;data_in = testData5[1901];
@(posedge clk);
#1;data_in = testData5[1902];
@(posedge clk);
#1;data_in = testData5[1903];
@(posedge clk);
#1;data_in = testData5[1904];
@(posedge clk);
#1;data_in = testData5[1905];
@(posedge clk);
#1;data_in = testData5[1906];
@(posedge clk);
#1;data_in = testData5[1907];
@(posedge clk);
#1;data_in = testData5[1908];
@(posedge clk);
#1;data_in = testData5[1909];
@(posedge clk);
#1;data_in = testData5[1910];
@(posedge clk);
#1;data_in = testData5[1911];
@(posedge clk);
#1;data_in = testData5[1912];
@(posedge clk);
#1;data_in = testData5[1913];
@(posedge clk);
#1;data_in = testData5[1914];
@(posedge clk);
#1;data_in = testData5[1915];
@(posedge clk);
#1;data_in = testData5[1916];
@(posedge clk);
#1;data_in = testData5[1917];
@(posedge clk);
#1;data_in = testData5[1918];
@(posedge clk);
#1;data_in = testData5[1919];
@(posedge clk);
#1;data_in = testData5[1920];
@(posedge clk);
#1;data_in = testData5[1921];
@(posedge clk);
#1;data_in = testData5[1922];
@(posedge clk);
#1;data_in = testData5[1923];
@(posedge clk);
#1;data_in = testData5[1924];
@(posedge clk);
#1;data_in = testData5[1925];
@(posedge clk);
#1;data_in = testData5[1926];
@(posedge clk);
#1;data_in = testData5[1927];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1928]; 
@(posedge clk);
#1;data_in = testData5[1929];
@(posedge clk);
#1;data_in = testData5[1930];
@(posedge clk);
#1;data_in = testData5[1931];
@(posedge clk);
#1;data_in = testData5[1932];
@(posedge clk);
#1;data_in = testData5[1933];
@(posedge clk);
#1;data_in = testData5[1934];
@(posedge clk);
#1;data_in = testData5[1935];
@(posedge clk);
#1;data_in = testData5[1936];
@(posedge clk);
#1;data_in = testData5[1937];
@(posedge clk);
#1;data_in = testData5[1938];
@(posedge clk);
#1;data_in = testData5[1939];
@(posedge clk);
#1;data_in = testData5[1940];
@(posedge clk);
#1;data_in = testData5[1941];
@(posedge clk);
#1;data_in = testData5[1942];
@(posedge clk);
#1;data_in = testData5[1943];
@(posedge clk);
#1;data_in = testData5[1944];
@(posedge clk);
#1;data_in = testData5[1945];
@(posedge clk);
#1;data_in = testData5[1946];
@(posedge clk);
#1;data_in = testData5[1947];
@(posedge clk);
#1;data_in = testData5[1948];
@(posedge clk);
#1;data_in = testData5[1949];
@(posedge clk);
#1;data_in = testData5[1950];
@(posedge clk);
#1;data_in = testData5[1951];
@(posedge clk);
#1;data_in = testData5[1952];
@(posedge clk);
#1;data_in = testData5[1953];
@(posedge clk);
#1;data_in = testData5[1954];
@(posedge clk);
#1;data_in = testData5[1955];
@(posedge clk);
#1;data_in = testData5[1956];
@(posedge clk);
#1;data_in = testData5[1957];
@(posedge clk);
#1;data_in = testData5[1958];
@(posedge clk);
#1;data_in = testData5[1959];
@(posedge clk);
#1;data_in = testData5[1960];
@(posedge clk);
#1;data_in = testData5[1961];
@(posedge clk);
#1;data_in = testData5[1962];
@(posedge clk);
#1;data_in = testData5[1963];
@(posedge clk);
#1;data_in = testData5[1964];
@(posedge clk);
#1;data_in = testData5[1965];
@(posedge clk);
#1;data_in = testData5[1966];
@(posedge clk);
#1;data_in = testData5[1967];
@(posedge clk);
#1;data_in = testData5[1968];
@(posedge clk);
#1;data_in = testData5[1969];
@(posedge clk);
#1;data_in = testData5[1970];
@(posedge clk);
#1;data_in = testData5[1971];
@(posedge clk);
#1;data_in = testData5[1972];
@(posedge clk);
#1;data_in = testData5[1973];
@(posedge clk);
#1;data_in = testData5[1974];
@(posedge clk);
#1;data_in = testData5[1975];
@(posedge clk);
#1;data_in = testData5[1976];
@(posedge clk);
#1;data_in = testData5[1977];
@(posedge clk);
#1;data_in = testData5[1978];
@(posedge clk);
#1;data_in = testData5[1979];
@(posedge clk);
#1;data_in = testData5[1980];
@(posedge clk);
#1;data_in = testData5[1981];
@(posedge clk);
#1;data_in = testData5[1982];
@(posedge clk);
#1;data_in = testData5[1983];
@(posedge clk);
#1;data_in = testData5[1984];
@(posedge clk);
#1;data_in = testData5[1985];
@(posedge clk);
#1;data_in = testData5[1986];
@(posedge clk);
#1;data_in = testData5[1987];
@(posedge clk);
#1;data_in = testData5[1988];
@(posedge clk);
#1;data_in = testData5[1989];
@(posedge clk);
#1;data_in = testData5[1990];
@(posedge clk);
#1;data_in = testData5[1991];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[1992]; 
@(posedge clk);
#1;data_in = testData5[1993];
@(posedge clk);
#1;data_in = testData5[1994];
@(posedge clk);
#1;data_in = testData5[1995];
@(posedge clk);
#1;data_in = testData5[1996];
@(posedge clk);
#1;data_in = testData5[1997];
@(posedge clk);
#1;data_in = testData5[1998];
@(posedge clk);
#1;data_in = testData5[1999];
@(posedge clk);
#1;data_in = testData5[2000];
@(posedge clk);
#1;data_in = testData5[2001];
@(posedge clk);
#1;data_in = testData5[2002];
@(posedge clk);
#1;data_in = testData5[2003];
@(posedge clk);
#1;data_in = testData5[2004];
@(posedge clk);
#1;data_in = testData5[2005];
@(posedge clk);
#1;data_in = testData5[2006];
@(posedge clk);
#1;data_in = testData5[2007];
@(posedge clk);
#1;data_in = testData5[2008];
@(posedge clk);
#1;data_in = testData5[2009];
@(posedge clk);
#1;data_in = testData5[2010];
@(posedge clk);
#1;data_in = testData5[2011];
@(posedge clk);
#1;data_in = testData5[2012];
@(posedge clk);
#1;data_in = testData5[2013];
@(posedge clk);
#1;data_in = testData5[2014];
@(posedge clk);
#1;data_in = testData5[2015];
@(posedge clk);
#1;data_in = testData5[2016];
@(posedge clk);
#1;data_in = testData5[2017];
@(posedge clk);
#1;data_in = testData5[2018];
@(posedge clk);
#1;data_in = testData5[2019];
@(posedge clk);
#1;data_in = testData5[2020];
@(posedge clk);
#1;data_in = testData5[2021];
@(posedge clk);
#1;data_in = testData5[2022];
@(posedge clk);
#1;data_in = testData5[2023];
@(posedge clk);
#1;data_in = testData5[2024];
@(posedge clk);
#1;data_in = testData5[2025];
@(posedge clk);
#1;data_in = testData5[2026];
@(posedge clk);
#1;data_in = testData5[2027];
@(posedge clk);
#1;data_in = testData5[2028];
@(posedge clk);
#1;data_in = testData5[2029];
@(posedge clk);
#1;data_in = testData5[2030];
@(posedge clk);
#1;data_in = testData5[2031];
@(posedge clk);
#1;data_in = testData5[2032];
@(posedge clk);
#1;data_in = testData5[2033];
@(posedge clk);
#1;data_in = testData5[2034];
@(posedge clk);
#1;data_in = testData5[2035];
@(posedge clk);
#1;data_in = testData5[2036];
@(posedge clk);
#1;data_in = testData5[2037];
@(posedge clk);
#1;data_in = testData5[2038];
@(posedge clk);
#1;data_in = testData5[2039];
@(posedge clk);
#1;data_in = testData5[2040];
@(posedge clk);
#1;data_in = testData5[2041];
@(posedge clk);
#1;data_in = testData5[2042];
@(posedge clk);
#1;data_in = testData5[2043];
@(posedge clk);
#1;data_in = testData5[2044];
@(posedge clk);
#1;data_in = testData5[2045];
@(posedge clk);
#1;data_in = testData5[2046];
@(posedge clk);
#1;data_in = testData5[2047];
@(posedge clk);
#1;data_in = testData5[2048];
@(posedge clk);
#1;data_in = testData5[2049];
@(posedge clk);
#1;data_in = testData5[2050];
@(posedge clk);
#1;data_in = testData5[2051];
@(posedge clk);
#1;data_in = testData5[2052];
@(posedge clk);
#1;data_in = testData5[2053];
@(posedge clk);
#1;data_in = testData5[2054];
@(posedge clk);
#1;data_in = testData5[2055];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2056]; 
@(posedge clk);
#1;data_in = testData5[2057];
@(posedge clk);
#1;data_in = testData5[2058];
@(posedge clk);
#1;data_in = testData5[2059];
@(posedge clk);
#1;data_in = testData5[2060];
@(posedge clk);
#1;data_in = testData5[2061];
@(posedge clk);
#1;data_in = testData5[2062];
@(posedge clk);
#1;data_in = testData5[2063];
@(posedge clk);
#1;data_in = testData5[2064];
@(posedge clk);
#1;data_in = testData5[2065];
@(posedge clk);
#1;data_in = testData5[2066];
@(posedge clk);
#1;data_in = testData5[2067];
@(posedge clk);
#1;data_in = testData5[2068];
@(posedge clk);
#1;data_in = testData5[2069];
@(posedge clk);
#1;data_in = testData5[2070];
@(posedge clk);
#1;data_in = testData5[2071];
@(posedge clk);
#1;data_in = testData5[2072];
@(posedge clk);
#1;data_in = testData5[2073];
@(posedge clk);
#1;data_in = testData5[2074];
@(posedge clk);
#1;data_in = testData5[2075];
@(posedge clk);
#1;data_in = testData5[2076];
@(posedge clk);
#1;data_in = testData5[2077];
@(posedge clk);
#1;data_in = testData5[2078];
@(posedge clk);
#1;data_in = testData5[2079];
@(posedge clk);
#1;data_in = testData5[2080];
@(posedge clk);
#1;data_in = testData5[2081];
@(posedge clk);
#1;data_in = testData5[2082];
@(posedge clk);
#1;data_in = testData5[2083];
@(posedge clk);
#1;data_in = testData5[2084];
@(posedge clk);
#1;data_in = testData5[2085];
@(posedge clk);
#1;data_in = testData5[2086];
@(posedge clk);
#1;data_in = testData5[2087];
@(posedge clk);
#1;data_in = testData5[2088];
@(posedge clk);
#1;data_in = testData5[2089];
@(posedge clk);
#1;data_in = testData5[2090];
@(posedge clk);
#1;data_in = testData5[2091];
@(posedge clk);
#1;data_in = testData5[2092];
@(posedge clk);
#1;data_in = testData5[2093];
@(posedge clk);
#1;data_in = testData5[2094];
@(posedge clk);
#1;data_in = testData5[2095];
@(posedge clk);
#1;data_in = testData5[2096];
@(posedge clk);
#1;data_in = testData5[2097];
@(posedge clk);
#1;data_in = testData5[2098];
@(posedge clk);
#1;data_in = testData5[2099];
@(posedge clk);
#1;data_in = testData5[2100];
@(posedge clk);
#1;data_in = testData5[2101];
@(posedge clk);
#1;data_in = testData5[2102];
@(posedge clk);
#1;data_in = testData5[2103];
@(posedge clk);
#1;data_in = testData5[2104];
@(posedge clk);
#1;data_in = testData5[2105];
@(posedge clk);
#1;data_in = testData5[2106];
@(posedge clk);
#1;data_in = testData5[2107];
@(posedge clk);
#1;data_in = testData5[2108];
@(posedge clk);
#1;data_in = testData5[2109];
@(posedge clk);
#1;data_in = testData5[2110];
@(posedge clk);
#1;data_in = testData5[2111];
@(posedge clk);
#1;data_in = testData5[2112];
@(posedge clk);
#1;data_in = testData5[2113];
@(posedge clk);
#1;data_in = testData5[2114];
@(posedge clk);
#1;data_in = testData5[2115];
@(posedge clk);
#1;data_in = testData5[2116];
@(posedge clk);
#1;data_in = testData5[2117];
@(posedge clk);
#1;data_in = testData5[2118];
@(posedge clk);
#1;data_in = testData5[2119];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2120]; 
@(posedge clk);
#1;data_in = testData5[2121];
@(posedge clk);
#1;data_in = testData5[2122];
@(posedge clk);
#1;data_in = testData5[2123];
@(posedge clk);
#1;data_in = testData5[2124];
@(posedge clk);
#1;data_in = testData5[2125];
@(posedge clk);
#1;data_in = testData5[2126];
@(posedge clk);
#1;data_in = testData5[2127];
@(posedge clk);
#1;data_in = testData5[2128];
@(posedge clk);
#1;data_in = testData5[2129];
@(posedge clk);
#1;data_in = testData5[2130];
@(posedge clk);
#1;data_in = testData5[2131];
@(posedge clk);
#1;data_in = testData5[2132];
@(posedge clk);
#1;data_in = testData5[2133];
@(posedge clk);
#1;data_in = testData5[2134];
@(posedge clk);
#1;data_in = testData5[2135];
@(posedge clk);
#1;data_in = testData5[2136];
@(posedge clk);
#1;data_in = testData5[2137];
@(posedge clk);
#1;data_in = testData5[2138];
@(posedge clk);
#1;data_in = testData5[2139];
@(posedge clk);
#1;data_in = testData5[2140];
@(posedge clk);
#1;data_in = testData5[2141];
@(posedge clk);
#1;data_in = testData5[2142];
@(posedge clk);
#1;data_in = testData5[2143];
@(posedge clk);
#1;data_in = testData5[2144];
@(posedge clk);
#1;data_in = testData5[2145];
@(posedge clk);
#1;data_in = testData5[2146];
@(posedge clk);
#1;data_in = testData5[2147];
@(posedge clk);
#1;data_in = testData5[2148];
@(posedge clk);
#1;data_in = testData5[2149];
@(posedge clk);
#1;data_in = testData5[2150];
@(posedge clk);
#1;data_in = testData5[2151];
@(posedge clk);
#1;data_in = testData5[2152];
@(posedge clk);
#1;data_in = testData5[2153];
@(posedge clk);
#1;data_in = testData5[2154];
@(posedge clk);
#1;data_in = testData5[2155];
@(posedge clk);
#1;data_in = testData5[2156];
@(posedge clk);
#1;data_in = testData5[2157];
@(posedge clk);
#1;data_in = testData5[2158];
@(posedge clk);
#1;data_in = testData5[2159];
@(posedge clk);
#1;data_in = testData5[2160];
@(posedge clk);
#1;data_in = testData5[2161];
@(posedge clk);
#1;data_in = testData5[2162];
@(posedge clk);
#1;data_in = testData5[2163];
@(posedge clk);
#1;data_in = testData5[2164];
@(posedge clk);
#1;data_in = testData5[2165];
@(posedge clk);
#1;data_in = testData5[2166];
@(posedge clk);
#1;data_in = testData5[2167];
@(posedge clk);
#1;data_in = testData5[2168];
@(posedge clk);
#1;data_in = testData5[2169];
@(posedge clk);
#1;data_in = testData5[2170];
@(posedge clk);
#1;data_in = testData5[2171];
@(posedge clk);
#1;data_in = testData5[2172];
@(posedge clk);
#1;data_in = testData5[2173];
@(posedge clk);
#1;data_in = testData5[2174];
@(posedge clk);
#1;data_in = testData5[2175];
@(posedge clk);
#1;data_in = testData5[2176];
@(posedge clk);
#1;data_in = testData5[2177];
@(posedge clk);
#1;data_in = testData5[2178];
@(posedge clk);
#1;data_in = testData5[2179];
@(posedge clk);
#1;data_in = testData5[2180];
@(posedge clk);
#1;data_in = testData5[2181];
@(posedge clk);
#1;data_in = testData5[2182];
@(posedge clk);
#1;data_in = testData5[2183];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2184]; 
@(posedge clk);
#1;data_in = testData5[2185];
@(posedge clk);
#1;data_in = testData5[2186];
@(posedge clk);
#1;data_in = testData5[2187];
@(posedge clk);
#1;data_in = testData5[2188];
@(posedge clk);
#1;data_in = testData5[2189];
@(posedge clk);
#1;data_in = testData5[2190];
@(posedge clk);
#1;data_in = testData5[2191];
@(posedge clk);
#1;data_in = testData5[2192];
@(posedge clk);
#1;data_in = testData5[2193];
@(posedge clk);
#1;data_in = testData5[2194];
@(posedge clk);
#1;data_in = testData5[2195];
@(posedge clk);
#1;data_in = testData5[2196];
@(posedge clk);
#1;data_in = testData5[2197];
@(posedge clk);
#1;data_in = testData5[2198];
@(posedge clk);
#1;data_in = testData5[2199];
@(posedge clk);
#1;data_in = testData5[2200];
@(posedge clk);
#1;data_in = testData5[2201];
@(posedge clk);
#1;data_in = testData5[2202];
@(posedge clk);
#1;data_in = testData5[2203];
@(posedge clk);
#1;data_in = testData5[2204];
@(posedge clk);
#1;data_in = testData5[2205];
@(posedge clk);
#1;data_in = testData5[2206];
@(posedge clk);
#1;data_in = testData5[2207];
@(posedge clk);
#1;data_in = testData5[2208];
@(posedge clk);
#1;data_in = testData5[2209];
@(posedge clk);
#1;data_in = testData5[2210];
@(posedge clk);
#1;data_in = testData5[2211];
@(posedge clk);
#1;data_in = testData5[2212];
@(posedge clk);
#1;data_in = testData5[2213];
@(posedge clk);
#1;data_in = testData5[2214];
@(posedge clk);
#1;data_in = testData5[2215];
@(posedge clk);
#1;data_in = testData5[2216];
@(posedge clk);
#1;data_in = testData5[2217];
@(posedge clk);
#1;data_in = testData5[2218];
@(posedge clk);
#1;data_in = testData5[2219];
@(posedge clk);
#1;data_in = testData5[2220];
@(posedge clk);
#1;data_in = testData5[2221];
@(posedge clk);
#1;data_in = testData5[2222];
@(posedge clk);
#1;data_in = testData5[2223];
@(posedge clk);
#1;data_in = testData5[2224];
@(posedge clk);
#1;data_in = testData5[2225];
@(posedge clk);
#1;data_in = testData5[2226];
@(posedge clk);
#1;data_in = testData5[2227];
@(posedge clk);
#1;data_in = testData5[2228];
@(posedge clk);
#1;data_in = testData5[2229];
@(posedge clk);
#1;data_in = testData5[2230];
@(posedge clk);
#1;data_in = testData5[2231];
@(posedge clk);
#1;data_in = testData5[2232];
@(posedge clk);
#1;data_in = testData5[2233];
@(posedge clk);
#1;data_in = testData5[2234];
@(posedge clk);
#1;data_in = testData5[2235];
@(posedge clk);
#1;data_in = testData5[2236];
@(posedge clk);
#1;data_in = testData5[2237];
@(posedge clk);
#1;data_in = testData5[2238];
@(posedge clk);
#1;data_in = testData5[2239];
@(posedge clk);
#1;data_in = testData5[2240];
@(posedge clk);
#1;data_in = testData5[2241];
@(posedge clk);
#1;data_in = testData5[2242];
@(posedge clk);
#1;data_in = testData5[2243];
@(posedge clk);
#1;data_in = testData5[2244];
@(posedge clk);
#1;data_in = testData5[2245];
@(posedge clk);
#1;data_in = testData5[2246];
@(posedge clk);
#1;data_in = testData5[2247];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2248]; 
@(posedge clk);
#1;data_in = testData5[2249];
@(posedge clk);
#1;data_in = testData5[2250];
@(posedge clk);
#1;data_in = testData5[2251];
@(posedge clk);
#1;data_in = testData5[2252];
@(posedge clk);
#1;data_in = testData5[2253];
@(posedge clk);
#1;data_in = testData5[2254];
@(posedge clk);
#1;data_in = testData5[2255];
@(posedge clk);
#1;data_in = testData5[2256];
@(posedge clk);
#1;data_in = testData5[2257];
@(posedge clk);
#1;data_in = testData5[2258];
@(posedge clk);
#1;data_in = testData5[2259];
@(posedge clk);
#1;data_in = testData5[2260];
@(posedge clk);
#1;data_in = testData5[2261];
@(posedge clk);
#1;data_in = testData5[2262];
@(posedge clk);
#1;data_in = testData5[2263];
@(posedge clk);
#1;data_in = testData5[2264];
@(posedge clk);
#1;data_in = testData5[2265];
@(posedge clk);
#1;data_in = testData5[2266];
@(posedge clk);
#1;data_in = testData5[2267];
@(posedge clk);
#1;data_in = testData5[2268];
@(posedge clk);
#1;data_in = testData5[2269];
@(posedge clk);
#1;data_in = testData5[2270];
@(posedge clk);
#1;data_in = testData5[2271];
@(posedge clk);
#1;data_in = testData5[2272];
@(posedge clk);
#1;data_in = testData5[2273];
@(posedge clk);
#1;data_in = testData5[2274];
@(posedge clk);
#1;data_in = testData5[2275];
@(posedge clk);
#1;data_in = testData5[2276];
@(posedge clk);
#1;data_in = testData5[2277];
@(posedge clk);
#1;data_in = testData5[2278];
@(posedge clk);
#1;data_in = testData5[2279];
@(posedge clk);
#1;data_in = testData5[2280];
@(posedge clk);
#1;data_in = testData5[2281];
@(posedge clk);
#1;data_in = testData5[2282];
@(posedge clk);
#1;data_in = testData5[2283];
@(posedge clk);
#1;data_in = testData5[2284];
@(posedge clk);
#1;data_in = testData5[2285];
@(posedge clk);
#1;data_in = testData5[2286];
@(posedge clk);
#1;data_in = testData5[2287];
@(posedge clk);
#1;data_in = testData5[2288];
@(posedge clk);
#1;data_in = testData5[2289];
@(posedge clk);
#1;data_in = testData5[2290];
@(posedge clk);
#1;data_in = testData5[2291];
@(posedge clk);
#1;data_in = testData5[2292];
@(posedge clk);
#1;data_in = testData5[2293];
@(posedge clk);
#1;data_in = testData5[2294];
@(posedge clk);
#1;data_in = testData5[2295];
@(posedge clk);
#1;data_in = testData5[2296];
@(posedge clk);
#1;data_in = testData5[2297];
@(posedge clk);
#1;data_in = testData5[2298];
@(posedge clk);
#1;data_in = testData5[2299];
@(posedge clk);
#1;data_in = testData5[2300];
@(posedge clk);
#1;data_in = testData5[2301];
@(posedge clk);
#1;data_in = testData5[2302];
@(posedge clk);
#1;data_in = testData5[2303];
@(posedge clk);
#1;data_in = testData5[2304];
@(posedge clk);
#1;data_in = testData5[2305];
@(posedge clk);
#1;data_in = testData5[2306];
@(posedge clk);
#1;data_in = testData5[2307];
@(posedge clk);
#1;data_in = testData5[2308];
@(posedge clk);
#1;data_in = testData5[2309];
@(posedge clk);
#1;data_in = testData5[2310];
@(posedge clk);
#1;data_in = testData5[2311];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2312]; 
@(posedge clk);
#1;data_in = testData5[2313];
@(posedge clk);
#1;data_in = testData5[2314];
@(posedge clk);
#1;data_in = testData5[2315];
@(posedge clk);
#1;data_in = testData5[2316];
@(posedge clk);
#1;data_in = testData5[2317];
@(posedge clk);
#1;data_in = testData5[2318];
@(posedge clk);
#1;data_in = testData5[2319];
@(posedge clk);
#1;data_in = testData5[2320];
@(posedge clk);
#1;data_in = testData5[2321];
@(posedge clk);
#1;data_in = testData5[2322];
@(posedge clk);
#1;data_in = testData5[2323];
@(posedge clk);
#1;data_in = testData5[2324];
@(posedge clk);
#1;data_in = testData5[2325];
@(posedge clk);
#1;data_in = testData5[2326];
@(posedge clk);
#1;data_in = testData5[2327];
@(posedge clk);
#1;data_in = testData5[2328];
@(posedge clk);
#1;data_in = testData5[2329];
@(posedge clk);
#1;data_in = testData5[2330];
@(posedge clk);
#1;data_in = testData5[2331];
@(posedge clk);
#1;data_in = testData5[2332];
@(posedge clk);
#1;data_in = testData5[2333];
@(posedge clk);
#1;data_in = testData5[2334];
@(posedge clk);
#1;data_in = testData5[2335];
@(posedge clk);
#1;data_in = testData5[2336];
@(posedge clk);
#1;data_in = testData5[2337];
@(posedge clk);
#1;data_in = testData5[2338];
@(posedge clk);
#1;data_in = testData5[2339];
@(posedge clk);
#1;data_in = testData5[2340];
@(posedge clk);
#1;data_in = testData5[2341];
@(posedge clk);
#1;data_in = testData5[2342];
@(posedge clk);
#1;data_in = testData5[2343];
@(posedge clk);
#1;data_in = testData5[2344];
@(posedge clk);
#1;data_in = testData5[2345];
@(posedge clk);
#1;data_in = testData5[2346];
@(posedge clk);
#1;data_in = testData5[2347];
@(posedge clk);
#1;data_in = testData5[2348];
@(posedge clk);
#1;data_in = testData5[2349];
@(posedge clk);
#1;data_in = testData5[2350];
@(posedge clk);
#1;data_in = testData5[2351];
@(posedge clk);
#1;data_in = testData5[2352];
@(posedge clk);
#1;data_in = testData5[2353];
@(posedge clk);
#1;data_in = testData5[2354];
@(posedge clk);
#1;data_in = testData5[2355];
@(posedge clk);
#1;data_in = testData5[2356];
@(posedge clk);
#1;data_in = testData5[2357];
@(posedge clk);
#1;data_in = testData5[2358];
@(posedge clk);
#1;data_in = testData5[2359];
@(posedge clk);
#1;data_in = testData5[2360];
@(posedge clk);
#1;data_in = testData5[2361];
@(posedge clk);
#1;data_in = testData5[2362];
@(posedge clk);
#1;data_in = testData5[2363];
@(posedge clk);
#1;data_in = testData5[2364];
@(posedge clk);
#1;data_in = testData5[2365];
@(posedge clk);
#1;data_in = testData5[2366];
@(posedge clk);
#1;data_in = testData5[2367];
@(posedge clk);
#1;data_in = testData5[2368];
@(posedge clk);
#1;data_in = testData5[2369];
@(posedge clk);
#1;data_in = testData5[2370];
@(posedge clk);
#1;data_in = testData5[2371];
@(posedge clk);
#1;data_in = testData5[2372];
@(posedge clk);
#1;data_in = testData5[2373];
@(posedge clk);
#1;data_in = testData5[2374];
@(posedge clk);
#1;data_in = testData5[2375];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2376]; 
@(posedge clk);
#1;data_in = testData5[2377];
@(posedge clk);
#1;data_in = testData5[2378];
@(posedge clk);
#1;data_in = testData5[2379];
@(posedge clk);
#1;data_in = testData5[2380];
@(posedge clk);
#1;data_in = testData5[2381];
@(posedge clk);
#1;data_in = testData5[2382];
@(posedge clk);
#1;data_in = testData5[2383];
@(posedge clk);
#1;data_in = testData5[2384];
@(posedge clk);
#1;data_in = testData5[2385];
@(posedge clk);
#1;data_in = testData5[2386];
@(posedge clk);
#1;data_in = testData5[2387];
@(posedge clk);
#1;data_in = testData5[2388];
@(posedge clk);
#1;data_in = testData5[2389];
@(posedge clk);
#1;data_in = testData5[2390];
@(posedge clk);
#1;data_in = testData5[2391];
@(posedge clk);
#1;data_in = testData5[2392];
@(posedge clk);
#1;data_in = testData5[2393];
@(posedge clk);
#1;data_in = testData5[2394];
@(posedge clk);
#1;data_in = testData5[2395];
@(posedge clk);
#1;data_in = testData5[2396];
@(posedge clk);
#1;data_in = testData5[2397];
@(posedge clk);
#1;data_in = testData5[2398];
@(posedge clk);
#1;data_in = testData5[2399];
@(posedge clk);
#1;data_in = testData5[2400];
@(posedge clk);
#1;data_in = testData5[2401];
@(posedge clk);
#1;data_in = testData5[2402];
@(posedge clk);
#1;data_in = testData5[2403];
@(posedge clk);
#1;data_in = testData5[2404];
@(posedge clk);
#1;data_in = testData5[2405];
@(posedge clk);
#1;data_in = testData5[2406];
@(posedge clk);
#1;data_in = testData5[2407];
@(posedge clk);
#1;data_in = testData5[2408];
@(posedge clk);
#1;data_in = testData5[2409];
@(posedge clk);
#1;data_in = testData5[2410];
@(posedge clk);
#1;data_in = testData5[2411];
@(posedge clk);
#1;data_in = testData5[2412];
@(posedge clk);
#1;data_in = testData5[2413];
@(posedge clk);
#1;data_in = testData5[2414];
@(posedge clk);
#1;data_in = testData5[2415];
@(posedge clk);
#1;data_in = testData5[2416];
@(posedge clk);
#1;data_in = testData5[2417];
@(posedge clk);
#1;data_in = testData5[2418];
@(posedge clk);
#1;data_in = testData5[2419];
@(posedge clk);
#1;data_in = testData5[2420];
@(posedge clk);
#1;data_in = testData5[2421];
@(posedge clk);
#1;data_in = testData5[2422];
@(posedge clk);
#1;data_in = testData5[2423];
@(posedge clk);
#1;data_in = testData5[2424];
@(posedge clk);
#1;data_in = testData5[2425];
@(posedge clk);
#1;data_in = testData5[2426];
@(posedge clk);
#1;data_in = testData5[2427];
@(posedge clk);
#1;data_in = testData5[2428];
@(posedge clk);
#1;data_in = testData5[2429];
@(posedge clk);
#1;data_in = testData5[2430];
@(posedge clk);
#1;data_in = testData5[2431];
@(posedge clk);
#1;data_in = testData5[2432];
@(posedge clk);
#1;data_in = testData5[2433];
@(posedge clk);
#1;data_in = testData5[2434];
@(posedge clk);
#1;data_in = testData5[2435];
@(posedge clk);
#1;data_in = testData5[2436];
@(posedge clk);
#1;data_in = testData5[2437];
@(posedge clk);
#1;data_in = testData5[2438];
@(posedge clk);
#1;data_in = testData5[2439];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2440]; 
@(posedge clk);
#1;data_in = testData5[2441];
@(posedge clk);
#1;data_in = testData5[2442];
@(posedge clk);
#1;data_in = testData5[2443];
@(posedge clk);
#1;data_in = testData5[2444];
@(posedge clk);
#1;data_in = testData5[2445];
@(posedge clk);
#1;data_in = testData5[2446];
@(posedge clk);
#1;data_in = testData5[2447];
@(posedge clk);
#1;data_in = testData5[2448];
@(posedge clk);
#1;data_in = testData5[2449];
@(posedge clk);
#1;data_in = testData5[2450];
@(posedge clk);
#1;data_in = testData5[2451];
@(posedge clk);
#1;data_in = testData5[2452];
@(posedge clk);
#1;data_in = testData5[2453];
@(posedge clk);
#1;data_in = testData5[2454];
@(posedge clk);
#1;data_in = testData5[2455];
@(posedge clk);
#1;data_in = testData5[2456];
@(posedge clk);
#1;data_in = testData5[2457];
@(posedge clk);
#1;data_in = testData5[2458];
@(posedge clk);
#1;data_in = testData5[2459];
@(posedge clk);
#1;data_in = testData5[2460];
@(posedge clk);
#1;data_in = testData5[2461];
@(posedge clk);
#1;data_in = testData5[2462];
@(posedge clk);
#1;data_in = testData5[2463];
@(posedge clk);
#1;data_in = testData5[2464];
@(posedge clk);
#1;data_in = testData5[2465];
@(posedge clk);
#1;data_in = testData5[2466];
@(posedge clk);
#1;data_in = testData5[2467];
@(posedge clk);
#1;data_in = testData5[2468];
@(posedge clk);
#1;data_in = testData5[2469];
@(posedge clk);
#1;data_in = testData5[2470];
@(posedge clk);
#1;data_in = testData5[2471];
@(posedge clk);
#1;data_in = testData5[2472];
@(posedge clk);
#1;data_in = testData5[2473];
@(posedge clk);
#1;data_in = testData5[2474];
@(posedge clk);
#1;data_in = testData5[2475];
@(posedge clk);
#1;data_in = testData5[2476];
@(posedge clk);
#1;data_in = testData5[2477];
@(posedge clk);
#1;data_in = testData5[2478];
@(posedge clk);
#1;data_in = testData5[2479];
@(posedge clk);
#1;data_in = testData5[2480];
@(posedge clk);
#1;data_in = testData5[2481];
@(posedge clk);
#1;data_in = testData5[2482];
@(posedge clk);
#1;data_in = testData5[2483];
@(posedge clk);
#1;data_in = testData5[2484];
@(posedge clk);
#1;data_in = testData5[2485];
@(posedge clk);
#1;data_in = testData5[2486];
@(posedge clk);
#1;data_in = testData5[2487];
@(posedge clk);
#1;data_in = testData5[2488];
@(posedge clk);
#1;data_in = testData5[2489];
@(posedge clk);
#1;data_in = testData5[2490];
@(posedge clk);
#1;data_in = testData5[2491];
@(posedge clk);
#1;data_in = testData5[2492];
@(posedge clk);
#1;data_in = testData5[2493];
@(posedge clk);
#1;data_in = testData5[2494];
@(posedge clk);
#1;data_in = testData5[2495];
@(posedge clk);
#1;data_in = testData5[2496];
@(posedge clk);
#1;data_in = testData5[2497];
@(posedge clk);
#1;data_in = testData5[2498];
@(posedge clk);
#1;data_in = testData5[2499];
@(posedge clk);
#1;data_in = testData5[2500];
@(posedge clk);
#1;data_in = testData5[2501];
@(posedge clk);
#1;data_in = testData5[2502];
@(posedge clk);
#1;data_in = testData5[2503];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2504]; 
@(posedge clk);
#1;data_in = testData5[2505];
@(posedge clk);
#1;data_in = testData5[2506];
@(posedge clk);
#1;data_in = testData5[2507];
@(posedge clk);
#1;data_in = testData5[2508];
@(posedge clk);
#1;data_in = testData5[2509];
@(posedge clk);
#1;data_in = testData5[2510];
@(posedge clk);
#1;data_in = testData5[2511];
@(posedge clk);
#1;data_in = testData5[2512];
@(posedge clk);
#1;data_in = testData5[2513];
@(posedge clk);
#1;data_in = testData5[2514];
@(posedge clk);
#1;data_in = testData5[2515];
@(posedge clk);
#1;data_in = testData5[2516];
@(posedge clk);
#1;data_in = testData5[2517];
@(posedge clk);
#1;data_in = testData5[2518];
@(posedge clk);
#1;data_in = testData5[2519];
@(posedge clk);
#1;data_in = testData5[2520];
@(posedge clk);
#1;data_in = testData5[2521];
@(posedge clk);
#1;data_in = testData5[2522];
@(posedge clk);
#1;data_in = testData5[2523];
@(posedge clk);
#1;data_in = testData5[2524];
@(posedge clk);
#1;data_in = testData5[2525];
@(posedge clk);
#1;data_in = testData5[2526];
@(posedge clk);
#1;data_in = testData5[2527];
@(posedge clk);
#1;data_in = testData5[2528];
@(posedge clk);
#1;data_in = testData5[2529];
@(posedge clk);
#1;data_in = testData5[2530];
@(posedge clk);
#1;data_in = testData5[2531];
@(posedge clk);
#1;data_in = testData5[2532];
@(posedge clk);
#1;data_in = testData5[2533];
@(posedge clk);
#1;data_in = testData5[2534];
@(posedge clk);
#1;data_in = testData5[2535];
@(posedge clk);
#1;data_in = testData5[2536];
@(posedge clk);
#1;data_in = testData5[2537];
@(posedge clk);
#1;data_in = testData5[2538];
@(posedge clk);
#1;data_in = testData5[2539];
@(posedge clk);
#1;data_in = testData5[2540];
@(posedge clk);
#1;data_in = testData5[2541];
@(posedge clk);
#1;data_in = testData5[2542];
@(posedge clk);
#1;data_in = testData5[2543];
@(posedge clk);
#1;data_in = testData5[2544];
@(posedge clk);
#1;data_in = testData5[2545];
@(posedge clk);
#1;data_in = testData5[2546];
@(posedge clk);
#1;data_in = testData5[2547];
@(posedge clk);
#1;data_in = testData5[2548];
@(posedge clk);
#1;data_in = testData5[2549];
@(posedge clk);
#1;data_in = testData5[2550];
@(posedge clk);
#1;data_in = testData5[2551];
@(posedge clk);
#1;data_in = testData5[2552];
@(posedge clk);
#1;data_in = testData5[2553];
@(posedge clk);
#1;data_in = testData5[2554];
@(posedge clk);
#1;data_in = testData5[2555];
@(posedge clk);
#1;data_in = testData5[2556];
@(posedge clk);
#1;data_in = testData5[2557];
@(posedge clk);
#1;data_in = testData5[2558];
@(posedge clk);
#1;data_in = testData5[2559];
@(posedge clk);
#1;data_in = testData5[2560];
@(posedge clk);
#1;data_in = testData5[2561];
@(posedge clk);
#1;data_in = testData5[2562];
@(posedge clk);
#1;data_in = testData5[2563];
@(posedge clk);
#1;data_in = testData5[2564];
@(posedge clk);
#1;data_in = testData5[2565];
@(posedge clk);
#1;data_in = testData5[2566];
@(posedge clk);
#1;data_in = testData5[2567];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2568]; 
@(posedge clk);
#1;data_in = testData5[2569];
@(posedge clk);
#1;data_in = testData5[2570];
@(posedge clk);
#1;data_in = testData5[2571];
@(posedge clk);
#1;data_in = testData5[2572];
@(posedge clk);
#1;data_in = testData5[2573];
@(posedge clk);
#1;data_in = testData5[2574];
@(posedge clk);
#1;data_in = testData5[2575];
@(posedge clk);
#1;data_in = testData5[2576];
@(posedge clk);
#1;data_in = testData5[2577];
@(posedge clk);
#1;data_in = testData5[2578];
@(posedge clk);
#1;data_in = testData5[2579];
@(posedge clk);
#1;data_in = testData5[2580];
@(posedge clk);
#1;data_in = testData5[2581];
@(posedge clk);
#1;data_in = testData5[2582];
@(posedge clk);
#1;data_in = testData5[2583];
@(posedge clk);
#1;data_in = testData5[2584];
@(posedge clk);
#1;data_in = testData5[2585];
@(posedge clk);
#1;data_in = testData5[2586];
@(posedge clk);
#1;data_in = testData5[2587];
@(posedge clk);
#1;data_in = testData5[2588];
@(posedge clk);
#1;data_in = testData5[2589];
@(posedge clk);
#1;data_in = testData5[2590];
@(posedge clk);
#1;data_in = testData5[2591];
@(posedge clk);
#1;data_in = testData5[2592];
@(posedge clk);
#1;data_in = testData5[2593];
@(posedge clk);
#1;data_in = testData5[2594];
@(posedge clk);
#1;data_in = testData5[2595];
@(posedge clk);
#1;data_in = testData5[2596];
@(posedge clk);
#1;data_in = testData5[2597];
@(posedge clk);
#1;data_in = testData5[2598];
@(posedge clk);
#1;data_in = testData5[2599];
@(posedge clk);
#1;data_in = testData5[2600];
@(posedge clk);
#1;data_in = testData5[2601];
@(posedge clk);
#1;data_in = testData5[2602];
@(posedge clk);
#1;data_in = testData5[2603];
@(posedge clk);
#1;data_in = testData5[2604];
@(posedge clk);
#1;data_in = testData5[2605];
@(posedge clk);
#1;data_in = testData5[2606];
@(posedge clk);
#1;data_in = testData5[2607];
@(posedge clk);
#1;data_in = testData5[2608];
@(posedge clk);
#1;data_in = testData5[2609];
@(posedge clk);
#1;data_in = testData5[2610];
@(posedge clk);
#1;data_in = testData5[2611];
@(posedge clk);
#1;data_in = testData5[2612];
@(posedge clk);
#1;data_in = testData5[2613];
@(posedge clk);
#1;data_in = testData5[2614];
@(posedge clk);
#1;data_in = testData5[2615];
@(posedge clk);
#1;data_in = testData5[2616];
@(posedge clk);
#1;data_in = testData5[2617];
@(posedge clk);
#1;data_in = testData5[2618];
@(posedge clk);
#1;data_in = testData5[2619];
@(posedge clk);
#1;data_in = testData5[2620];
@(posedge clk);
#1;data_in = testData5[2621];
@(posedge clk);
#1;data_in = testData5[2622];
@(posedge clk);
#1;data_in = testData5[2623];
@(posedge clk);
#1;data_in = testData5[2624];
@(posedge clk);
#1;data_in = testData5[2625];
@(posedge clk);
#1;data_in = testData5[2626];
@(posedge clk);
#1;data_in = testData5[2627];
@(posedge clk);
#1;data_in = testData5[2628];
@(posedge clk);
#1;data_in = testData5[2629];
@(posedge clk);
#1;data_in = testData5[2630];
@(posedge clk);
#1;data_in = testData5[2631];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2632]; 
@(posedge clk);
#1;data_in = testData5[2633];
@(posedge clk);
#1;data_in = testData5[2634];
@(posedge clk);
#1;data_in = testData5[2635];
@(posedge clk);
#1;data_in = testData5[2636];
@(posedge clk);
#1;data_in = testData5[2637];
@(posedge clk);
#1;data_in = testData5[2638];
@(posedge clk);
#1;data_in = testData5[2639];
@(posedge clk);
#1;data_in = testData5[2640];
@(posedge clk);
#1;data_in = testData5[2641];
@(posedge clk);
#1;data_in = testData5[2642];
@(posedge clk);
#1;data_in = testData5[2643];
@(posedge clk);
#1;data_in = testData5[2644];
@(posedge clk);
#1;data_in = testData5[2645];
@(posedge clk);
#1;data_in = testData5[2646];
@(posedge clk);
#1;data_in = testData5[2647];
@(posedge clk);
#1;data_in = testData5[2648];
@(posedge clk);
#1;data_in = testData5[2649];
@(posedge clk);
#1;data_in = testData5[2650];
@(posedge clk);
#1;data_in = testData5[2651];
@(posedge clk);
#1;data_in = testData5[2652];
@(posedge clk);
#1;data_in = testData5[2653];
@(posedge clk);
#1;data_in = testData5[2654];
@(posedge clk);
#1;data_in = testData5[2655];
@(posedge clk);
#1;data_in = testData5[2656];
@(posedge clk);
#1;data_in = testData5[2657];
@(posedge clk);
#1;data_in = testData5[2658];
@(posedge clk);
#1;data_in = testData5[2659];
@(posedge clk);
#1;data_in = testData5[2660];
@(posedge clk);
#1;data_in = testData5[2661];
@(posedge clk);
#1;data_in = testData5[2662];
@(posedge clk);
#1;data_in = testData5[2663];
@(posedge clk);
#1;data_in = testData5[2664];
@(posedge clk);
#1;data_in = testData5[2665];
@(posedge clk);
#1;data_in = testData5[2666];
@(posedge clk);
#1;data_in = testData5[2667];
@(posedge clk);
#1;data_in = testData5[2668];
@(posedge clk);
#1;data_in = testData5[2669];
@(posedge clk);
#1;data_in = testData5[2670];
@(posedge clk);
#1;data_in = testData5[2671];
@(posedge clk);
#1;data_in = testData5[2672];
@(posedge clk);
#1;data_in = testData5[2673];
@(posedge clk);
#1;data_in = testData5[2674];
@(posedge clk);
#1;data_in = testData5[2675];
@(posedge clk);
#1;data_in = testData5[2676];
@(posedge clk);
#1;data_in = testData5[2677];
@(posedge clk);
#1;data_in = testData5[2678];
@(posedge clk);
#1;data_in = testData5[2679];
@(posedge clk);
#1;data_in = testData5[2680];
@(posedge clk);
#1;data_in = testData5[2681];
@(posedge clk);
#1;data_in = testData5[2682];
@(posedge clk);
#1;data_in = testData5[2683];
@(posedge clk);
#1;data_in = testData5[2684];
@(posedge clk);
#1;data_in = testData5[2685];
@(posedge clk);
#1;data_in = testData5[2686];
@(posedge clk);
#1;data_in = testData5[2687];
@(posedge clk);
#1;data_in = testData5[2688];
@(posedge clk);
#1;data_in = testData5[2689];
@(posedge clk);
#1;data_in = testData5[2690];
@(posedge clk);
#1;data_in = testData5[2691];
@(posedge clk);
#1;data_in = testData5[2692];
@(posedge clk);
#1;data_in = testData5[2693];
@(posedge clk);
#1;data_in = testData5[2694];
@(posedge clk);
#1;data_in = testData5[2695];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2696]; 
@(posedge clk);
#1;data_in = testData5[2697];
@(posedge clk);
#1;data_in = testData5[2698];
@(posedge clk);
#1;data_in = testData5[2699];
@(posedge clk);
#1;data_in = testData5[2700];
@(posedge clk);
#1;data_in = testData5[2701];
@(posedge clk);
#1;data_in = testData5[2702];
@(posedge clk);
#1;data_in = testData5[2703];
@(posedge clk);
#1;data_in = testData5[2704];
@(posedge clk);
#1;data_in = testData5[2705];
@(posedge clk);
#1;data_in = testData5[2706];
@(posedge clk);
#1;data_in = testData5[2707];
@(posedge clk);
#1;data_in = testData5[2708];
@(posedge clk);
#1;data_in = testData5[2709];
@(posedge clk);
#1;data_in = testData5[2710];
@(posedge clk);
#1;data_in = testData5[2711];
@(posedge clk);
#1;data_in = testData5[2712];
@(posedge clk);
#1;data_in = testData5[2713];
@(posedge clk);
#1;data_in = testData5[2714];
@(posedge clk);
#1;data_in = testData5[2715];
@(posedge clk);
#1;data_in = testData5[2716];
@(posedge clk);
#1;data_in = testData5[2717];
@(posedge clk);
#1;data_in = testData5[2718];
@(posedge clk);
#1;data_in = testData5[2719];
@(posedge clk);
#1;data_in = testData5[2720];
@(posedge clk);
#1;data_in = testData5[2721];
@(posedge clk);
#1;data_in = testData5[2722];
@(posedge clk);
#1;data_in = testData5[2723];
@(posedge clk);
#1;data_in = testData5[2724];
@(posedge clk);
#1;data_in = testData5[2725];
@(posedge clk);
#1;data_in = testData5[2726];
@(posedge clk);
#1;data_in = testData5[2727];
@(posedge clk);
#1;data_in = testData5[2728];
@(posedge clk);
#1;data_in = testData5[2729];
@(posedge clk);
#1;data_in = testData5[2730];
@(posedge clk);
#1;data_in = testData5[2731];
@(posedge clk);
#1;data_in = testData5[2732];
@(posedge clk);
#1;data_in = testData5[2733];
@(posedge clk);
#1;data_in = testData5[2734];
@(posedge clk);
#1;data_in = testData5[2735];
@(posedge clk);
#1;data_in = testData5[2736];
@(posedge clk);
#1;data_in = testData5[2737];
@(posedge clk);
#1;data_in = testData5[2738];
@(posedge clk);
#1;data_in = testData5[2739];
@(posedge clk);
#1;data_in = testData5[2740];
@(posedge clk);
#1;data_in = testData5[2741];
@(posedge clk);
#1;data_in = testData5[2742];
@(posedge clk);
#1;data_in = testData5[2743];
@(posedge clk);
#1;data_in = testData5[2744];
@(posedge clk);
#1;data_in = testData5[2745];
@(posedge clk);
#1;data_in = testData5[2746];
@(posedge clk);
#1;data_in = testData5[2747];
@(posedge clk);
#1;data_in = testData5[2748];
@(posedge clk);
#1;data_in = testData5[2749];
@(posedge clk);
#1;data_in = testData5[2750];
@(posedge clk);
#1;data_in = testData5[2751];
@(posedge clk);
#1;data_in = testData5[2752];
@(posedge clk);
#1;data_in = testData5[2753];
@(posedge clk);
#1;data_in = testData5[2754];
@(posedge clk);
#1;data_in = testData5[2755];
@(posedge clk);
#1;data_in = testData5[2756];
@(posedge clk);
#1;data_in = testData5[2757];
@(posedge clk);
#1;data_in = testData5[2758];
@(posedge clk);
#1;data_in = testData5[2759];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2760]; 
@(posedge clk);
#1;data_in = testData5[2761];
@(posedge clk);
#1;data_in = testData5[2762];
@(posedge clk);
#1;data_in = testData5[2763];
@(posedge clk);
#1;data_in = testData5[2764];
@(posedge clk);
#1;data_in = testData5[2765];
@(posedge clk);
#1;data_in = testData5[2766];
@(posedge clk);
#1;data_in = testData5[2767];
@(posedge clk);
#1;data_in = testData5[2768];
@(posedge clk);
#1;data_in = testData5[2769];
@(posedge clk);
#1;data_in = testData5[2770];
@(posedge clk);
#1;data_in = testData5[2771];
@(posedge clk);
#1;data_in = testData5[2772];
@(posedge clk);
#1;data_in = testData5[2773];
@(posedge clk);
#1;data_in = testData5[2774];
@(posedge clk);
#1;data_in = testData5[2775];
@(posedge clk);
#1;data_in = testData5[2776];
@(posedge clk);
#1;data_in = testData5[2777];
@(posedge clk);
#1;data_in = testData5[2778];
@(posedge clk);
#1;data_in = testData5[2779];
@(posedge clk);
#1;data_in = testData5[2780];
@(posedge clk);
#1;data_in = testData5[2781];
@(posedge clk);
#1;data_in = testData5[2782];
@(posedge clk);
#1;data_in = testData5[2783];
@(posedge clk);
#1;data_in = testData5[2784];
@(posedge clk);
#1;data_in = testData5[2785];
@(posedge clk);
#1;data_in = testData5[2786];
@(posedge clk);
#1;data_in = testData5[2787];
@(posedge clk);
#1;data_in = testData5[2788];
@(posedge clk);
#1;data_in = testData5[2789];
@(posedge clk);
#1;data_in = testData5[2790];
@(posedge clk);
#1;data_in = testData5[2791];
@(posedge clk);
#1;data_in = testData5[2792];
@(posedge clk);
#1;data_in = testData5[2793];
@(posedge clk);
#1;data_in = testData5[2794];
@(posedge clk);
#1;data_in = testData5[2795];
@(posedge clk);
#1;data_in = testData5[2796];
@(posedge clk);
#1;data_in = testData5[2797];
@(posedge clk);
#1;data_in = testData5[2798];
@(posedge clk);
#1;data_in = testData5[2799];
@(posedge clk);
#1;data_in = testData5[2800];
@(posedge clk);
#1;data_in = testData5[2801];
@(posedge clk);
#1;data_in = testData5[2802];
@(posedge clk);
#1;data_in = testData5[2803];
@(posedge clk);
#1;data_in = testData5[2804];
@(posedge clk);
#1;data_in = testData5[2805];
@(posedge clk);
#1;data_in = testData5[2806];
@(posedge clk);
#1;data_in = testData5[2807];
@(posedge clk);
#1;data_in = testData5[2808];
@(posedge clk);
#1;data_in = testData5[2809];
@(posedge clk);
#1;data_in = testData5[2810];
@(posedge clk);
#1;data_in = testData5[2811];
@(posedge clk);
#1;data_in = testData5[2812];
@(posedge clk);
#1;data_in = testData5[2813];
@(posedge clk);
#1;data_in = testData5[2814];
@(posedge clk);
#1;data_in = testData5[2815];
@(posedge clk);
#1;data_in = testData5[2816];
@(posedge clk);
#1;data_in = testData5[2817];
@(posedge clk);
#1;data_in = testData5[2818];
@(posedge clk);
#1;data_in = testData5[2819];
@(posedge clk);
#1;data_in = testData5[2820];
@(posedge clk);
#1;data_in = testData5[2821];
@(posedge clk);
#1;data_in = testData5[2822];
@(posedge clk);
#1;data_in = testData5[2823];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2824]; 
@(posedge clk);
#1;data_in = testData5[2825];
@(posedge clk);
#1;data_in = testData5[2826];
@(posedge clk);
#1;data_in = testData5[2827];
@(posedge clk);
#1;data_in = testData5[2828];
@(posedge clk);
#1;data_in = testData5[2829];
@(posedge clk);
#1;data_in = testData5[2830];
@(posedge clk);
#1;data_in = testData5[2831];
@(posedge clk);
#1;data_in = testData5[2832];
@(posedge clk);
#1;data_in = testData5[2833];
@(posedge clk);
#1;data_in = testData5[2834];
@(posedge clk);
#1;data_in = testData5[2835];
@(posedge clk);
#1;data_in = testData5[2836];
@(posedge clk);
#1;data_in = testData5[2837];
@(posedge clk);
#1;data_in = testData5[2838];
@(posedge clk);
#1;data_in = testData5[2839];
@(posedge clk);
#1;data_in = testData5[2840];
@(posedge clk);
#1;data_in = testData5[2841];
@(posedge clk);
#1;data_in = testData5[2842];
@(posedge clk);
#1;data_in = testData5[2843];
@(posedge clk);
#1;data_in = testData5[2844];
@(posedge clk);
#1;data_in = testData5[2845];
@(posedge clk);
#1;data_in = testData5[2846];
@(posedge clk);
#1;data_in = testData5[2847];
@(posedge clk);
#1;data_in = testData5[2848];
@(posedge clk);
#1;data_in = testData5[2849];
@(posedge clk);
#1;data_in = testData5[2850];
@(posedge clk);
#1;data_in = testData5[2851];
@(posedge clk);
#1;data_in = testData5[2852];
@(posedge clk);
#1;data_in = testData5[2853];
@(posedge clk);
#1;data_in = testData5[2854];
@(posedge clk);
#1;data_in = testData5[2855];
@(posedge clk);
#1;data_in = testData5[2856];
@(posedge clk);
#1;data_in = testData5[2857];
@(posedge clk);
#1;data_in = testData5[2858];
@(posedge clk);
#1;data_in = testData5[2859];
@(posedge clk);
#1;data_in = testData5[2860];
@(posedge clk);
#1;data_in = testData5[2861];
@(posedge clk);
#1;data_in = testData5[2862];
@(posedge clk);
#1;data_in = testData5[2863];
@(posedge clk);
#1;data_in = testData5[2864];
@(posedge clk);
#1;data_in = testData5[2865];
@(posedge clk);
#1;data_in = testData5[2866];
@(posedge clk);
#1;data_in = testData5[2867];
@(posedge clk);
#1;data_in = testData5[2868];
@(posedge clk);
#1;data_in = testData5[2869];
@(posedge clk);
#1;data_in = testData5[2870];
@(posedge clk);
#1;data_in = testData5[2871];
@(posedge clk);
#1;data_in = testData5[2872];
@(posedge clk);
#1;data_in = testData5[2873];
@(posedge clk);
#1;data_in = testData5[2874];
@(posedge clk);
#1;data_in = testData5[2875];
@(posedge clk);
#1;data_in = testData5[2876];
@(posedge clk);
#1;data_in = testData5[2877];
@(posedge clk);
#1;data_in = testData5[2878];
@(posedge clk);
#1;data_in = testData5[2879];
@(posedge clk);
#1;data_in = testData5[2880];
@(posedge clk);
#1;data_in = testData5[2881];
@(posedge clk);
#1;data_in = testData5[2882];
@(posedge clk);
#1;data_in = testData5[2883];
@(posedge clk);
#1;data_in = testData5[2884];
@(posedge clk);
#1;data_in = testData5[2885];
@(posedge clk);
#1;data_in = testData5[2886];
@(posedge clk);
#1;data_in = testData5[2887];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2888]; 
@(posedge clk);
#1;data_in = testData5[2889];
@(posedge clk);
#1;data_in = testData5[2890];
@(posedge clk);
#1;data_in = testData5[2891];
@(posedge clk);
#1;data_in = testData5[2892];
@(posedge clk);
#1;data_in = testData5[2893];
@(posedge clk);
#1;data_in = testData5[2894];
@(posedge clk);
#1;data_in = testData5[2895];
@(posedge clk);
#1;data_in = testData5[2896];
@(posedge clk);
#1;data_in = testData5[2897];
@(posedge clk);
#1;data_in = testData5[2898];
@(posedge clk);
#1;data_in = testData5[2899];
@(posedge clk);
#1;data_in = testData5[2900];
@(posedge clk);
#1;data_in = testData5[2901];
@(posedge clk);
#1;data_in = testData5[2902];
@(posedge clk);
#1;data_in = testData5[2903];
@(posedge clk);
#1;data_in = testData5[2904];
@(posedge clk);
#1;data_in = testData5[2905];
@(posedge clk);
#1;data_in = testData5[2906];
@(posedge clk);
#1;data_in = testData5[2907];
@(posedge clk);
#1;data_in = testData5[2908];
@(posedge clk);
#1;data_in = testData5[2909];
@(posedge clk);
#1;data_in = testData5[2910];
@(posedge clk);
#1;data_in = testData5[2911];
@(posedge clk);
#1;data_in = testData5[2912];
@(posedge clk);
#1;data_in = testData5[2913];
@(posedge clk);
#1;data_in = testData5[2914];
@(posedge clk);
#1;data_in = testData5[2915];
@(posedge clk);
#1;data_in = testData5[2916];
@(posedge clk);
#1;data_in = testData5[2917];
@(posedge clk);
#1;data_in = testData5[2918];
@(posedge clk);
#1;data_in = testData5[2919];
@(posedge clk);
#1;data_in = testData5[2920];
@(posedge clk);
#1;data_in = testData5[2921];
@(posedge clk);
#1;data_in = testData5[2922];
@(posedge clk);
#1;data_in = testData5[2923];
@(posedge clk);
#1;data_in = testData5[2924];
@(posedge clk);
#1;data_in = testData5[2925];
@(posedge clk);
#1;data_in = testData5[2926];
@(posedge clk);
#1;data_in = testData5[2927];
@(posedge clk);
#1;data_in = testData5[2928];
@(posedge clk);
#1;data_in = testData5[2929];
@(posedge clk);
#1;data_in = testData5[2930];
@(posedge clk);
#1;data_in = testData5[2931];
@(posedge clk);
#1;data_in = testData5[2932];
@(posedge clk);
#1;data_in = testData5[2933];
@(posedge clk);
#1;data_in = testData5[2934];
@(posedge clk);
#1;data_in = testData5[2935];
@(posedge clk);
#1;data_in = testData5[2936];
@(posedge clk);
#1;data_in = testData5[2937];
@(posedge clk);
#1;data_in = testData5[2938];
@(posedge clk);
#1;data_in = testData5[2939];
@(posedge clk);
#1;data_in = testData5[2940];
@(posedge clk);
#1;data_in = testData5[2941];
@(posedge clk);
#1;data_in = testData5[2942];
@(posedge clk);
#1;data_in = testData5[2943];
@(posedge clk);
#1;data_in = testData5[2944];
@(posedge clk);
#1;data_in = testData5[2945];
@(posedge clk);
#1;data_in = testData5[2946];
@(posedge clk);
#1;data_in = testData5[2947];
@(posedge clk);
#1;data_in = testData5[2948];
@(posedge clk);
#1;data_in = testData5[2949];
@(posedge clk);
#1;data_in = testData5[2950];
@(posedge clk);
#1;data_in = testData5[2951];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[2952]; 
@(posedge clk);
#1;data_in = testData5[2953];
@(posedge clk);
#1;data_in = testData5[2954];
@(posedge clk);
#1;data_in = testData5[2955];
@(posedge clk);
#1;data_in = testData5[2956];
@(posedge clk);
#1;data_in = testData5[2957];
@(posedge clk);
#1;data_in = testData5[2958];
@(posedge clk);
#1;data_in = testData5[2959];
@(posedge clk);
#1;data_in = testData5[2960];
@(posedge clk);
#1;data_in = testData5[2961];
@(posedge clk);
#1;data_in = testData5[2962];
@(posedge clk);
#1;data_in = testData5[2963];
@(posedge clk);
#1;data_in = testData5[2964];
@(posedge clk);
#1;data_in = testData5[2965];
@(posedge clk);
#1;data_in = testData5[2966];
@(posedge clk);
#1;data_in = testData5[2967];
@(posedge clk);
#1;data_in = testData5[2968];
@(posedge clk);
#1;data_in = testData5[2969];
@(posedge clk);
#1;data_in = testData5[2970];
@(posedge clk);
#1;data_in = testData5[2971];
@(posedge clk);
#1;data_in = testData5[2972];
@(posedge clk);
#1;data_in = testData5[2973];
@(posedge clk);
#1;data_in = testData5[2974];
@(posedge clk);
#1;data_in = testData5[2975];
@(posedge clk);
#1;data_in = testData5[2976];
@(posedge clk);
#1;data_in = testData5[2977];
@(posedge clk);
#1;data_in = testData5[2978];
@(posedge clk);
#1;data_in = testData5[2979];
@(posedge clk);
#1;data_in = testData5[2980];
@(posedge clk);
#1;data_in = testData5[2981];
@(posedge clk);
#1;data_in = testData5[2982];
@(posedge clk);
#1;data_in = testData5[2983];
@(posedge clk);
#1;data_in = testData5[2984];
@(posedge clk);
#1;data_in = testData5[2985];
@(posedge clk);
#1;data_in = testData5[2986];
@(posedge clk);
#1;data_in = testData5[2987];
@(posedge clk);
#1;data_in = testData5[2988];
@(posedge clk);
#1;data_in = testData5[2989];
@(posedge clk);
#1;data_in = testData5[2990];
@(posedge clk);
#1;data_in = testData5[2991];
@(posedge clk);
#1;data_in = testData5[2992];
@(posedge clk);
#1;data_in = testData5[2993];
@(posedge clk);
#1;data_in = testData5[2994];
@(posedge clk);
#1;data_in = testData5[2995];
@(posedge clk);
#1;data_in = testData5[2996];
@(posedge clk);
#1;data_in = testData5[2997];
@(posedge clk);
#1;data_in = testData5[2998];
@(posedge clk);
#1;data_in = testData5[2999];
@(posedge clk);
#1;data_in = testData5[3000];
@(posedge clk);
#1;data_in = testData5[3001];
@(posedge clk);
#1;data_in = testData5[3002];
@(posedge clk);
#1;data_in = testData5[3003];
@(posedge clk);
#1;data_in = testData5[3004];
@(posedge clk);
#1;data_in = testData5[3005];
@(posedge clk);
#1;data_in = testData5[3006];
@(posedge clk);
#1;data_in = testData5[3007];
@(posedge clk);
#1;data_in = testData5[3008];
@(posedge clk);
#1;data_in = testData5[3009];
@(posedge clk);
#1;data_in = testData5[3010];
@(posedge clk);
#1;data_in = testData5[3011];
@(posedge clk);
#1;data_in = testData5[3012];
@(posedge clk);
#1;data_in = testData5[3013];
@(posedge clk);
#1;data_in = testData5[3014];
@(posedge clk);
#1;data_in = testData5[3015];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[3016]; 
@(posedge clk);
#1;data_in = testData5[3017];
@(posedge clk);
#1;data_in = testData5[3018];
@(posedge clk);
#1;data_in = testData5[3019];
@(posedge clk);
#1;data_in = testData5[3020];
@(posedge clk);
#1;data_in = testData5[3021];
@(posedge clk);
#1;data_in = testData5[3022];
@(posedge clk);
#1;data_in = testData5[3023];
@(posedge clk);
#1;data_in = testData5[3024];
@(posedge clk);
#1;data_in = testData5[3025];
@(posedge clk);
#1;data_in = testData5[3026];
@(posedge clk);
#1;data_in = testData5[3027];
@(posedge clk);
#1;data_in = testData5[3028];
@(posedge clk);
#1;data_in = testData5[3029];
@(posedge clk);
#1;data_in = testData5[3030];
@(posedge clk);
#1;data_in = testData5[3031];
@(posedge clk);
#1;data_in = testData5[3032];
@(posedge clk);
#1;data_in = testData5[3033];
@(posedge clk);
#1;data_in = testData5[3034];
@(posedge clk);
#1;data_in = testData5[3035];
@(posedge clk);
#1;data_in = testData5[3036];
@(posedge clk);
#1;data_in = testData5[3037];
@(posedge clk);
#1;data_in = testData5[3038];
@(posedge clk);
#1;data_in = testData5[3039];
@(posedge clk);
#1;data_in = testData5[3040];
@(posedge clk);
#1;data_in = testData5[3041];
@(posedge clk);
#1;data_in = testData5[3042];
@(posedge clk);
#1;data_in = testData5[3043];
@(posedge clk);
#1;data_in = testData5[3044];
@(posedge clk);
#1;data_in = testData5[3045];
@(posedge clk);
#1;data_in = testData5[3046];
@(posedge clk);
#1;data_in = testData5[3047];
@(posedge clk);
#1;data_in = testData5[3048];
@(posedge clk);
#1;data_in = testData5[3049];
@(posedge clk);
#1;data_in = testData5[3050];
@(posedge clk);
#1;data_in = testData5[3051];
@(posedge clk);
#1;data_in = testData5[3052];
@(posedge clk);
#1;data_in = testData5[3053];
@(posedge clk);
#1;data_in = testData5[3054];
@(posedge clk);
#1;data_in = testData5[3055];
@(posedge clk);
#1;data_in = testData5[3056];
@(posedge clk);
#1;data_in = testData5[3057];
@(posedge clk);
#1;data_in = testData5[3058];
@(posedge clk);
#1;data_in = testData5[3059];
@(posedge clk);
#1;data_in = testData5[3060];
@(posedge clk);
#1;data_in = testData5[3061];
@(posedge clk);
#1;data_in = testData5[3062];
@(posedge clk);
#1;data_in = testData5[3063];
@(posedge clk);
#1;data_in = testData5[3064];
@(posedge clk);
#1;data_in = testData5[3065];
@(posedge clk);
#1;data_in = testData5[3066];
@(posedge clk);
#1;data_in = testData5[3067];
@(posedge clk);
#1;data_in = testData5[3068];
@(posedge clk);
#1;data_in = testData5[3069];
@(posedge clk);
#1;data_in = testData5[3070];
@(posedge clk);
#1;data_in = testData5[3071];
@(posedge clk);
#1;data_in = testData5[3072];
@(posedge clk);
#1;data_in = testData5[3073];
@(posedge clk);
#1;data_in = testData5[3074];
@(posedge clk);
#1;data_in = testData5[3075];
@(posedge clk);
#1;data_in = testData5[3076];
@(posedge clk);
#1;data_in = testData5[3077];
@(posedge clk);
#1;data_in = testData5[3078];
@(posedge clk);
#1;data_in = testData5[3079];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[3080]; 
@(posedge clk);
#1;data_in = testData5[3081];
@(posedge clk);
#1;data_in = testData5[3082];
@(posedge clk);
#1;data_in = testData5[3083];
@(posedge clk);
#1;data_in = testData5[3084];
@(posedge clk);
#1;data_in = testData5[3085];
@(posedge clk);
#1;data_in = testData5[3086];
@(posedge clk);
#1;data_in = testData5[3087];
@(posedge clk);
#1;data_in = testData5[3088];
@(posedge clk);
#1;data_in = testData5[3089];
@(posedge clk);
#1;data_in = testData5[3090];
@(posedge clk);
#1;data_in = testData5[3091];
@(posedge clk);
#1;data_in = testData5[3092];
@(posedge clk);
#1;data_in = testData5[3093];
@(posedge clk);
#1;data_in = testData5[3094];
@(posedge clk);
#1;data_in = testData5[3095];
@(posedge clk);
#1;data_in = testData5[3096];
@(posedge clk);
#1;data_in = testData5[3097];
@(posedge clk);
#1;data_in = testData5[3098];
@(posedge clk);
#1;data_in = testData5[3099];
@(posedge clk);
#1;data_in = testData5[3100];
@(posedge clk);
#1;data_in = testData5[3101];
@(posedge clk);
#1;data_in = testData5[3102];
@(posedge clk);
#1;data_in = testData5[3103];
@(posedge clk);
#1;data_in = testData5[3104];
@(posedge clk);
#1;data_in = testData5[3105];
@(posedge clk);
#1;data_in = testData5[3106];
@(posedge clk);
#1;data_in = testData5[3107];
@(posedge clk);
#1;data_in = testData5[3108];
@(posedge clk);
#1;data_in = testData5[3109];
@(posedge clk);
#1;data_in = testData5[3110];
@(posedge clk);
#1;data_in = testData5[3111];
@(posedge clk);
#1;data_in = testData5[3112];
@(posedge clk);
#1;data_in = testData5[3113];
@(posedge clk);
#1;data_in = testData5[3114];
@(posedge clk);
#1;data_in = testData5[3115];
@(posedge clk);
#1;data_in = testData5[3116];
@(posedge clk);
#1;data_in = testData5[3117];
@(posedge clk);
#1;data_in = testData5[3118];
@(posedge clk);
#1;data_in = testData5[3119];
@(posedge clk);
#1;data_in = testData5[3120];
@(posedge clk);
#1;data_in = testData5[3121];
@(posedge clk);
#1;data_in = testData5[3122];
@(posedge clk);
#1;data_in = testData5[3123];
@(posedge clk);
#1;data_in = testData5[3124];
@(posedge clk);
#1;data_in = testData5[3125];
@(posedge clk);
#1;data_in = testData5[3126];
@(posedge clk);
#1;data_in = testData5[3127];
@(posedge clk);
#1;data_in = testData5[3128];
@(posedge clk);
#1;data_in = testData5[3129];
@(posedge clk);
#1;data_in = testData5[3130];
@(posedge clk);
#1;data_in = testData5[3131];
@(posedge clk);
#1;data_in = testData5[3132];
@(posedge clk);
#1;data_in = testData5[3133];
@(posedge clk);
#1;data_in = testData5[3134];
@(posedge clk);
#1;data_in = testData5[3135];
@(posedge clk);
#1;data_in = testData5[3136];
@(posedge clk);
#1;data_in = testData5[3137];
@(posedge clk);
#1;data_in = testData5[3138];
@(posedge clk);
#1;data_in = testData5[3139];
@(posedge clk);
#1;data_in = testData5[3140];
@(posedge clk);
#1;data_in = testData5[3141];
@(posedge clk);
#1;data_in = testData5[3142];
@(posedge clk);
#1;data_in = testData5[3143];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[3144]; 
@(posedge clk);
#1;data_in = testData5[3145];
@(posedge clk);
#1;data_in = testData5[3146];
@(posedge clk);
#1;data_in = testData5[3147];
@(posedge clk);
#1;data_in = testData5[3148];
@(posedge clk);
#1;data_in = testData5[3149];
@(posedge clk);
#1;data_in = testData5[3150];
@(posedge clk);
#1;data_in = testData5[3151];
@(posedge clk);
#1;data_in = testData5[3152];
@(posedge clk);
#1;data_in = testData5[3153];
@(posedge clk);
#1;data_in = testData5[3154];
@(posedge clk);
#1;data_in = testData5[3155];
@(posedge clk);
#1;data_in = testData5[3156];
@(posedge clk);
#1;data_in = testData5[3157];
@(posedge clk);
#1;data_in = testData5[3158];
@(posedge clk);
#1;data_in = testData5[3159];
@(posedge clk);
#1;data_in = testData5[3160];
@(posedge clk);
#1;data_in = testData5[3161];
@(posedge clk);
#1;data_in = testData5[3162];
@(posedge clk);
#1;data_in = testData5[3163];
@(posedge clk);
#1;data_in = testData5[3164];
@(posedge clk);
#1;data_in = testData5[3165];
@(posedge clk);
#1;data_in = testData5[3166];
@(posedge clk);
#1;data_in = testData5[3167];
@(posedge clk);
#1;data_in = testData5[3168];
@(posedge clk);
#1;data_in = testData5[3169];
@(posedge clk);
#1;data_in = testData5[3170];
@(posedge clk);
#1;data_in = testData5[3171];
@(posedge clk);
#1;data_in = testData5[3172];
@(posedge clk);
#1;data_in = testData5[3173];
@(posedge clk);
#1;data_in = testData5[3174];
@(posedge clk);
#1;data_in = testData5[3175];
@(posedge clk);
#1;data_in = testData5[3176];
@(posedge clk);
#1;data_in = testData5[3177];
@(posedge clk);
#1;data_in = testData5[3178];
@(posedge clk);
#1;data_in = testData5[3179];
@(posedge clk);
#1;data_in = testData5[3180];
@(posedge clk);
#1;data_in = testData5[3181];
@(posedge clk);
#1;data_in = testData5[3182];
@(posedge clk);
#1;data_in = testData5[3183];
@(posedge clk);
#1;data_in = testData5[3184];
@(posedge clk);
#1;data_in = testData5[3185];
@(posedge clk);
#1;data_in = testData5[3186];
@(posedge clk);
#1;data_in = testData5[3187];
@(posedge clk);
#1;data_in = testData5[3188];
@(posedge clk);
#1;data_in = testData5[3189];
@(posedge clk);
#1;data_in = testData5[3190];
@(posedge clk);
#1;data_in = testData5[3191];
@(posedge clk);
#1;data_in = testData5[3192];
@(posedge clk);
#1;data_in = testData5[3193];
@(posedge clk);
#1;data_in = testData5[3194];
@(posedge clk);
#1;data_in = testData5[3195];
@(posedge clk);
#1;data_in = testData5[3196];
@(posedge clk);
#1;data_in = testData5[3197];
@(posedge clk);
#1;data_in = testData5[3198];
@(posedge clk);
#1;data_in = testData5[3199];
@(posedge clk);
#1;data_in = testData5[3200];
@(posedge clk);
#1;data_in = testData5[3201];
@(posedge clk);
#1;data_in = testData5[3202];
@(posedge clk);
#1;data_in = testData5[3203];
@(posedge clk);
#1;data_in = testData5[3204];
@(posedge clk);
#1;data_in = testData5[3205];
@(posedge clk);
#1;data_in = testData5[3206];
@(posedge clk);
#1;data_in = testData5[3207];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[3208]; 
@(posedge clk);
#1;data_in = testData5[3209];
@(posedge clk);
#1;data_in = testData5[3210];
@(posedge clk);
#1;data_in = testData5[3211];
@(posedge clk);
#1;data_in = testData5[3212];
@(posedge clk);
#1;data_in = testData5[3213];
@(posedge clk);
#1;data_in = testData5[3214];
@(posedge clk);
#1;data_in = testData5[3215];
@(posedge clk);
#1;data_in = testData5[3216];
@(posedge clk);
#1;data_in = testData5[3217];
@(posedge clk);
#1;data_in = testData5[3218];
@(posedge clk);
#1;data_in = testData5[3219];
@(posedge clk);
#1;data_in = testData5[3220];
@(posedge clk);
#1;data_in = testData5[3221];
@(posedge clk);
#1;data_in = testData5[3222];
@(posedge clk);
#1;data_in = testData5[3223];
@(posedge clk);
#1;data_in = testData5[3224];
@(posedge clk);
#1;data_in = testData5[3225];
@(posedge clk);
#1;data_in = testData5[3226];
@(posedge clk);
#1;data_in = testData5[3227];
@(posedge clk);
#1;data_in = testData5[3228];
@(posedge clk);
#1;data_in = testData5[3229];
@(posedge clk);
#1;data_in = testData5[3230];
@(posedge clk);
#1;data_in = testData5[3231];
@(posedge clk);
#1;data_in = testData5[3232];
@(posedge clk);
#1;data_in = testData5[3233];
@(posedge clk);
#1;data_in = testData5[3234];
@(posedge clk);
#1;data_in = testData5[3235];
@(posedge clk);
#1;data_in = testData5[3236];
@(posedge clk);
#1;data_in = testData5[3237];
@(posedge clk);
#1;data_in = testData5[3238];
@(posedge clk);
#1;data_in = testData5[3239];
@(posedge clk);
#1;data_in = testData5[3240];
@(posedge clk);
#1;data_in = testData5[3241];
@(posedge clk);
#1;data_in = testData5[3242];
@(posedge clk);
#1;data_in = testData5[3243];
@(posedge clk);
#1;data_in = testData5[3244];
@(posedge clk);
#1;data_in = testData5[3245];
@(posedge clk);
#1;data_in = testData5[3246];
@(posedge clk);
#1;data_in = testData5[3247];
@(posedge clk);
#1;data_in = testData5[3248];
@(posedge clk);
#1;data_in = testData5[3249];
@(posedge clk);
#1;data_in = testData5[3250];
@(posedge clk);
#1;data_in = testData5[3251];
@(posedge clk);
#1;data_in = testData5[3252];
@(posedge clk);
#1;data_in = testData5[3253];
@(posedge clk);
#1;data_in = testData5[3254];
@(posedge clk);
#1;data_in = testData5[3255];
@(posedge clk);
#1;data_in = testData5[3256];
@(posedge clk);
#1;data_in = testData5[3257];
@(posedge clk);
#1;data_in = testData5[3258];
@(posedge clk);
#1;data_in = testData5[3259];
@(posedge clk);
#1;data_in = testData5[3260];
@(posedge clk);
#1;data_in = testData5[3261];
@(posedge clk);
#1;data_in = testData5[3262];
@(posedge clk);
#1;data_in = testData5[3263];
@(posedge clk);
#1;data_in = testData5[3264];
@(posedge clk);
#1;data_in = testData5[3265];
@(posedge clk);
#1;data_in = testData5[3266];
@(posedge clk);
#1;data_in = testData5[3267];
@(posedge clk);
#1;data_in = testData5[3268];
@(posedge clk);
#1;data_in = testData5[3269];
@(posedge clk);
#1;data_in = testData5[3270];
@(posedge clk);
#1;data_in = testData5[3271];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[4] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[5] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[6] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[7] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
