
module memory_WIDTH8_SIZE32_LOGSIZE5_0 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n253), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n254), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n255), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n256), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n257), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n258), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n259), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n260), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n261), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n262), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n263), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n264), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n265), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n266), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n267), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n268), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n269), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n270), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n271), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n272), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n273), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n274), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n275), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n276), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n277), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n278), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n279), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n280), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n281), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n282), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n283), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n284), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n285), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n286), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n287), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n288), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n289), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n290), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n291), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n292), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n293), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n594), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n595), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n596), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n597), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n598), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n599), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n600), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n601), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n602), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n603), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n604), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n605), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n606), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n607), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n608), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n609), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n610), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n611), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n612), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n613), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n614), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n615), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n616), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n617), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n618), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n619), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n620), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n621), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n622), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n623), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n624), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n625), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n626), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n627), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n628), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n629), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n630), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n631), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n632), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n633), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n634), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n635), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n636), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n637), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n638), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n639), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n640), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n641), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n642), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n643), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n644), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n645), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n646), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n647), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n648), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n649), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n650), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n651), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n652), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n653), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n654), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n655), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n656), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n657), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n658), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n659), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n660), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n661), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n662), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n663), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n664), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n665), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n666), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n667), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n668), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n669), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n670), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n671), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n672), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n673), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n674), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n675), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n676), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n677), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n678), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n679), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n680), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n681), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n682), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n683), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n684), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n685), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n686), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n687), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n688), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n689), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n690), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n691), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n692), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n693), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n694), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n695), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n696), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n697), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n698), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n699), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n700), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n701), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n702), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n703), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n704), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n705), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n706), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n707), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n708), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n709), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n710), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n711), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n712), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n713), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n714), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n715), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n716), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n717), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n718), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n719), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n720), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n721), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n722), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n723), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n724), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n725), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n726), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n727), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n728), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n729), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n730), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n731), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n732), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n733), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n734), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n735), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n736), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n737), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n738), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n739), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n740), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n741), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n742), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n743), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n744), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n745), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n746), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n747), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n748), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n749), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n750), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n751), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n752), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n753), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n754), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n755), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n756), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n757), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n758), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n759), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n760), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n761), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n762), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n763), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n764), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n765), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n766), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n767), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n768), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n769), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n770), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n771), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n772), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n773), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n774), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n775), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n776), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n777), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n778), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n779), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n780), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n781), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n782), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n783), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n784), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n785), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n786), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n787), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n788), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n789), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n790), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n791), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n792), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n793), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n794), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n795), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n796), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n797), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n798), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n799), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n800), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n801), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n802), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n803), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n804), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n805), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n806), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n807), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n808), .CK(clk), .Q(\mem[0][0] ) );
  BUF_X1 U3 ( .A(n249), .Z(n247) );
  BUF_X1 U4 ( .A(N10), .Z(n248) );
  BUF_X1 U5 ( .A(n249), .Z(n245) );
  BUF_X1 U6 ( .A(n249), .Z(n246) );
  BUF_X1 U7 ( .A(N10), .Z(n249) );
  INV_X1 U8 ( .A(n326), .ZN(n840) );
  INV_X1 U9 ( .A(n337), .ZN(n839) );
  INV_X1 U10 ( .A(n347), .ZN(n838) );
  INV_X1 U11 ( .A(n357), .ZN(n837) );
  INV_X1 U12 ( .A(n367), .ZN(n836) );
  INV_X1 U13 ( .A(n377), .ZN(n835) );
  INV_X1 U14 ( .A(n386), .ZN(n834) );
  INV_X1 U15 ( .A(n395), .ZN(n833) );
  NOR3_X1 U16 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n334) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(n250), .ZN(n345) );
  NAND2_X1 U18 ( .A1(n335), .A2(n303), .ZN(n377) );
  NAND2_X1 U19 ( .A1(n334), .A2(n335), .ZN(n326) );
  NAND2_X1 U20 ( .A1(n345), .A2(n335), .ZN(n337) );
  NAND2_X1 U21 ( .A1(n355), .A2(n335), .ZN(n347) );
  NAND2_X1 U22 ( .A1(n365), .A2(n335), .ZN(n357) );
  NAND2_X1 U23 ( .A1(n375), .A2(n335), .ZN(n367) );
  NAND2_X1 U24 ( .A1(n335), .A2(n314), .ZN(n386) );
  NAND2_X1 U25 ( .A1(n335), .A2(n324), .ZN(n395) );
  INV_X1 U26 ( .A(n306), .ZN(n815) );
  INV_X1 U27 ( .A(n316), .ZN(n814) );
  INV_X1 U28 ( .A(n550), .ZN(n813) );
  INV_X1 U29 ( .A(n559), .ZN(n812) );
  INV_X1 U30 ( .A(n568), .ZN(n811) );
  INV_X1 U31 ( .A(n577), .ZN(n810) );
  INV_X1 U32 ( .A(n586), .ZN(n809) );
  INV_X1 U33 ( .A(n450), .ZN(n827) );
  INV_X1 U34 ( .A(n459), .ZN(n826) );
  INV_X1 U35 ( .A(n468), .ZN(n825) );
  INV_X1 U36 ( .A(n523), .ZN(n819) );
  INV_X1 U37 ( .A(n532), .ZN(n818) );
  INV_X1 U38 ( .A(n541), .ZN(n817) );
  INV_X1 U39 ( .A(n404), .ZN(n832) );
  INV_X1 U40 ( .A(n414), .ZN(n831) );
  INV_X1 U41 ( .A(n423), .ZN(n830) );
  INV_X1 U42 ( .A(n432), .ZN(n829) );
  INV_X1 U43 ( .A(n441), .ZN(n828) );
  INV_X1 U44 ( .A(n477), .ZN(n824) );
  INV_X1 U45 ( .A(n487), .ZN(n823) );
  INV_X1 U46 ( .A(n496), .ZN(n822) );
  INV_X1 U47 ( .A(n505), .ZN(n821) );
  INV_X1 U48 ( .A(n514), .ZN(n820) );
  INV_X1 U49 ( .A(n295), .ZN(n816) );
  BUF_X1 U50 ( .A(N11), .Z(n242) );
  BUF_X1 U51 ( .A(N11), .Z(n243) );
  BUF_X1 U52 ( .A(N11), .Z(n244) );
  INV_X1 U53 ( .A(N10), .ZN(n250) );
  BUF_X1 U54 ( .A(N12), .Z(n241) );
  NOR3_X1 U55 ( .A1(n252), .A2(N10), .A3(n251), .ZN(n314) );
  NOR3_X1 U56 ( .A1(n252), .A2(n250), .A3(n251), .ZN(n324) );
  NOR3_X1 U57 ( .A1(n250), .A2(N11), .A3(n252), .ZN(n303) );
  NOR3_X1 U58 ( .A1(N10), .A2(N12), .A3(n251), .ZN(n355) );
  NOR3_X1 U59 ( .A1(N10), .A2(N11), .A3(n252), .ZN(n375) );
  NAND2_X1 U60 ( .A1(n412), .A2(n303), .ZN(n450) );
  NAND2_X1 U61 ( .A1(n485), .A2(n303), .ZN(n523) );
  NAND2_X1 U62 ( .A1(n412), .A2(n375), .ZN(n441) );
  NAND2_X1 U63 ( .A1(n485), .A2(n375), .ZN(n514) );
  NAND2_X1 U64 ( .A1(n412), .A2(n334), .ZN(n404) );
  NAND2_X1 U65 ( .A1(n412), .A2(n345), .ZN(n414) );
  NAND2_X1 U66 ( .A1(n485), .A2(n334), .ZN(n477) );
  NAND2_X1 U67 ( .A1(n485), .A2(n345), .ZN(n487) );
  NAND2_X1 U68 ( .A1(n334), .A2(n304), .ZN(n550) );
  NAND2_X1 U69 ( .A1(n345), .A2(n304), .ZN(n559) );
  NAND2_X1 U70 ( .A1(n355), .A2(n304), .ZN(n568) );
  NAND2_X1 U71 ( .A1(n365), .A2(n304), .ZN(n577) );
  NAND2_X1 U72 ( .A1(n375), .A2(n304), .ZN(n586) );
  NAND2_X1 U73 ( .A1(n303), .A2(n304), .ZN(n295) );
  NAND2_X1 U74 ( .A1(n314), .A2(n304), .ZN(n306) );
  NAND2_X1 U75 ( .A1(n324), .A2(n304), .ZN(n316) );
  NAND2_X1 U76 ( .A1(n412), .A2(n355), .ZN(n423) );
  NAND2_X1 U77 ( .A1(n412), .A2(n365), .ZN(n432) );
  NAND2_X1 U78 ( .A1(n485), .A2(n355), .ZN(n496) );
  NAND2_X1 U79 ( .A1(n485), .A2(n365), .ZN(n505) );
  NAND2_X1 U80 ( .A1(n412), .A2(n314), .ZN(n459) );
  NAND2_X1 U81 ( .A1(n485), .A2(n314), .ZN(n532) );
  NAND2_X1 U82 ( .A1(n412), .A2(n324), .ZN(n468) );
  NAND2_X1 U83 ( .A1(n485), .A2(n324), .ZN(n541) );
  AND3_X1 U84 ( .A1(n841), .A2(n842), .A3(wr_en), .ZN(n335) );
  NOR3_X1 U85 ( .A1(n250), .A2(N12), .A3(n251), .ZN(n365) );
  AND3_X1 U86 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n304) );
  AND3_X1 U87 ( .A1(N13), .A2(n842), .A3(wr_en), .ZN(n412) );
  AND3_X1 U88 ( .A1(N14), .A2(n841), .A3(wr_en), .ZN(n485) );
  INV_X1 U89 ( .A(n376), .ZN(n768) );
  AOI22_X1 U90 ( .A1(data_in[0]), .A2(n835), .B1(n377), .B2(\mem[5][0] ), .ZN(
        n376) );
  INV_X1 U91 ( .A(n378), .ZN(n767) );
  AOI22_X1 U92 ( .A1(data_in[1]), .A2(n835), .B1(n377), .B2(\mem[5][1] ), .ZN(
        n378) );
  INV_X1 U93 ( .A(n379), .ZN(n766) );
  AOI22_X1 U94 ( .A1(data_in[2]), .A2(n835), .B1(n377), .B2(\mem[5][2] ), .ZN(
        n379) );
  INV_X1 U95 ( .A(n380), .ZN(n765) );
  AOI22_X1 U96 ( .A1(data_in[3]), .A2(n835), .B1(n377), .B2(\mem[5][3] ), .ZN(
        n380) );
  INV_X1 U97 ( .A(n381), .ZN(n764) );
  AOI22_X1 U98 ( .A1(data_in[4]), .A2(n835), .B1(n377), .B2(\mem[5][4] ), .ZN(
        n381) );
  INV_X1 U99 ( .A(n382), .ZN(n763) );
  AOI22_X1 U100 ( .A1(data_in[5]), .A2(n835), .B1(n377), .B2(\mem[5][5] ), 
        .ZN(n382) );
  INV_X1 U101 ( .A(n383), .ZN(n762) );
  AOI22_X1 U102 ( .A1(data_in[6]), .A2(n835), .B1(n377), .B2(\mem[5][6] ), 
        .ZN(n383) );
  INV_X1 U103 ( .A(n449), .ZN(n704) );
  AOI22_X1 U104 ( .A1(data_in[0]), .A2(n827), .B1(n450), .B2(\mem[13][0] ), 
        .ZN(n449) );
  INV_X1 U105 ( .A(n453), .ZN(n701) );
  AOI22_X1 U106 ( .A1(data_in[3]), .A2(n827), .B1(n450), .B2(\mem[13][3] ), 
        .ZN(n453) );
  INV_X1 U107 ( .A(n524), .ZN(n639) );
  AOI22_X1 U108 ( .A1(data_in[1]), .A2(n819), .B1(n523), .B2(\mem[21][1] ), 
        .ZN(n524) );
  INV_X1 U109 ( .A(n525), .ZN(n638) );
  AOI22_X1 U110 ( .A1(data_in[2]), .A2(n819), .B1(n523), .B2(\mem[21][2] ), 
        .ZN(n525) );
  INV_X1 U111 ( .A(n527), .ZN(n636) );
  AOI22_X1 U112 ( .A1(data_in[4]), .A2(n819), .B1(n523), .B2(\mem[21][4] ), 
        .ZN(n527) );
  INV_X1 U113 ( .A(n528), .ZN(n635) );
  AOI22_X1 U114 ( .A1(data_in[5]), .A2(n819), .B1(n523), .B2(\mem[21][5] ), 
        .ZN(n528) );
  INV_X1 U115 ( .A(n529), .ZN(n634) );
  AOI22_X1 U116 ( .A1(data_in[6]), .A2(n819), .B1(n523), .B2(\mem[21][6] ), 
        .ZN(n529) );
  INV_X1 U117 ( .A(n530), .ZN(n633) );
  AOI22_X1 U118 ( .A1(data_in[7]), .A2(n819), .B1(n523), .B2(\mem[21][7] ), 
        .ZN(n530) );
  INV_X1 U119 ( .A(n416), .ZN(n734) );
  AOI22_X1 U120 ( .A1(data_in[2]), .A2(n831), .B1(n414), .B2(\mem[9][2] ), 
        .ZN(n416) );
  INV_X1 U121 ( .A(n417), .ZN(n733) );
  AOI22_X1 U122 ( .A1(data_in[3]), .A2(n831), .B1(n414), .B2(\mem[9][3] ), 
        .ZN(n417) );
  INV_X1 U123 ( .A(n418), .ZN(n732) );
  AOI22_X1 U124 ( .A1(data_in[4]), .A2(n831), .B1(n414), .B2(\mem[9][4] ), 
        .ZN(n418) );
  INV_X1 U125 ( .A(n419), .ZN(n731) );
  AOI22_X1 U126 ( .A1(data_in[5]), .A2(n831), .B1(n414), .B2(\mem[9][5] ), 
        .ZN(n419) );
  INV_X1 U127 ( .A(n420), .ZN(n730) );
  AOI22_X1 U128 ( .A1(data_in[6]), .A2(n831), .B1(n414), .B2(\mem[9][6] ), 
        .ZN(n420) );
  INV_X1 U129 ( .A(n421), .ZN(n729) );
  AOI22_X1 U130 ( .A1(data_in[7]), .A2(n831), .B1(n414), .B2(\mem[9][7] ), 
        .ZN(n421) );
  INV_X1 U131 ( .A(n526), .ZN(n637) );
  AOI22_X1 U132 ( .A1(data_in[3]), .A2(n819), .B1(n523), .B2(\mem[21][3] ), 
        .ZN(n526) );
  INV_X1 U133 ( .A(n384), .ZN(n761) );
  AOI22_X1 U134 ( .A1(data_in[7]), .A2(n835), .B1(n377), .B2(\mem[5][7] ), 
        .ZN(n384) );
  INV_X1 U135 ( .A(n452), .ZN(n702) );
  AOI22_X1 U136 ( .A1(data_in[2]), .A2(n827), .B1(n450), .B2(\mem[13][2] ), 
        .ZN(n452) );
  INV_X1 U137 ( .A(n454), .ZN(n700) );
  AOI22_X1 U138 ( .A1(data_in[4]), .A2(n827), .B1(n450), .B2(\mem[13][4] ), 
        .ZN(n454) );
  INV_X1 U139 ( .A(n455), .ZN(n699) );
  AOI22_X1 U140 ( .A1(data_in[5]), .A2(n827), .B1(n450), .B2(\mem[13][5] ), 
        .ZN(n455) );
  INV_X1 U141 ( .A(n456), .ZN(n698) );
  AOI22_X1 U142 ( .A1(data_in[6]), .A2(n827), .B1(n450), .B2(\mem[13][6] ), 
        .ZN(n456) );
  INV_X1 U143 ( .A(n457), .ZN(n697) );
  AOI22_X1 U144 ( .A1(data_in[7]), .A2(n827), .B1(n450), .B2(\mem[13][7] ), 
        .ZN(n457) );
  INV_X1 U145 ( .A(n451), .ZN(n703) );
  AOI22_X1 U146 ( .A1(data_in[1]), .A2(n827), .B1(n450), .B2(\mem[13][1] ), 
        .ZN(n451) );
  INV_X1 U147 ( .A(n413), .ZN(n736) );
  AOI22_X1 U148 ( .A1(data_in[0]), .A2(n831), .B1(n414), .B2(\mem[9][0] ), 
        .ZN(n413) );
  INV_X1 U149 ( .A(n415), .ZN(n735) );
  AOI22_X1 U150 ( .A1(data_in[1]), .A2(n831), .B1(n414), .B2(\mem[9][1] ), 
        .ZN(n415) );
  INV_X1 U151 ( .A(n385), .ZN(n760) );
  AOI22_X1 U152 ( .A1(data_in[0]), .A2(n834), .B1(n386), .B2(\mem[6][0] ), 
        .ZN(n385) );
  INV_X1 U153 ( .A(n387), .ZN(n759) );
  AOI22_X1 U154 ( .A1(data_in[1]), .A2(n834), .B1(n386), .B2(\mem[6][1] ), 
        .ZN(n387) );
  INV_X1 U155 ( .A(n388), .ZN(n758) );
  AOI22_X1 U156 ( .A1(data_in[2]), .A2(n834), .B1(n386), .B2(\mem[6][2] ), 
        .ZN(n388) );
  INV_X1 U157 ( .A(n389), .ZN(n757) );
  AOI22_X1 U158 ( .A1(data_in[3]), .A2(n834), .B1(n386), .B2(\mem[6][3] ), 
        .ZN(n389) );
  INV_X1 U159 ( .A(n390), .ZN(n756) );
  AOI22_X1 U160 ( .A1(data_in[4]), .A2(n834), .B1(n386), .B2(\mem[6][4] ), 
        .ZN(n390) );
  INV_X1 U161 ( .A(n391), .ZN(n755) );
  AOI22_X1 U162 ( .A1(data_in[5]), .A2(n834), .B1(n386), .B2(\mem[6][5] ), 
        .ZN(n391) );
  INV_X1 U163 ( .A(n392), .ZN(n754) );
  AOI22_X1 U164 ( .A1(data_in[6]), .A2(n834), .B1(n386), .B2(\mem[6][6] ), 
        .ZN(n392) );
  INV_X1 U165 ( .A(n393), .ZN(n753) );
  AOI22_X1 U166 ( .A1(data_in[7]), .A2(n834), .B1(n386), .B2(\mem[6][7] ), 
        .ZN(n393) );
  INV_X1 U167 ( .A(n394), .ZN(n752) );
  AOI22_X1 U168 ( .A1(data_in[0]), .A2(n833), .B1(n395), .B2(\mem[7][0] ), 
        .ZN(n394) );
  INV_X1 U169 ( .A(n396), .ZN(n751) );
  AOI22_X1 U170 ( .A1(data_in[1]), .A2(n833), .B1(n395), .B2(\mem[7][1] ), 
        .ZN(n396) );
  INV_X1 U171 ( .A(n397), .ZN(n750) );
  AOI22_X1 U172 ( .A1(data_in[2]), .A2(n833), .B1(n395), .B2(\mem[7][2] ), 
        .ZN(n397) );
  INV_X1 U173 ( .A(n398), .ZN(n749) );
  AOI22_X1 U174 ( .A1(data_in[3]), .A2(n833), .B1(n395), .B2(\mem[7][3] ), 
        .ZN(n398) );
  INV_X1 U175 ( .A(n399), .ZN(n748) );
  AOI22_X1 U176 ( .A1(data_in[4]), .A2(n833), .B1(n395), .B2(\mem[7][4] ), 
        .ZN(n399) );
  INV_X1 U177 ( .A(n400), .ZN(n747) );
  AOI22_X1 U178 ( .A1(data_in[5]), .A2(n833), .B1(n395), .B2(\mem[7][5] ), 
        .ZN(n400) );
  INV_X1 U179 ( .A(n401), .ZN(n746) );
  AOI22_X1 U180 ( .A1(data_in[6]), .A2(n833), .B1(n395), .B2(\mem[7][6] ), 
        .ZN(n401) );
  INV_X1 U181 ( .A(n402), .ZN(n745) );
  AOI22_X1 U182 ( .A1(data_in[7]), .A2(n833), .B1(n395), .B2(\mem[7][7] ), 
        .ZN(n402) );
  INV_X1 U183 ( .A(n422), .ZN(n728) );
  AOI22_X1 U184 ( .A1(data_in[0]), .A2(n830), .B1(n423), .B2(\mem[10][0] ), 
        .ZN(n422) );
  INV_X1 U185 ( .A(n424), .ZN(n727) );
  AOI22_X1 U186 ( .A1(data_in[1]), .A2(n830), .B1(n423), .B2(\mem[10][1] ), 
        .ZN(n424) );
  INV_X1 U187 ( .A(n425), .ZN(n726) );
  AOI22_X1 U188 ( .A1(data_in[2]), .A2(n830), .B1(n423), .B2(\mem[10][2] ), 
        .ZN(n425) );
  INV_X1 U189 ( .A(n426), .ZN(n725) );
  AOI22_X1 U190 ( .A1(data_in[3]), .A2(n830), .B1(n423), .B2(\mem[10][3] ), 
        .ZN(n426) );
  INV_X1 U191 ( .A(n427), .ZN(n724) );
  AOI22_X1 U192 ( .A1(data_in[4]), .A2(n830), .B1(n423), .B2(\mem[10][4] ), 
        .ZN(n427) );
  INV_X1 U193 ( .A(n428), .ZN(n723) );
  AOI22_X1 U194 ( .A1(data_in[5]), .A2(n830), .B1(n423), .B2(\mem[10][5] ), 
        .ZN(n428) );
  INV_X1 U195 ( .A(n429), .ZN(n722) );
  AOI22_X1 U196 ( .A1(data_in[6]), .A2(n830), .B1(n423), .B2(\mem[10][6] ), 
        .ZN(n429) );
  INV_X1 U197 ( .A(n430), .ZN(n721) );
  AOI22_X1 U198 ( .A1(data_in[7]), .A2(n830), .B1(n423), .B2(\mem[10][7] ), 
        .ZN(n430) );
  INV_X1 U199 ( .A(n431), .ZN(n720) );
  AOI22_X1 U200 ( .A1(data_in[0]), .A2(n829), .B1(n432), .B2(\mem[11][0] ), 
        .ZN(n431) );
  INV_X1 U201 ( .A(n433), .ZN(n719) );
  AOI22_X1 U202 ( .A1(data_in[1]), .A2(n829), .B1(n432), .B2(\mem[11][1] ), 
        .ZN(n433) );
  INV_X1 U203 ( .A(n434), .ZN(n718) );
  AOI22_X1 U204 ( .A1(data_in[2]), .A2(n829), .B1(n432), .B2(\mem[11][2] ), 
        .ZN(n434) );
  INV_X1 U205 ( .A(n435), .ZN(n717) );
  AOI22_X1 U206 ( .A1(data_in[3]), .A2(n829), .B1(n432), .B2(\mem[11][3] ), 
        .ZN(n435) );
  INV_X1 U207 ( .A(n436), .ZN(n716) );
  AOI22_X1 U208 ( .A1(data_in[4]), .A2(n829), .B1(n432), .B2(\mem[11][4] ), 
        .ZN(n436) );
  INV_X1 U209 ( .A(n437), .ZN(n715) );
  AOI22_X1 U210 ( .A1(data_in[5]), .A2(n829), .B1(n432), .B2(\mem[11][5] ), 
        .ZN(n437) );
  INV_X1 U211 ( .A(n438), .ZN(n714) );
  AOI22_X1 U212 ( .A1(data_in[6]), .A2(n829), .B1(n432), .B2(\mem[11][6] ), 
        .ZN(n438) );
  INV_X1 U213 ( .A(n486), .ZN(n672) );
  AOI22_X1 U214 ( .A1(data_in[0]), .A2(n823), .B1(n487), .B2(\mem[17][0] ), 
        .ZN(n486) );
  INV_X1 U215 ( .A(n490), .ZN(n669) );
  AOI22_X1 U216 ( .A1(data_in[3]), .A2(n823), .B1(n487), .B2(\mem[17][3] ), 
        .ZN(n490) );
  INV_X1 U217 ( .A(n522), .ZN(n640) );
  AOI22_X1 U218 ( .A1(data_in[0]), .A2(n819), .B1(n523), .B2(\mem[21][0] ), 
        .ZN(n522) );
  INV_X1 U219 ( .A(n439), .ZN(n713) );
  AOI22_X1 U220 ( .A1(data_in[7]), .A2(n829), .B1(n432), .B2(\mem[11][7] ), 
        .ZN(n439) );
  INV_X1 U221 ( .A(n488), .ZN(n671) );
  AOI22_X1 U222 ( .A1(data_in[1]), .A2(n823), .B1(n487), .B2(\mem[17][1] ), 
        .ZN(n488) );
  INV_X1 U223 ( .A(n489), .ZN(n670) );
  AOI22_X1 U224 ( .A1(data_in[2]), .A2(n823), .B1(n487), .B2(\mem[17][2] ), 
        .ZN(n489) );
  INV_X1 U225 ( .A(n491), .ZN(n668) );
  AOI22_X1 U226 ( .A1(data_in[4]), .A2(n823), .B1(n487), .B2(\mem[17][4] ), 
        .ZN(n491) );
  INV_X1 U227 ( .A(n492), .ZN(n667) );
  AOI22_X1 U228 ( .A1(data_in[5]), .A2(n823), .B1(n487), .B2(\mem[17][5] ), 
        .ZN(n492) );
  INV_X1 U229 ( .A(n493), .ZN(n666) );
  AOI22_X1 U230 ( .A1(data_in[6]), .A2(n823), .B1(n487), .B2(\mem[17][6] ), 
        .ZN(n493) );
  INV_X1 U231 ( .A(n494), .ZN(n665) );
  AOI22_X1 U232 ( .A1(data_in[7]), .A2(n823), .B1(n487), .B2(\mem[17][7] ), 
        .ZN(n494) );
  INV_X1 U233 ( .A(n458), .ZN(n696) );
  AOI22_X1 U234 ( .A1(data_in[0]), .A2(n826), .B1(n459), .B2(\mem[14][0] ), 
        .ZN(n458) );
  INV_X1 U235 ( .A(n460), .ZN(n695) );
  AOI22_X1 U236 ( .A1(data_in[1]), .A2(n826), .B1(n459), .B2(\mem[14][1] ), 
        .ZN(n460) );
  INV_X1 U237 ( .A(n461), .ZN(n694) );
  AOI22_X1 U238 ( .A1(data_in[2]), .A2(n826), .B1(n459), .B2(\mem[14][2] ), 
        .ZN(n461) );
  INV_X1 U239 ( .A(n462), .ZN(n693) );
  AOI22_X1 U240 ( .A1(data_in[3]), .A2(n826), .B1(n459), .B2(\mem[14][3] ), 
        .ZN(n462) );
  INV_X1 U241 ( .A(n463), .ZN(n692) );
  AOI22_X1 U242 ( .A1(data_in[4]), .A2(n826), .B1(n459), .B2(\mem[14][4] ), 
        .ZN(n463) );
  INV_X1 U243 ( .A(n464), .ZN(n691) );
  AOI22_X1 U244 ( .A1(data_in[5]), .A2(n826), .B1(n459), .B2(\mem[14][5] ), 
        .ZN(n464) );
  INV_X1 U245 ( .A(n465), .ZN(n690) );
  AOI22_X1 U246 ( .A1(data_in[6]), .A2(n826), .B1(n459), .B2(\mem[14][6] ), 
        .ZN(n465) );
  INV_X1 U247 ( .A(n466), .ZN(n689) );
  AOI22_X1 U248 ( .A1(data_in[7]), .A2(n826), .B1(n459), .B2(\mem[14][7] ), 
        .ZN(n466) );
  INV_X1 U249 ( .A(n467), .ZN(n688) );
  AOI22_X1 U250 ( .A1(data_in[0]), .A2(n825), .B1(n468), .B2(\mem[15][0] ), 
        .ZN(n467) );
  INV_X1 U251 ( .A(n469), .ZN(n687) );
  AOI22_X1 U252 ( .A1(data_in[1]), .A2(n825), .B1(n468), .B2(\mem[15][1] ), 
        .ZN(n469) );
  INV_X1 U253 ( .A(n470), .ZN(n686) );
  AOI22_X1 U254 ( .A1(data_in[2]), .A2(n825), .B1(n468), .B2(\mem[15][2] ), 
        .ZN(n470) );
  INV_X1 U255 ( .A(n471), .ZN(n685) );
  AOI22_X1 U256 ( .A1(data_in[3]), .A2(n825), .B1(n468), .B2(\mem[15][3] ), 
        .ZN(n471) );
  INV_X1 U257 ( .A(n472), .ZN(n684) );
  AOI22_X1 U258 ( .A1(data_in[4]), .A2(n825), .B1(n468), .B2(\mem[15][4] ), 
        .ZN(n472) );
  INV_X1 U259 ( .A(n473), .ZN(n683) );
  AOI22_X1 U260 ( .A1(data_in[5]), .A2(n825), .B1(n468), .B2(\mem[15][5] ), 
        .ZN(n473) );
  INV_X1 U261 ( .A(n474), .ZN(n682) );
  AOI22_X1 U262 ( .A1(data_in[6]), .A2(n825), .B1(n468), .B2(\mem[15][6] ), 
        .ZN(n474) );
  INV_X1 U263 ( .A(n475), .ZN(n681) );
  AOI22_X1 U264 ( .A1(data_in[7]), .A2(n825), .B1(n468), .B2(\mem[15][7] ), 
        .ZN(n475) );
  INV_X1 U265 ( .A(n495), .ZN(n664) );
  AOI22_X1 U266 ( .A1(data_in[0]), .A2(n822), .B1(n496), .B2(\mem[18][0] ), 
        .ZN(n495) );
  INV_X1 U267 ( .A(n497), .ZN(n663) );
  AOI22_X1 U268 ( .A1(data_in[1]), .A2(n822), .B1(n496), .B2(\mem[18][1] ), 
        .ZN(n497) );
  INV_X1 U269 ( .A(n498), .ZN(n662) );
  AOI22_X1 U270 ( .A1(data_in[2]), .A2(n822), .B1(n496), .B2(\mem[18][2] ), 
        .ZN(n498) );
  INV_X1 U271 ( .A(n499), .ZN(n661) );
  AOI22_X1 U272 ( .A1(data_in[3]), .A2(n822), .B1(n496), .B2(\mem[18][3] ), 
        .ZN(n499) );
  INV_X1 U273 ( .A(n500), .ZN(n660) );
  AOI22_X1 U274 ( .A1(data_in[4]), .A2(n822), .B1(n496), .B2(\mem[18][4] ), 
        .ZN(n500) );
  INV_X1 U275 ( .A(n501), .ZN(n659) );
  AOI22_X1 U276 ( .A1(data_in[5]), .A2(n822), .B1(n496), .B2(\mem[18][5] ), 
        .ZN(n501) );
  INV_X1 U277 ( .A(n502), .ZN(n658) );
  AOI22_X1 U278 ( .A1(data_in[6]), .A2(n822), .B1(n496), .B2(\mem[18][6] ), 
        .ZN(n502) );
  INV_X1 U279 ( .A(n503), .ZN(n657) );
  AOI22_X1 U280 ( .A1(data_in[7]), .A2(n822), .B1(n496), .B2(\mem[18][7] ), 
        .ZN(n503) );
  INV_X1 U281 ( .A(n504), .ZN(n656) );
  AOI22_X1 U282 ( .A1(data_in[0]), .A2(n821), .B1(n505), .B2(\mem[19][0] ), 
        .ZN(n504) );
  INV_X1 U283 ( .A(n506), .ZN(n655) );
  AOI22_X1 U284 ( .A1(data_in[1]), .A2(n821), .B1(n505), .B2(\mem[19][1] ), 
        .ZN(n506) );
  INV_X1 U285 ( .A(n507), .ZN(n654) );
  AOI22_X1 U286 ( .A1(data_in[2]), .A2(n821), .B1(n505), .B2(\mem[19][2] ), 
        .ZN(n507) );
  INV_X1 U287 ( .A(n508), .ZN(n653) );
  AOI22_X1 U288 ( .A1(data_in[3]), .A2(n821), .B1(n505), .B2(\mem[19][3] ), 
        .ZN(n508) );
  INV_X1 U289 ( .A(n509), .ZN(n652) );
  AOI22_X1 U290 ( .A1(data_in[4]), .A2(n821), .B1(n505), .B2(\mem[19][4] ), 
        .ZN(n509) );
  INV_X1 U291 ( .A(n510), .ZN(n651) );
  AOI22_X1 U292 ( .A1(data_in[5]), .A2(n821), .B1(n505), .B2(\mem[19][5] ), 
        .ZN(n510) );
  INV_X1 U293 ( .A(n511), .ZN(n650) );
  AOI22_X1 U294 ( .A1(data_in[6]), .A2(n821), .B1(n505), .B2(\mem[19][6] ), 
        .ZN(n511) );
  INV_X1 U295 ( .A(n512), .ZN(n649) );
  AOI22_X1 U296 ( .A1(data_in[7]), .A2(n821), .B1(n505), .B2(\mem[19][7] ), 
        .ZN(n512) );
  INV_X1 U297 ( .A(n531), .ZN(n632) );
  AOI22_X1 U298 ( .A1(data_in[0]), .A2(n818), .B1(n532), .B2(\mem[22][0] ), 
        .ZN(n531) );
  INV_X1 U299 ( .A(n533), .ZN(n631) );
  AOI22_X1 U300 ( .A1(data_in[1]), .A2(n818), .B1(n532), .B2(\mem[22][1] ), 
        .ZN(n533) );
  INV_X1 U301 ( .A(n534), .ZN(n630) );
  AOI22_X1 U302 ( .A1(data_in[2]), .A2(n818), .B1(n532), .B2(\mem[22][2] ), 
        .ZN(n534) );
  INV_X1 U303 ( .A(n535), .ZN(n629) );
  AOI22_X1 U304 ( .A1(data_in[3]), .A2(n818), .B1(n532), .B2(\mem[22][3] ), 
        .ZN(n535) );
  INV_X1 U305 ( .A(n536), .ZN(n628) );
  AOI22_X1 U306 ( .A1(data_in[4]), .A2(n818), .B1(n532), .B2(\mem[22][4] ), 
        .ZN(n536) );
  INV_X1 U307 ( .A(n537), .ZN(n627) );
  AOI22_X1 U308 ( .A1(data_in[5]), .A2(n818), .B1(n532), .B2(\mem[22][5] ), 
        .ZN(n537) );
  INV_X1 U309 ( .A(n538), .ZN(n626) );
  AOI22_X1 U310 ( .A1(data_in[6]), .A2(n818), .B1(n532), .B2(\mem[22][6] ), 
        .ZN(n538) );
  INV_X1 U311 ( .A(n539), .ZN(n625) );
  AOI22_X1 U312 ( .A1(data_in[7]), .A2(n818), .B1(n532), .B2(\mem[22][7] ), 
        .ZN(n539) );
  INV_X1 U313 ( .A(n540), .ZN(n624) );
  AOI22_X1 U314 ( .A1(data_in[0]), .A2(n817), .B1(n541), .B2(\mem[23][0] ), 
        .ZN(n540) );
  INV_X1 U315 ( .A(n542), .ZN(n623) );
  AOI22_X1 U316 ( .A1(data_in[1]), .A2(n817), .B1(n541), .B2(\mem[23][1] ), 
        .ZN(n542) );
  INV_X1 U317 ( .A(n543), .ZN(n622) );
  AOI22_X1 U318 ( .A1(data_in[2]), .A2(n817), .B1(n541), .B2(\mem[23][2] ), 
        .ZN(n543) );
  INV_X1 U319 ( .A(n544), .ZN(n621) );
  AOI22_X1 U320 ( .A1(data_in[3]), .A2(n817), .B1(n541), .B2(\mem[23][3] ), 
        .ZN(n544) );
  INV_X1 U321 ( .A(n545), .ZN(n620) );
  AOI22_X1 U322 ( .A1(data_in[4]), .A2(n817), .B1(n541), .B2(\mem[23][4] ), 
        .ZN(n545) );
  INV_X1 U323 ( .A(n546), .ZN(n619) );
  AOI22_X1 U324 ( .A1(data_in[5]), .A2(n817), .B1(n541), .B2(\mem[23][5] ), 
        .ZN(n546) );
  INV_X1 U325 ( .A(n547), .ZN(n618) );
  AOI22_X1 U326 ( .A1(data_in[6]), .A2(n817), .B1(n541), .B2(\mem[23][6] ), 
        .ZN(n547) );
  INV_X1 U327 ( .A(n548), .ZN(n617) );
  AOI22_X1 U328 ( .A1(data_in[7]), .A2(n817), .B1(n541), .B2(\mem[23][7] ), 
        .ZN(n548) );
  INV_X1 U329 ( .A(N11), .ZN(n251) );
  INV_X1 U330 ( .A(n440), .ZN(n712) );
  AOI22_X1 U331 ( .A1(data_in[0]), .A2(n828), .B1(n441), .B2(\mem[12][0] ), 
        .ZN(n440) );
  INV_X1 U332 ( .A(n442), .ZN(n711) );
  AOI22_X1 U333 ( .A1(data_in[1]), .A2(n828), .B1(n441), .B2(\mem[12][1] ), 
        .ZN(n442) );
  INV_X1 U334 ( .A(n443), .ZN(n710) );
  AOI22_X1 U335 ( .A1(data_in[2]), .A2(n828), .B1(n441), .B2(\mem[12][2] ), 
        .ZN(n443) );
  INV_X1 U336 ( .A(n444), .ZN(n709) );
  AOI22_X1 U337 ( .A1(data_in[3]), .A2(n828), .B1(n441), .B2(\mem[12][3] ), 
        .ZN(n444) );
  INV_X1 U338 ( .A(n445), .ZN(n708) );
  AOI22_X1 U339 ( .A1(data_in[4]), .A2(n828), .B1(n441), .B2(\mem[12][4] ), 
        .ZN(n445) );
  INV_X1 U340 ( .A(n446), .ZN(n707) );
  AOI22_X1 U341 ( .A1(data_in[5]), .A2(n828), .B1(n441), .B2(\mem[12][5] ), 
        .ZN(n446) );
  INV_X1 U342 ( .A(n447), .ZN(n706) );
  AOI22_X1 U343 ( .A1(data_in[6]), .A2(n828), .B1(n441), .B2(\mem[12][6] ), 
        .ZN(n447) );
  INV_X1 U344 ( .A(n448), .ZN(n705) );
  AOI22_X1 U345 ( .A1(data_in[7]), .A2(n828), .B1(n441), .B2(\mem[12][7] ), 
        .ZN(n448) );
  INV_X1 U346 ( .A(n513), .ZN(n648) );
  AOI22_X1 U347 ( .A1(data_in[0]), .A2(n820), .B1(n514), .B2(\mem[20][0] ), 
        .ZN(n513) );
  INV_X1 U348 ( .A(n515), .ZN(n647) );
  AOI22_X1 U349 ( .A1(data_in[1]), .A2(n820), .B1(n514), .B2(\mem[20][1] ), 
        .ZN(n515) );
  INV_X1 U350 ( .A(n516), .ZN(n646) );
  AOI22_X1 U351 ( .A1(data_in[2]), .A2(n820), .B1(n514), .B2(\mem[20][2] ), 
        .ZN(n516) );
  INV_X1 U352 ( .A(n517), .ZN(n645) );
  AOI22_X1 U353 ( .A1(data_in[3]), .A2(n820), .B1(n514), .B2(\mem[20][3] ), 
        .ZN(n517) );
  INV_X1 U354 ( .A(n518), .ZN(n644) );
  AOI22_X1 U355 ( .A1(data_in[4]), .A2(n820), .B1(n514), .B2(\mem[20][4] ), 
        .ZN(n518) );
  INV_X1 U356 ( .A(n519), .ZN(n643) );
  AOI22_X1 U357 ( .A1(data_in[5]), .A2(n820), .B1(n514), .B2(\mem[20][5] ), 
        .ZN(n519) );
  INV_X1 U358 ( .A(n520), .ZN(n642) );
  AOI22_X1 U359 ( .A1(data_in[6]), .A2(n820), .B1(n514), .B2(\mem[20][6] ), 
        .ZN(n520) );
  INV_X1 U360 ( .A(n521), .ZN(n641) );
  AOI22_X1 U361 ( .A1(data_in[7]), .A2(n820), .B1(n514), .B2(\mem[20][7] ), 
        .ZN(n521) );
  INV_X1 U362 ( .A(n403), .ZN(n744) );
  AOI22_X1 U363 ( .A1(data_in[0]), .A2(n832), .B1(n404), .B2(\mem[8][0] ), 
        .ZN(n403) );
  INV_X1 U364 ( .A(n405), .ZN(n743) );
  AOI22_X1 U365 ( .A1(data_in[1]), .A2(n832), .B1(n404), .B2(\mem[8][1] ), 
        .ZN(n405) );
  INV_X1 U366 ( .A(n406), .ZN(n742) );
  AOI22_X1 U367 ( .A1(data_in[2]), .A2(n832), .B1(n404), .B2(\mem[8][2] ), 
        .ZN(n406) );
  INV_X1 U368 ( .A(n407), .ZN(n741) );
  AOI22_X1 U369 ( .A1(data_in[3]), .A2(n832), .B1(n404), .B2(\mem[8][3] ), 
        .ZN(n407) );
  INV_X1 U370 ( .A(n408), .ZN(n740) );
  AOI22_X1 U371 ( .A1(data_in[4]), .A2(n832), .B1(n404), .B2(\mem[8][4] ), 
        .ZN(n408) );
  INV_X1 U372 ( .A(n409), .ZN(n739) );
  AOI22_X1 U373 ( .A1(data_in[5]), .A2(n832), .B1(n404), .B2(\mem[8][5] ), 
        .ZN(n409) );
  INV_X1 U374 ( .A(n410), .ZN(n738) );
  AOI22_X1 U375 ( .A1(data_in[6]), .A2(n832), .B1(n404), .B2(\mem[8][6] ), 
        .ZN(n410) );
  INV_X1 U376 ( .A(n411), .ZN(n737) );
  AOI22_X1 U377 ( .A1(data_in[7]), .A2(n832), .B1(n404), .B2(\mem[8][7] ), 
        .ZN(n411) );
  INV_X1 U378 ( .A(n476), .ZN(n680) );
  AOI22_X1 U379 ( .A1(data_in[0]), .A2(n824), .B1(n477), .B2(\mem[16][0] ), 
        .ZN(n476) );
  INV_X1 U380 ( .A(n478), .ZN(n679) );
  AOI22_X1 U381 ( .A1(data_in[1]), .A2(n824), .B1(n477), .B2(\mem[16][1] ), 
        .ZN(n478) );
  INV_X1 U382 ( .A(n479), .ZN(n678) );
  AOI22_X1 U383 ( .A1(data_in[2]), .A2(n824), .B1(n477), .B2(\mem[16][2] ), 
        .ZN(n479) );
  INV_X1 U384 ( .A(n480), .ZN(n677) );
  AOI22_X1 U385 ( .A1(data_in[3]), .A2(n824), .B1(n477), .B2(\mem[16][3] ), 
        .ZN(n480) );
  INV_X1 U386 ( .A(n481), .ZN(n676) );
  AOI22_X1 U387 ( .A1(data_in[4]), .A2(n824), .B1(n477), .B2(\mem[16][4] ), 
        .ZN(n481) );
  INV_X1 U388 ( .A(n482), .ZN(n675) );
  AOI22_X1 U389 ( .A1(data_in[5]), .A2(n824), .B1(n477), .B2(\mem[16][5] ), 
        .ZN(n482) );
  INV_X1 U390 ( .A(n483), .ZN(n674) );
  AOI22_X1 U391 ( .A1(data_in[6]), .A2(n824), .B1(n477), .B2(\mem[16][6] ), 
        .ZN(n483) );
  INV_X1 U392 ( .A(n484), .ZN(n673) );
  AOI22_X1 U393 ( .A1(data_in[7]), .A2(n824), .B1(n477), .B2(\mem[16][7] ), 
        .ZN(n484) );
  INV_X1 U394 ( .A(n549), .ZN(n616) );
  AOI22_X1 U395 ( .A1(data_in[0]), .A2(n813), .B1(n550), .B2(\mem[24][0] ), 
        .ZN(n549) );
  INV_X1 U396 ( .A(n551), .ZN(n615) );
  AOI22_X1 U397 ( .A1(data_in[1]), .A2(n813), .B1(n550), .B2(\mem[24][1] ), 
        .ZN(n551) );
  INV_X1 U398 ( .A(n552), .ZN(n614) );
  AOI22_X1 U399 ( .A1(data_in[2]), .A2(n813), .B1(n550), .B2(\mem[24][2] ), 
        .ZN(n552) );
  INV_X1 U400 ( .A(n553), .ZN(n613) );
  AOI22_X1 U401 ( .A1(data_in[3]), .A2(n813), .B1(n550), .B2(\mem[24][3] ), 
        .ZN(n553) );
  INV_X1 U402 ( .A(n554), .ZN(n612) );
  AOI22_X1 U403 ( .A1(data_in[4]), .A2(n813), .B1(n550), .B2(\mem[24][4] ), 
        .ZN(n554) );
  INV_X1 U404 ( .A(n555), .ZN(n611) );
  AOI22_X1 U405 ( .A1(data_in[5]), .A2(n813), .B1(n550), .B2(\mem[24][5] ), 
        .ZN(n555) );
  INV_X1 U406 ( .A(n556), .ZN(n610) );
  AOI22_X1 U407 ( .A1(data_in[6]), .A2(n813), .B1(n550), .B2(\mem[24][6] ), 
        .ZN(n556) );
  INV_X1 U408 ( .A(n557), .ZN(n609) );
  AOI22_X1 U409 ( .A1(data_in[7]), .A2(n813), .B1(n550), .B2(\mem[24][7] ), 
        .ZN(n557) );
  INV_X1 U410 ( .A(n558), .ZN(n608) );
  AOI22_X1 U411 ( .A1(data_in[0]), .A2(n812), .B1(n559), .B2(\mem[25][0] ), 
        .ZN(n558) );
  INV_X1 U412 ( .A(n560), .ZN(n607) );
  AOI22_X1 U413 ( .A1(data_in[1]), .A2(n812), .B1(n559), .B2(\mem[25][1] ), 
        .ZN(n560) );
  INV_X1 U414 ( .A(n561), .ZN(n606) );
  AOI22_X1 U415 ( .A1(data_in[2]), .A2(n812), .B1(n559), .B2(\mem[25][2] ), 
        .ZN(n561) );
  INV_X1 U416 ( .A(n562), .ZN(n605) );
  AOI22_X1 U417 ( .A1(data_in[3]), .A2(n812), .B1(n559), .B2(\mem[25][3] ), 
        .ZN(n562) );
  INV_X1 U418 ( .A(n563), .ZN(n604) );
  AOI22_X1 U419 ( .A1(data_in[4]), .A2(n812), .B1(n559), .B2(\mem[25][4] ), 
        .ZN(n563) );
  INV_X1 U420 ( .A(n564), .ZN(n603) );
  AOI22_X1 U421 ( .A1(data_in[5]), .A2(n812), .B1(n559), .B2(\mem[25][5] ), 
        .ZN(n564) );
  INV_X1 U422 ( .A(n565), .ZN(n602) );
  AOI22_X1 U423 ( .A1(data_in[6]), .A2(n812), .B1(n559), .B2(\mem[25][6] ), 
        .ZN(n565) );
  INV_X1 U424 ( .A(n566), .ZN(n601) );
  AOI22_X1 U425 ( .A1(data_in[7]), .A2(n812), .B1(n559), .B2(\mem[25][7] ), 
        .ZN(n566) );
  INV_X1 U426 ( .A(n567), .ZN(n600) );
  AOI22_X1 U427 ( .A1(data_in[0]), .A2(n811), .B1(n568), .B2(\mem[26][0] ), 
        .ZN(n567) );
  INV_X1 U428 ( .A(n569), .ZN(n599) );
  AOI22_X1 U429 ( .A1(data_in[1]), .A2(n811), .B1(n568), .B2(\mem[26][1] ), 
        .ZN(n569) );
  INV_X1 U430 ( .A(n570), .ZN(n598) );
  AOI22_X1 U431 ( .A1(data_in[2]), .A2(n811), .B1(n568), .B2(\mem[26][2] ), 
        .ZN(n570) );
  INV_X1 U432 ( .A(n571), .ZN(n597) );
  AOI22_X1 U433 ( .A1(data_in[3]), .A2(n811), .B1(n568), .B2(\mem[26][3] ), 
        .ZN(n571) );
  INV_X1 U434 ( .A(n572), .ZN(n596) );
  AOI22_X1 U435 ( .A1(data_in[4]), .A2(n811), .B1(n568), .B2(\mem[26][4] ), 
        .ZN(n572) );
  INV_X1 U436 ( .A(n573), .ZN(n595) );
  AOI22_X1 U437 ( .A1(data_in[5]), .A2(n811), .B1(n568), .B2(\mem[26][5] ), 
        .ZN(n573) );
  INV_X1 U438 ( .A(n574), .ZN(n594) );
  AOI22_X1 U439 ( .A1(data_in[6]), .A2(n811), .B1(n568), .B2(\mem[26][6] ), 
        .ZN(n574) );
  INV_X1 U440 ( .A(n575), .ZN(n293) );
  AOI22_X1 U441 ( .A1(data_in[7]), .A2(n811), .B1(n568), .B2(\mem[26][7] ), 
        .ZN(n575) );
  INV_X1 U442 ( .A(n576), .ZN(n292) );
  AOI22_X1 U443 ( .A1(data_in[0]), .A2(n810), .B1(n577), .B2(\mem[27][0] ), 
        .ZN(n576) );
  INV_X1 U444 ( .A(n578), .ZN(n291) );
  AOI22_X1 U445 ( .A1(data_in[1]), .A2(n810), .B1(n577), .B2(\mem[27][1] ), 
        .ZN(n578) );
  INV_X1 U446 ( .A(n579), .ZN(n290) );
  AOI22_X1 U447 ( .A1(data_in[2]), .A2(n810), .B1(n577), .B2(\mem[27][2] ), 
        .ZN(n579) );
  INV_X1 U448 ( .A(n580), .ZN(n289) );
  AOI22_X1 U449 ( .A1(data_in[3]), .A2(n810), .B1(n577), .B2(\mem[27][3] ), 
        .ZN(n580) );
  INV_X1 U450 ( .A(n581), .ZN(n288) );
  AOI22_X1 U451 ( .A1(data_in[4]), .A2(n810), .B1(n577), .B2(\mem[27][4] ), 
        .ZN(n581) );
  INV_X1 U452 ( .A(n582), .ZN(n287) );
  AOI22_X1 U453 ( .A1(data_in[5]), .A2(n810), .B1(n577), .B2(\mem[27][5] ), 
        .ZN(n582) );
  INV_X1 U454 ( .A(n583), .ZN(n286) );
  AOI22_X1 U455 ( .A1(data_in[6]), .A2(n810), .B1(n577), .B2(\mem[27][6] ), 
        .ZN(n583) );
  INV_X1 U456 ( .A(n584), .ZN(n285) );
  AOI22_X1 U457 ( .A1(data_in[7]), .A2(n810), .B1(n577), .B2(\mem[27][7] ), 
        .ZN(n584) );
  INV_X1 U458 ( .A(n585), .ZN(n284) );
  AOI22_X1 U459 ( .A1(data_in[0]), .A2(n809), .B1(n586), .B2(\mem[28][0] ), 
        .ZN(n585) );
  INV_X1 U460 ( .A(n587), .ZN(n283) );
  AOI22_X1 U461 ( .A1(data_in[1]), .A2(n809), .B1(n586), .B2(\mem[28][1] ), 
        .ZN(n587) );
  INV_X1 U462 ( .A(n588), .ZN(n282) );
  AOI22_X1 U463 ( .A1(data_in[2]), .A2(n809), .B1(n586), .B2(\mem[28][2] ), 
        .ZN(n588) );
  INV_X1 U464 ( .A(n589), .ZN(n281) );
  AOI22_X1 U465 ( .A1(data_in[3]), .A2(n809), .B1(n586), .B2(\mem[28][3] ), 
        .ZN(n589) );
  INV_X1 U466 ( .A(n590), .ZN(n280) );
  AOI22_X1 U467 ( .A1(data_in[4]), .A2(n809), .B1(n586), .B2(\mem[28][4] ), 
        .ZN(n590) );
  INV_X1 U468 ( .A(n591), .ZN(n279) );
  AOI22_X1 U469 ( .A1(data_in[5]), .A2(n809), .B1(n586), .B2(\mem[28][5] ), 
        .ZN(n591) );
  INV_X1 U470 ( .A(n592), .ZN(n278) );
  AOI22_X1 U471 ( .A1(data_in[6]), .A2(n809), .B1(n586), .B2(\mem[28][6] ), 
        .ZN(n592) );
  INV_X1 U472 ( .A(n593), .ZN(n277) );
  AOI22_X1 U473 ( .A1(data_in[7]), .A2(n809), .B1(n586), .B2(\mem[28][7] ), 
        .ZN(n593) );
  INV_X1 U474 ( .A(n294), .ZN(n276) );
  AOI22_X1 U475 ( .A1(n816), .A2(data_in[0]), .B1(n295), .B2(\mem[29][0] ), 
        .ZN(n294) );
  INV_X1 U476 ( .A(n296), .ZN(n275) );
  AOI22_X1 U477 ( .A1(n816), .A2(data_in[1]), .B1(n295), .B2(\mem[29][1] ), 
        .ZN(n296) );
  INV_X1 U478 ( .A(n297), .ZN(n274) );
  AOI22_X1 U479 ( .A1(n816), .A2(data_in[2]), .B1(n295), .B2(\mem[29][2] ), 
        .ZN(n297) );
  INV_X1 U480 ( .A(n298), .ZN(n273) );
  AOI22_X1 U481 ( .A1(n816), .A2(data_in[3]), .B1(n295), .B2(\mem[29][3] ), 
        .ZN(n298) );
  INV_X1 U482 ( .A(n299), .ZN(n272) );
  AOI22_X1 U483 ( .A1(n816), .A2(data_in[4]), .B1(n295), .B2(\mem[29][4] ), 
        .ZN(n299) );
  INV_X1 U484 ( .A(n300), .ZN(n271) );
  AOI22_X1 U485 ( .A1(n816), .A2(data_in[5]), .B1(n295), .B2(\mem[29][5] ), 
        .ZN(n300) );
  INV_X1 U486 ( .A(n301), .ZN(n270) );
  AOI22_X1 U487 ( .A1(n816), .A2(data_in[6]), .B1(n295), .B2(\mem[29][6] ), 
        .ZN(n301) );
  INV_X1 U488 ( .A(n302), .ZN(n269) );
  AOI22_X1 U489 ( .A1(n816), .A2(data_in[7]), .B1(n295), .B2(\mem[29][7] ), 
        .ZN(n302) );
  INV_X1 U490 ( .A(n305), .ZN(n268) );
  AOI22_X1 U491 ( .A1(data_in[0]), .A2(n815), .B1(n306), .B2(\mem[30][0] ), 
        .ZN(n305) );
  INV_X1 U492 ( .A(n307), .ZN(n267) );
  AOI22_X1 U493 ( .A1(data_in[1]), .A2(n815), .B1(n306), .B2(\mem[30][1] ), 
        .ZN(n307) );
  INV_X1 U494 ( .A(n308), .ZN(n266) );
  AOI22_X1 U495 ( .A1(data_in[2]), .A2(n815), .B1(n306), .B2(\mem[30][2] ), 
        .ZN(n308) );
  INV_X1 U496 ( .A(n309), .ZN(n265) );
  AOI22_X1 U497 ( .A1(data_in[3]), .A2(n815), .B1(n306), .B2(\mem[30][3] ), 
        .ZN(n309) );
  INV_X1 U498 ( .A(n310), .ZN(n264) );
  AOI22_X1 U499 ( .A1(data_in[4]), .A2(n815), .B1(n306), .B2(\mem[30][4] ), 
        .ZN(n310) );
  INV_X1 U500 ( .A(n311), .ZN(n263) );
  AOI22_X1 U501 ( .A1(data_in[5]), .A2(n815), .B1(n306), .B2(\mem[30][5] ), 
        .ZN(n311) );
  INV_X1 U502 ( .A(n312), .ZN(n262) );
  AOI22_X1 U503 ( .A1(data_in[6]), .A2(n815), .B1(n306), .B2(\mem[30][6] ), 
        .ZN(n312) );
  INV_X1 U504 ( .A(n313), .ZN(n261) );
  AOI22_X1 U505 ( .A1(data_in[7]), .A2(n815), .B1(n306), .B2(\mem[30][7] ), 
        .ZN(n313) );
  INV_X1 U506 ( .A(n315), .ZN(n260) );
  AOI22_X1 U507 ( .A1(data_in[0]), .A2(n814), .B1(n316), .B2(\mem[31][0] ), 
        .ZN(n315) );
  INV_X1 U508 ( .A(n317), .ZN(n259) );
  AOI22_X1 U509 ( .A1(data_in[1]), .A2(n814), .B1(n316), .B2(\mem[31][1] ), 
        .ZN(n317) );
  INV_X1 U510 ( .A(n318), .ZN(n258) );
  AOI22_X1 U511 ( .A1(data_in[2]), .A2(n814), .B1(n316), .B2(\mem[31][2] ), 
        .ZN(n318) );
  INV_X1 U512 ( .A(n319), .ZN(n257) );
  AOI22_X1 U513 ( .A1(data_in[3]), .A2(n814), .B1(n316), .B2(\mem[31][3] ), 
        .ZN(n319) );
  INV_X1 U514 ( .A(n320), .ZN(n256) );
  AOI22_X1 U515 ( .A1(data_in[4]), .A2(n814), .B1(n316), .B2(\mem[31][4] ), 
        .ZN(n320) );
  INV_X1 U516 ( .A(n321), .ZN(n255) );
  AOI22_X1 U517 ( .A1(data_in[5]), .A2(n814), .B1(n316), .B2(\mem[31][5] ), 
        .ZN(n321) );
  INV_X1 U518 ( .A(n322), .ZN(n254) );
  AOI22_X1 U519 ( .A1(data_in[6]), .A2(n814), .B1(n316), .B2(\mem[31][6] ), 
        .ZN(n322) );
  INV_X1 U520 ( .A(n323), .ZN(n253) );
  AOI22_X1 U521 ( .A1(data_in[7]), .A2(n814), .B1(n316), .B2(\mem[31][7] ), 
        .ZN(n323) );
  INV_X1 U522 ( .A(n325), .ZN(n808) );
  AOI22_X1 U523 ( .A1(data_in[0]), .A2(n840), .B1(n326), .B2(\mem[0][0] ), 
        .ZN(n325) );
  INV_X1 U524 ( .A(n327), .ZN(n807) );
  AOI22_X1 U525 ( .A1(data_in[1]), .A2(n840), .B1(n326), .B2(\mem[0][1] ), 
        .ZN(n327) );
  INV_X1 U526 ( .A(n328), .ZN(n806) );
  AOI22_X1 U527 ( .A1(data_in[2]), .A2(n840), .B1(n326), .B2(\mem[0][2] ), 
        .ZN(n328) );
  INV_X1 U528 ( .A(n329), .ZN(n805) );
  AOI22_X1 U529 ( .A1(data_in[3]), .A2(n840), .B1(n326), .B2(\mem[0][3] ), 
        .ZN(n329) );
  INV_X1 U530 ( .A(n330), .ZN(n804) );
  AOI22_X1 U531 ( .A1(data_in[4]), .A2(n840), .B1(n326), .B2(\mem[0][4] ), 
        .ZN(n330) );
  INV_X1 U532 ( .A(n331), .ZN(n803) );
  AOI22_X1 U533 ( .A1(data_in[5]), .A2(n840), .B1(n326), .B2(\mem[0][5] ), 
        .ZN(n331) );
  INV_X1 U534 ( .A(n332), .ZN(n802) );
  AOI22_X1 U535 ( .A1(data_in[6]), .A2(n840), .B1(n326), .B2(\mem[0][6] ), 
        .ZN(n332) );
  INV_X1 U536 ( .A(n333), .ZN(n801) );
  AOI22_X1 U537 ( .A1(data_in[7]), .A2(n840), .B1(n326), .B2(\mem[0][7] ), 
        .ZN(n333) );
  INV_X1 U538 ( .A(n336), .ZN(n800) );
  AOI22_X1 U539 ( .A1(data_in[0]), .A2(n839), .B1(n337), .B2(\mem[1][0] ), 
        .ZN(n336) );
  INV_X1 U540 ( .A(n338), .ZN(n799) );
  AOI22_X1 U541 ( .A1(data_in[1]), .A2(n839), .B1(n337), .B2(\mem[1][1] ), 
        .ZN(n338) );
  INV_X1 U542 ( .A(n339), .ZN(n798) );
  AOI22_X1 U543 ( .A1(data_in[2]), .A2(n839), .B1(n337), .B2(\mem[1][2] ), 
        .ZN(n339) );
  INV_X1 U544 ( .A(n340), .ZN(n797) );
  AOI22_X1 U545 ( .A1(data_in[3]), .A2(n839), .B1(n337), .B2(\mem[1][3] ), 
        .ZN(n340) );
  INV_X1 U546 ( .A(n341), .ZN(n796) );
  AOI22_X1 U547 ( .A1(data_in[4]), .A2(n839), .B1(n337), .B2(\mem[1][4] ), 
        .ZN(n341) );
  INV_X1 U548 ( .A(n342), .ZN(n795) );
  AOI22_X1 U549 ( .A1(data_in[5]), .A2(n839), .B1(n337), .B2(\mem[1][5] ), 
        .ZN(n342) );
  INV_X1 U550 ( .A(n343), .ZN(n794) );
  AOI22_X1 U551 ( .A1(data_in[6]), .A2(n839), .B1(n337), .B2(\mem[1][6] ), 
        .ZN(n343) );
  INV_X1 U552 ( .A(n344), .ZN(n793) );
  AOI22_X1 U553 ( .A1(data_in[7]), .A2(n839), .B1(n337), .B2(\mem[1][7] ), 
        .ZN(n344) );
  INV_X1 U554 ( .A(n346), .ZN(n792) );
  AOI22_X1 U555 ( .A1(data_in[0]), .A2(n838), .B1(n347), .B2(\mem[2][0] ), 
        .ZN(n346) );
  INV_X1 U556 ( .A(n348), .ZN(n791) );
  AOI22_X1 U557 ( .A1(data_in[1]), .A2(n838), .B1(n347), .B2(\mem[2][1] ), 
        .ZN(n348) );
  INV_X1 U558 ( .A(n349), .ZN(n790) );
  AOI22_X1 U559 ( .A1(data_in[2]), .A2(n838), .B1(n347), .B2(\mem[2][2] ), 
        .ZN(n349) );
  INV_X1 U560 ( .A(n350), .ZN(n789) );
  AOI22_X1 U561 ( .A1(data_in[3]), .A2(n838), .B1(n347), .B2(\mem[2][3] ), 
        .ZN(n350) );
  INV_X1 U562 ( .A(n351), .ZN(n788) );
  AOI22_X1 U563 ( .A1(data_in[4]), .A2(n838), .B1(n347), .B2(\mem[2][4] ), 
        .ZN(n351) );
  INV_X1 U564 ( .A(n352), .ZN(n787) );
  AOI22_X1 U565 ( .A1(data_in[5]), .A2(n838), .B1(n347), .B2(\mem[2][5] ), 
        .ZN(n352) );
  INV_X1 U566 ( .A(n353), .ZN(n786) );
  AOI22_X1 U567 ( .A1(data_in[6]), .A2(n838), .B1(n347), .B2(\mem[2][6] ), 
        .ZN(n353) );
  INV_X1 U568 ( .A(n354), .ZN(n785) );
  AOI22_X1 U569 ( .A1(data_in[7]), .A2(n838), .B1(n347), .B2(\mem[2][7] ), 
        .ZN(n354) );
  INV_X1 U570 ( .A(n356), .ZN(n784) );
  AOI22_X1 U571 ( .A1(data_in[0]), .A2(n837), .B1(n357), .B2(\mem[3][0] ), 
        .ZN(n356) );
  INV_X1 U572 ( .A(n358), .ZN(n783) );
  AOI22_X1 U573 ( .A1(data_in[1]), .A2(n837), .B1(n357), .B2(\mem[3][1] ), 
        .ZN(n358) );
  INV_X1 U574 ( .A(n359), .ZN(n782) );
  AOI22_X1 U575 ( .A1(data_in[2]), .A2(n837), .B1(n357), .B2(\mem[3][2] ), 
        .ZN(n359) );
  INV_X1 U576 ( .A(n360), .ZN(n781) );
  AOI22_X1 U577 ( .A1(data_in[3]), .A2(n837), .B1(n357), .B2(\mem[3][3] ), 
        .ZN(n360) );
  INV_X1 U578 ( .A(n361), .ZN(n780) );
  AOI22_X1 U579 ( .A1(data_in[4]), .A2(n837), .B1(n357), .B2(\mem[3][4] ), 
        .ZN(n361) );
  INV_X1 U580 ( .A(n362), .ZN(n779) );
  AOI22_X1 U581 ( .A1(data_in[5]), .A2(n837), .B1(n357), .B2(\mem[3][5] ), 
        .ZN(n362) );
  INV_X1 U582 ( .A(n363), .ZN(n778) );
  AOI22_X1 U583 ( .A1(data_in[6]), .A2(n837), .B1(n357), .B2(\mem[3][6] ), 
        .ZN(n363) );
  INV_X1 U584 ( .A(n364), .ZN(n777) );
  AOI22_X1 U585 ( .A1(data_in[7]), .A2(n837), .B1(n357), .B2(\mem[3][7] ), 
        .ZN(n364) );
  INV_X1 U586 ( .A(n366), .ZN(n776) );
  AOI22_X1 U587 ( .A1(data_in[0]), .A2(n836), .B1(n367), .B2(\mem[4][0] ), 
        .ZN(n366) );
  INV_X1 U588 ( .A(n368), .ZN(n775) );
  AOI22_X1 U589 ( .A1(data_in[1]), .A2(n836), .B1(n367), .B2(\mem[4][1] ), 
        .ZN(n368) );
  INV_X1 U590 ( .A(n369), .ZN(n774) );
  AOI22_X1 U591 ( .A1(data_in[2]), .A2(n836), .B1(n367), .B2(\mem[4][2] ), 
        .ZN(n369) );
  INV_X1 U592 ( .A(n370), .ZN(n773) );
  AOI22_X1 U593 ( .A1(data_in[3]), .A2(n836), .B1(n367), .B2(\mem[4][3] ), 
        .ZN(n370) );
  INV_X1 U594 ( .A(n371), .ZN(n772) );
  AOI22_X1 U595 ( .A1(data_in[4]), .A2(n836), .B1(n367), .B2(\mem[4][4] ), 
        .ZN(n371) );
  INV_X1 U596 ( .A(n372), .ZN(n771) );
  AOI22_X1 U597 ( .A1(data_in[5]), .A2(n836), .B1(n367), .B2(\mem[4][5] ), 
        .ZN(n372) );
  INV_X1 U598 ( .A(n373), .ZN(n770) );
  AOI22_X1 U599 ( .A1(data_in[6]), .A2(n836), .B1(n367), .B2(\mem[4][6] ), 
        .ZN(n373) );
  INV_X1 U600 ( .A(n374), .ZN(n769) );
  AOI22_X1 U601 ( .A1(data_in[7]), .A2(n836), .B1(n367), .B2(\mem[4][7] ), 
        .ZN(n374) );
  INV_X1 U602 ( .A(N13), .ZN(n841) );
  INV_X1 U603 ( .A(N14), .ZN(n842) );
  INV_X1 U604 ( .A(N12), .ZN(n252) );
  MUX2_X1 U605 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n248), .Z(n1) );
  MUX2_X1 U606 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n248), .Z(n2) );
  MUX2_X1 U607 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U608 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n248), .Z(n4) );
  MUX2_X1 U609 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n247), .Z(n5) );
  MUX2_X1 U610 ( .A(n5), .B(n4), .S(n242), .Z(n6) );
  MUX2_X1 U611 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U612 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n248), .Z(n8) );
  MUX2_X1 U613 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n248), .Z(n9) );
  MUX2_X1 U614 ( .A(n9), .B(n8), .S(N11), .Z(n10) );
  MUX2_X1 U615 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n248), .Z(n11) );
  MUX2_X1 U616 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n247), .Z(n12) );
  MUX2_X1 U617 ( .A(n12), .B(n11), .S(n244), .Z(n13) );
  MUX2_X1 U618 ( .A(n13), .B(n10), .S(n241), .Z(n14) );
  MUX2_X1 U619 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U620 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n245), .Z(n16) );
  MUX2_X1 U621 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n245), .Z(n17) );
  MUX2_X1 U622 ( .A(n17), .B(n16), .S(n243), .Z(n18) );
  MUX2_X1 U623 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U624 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n245), .Z(n20) );
  MUX2_X1 U625 ( .A(n20), .B(n19), .S(N11), .Z(n21) );
  MUX2_X1 U626 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U627 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n245), .Z(n23) );
  MUX2_X1 U628 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n245), .Z(n24) );
  MUX2_X1 U629 ( .A(n24), .B(n23), .S(n243), .Z(n25) );
  MUX2_X1 U630 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n245), .Z(n26) );
  MUX2_X1 U631 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n245), .Z(n27) );
  MUX2_X1 U632 ( .A(n27), .B(n26), .S(N11), .Z(n28) );
  MUX2_X1 U633 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U634 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U635 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U636 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n245), .Z(n31) );
  MUX2_X1 U637 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n245), .Z(n32) );
  MUX2_X1 U638 ( .A(n32), .B(n31), .S(n242), .Z(n33) );
  MUX2_X1 U639 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U640 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U641 ( .A(n35), .B(n34), .S(n242), .Z(n36) );
  MUX2_X1 U642 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U643 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n246), .Z(n38) );
  MUX2_X1 U644 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n246), .Z(n39) );
  MUX2_X1 U645 ( .A(n39), .B(n38), .S(n244), .Z(n40) );
  MUX2_X1 U646 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n246), .Z(n41) );
  MUX2_X1 U647 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n246), .Z(n42) );
  MUX2_X1 U648 ( .A(n42), .B(n41), .S(N11), .Z(n43) );
  MUX2_X1 U649 ( .A(n43), .B(n40), .S(N12), .Z(n44) );
  MUX2_X1 U650 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U651 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n246), .Z(n46) );
  MUX2_X1 U652 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n246), .Z(n47) );
  MUX2_X1 U653 ( .A(n47), .B(n46), .S(n244), .Z(n48) );
  MUX2_X1 U654 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n246), .Z(n49) );
  MUX2_X1 U655 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n246), .Z(n50) );
  MUX2_X1 U656 ( .A(n50), .B(n49), .S(N11), .Z(n51) );
  MUX2_X1 U657 ( .A(n51), .B(n48), .S(N12), .Z(n52) );
  MUX2_X1 U658 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n246), .Z(n53) );
  MUX2_X1 U659 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n246), .Z(n54) );
  MUX2_X1 U660 ( .A(n54), .B(n53), .S(n244), .Z(n55) );
  MUX2_X1 U661 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n246), .Z(n56) );
  MUX2_X1 U662 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n246), .Z(n57) );
  MUX2_X1 U663 ( .A(n57), .B(n56), .S(N11), .Z(n58) );
  MUX2_X1 U664 ( .A(n58), .B(n55), .S(N12), .Z(n59) );
  MUX2_X1 U665 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U666 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U667 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n246), .Z(n61) );
  MUX2_X1 U668 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n245), .Z(n62) );
  MUX2_X1 U669 ( .A(n62), .B(n61), .S(N11), .Z(n63) );
  MUX2_X1 U670 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n247), .Z(n64) );
  MUX2_X1 U671 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n246), .Z(n65) );
  MUX2_X1 U672 ( .A(n65), .B(n64), .S(N11), .Z(n66) );
  MUX2_X1 U673 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U674 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n245), .Z(n68) );
  MUX2_X1 U675 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n247), .Z(n69) );
  MUX2_X1 U676 ( .A(n69), .B(n68), .S(N11), .Z(n70) );
  MUX2_X1 U677 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n247), .Z(n71) );
  MUX2_X1 U678 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n246), .Z(n72) );
  MUX2_X1 U679 ( .A(n72), .B(n71), .S(n243), .Z(n73) );
  MUX2_X1 U680 ( .A(n73), .B(n70), .S(n241), .Z(n74) );
  MUX2_X1 U681 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U682 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n246), .Z(n76) );
  MUX2_X1 U683 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n245), .Z(n77) );
  MUX2_X1 U684 ( .A(n77), .B(n76), .S(N11), .Z(n78) );
  MUX2_X1 U685 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n245), .Z(n79) );
  MUX2_X1 U686 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n247), .Z(n80) );
  MUX2_X1 U687 ( .A(n80), .B(n79), .S(n242), .Z(n81) );
  MUX2_X1 U688 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U689 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n246), .Z(n83) );
  MUX2_X1 U690 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n247), .Z(n84) );
  MUX2_X1 U691 ( .A(n84), .B(n83), .S(n243), .Z(n85) );
  MUX2_X1 U692 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n245), .Z(n86) );
  MUX2_X1 U693 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n247), .Z(n87) );
  MUX2_X1 U694 ( .A(n87), .B(n86), .S(n243), .Z(n88) );
  MUX2_X1 U695 ( .A(n88), .B(n85), .S(n241), .Z(n89) );
  MUX2_X1 U696 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U697 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U698 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n249), .Z(n91) );
  MUX2_X1 U699 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n249), .Z(n92) );
  MUX2_X1 U700 ( .A(n92), .B(n91), .S(N11), .Z(n93) );
  MUX2_X1 U701 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n246), .Z(n94) );
  MUX2_X1 U702 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n247), .Z(n95) );
  MUX2_X1 U703 ( .A(n95), .B(n94), .S(N11), .Z(n96) );
  MUX2_X1 U704 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U705 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n247), .Z(n98) );
  MUX2_X1 U706 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n245), .Z(n99) );
  MUX2_X1 U707 ( .A(n99), .B(n98), .S(N11), .Z(n100) );
  MUX2_X1 U708 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n246), .Z(n101) );
  MUX2_X1 U709 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n246), .Z(n102) );
  MUX2_X1 U710 ( .A(n102), .B(n101), .S(n244), .Z(n103) );
  MUX2_X1 U711 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U712 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U713 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n248), .Z(n106) );
  MUX2_X1 U714 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n249), .Z(n107) );
  MUX2_X1 U715 ( .A(n107), .B(n106), .S(n242), .Z(n108) );
  MUX2_X1 U716 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n248), .Z(n109) );
  MUX2_X1 U717 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n110) );
  MUX2_X1 U718 ( .A(n110), .B(n109), .S(n242), .Z(n111) );
  MUX2_X1 U719 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U720 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(N10), .Z(n113) );
  MUX2_X1 U721 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n114) );
  MUX2_X1 U722 ( .A(n114), .B(n113), .S(n242), .Z(n115) );
  MUX2_X1 U723 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n116) );
  MUX2_X1 U724 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n117) );
  MUX2_X1 U725 ( .A(n117), .B(n116), .S(n242), .Z(n118) );
  MUX2_X1 U726 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U727 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U728 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U729 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n248), .Z(n121) );
  MUX2_X1 U730 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(N10), .Z(n122) );
  MUX2_X1 U731 ( .A(n122), .B(n121), .S(n242), .Z(n123) );
  MUX2_X1 U732 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n248), .Z(n124) );
  MUX2_X1 U733 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n249), .Z(n125) );
  MUX2_X1 U734 ( .A(n125), .B(n124), .S(n242), .Z(n126) );
  MUX2_X1 U735 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U736 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n247), .Z(n128) );
  MUX2_X1 U737 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n247), .Z(n129) );
  MUX2_X1 U738 ( .A(n129), .B(n128), .S(n242), .Z(n130) );
  MUX2_X1 U739 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n247), .Z(n131) );
  MUX2_X1 U740 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n247), .Z(n132) );
  MUX2_X1 U741 ( .A(n132), .B(n131), .S(n242), .Z(n133) );
  MUX2_X1 U742 ( .A(n133), .B(n130), .S(n241), .Z(n134) );
  MUX2_X1 U743 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U744 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n247), .Z(n136) );
  MUX2_X1 U745 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n247), .Z(n137) );
  MUX2_X1 U746 ( .A(n137), .B(n136), .S(n242), .Z(n138) );
  MUX2_X1 U747 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n247), .Z(n139) );
  MUX2_X1 U748 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n247), .Z(n140) );
  MUX2_X1 U749 ( .A(n140), .B(n139), .S(n242), .Z(n141) );
  MUX2_X1 U750 ( .A(n141), .B(n138), .S(n241), .Z(n142) );
  MUX2_X1 U751 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n247), .Z(n143) );
  MUX2_X1 U752 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n247), .Z(n144) );
  MUX2_X1 U753 ( .A(n144), .B(n143), .S(n242), .Z(n145) );
  MUX2_X1 U754 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n247), .Z(n146) );
  MUX2_X1 U755 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n247), .Z(n147) );
  MUX2_X1 U756 ( .A(n147), .B(n146), .S(n242), .Z(n148) );
  MUX2_X1 U757 ( .A(n148), .B(n145), .S(n241), .Z(n149) );
  MUX2_X1 U758 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U759 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U760 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n248), .Z(n151) );
  MUX2_X1 U761 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n248), .Z(n152) );
  MUX2_X1 U762 ( .A(n152), .B(n151), .S(n243), .Z(n153) );
  MUX2_X1 U763 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n248), .Z(n154) );
  MUX2_X1 U764 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n248), .Z(n155) );
  MUX2_X1 U765 ( .A(n155), .B(n154), .S(n243), .Z(n156) );
  MUX2_X1 U766 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U767 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n248), .Z(n158) );
  MUX2_X1 U768 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n248), .Z(n159) );
  MUX2_X1 U769 ( .A(n159), .B(n158), .S(n243), .Z(n160) );
  MUX2_X1 U770 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n248), .Z(n161) );
  MUX2_X1 U771 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n248), .Z(n162) );
  MUX2_X1 U772 ( .A(n162), .B(n161), .S(n243), .Z(n163) );
  MUX2_X1 U773 ( .A(n163), .B(n160), .S(N12), .Z(n164) );
  MUX2_X1 U774 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U775 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n248), .Z(n166) );
  MUX2_X1 U776 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n248), .Z(n167) );
  MUX2_X1 U777 ( .A(n167), .B(n166), .S(n243), .Z(n168) );
  MUX2_X1 U778 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n248), .Z(n169) );
  MUX2_X1 U779 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n248), .Z(n170) );
  MUX2_X1 U780 ( .A(n170), .B(n169), .S(n243), .Z(n171) );
  MUX2_X1 U781 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U782 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n246), .Z(n173) );
  MUX2_X1 U783 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n249), .Z(n174) );
  MUX2_X1 U784 ( .A(n174), .B(n173), .S(n243), .Z(n175) );
  MUX2_X1 U785 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n249), .Z(n176) );
  MUX2_X1 U786 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n249), .Z(n177) );
  MUX2_X1 U787 ( .A(n177), .B(n176), .S(n243), .Z(n178) );
  MUX2_X1 U788 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U789 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U790 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U791 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n248), .Z(n181) );
  MUX2_X1 U792 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n249), .Z(n182) );
  MUX2_X1 U793 ( .A(n182), .B(n181), .S(n243), .Z(n183) );
  MUX2_X1 U794 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n249), .Z(n184) );
  MUX2_X1 U795 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n245), .Z(n185) );
  MUX2_X1 U796 ( .A(n185), .B(n184), .S(n243), .Z(n186) );
  MUX2_X1 U797 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U798 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n246), .Z(n188) );
  MUX2_X1 U799 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n249), .Z(n189) );
  MUX2_X1 U800 ( .A(n189), .B(n188), .S(n243), .Z(n190) );
  MUX2_X1 U801 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n245), .Z(n191) );
  MUX2_X1 U802 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n245), .Z(n192) );
  MUX2_X1 U803 ( .A(n192), .B(n191), .S(n243), .Z(n193) );
  MUX2_X1 U804 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U805 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U806 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n249), .Z(n196) );
  MUX2_X1 U807 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(N10), .Z(n197) );
  MUX2_X1 U808 ( .A(n197), .B(n196), .S(n244), .Z(n198) );
  MUX2_X1 U809 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(N10), .Z(n199) );
  MUX2_X1 U810 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n249), .Z(n200) );
  MUX2_X1 U811 ( .A(n200), .B(n199), .S(n244), .Z(n201) );
  MUX2_X1 U812 ( .A(n201), .B(n198), .S(n241), .Z(n202) );
  MUX2_X1 U813 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n249), .Z(n203) );
  MUX2_X1 U814 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n249), .Z(n204) );
  MUX2_X1 U815 ( .A(n204), .B(n203), .S(n244), .Z(n205) );
  MUX2_X1 U816 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n249), .Z(n206) );
  MUX2_X1 U817 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n249), .Z(n207) );
  MUX2_X1 U818 ( .A(n207), .B(n206), .S(n244), .Z(n208) );
  MUX2_X1 U819 ( .A(n208), .B(n205), .S(N12), .Z(n209) );
  MUX2_X1 U820 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U821 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U822 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n249), .Z(n211) );
  MUX2_X1 U823 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(N10), .Z(n212) );
  MUX2_X1 U824 ( .A(n212), .B(n211), .S(n244), .Z(n213) );
  MUX2_X1 U825 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(N10), .Z(n214) );
  MUX2_X1 U826 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n249), .Z(n215) );
  MUX2_X1 U827 ( .A(n215), .B(n214), .S(n244), .Z(n216) );
  MUX2_X1 U828 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U829 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n247), .Z(n218) );
  MUX2_X1 U830 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(N10), .Z(n219) );
  MUX2_X1 U831 ( .A(n219), .B(n218), .S(n244), .Z(n220) );
  MUX2_X1 U832 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n249), .Z(n221) );
  MUX2_X1 U833 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n222) );
  MUX2_X1 U834 ( .A(n222), .B(n221), .S(n244), .Z(n223) );
  MUX2_X1 U835 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U836 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U837 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n249), .Z(n226) );
  MUX2_X1 U838 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n246), .Z(n227) );
  MUX2_X1 U839 ( .A(n227), .B(n226), .S(n244), .Z(n228) );
  MUX2_X1 U840 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n245), .Z(n229) );
  MUX2_X1 U841 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n245), .Z(n230) );
  MUX2_X1 U842 ( .A(n230), .B(n229), .S(n244), .Z(n231) );
  MUX2_X1 U843 ( .A(n231), .B(n228), .S(n241), .Z(n232) );
  MUX2_X1 U844 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n249), .Z(n233) );
  MUX2_X1 U845 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n234) );
  MUX2_X1 U846 ( .A(n234), .B(n233), .S(n244), .Z(n235) );
  MUX2_X1 U847 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n236) );
  MUX2_X1 U848 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n237) );
  MUX2_X1 U849 ( .A(n237), .B(n236), .S(n244), .Z(n238) );
  MUX2_X1 U850 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U851 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U852 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_32 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(n250), .Z(n249) );
  BUF_X1 U4 ( .A(n250), .Z(n246) );
  BUF_X1 U5 ( .A(n250), .Z(n247) );
  BUF_X1 U6 ( .A(N10), .Z(n248) );
  BUF_X1 U7 ( .A(n250), .Z(n245) );
  BUF_X1 U8 ( .A(N10), .Z(n250) );
  INV_X1 U9 ( .A(n1111), .ZN(n841) );
  INV_X1 U10 ( .A(n1100), .ZN(n840) );
  INV_X1 U11 ( .A(n1090), .ZN(n839) );
  INV_X1 U12 ( .A(n1080), .ZN(n838) );
  INV_X1 U13 ( .A(n1070), .ZN(n837) );
  INV_X1 U14 ( .A(n1060), .ZN(n836) );
  INV_X1 U15 ( .A(n1051), .ZN(n835) );
  INV_X1 U16 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U19 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U20 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U21 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U22 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U23 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U24 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U26 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U27 ( .A(n1131), .ZN(n816) );
  INV_X1 U28 ( .A(n1121), .ZN(n815) );
  INV_X1 U29 ( .A(n887), .ZN(n814) );
  INV_X1 U30 ( .A(n878), .ZN(n813) );
  INV_X1 U31 ( .A(n869), .ZN(n812) );
  INV_X1 U32 ( .A(n860), .ZN(n811) );
  INV_X1 U33 ( .A(n851), .ZN(n810) );
  INV_X1 U34 ( .A(n987), .ZN(n828) );
  INV_X1 U35 ( .A(n978), .ZN(n827) );
  INV_X1 U36 ( .A(n969), .ZN(n826) );
  INV_X1 U37 ( .A(n914), .ZN(n820) );
  INV_X1 U38 ( .A(n905), .ZN(n819) );
  INV_X1 U39 ( .A(n896), .ZN(n818) );
  INV_X1 U40 ( .A(n1033), .ZN(n833) );
  INV_X1 U41 ( .A(n1023), .ZN(n832) );
  INV_X1 U42 ( .A(n1014), .ZN(n831) );
  INV_X1 U43 ( .A(n1005), .ZN(n830) );
  INV_X1 U44 ( .A(n996), .ZN(n829) );
  INV_X1 U45 ( .A(n960), .ZN(n825) );
  INV_X1 U46 ( .A(n950), .ZN(n824) );
  INV_X1 U47 ( .A(n941), .ZN(n823) );
  INV_X1 U48 ( .A(n932), .ZN(n822) );
  INV_X1 U49 ( .A(n923), .ZN(n821) );
  INV_X1 U50 ( .A(n1142), .ZN(n817) );
  BUF_X1 U51 ( .A(N11), .Z(n242) );
  BUF_X1 U52 ( .A(N11), .Z(n243) );
  BUF_X1 U53 ( .A(N11), .Z(n244) );
  INV_X1 U54 ( .A(N10), .ZN(n251) );
  BUF_X1 U55 ( .A(N12), .Z(n241) );
  NOR3_X1 U56 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U57 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U58 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U60 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U62 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U63 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U64 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U65 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U67 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U69 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U70 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U71 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U72 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U73 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U74 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U75 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U76 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U77 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U79 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U81 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U82 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U83 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U84 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U85 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U86 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U88 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U89 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U90 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U92 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U94 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U95 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U96 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U97 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U98 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U99 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U100 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U101 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U102 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U103 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U104 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U105 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U106 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U107 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U108 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U109 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U110 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U111 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U112 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U113 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U114 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U115 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U116 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U117 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U118 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U119 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U120 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U121 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U122 ( .A(n988), .ZN(n705) );
  AOI22_X1 U123 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U124 ( .A(n986), .ZN(n704) );
  AOI22_X1 U125 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U126 ( .A(n985), .ZN(n703) );
  AOI22_X1 U127 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U128 ( .A(n984), .ZN(n702) );
  AOI22_X1 U129 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U130 ( .A(n983), .ZN(n701) );
  AOI22_X1 U131 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U132 ( .A(n982), .ZN(n700) );
  AOI22_X1 U133 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U134 ( .A(n981), .ZN(n699) );
  AOI22_X1 U135 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U136 ( .A(n980), .ZN(n698) );
  AOI22_X1 U137 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U138 ( .A(n913), .ZN(n640) );
  AOI22_X1 U139 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U140 ( .A(n912), .ZN(n639) );
  AOI22_X1 U141 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U142 ( .A(n911), .ZN(n638) );
  AOI22_X1 U143 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U144 ( .A(n910), .ZN(n637) );
  AOI22_X1 U145 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U146 ( .A(n909), .ZN(n636) );
  AOI22_X1 U147 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U148 ( .A(n908), .ZN(n635) );
  AOI22_X1 U149 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U150 ( .A(n907), .ZN(n634) );
  AOI22_X1 U151 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U152 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U153 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U154 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U155 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U156 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U157 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U158 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U159 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U160 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U161 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U162 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U163 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U164 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U165 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U166 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U167 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U168 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U169 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U170 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U171 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U172 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U173 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U174 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U175 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U176 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U177 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U178 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U179 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U180 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U181 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U182 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U183 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U184 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U185 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U186 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U187 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U188 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U189 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U190 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U191 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U192 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U193 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U194 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U195 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U196 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U197 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U198 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U199 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U200 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U201 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U202 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U203 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U204 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U205 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U206 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U207 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U208 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U209 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U210 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U211 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U212 ( .A(n999), .ZN(n715) );
  AOI22_X1 U213 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U214 ( .A(n998), .ZN(n714) );
  AOI22_X1 U215 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U216 ( .A(n951), .ZN(n673) );
  AOI22_X1 U217 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U218 ( .A(n949), .ZN(n672) );
  AOI22_X1 U219 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U220 ( .A(n948), .ZN(n671) );
  AOI22_X1 U221 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U222 ( .A(n947), .ZN(n670) );
  AOI22_X1 U223 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U224 ( .A(n946), .ZN(n669) );
  AOI22_X1 U225 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U226 ( .A(n945), .ZN(n668) );
  AOI22_X1 U227 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U228 ( .A(n944), .ZN(n667) );
  AOI22_X1 U229 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U230 ( .A(n943), .ZN(n666) );
  AOI22_X1 U231 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U232 ( .A(n915), .ZN(n641) );
  AOI22_X1 U233 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U234 ( .A(n979), .ZN(n697) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U236 ( .A(n977), .ZN(n696) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U238 ( .A(n976), .ZN(n695) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U240 ( .A(n975), .ZN(n694) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U242 ( .A(n974), .ZN(n693) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U244 ( .A(n973), .ZN(n692) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U246 ( .A(n972), .ZN(n691) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U248 ( .A(n971), .ZN(n690) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U250 ( .A(n970), .ZN(n689) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U252 ( .A(n968), .ZN(n688) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U254 ( .A(n967), .ZN(n687) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U256 ( .A(n966), .ZN(n686) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U258 ( .A(n965), .ZN(n685) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U260 ( .A(n964), .ZN(n684) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U262 ( .A(n963), .ZN(n683) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U264 ( .A(n962), .ZN(n682) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U266 ( .A(n942), .ZN(n665) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U268 ( .A(n940), .ZN(n664) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U270 ( .A(n939), .ZN(n663) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U272 ( .A(n938), .ZN(n662) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U274 ( .A(n937), .ZN(n661) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U276 ( .A(n936), .ZN(n660) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U278 ( .A(n935), .ZN(n659) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U280 ( .A(n934), .ZN(n658) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U282 ( .A(n933), .ZN(n657) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U284 ( .A(n931), .ZN(n656) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U286 ( .A(n930), .ZN(n655) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U288 ( .A(n929), .ZN(n654) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U290 ( .A(n928), .ZN(n653) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U292 ( .A(n927), .ZN(n652) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U294 ( .A(n926), .ZN(n651) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U296 ( .A(n925), .ZN(n650) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U298 ( .A(n906), .ZN(n633) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U300 ( .A(n904), .ZN(n632) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U302 ( .A(n903), .ZN(n631) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U304 ( .A(n902), .ZN(n630) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U306 ( .A(n901), .ZN(n629) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U308 ( .A(n900), .ZN(n628) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U310 ( .A(n899), .ZN(n627) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U312 ( .A(n898), .ZN(n626) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U314 ( .A(n897), .ZN(n625) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U316 ( .A(n895), .ZN(n624) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U318 ( .A(n894), .ZN(n623) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U320 ( .A(n893), .ZN(n622) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U322 ( .A(n892), .ZN(n621) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U324 ( .A(n891), .ZN(n620) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U326 ( .A(n890), .ZN(n619) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U328 ( .A(n889), .ZN(n618) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U330 ( .A(N12), .ZN(n253) );
  INV_X1 U331 ( .A(N11), .ZN(n252) );
  INV_X1 U332 ( .A(n997), .ZN(n713) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U334 ( .A(n995), .ZN(n712) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U336 ( .A(n994), .ZN(n711) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U338 ( .A(n993), .ZN(n710) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U340 ( .A(n992), .ZN(n709) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U342 ( .A(n991), .ZN(n708) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U344 ( .A(n990), .ZN(n707) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U346 ( .A(n989), .ZN(n706) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U348 ( .A(n924), .ZN(n649) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U350 ( .A(n922), .ZN(n648) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U352 ( .A(n921), .ZN(n647) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U354 ( .A(n920), .ZN(n646) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U356 ( .A(n919), .ZN(n645) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U358 ( .A(n918), .ZN(n644) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U360 ( .A(n917), .ZN(n643) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U362 ( .A(n916), .ZN(n642) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U364 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U366 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U368 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U370 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U372 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U374 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U376 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U378 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U380 ( .A(n961), .ZN(n681) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U382 ( .A(n959), .ZN(n680) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U384 ( .A(n958), .ZN(n679) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U386 ( .A(n957), .ZN(n678) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U388 ( .A(n956), .ZN(n677) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U390 ( .A(n955), .ZN(n676) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U392 ( .A(n954), .ZN(n675) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U394 ( .A(n953), .ZN(n674) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U396 ( .A(n888), .ZN(n617) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U398 ( .A(n886), .ZN(n616) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U400 ( .A(n885), .ZN(n615) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U402 ( .A(n884), .ZN(n614) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U404 ( .A(n883), .ZN(n613) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U406 ( .A(n882), .ZN(n612) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U408 ( .A(n881), .ZN(n611) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U410 ( .A(n880), .ZN(n610) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U412 ( .A(n879), .ZN(n609) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U414 ( .A(n877), .ZN(n608) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U416 ( .A(n876), .ZN(n607) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U418 ( .A(n875), .ZN(n606) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U420 ( .A(n874), .ZN(n605) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U422 ( .A(n873), .ZN(n604) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U424 ( .A(n872), .ZN(n603) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U426 ( .A(n871), .ZN(n602) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U428 ( .A(n870), .ZN(n601) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U430 ( .A(n868), .ZN(n600) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U432 ( .A(n867), .ZN(n599) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U434 ( .A(n866), .ZN(n598) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U436 ( .A(n865), .ZN(n597) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U438 ( .A(n864), .ZN(n596) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U440 ( .A(n863), .ZN(n595) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U442 ( .A(n862), .ZN(n594) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U444 ( .A(n861), .ZN(n293) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U446 ( .A(n859), .ZN(n292) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U448 ( .A(n858), .ZN(n291) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U450 ( .A(n857), .ZN(n290) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U452 ( .A(n856), .ZN(n289) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U454 ( .A(n855), .ZN(n288) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U456 ( .A(n854), .ZN(n287) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U458 ( .A(n853), .ZN(n286) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U460 ( .A(n852), .ZN(n285) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U462 ( .A(n850), .ZN(n284) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U464 ( .A(n849), .ZN(n283) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U466 ( .A(n848), .ZN(n282) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U468 ( .A(n847), .ZN(n281) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U470 ( .A(n846), .ZN(n280) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U472 ( .A(n845), .ZN(n279) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U474 ( .A(n844), .ZN(n278) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U476 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U477 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U478 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U479 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U480 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U481 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U482 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U483 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U484 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U485 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U486 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U487 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U488 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U489 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U490 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U491 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U492 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U494 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U496 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U498 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U500 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U502 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U504 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U506 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U508 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U510 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U512 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U514 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U516 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U518 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U520 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U522 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U524 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U526 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U528 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U530 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U532 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U534 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U536 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U538 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U540 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U542 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U544 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U546 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U548 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U550 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U552 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U554 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U556 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U558 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U560 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U562 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U564 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U566 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U568 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U570 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U572 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U574 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U576 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U578 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U580 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U582 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U584 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U586 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U588 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U590 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U592 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U594 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U596 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U598 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U600 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U602 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U604 ( .A(N13), .ZN(n842) );
  INV_X1 U605 ( .A(N14), .ZN(n843) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n248), .Z(n1) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n248), .Z(n2) );
  MUX2_X1 U608 ( .A(n2), .B(n1), .S(n243), .Z(n3) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n248), .Z(n4) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n248), .Z(n5) );
  MUX2_X1 U611 ( .A(n5), .B(n4), .S(n243), .Z(n6) );
  MUX2_X1 U612 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n248), .Z(n8) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n248), .Z(n9) );
  MUX2_X1 U615 ( .A(n9), .B(n8), .S(N11), .Z(n10) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n248), .Z(n11) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n248), .Z(n12) );
  MUX2_X1 U618 ( .A(n12), .B(n11), .S(N11), .Z(n13) );
  MUX2_X1 U619 ( .A(n13), .B(n10), .S(n241), .Z(n14) );
  MUX2_X1 U620 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n245), .Z(n16) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n245), .Z(n17) );
  MUX2_X1 U623 ( .A(n17), .B(n16), .S(n244), .Z(n18) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n245), .Z(n20) );
  MUX2_X1 U626 ( .A(n20), .B(n19), .S(n242), .Z(n21) );
  MUX2_X1 U627 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n245), .Z(n23) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n245), .Z(n24) );
  MUX2_X1 U630 ( .A(n24), .B(n23), .S(N11), .Z(n25) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n245), .Z(n26) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n245), .Z(n27) );
  MUX2_X1 U633 ( .A(n27), .B(n26), .S(n244), .Z(n28) );
  MUX2_X1 U634 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U635 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U636 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n245), .Z(n31) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n245), .Z(n32) );
  MUX2_X1 U639 ( .A(n32), .B(n31), .S(n242), .Z(n33) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U642 ( .A(n35), .B(n34), .S(n242), .Z(n36) );
  MUX2_X1 U643 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n247), .Z(n38) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n246), .Z(n39) );
  MUX2_X1 U646 ( .A(n39), .B(n38), .S(n244), .Z(n40) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n249), .Z(n41) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n247), .Z(n42) );
  MUX2_X1 U649 ( .A(n42), .B(n41), .S(n244), .Z(n43) );
  MUX2_X1 U650 ( .A(n43), .B(n40), .S(n241), .Z(n44) );
  MUX2_X1 U651 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n249), .Z(n46) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n245), .Z(n47) );
  MUX2_X1 U654 ( .A(n47), .B(n46), .S(N11), .Z(n48) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n247), .Z(n49) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n246), .Z(n50) );
  MUX2_X1 U657 ( .A(n50), .B(n49), .S(n243), .Z(n51) );
  MUX2_X1 U658 ( .A(n51), .B(n48), .S(n241), .Z(n52) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n246), .Z(n53) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n245), .Z(n54) );
  MUX2_X1 U661 ( .A(n54), .B(n53), .S(N11), .Z(n55) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n246), .Z(n56) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n249), .Z(n57) );
  MUX2_X1 U664 ( .A(n57), .B(n56), .S(N11), .Z(n58) );
  MUX2_X1 U665 ( .A(n58), .B(n55), .S(n241), .Z(n59) );
  MUX2_X1 U666 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U667 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n250), .Z(n61) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n245), .Z(n62) );
  MUX2_X1 U670 ( .A(n62), .B(n61), .S(n242), .Z(n63) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n246), .Z(n64) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n247), .Z(n65) );
  MUX2_X1 U673 ( .A(n65), .B(n64), .S(n242), .Z(n66) );
  MUX2_X1 U674 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n246), .Z(n68) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n245), .Z(n69) );
  MUX2_X1 U677 ( .A(n69), .B(n68), .S(n242), .Z(n70) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n249), .Z(n71) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n247), .Z(n72) );
  MUX2_X1 U680 ( .A(n72), .B(n71), .S(n242), .Z(n73) );
  MUX2_X1 U681 ( .A(n73), .B(n70), .S(N12), .Z(n74) );
  MUX2_X1 U682 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n247), .Z(n76) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n245), .Z(n77) );
  MUX2_X1 U685 ( .A(n77), .B(n76), .S(n242), .Z(n78) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n249), .Z(n79) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n245), .Z(n80) );
  MUX2_X1 U688 ( .A(n80), .B(n79), .S(n242), .Z(n81) );
  MUX2_X1 U689 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n250), .Z(n83) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n250), .Z(n84) );
  MUX2_X1 U692 ( .A(n84), .B(n83), .S(n242), .Z(n85) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n250), .Z(n86) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n250), .Z(n87) );
  MUX2_X1 U695 ( .A(n87), .B(n86), .S(n242), .Z(n88) );
  MUX2_X1 U696 ( .A(n88), .B(n85), .S(N12), .Z(n89) );
  MUX2_X1 U697 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U698 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n250), .Z(n91) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n92) );
  MUX2_X1 U701 ( .A(n92), .B(n91), .S(n242), .Z(n93) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n250), .Z(n95) );
  MUX2_X1 U704 ( .A(n95), .B(n94), .S(n242), .Z(n96) );
  MUX2_X1 U705 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n98) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n250), .Z(n99) );
  MUX2_X1 U708 ( .A(n99), .B(n98), .S(n242), .Z(n100) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n250), .Z(n101) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n250), .Z(n102) );
  MUX2_X1 U711 ( .A(n102), .B(n101), .S(n242), .Z(n103) );
  MUX2_X1 U712 ( .A(n103), .B(n100), .S(N12), .Z(n104) );
  MUX2_X1 U713 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n246), .Z(n106) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n246), .Z(n107) );
  MUX2_X1 U716 ( .A(n107), .B(n106), .S(n243), .Z(n108) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n246), .Z(n109) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n246), .Z(n110) );
  MUX2_X1 U719 ( .A(n110), .B(n109), .S(n243), .Z(n111) );
  MUX2_X1 U720 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n246), .Z(n113) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n246), .Z(n114) );
  MUX2_X1 U723 ( .A(n114), .B(n113), .S(n243), .Z(n115) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n246), .Z(n116) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n246), .Z(n117) );
  MUX2_X1 U726 ( .A(n117), .B(n116), .S(n243), .Z(n118) );
  MUX2_X1 U727 ( .A(n118), .B(n115), .S(N12), .Z(n119) );
  MUX2_X1 U728 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U729 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n246), .Z(n121) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n246), .Z(n122) );
  MUX2_X1 U732 ( .A(n122), .B(n121), .S(n243), .Z(n123) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n246), .Z(n124) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n246), .Z(n125) );
  MUX2_X1 U735 ( .A(n125), .B(n124), .S(n243), .Z(n126) );
  MUX2_X1 U736 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n247), .Z(n128) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n247), .Z(n129) );
  MUX2_X1 U739 ( .A(n129), .B(n128), .S(n243), .Z(n130) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n247), .Z(n131) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n247), .Z(n132) );
  MUX2_X1 U742 ( .A(n132), .B(n131), .S(n243), .Z(n133) );
  MUX2_X1 U743 ( .A(n133), .B(n130), .S(N12), .Z(n134) );
  MUX2_X1 U744 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n247), .Z(n136) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n247), .Z(n137) );
  MUX2_X1 U747 ( .A(n137), .B(n136), .S(n243), .Z(n138) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n247), .Z(n139) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n247), .Z(n140) );
  MUX2_X1 U750 ( .A(n140), .B(n139), .S(n243), .Z(n141) );
  MUX2_X1 U751 ( .A(n141), .B(n138), .S(n241), .Z(n142) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n247), .Z(n143) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n247), .Z(n144) );
  MUX2_X1 U754 ( .A(n144), .B(n143), .S(n243), .Z(n145) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n247), .Z(n146) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n247), .Z(n147) );
  MUX2_X1 U757 ( .A(n147), .B(n146), .S(n243), .Z(n148) );
  MUX2_X1 U758 ( .A(n148), .B(n145), .S(N12), .Z(n149) );
  MUX2_X1 U759 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U760 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n248), .Z(n151) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n248), .Z(n152) );
  MUX2_X1 U763 ( .A(n152), .B(n151), .S(n244), .Z(n153) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n248), .Z(n154) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n248), .Z(n155) );
  MUX2_X1 U766 ( .A(n155), .B(n154), .S(n244), .Z(n156) );
  MUX2_X1 U767 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n248), .Z(n158) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n248), .Z(n159) );
  MUX2_X1 U770 ( .A(n159), .B(n158), .S(n244), .Z(n160) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n248), .Z(n161) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n248), .Z(n162) );
  MUX2_X1 U773 ( .A(n162), .B(n161), .S(n244), .Z(n163) );
  MUX2_X1 U774 ( .A(n163), .B(n160), .S(N12), .Z(n164) );
  MUX2_X1 U775 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n248), .Z(n166) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n248), .Z(n167) );
  MUX2_X1 U778 ( .A(n167), .B(n166), .S(n244), .Z(n168) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n248), .Z(n169) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n248), .Z(n170) );
  MUX2_X1 U781 ( .A(n170), .B(n169), .S(n244), .Z(n171) );
  MUX2_X1 U782 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(N10), .Z(n173) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n250), .Z(n174) );
  MUX2_X1 U785 ( .A(n174), .B(n173), .S(n244), .Z(n175) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n176) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n250), .Z(n177) );
  MUX2_X1 U788 ( .A(n177), .B(n176), .S(n244), .Z(n178) );
  MUX2_X1 U789 ( .A(n178), .B(n175), .S(n241), .Z(n179) );
  MUX2_X1 U790 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U791 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n250), .Z(n181) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(N10), .Z(n182) );
  MUX2_X1 U794 ( .A(n182), .B(n181), .S(n244), .Z(n183) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(N10), .Z(n184) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(N10), .Z(n185) );
  MUX2_X1 U797 ( .A(n185), .B(n184), .S(n244), .Z(n186) );
  MUX2_X1 U798 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n250), .Z(n188) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(N10), .Z(n189) );
  MUX2_X1 U801 ( .A(n189), .B(n188), .S(n244), .Z(n190) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(N10), .Z(n191) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n250), .Z(n192) );
  MUX2_X1 U804 ( .A(n192), .B(n191), .S(n244), .Z(n193) );
  MUX2_X1 U805 ( .A(n193), .B(n190), .S(n241), .Z(n194) );
  MUX2_X1 U806 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n248), .Z(n196) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n250), .Z(n197) );
  MUX2_X1 U809 ( .A(n197), .B(n196), .S(N11), .Z(n198) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(N10), .Z(n199) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n200) );
  MUX2_X1 U812 ( .A(n200), .B(n199), .S(n244), .Z(n201) );
  MUX2_X1 U813 ( .A(n201), .B(n198), .S(n241), .Z(n202) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n203) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n204) );
  MUX2_X1 U816 ( .A(n204), .B(n203), .S(N11), .Z(n205) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n206) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n207) );
  MUX2_X1 U819 ( .A(n207), .B(n206), .S(n242), .Z(n208) );
  MUX2_X1 U820 ( .A(n208), .B(n205), .S(N12), .Z(n209) );
  MUX2_X1 U821 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U822 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n248), .Z(n211) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(N10), .Z(n212) );
  MUX2_X1 U825 ( .A(n212), .B(n211), .S(N11), .Z(n213) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n248), .Z(n214) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n250), .Z(n215) );
  MUX2_X1 U828 ( .A(n215), .B(n214), .S(N11), .Z(n216) );
  MUX2_X1 U829 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n249), .Z(n218) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n249), .Z(n219) );
  MUX2_X1 U832 ( .A(n219), .B(n218), .S(N11), .Z(n220) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n249), .Z(n221) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n249), .Z(n222) );
  MUX2_X1 U835 ( .A(n222), .B(n221), .S(n243), .Z(n223) );
  MUX2_X1 U836 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U837 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n249), .Z(n226) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n249), .Z(n227) );
  MUX2_X1 U840 ( .A(n227), .B(n226), .S(N11), .Z(n228) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n249), .Z(n229) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n249), .Z(n230) );
  MUX2_X1 U843 ( .A(n230), .B(n229), .S(n242), .Z(n231) );
  MUX2_X1 U844 ( .A(n231), .B(n228), .S(n241), .Z(n232) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n249), .Z(n233) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n249), .Z(n234) );
  MUX2_X1 U847 ( .A(n234), .B(n233), .S(N11), .Z(n235) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n249), .Z(n236) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n249), .Z(n237) );
  MUX2_X1 U850 ( .A(n237), .B(n236), .S(n243), .Z(n238) );
  MUX2_X1 U851 ( .A(n238), .B(n235), .S(n241), .Z(n239) );
  MUX2_X1 U852 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U853 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_31 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n256), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n257), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n258), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n259), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n260), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n261), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n262), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n263), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n264), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n265), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n266), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n267), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n268), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n269), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n270), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n271), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n272), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n273), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n274), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n275), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n276), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n277), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n278), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n279), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n280), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n281), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n282), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n283), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n284), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n285), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n286), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n287), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n288), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n289), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n290), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n291), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n292), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n293), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n594), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n595), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n596), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n597), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n598), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n599), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n600), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n601), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n602), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n603), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n604), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n605), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n606), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n607), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n608), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n609), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n610), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n611), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n612), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n613), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n614), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n615), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n616), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n617), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n618), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n619), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n620), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n621), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n622), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n623), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n624), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n625), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n626), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n627), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n628), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n629), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n630), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n631), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n632), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n633), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n634), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n635), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n636), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n637), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n638), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n639), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n640), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n641), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n642), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n643), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n644), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n645), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n646), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n647), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n648), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n649), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n650), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n651), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n652), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n653), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n654), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n655), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n656), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n657), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n658), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n659), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n660), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n661), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n662), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n663), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n664), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n665), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n666), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n667), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n668), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n669), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n670), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n671), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n672), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n673), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n674), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n675), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n676), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n677), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n678), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n679), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n680), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n681), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n682), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n683), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n684), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n685), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n686), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n687), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n688), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n689), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n690), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n691), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n692), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n693), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n694), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n695), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n696), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n697), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n698), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n699), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n700), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n701), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n702), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n703), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n704), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n705), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n706), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n707), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n708), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n709), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n710), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n711), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n712), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n713), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n714), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n715), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n716), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n717), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n718), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n719), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n720), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n721), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n722), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n723), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n724), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n725), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n726), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n727), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n728), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n729), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n730), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n731), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n732), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n733), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n734), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n735), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n736), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n737), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n738), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n739), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n740), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n741), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n742), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n743), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n744), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n745), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n746), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n747), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n748), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n749), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n750), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n751), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n752), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n753), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n754), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n755), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n756), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n757), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n758), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n759), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n760), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n761), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n762), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n763), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n764), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n765), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n766), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n767), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n768), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n769), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n770), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n771), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n772), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n773), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n774), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n775), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n776), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n777), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n778), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n779), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n780), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n781), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n782), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n783), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n784), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n785), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n786), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n787), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n788), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n789), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n790), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n791), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n792), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n793), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n794), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n795), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n796), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n797), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n798), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n799), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n800), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n801), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n802), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n803), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n804), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n805), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n806), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n807), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n808), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n809), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n810), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n811), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(n252), .Z(n251) );
  BUF_X1 U5 ( .A(n252), .Z(n247) );
  BUF_X1 U6 ( .A(n252), .Z(n248) );
  BUF_X1 U7 ( .A(n252), .Z(n249) );
  BUF_X1 U8 ( .A(n252), .Z(n250) );
  BUF_X1 U9 ( .A(N10), .Z(n252) );
  INV_X1 U10 ( .A(n1113), .ZN(n843) );
  INV_X1 U11 ( .A(n1102), .ZN(n842) );
  INV_X1 U12 ( .A(n1092), .ZN(n841) );
  INV_X1 U13 ( .A(n1082), .ZN(n840) );
  INV_X1 U14 ( .A(n1072), .ZN(n839) );
  INV_X1 U15 ( .A(n1062), .ZN(n838) );
  INV_X1 U16 ( .A(n1053), .ZN(n837) );
  INV_X1 U17 ( .A(n1044), .ZN(n836) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1105) );
  NOR3_X1 U19 ( .A1(N11), .A2(N12), .A3(n253), .ZN(n1094) );
  NAND2_X1 U20 ( .A1(n1104), .A2(n1136), .ZN(n1062) );
  NAND2_X1 U21 ( .A1(n1105), .A2(n1104), .ZN(n1113) );
  NAND2_X1 U22 ( .A1(n1094), .A2(n1104), .ZN(n1102) );
  NAND2_X1 U23 ( .A1(n1084), .A2(n1104), .ZN(n1092) );
  NAND2_X1 U24 ( .A1(n1074), .A2(n1104), .ZN(n1082) );
  NAND2_X1 U25 ( .A1(n1064), .A2(n1104), .ZN(n1072) );
  NAND2_X1 U26 ( .A1(n1104), .A2(n1125), .ZN(n1053) );
  NAND2_X1 U27 ( .A1(n1104), .A2(n1115), .ZN(n1044) );
  INV_X1 U28 ( .A(n1133), .ZN(n818) );
  INV_X1 U29 ( .A(n1123), .ZN(n817) );
  INV_X1 U30 ( .A(n889), .ZN(n816) );
  INV_X1 U31 ( .A(n880), .ZN(n815) );
  INV_X1 U32 ( .A(n871), .ZN(n814) );
  INV_X1 U33 ( .A(n862), .ZN(n813) );
  INV_X1 U34 ( .A(n853), .ZN(n812) );
  INV_X1 U35 ( .A(n989), .ZN(n830) );
  INV_X1 U36 ( .A(n980), .ZN(n829) );
  INV_X1 U37 ( .A(n971), .ZN(n828) );
  INV_X1 U38 ( .A(n916), .ZN(n822) );
  INV_X1 U39 ( .A(n907), .ZN(n821) );
  INV_X1 U40 ( .A(n898), .ZN(n820) );
  INV_X1 U41 ( .A(n1035), .ZN(n835) );
  INV_X1 U42 ( .A(n1025), .ZN(n834) );
  INV_X1 U43 ( .A(n1016), .ZN(n833) );
  INV_X1 U44 ( .A(n1007), .ZN(n832) );
  INV_X1 U45 ( .A(n998), .ZN(n831) );
  INV_X1 U46 ( .A(n962), .ZN(n827) );
  INV_X1 U47 ( .A(n952), .ZN(n826) );
  INV_X1 U48 ( .A(n943), .ZN(n825) );
  INV_X1 U49 ( .A(n934), .ZN(n824) );
  INV_X1 U50 ( .A(n925), .ZN(n823) );
  INV_X1 U51 ( .A(n1144), .ZN(n819) );
  BUF_X1 U52 ( .A(N11), .Z(n244) );
  BUF_X1 U53 ( .A(N11), .Z(n245) );
  BUF_X1 U54 ( .A(N11), .Z(n246) );
  INV_X1 U55 ( .A(N10), .ZN(n253) );
  BUF_X1 U56 ( .A(N12), .Z(n243) );
  NOR3_X1 U57 ( .A1(n255), .A2(N10), .A3(n254), .ZN(n1125) );
  NOR3_X1 U58 ( .A1(n255), .A2(n253), .A3(n254), .ZN(n1115) );
  NOR3_X1 U59 ( .A1(n253), .A2(N11), .A3(n255), .ZN(n1136) );
  NOR3_X1 U60 ( .A1(N10), .A2(N12), .A3(n254), .ZN(n1084) );
  NOR3_X1 U61 ( .A1(n253), .A2(N12), .A3(n254), .ZN(n1074) );
  NOR3_X1 U62 ( .A1(N10), .A2(N11), .A3(n255), .ZN(n1064) );
  NAND2_X1 U63 ( .A1(n1027), .A2(n1136), .ZN(n989) );
  NAND2_X1 U64 ( .A1(n954), .A2(n1136), .ZN(n916) );
  NAND2_X1 U65 ( .A1(n1027), .A2(n1064), .ZN(n998) );
  NAND2_X1 U66 ( .A1(n954), .A2(n1064), .ZN(n925) );
  NAND2_X1 U67 ( .A1(n1027), .A2(n1105), .ZN(n1035) );
  NAND2_X1 U68 ( .A1(n1027), .A2(n1094), .ZN(n1025) );
  NAND2_X1 U69 ( .A1(n954), .A2(n1105), .ZN(n962) );
  NAND2_X1 U70 ( .A1(n954), .A2(n1094), .ZN(n952) );
  NAND2_X1 U71 ( .A1(n1105), .A2(n1135), .ZN(n889) );
  NAND2_X1 U72 ( .A1(n1094), .A2(n1135), .ZN(n880) );
  NAND2_X1 U73 ( .A1(n1084), .A2(n1135), .ZN(n871) );
  NAND2_X1 U74 ( .A1(n1074), .A2(n1135), .ZN(n862) );
  NAND2_X1 U75 ( .A1(n1064), .A2(n1135), .ZN(n853) );
  NAND2_X1 U76 ( .A1(n1136), .A2(n1135), .ZN(n1144) );
  NAND2_X1 U77 ( .A1(n1125), .A2(n1135), .ZN(n1133) );
  NAND2_X1 U78 ( .A1(n1115), .A2(n1135), .ZN(n1123) );
  NAND2_X1 U79 ( .A1(n1027), .A2(n1084), .ZN(n1016) );
  NAND2_X1 U80 ( .A1(n1027), .A2(n1074), .ZN(n1007) );
  NAND2_X1 U81 ( .A1(n954), .A2(n1084), .ZN(n943) );
  NAND2_X1 U82 ( .A1(n954), .A2(n1074), .ZN(n934) );
  NAND2_X1 U83 ( .A1(n1027), .A2(n1125), .ZN(n980) );
  NAND2_X1 U84 ( .A1(n954), .A2(n1125), .ZN(n907) );
  NAND2_X1 U85 ( .A1(n1027), .A2(n1115), .ZN(n971) );
  NAND2_X1 U86 ( .A1(n954), .A2(n1115), .ZN(n898) );
  AND3_X1 U87 ( .A1(n844), .A2(n845), .A3(wr_en), .ZN(n1104) );
  AND3_X1 U88 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1135) );
  AND3_X1 U89 ( .A1(N13), .A2(n845), .A3(wr_en), .ZN(n1027) );
  AND3_X1 U90 ( .A1(N14), .A2(n844), .A3(wr_en), .ZN(n954) );
  INV_X1 U91 ( .A(n1063), .ZN(n771) );
  AOI22_X1 U92 ( .A1(data_in[0]), .A2(n838), .B1(n1062), .B2(\mem[5][0] ), 
        .ZN(n1063) );
  INV_X1 U93 ( .A(n1061), .ZN(n770) );
  AOI22_X1 U94 ( .A1(data_in[1]), .A2(n838), .B1(n1062), .B2(\mem[5][1] ), 
        .ZN(n1061) );
  INV_X1 U95 ( .A(n1060), .ZN(n769) );
  AOI22_X1 U96 ( .A1(data_in[2]), .A2(n838), .B1(n1062), .B2(\mem[5][2] ), 
        .ZN(n1060) );
  INV_X1 U97 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U98 ( .A1(data_in[3]), .A2(n838), .B1(n1062), .B2(\mem[5][3] ), 
        .ZN(n1059) );
  INV_X1 U99 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U100 ( .A1(data_in[4]), .A2(n838), .B1(n1062), .B2(\mem[5][4] ), 
        .ZN(n1058) );
  INV_X1 U101 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U102 ( .A1(data_in[5]), .A2(n838), .B1(n1062), .B2(\mem[5][5] ), 
        .ZN(n1057) );
  INV_X1 U103 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U104 ( .A1(data_in[6]), .A2(n838), .B1(n1062), .B2(\mem[5][6] ), 
        .ZN(n1056) );
  INV_X1 U105 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U106 ( .A1(data_in[7]), .A2(n838), .B1(n1062), .B2(\mem[5][7] ), 
        .ZN(n1055) );
  INV_X1 U107 ( .A(n1026), .ZN(n739) );
  AOI22_X1 U108 ( .A1(data_in[0]), .A2(n834), .B1(n1025), .B2(\mem[9][0] ), 
        .ZN(n1026) );
  INV_X1 U109 ( .A(n1024), .ZN(n738) );
  AOI22_X1 U110 ( .A1(data_in[1]), .A2(n834), .B1(n1025), .B2(\mem[9][1] ), 
        .ZN(n1024) );
  INV_X1 U111 ( .A(n1023), .ZN(n737) );
  AOI22_X1 U112 ( .A1(data_in[2]), .A2(n834), .B1(n1025), .B2(\mem[9][2] ), 
        .ZN(n1023) );
  INV_X1 U113 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U114 ( .A1(data_in[3]), .A2(n834), .B1(n1025), .B2(\mem[9][3] ), 
        .ZN(n1022) );
  INV_X1 U115 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U116 ( .A1(data_in[4]), .A2(n834), .B1(n1025), .B2(\mem[9][4] ), 
        .ZN(n1021) );
  INV_X1 U117 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U118 ( .A1(data_in[5]), .A2(n834), .B1(n1025), .B2(\mem[9][5] ), 
        .ZN(n1020) );
  INV_X1 U119 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U120 ( .A1(data_in[6]), .A2(n834), .B1(n1025), .B2(\mem[9][6] ), 
        .ZN(n1019) );
  INV_X1 U121 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U122 ( .A1(data_in[7]), .A2(n834), .B1(n1025), .B2(\mem[9][7] ), 
        .ZN(n1018) );
  INV_X1 U123 ( .A(n990), .ZN(n707) );
  AOI22_X1 U124 ( .A1(data_in[0]), .A2(n830), .B1(n989), .B2(\mem[13][0] ), 
        .ZN(n990) );
  INV_X1 U125 ( .A(n988), .ZN(n706) );
  AOI22_X1 U126 ( .A1(data_in[1]), .A2(n830), .B1(n989), .B2(\mem[13][1] ), 
        .ZN(n988) );
  INV_X1 U127 ( .A(n987), .ZN(n705) );
  AOI22_X1 U128 ( .A1(data_in[2]), .A2(n830), .B1(n989), .B2(\mem[13][2] ), 
        .ZN(n987) );
  INV_X1 U129 ( .A(n986), .ZN(n704) );
  AOI22_X1 U130 ( .A1(data_in[3]), .A2(n830), .B1(n989), .B2(\mem[13][3] ), 
        .ZN(n986) );
  INV_X1 U131 ( .A(n985), .ZN(n703) );
  AOI22_X1 U132 ( .A1(data_in[4]), .A2(n830), .B1(n989), .B2(\mem[13][4] ), 
        .ZN(n985) );
  INV_X1 U133 ( .A(n984), .ZN(n702) );
  AOI22_X1 U134 ( .A1(data_in[5]), .A2(n830), .B1(n989), .B2(\mem[13][5] ), 
        .ZN(n984) );
  INV_X1 U135 ( .A(n983), .ZN(n701) );
  AOI22_X1 U136 ( .A1(data_in[6]), .A2(n830), .B1(n989), .B2(\mem[13][6] ), 
        .ZN(n983) );
  INV_X1 U137 ( .A(n982), .ZN(n700) );
  AOI22_X1 U138 ( .A1(data_in[7]), .A2(n830), .B1(n989), .B2(\mem[13][7] ), 
        .ZN(n982) );
  INV_X1 U139 ( .A(n953), .ZN(n675) );
  AOI22_X1 U140 ( .A1(data_in[0]), .A2(n826), .B1(n952), .B2(\mem[17][0] ), 
        .ZN(n953) );
  INV_X1 U141 ( .A(n951), .ZN(n674) );
  AOI22_X1 U142 ( .A1(data_in[1]), .A2(n826), .B1(n952), .B2(\mem[17][1] ), 
        .ZN(n951) );
  INV_X1 U143 ( .A(n950), .ZN(n673) );
  AOI22_X1 U144 ( .A1(data_in[2]), .A2(n826), .B1(n952), .B2(\mem[17][2] ), 
        .ZN(n950) );
  INV_X1 U145 ( .A(n949), .ZN(n672) );
  AOI22_X1 U146 ( .A1(data_in[3]), .A2(n826), .B1(n952), .B2(\mem[17][3] ), 
        .ZN(n949) );
  INV_X1 U147 ( .A(n948), .ZN(n671) );
  AOI22_X1 U148 ( .A1(data_in[4]), .A2(n826), .B1(n952), .B2(\mem[17][4] ), 
        .ZN(n948) );
  INV_X1 U149 ( .A(n947), .ZN(n670) );
  AOI22_X1 U150 ( .A1(data_in[5]), .A2(n826), .B1(n952), .B2(\mem[17][5] ), 
        .ZN(n947) );
  INV_X1 U151 ( .A(n946), .ZN(n669) );
  AOI22_X1 U152 ( .A1(data_in[6]), .A2(n826), .B1(n952), .B2(\mem[17][6] ), 
        .ZN(n946) );
  INV_X1 U153 ( .A(n945), .ZN(n668) );
  AOI22_X1 U154 ( .A1(data_in[7]), .A2(n826), .B1(n952), .B2(\mem[17][7] ), 
        .ZN(n945) );
  INV_X1 U155 ( .A(n917), .ZN(n643) );
  AOI22_X1 U156 ( .A1(data_in[0]), .A2(n822), .B1(n916), .B2(\mem[21][0] ), 
        .ZN(n917) );
  INV_X1 U157 ( .A(n915), .ZN(n642) );
  AOI22_X1 U158 ( .A1(data_in[1]), .A2(n822), .B1(n916), .B2(\mem[21][1] ), 
        .ZN(n915) );
  INV_X1 U159 ( .A(n914), .ZN(n641) );
  AOI22_X1 U160 ( .A1(data_in[2]), .A2(n822), .B1(n916), .B2(\mem[21][2] ), 
        .ZN(n914) );
  INV_X1 U161 ( .A(n913), .ZN(n640) );
  AOI22_X1 U162 ( .A1(data_in[3]), .A2(n822), .B1(n916), .B2(\mem[21][3] ), 
        .ZN(n913) );
  INV_X1 U163 ( .A(n912), .ZN(n639) );
  AOI22_X1 U164 ( .A1(data_in[4]), .A2(n822), .B1(n916), .B2(\mem[21][4] ), 
        .ZN(n912) );
  INV_X1 U165 ( .A(n911), .ZN(n638) );
  AOI22_X1 U166 ( .A1(data_in[5]), .A2(n822), .B1(n916), .B2(\mem[21][5] ), 
        .ZN(n911) );
  INV_X1 U167 ( .A(n910), .ZN(n637) );
  AOI22_X1 U168 ( .A1(data_in[6]), .A2(n822), .B1(n916), .B2(\mem[21][6] ), 
        .ZN(n910) );
  INV_X1 U169 ( .A(n909), .ZN(n636) );
  AOI22_X1 U170 ( .A1(data_in[7]), .A2(n822), .B1(n916), .B2(\mem[21][7] ), 
        .ZN(n909) );
  INV_X1 U171 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U172 ( .A1(data_in[0]), .A2(n837), .B1(n1053), .B2(\mem[6][0] ), 
        .ZN(n1054) );
  INV_X1 U173 ( .A(n1052), .ZN(n762) );
  AOI22_X1 U174 ( .A1(data_in[1]), .A2(n837), .B1(n1053), .B2(\mem[6][1] ), 
        .ZN(n1052) );
  INV_X1 U175 ( .A(n1051), .ZN(n761) );
  AOI22_X1 U176 ( .A1(data_in[2]), .A2(n837), .B1(n1053), .B2(\mem[6][2] ), 
        .ZN(n1051) );
  INV_X1 U177 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U178 ( .A1(data_in[3]), .A2(n837), .B1(n1053), .B2(\mem[6][3] ), 
        .ZN(n1050) );
  INV_X1 U179 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U180 ( .A1(data_in[4]), .A2(n837), .B1(n1053), .B2(\mem[6][4] ), 
        .ZN(n1049) );
  INV_X1 U181 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U182 ( .A1(data_in[5]), .A2(n837), .B1(n1053), .B2(\mem[6][5] ), 
        .ZN(n1048) );
  INV_X1 U183 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U184 ( .A1(data_in[6]), .A2(n837), .B1(n1053), .B2(\mem[6][6] ), 
        .ZN(n1047) );
  INV_X1 U185 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U186 ( .A1(data_in[7]), .A2(n837), .B1(n1053), .B2(\mem[6][7] ), 
        .ZN(n1046) );
  INV_X1 U187 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U188 ( .A1(data_in[0]), .A2(n836), .B1(n1044), .B2(\mem[7][0] ), 
        .ZN(n1045) );
  INV_X1 U189 ( .A(n1043), .ZN(n754) );
  AOI22_X1 U190 ( .A1(data_in[1]), .A2(n836), .B1(n1044), .B2(\mem[7][1] ), 
        .ZN(n1043) );
  INV_X1 U191 ( .A(n1042), .ZN(n753) );
  AOI22_X1 U192 ( .A1(data_in[2]), .A2(n836), .B1(n1044), .B2(\mem[7][2] ), 
        .ZN(n1042) );
  INV_X1 U193 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U194 ( .A1(data_in[3]), .A2(n836), .B1(n1044), .B2(\mem[7][3] ), 
        .ZN(n1041) );
  INV_X1 U195 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U196 ( .A1(data_in[4]), .A2(n836), .B1(n1044), .B2(\mem[7][4] ), 
        .ZN(n1040) );
  INV_X1 U197 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U198 ( .A1(data_in[5]), .A2(n836), .B1(n1044), .B2(\mem[7][5] ), 
        .ZN(n1039) );
  INV_X1 U199 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U200 ( .A1(data_in[6]), .A2(n836), .B1(n1044), .B2(\mem[7][6] ), 
        .ZN(n1038) );
  INV_X1 U201 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U202 ( .A1(data_in[7]), .A2(n836), .B1(n1044), .B2(\mem[7][7] ), 
        .ZN(n1037) );
  INV_X1 U203 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U204 ( .A1(data_in[0]), .A2(n833), .B1(n1016), .B2(\mem[10][0] ), 
        .ZN(n1017) );
  INV_X1 U205 ( .A(n1015), .ZN(n730) );
  AOI22_X1 U206 ( .A1(data_in[1]), .A2(n833), .B1(n1016), .B2(\mem[10][1] ), 
        .ZN(n1015) );
  INV_X1 U207 ( .A(n1014), .ZN(n729) );
  AOI22_X1 U208 ( .A1(data_in[2]), .A2(n833), .B1(n1016), .B2(\mem[10][2] ), 
        .ZN(n1014) );
  INV_X1 U209 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U210 ( .A1(data_in[3]), .A2(n833), .B1(n1016), .B2(\mem[10][3] ), 
        .ZN(n1013) );
  INV_X1 U211 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U212 ( .A1(data_in[4]), .A2(n833), .B1(n1016), .B2(\mem[10][4] ), 
        .ZN(n1012) );
  INV_X1 U213 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U214 ( .A1(data_in[5]), .A2(n833), .B1(n1016), .B2(\mem[10][5] ), 
        .ZN(n1011) );
  INV_X1 U215 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U216 ( .A1(data_in[6]), .A2(n833), .B1(n1016), .B2(\mem[10][6] ), 
        .ZN(n1010) );
  INV_X1 U217 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U218 ( .A1(data_in[7]), .A2(n833), .B1(n1016), .B2(\mem[10][7] ), 
        .ZN(n1009) );
  INV_X1 U219 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U220 ( .A1(data_in[0]), .A2(n832), .B1(n1007), .B2(\mem[11][0] ), 
        .ZN(n1008) );
  INV_X1 U221 ( .A(n1006), .ZN(n722) );
  AOI22_X1 U222 ( .A1(data_in[1]), .A2(n832), .B1(n1007), .B2(\mem[11][1] ), 
        .ZN(n1006) );
  INV_X1 U223 ( .A(n1005), .ZN(n721) );
  AOI22_X1 U224 ( .A1(data_in[2]), .A2(n832), .B1(n1007), .B2(\mem[11][2] ), 
        .ZN(n1005) );
  INV_X1 U225 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U226 ( .A1(data_in[3]), .A2(n832), .B1(n1007), .B2(\mem[11][3] ), 
        .ZN(n1004) );
  INV_X1 U227 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U228 ( .A1(data_in[4]), .A2(n832), .B1(n1007), .B2(\mem[11][4] ), 
        .ZN(n1003) );
  INV_X1 U229 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U230 ( .A1(data_in[5]), .A2(n832), .B1(n1007), .B2(\mem[11][5] ), 
        .ZN(n1002) );
  INV_X1 U231 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U232 ( .A1(data_in[6]), .A2(n832), .B1(n1007), .B2(\mem[11][6] ), 
        .ZN(n1001) );
  INV_X1 U233 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U234 ( .A1(data_in[7]), .A2(n832), .B1(n1007), .B2(\mem[11][7] ), 
        .ZN(n1000) );
  INV_X1 U235 ( .A(n937), .ZN(n661) );
  AOI22_X1 U236 ( .A1(data_in[6]), .A2(n825), .B1(n943), .B2(\mem[18][6] ), 
        .ZN(n937) );
  INV_X1 U237 ( .A(n936), .ZN(n660) );
  AOI22_X1 U238 ( .A1(data_in[7]), .A2(n825), .B1(n943), .B2(\mem[18][7] ), 
        .ZN(n936) );
  INV_X1 U239 ( .A(n935), .ZN(n659) );
  AOI22_X1 U240 ( .A1(data_in[0]), .A2(n824), .B1(n934), .B2(\mem[19][0] ), 
        .ZN(n935) );
  INV_X1 U241 ( .A(n933), .ZN(n658) );
  AOI22_X1 U242 ( .A1(data_in[1]), .A2(n824), .B1(n934), .B2(\mem[19][1] ), 
        .ZN(n933) );
  INV_X1 U243 ( .A(n932), .ZN(n657) );
  AOI22_X1 U244 ( .A1(data_in[2]), .A2(n824), .B1(n934), .B2(\mem[19][2] ), 
        .ZN(n932) );
  INV_X1 U245 ( .A(n931), .ZN(n656) );
  AOI22_X1 U246 ( .A1(data_in[3]), .A2(n824), .B1(n934), .B2(\mem[19][3] ), 
        .ZN(n931) );
  INV_X1 U247 ( .A(n930), .ZN(n655) );
  AOI22_X1 U248 ( .A1(data_in[4]), .A2(n824), .B1(n934), .B2(\mem[19][4] ), 
        .ZN(n930) );
  INV_X1 U249 ( .A(n929), .ZN(n654) );
  AOI22_X1 U250 ( .A1(data_in[5]), .A2(n824), .B1(n934), .B2(\mem[19][5] ), 
        .ZN(n929) );
  INV_X1 U251 ( .A(n981), .ZN(n699) );
  AOI22_X1 U252 ( .A1(data_in[0]), .A2(n829), .B1(n980), .B2(\mem[14][0] ), 
        .ZN(n981) );
  INV_X1 U253 ( .A(n979), .ZN(n698) );
  AOI22_X1 U254 ( .A1(data_in[1]), .A2(n829), .B1(n980), .B2(\mem[14][1] ), 
        .ZN(n979) );
  INV_X1 U255 ( .A(n978), .ZN(n697) );
  AOI22_X1 U256 ( .A1(data_in[2]), .A2(n829), .B1(n980), .B2(\mem[14][2] ), 
        .ZN(n978) );
  INV_X1 U257 ( .A(n977), .ZN(n696) );
  AOI22_X1 U258 ( .A1(data_in[3]), .A2(n829), .B1(n980), .B2(\mem[14][3] ), 
        .ZN(n977) );
  INV_X1 U259 ( .A(n976), .ZN(n695) );
  AOI22_X1 U260 ( .A1(data_in[4]), .A2(n829), .B1(n980), .B2(\mem[14][4] ), 
        .ZN(n976) );
  INV_X1 U261 ( .A(n975), .ZN(n694) );
  AOI22_X1 U262 ( .A1(data_in[5]), .A2(n829), .B1(n980), .B2(\mem[14][5] ), 
        .ZN(n975) );
  INV_X1 U263 ( .A(n974), .ZN(n693) );
  AOI22_X1 U264 ( .A1(data_in[6]), .A2(n829), .B1(n980), .B2(\mem[14][6] ), 
        .ZN(n974) );
  INV_X1 U265 ( .A(n973), .ZN(n692) );
  AOI22_X1 U266 ( .A1(data_in[7]), .A2(n829), .B1(n980), .B2(\mem[14][7] ), 
        .ZN(n973) );
  INV_X1 U267 ( .A(n972), .ZN(n691) );
  AOI22_X1 U268 ( .A1(data_in[0]), .A2(n828), .B1(n971), .B2(\mem[15][0] ), 
        .ZN(n972) );
  INV_X1 U269 ( .A(n970), .ZN(n690) );
  AOI22_X1 U270 ( .A1(data_in[1]), .A2(n828), .B1(n971), .B2(\mem[15][1] ), 
        .ZN(n970) );
  INV_X1 U271 ( .A(n969), .ZN(n689) );
  AOI22_X1 U272 ( .A1(data_in[2]), .A2(n828), .B1(n971), .B2(\mem[15][2] ), 
        .ZN(n969) );
  INV_X1 U273 ( .A(n968), .ZN(n688) );
  AOI22_X1 U274 ( .A1(data_in[3]), .A2(n828), .B1(n971), .B2(\mem[15][3] ), 
        .ZN(n968) );
  INV_X1 U275 ( .A(n967), .ZN(n687) );
  AOI22_X1 U276 ( .A1(data_in[4]), .A2(n828), .B1(n971), .B2(\mem[15][4] ), 
        .ZN(n967) );
  INV_X1 U277 ( .A(n966), .ZN(n686) );
  AOI22_X1 U278 ( .A1(data_in[5]), .A2(n828), .B1(n971), .B2(\mem[15][5] ), 
        .ZN(n966) );
  INV_X1 U279 ( .A(n965), .ZN(n685) );
  AOI22_X1 U280 ( .A1(data_in[6]), .A2(n828), .B1(n971), .B2(\mem[15][6] ), 
        .ZN(n965) );
  INV_X1 U281 ( .A(n964), .ZN(n684) );
  AOI22_X1 U282 ( .A1(data_in[7]), .A2(n828), .B1(n971), .B2(\mem[15][7] ), 
        .ZN(n964) );
  INV_X1 U283 ( .A(n944), .ZN(n667) );
  AOI22_X1 U284 ( .A1(data_in[0]), .A2(n825), .B1(n943), .B2(\mem[18][0] ), 
        .ZN(n944) );
  INV_X1 U285 ( .A(n942), .ZN(n666) );
  AOI22_X1 U286 ( .A1(data_in[1]), .A2(n825), .B1(n943), .B2(\mem[18][1] ), 
        .ZN(n942) );
  INV_X1 U287 ( .A(n941), .ZN(n665) );
  AOI22_X1 U288 ( .A1(data_in[2]), .A2(n825), .B1(n943), .B2(\mem[18][2] ), 
        .ZN(n941) );
  INV_X1 U289 ( .A(n940), .ZN(n664) );
  AOI22_X1 U290 ( .A1(data_in[3]), .A2(n825), .B1(n943), .B2(\mem[18][3] ), 
        .ZN(n940) );
  INV_X1 U291 ( .A(n939), .ZN(n663) );
  AOI22_X1 U292 ( .A1(data_in[4]), .A2(n825), .B1(n943), .B2(\mem[18][4] ), 
        .ZN(n939) );
  INV_X1 U293 ( .A(n938), .ZN(n662) );
  AOI22_X1 U294 ( .A1(data_in[5]), .A2(n825), .B1(n943), .B2(\mem[18][5] ), 
        .ZN(n938) );
  INV_X1 U295 ( .A(n928), .ZN(n653) );
  AOI22_X1 U296 ( .A1(data_in[6]), .A2(n824), .B1(n934), .B2(\mem[19][6] ), 
        .ZN(n928) );
  INV_X1 U297 ( .A(n927), .ZN(n652) );
  AOI22_X1 U298 ( .A1(data_in[7]), .A2(n824), .B1(n934), .B2(\mem[19][7] ), 
        .ZN(n927) );
  INV_X1 U299 ( .A(n908), .ZN(n635) );
  AOI22_X1 U300 ( .A1(data_in[0]), .A2(n821), .B1(n907), .B2(\mem[22][0] ), 
        .ZN(n908) );
  INV_X1 U301 ( .A(n906), .ZN(n634) );
  AOI22_X1 U302 ( .A1(data_in[1]), .A2(n821), .B1(n907), .B2(\mem[22][1] ), 
        .ZN(n906) );
  INV_X1 U303 ( .A(n905), .ZN(n633) );
  AOI22_X1 U304 ( .A1(data_in[2]), .A2(n821), .B1(n907), .B2(\mem[22][2] ), 
        .ZN(n905) );
  INV_X1 U305 ( .A(n904), .ZN(n632) );
  AOI22_X1 U306 ( .A1(data_in[3]), .A2(n821), .B1(n907), .B2(\mem[22][3] ), 
        .ZN(n904) );
  INV_X1 U307 ( .A(n903), .ZN(n631) );
  AOI22_X1 U308 ( .A1(data_in[4]), .A2(n821), .B1(n907), .B2(\mem[22][4] ), 
        .ZN(n903) );
  INV_X1 U309 ( .A(n902), .ZN(n630) );
  AOI22_X1 U310 ( .A1(data_in[5]), .A2(n821), .B1(n907), .B2(\mem[22][5] ), 
        .ZN(n902) );
  INV_X1 U311 ( .A(n901), .ZN(n629) );
  AOI22_X1 U312 ( .A1(data_in[6]), .A2(n821), .B1(n907), .B2(\mem[22][6] ), 
        .ZN(n901) );
  INV_X1 U313 ( .A(n900), .ZN(n628) );
  AOI22_X1 U314 ( .A1(data_in[7]), .A2(n821), .B1(n907), .B2(\mem[22][7] ), 
        .ZN(n900) );
  INV_X1 U315 ( .A(n899), .ZN(n627) );
  AOI22_X1 U316 ( .A1(data_in[0]), .A2(n820), .B1(n898), .B2(\mem[23][0] ), 
        .ZN(n899) );
  INV_X1 U317 ( .A(n897), .ZN(n626) );
  AOI22_X1 U318 ( .A1(data_in[1]), .A2(n820), .B1(n898), .B2(\mem[23][1] ), 
        .ZN(n897) );
  INV_X1 U319 ( .A(n896), .ZN(n625) );
  AOI22_X1 U320 ( .A1(data_in[2]), .A2(n820), .B1(n898), .B2(\mem[23][2] ), 
        .ZN(n896) );
  INV_X1 U321 ( .A(n895), .ZN(n624) );
  AOI22_X1 U322 ( .A1(data_in[3]), .A2(n820), .B1(n898), .B2(\mem[23][3] ), 
        .ZN(n895) );
  INV_X1 U323 ( .A(n894), .ZN(n623) );
  AOI22_X1 U324 ( .A1(data_in[4]), .A2(n820), .B1(n898), .B2(\mem[23][4] ), 
        .ZN(n894) );
  INV_X1 U325 ( .A(n893), .ZN(n622) );
  AOI22_X1 U326 ( .A1(data_in[5]), .A2(n820), .B1(n898), .B2(\mem[23][5] ), 
        .ZN(n893) );
  INV_X1 U327 ( .A(n892), .ZN(n621) );
  AOI22_X1 U328 ( .A1(data_in[6]), .A2(n820), .B1(n898), .B2(\mem[23][6] ), 
        .ZN(n892) );
  INV_X1 U329 ( .A(n891), .ZN(n620) );
  AOI22_X1 U330 ( .A1(data_in[7]), .A2(n820), .B1(n898), .B2(\mem[23][7] ), 
        .ZN(n891) );
  INV_X1 U331 ( .A(N12), .ZN(n255) );
  INV_X1 U332 ( .A(N11), .ZN(n254) );
  INV_X1 U333 ( .A(n999), .ZN(n715) );
  AOI22_X1 U334 ( .A1(data_in[0]), .A2(n831), .B1(n998), .B2(\mem[12][0] ), 
        .ZN(n999) );
  INV_X1 U335 ( .A(n997), .ZN(n714) );
  AOI22_X1 U336 ( .A1(data_in[1]), .A2(n831), .B1(n998), .B2(\mem[12][1] ), 
        .ZN(n997) );
  INV_X1 U337 ( .A(n996), .ZN(n713) );
  AOI22_X1 U338 ( .A1(data_in[2]), .A2(n831), .B1(n998), .B2(\mem[12][2] ), 
        .ZN(n996) );
  INV_X1 U339 ( .A(n995), .ZN(n712) );
  AOI22_X1 U340 ( .A1(data_in[3]), .A2(n831), .B1(n998), .B2(\mem[12][3] ), 
        .ZN(n995) );
  INV_X1 U341 ( .A(n994), .ZN(n711) );
  AOI22_X1 U342 ( .A1(data_in[4]), .A2(n831), .B1(n998), .B2(\mem[12][4] ), 
        .ZN(n994) );
  INV_X1 U343 ( .A(n993), .ZN(n710) );
  AOI22_X1 U344 ( .A1(data_in[5]), .A2(n831), .B1(n998), .B2(\mem[12][5] ), 
        .ZN(n993) );
  INV_X1 U345 ( .A(n992), .ZN(n709) );
  AOI22_X1 U346 ( .A1(data_in[6]), .A2(n831), .B1(n998), .B2(\mem[12][6] ), 
        .ZN(n992) );
  INV_X1 U347 ( .A(n991), .ZN(n708) );
  AOI22_X1 U348 ( .A1(data_in[7]), .A2(n831), .B1(n998), .B2(\mem[12][7] ), 
        .ZN(n991) );
  INV_X1 U349 ( .A(n926), .ZN(n651) );
  AOI22_X1 U350 ( .A1(data_in[0]), .A2(n823), .B1(n925), .B2(\mem[20][0] ), 
        .ZN(n926) );
  INV_X1 U351 ( .A(n924), .ZN(n650) );
  AOI22_X1 U352 ( .A1(data_in[1]), .A2(n823), .B1(n925), .B2(\mem[20][1] ), 
        .ZN(n924) );
  INV_X1 U353 ( .A(n923), .ZN(n649) );
  AOI22_X1 U354 ( .A1(data_in[2]), .A2(n823), .B1(n925), .B2(\mem[20][2] ), 
        .ZN(n923) );
  INV_X1 U355 ( .A(n922), .ZN(n648) );
  AOI22_X1 U356 ( .A1(data_in[3]), .A2(n823), .B1(n925), .B2(\mem[20][3] ), 
        .ZN(n922) );
  INV_X1 U357 ( .A(n921), .ZN(n647) );
  AOI22_X1 U358 ( .A1(data_in[4]), .A2(n823), .B1(n925), .B2(\mem[20][4] ), 
        .ZN(n921) );
  INV_X1 U359 ( .A(n920), .ZN(n646) );
  AOI22_X1 U360 ( .A1(data_in[5]), .A2(n823), .B1(n925), .B2(\mem[20][5] ), 
        .ZN(n920) );
  INV_X1 U361 ( .A(n919), .ZN(n645) );
  AOI22_X1 U362 ( .A1(data_in[6]), .A2(n823), .B1(n925), .B2(\mem[20][6] ), 
        .ZN(n919) );
  INV_X1 U363 ( .A(n918), .ZN(n644) );
  AOI22_X1 U364 ( .A1(data_in[7]), .A2(n823), .B1(n925), .B2(\mem[20][7] ), 
        .ZN(n918) );
  INV_X1 U365 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U366 ( .A1(data_in[0]), .A2(n835), .B1(n1035), .B2(\mem[8][0] ), 
        .ZN(n1036) );
  INV_X1 U367 ( .A(n1034), .ZN(n746) );
  AOI22_X1 U368 ( .A1(data_in[1]), .A2(n835), .B1(n1035), .B2(\mem[8][1] ), 
        .ZN(n1034) );
  INV_X1 U369 ( .A(n1033), .ZN(n745) );
  AOI22_X1 U370 ( .A1(data_in[2]), .A2(n835), .B1(n1035), .B2(\mem[8][2] ), 
        .ZN(n1033) );
  INV_X1 U371 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U372 ( .A1(data_in[3]), .A2(n835), .B1(n1035), .B2(\mem[8][3] ), 
        .ZN(n1032) );
  INV_X1 U373 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U374 ( .A1(data_in[4]), .A2(n835), .B1(n1035), .B2(\mem[8][4] ), 
        .ZN(n1031) );
  INV_X1 U375 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U376 ( .A1(data_in[5]), .A2(n835), .B1(n1035), .B2(\mem[8][5] ), 
        .ZN(n1030) );
  INV_X1 U377 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U378 ( .A1(data_in[6]), .A2(n835), .B1(n1035), .B2(\mem[8][6] ), 
        .ZN(n1029) );
  INV_X1 U379 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U380 ( .A1(data_in[7]), .A2(n835), .B1(n1035), .B2(\mem[8][7] ), 
        .ZN(n1028) );
  INV_X1 U381 ( .A(n963), .ZN(n683) );
  AOI22_X1 U382 ( .A1(data_in[0]), .A2(n827), .B1(n962), .B2(\mem[16][0] ), 
        .ZN(n963) );
  INV_X1 U383 ( .A(n961), .ZN(n682) );
  AOI22_X1 U384 ( .A1(data_in[1]), .A2(n827), .B1(n962), .B2(\mem[16][1] ), 
        .ZN(n961) );
  INV_X1 U385 ( .A(n960), .ZN(n681) );
  AOI22_X1 U386 ( .A1(data_in[2]), .A2(n827), .B1(n962), .B2(\mem[16][2] ), 
        .ZN(n960) );
  INV_X1 U387 ( .A(n959), .ZN(n680) );
  AOI22_X1 U388 ( .A1(data_in[3]), .A2(n827), .B1(n962), .B2(\mem[16][3] ), 
        .ZN(n959) );
  INV_X1 U389 ( .A(n958), .ZN(n679) );
  AOI22_X1 U390 ( .A1(data_in[4]), .A2(n827), .B1(n962), .B2(\mem[16][4] ), 
        .ZN(n958) );
  INV_X1 U391 ( .A(n957), .ZN(n678) );
  AOI22_X1 U392 ( .A1(data_in[5]), .A2(n827), .B1(n962), .B2(\mem[16][5] ), 
        .ZN(n957) );
  INV_X1 U393 ( .A(n956), .ZN(n677) );
  AOI22_X1 U394 ( .A1(data_in[6]), .A2(n827), .B1(n962), .B2(\mem[16][6] ), 
        .ZN(n956) );
  INV_X1 U395 ( .A(n955), .ZN(n676) );
  AOI22_X1 U396 ( .A1(data_in[7]), .A2(n827), .B1(n962), .B2(\mem[16][7] ), 
        .ZN(n955) );
  INV_X1 U397 ( .A(n890), .ZN(n619) );
  AOI22_X1 U398 ( .A1(data_in[0]), .A2(n816), .B1(n889), .B2(\mem[24][0] ), 
        .ZN(n890) );
  INV_X1 U399 ( .A(n888), .ZN(n618) );
  AOI22_X1 U400 ( .A1(data_in[1]), .A2(n816), .B1(n889), .B2(\mem[24][1] ), 
        .ZN(n888) );
  INV_X1 U401 ( .A(n887), .ZN(n617) );
  AOI22_X1 U402 ( .A1(data_in[2]), .A2(n816), .B1(n889), .B2(\mem[24][2] ), 
        .ZN(n887) );
  INV_X1 U403 ( .A(n886), .ZN(n616) );
  AOI22_X1 U404 ( .A1(data_in[3]), .A2(n816), .B1(n889), .B2(\mem[24][3] ), 
        .ZN(n886) );
  INV_X1 U405 ( .A(n885), .ZN(n615) );
  AOI22_X1 U406 ( .A1(data_in[4]), .A2(n816), .B1(n889), .B2(\mem[24][4] ), 
        .ZN(n885) );
  INV_X1 U407 ( .A(n884), .ZN(n614) );
  AOI22_X1 U408 ( .A1(data_in[5]), .A2(n816), .B1(n889), .B2(\mem[24][5] ), 
        .ZN(n884) );
  INV_X1 U409 ( .A(n883), .ZN(n613) );
  AOI22_X1 U410 ( .A1(data_in[6]), .A2(n816), .B1(n889), .B2(\mem[24][6] ), 
        .ZN(n883) );
  INV_X1 U411 ( .A(n882), .ZN(n612) );
  AOI22_X1 U412 ( .A1(data_in[7]), .A2(n816), .B1(n889), .B2(\mem[24][7] ), 
        .ZN(n882) );
  INV_X1 U413 ( .A(n881), .ZN(n611) );
  AOI22_X1 U414 ( .A1(data_in[0]), .A2(n815), .B1(n880), .B2(\mem[25][0] ), 
        .ZN(n881) );
  INV_X1 U415 ( .A(n879), .ZN(n610) );
  AOI22_X1 U416 ( .A1(data_in[1]), .A2(n815), .B1(n880), .B2(\mem[25][1] ), 
        .ZN(n879) );
  INV_X1 U417 ( .A(n878), .ZN(n609) );
  AOI22_X1 U418 ( .A1(data_in[2]), .A2(n815), .B1(n880), .B2(\mem[25][2] ), 
        .ZN(n878) );
  INV_X1 U419 ( .A(n877), .ZN(n608) );
  AOI22_X1 U420 ( .A1(data_in[3]), .A2(n815), .B1(n880), .B2(\mem[25][3] ), 
        .ZN(n877) );
  INV_X1 U421 ( .A(n876), .ZN(n607) );
  AOI22_X1 U422 ( .A1(data_in[4]), .A2(n815), .B1(n880), .B2(\mem[25][4] ), 
        .ZN(n876) );
  INV_X1 U423 ( .A(n875), .ZN(n606) );
  AOI22_X1 U424 ( .A1(data_in[5]), .A2(n815), .B1(n880), .B2(\mem[25][5] ), 
        .ZN(n875) );
  INV_X1 U425 ( .A(n874), .ZN(n605) );
  AOI22_X1 U426 ( .A1(data_in[6]), .A2(n815), .B1(n880), .B2(\mem[25][6] ), 
        .ZN(n874) );
  INV_X1 U427 ( .A(n873), .ZN(n604) );
  AOI22_X1 U428 ( .A1(data_in[7]), .A2(n815), .B1(n880), .B2(\mem[25][7] ), 
        .ZN(n873) );
  INV_X1 U429 ( .A(n872), .ZN(n603) );
  AOI22_X1 U430 ( .A1(data_in[0]), .A2(n814), .B1(n871), .B2(\mem[26][0] ), 
        .ZN(n872) );
  INV_X1 U431 ( .A(n870), .ZN(n602) );
  AOI22_X1 U432 ( .A1(data_in[1]), .A2(n814), .B1(n871), .B2(\mem[26][1] ), 
        .ZN(n870) );
  INV_X1 U433 ( .A(n869), .ZN(n601) );
  AOI22_X1 U434 ( .A1(data_in[2]), .A2(n814), .B1(n871), .B2(\mem[26][2] ), 
        .ZN(n869) );
  INV_X1 U435 ( .A(n868), .ZN(n600) );
  AOI22_X1 U436 ( .A1(data_in[3]), .A2(n814), .B1(n871), .B2(\mem[26][3] ), 
        .ZN(n868) );
  INV_X1 U437 ( .A(n867), .ZN(n599) );
  AOI22_X1 U438 ( .A1(data_in[4]), .A2(n814), .B1(n871), .B2(\mem[26][4] ), 
        .ZN(n867) );
  INV_X1 U439 ( .A(n866), .ZN(n598) );
  AOI22_X1 U440 ( .A1(data_in[5]), .A2(n814), .B1(n871), .B2(\mem[26][5] ), 
        .ZN(n866) );
  INV_X1 U441 ( .A(n865), .ZN(n597) );
  AOI22_X1 U442 ( .A1(data_in[6]), .A2(n814), .B1(n871), .B2(\mem[26][6] ), 
        .ZN(n865) );
  INV_X1 U443 ( .A(n864), .ZN(n596) );
  AOI22_X1 U444 ( .A1(data_in[7]), .A2(n814), .B1(n871), .B2(\mem[26][7] ), 
        .ZN(n864) );
  INV_X1 U445 ( .A(n863), .ZN(n595) );
  AOI22_X1 U446 ( .A1(data_in[0]), .A2(n813), .B1(n862), .B2(\mem[27][0] ), 
        .ZN(n863) );
  INV_X1 U447 ( .A(n861), .ZN(n594) );
  AOI22_X1 U448 ( .A1(data_in[1]), .A2(n813), .B1(n862), .B2(\mem[27][1] ), 
        .ZN(n861) );
  INV_X1 U449 ( .A(n860), .ZN(n293) );
  AOI22_X1 U450 ( .A1(data_in[2]), .A2(n813), .B1(n862), .B2(\mem[27][2] ), 
        .ZN(n860) );
  INV_X1 U451 ( .A(n859), .ZN(n292) );
  AOI22_X1 U452 ( .A1(data_in[3]), .A2(n813), .B1(n862), .B2(\mem[27][3] ), 
        .ZN(n859) );
  INV_X1 U453 ( .A(n858), .ZN(n291) );
  AOI22_X1 U454 ( .A1(data_in[4]), .A2(n813), .B1(n862), .B2(\mem[27][4] ), 
        .ZN(n858) );
  INV_X1 U455 ( .A(n857), .ZN(n290) );
  AOI22_X1 U456 ( .A1(data_in[5]), .A2(n813), .B1(n862), .B2(\mem[27][5] ), 
        .ZN(n857) );
  INV_X1 U457 ( .A(n856), .ZN(n289) );
  AOI22_X1 U458 ( .A1(data_in[6]), .A2(n813), .B1(n862), .B2(\mem[27][6] ), 
        .ZN(n856) );
  INV_X1 U459 ( .A(n855), .ZN(n288) );
  AOI22_X1 U460 ( .A1(data_in[7]), .A2(n813), .B1(n862), .B2(\mem[27][7] ), 
        .ZN(n855) );
  INV_X1 U461 ( .A(n854), .ZN(n287) );
  AOI22_X1 U462 ( .A1(data_in[0]), .A2(n812), .B1(n853), .B2(\mem[28][0] ), 
        .ZN(n854) );
  INV_X1 U463 ( .A(n852), .ZN(n286) );
  AOI22_X1 U464 ( .A1(data_in[1]), .A2(n812), .B1(n853), .B2(\mem[28][1] ), 
        .ZN(n852) );
  INV_X1 U465 ( .A(n851), .ZN(n285) );
  AOI22_X1 U466 ( .A1(data_in[2]), .A2(n812), .B1(n853), .B2(\mem[28][2] ), 
        .ZN(n851) );
  INV_X1 U467 ( .A(n850), .ZN(n284) );
  AOI22_X1 U468 ( .A1(data_in[3]), .A2(n812), .B1(n853), .B2(\mem[28][3] ), 
        .ZN(n850) );
  INV_X1 U469 ( .A(n849), .ZN(n283) );
  AOI22_X1 U470 ( .A1(data_in[4]), .A2(n812), .B1(n853), .B2(\mem[28][4] ), 
        .ZN(n849) );
  INV_X1 U471 ( .A(n848), .ZN(n282) );
  AOI22_X1 U472 ( .A1(data_in[5]), .A2(n812), .B1(n853), .B2(\mem[28][5] ), 
        .ZN(n848) );
  INV_X1 U473 ( .A(n847), .ZN(n281) );
  AOI22_X1 U474 ( .A1(data_in[6]), .A2(n812), .B1(n853), .B2(\mem[28][6] ), 
        .ZN(n847) );
  INV_X1 U475 ( .A(n846), .ZN(n280) );
  AOI22_X1 U476 ( .A1(data_in[7]), .A2(n812), .B1(n853), .B2(\mem[28][7] ), 
        .ZN(n846) );
  INV_X1 U477 ( .A(n1145), .ZN(n279) );
  AOI22_X1 U478 ( .A1(n819), .A2(data_in[0]), .B1(n1144), .B2(\mem[29][0] ), 
        .ZN(n1145) );
  INV_X1 U479 ( .A(n1143), .ZN(n278) );
  AOI22_X1 U480 ( .A1(n819), .A2(data_in[1]), .B1(n1144), .B2(\mem[29][1] ), 
        .ZN(n1143) );
  INV_X1 U481 ( .A(n1142), .ZN(n277) );
  AOI22_X1 U482 ( .A1(n819), .A2(data_in[2]), .B1(n1144), .B2(\mem[29][2] ), 
        .ZN(n1142) );
  INV_X1 U483 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U484 ( .A1(n819), .A2(data_in[3]), .B1(n1144), .B2(\mem[29][3] ), 
        .ZN(n1141) );
  INV_X1 U485 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U486 ( .A1(n819), .A2(data_in[4]), .B1(n1144), .B2(\mem[29][4] ), 
        .ZN(n1140) );
  INV_X1 U487 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U488 ( .A1(n819), .A2(data_in[5]), .B1(n1144), .B2(\mem[29][5] ), 
        .ZN(n1139) );
  INV_X1 U489 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U490 ( .A1(n819), .A2(data_in[6]), .B1(n1144), .B2(\mem[29][6] ), 
        .ZN(n1138) );
  INV_X1 U491 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U492 ( .A1(n819), .A2(data_in[7]), .B1(n1144), .B2(\mem[29][7] ), 
        .ZN(n1137) );
  INV_X1 U493 ( .A(n1134), .ZN(n271) );
  AOI22_X1 U494 ( .A1(data_in[0]), .A2(n818), .B1(n1133), .B2(\mem[30][0] ), 
        .ZN(n1134) );
  INV_X1 U495 ( .A(n1132), .ZN(n270) );
  AOI22_X1 U496 ( .A1(data_in[1]), .A2(n818), .B1(n1133), .B2(\mem[30][1] ), 
        .ZN(n1132) );
  INV_X1 U497 ( .A(n1131), .ZN(n269) );
  AOI22_X1 U498 ( .A1(data_in[2]), .A2(n818), .B1(n1133), .B2(\mem[30][2] ), 
        .ZN(n1131) );
  INV_X1 U499 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U500 ( .A1(data_in[3]), .A2(n818), .B1(n1133), .B2(\mem[30][3] ), 
        .ZN(n1130) );
  INV_X1 U501 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U502 ( .A1(data_in[4]), .A2(n818), .B1(n1133), .B2(\mem[30][4] ), 
        .ZN(n1129) );
  INV_X1 U503 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U504 ( .A1(data_in[5]), .A2(n818), .B1(n1133), .B2(\mem[30][5] ), 
        .ZN(n1128) );
  INV_X1 U505 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U506 ( .A1(data_in[6]), .A2(n818), .B1(n1133), .B2(\mem[30][6] ), 
        .ZN(n1127) );
  INV_X1 U507 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U508 ( .A1(data_in[7]), .A2(n818), .B1(n1133), .B2(\mem[30][7] ), 
        .ZN(n1126) );
  INV_X1 U509 ( .A(n1124), .ZN(n263) );
  AOI22_X1 U510 ( .A1(data_in[0]), .A2(n817), .B1(n1123), .B2(\mem[31][0] ), 
        .ZN(n1124) );
  INV_X1 U511 ( .A(n1122), .ZN(n262) );
  AOI22_X1 U512 ( .A1(data_in[1]), .A2(n817), .B1(n1123), .B2(\mem[31][1] ), 
        .ZN(n1122) );
  INV_X1 U513 ( .A(n1121), .ZN(n261) );
  AOI22_X1 U514 ( .A1(data_in[2]), .A2(n817), .B1(n1123), .B2(\mem[31][2] ), 
        .ZN(n1121) );
  INV_X1 U515 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U516 ( .A1(data_in[3]), .A2(n817), .B1(n1123), .B2(\mem[31][3] ), 
        .ZN(n1120) );
  INV_X1 U517 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U518 ( .A1(data_in[4]), .A2(n817), .B1(n1123), .B2(\mem[31][4] ), 
        .ZN(n1119) );
  INV_X1 U519 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U520 ( .A1(data_in[5]), .A2(n817), .B1(n1123), .B2(\mem[31][5] ), 
        .ZN(n1118) );
  INV_X1 U521 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U522 ( .A1(data_in[6]), .A2(n817), .B1(n1123), .B2(\mem[31][6] ), 
        .ZN(n1117) );
  INV_X1 U523 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U524 ( .A1(data_in[7]), .A2(n817), .B1(n1123), .B2(\mem[31][7] ), 
        .ZN(n1116) );
  INV_X1 U525 ( .A(n1114), .ZN(n811) );
  AOI22_X1 U526 ( .A1(data_in[0]), .A2(n843), .B1(n1113), .B2(\mem[0][0] ), 
        .ZN(n1114) );
  INV_X1 U527 ( .A(n1112), .ZN(n810) );
  AOI22_X1 U528 ( .A1(data_in[1]), .A2(n843), .B1(n1113), .B2(\mem[0][1] ), 
        .ZN(n1112) );
  INV_X1 U529 ( .A(n1111), .ZN(n809) );
  AOI22_X1 U530 ( .A1(data_in[2]), .A2(n843), .B1(n1113), .B2(\mem[0][2] ), 
        .ZN(n1111) );
  INV_X1 U531 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U532 ( .A1(data_in[3]), .A2(n843), .B1(n1113), .B2(\mem[0][3] ), 
        .ZN(n1110) );
  INV_X1 U533 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U534 ( .A1(data_in[4]), .A2(n843), .B1(n1113), .B2(\mem[0][4] ), 
        .ZN(n1109) );
  INV_X1 U535 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U536 ( .A1(data_in[5]), .A2(n843), .B1(n1113), .B2(\mem[0][5] ), 
        .ZN(n1108) );
  INV_X1 U537 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U538 ( .A1(data_in[6]), .A2(n843), .B1(n1113), .B2(\mem[0][6] ), 
        .ZN(n1107) );
  INV_X1 U539 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U540 ( .A1(data_in[7]), .A2(n843), .B1(n1113), .B2(\mem[0][7] ), 
        .ZN(n1106) );
  INV_X1 U541 ( .A(n1103), .ZN(n803) );
  AOI22_X1 U542 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[1][0] ), 
        .ZN(n1103) );
  INV_X1 U543 ( .A(n1101), .ZN(n802) );
  AOI22_X1 U544 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[1][1] ), 
        .ZN(n1101) );
  INV_X1 U545 ( .A(n1100), .ZN(n801) );
  AOI22_X1 U546 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[1][2] ), 
        .ZN(n1100) );
  INV_X1 U547 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U548 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[1][3] ), 
        .ZN(n1099) );
  INV_X1 U549 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U550 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[1][4] ), 
        .ZN(n1098) );
  INV_X1 U551 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U552 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[1][5] ), 
        .ZN(n1097) );
  INV_X1 U553 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U554 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[1][6] ), 
        .ZN(n1096) );
  INV_X1 U555 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U556 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[1][7] ), 
        .ZN(n1095) );
  INV_X1 U557 ( .A(n1093), .ZN(n795) );
  AOI22_X1 U558 ( .A1(data_in[0]), .A2(n841), .B1(n1092), .B2(\mem[2][0] ), 
        .ZN(n1093) );
  INV_X1 U559 ( .A(n1091), .ZN(n794) );
  AOI22_X1 U560 ( .A1(data_in[1]), .A2(n841), .B1(n1092), .B2(\mem[2][1] ), 
        .ZN(n1091) );
  INV_X1 U561 ( .A(n1090), .ZN(n793) );
  AOI22_X1 U562 ( .A1(data_in[2]), .A2(n841), .B1(n1092), .B2(\mem[2][2] ), 
        .ZN(n1090) );
  INV_X1 U563 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U564 ( .A1(data_in[3]), .A2(n841), .B1(n1092), .B2(\mem[2][3] ), 
        .ZN(n1089) );
  INV_X1 U565 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U566 ( .A1(data_in[4]), .A2(n841), .B1(n1092), .B2(\mem[2][4] ), 
        .ZN(n1088) );
  INV_X1 U567 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U568 ( .A1(data_in[5]), .A2(n841), .B1(n1092), .B2(\mem[2][5] ), 
        .ZN(n1087) );
  INV_X1 U569 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U570 ( .A1(data_in[6]), .A2(n841), .B1(n1092), .B2(\mem[2][6] ), 
        .ZN(n1086) );
  INV_X1 U571 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U572 ( .A1(data_in[7]), .A2(n841), .B1(n1092), .B2(\mem[2][7] ), 
        .ZN(n1085) );
  INV_X1 U573 ( .A(n1083), .ZN(n787) );
  AOI22_X1 U574 ( .A1(data_in[0]), .A2(n840), .B1(n1082), .B2(\mem[3][0] ), 
        .ZN(n1083) );
  INV_X1 U575 ( .A(n1081), .ZN(n786) );
  AOI22_X1 U576 ( .A1(data_in[1]), .A2(n840), .B1(n1082), .B2(\mem[3][1] ), 
        .ZN(n1081) );
  INV_X1 U577 ( .A(n1080), .ZN(n785) );
  AOI22_X1 U578 ( .A1(data_in[2]), .A2(n840), .B1(n1082), .B2(\mem[3][2] ), 
        .ZN(n1080) );
  INV_X1 U579 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U580 ( .A1(data_in[3]), .A2(n840), .B1(n1082), .B2(\mem[3][3] ), 
        .ZN(n1079) );
  INV_X1 U581 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U582 ( .A1(data_in[4]), .A2(n840), .B1(n1082), .B2(\mem[3][4] ), 
        .ZN(n1078) );
  INV_X1 U583 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U584 ( .A1(data_in[5]), .A2(n840), .B1(n1082), .B2(\mem[3][5] ), 
        .ZN(n1077) );
  INV_X1 U585 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U586 ( .A1(data_in[6]), .A2(n840), .B1(n1082), .B2(\mem[3][6] ), 
        .ZN(n1076) );
  INV_X1 U587 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U588 ( .A1(data_in[7]), .A2(n840), .B1(n1082), .B2(\mem[3][7] ), 
        .ZN(n1075) );
  INV_X1 U589 ( .A(n1073), .ZN(n779) );
  AOI22_X1 U590 ( .A1(data_in[0]), .A2(n839), .B1(n1072), .B2(\mem[4][0] ), 
        .ZN(n1073) );
  INV_X1 U591 ( .A(n1071), .ZN(n778) );
  AOI22_X1 U592 ( .A1(data_in[1]), .A2(n839), .B1(n1072), .B2(\mem[4][1] ), 
        .ZN(n1071) );
  INV_X1 U593 ( .A(n1070), .ZN(n777) );
  AOI22_X1 U594 ( .A1(data_in[2]), .A2(n839), .B1(n1072), .B2(\mem[4][2] ), 
        .ZN(n1070) );
  INV_X1 U595 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U596 ( .A1(data_in[3]), .A2(n839), .B1(n1072), .B2(\mem[4][3] ), 
        .ZN(n1069) );
  INV_X1 U597 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U598 ( .A1(data_in[4]), .A2(n839), .B1(n1072), .B2(\mem[4][4] ), 
        .ZN(n1068) );
  INV_X1 U599 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U600 ( .A1(data_in[5]), .A2(n839), .B1(n1072), .B2(\mem[4][5] ), 
        .ZN(n1067) );
  INV_X1 U601 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U602 ( .A1(data_in[6]), .A2(n839), .B1(n1072), .B2(\mem[4][6] ), 
        .ZN(n1066) );
  INV_X1 U603 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U604 ( .A1(data_in[7]), .A2(n839), .B1(n1072), .B2(\mem[4][7] ), 
        .ZN(n1065) );
  INV_X1 U605 ( .A(N13), .ZN(n844) );
  INV_X1 U606 ( .A(N14), .ZN(n845) );
  MUX2_X1 U607 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n251), .Z(n3) );
  MUX2_X1 U608 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n247), .Z(n4) );
  MUX2_X1 U609 ( .A(n4), .B(n3), .S(n245), .Z(n5) );
  MUX2_X1 U610 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n251), .Z(n6) );
  MUX2_X1 U611 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n251), .Z(n7) );
  MUX2_X1 U612 ( .A(n7), .B(n6), .S(n245), .Z(n8) );
  MUX2_X1 U613 ( .A(n8), .B(n5), .S(n243), .Z(n9) );
  MUX2_X1 U614 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n252), .Z(n10) );
  MUX2_X1 U615 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n250), .Z(n11) );
  MUX2_X1 U616 ( .A(n11), .B(n10), .S(N11), .Z(n12) );
  MUX2_X1 U617 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n249), .Z(n13) );
  MUX2_X1 U618 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n249), .Z(n14) );
  MUX2_X1 U619 ( .A(n14), .B(n13), .S(N11), .Z(n15) );
  MUX2_X1 U620 ( .A(n15), .B(n12), .S(n243), .Z(n16) );
  MUX2_X1 U621 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U622 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n247), .Z(n18) );
  MUX2_X1 U623 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n247), .Z(n19) );
  MUX2_X1 U624 ( .A(n19), .B(n18), .S(n246), .Z(n20) );
  MUX2_X1 U625 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n247), .Z(n21) );
  MUX2_X1 U626 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n247), .Z(n22) );
  MUX2_X1 U627 ( .A(n22), .B(n21), .S(n244), .Z(n23) );
  MUX2_X1 U628 ( .A(n23), .B(n20), .S(n243), .Z(n24) );
  MUX2_X1 U629 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n247), .Z(n25) );
  MUX2_X1 U630 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n247), .Z(n26) );
  MUX2_X1 U631 ( .A(n26), .B(n25), .S(N11), .Z(n27) );
  MUX2_X1 U632 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n247), .Z(n28) );
  MUX2_X1 U633 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n247), .Z(n29) );
  MUX2_X1 U634 ( .A(n29), .B(n28), .S(n246), .Z(n30) );
  MUX2_X1 U635 ( .A(n30), .B(n27), .S(n243), .Z(n31) );
  MUX2_X1 U636 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U637 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U638 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n247), .Z(n33) );
  MUX2_X1 U639 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n247), .Z(n34) );
  MUX2_X1 U640 ( .A(n34), .B(n33), .S(n244), .Z(n35) );
  MUX2_X1 U641 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n247), .Z(n36) );
  MUX2_X1 U642 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n247), .Z(n37) );
  MUX2_X1 U643 ( .A(n37), .B(n36), .S(n244), .Z(n38) );
  MUX2_X1 U644 ( .A(n38), .B(n35), .S(n243), .Z(n39) );
  MUX2_X1 U645 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n248), .Z(n40) );
  MUX2_X1 U646 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n248), .Z(n41) );
  MUX2_X1 U647 ( .A(n41), .B(n40), .S(n246), .Z(n42) );
  MUX2_X1 U648 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n248), .Z(n43) );
  MUX2_X1 U649 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n248), .Z(n44) );
  MUX2_X1 U650 ( .A(n44), .B(n43), .S(n246), .Z(n45) );
  MUX2_X1 U651 ( .A(n45), .B(n42), .S(N12), .Z(n46) );
  MUX2_X1 U652 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U653 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n248), .Z(n48) );
  MUX2_X1 U654 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n248), .Z(n49) );
  MUX2_X1 U655 ( .A(n49), .B(n48), .S(N11), .Z(n50) );
  MUX2_X1 U656 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n248), .Z(n51) );
  MUX2_X1 U657 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n248), .Z(n52) );
  MUX2_X1 U658 ( .A(n52), .B(n51), .S(n245), .Z(n53) );
  MUX2_X1 U659 ( .A(n53), .B(n50), .S(N12), .Z(n54) );
  MUX2_X1 U660 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n248), .Z(n55) );
  MUX2_X1 U661 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n248), .Z(n56) );
  MUX2_X1 U662 ( .A(n56), .B(n55), .S(N11), .Z(n57) );
  MUX2_X1 U663 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n248), .Z(n58) );
  MUX2_X1 U664 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n248), .Z(n59) );
  MUX2_X1 U665 ( .A(n59), .B(n58), .S(N11), .Z(n60) );
  MUX2_X1 U666 ( .A(n60), .B(n57), .S(N12), .Z(n61) );
  MUX2_X1 U667 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U668 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U669 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n249), .Z(n63) );
  MUX2_X1 U670 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n249), .Z(n64) );
  MUX2_X1 U671 ( .A(n64), .B(n63), .S(n244), .Z(n65) );
  MUX2_X1 U672 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n249), .Z(n66) );
  MUX2_X1 U673 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n249), .Z(n67) );
  MUX2_X1 U674 ( .A(n67), .B(n66), .S(n244), .Z(n68) );
  MUX2_X1 U675 ( .A(n68), .B(n65), .S(n243), .Z(n69) );
  MUX2_X1 U676 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n249), .Z(n70) );
  MUX2_X1 U677 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n249), .Z(n71) );
  MUX2_X1 U678 ( .A(n71), .B(n70), .S(n244), .Z(n72) );
  MUX2_X1 U679 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n249), .Z(n73) );
  MUX2_X1 U680 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n249), .Z(n74) );
  MUX2_X1 U681 ( .A(n74), .B(n73), .S(n244), .Z(n75) );
  MUX2_X1 U682 ( .A(n75), .B(n72), .S(n243), .Z(n76) );
  MUX2_X1 U683 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U684 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n249), .Z(n78) );
  MUX2_X1 U685 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n249), .Z(n79) );
  MUX2_X1 U686 ( .A(n79), .B(n78), .S(n244), .Z(n80) );
  MUX2_X1 U687 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n249), .Z(n81) );
  MUX2_X1 U688 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n249), .Z(n82) );
  MUX2_X1 U689 ( .A(n82), .B(n81), .S(n244), .Z(n83) );
  MUX2_X1 U690 ( .A(n83), .B(n80), .S(n243), .Z(n84) );
  MUX2_X1 U691 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n250), .Z(n85) );
  MUX2_X1 U692 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n250), .Z(n86) );
  MUX2_X1 U693 ( .A(n86), .B(n85), .S(n244), .Z(n87) );
  MUX2_X1 U694 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n250), .Z(n88) );
  MUX2_X1 U695 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n250), .Z(n89) );
  MUX2_X1 U696 ( .A(n89), .B(n88), .S(n244), .Z(n90) );
  MUX2_X1 U697 ( .A(n90), .B(n87), .S(n243), .Z(n91) );
  MUX2_X1 U698 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U699 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U700 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n250), .Z(n93) );
  MUX2_X1 U701 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U702 ( .A(n94), .B(n93), .S(n244), .Z(n95) );
  MUX2_X1 U703 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n250), .Z(n96) );
  MUX2_X1 U704 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n250), .Z(n97) );
  MUX2_X1 U705 ( .A(n97), .B(n96), .S(n244), .Z(n98) );
  MUX2_X1 U706 ( .A(n98), .B(n95), .S(n243), .Z(n99) );
  MUX2_X1 U707 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n100) );
  MUX2_X1 U708 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n250), .Z(n101) );
  MUX2_X1 U709 ( .A(n101), .B(n100), .S(n244), .Z(n102) );
  MUX2_X1 U710 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n250), .Z(n103) );
  MUX2_X1 U711 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n250), .Z(n104) );
  MUX2_X1 U712 ( .A(n104), .B(n103), .S(n244), .Z(n105) );
  MUX2_X1 U713 ( .A(n105), .B(n102), .S(n243), .Z(n106) );
  MUX2_X1 U714 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U715 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n252), .Z(n108) );
  MUX2_X1 U716 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(N10), .Z(n109) );
  MUX2_X1 U717 ( .A(n109), .B(n108), .S(n245), .Z(n110) );
  MUX2_X1 U718 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(N10), .Z(n111) );
  MUX2_X1 U719 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n248), .Z(n112) );
  MUX2_X1 U720 ( .A(n112), .B(n111), .S(n245), .Z(n113) );
  MUX2_X1 U721 ( .A(n113), .B(n110), .S(n243), .Z(n114) );
  MUX2_X1 U722 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(N10), .Z(n115) );
  MUX2_X1 U723 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n252), .Z(n116) );
  MUX2_X1 U724 ( .A(n116), .B(n115), .S(n245), .Z(n117) );
  MUX2_X1 U725 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n118) );
  MUX2_X1 U726 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n248), .Z(n119) );
  MUX2_X1 U727 ( .A(n119), .B(n118), .S(n245), .Z(n120) );
  MUX2_X1 U728 ( .A(n120), .B(n117), .S(n243), .Z(n121) );
  MUX2_X1 U729 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U730 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U731 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n248), .Z(n123) );
  MUX2_X1 U732 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(N10), .Z(n124) );
  MUX2_X1 U733 ( .A(n124), .B(n123), .S(n245), .Z(n125) );
  MUX2_X1 U734 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(N10), .Z(n126) );
  MUX2_X1 U735 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n127) );
  MUX2_X1 U736 ( .A(n127), .B(n126), .S(n245), .Z(n128) );
  MUX2_X1 U737 ( .A(n128), .B(n125), .S(n243), .Z(n129) );
  MUX2_X1 U738 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n251), .Z(n130) );
  MUX2_X1 U739 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(N10), .Z(n131) );
  MUX2_X1 U740 ( .A(n131), .B(n130), .S(n245), .Z(n132) );
  MUX2_X1 U741 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n252), .Z(n133) );
  MUX2_X1 U742 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(N10), .Z(n134) );
  MUX2_X1 U743 ( .A(n134), .B(n133), .S(n245), .Z(n135) );
  MUX2_X1 U744 ( .A(n135), .B(n132), .S(n243), .Z(n136) );
  MUX2_X1 U745 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U746 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n251), .Z(n138) );
  MUX2_X1 U747 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n252), .Z(n139) );
  MUX2_X1 U748 ( .A(n139), .B(n138), .S(n245), .Z(n140) );
  MUX2_X1 U749 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n248), .Z(n141) );
  MUX2_X1 U750 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(N10), .Z(n142) );
  MUX2_X1 U751 ( .A(n142), .B(n141), .S(n245), .Z(n143) );
  MUX2_X1 U752 ( .A(n143), .B(n140), .S(n243), .Z(n144) );
  MUX2_X1 U753 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(N10), .Z(n145) );
  MUX2_X1 U754 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(N10), .Z(n146) );
  MUX2_X1 U755 ( .A(n146), .B(n145), .S(n245), .Z(n147) );
  MUX2_X1 U756 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(N10), .Z(n148) );
  MUX2_X1 U757 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n149) );
  MUX2_X1 U758 ( .A(n149), .B(n148), .S(n245), .Z(n150) );
  MUX2_X1 U759 ( .A(n150), .B(n147), .S(n243), .Z(n151) );
  MUX2_X1 U760 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U761 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U762 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n251), .Z(n153) );
  MUX2_X1 U763 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n251), .Z(n154) );
  MUX2_X1 U764 ( .A(n154), .B(n153), .S(n246), .Z(n155) );
  MUX2_X1 U765 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n251), .Z(n156) );
  MUX2_X1 U766 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n251), .Z(n157) );
  MUX2_X1 U767 ( .A(n157), .B(n156), .S(n246), .Z(n158) );
  MUX2_X1 U768 ( .A(n158), .B(n155), .S(n243), .Z(n159) );
  MUX2_X1 U769 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n251), .Z(n160) );
  MUX2_X1 U770 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n251), .Z(n161) );
  MUX2_X1 U771 ( .A(n161), .B(n160), .S(n246), .Z(n162) );
  MUX2_X1 U772 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n251), .Z(n163) );
  MUX2_X1 U773 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n251), .Z(n164) );
  MUX2_X1 U774 ( .A(n164), .B(n163), .S(n246), .Z(n165) );
  MUX2_X1 U775 ( .A(n165), .B(n162), .S(N12), .Z(n166) );
  MUX2_X1 U776 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U777 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n251), .Z(n168) );
  MUX2_X1 U778 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n251), .Z(n169) );
  MUX2_X1 U779 ( .A(n169), .B(n168), .S(n246), .Z(n170) );
  MUX2_X1 U780 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n251), .Z(n171) );
  MUX2_X1 U781 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n251), .Z(n172) );
  MUX2_X1 U782 ( .A(n172), .B(n171), .S(n246), .Z(n173) );
  MUX2_X1 U783 ( .A(n173), .B(n170), .S(n243), .Z(n174) );
  MUX2_X1 U784 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n252), .Z(n175) );
  MUX2_X1 U785 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n247), .Z(n176) );
  MUX2_X1 U786 ( .A(n176), .B(n175), .S(n246), .Z(n177) );
  MUX2_X1 U787 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n252), .Z(n178) );
  MUX2_X1 U788 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n247), .Z(n179) );
  MUX2_X1 U789 ( .A(n179), .B(n178), .S(n246), .Z(n180) );
  MUX2_X1 U790 ( .A(n180), .B(n177), .S(N12), .Z(n181) );
  MUX2_X1 U791 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U792 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U793 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n247), .Z(n183) );
  MUX2_X1 U794 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n250), .Z(n184) );
  MUX2_X1 U795 ( .A(n184), .B(n183), .S(n246), .Z(n185) );
  MUX2_X1 U796 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n251), .Z(n186) );
  MUX2_X1 U797 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n252), .Z(n187) );
  MUX2_X1 U798 ( .A(n187), .B(n186), .S(n246), .Z(n188) );
  MUX2_X1 U799 ( .A(n188), .B(n185), .S(n243), .Z(n189) );
  MUX2_X1 U800 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n252), .Z(n190) );
  MUX2_X1 U801 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n252), .Z(n191) );
  MUX2_X1 U802 ( .A(n191), .B(n190), .S(n246), .Z(n192) );
  MUX2_X1 U803 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n249), .Z(n193) );
  MUX2_X1 U804 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n252), .Z(n194) );
  MUX2_X1 U805 ( .A(n194), .B(n193), .S(n246), .Z(n195) );
  MUX2_X1 U806 ( .A(n195), .B(n192), .S(N12), .Z(n196) );
  MUX2_X1 U807 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U808 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n250), .Z(n198) );
  MUX2_X1 U809 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n252), .Z(n199) );
  MUX2_X1 U810 ( .A(n199), .B(n198), .S(N11), .Z(n200) );
  MUX2_X1 U811 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n248), .Z(n201) );
  MUX2_X1 U812 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n249), .Z(n202) );
  MUX2_X1 U813 ( .A(n202), .B(n201), .S(n246), .Z(n203) );
  MUX2_X1 U814 ( .A(n203), .B(n200), .S(n243), .Z(n204) );
  MUX2_X1 U815 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n250), .Z(n205) );
  MUX2_X1 U816 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n252), .Z(n206) );
  MUX2_X1 U817 ( .A(n206), .B(n205), .S(N11), .Z(n207) );
  MUX2_X1 U818 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n252), .Z(n208) );
  MUX2_X1 U819 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n249), .Z(n209) );
  MUX2_X1 U820 ( .A(n209), .B(n208), .S(n244), .Z(n210) );
  MUX2_X1 U821 ( .A(n210), .B(n207), .S(N12), .Z(n211) );
  MUX2_X1 U822 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U823 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U824 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n249), .Z(n213) );
  MUX2_X1 U825 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n249), .Z(n214) );
  MUX2_X1 U826 ( .A(n214), .B(n213), .S(N11), .Z(n215) );
  MUX2_X1 U827 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n247), .Z(n216) );
  MUX2_X1 U828 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n250), .Z(n217) );
  MUX2_X1 U829 ( .A(n217), .B(n216), .S(N11), .Z(n218) );
  MUX2_X1 U830 ( .A(n218), .B(n215), .S(n243), .Z(n219) );
  MUX2_X1 U831 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n252), .Z(n220) );
  MUX2_X1 U832 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n250), .Z(n221) );
  MUX2_X1 U833 ( .A(n221), .B(n220), .S(N11), .Z(n222) );
  MUX2_X1 U834 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n252), .Z(n223) );
  MUX2_X1 U835 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n250), .Z(n224) );
  MUX2_X1 U836 ( .A(n224), .B(n223), .S(n245), .Z(n225) );
  MUX2_X1 U837 ( .A(n225), .B(n222), .S(N12), .Z(n226) );
  MUX2_X1 U838 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U839 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(N10), .Z(n228) );
  MUX2_X1 U840 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n248), .Z(n229) );
  MUX2_X1 U841 ( .A(n229), .B(n228), .S(N11), .Z(n230) );
  MUX2_X1 U842 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n252), .Z(n231) );
  MUX2_X1 U843 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n248), .Z(n232) );
  MUX2_X1 U844 ( .A(n232), .B(n231), .S(n244), .Z(n233) );
  MUX2_X1 U845 ( .A(n233), .B(n230), .S(n243), .Z(n234) );
  MUX2_X1 U846 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n247), .Z(n235) );
  MUX2_X1 U847 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n252), .Z(n236) );
  MUX2_X1 U848 ( .A(n236), .B(n235), .S(N11), .Z(n237) );
  MUX2_X1 U849 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n252), .Z(n238) );
  MUX2_X1 U850 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n252), .Z(n239) );
  MUX2_X1 U851 ( .A(n239), .B(n238), .S(n245), .Z(n240) );
  MUX2_X1 U852 ( .A(n240), .B(n237), .S(N12), .Z(n241) );
  MUX2_X1 U853 ( .A(n241), .B(n234), .S(N13), .Z(n242) );
  MUX2_X1 U854 ( .A(n242), .B(n227), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_30 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n256), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n257), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n258), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n259), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n260), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n261), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n262), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n263), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n264), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n265), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n266), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n267), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n268), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n269), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n270), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n271), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n272), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n273), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n274), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n275), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n276), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n277), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n278), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n279), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n280), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n281), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n282), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n283), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n284), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n285), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n286), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n287), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n288), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n289), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n290), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n291), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n292), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n293), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n594), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n595), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n596), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n597), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n598), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n599), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n600), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n601), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n602), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n603), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n604), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n605), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n606), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n607), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n608), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n609), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n610), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n611), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n612), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n613), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n614), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n615), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n616), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n617), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n618), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n619), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n620), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n621), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n622), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n623), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n624), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n625), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n626), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n627), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n628), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n629), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n630), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n631), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n632), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n633), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n634), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n635), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n636), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n637), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n638), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n639), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n640), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n641), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n642), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n643), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n644), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n645), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n646), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n647), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n648), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n649), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n650), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n651), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n652), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n653), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n654), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n655), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n656), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n657), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n658), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n659), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n660), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n661), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n662), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n663), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n664), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n665), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n666), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n667), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n668), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n669), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n670), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n671), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n672), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n673), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n674), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n675), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n676), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n677), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n678), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n679), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n680), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n681), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n682), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n683), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n684), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n685), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n686), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n687), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n688), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n689), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n690), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n691), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n692), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n693), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n694), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n695), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n696), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n697), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n698), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n699), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n700), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n701), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n702), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n703), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n704), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n705), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n706), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n707), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n708), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n709), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n710), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n711), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n712), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n713), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n714), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n715), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n716), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n717), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n718), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n719), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n720), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n721), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n722), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n723), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n724), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n725), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n726), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n727), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n728), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n729), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n730), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n731), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n732), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n733), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n734), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n735), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n736), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n737), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n738), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n739), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n740), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n741), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n742), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n743), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n744), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n745), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n746), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n747), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n748), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n749), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n750), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n751), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n752), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n753), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n754), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n755), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n756), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n757), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n758), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n759), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n760), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n761), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n762), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n763), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n764), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n765), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n766), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n767), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n768), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n769), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n770), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n771), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n772), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n773), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n774), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n775), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n776), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n777), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n778), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n779), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n780), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n781), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n782), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n783), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n784), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n785), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n786), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n787), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n788), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n789), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n790), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n791), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n792), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n793), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n794), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n795), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n796), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n797), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n798), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n799), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n800), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n801), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n802), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n803), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n804), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n805), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n806), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n807), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n808), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n809), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n810), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n811), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(n252), .Z(n249) );
  BUF_X1 U5 ( .A(n252), .Z(n250) );
  BUF_X1 U6 ( .A(N10), .Z(n251) );
  BUF_X1 U7 ( .A(n252), .Z(n248) );
  BUF_X1 U8 ( .A(n252), .Z(n247) );
  BUF_X1 U9 ( .A(N10), .Z(n252) );
  INV_X1 U10 ( .A(n1113), .ZN(n843) );
  INV_X1 U11 ( .A(n1102), .ZN(n842) );
  INV_X1 U12 ( .A(n1092), .ZN(n841) );
  INV_X1 U13 ( .A(n1082), .ZN(n840) );
  INV_X1 U14 ( .A(n1072), .ZN(n839) );
  INV_X1 U15 ( .A(n1062), .ZN(n838) );
  INV_X1 U16 ( .A(n1053), .ZN(n837) );
  INV_X1 U17 ( .A(n1044), .ZN(n836) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1105) );
  NOR3_X1 U19 ( .A1(N11), .A2(N12), .A3(n253), .ZN(n1094) );
  NAND2_X1 U20 ( .A1(n1104), .A2(n1136), .ZN(n1062) );
  NAND2_X1 U21 ( .A1(n1105), .A2(n1104), .ZN(n1113) );
  NAND2_X1 U22 ( .A1(n1094), .A2(n1104), .ZN(n1102) );
  NAND2_X1 U23 ( .A1(n1084), .A2(n1104), .ZN(n1092) );
  NAND2_X1 U24 ( .A1(n1074), .A2(n1104), .ZN(n1082) );
  NAND2_X1 U25 ( .A1(n1064), .A2(n1104), .ZN(n1072) );
  NAND2_X1 U26 ( .A1(n1104), .A2(n1125), .ZN(n1053) );
  NAND2_X1 U27 ( .A1(n1104), .A2(n1115), .ZN(n1044) );
  INV_X1 U28 ( .A(n1133), .ZN(n818) );
  INV_X1 U29 ( .A(n1123), .ZN(n817) );
  INV_X1 U30 ( .A(n889), .ZN(n816) );
  INV_X1 U31 ( .A(n880), .ZN(n815) );
  INV_X1 U32 ( .A(n871), .ZN(n814) );
  INV_X1 U33 ( .A(n862), .ZN(n813) );
  INV_X1 U34 ( .A(n853), .ZN(n812) );
  INV_X1 U35 ( .A(n989), .ZN(n830) );
  INV_X1 U36 ( .A(n980), .ZN(n829) );
  INV_X1 U37 ( .A(n971), .ZN(n828) );
  INV_X1 U38 ( .A(n916), .ZN(n822) );
  INV_X1 U39 ( .A(n907), .ZN(n821) );
  INV_X1 U40 ( .A(n898), .ZN(n820) );
  INV_X1 U41 ( .A(n1035), .ZN(n835) );
  INV_X1 U42 ( .A(n1025), .ZN(n834) );
  INV_X1 U43 ( .A(n1016), .ZN(n833) );
  INV_X1 U44 ( .A(n1007), .ZN(n832) );
  INV_X1 U45 ( .A(n998), .ZN(n831) );
  INV_X1 U46 ( .A(n962), .ZN(n827) );
  INV_X1 U47 ( .A(n952), .ZN(n826) );
  INV_X1 U48 ( .A(n943), .ZN(n825) );
  INV_X1 U49 ( .A(n934), .ZN(n824) );
  INV_X1 U50 ( .A(n925), .ZN(n823) );
  INV_X1 U51 ( .A(n1144), .ZN(n819) );
  BUF_X1 U52 ( .A(N11), .Z(n244) );
  BUF_X1 U53 ( .A(N11), .Z(n245) );
  BUF_X1 U54 ( .A(N11), .Z(n246) );
  INV_X1 U55 ( .A(N10), .ZN(n253) );
  BUF_X1 U56 ( .A(N12), .Z(n243) );
  NOR3_X1 U57 ( .A1(n255), .A2(N10), .A3(n254), .ZN(n1125) );
  NOR3_X1 U58 ( .A1(n255), .A2(n253), .A3(n254), .ZN(n1115) );
  NOR3_X1 U59 ( .A1(n253), .A2(N11), .A3(n255), .ZN(n1136) );
  NOR3_X1 U60 ( .A1(N10), .A2(N12), .A3(n254), .ZN(n1084) );
  NOR3_X1 U61 ( .A1(n253), .A2(N12), .A3(n254), .ZN(n1074) );
  NOR3_X1 U62 ( .A1(N10), .A2(N11), .A3(n255), .ZN(n1064) );
  NAND2_X1 U63 ( .A1(n1027), .A2(n1136), .ZN(n989) );
  NAND2_X1 U64 ( .A1(n954), .A2(n1136), .ZN(n916) );
  NAND2_X1 U65 ( .A1(n1027), .A2(n1064), .ZN(n998) );
  NAND2_X1 U66 ( .A1(n954), .A2(n1064), .ZN(n925) );
  NAND2_X1 U67 ( .A1(n1027), .A2(n1105), .ZN(n1035) );
  NAND2_X1 U68 ( .A1(n1027), .A2(n1094), .ZN(n1025) );
  NAND2_X1 U69 ( .A1(n954), .A2(n1105), .ZN(n962) );
  NAND2_X1 U70 ( .A1(n954), .A2(n1094), .ZN(n952) );
  NAND2_X1 U71 ( .A1(n1105), .A2(n1135), .ZN(n889) );
  NAND2_X1 U72 ( .A1(n1094), .A2(n1135), .ZN(n880) );
  NAND2_X1 U73 ( .A1(n1084), .A2(n1135), .ZN(n871) );
  NAND2_X1 U74 ( .A1(n1074), .A2(n1135), .ZN(n862) );
  NAND2_X1 U75 ( .A1(n1064), .A2(n1135), .ZN(n853) );
  NAND2_X1 U76 ( .A1(n1136), .A2(n1135), .ZN(n1144) );
  NAND2_X1 U77 ( .A1(n1125), .A2(n1135), .ZN(n1133) );
  NAND2_X1 U78 ( .A1(n1115), .A2(n1135), .ZN(n1123) );
  NAND2_X1 U79 ( .A1(n1027), .A2(n1084), .ZN(n1016) );
  NAND2_X1 U80 ( .A1(n1027), .A2(n1074), .ZN(n1007) );
  NAND2_X1 U81 ( .A1(n954), .A2(n1084), .ZN(n943) );
  NAND2_X1 U82 ( .A1(n954), .A2(n1074), .ZN(n934) );
  NAND2_X1 U83 ( .A1(n1027), .A2(n1125), .ZN(n980) );
  NAND2_X1 U84 ( .A1(n954), .A2(n1125), .ZN(n907) );
  NAND2_X1 U85 ( .A1(n1027), .A2(n1115), .ZN(n971) );
  NAND2_X1 U86 ( .A1(n954), .A2(n1115), .ZN(n898) );
  AND3_X1 U87 ( .A1(n844), .A2(n845), .A3(wr_en), .ZN(n1104) );
  AND3_X1 U88 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1135) );
  AND3_X1 U89 ( .A1(N13), .A2(n845), .A3(wr_en), .ZN(n1027) );
  AND3_X1 U90 ( .A1(N14), .A2(n844), .A3(wr_en), .ZN(n954) );
  INV_X1 U91 ( .A(n1063), .ZN(n771) );
  AOI22_X1 U92 ( .A1(data_in[0]), .A2(n838), .B1(n1062), .B2(\mem[5][0] ), 
        .ZN(n1063) );
  INV_X1 U93 ( .A(n1061), .ZN(n770) );
  AOI22_X1 U94 ( .A1(data_in[1]), .A2(n838), .B1(n1062), .B2(\mem[5][1] ), 
        .ZN(n1061) );
  INV_X1 U95 ( .A(n1060), .ZN(n769) );
  AOI22_X1 U96 ( .A1(data_in[2]), .A2(n838), .B1(n1062), .B2(\mem[5][2] ), 
        .ZN(n1060) );
  INV_X1 U97 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U98 ( .A1(data_in[3]), .A2(n838), .B1(n1062), .B2(\mem[5][3] ), 
        .ZN(n1059) );
  INV_X1 U99 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U100 ( .A1(data_in[4]), .A2(n838), .B1(n1062), .B2(\mem[5][4] ), 
        .ZN(n1058) );
  INV_X1 U101 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U102 ( .A1(data_in[5]), .A2(n838), .B1(n1062), .B2(\mem[5][5] ), 
        .ZN(n1057) );
  INV_X1 U103 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U104 ( .A1(data_in[6]), .A2(n838), .B1(n1062), .B2(\mem[5][6] ), 
        .ZN(n1056) );
  INV_X1 U105 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U106 ( .A1(data_in[7]), .A2(n838), .B1(n1062), .B2(\mem[5][7] ), 
        .ZN(n1055) );
  INV_X1 U107 ( .A(n1026), .ZN(n739) );
  AOI22_X1 U108 ( .A1(data_in[0]), .A2(n834), .B1(n1025), .B2(\mem[9][0] ), 
        .ZN(n1026) );
  INV_X1 U109 ( .A(n1024), .ZN(n738) );
  AOI22_X1 U110 ( .A1(data_in[1]), .A2(n834), .B1(n1025), .B2(\mem[9][1] ), 
        .ZN(n1024) );
  INV_X1 U111 ( .A(n1023), .ZN(n737) );
  AOI22_X1 U112 ( .A1(data_in[2]), .A2(n834), .B1(n1025), .B2(\mem[9][2] ), 
        .ZN(n1023) );
  INV_X1 U113 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U114 ( .A1(data_in[3]), .A2(n834), .B1(n1025), .B2(\mem[9][3] ), 
        .ZN(n1022) );
  INV_X1 U115 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U116 ( .A1(data_in[4]), .A2(n834), .B1(n1025), .B2(\mem[9][4] ), 
        .ZN(n1021) );
  INV_X1 U117 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U118 ( .A1(data_in[5]), .A2(n834), .B1(n1025), .B2(\mem[9][5] ), 
        .ZN(n1020) );
  INV_X1 U119 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U120 ( .A1(data_in[6]), .A2(n834), .B1(n1025), .B2(\mem[9][6] ), 
        .ZN(n1019) );
  INV_X1 U121 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U122 ( .A1(data_in[7]), .A2(n834), .B1(n1025), .B2(\mem[9][7] ), 
        .ZN(n1018) );
  INV_X1 U123 ( .A(n990), .ZN(n707) );
  AOI22_X1 U124 ( .A1(data_in[0]), .A2(n830), .B1(n989), .B2(\mem[13][0] ), 
        .ZN(n990) );
  INV_X1 U125 ( .A(n988), .ZN(n706) );
  AOI22_X1 U126 ( .A1(data_in[1]), .A2(n830), .B1(n989), .B2(\mem[13][1] ), 
        .ZN(n988) );
  INV_X1 U127 ( .A(n987), .ZN(n705) );
  AOI22_X1 U128 ( .A1(data_in[2]), .A2(n830), .B1(n989), .B2(\mem[13][2] ), 
        .ZN(n987) );
  INV_X1 U129 ( .A(n986), .ZN(n704) );
  AOI22_X1 U130 ( .A1(data_in[3]), .A2(n830), .B1(n989), .B2(\mem[13][3] ), 
        .ZN(n986) );
  INV_X1 U131 ( .A(n985), .ZN(n703) );
  AOI22_X1 U132 ( .A1(data_in[4]), .A2(n830), .B1(n989), .B2(\mem[13][4] ), 
        .ZN(n985) );
  INV_X1 U133 ( .A(n984), .ZN(n702) );
  AOI22_X1 U134 ( .A1(data_in[5]), .A2(n830), .B1(n989), .B2(\mem[13][5] ), 
        .ZN(n984) );
  INV_X1 U135 ( .A(n983), .ZN(n701) );
  AOI22_X1 U136 ( .A1(data_in[6]), .A2(n830), .B1(n989), .B2(\mem[13][6] ), 
        .ZN(n983) );
  INV_X1 U137 ( .A(n982), .ZN(n700) );
  AOI22_X1 U138 ( .A1(data_in[7]), .A2(n830), .B1(n989), .B2(\mem[13][7] ), 
        .ZN(n982) );
  INV_X1 U139 ( .A(n915), .ZN(n642) );
  AOI22_X1 U140 ( .A1(data_in[1]), .A2(n822), .B1(n916), .B2(\mem[21][1] ), 
        .ZN(n915) );
  INV_X1 U141 ( .A(n914), .ZN(n641) );
  AOI22_X1 U142 ( .A1(data_in[2]), .A2(n822), .B1(n916), .B2(\mem[21][2] ), 
        .ZN(n914) );
  INV_X1 U143 ( .A(n913), .ZN(n640) );
  AOI22_X1 U144 ( .A1(data_in[3]), .A2(n822), .B1(n916), .B2(\mem[21][3] ), 
        .ZN(n913) );
  INV_X1 U145 ( .A(n912), .ZN(n639) );
  AOI22_X1 U146 ( .A1(data_in[4]), .A2(n822), .B1(n916), .B2(\mem[21][4] ), 
        .ZN(n912) );
  INV_X1 U147 ( .A(n911), .ZN(n638) );
  AOI22_X1 U148 ( .A1(data_in[5]), .A2(n822), .B1(n916), .B2(\mem[21][5] ), 
        .ZN(n911) );
  INV_X1 U149 ( .A(n910), .ZN(n637) );
  AOI22_X1 U150 ( .A1(data_in[6]), .A2(n822), .B1(n916), .B2(\mem[21][6] ), 
        .ZN(n910) );
  INV_X1 U151 ( .A(n909), .ZN(n636) );
  AOI22_X1 U152 ( .A1(data_in[7]), .A2(n822), .B1(n916), .B2(\mem[21][7] ), 
        .ZN(n909) );
  INV_X1 U153 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U154 ( .A1(data_in[0]), .A2(n837), .B1(n1053), .B2(\mem[6][0] ), 
        .ZN(n1054) );
  INV_X1 U155 ( .A(n1052), .ZN(n762) );
  AOI22_X1 U156 ( .A1(data_in[1]), .A2(n837), .B1(n1053), .B2(\mem[6][1] ), 
        .ZN(n1052) );
  INV_X1 U157 ( .A(n1051), .ZN(n761) );
  AOI22_X1 U158 ( .A1(data_in[2]), .A2(n837), .B1(n1053), .B2(\mem[6][2] ), 
        .ZN(n1051) );
  INV_X1 U159 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U160 ( .A1(data_in[3]), .A2(n837), .B1(n1053), .B2(\mem[6][3] ), 
        .ZN(n1050) );
  INV_X1 U161 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U162 ( .A1(data_in[4]), .A2(n837), .B1(n1053), .B2(\mem[6][4] ), 
        .ZN(n1049) );
  INV_X1 U163 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U164 ( .A1(data_in[5]), .A2(n837), .B1(n1053), .B2(\mem[6][5] ), 
        .ZN(n1048) );
  INV_X1 U165 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U166 ( .A1(data_in[6]), .A2(n837), .B1(n1053), .B2(\mem[6][6] ), 
        .ZN(n1047) );
  INV_X1 U167 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U168 ( .A1(data_in[7]), .A2(n837), .B1(n1053), .B2(\mem[6][7] ), 
        .ZN(n1046) );
  INV_X1 U169 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U170 ( .A1(data_in[0]), .A2(n836), .B1(n1044), .B2(\mem[7][0] ), 
        .ZN(n1045) );
  INV_X1 U171 ( .A(n1043), .ZN(n754) );
  AOI22_X1 U172 ( .A1(data_in[1]), .A2(n836), .B1(n1044), .B2(\mem[7][1] ), 
        .ZN(n1043) );
  INV_X1 U173 ( .A(n1042), .ZN(n753) );
  AOI22_X1 U174 ( .A1(data_in[2]), .A2(n836), .B1(n1044), .B2(\mem[7][2] ), 
        .ZN(n1042) );
  INV_X1 U175 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U176 ( .A1(data_in[3]), .A2(n836), .B1(n1044), .B2(\mem[7][3] ), 
        .ZN(n1041) );
  INV_X1 U177 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U178 ( .A1(data_in[4]), .A2(n836), .B1(n1044), .B2(\mem[7][4] ), 
        .ZN(n1040) );
  INV_X1 U179 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U180 ( .A1(data_in[5]), .A2(n836), .B1(n1044), .B2(\mem[7][5] ), 
        .ZN(n1039) );
  INV_X1 U181 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U182 ( .A1(data_in[6]), .A2(n836), .B1(n1044), .B2(\mem[7][6] ), 
        .ZN(n1038) );
  INV_X1 U183 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U184 ( .A1(data_in[7]), .A2(n836), .B1(n1044), .B2(\mem[7][7] ), 
        .ZN(n1037) );
  INV_X1 U185 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U186 ( .A1(data_in[0]), .A2(n833), .B1(n1016), .B2(\mem[10][0] ), 
        .ZN(n1017) );
  INV_X1 U187 ( .A(n1015), .ZN(n730) );
  AOI22_X1 U188 ( .A1(data_in[1]), .A2(n833), .B1(n1016), .B2(\mem[10][1] ), 
        .ZN(n1015) );
  INV_X1 U189 ( .A(n1014), .ZN(n729) );
  AOI22_X1 U190 ( .A1(data_in[2]), .A2(n833), .B1(n1016), .B2(\mem[10][2] ), 
        .ZN(n1014) );
  INV_X1 U191 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U192 ( .A1(data_in[3]), .A2(n833), .B1(n1016), .B2(\mem[10][3] ), 
        .ZN(n1013) );
  INV_X1 U193 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U194 ( .A1(data_in[4]), .A2(n833), .B1(n1016), .B2(\mem[10][4] ), 
        .ZN(n1012) );
  INV_X1 U195 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U196 ( .A1(data_in[5]), .A2(n833), .B1(n1016), .B2(\mem[10][5] ), 
        .ZN(n1011) );
  INV_X1 U197 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U198 ( .A1(data_in[6]), .A2(n833), .B1(n1016), .B2(\mem[10][6] ), 
        .ZN(n1010) );
  INV_X1 U199 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U200 ( .A1(data_in[7]), .A2(n833), .B1(n1016), .B2(\mem[10][7] ), 
        .ZN(n1009) );
  INV_X1 U201 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U202 ( .A1(data_in[0]), .A2(n832), .B1(n1007), .B2(\mem[11][0] ), 
        .ZN(n1008) );
  INV_X1 U203 ( .A(n1006), .ZN(n722) );
  AOI22_X1 U204 ( .A1(data_in[1]), .A2(n832), .B1(n1007), .B2(\mem[11][1] ), 
        .ZN(n1006) );
  INV_X1 U205 ( .A(n1005), .ZN(n721) );
  AOI22_X1 U206 ( .A1(data_in[2]), .A2(n832), .B1(n1007), .B2(\mem[11][2] ), 
        .ZN(n1005) );
  INV_X1 U207 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U208 ( .A1(data_in[3]), .A2(n832), .B1(n1007), .B2(\mem[11][3] ), 
        .ZN(n1004) );
  INV_X1 U209 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U210 ( .A1(data_in[4]), .A2(n832), .B1(n1007), .B2(\mem[11][4] ), 
        .ZN(n1003) );
  INV_X1 U211 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U212 ( .A1(data_in[5]), .A2(n832), .B1(n1007), .B2(\mem[11][5] ), 
        .ZN(n1002) );
  INV_X1 U213 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U214 ( .A1(data_in[6]), .A2(n832), .B1(n1007), .B2(\mem[11][6] ), 
        .ZN(n1001) );
  INV_X1 U215 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U216 ( .A1(data_in[7]), .A2(n832), .B1(n1007), .B2(\mem[11][7] ), 
        .ZN(n1000) );
  INV_X1 U217 ( .A(n953), .ZN(n675) );
  AOI22_X1 U218 ( .A1(data_in[0]), .A2(n826), .B1(n952), .B2(\mem[17][0] ), 
        .ZN(n953) );
  INV_X1 U219 ( .A(n951), .ZN(n674) );
  AOI22_X1 U220 ( .A1(data_in[1]), .A2(n826), .B1(n952), .B2(\mem[17][1] ), 
        .ZN(n951) );
  INV_X1 U221 ( .A(n950), .ZN(n673) );
  AOI22_X1 U222 ( .A1(data_in[2]), .A2(n826), .B1(n952), .B2(\mem[17][2] ), 
        .ZN(n950) );
  INV_X1 U223 ( .A(n949), .ZN(n672) );
  AOI22_X1 U224 ( .A1(data_in[3]), .A2(n826), .B1(n952), .B2(\mem[17][3] ), 
        .ZN(n949) );
  INV_X1 U225 ( .A(n948), .ZN(n671) );
  AOI22_X1 U226 ( .A1(data_in[4]), .A2(n826), .B1(n952), .B2(\mem[17][4] ), 
        .ZN(n948) );
  INV_X1 U227 ( .A(n947), .ZN(n670) );
  AOI22_X1 U228 ( .A1(data_in[5]), .A2(n826), .B1(n952), .B2(\mem[17][5] ), 
        .ZN(n947) );
  INV_X1 U229 ( .A(n946), .ZN(n669) );
  AOI22_X1 U230 ( .A1(data_in[6]), .A2(n826), .B1(n952), .B2(\mem[17][6] ), 
        .ZN(n946) );
  INV_X1 U231 ( .A(n945), .ZN(n668) );
  AOI22_X1 U232 ( .A1(data_in[7]), .A2(n826), .B1(n952), .B2(\mem[17][7] ), 
        .ZN(n945) );
  INV_X1 U233 ( .A(n917), .ZN(n643) );
  AOI22_X1 U234 ( .A1(data_in[0]), .A2(n822), .B1(n916), .B2(\mem[21][0] ), 
        .ZN(n917) );
  INV_X1 U235 ( .A(n981), .ZN(n699) );
  AOI22_X1 U236 ( .A1(data_in[0]), .A2(n829), .B1(n980), .B2(\mem[14][0] ), 
        .ZN(n981) );
  INV_X1 U237 ( .A(n979), .ZN(n698) );
  AOI22_X1 U238 ( .A1(data_in[1]), .A2(n829), .B1(n980), .B2(\mem[14][1] ), 
        .ZN(n979) );
  INV_X1 U239 ( .A(n978), .ZN(n697) );
  AOI22_X1 U240 ( .A1(data_in[2]), .A2(n829), .B1(n980), .B2(\mem[14][2] ), 
        .ZN(n978) );
  INV_X1 U241 ( .A(n977), .ZN(n696) );
  AOI22_X1 U242 ( .A1(data_in[3]), .A2(n829), .B1(n980), .B2(\mem[14][3] ), 
        .ZN(n977) );
  INV_X1 U243 ( .A(n976), .ZN(n695) );
  AOI22_X1 U244 ( .A1(data_in[4]), .A2(n829), .B1(n980), .B2(\mem[14][4] ), 
        .ZN(n976) );
  INV_X1 U245 ( .A(n975), .ZN(n694) );
  AOI22_X1 U246 ( .A1(data_in[5]), .A2(n829), .B1(n980), .B2(\mem[14][5] ), 
        .ZN(n975) );
  INV_X1 U247 ( .A(n974), .ZN(n693) );
  AOI22_X1 U248 ( .A1(data_in[6]), .A2(n829), .B1(n980), .B2(\mem[14][6] ), 
        .ZN(n974) );
  INV_X1 U249 ( .A(n973), .ZN(n692) );
  AOI22_X1 U250 ( .A1(data_in[7]), .A2(n829), .B1(n980), .B2(\mem[14][7] ), 
        .ZN(n973) );
  INV_X1 U251 ( .A(n972), .ZN(n691) );
  AOI22_X1 U252 ( .A1(data_in[0]), .A2(n828), .B1(n971), .B2(\mem[15][0] ), 
        .ZN(n972) );
  INV_X1 U253 ( .A(n970), .ZN(n690) );
  AOI22_X1 U254 ( .A1(data_in[1]), .A2(n828), .B1(n971), .B2(\mem[15][1] ), 
        .ZN(n970) );
  INV_X1 U255 ( .A(n969), .ZN(n689) );
  AOI22_X1 U256 ( .A1(data_in[2]), .A2(n828), .B1(n971), .B2(\mem[15][2] ), 
        .ZN(n969) );
  INV_X1 U257 ( .A(n968), .ZN(n688) );
  AOI22_X1 U258 ( .A1(data_in[3]), .A2(n828), .B1(n971), .B2(\mem[15][3] ), 
        .ZN(n968) );
  INV_X1 U259 ( .A(n967), .ZN(n687) );
  AOI22_X1 U260 ( .A1(data_in[4]), .A2(n828), .B1(n971), .B2(\mem[15][4] ), 
        .ZN(n967) );
  INV_X1 U261 ( .A(n966), .ZN(n686) );
  AOI22_X1 U262 ( .A1(data_in[5]), .A2(n828), .B1(n971), .B2(\mem[15][5] ), 
        .ZN(n966) );
  INV_X1 U263 ( .A(n965), .ZN(n685) );
  AOI22_X1 U264 ( .A1(data_in[6]), .A2(n828), .B1(n971), .B2(\mem[15][6] ), 
        .ZN(n965) );
  INV_X1 U265 ( .A(n964), .ZN(n684) );
  AOI22_X1 U266 ( .A1(data_in[7]), .A2(n828), .B1(n971), .B2(\mem[15][7] ), 
        .ZN(n964) );
  INV_X1 U267 ( .A(n944), .ZN(n667) );
  AOI22_X1 U268 ( .A1(data_in[0]), .A2(n825), .B1(n943), .B2(\mem[18][0] ), 
        .ZN(n944) );
  INV_X1 U269 ( .A(n942), .ZN(n666) );
  AOI22_X1 U270 ( .A1(data_in[1]), .A2(n825), .B1(n943), .B2(\mem[18][1] ), 
        .ZN(n942) );
  INV_X1 U271 ( .A(n941), .ZN(n665) );
  AOI22_X1 U272 ( .A1(data_in[2]), .A2(n825), .B1(n943), .B2(\mem[18][2] ), 
        .ZN(n941) );
  INV_X1 U273 ( .A(n940), .ZN(n664) );
  AOI22_X1 U274 ( .A1(data_in[3]), .A2(n825), .B1(n943), .B2(\mem[18][3] ), 
        .ZN(n940) );
  INV_X1 U275 ( .A(n939), .ZN(n663) );
  AOI22_X1 U276 ( .A1(data_in[4]), .A2(n825), .B1(n943), .B2(\mem[18][4] ), 
        .ZN(n939) );
  INV_X1 U277 ( .A(n938), .ZN(n662) );
  AOI22_X1 U278 ( .A1(data_in[5]), .A2(n825), .B1(n943), .B2(\mem[18][5] ), 
        .ZN(n938) );
  INV_X1 U279 ( .A(n937), .ZN(n661) );
  AOI22_X1 U280 ( .A1(data_in[6]), .A2(n825), .B1(n943), .B2(\mem[18][6] ), 
        .ZN(n937) );
  INV_X1 U281 ( .A(n936), .ZN(n660) );
  AOI22_X1 U282 ( .A1(data_in[7]), .A2(n825), .B1(n943), .B2(\mem[18][7] ), 
        .ZN(n936) );
  INV_X1 U283 ( .A(n935), .ZN(n659) );
  AOI22_X1 U284 ( .A1(data_in[0]), .A2(n824), .B1(n934), .B2(\mem[19][0] ), 
        .ZN(n935) );
  INV_X1 U285 ( .A(n933), .ZN(n658) );
  AOI22_X1 U286 ( .A1(data_in[1]), .A2(n824), .B1(n934), .B2(\mem[19][1] ), 
        .ZN(n933) );
  INV_X1 U287 ( .A(n932), .ZN(n657) );
  AOI22_X1 U288 ( .A1(data_in[2]), .A2(n824), .B1(n934), .B2(\mem[19][2] ), 
        .ZN(n932) );
  INV_X1 U289 ( .A(n931), .ZN(n656) );
  AOI22_X1 U290 ( .A1(data_in[3]), .A2(n824), .B1(n934), .B2(\mem[19][3] ), 
        .ZN(n931) );
  INV_X1 U291 ( .A(n930), .ZN(n655) );
  AOI22_X1 U292 ( .A1(data_in[4]), .A2(n824), .B1(n934), .B2(\mem[19][4] ), 
        .ZN(n930) );
  INV_X1 U293 ( .A(n929), .ZN(n654) );
  AOI22_X1 U294 ( .A1(data_in[5]), .A2(n824), .B1(n934), .B2(\mem[19][5] ), 
        .ZN(n929) );
  INV_X1 U295 ( .A(n928), .ZN(n653) );
  AOI22_X1 U296 ( .A1(data_in[6]), .A2(n824), .B1(n934), .B2(\mem[19][6] ), 
        .ZN(n928) );
  INV_X1 U297 ( .A(n927), .ZN(n652) );
  AOI22_X1 U298 ( .A1(data_in[7]), .A2(n824), .B1(n934), .B2(\mem[19][7] ), 
        .ZN(n927) );
  INV_X1 U299 ( .A(n908), .ZN(n635) );
  AOI22_X1 U300 ( .A1(data_in[0]), .A2(n821), .B1(n907), .B2(\mem[22][0] ), 
        .ZN(n908) );
  INV_X1 U301 ( .A(n906), .ZN(n634) );
  AOI22_X1 U302 ( .A1(data_in[1]), .A2(n821), .B1(n907), .B2(\mem[22][1] ), 
        .ZN(n906) );
  INV_X1 U303 ( .A(n905), .ZN(n633) );
  AOI22_X1 U304 ( .A1(data_in[2]), .A2(n821), .B1(n907), .B2(\mem[22][2] ), 
        .ZN(n905) );
  INV_X1 U305 ( .A(n904), .ZN(n632) );
  AOI22_X1 U306 ( .A1(data_in[3]), .A2(n821), .B1(n907), .B2(\mem[22][3] ), 
        .ZN(n904) );
  INV_X1 U307 ( .A(n903), .ZN(n631) );
  AOI22_X1 U308 ( .A1(data_in[4]), .A2(n821), .B1(n907), .B2(\mem[22][4] ), 
        .ZN(n903) );
  INV_X1 U309 ( .A(n902), .ZN(n630) );
  AOI22_X1 U310 ( .A1(data_in[5]), .A2(n821), .B1(n907), .B2(\mem[22][5] ), 
        .ZN(n902) );
  INV_X1 U311 ( .A(n901), .ZN(n629) );
  AOI22_X1 U312 ( .A1(data_in[6]), .A2(n821), .B1(n907), .B2(\mem[22][6] ), 
        .ZN(n901) );
  INV_X1 U313 ( .A(n900), .ZN(n628) );
  AOI22_X1 U314 ( .A1(data_in[7]), .A2(n821), .B1(n907), .B2(\mem[22][7] ), 
        .ZN(n900) );
  INV_X1 U315 ( .A(n899), .ZN(n627) );
  AOI22_X1 U316 ( .A1(data_in[0]), .A2(n820), .B1(n898), .B2(\mem[23][0] ), 
        .ZN(n899) );
  INV_X1 U317 ( .A(n897), .ZN(n626) );
  AOI22_X1 U318 ( .A1(data_in[1]), .A2(n820), .B1(n898), .B2(\mem[23][1] ), 
        .ZN(n897) );
  INV_X1 U319 ( .A(n896), .ZN(n625) );
  AOI22_X1 U320 ( .A1(data_in[2]), .A2(n820), .B1(n898), .B2(\mem[23][2] ), 
        .ZN(n896) );
  INV_X1 U321 ( .A(n895), .ZN(n624) );
  AOI22_X1 U322 ( .A1(data_in[3]), .A2(n820), .B1(n898), .B2(\mem[23][3] ), 
        .ZN(n895) );
  INV_X1 U323 ( .A(n894), .ZN(n623) );
  AOI22_X1 U324 ( .A1(data_in[4]), .A2(n820), .B1(n898), .B2(\mem[23][4] ), 
        .ZN(n894) );
  INV_X1 U325 ( .A(n893), .ZN(n622) );
  AOI22_X1 U326 ( .A1(data_in[5]), .A2(n820), .B1(n898), .B2(\mem[23][5] ), 
        .ZN(n893) );
  INV_X1 U327 ( .A(n892), .ZN(n621) );
  AOI22_X1 U328 ( .A1(data_in[6]), .A2(n820), .B1(n898), .B2(\mem[23][6] ), 
        .ZN(n892) );
  INV_X1 U329 ( .A(n891), .ZN(n620) );
  AOI22_X1 U330 ( .A1(data_in[7]), .A2(n820), .B1(n898), .B2(\mem[23][7] ), 
        .ZN(n891) );
  INV_X1 U331 ( .A(N12), .ZN(n255) );
  INV_X1 U332 ( .A(N11), .ZN(n254) );
  INV_X1 U333 ( .A(n999), .ZN(n715) );
  AOI22_X1 U334 ( .A1(data_in[0]), .A2(n831), .B1(n998), .B2(\mem[12][0] ), 
        .ZN(n999) );
  INV_X1 U335 ( .A(n997), .ZN(n714) );
  AOI22_X1 U336 ( .A1(data_in[1]), .A2(n831), .B1(n998), .B2(\mem[12][1] ), 
        .ZN(n997) );
  INV_X1 U337 ( .A(n996), .ZN(n713) );
  AOI22_X1 U338 ( .A1(data_in[2]), .A2(n831), .B1(n998), .B2(\mem[12][2] ), 
        .ZN(n996) );
  INV_X1 U339 ( .A(n995), .ZN(n712) );
  AOI22_X1 U340 ( .A1(data_in[3]), .A2(n831), .B1(n998), .B2(\mem[12][3] ), 
        .ZN(n995) );
  INV_X1 U341 ( .A(n994), .ZN(n711) );
  AOI22_X1 U342 ( .A1(data_in[4]), .A2(n831), .B1(n998), .B2(\mem[12][4] ), 
        .ZN(n994) );
  INV_X1 U343 ( .A(n993), .ZN(n710) );
  AOI22_X1 U344 ( .A1(data_in[5]), .A2(n831), .B1(n998), .B2(\mem[12][5] ), 
        .ZN(n993) );
  INV_X1 U345 ( .A(n992), .ZN(n709) );
  AOI22_X1 U346 ( .A1(data_in[6]), .A2(n831), .B1(n998), .B2(\mem[12][6] ), 
        .ZN(n992) );
  INV_X1 U347 ( .A(n991), .ZN(n708) );
  AOI22_X1 U348 ( .A1(data_in[7]), .A2(n831), .B1(n998), .B2(\mem[12][7] ), 
        .ZN(n991) );
  INV_X1 U349 ( .A(n926), .ZN(n651) );
  AOI22_X1 U350 ( .A1(data_in[0]), .A2(n823), .B1(n925), .B2(\mem[20][0] ), 
        .ZN(n926) );
  INV_X1 U351 ( .A(n924), .ZN(n650) );
  AOI22_X1 U352 ( .A1(data_in[1]), .A2(n823), .B1(n925), .B2(\mem[20][1] ), 
        .ZN(n924) );
  INV_X1 U353 ( .A(n923), .ZN(n649) );
  AOI22_X1 U354 ( .A1(data_in[2]), .A2(n823), .B1(n925), .B2(\mem[20][2] ), 
        .ZN(n923) );
  INV_X1 U355 ( .A(n922), .ZN(n648) );
  AOI22_X1 U356 ( .A1(data_in[3]), .A2(n823), .B1(n925), .B2(\mem[20][3] ), 
        .ZN(n922) );
  INV_X1 U357 ( .A(n921), .ZN(n647) );
  AOI22_X1 U358 ( .A1(data_in[4]), .A2(n823), .B1(n925), .B2(\mem[20][4] ), 
        .ZN(n921) );
  INV_X1 U359 ( .A(n920), .ZN(n646) );
  AOI22_X1 U360 ( .A1(data_in[5]), .A2(n823), .B1(n925), .B2(\mem[20][5] ), 
        .ZN(n920) );
  INV_X1 U361 ( .A(n919), .ZN(n645) );
  AOI22_X1 U362 ( .A1(data_in[6]), .A2(n823), .B1(n925), .B2(\mem[20][6] ), 
        .ZN(n919) );
  INV_X1 U363 ( .A(n918), .ZN(n644) );
  AOI22_X1 U364 ( .A1(data_in[7]), .A2(n823), .B1(n925), .B2(\mem[20][7] ), 
        .ZN(n918) );
  INV_X1 U365 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U366 ( .A1(data_in[0]), .A2(n835), .B1(n1035), .B2(\mem[8][0] ), 
        .ZN(n1036) );
  INV_X1 U367 ( .A(n1034), .ZN(n746) );
  AOI22_X1 U368 ( .A1(data_in[1]), .A2(n835), .B1(n1035), .B2(\mem[8][1] ), 
        .ZN(n1034) );
  INV_X1 U369 ( .A(n1033), .ZN(n745) );
  AOI22_X1 U370 ( .A1(data_in[2]), .A2(n835), .B1(n1035), .B2(\mem[8][2] ), 
        .ZN(n1033) );
  INV_X1 U371 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U372 ( .A1(data_in[3]), .A2(n835), .B1(n1035), .B2(\mem[8][3] ), 
        .ZN(n1032) );
  INV_X1 U373 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U374 ( .A1(data_in[4]), .A2(n835), .B1(n1035), .B2(\mem[8][4] ), 
        .ZN(n1031) );
  INV_X1 U375 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U376 ( .A1(data_in[5]), .A2(n835), .B1(n1035), .B2(\mem[8][5] ), 
        .ZN(n1030) );
  INV_X1 U377 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U378 ( .A1(data_in[6]), .A2(n835), .B1(n1035), .B2(\mem[8][6] ), 
        .ZN(n1029) );
  INV_X1 U379 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U380 ( .A1(data_in[7]), .A2(n835), .B1(n1035), .B2(\mem[8][7] ), 
        .ZN(n1028) );
  INV_X1 U381 ( .A(n963), .ZN(n683) );
  AOI22_X1 U382 ( .A1(data_in[0]), .A2(n827), .B1(n962), .B2(\mem[16][0] ), 
        .ZN(n963) );
  INV_X1 U383 ( .A(n961), .ZN(n682) );
  AOI22_X1 U384 ( .A1(data_in[1]), .A2(n827), .B1(n962), .B2(\mem[16][1] ), 
        .ZN(n961) );
  INV_X1 U385 ( .A(n960), .ZN(n681) );
  AOI22_X1 U386 ( .A1(data_in[2]), .A2(n827), .B1(n962), .B2(\mem[16][2] ), 
        .ZN(n960) );
  INV_X1 U387 ( .A(n959), .ZN(n680) );
  AOI22_X1 U388 ( .A1(data_in[3]), .A2(n827), .B1(n962), .B2(\mem[16][3] ), 
        .ZN(n959) );
  INV_X1 U389 ( .A(n958), .ZN(n679) );
  AOI22_X1 U390 ( .A1(data_in[4]), .A2(n827), .B1(n962), .B2(\mem[16][4] ), 
        .ZN(n958) );
  INV_X1 U391 ( .A(n957), .ZN(n678) );
  AOI22_X1 U392 ( .A1(data_in[5]), .A2(n827), .B1(n962), .B2(\mem[16][5] ), 
        .ZN(n957) );
  INV_X1 U393 ( .A(n956), .ZN(n677) );
  AOI22_X1 U394 ( .A1(data_in[6]), .A2(n827), .B1(n962), .B2(\mem[16][6] ), 
        .ZN(n956) );
  INV_X1 U395 ( .A(n955), .ZN(n676) );
  AOI22_X1 U396 ( .A1(data_in[7]), .A2(n827), .B1(n962), .B2(\mem[16][7] ), 
        .ZN(n955) );
  INV_X1 U397 ( .A(n890), .ZN(n619) );
  AOI22_X1 U398 ( .A1(data_in[0]), .A2(n816), .B1(n889), .B2(\mem[24][0] ), 
        .ZN(n890) );
  INV_X1 U399 ( .A(n888), .ZN(n618) );
  AOI22_X1 U400 ( .A1(data_in[1]), .A2(n816), .B1(n889), .B2(\mem[24][1] ), 
        .ZN(n888) );
  INV_X1 U401 ( .A(n887), .ZN(n617) );
  AOI22_X1 U402 ( .A1(data_in[2]), .A2(n816), .B1(n889), .B2(\mem[24][2] ), 
        .ZN(n887) );
  INV_X1 U403 ( .A(n886), .ZN(n616) );
  AOI22_X1 U404 ( .A1(data_in[3]), .A2(n816), .B1(n889), .B2(\mem[24][3] ), 
        .ZN(n886) );
  INV_X1 U405 ( .A(n885), .ZN(n615) );
  AOI22_X1 U406 ( .A1(data_in[4]), .A2(n816), .B1(n889), .B2(\mem[24][4] ), 
        .ZN(n885) );
  INV_X1 U407 ( .A(n884), .ZN(n614) );
  AOI22_X1 U408 ( .A1(data_in[5]), .A2(n816), .B1(n889), .B2(\mem[24][5] ), 
        .ZN(n884) );
  INV_X1 U409 ( .A(n883), .ZN(n613) );
  AOI22_X1 U410 ( .A1(data_in[6]), .A2(n816), .B1(n889), .B2(\mem[24][6] ), 
        .ZN(n883) );
  INV_X1 U411 ( .A(n882), .ZN(n612) );
  AOI22_X1 U412 ( .A1(data_in[7]), .A2(n816), .B1(n889), .B2(\mem[24][7] ), 
        .ZN(n882) );
  INV_X1 U413 ( .A(n881), .ZN(n611) );
  AOI22_X1 U414 ( .A1(data_in[0]), .A2(n815), .B1(n880), .B2(\mem[25][0] ), 
        .ZN(n881) );
  INV_X1 U415 ( .A(n879), .ZN(n610) );
  AOI22_X1 U416 ( .A1(data_in[1]), .A2(n815), .B1(n880), .B2(\mem[25][1] ), 
        .ZN(n879) );
  INV_X1 U417 ( .A(n878), .ZN(n609) );
  AOI22_X1 U418 ( .A1(data_in[2]), .A2(n815), .B1(n880), .B2(\mem[25][2] ), 
        .ZN(n878) );
  INV_X1 U419 ( .A(n877), .ZN(n608) );
  AOI22_X1 U420 ( .A1(data_in[3]), .A2(n815), .B1(n880), .B2(\mem[25][3] ), 
        .ZN(n877) );
  INV_X1 U421 ( .A(n876), .ZN(n607) );
  AOI22_X1 U422 ( .A1(data_in[4]), .A2(n815), .B1(n880), .B2(\mem[25][4] ), 
        .ZN(n876) );
  INV_X1 U423 ( .A(n875), .ZN(n606) );
  AOI22_X1 U424 ( .A1(data_in[5]), .A2(n815), .B1(n880), .B2(\mem[25][5] ), 
        .ZN(n875) );
  INV_X1 U425 ( .A(n874), .ZN(n605) );
  AOI22_X1 U426 ( .A1(data_in[6]), .A2(n815), .B1(n880), .B2(\mem[25][6] ), 
        .ZN(n874) );
  INV_X1 U427 ( .A(n873), .ZN(n604) );
  AOI22_X1 U428 ( .A1(data_in[7]), .A2(n815), .B1(n880), .B2(\mem[25][7] ), 
        .ZN(n873) );
  INV_X1 U429 ( .A(n872), .ZN(n603) );
  AOI22_X1 U430 ( .A1(data_in[0]), .A2(n814), .B1(n871), .B2(\mem[26][0] ), 
        .ZN(n872) );
  INV_X1 U431 ( .A(n870), .ZN(n602) );
  AOI22_X1 U432 ( .A1(data_in[1]), .A2(n814), .B1(n871), .B2(\mem[26][1] ), 
        .ZN(n870) );
  INV_X1 U433 ( .A(n869), .ZN(n601) );
  AOI22_X1 U434 ( .A1(data_in[2]), .A2(n814), .B1(n871), .B2(\mem[26][2] ), 
        .ZN(n869) );
  INV_X1 U435 ( .A(n868), .ZN(n600) );
  AOI22_X1 U436 ( .A1(data_in[3]), .A2(n814), .B1(n871), .B2(\mem[26][3] ), 
        .ZN(n868) );
  INV_X1 U437 ( .A(n867), .ZN(n599) );
  AOI22_X1 U438 ( .A1(data_in[4]), .A2(n814), .B1(n871), .B2(\mem[26][4] ), 
        .ZN(n867) );
  INV_X1 U439 ( .A(n866), .ZN(n598) );
  AOI22_X1 U440 ( .A1(data_in[5]), .A2(n814), .B1(n871), .B2(\mem[26][5] ), 
        .ZN(n866) );
  INV_X1 U441 ( .A(n865), .ZN(n597) );
  AOI22_X1 U442 ( .A1(data_in[6]), .A2(n814), .B1(n871), .B2(\mem[26][6] ), 
        .ZN(n865) );
  INV_X1 U443 ( .A(n864), .ZN(n596) );
  AOI22_X1 U444 ( .A1(data_in[7]), .A2(n814), .B1(n871), .B2(\mem[26][7] ), 
        .ZN(n864) );
  INV_X1 U445 ( .A(n863), .ZN(n595) );
  AOI22_X1 U446 ( .A1(data_in[0]), .A2(n813), .B1(n862), .B2(\mem[27][0] ), 
        .ZN(n863) );
  INV_X1 U447 ( .A(n861), .ZN(n594) );
  AOI22_X1 U448 ( .A1(data_in[1]), .A2(n813), .B1(n862), .B2(\mem[27][1] ), 
        .ZN(n861) );
  INV_X1 U449 ( .A(n860), .ZN(n293) );
  AOI22_X1 U450 ( .A1(data_in[2]), .A2(n813), .B1(n862), .B2(\mem[27][2] ), 
        .ZN(n860) );
  INV_X1 U451 ( .A(n859), .ZN(n292) );
  AOI22_X1 U452 ( .A1(data_in[3]), .A2(n813), .B1(n862), .B2(\mem[27][3] ), 
        .ZN(n859) );
  INV_X1 U453 ( .A(n858), .ZN(n291) );
  AOI22_X1 U454 ( .A1(data_in[4]), .A2(n813), .B1(n862), .B2(\mem[27][4] ), 
        .ZN(n858) );
  INV_X1 U455 ( .A(n857), .ZN(n290) );
  AOI22_X1 U456 ( .A1(data_in[5]), .A2(n813), .B1(n862), .B2(\mem[27][5] ), 
        .ZN(n857) );
  INV_X1 U457 ( .A(n856), .ZN(n289) );
  AOI22_X1 U458 ( .A1(data_in[6]), .A2(n813), .B1(n862), .B2(\mem[27][6] ), 
        .ZN(n856) );
  INV_X1 U459 ( .A(n855), .ZN(n288) );
  AOI22_X1 U460 ( .A1(data_in[7]), .A2(n813), .B1(n862), .B2(\mem[27][7] ), 
        .ZN(n855) );
  INV_X1 U461 ( .A(n854), .ZN(n287) );
  AOI22_X1 U462 ( .A1(data_in[0]), .A2(n812), .B1(n853), .B2(\mem[28][0] ), 
        .ZN(n854) );
  INV_X1 U463 ( .A(n852), .ZN(n286) );
  AOI22_X1 U464 ( .A1(data_in[1]), .A2(n812), .B1(n853), .B2(\mem[28][1] ), 
        .ZN(n852) );
  INV_X1 U465 ( .A(n851), .ZN(n285) );
  AOI22_X1 U466 ( .A1(data_in[2]), .A2(n812), .B1(n853), .B2(\mem[28][2] ), 
        .ZN(n851) );
  INV_X1 U467 ( .A(n850), .ZN(n284) );
  AOI22_X1 U468 ( .A1(data_in[3]), .A2(n812), .B1(n853), .B2(\mem[28][3] ), 
        .ZN(n850) );
  INV_X1 U469 ( .A(n849), .ZN(n283) );
  AOI22_X1 U470 ( .A1(data_in[4]), .A2(n812), .B1(n853), .B2(\mem[28][4] ), 
        .ZN(n849) );
  INV_X1 U471 ( .A(n848), .ZN(n282) );
  AOI22_X1 U472 ( .A1(data_in[5]), .A2(n812), .B1(n853), .B2(\mem[28][5] ), 
        .ZN(n848) );
  INV_X1 U473 ( .A(n847), .ZN(n281) );
  AOI22_X1 U474 ( .A1(data_in[6]), .A2(n812), .B1(n853), .B2(\mem[28][6] ), 
        .ZN(n847) );
  INV_X1 U475 ( .A(n846), .ZN(n280) );
  AOI22_X1 U476 ( .A1(data_in[7]), .A2(n812), .B1(n853), .B2(\mem[28][7] ), 
        .ZN(n846) );
  INV_X1 U477 ( .A(n1145), .ZN(n279) );
  AOI22_X1 U478 ( .A1(n819), .A2(data_in[0]), .B1(n1144), .B2(\mem[29][0] ), 
        .ZN(n1145) );
  INV_X1 U479 ( .A(n1143), .ZN(n278) );
  AOI22_X1 U480 ( .A1(n819), .A2(data_in[1]), .B1(n1144), .B2(\mem[29][1] ), 
        .ZN(n1143) );
  INV_X1 U481 ( .A(n1142), .ZN(n277) );
  AOI22_X1 U482 ( .A1(n819), .A2(data_in[2]), .B1(n1144), .B2(\mem[29][2] ), 
        .ZN(n1142) );
  INV_X1 U483 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U484 ( .A1(n819), .A2(data_in[3]), .B1(n1144), .B2(\mem[29][3] ), 
        .ZN(n1141) );
  INV_X1 U485 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U486 ( .A1(n819), .A2(data_in[4]), .B1(n1144), .B2(\mem[29][4] ), 
        .ZN(n1140) );
  INV_X1 U487 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U488 ( .A1(n819), .A2(data_in[5]), .B1(n1144), .B2(\mem[29][5] ), 
        .ZN(n1139) );
  INV_X1 U489 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U490 ( .A1(n819), .A2(data_in[6]), .B1(n1144), .B2(\mem[29][6] ), 
        .ZN(n1138) );
  INV_X1 U491 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U492 ( .A1(n819), .A2(data_in[7]), .B1(n1144), .B2(\mem[29][7] ), 
        .ZN(n1137) );
  INV_X1 U493 ( .A(n1134), .ZN(n271) );
  AOI22_X1 U494 ( .A1(data_in[0]), .A2(n818), .B1(n1133), .B2(\mem[30][0] ), 
        .ZN(n1134) );
  INV_X1 U495 ( .A(n1132), .ZN(n270) );
  AOI22_X1 U496 ( .A1(data_in[1]), .A2(n818), .B1(n1133), .B2(\mem[30][1] ), 
        .ZN(n1132) );
  INV_X1 U497 ( .A(n1131), .ZN(n269) );
  AOI22_X1 U498 ( .A1(data_in[2]), .A2(n818), .B1(n1133), .B2(\mem[30][2] ), 
        .ZN(n1131) );
  INV_X1 U499 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U500 ( .A1(data_in[3]), .A2(n818), .B1(n1133), .B2(\mem[30][3] ), 
        .ZN(n1130) );
  INV_X1 U501 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U502 ( .A1(data_in[4]), .A2(n818), .B1(n1133), .B2(\mem[30][4] ), 
        .ZN(n1129) );
  INV_X1 U503 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U504 ( .A1(data_in[5]), .A2(n818), .B1(n1133), .B2(\mem[30][5] ), 
        .ZN(n1128) );
  INV_X1 U505 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U506 ( .A1(data_in[6]), .A2(n818), .B1(n1133), .B2(\mem[30][6] ), 
        .ZN(n1127) );
  INV_X1 U507 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U508 ( .A1(data_in[7]), .A2(n818), .B1(n1133), .B2(\mem[30][7] ), 
        .ZN(n1126) );
  INV_X1 U509 ( .A(n1124), .ZN(n263) );
  AOI22_X1 U510 ( .A1(data_in[0]), .A2(n817), .B1(n1123), .B2(\mem[31][0] ), 
        .ZN(n1124) );
  INV_X1 U511 ( .A(n1122), .ZN(n262) );
  AOI22_X1 U512 ( .A1(data_in[1]), .A2(n817), .B1(n1123), .B2(\mem[31][1] ), 
        .ZN(n1122) );
  INV_X1 U513 ( .A(n1121), .ZN(n261) );
  AOI22_X1 U514 ( .A1(data_in[2]), .A2(n817), .B1(n1123), .B2(\mem[31][2] ), 
        .ZN(n1121) );
  INV_X1 U515 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U516 ( .A1(data_in[3]), .A2(n817), .B1(n1123), .B2(\mem[31][3] ), 
        .ZN(n1120) );
  INV_X1 U517 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U518 ( .A1(data_in[4]), .A2(n817), .B1(n1123), .B2(\mem[31][4] ), 
        .ZN(n1119) );
  INV_X1 U519 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U520 ( .A1(data_in[5]), .A2(n817), .B1(n1123), .B2(\mem[31][5] ), 
        .ZN(n1118) );
  INV_X1 U521 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U522 ( .A1(data_in[6]), .A2(n817), .B1(n1123), .B2(\mem[31][6] ), 
        .ZN(n1117) );
  INV_X1 U523 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U524 ( .A1(data_in[7]), .A2(n817), .B1(n1123), .B2(\mem[31][7] ), 
        .ZN(n1116) );
  INV_X1 U525 ( .A(n1114), .ZN(n811) );
  AOI22_X1 U526 ( .A1(data_in[0]), .A2(n843), .B1(n1113), .B2(\mem[0][0] ), 
        .ZN(n1114) );
  INV_X1 U527 ( .A(n1112), .ZN(n810) );
  AOI22_X1 U528 ( .A1(data_in[1]), .A2(n843), .B1(n1113), .B2(\mem[0][1] ), 
        .ZN(n1112) );
  INV_X1 U529 ( .A(n1111), .ZN(n809) );
  AOI22_X1 U530 ( .A1(data_in[2]), .A2(n843), .B1(n1113), .B2(\mem[0][2] ), 
        .ZN(n1111) );
  INV_X1 U531 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U532 ( .A1(data_in[3]), .A2(n843), .B1(n1113), .B2(\mem[0][3] ), 
        .ZN(n1110) );
  INV_X1 U533 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U534 ( .A1(data_in[4]), .A2(n843), .B1(n1113), .B2(\mem[0][4] ), 
        .ZN(n1109) );
  INV_X1 U535 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U536 ( .A1(data_in[5]), .A2(n843), .B1(n1113), .B2(\mem[0][5] ), 
        .ZN(n1108) );
  INV_X1 U537 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U538 ( .A1(data_in[6]), .A2(n843), .B1(n1113), .B2(\mem[0][6] ), 
        .ZN(n1107) );
  INV_X1 U539 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U540 ( .A1(data_in[7]), .A2(n843), .B1(n1113), .B2(\mem[0][7] ), 
        .ZN(n1106) );
  INV_X1 U541 ( .A(n1103), .ZN(n803) );
  AOI22_X1 U542 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[1][0] ), 
        .ZN(n1103) );
  INV_X1 U543 ( .A(n1101), .ZN(n802) );
  AOI22_X1 U544 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[1][1] ), 
        .ZN(n1101) );
  INV_X1 U545 ( .A(n1100), .ZN(n801) );
  AOI22_X1 U546 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[1][2] ), 
        .ZN(n1100) );
  INV_X1 U547 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U548 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[1][3] ), 
        .ZN(n1099) );
  INV_X1 U549 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U550 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[1][4] ), 
        .ZN(n1098) );
  INV_X1 U551 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U552 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[1][5] ), 
        .ZN(n1097) );
  INV_X1 U553 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U554 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[1][6] ), 
        .ZN(n1096) );
  INV_X1 U555 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U556 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[1][7] ), 
        .ZN(n1095) );
  INV_X1 U557 ( .A(n1093), .ZN(n795) );
  AOI22_X1 U558 ( .A1(data_in[0]), .A2(n841), .B1(n1092), .B2(\mem[2][0] ), 
        .ZN(n1093) );
  INV_X1 U559 ( .A(n1091), .ZN(n794) );
  AOI22_X1 U560 ( .A1(data_in[1]), .A2(n841), .B1(n1092), .B2(\mem[2][1] ), 
        .ZN(n1091) );
  INV_X1 U561 ( .A(n1090), .ZN(n793) );
  AOI22_X1 U562 ( .A1(data_in[2]), .A2(n841), .B1(n1092), .B2(\mem[2][2] ), 
        .ZN(n1090) );
  INV_X1 U563 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U564 ( .A1(data_in[3]), .A2(n841), .B1(n1092), .B2(\mem[2][3] ), 
        .ZN(n1089) );
  INV_X1 U565 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U566 ( .A1(data_in[4]), .A2(n841), .B1(n1092), .B2(\mem[2][4] ), 
        .ZN(n1088) );
  INV_X1 U567 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U568 ( .A1(data_in[5]), .A2(n841), .B1(n1092), .B2(\mem[2][5] ), 
        .ZN(n1087) );
  INV_X1 U569 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U570 ( .A1(data_in[6]), .A2(n841), .B1(n1092), .B2(\mem[2][6] ), 
        .ZN(n1086) );
  INV_X1 U571 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U572 ( .A1(data_in[7]), .A2(n841), .B1(n1092), .B2(\mem[2][7] ), 
        .ZN(n1085) );
  INV_X1 U573 ( .A(n1083), .ZN(n787) );
  AOI22_X1 U574 ( .A1(data_in[0]), .A2(n840), .B1(n1082), .B2(\mem[3][0] ), 
        .ZN(n1083) );
  INV_X1 U575 ( .A(n1081), .ZN(n786) );
  AOI22_X1 U576 ( .A1(data_in[1]), .A2(n840), .B1(n1082), .B2(\mem[3][1] ), 
        .ZN(n1081) );
  INV_X1 U577 ( .A(n1080), .ZN(n785) );
  AOI22_X1 U578 ( .A1(data_in[2]), .A2(n840), .B1(n1082), .B2(\mem[3][2] ), 
        .ZN(n1080) );
  INV_X1 U579 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U580 ( .A1(data_in[3]), .A2(n840), .B1(n1082), .B2(\mem[3][3] ), 
        .ZN(n1079) );
  INV_X1 U581 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U582 ( .A1(data_in[4]), .A2(n840), .B1(n1082), .B2(\mem[3][4] ), 
        .ZN(n1078) );
  INV_X1 U583 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U584 ( .A1(data_in[5]), .A2(n840), .B1(n1082), .B2(\mem[3][5] ), 
        .ZN(n1077) );
  INV_X1 U585 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U586 ( .A1(data_in[6]), .A2(n840), .B1(n1082), .B2(\mem[3][6] ), 
        .ZN(n1076) );
  INV_X1 U587 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U588 ( .A1(data_in[7]), .A2(n840), .B1(n1082), .B2(\mem[3][7] ), 
        .ZN(n1075) );
  INV_X1 U589 ( .A(n1073), .ZN(n779) );
  AOI22_X1 U590 ( .A1(data_in[0]), .A2(n839), .B1(n1072), .B2(\mem[4][0] ), 
        .ZN(n1073) );
  INV_X1 U591 ( .A(n1071), .ZN(n778) );
  AOI22_X1 U592 ( .A1(data_in[1]), .A2(n839), .B1(n1072), .B2(\mem[4][1] ), 
        .ZN(n1071) );
  INV_X1 U593 ( .A(n1070), .ZN(n777) );
  AOI22_X1 U594 ( .A1(data_in[2]), .A2(n839), .B1(n1072), .B2(\mem[4][2] ), 
        .ZN(n1070) );
  INV_X1 U595 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U596 ( .A1(data_in[3]), .A2(n839), .B1(n1072), .B2(\mem[4][3] ), 
        .ZN(n1069) );
  INV_X1 U597 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U598 ( .A1(data_in[4]), .A2(n839), .B1(n1072), .B2(\mem[4][4] ), 
        .ZN(n1068) );
  INV_X1 U599 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U600 ( .A1(data_in[5]), .A2(n839), .B1(n1072), .B2(\mem[4][5] ), 
        .ZN(n1067) );
  INV_X1 U601 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U602 ( .A1(data_in[6]), .A2(n839), .B1(n1072), .B2(\mem[4][6] ), 
        .ZN(n1066) );
  INV_X1 U603 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U604 ( .A1(data_in[7]), .A2(n839), .B1(n1072), .B2(\mem[4][7] ), 
        .ZN(n1065) );
  INV_X1 U605 ( .A(N13), .ZN(n844) );
  INV_X1 U606 ( .A(N14), .ZN(n845) );
  MUX2_X1 U607 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n251), .Z(n3) );
  MUX2_X1 U608 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n251), .Z(n4) );
  MUX2_X1 U609 ( .A(n4), .B(n3), .S(n244), .Z(n5) );
  MUX2_X1 U610 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n251), .Z(n6) );
  MUX2_X1 U611 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n251), .Z(n7) );
  MUX2_X1 U612 ( .A(n7), .B(n6), .S(n246), .Z(n8) );
  MUX2_X1 U613 ( .A(n8), .B(n5), .S(n243), .Z(n9) );
  MUX2_X1 U614 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n251), .Z(n10) );
  MUX2_X1 U615 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n251), .Z(n11) );
  MUX2_X1 U616 ( .A(n11), .B(n10), .S(n245), .Z(n12) );
  MUX2_X1 U617 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n251), .Z(n13) );
  MUX2_X1 U618 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n251), .Z(n14) );
  MUX2_X1 U619 ( .A(n14), .B(n13), .S(n245), .Z(n15) );
  MUX2_X1 U620 ( .A(n15), .B(n12), .S(n243), .Z(n16) );
  MUX2_X1 U621 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U622 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n247), .Z(n18) );
  MUX2_X1 U623 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n247), .Z(n19) );
  MUX2_X1 U624 ( .A(n19), .B(n18), .S(n244), .Z(n20) );
  MUX2_X1 U625 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n247), .Z(n21) );
  MUX2_X1 U626 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n247), .Z(n22) );
  MUX2_X1 U627 ( .A(n22), .B(n21), .S(n244), .Z(n23) );
  MUX2_X1 U628 ( .A(n23), .B(n20), .S(n243), .Z(n24) );
  MUX2_X1 U629 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n247), .Z(n25) );
  MUX2_X1 U630 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n247), .Z(n26) );
  MUX2_X1 U631 ( .A(n26), .B(n25), .S(n244), .Z(n27) );
  MUX2_X1 U632 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n247), .Z(n28) );
  MUX2_X1 U633 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n247), .Z(n29) );
  MUX2_X1 U634 ( .A(n29), .B(n28), .S(n244), .Z(n30) );
  MUX2_X1 U635 ( .A(n30), .B(n27), .S(n243), .Z(n31) );
  MUX2_X1 U636 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U637 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U638 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n247), .Z(n33) );
  MUX2_X1 U639 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n247), .Z(n34) );
  MUX2_X1 U640 ( .A(n34), .B(n33), .S(n244), .Z(n35) );
  MUX2_X1 U641 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n247), .Z(n36) );
  MUX2_X1 U642 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n247), .Z(n37) );
  MUX2_X1 U643 ( .A(n37), .B(n36), .S(n244), .Z(n38) );
  MUX2_X1 U644 ( .A(n38), .B(n35), .S(n243), .Z(n39) );
  MUX2_X1 U645 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n248), .Z(n40) );
  MUX2_X1 U646 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n248), .Z(n41) );
  MUX2_X1 U647 ( .A(n41), .B(n40), .S(n244), .Z(n42) );
  MUX2_X1 U648 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n248), .Z(n43) );
  MUX2_X1 U649 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n248), .Z(n44) );
  MUX2_X1 U650 ( .A(n44), .B(n43), .S(n244), .Z(n45) );
  MUX2_X1 U651 ( .A(n45), .B(n42), .S(N12), .Z(n46) );
  MUX2_X1 U652 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U653 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n248), .Z(n48) );
  MUX2_X1 U654 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n248), .Z(n49) );
  MUX2_X1 U655 ( .A(n49), .B(n48), .S(n244), .Z(n50) );
  MUX2_X1 U656 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n248), .Z(n51) );
  MUX2_X1 U657 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n248), .Z(n52) );
  MUX2_X1 U658 ( .A(n52), .B(n51), .S(n244), .Z(n53) );
  MUX2_X1 U659 ( .A(n53), .B(n50), .S(N12), .Z(n54) );
  MUX2_X1 U660 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n248), .Z(n55) );
  MUX2_X1 U661 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n248), .Z(n56) );
  MUX2_X1 U662 ( .A(n56), .B(n55), .S(n244), .Z(n57) );
  MUX2_X1 U663 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n248), .Z(n58) );
  MUX2_X1 U664 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n248), .Z(n59) );
  MUX2_X1 U665 ( .A(n59), .B(n58), .S(n244), .Z(n60) );
  MUX2_X1 U666 ( .A(n60), .B(n57), .S(N12), .Z(n61) );
  MUX2_X1 U667 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U668 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U669 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n250), .Z(n63) );
  MUX2_X1 U670 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n250), .Z(n64) );
  MUX2_X1 U671 ( .A(n64), .B(n63), .S(n245), .Z(n65) );
  MUX2_X1 U672 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n249), .Z(n66) );
  MUX2_X1 U673 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n247), .Z(n67) );
  MUX2_X1 U674 ( .A(n67), .B(n66), .S(n245), .Z(n68) );
  MUX2_X1 U675 ( .A(n68), .B(n65), .S(n243), .Z(n69) );
  MUX2_X1 U676 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n247), .Z(n70) );
  MUX2_X1 U677 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n249), .Z(n71) );
  MUX2_X1 U678 ( .A(n71), .B(n70), .S(n245), .Z(n72) );
  MUX2_X1 U679 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n247), .Z(n73) );
  MUX2_X1 U680 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n249), .Z(n74) );
  MUX2_X1 U681 ( .A(n74), .B(n73), .S(n245), .Z(n75) );
  MUX2_X1 U682 ( .A(n75), .B(n72), .S(n243), .Z(n76) );
  MUX2_X1 U683 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U684 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n248), .Z(n78) );
  MUX2_X1 U685 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n250), .Z(n79) );
  MUX2_X1 U686 ( .A(n79), .B(n78), .S(n245), .Z(n80) );
  MUX2_X1 U687 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n248), .Z(n81) );
  MUX2_X1 U688 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n250), .Z(n82) );
  MUX2_X1 U689 ( .A(n82), .B(n81), .S(n245), .Z(n83) );
  MUX2_X1 U690 ( .A(n83), .B(n80), .S(n243), .Z(n84) );
  MUX2_X1 U691 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n252), .Z(n85) );
  MUX2_X1 U692 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n249), .Z(n86) );
  MUX2_X1 U693 ( .A(n86), .B(n85), .S(n245), .Z(n87) );
  MUX2_X1 U694 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n248), .Z(n88) );
  MUX2_X1 U695 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n248), .Z(n89) );
  MUX2_X1 U696 ( .A(n89), .B(n88), .S(n245), .Z(n90) );
  MUX2_X1 U697 ( .A(n90), .B(n87), .S(n243), .Z(n91) );
  MUX2_X1 U698 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U699 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U700 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n249), .Z(n93) );
  MUX2_X1 U701 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n252), .Z(n94) );
  MUX2_X1 U702 ( .A(n94), .B(n93), .S(n245), .Z(n95) );
  MUX2_X1 U703 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n252), .Z(n96) );
  MUX2_X1 U704 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n250), .Z(n97) );
  MUX2_X1 U705 ( .A(n97), .B(n96), .S(n245), .Z(n98) );
  MUX2_X1 U706 ( .A(n98), .B(n95), .S(n243), .Z(n99) );
  MUX2_X1 U707 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n252), .Z(n100) );
  MUX2_X1 U708 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n248), .Z(n101) );
  MUX2_X1 U709 ( .A(n101), .B(n100), .S(n245), .Z(n102) );
  MUX2_X1 U710 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n252), .Z(n103) );
  MUX2_X1 U711 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n247), .Z(n104) );
  MUX2_X1 U712 ( .A(n104), .B(n103), .S(n245), .Z(n105) );
  MUX2_X1 U713 ( .A(n105), .B(n102), .S(n243), .Z(n106) );
  MUX2_X1 U714 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U715 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n249), .Z(n108) );
  MUX2_X1 U716 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n249), .Z(n109) );
  MUX2_X1 U717 ( .A(n109), .B(n108), .S(n246), .Z(n110) );
  MUX2_X1 U718 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n249), .Z(n111) );
  MUX2_X1 U719 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n249), .Z(n112) );
  MUX2_X1 U720 ( .A(n112), .B(n111), .S(n246), .Z(n113) );
  MUX2_X1 U721 ( .A(n113), .B(n110), .S(n243), .Z(n114) );
  MUX2_X1 U722 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n249), .Z(n115) );
  MUX2_X1 U723 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n249), .Z(n116) );
  MUX2_X1 U724 ( .A(n116), .B(n115), .S(n246), .Z(n117) );
  MUX2_X1 U725 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n249), .Z(n118) );
  MUX2_X1 U726 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n249), .Z(n119) );
  MUX2_X1 U727 ( .A(n119), .B(n118), .S(n246), .Z(n120) );
  MUX2_X1 U728 ( .A(n120), .B(n117), .S(n243), .Z(n121) );
  MUX2_X1 U729 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U730 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U731 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n249), .Z(n123) );
  MUX2_X1 U732 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n249), .Z(n124) );
  MUX2_X1 U733 ( .A(n124), .B(n123), .S(n246), .Z(n125) );
  MUX2_X1 U734 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n249), .Z(n126) );
  MUX2_X1 U735 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n249), .Z(n127) );
  MUX2_X1 U736 ( .A(n127), .B(n126), .S(n246), .Z(n128) );
  MUX2_X1 U737 ( .A(n128), .B(n125), .S(n243), .Z(n129) );
  MUX2_X1 U738 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n250), .Z(n130) );
  MUX2_X1 U739 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n250), .Z(n131) );
  MUX2_X1 U740 ( .A(n131), .B(n130), .S(n246), .Z(n132) );
  MUX2_X1 U741 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n250), .Z(n133) );
  MUX2_X1 U742 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n250), .Z(n134) );
  MUX2_X1 U743 ( .A(n134), .B(n133), .S(n246), .Z(n135) );
  MUX2_X1 U744 ( .A(n135), .B(n132), .S(n243), .Z(n136) );
  MUX2_X1 U745 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U746 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n250), .Z(n138) );
  MUX2_X1 U747 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n250), .Z(n139) );
  MUX2_X1 U748 ( .A(n139), .B(n138), .S(n246), .Z(n140) );
  MUX2_X1 U749 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n250), .Z(n141) );
  MUX2_X1 U750 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n250), .Z(n142) );
  MUX2_X1 U751 ( .A(n142), .B(n141), .S(n246), .Z(n143) );
  MUX2_X1 U752 ( .A(n143), .B(n140), .S(n243), .Z(n144) );
  MUX2_X1 U753 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n250), .Z(n145) );
  MUX2_X1 U754 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n250), .Z(n146) );
  MUX2_X1 U755 ( .A(n146), .B(n145), .S(n246), .Z(n147) );
  MUX2_X1 U756 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n250), .Z(n148) );
  MUX2_X1 U757 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n250), .Z(n149) );
  MUX2_X1 U758 ( .A(n149), .B(n148), .S(n246), .Z(n150) );
  MUX2_X1 U759 ( .A(n150), .B(n147), .S(n243), .Z(n151) );
  MUX2_X1 U760 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U761 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U762 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n251), .Z(n153) );
  MUX2_X1 U763 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n251), .Z(n154) );
  MUX2_X1 U764 ( .A(n154), .B(n153), .S(N11), .Z(n155) );
  MUX2_X1 U765 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n251), .Z(n156) );
  MUX2_X1 U766 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n251), .Z(n157) );
  MUX2_X1 U767 ( .A(n157), .B(n156), .S(N11), .Z(n158) );
  MUX2_X1 U768 ( .A(n158), .B(n155), .S(n243), .Z(n159) );
  MUX2_X1 U769 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n251), .Z(n160) );
  MUX2_X1 U770 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n251), .Z(n161) );
  MUX2_X1 U771 ( .A(n161), .B(n160), .S(N11), .Z(n162) );
  MUX2_X1 U772 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n251), .Z(n163) );
  MUX2_X1 U773 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n251), .Z(n164) );
  MUX2_X1 U774 ( .A(n164), .B(n163), .S(n246), .Z(n165) );
  MUX2_X1 U775 ( .A(n165), .B(n162), .S(N12), .Z(n166) );
  MUX2_X1 U776 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U777 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n251), .Z(n168) );
  MUX2_X1 U778 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n251), .Z(n169) );
  MUX2_X1 U779 ( .A(n169), .B(n168), .S(N11), .Z(n170) );
  MUX2_X1 U780 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n251), .Z(n171) );
  MUX2_X1 U781 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n251), .Z(n172) );
  MUX2_X1 U782 ( .A(n172), .B(n171), .S(n244), .Z(n173) );
  MUX2_X1 U783 ( .A(n173), .B(n170), .S(n243), .Z(n174) );
  MUX2_X1 U784 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n248), .Z(n175) );
  MUX2_X1 U785 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n252), .Z(n176) );
  MUX2_X1 U786 ( .A(n176), .B(n175), .S(N11), .Z(n177) );
  MUX2_X1 U787 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n252), .Z(n178) );
  MUX2_X1 U788 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n252), .Z(n179) );
  MUX2_X1 U789 ( .A(n179), .B(n178), .S(n246), .Z(n180) );
  MUX2_X1 U790 ( .A(n180), .B(n177), .S(N12), .Z(n181) );
  MUX2_X1 U791 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U792 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U793 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n247), .Z(n183) );
  MUX2_X1 U794 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n252), .Z(n184) );
  MUX2_X1 U795 ( .A(n184), .B(n183), .S(N11), .Z(n185) );
  MUX2_X1 U796 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n252), .Z(n186) );
  MUX2_X1 U797 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n250), .Z(n187) );
  MUX2_X1 U798 ( .A(n187), .B(n186), .S(N11), .Z(n188) );
  MUX2_X1 U799 ( .A(n188), .B(n185), .S(n243), .Z(n189) );
  MUX2_X1 U800 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n252), .Z(n190) );
  MUX2_X1 U801 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n252), .Z(n191) );
  MUX2_X1 U802 ( .A(n191), .B(n190), .S(N11), .Z(n192) );
  MUX2_X1 U803 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n252), .Z(n193) );
  MUX2_X1 U804 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n252), .Z(n194) );
  MUX2_X1 U805 ( .A(n194), .B(n193), .S(n244), .Z(n195) );
  MUX2_X1 U806 ( .A(n195), .B(n192), .S(N12), .Z(n196) );
  MUX2_X1 U807 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U808 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n252), .Z(n198) );
  MUX2_X1 U809 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(N10), .Z(n199) );
  MUX2_X1 U810 ( .A(n199), .B(n198), .S(n245), .Z(n200) );
  MUX2_X1 U811 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(N10), .Z(n201) );
  MUX2_X1 U812 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n202) );
  MUX2_X1 U813 ( .A(n202), .B(n201), .S(n245), .Z(n203) );
  MUX2_X1 U814 ( .A(n203), .B(n200), .S(n243), .Z(n204) );
  MUX2_X1 U815 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n252), .Z(n205) );
  MUX2_X1 U816 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n252), .Z(n206) );
  MUX2_X1 U817 ( .A(n206), .B(n205), .S(n245), .Z(n207) );
  MUX2_X1 U818 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n208) );
  MUX2_X1 U819 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n252), .Z(n209) );
  MUX2_X1 U820 ( .A(n209), .B(n208), .S(N11), .Z(n210) );
  MUX2_X1 U821 ( .A(n210), .B(n207), .S(N12), .Z(n211) );
  MUX2_X1 U822 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U823 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U824 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n249), .Z(n213) );
  MUX2_X1 U825 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(N10), .Z(n214) );
  MUX2_X1 U826 ( .A(n214), .B(n213), .S(n244), .Z(n215) );
  MUX2_X1 U827 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(N10), .Z(n216) );
  MUX2_X1 U828 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(N10), .Z(n217) );
  MUX2_X1 U829 ( .A(n217), .B(n216), .S(n244), .Z(n218) );
  MUX2_X1 U830 ( .A(n218), .B(n215), .S(n243), .Z(n219) );
  MUX2_X1 U831 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n251), .Z(n220) );
  MUX2_X1 U832 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(N10), .Z(n221) );
  MUX2_X1 U833 ( .A(n221), .B(n220), .S(N11), .Z(n222) );
  MUX2_X1 U834 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n252), .Z(n223) );
  MUX2_X1 U835 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n224) );
  MUX2_X1 U836 ( .A(n224), .B(n223), .S(N11), .Z(n225) );
  MUX2_X1 U837 ( .A(n225), .B(n222), .S(N12), .Z(n226) );
  MUX2_X1 U838 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U839 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n251), .Z(n228) );
  MUX2_X1 U840 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n252), .Z(n229) );
  MUX2_X1 U841 ( .A(n229), .B(n228), .S(n246), .Z(n230) );
  MUX2_X1 U842 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n251), .Z(n231) );
  MUX2_X1 U843 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n232) );
  MUX2_X1 U844 ( .A(n232), .B(n231), .S(N11), .Z(n233) );
  MUX2_X1 U845 ( .A(n233), .B(n230), .S(n243), .Z(n234) );
  MUX2_X1 U846 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n235) );
  MUX2_X1 U847 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n236) );
  MUX2_X1 U848 ( .A(n236), .B(n235), .S(n246), .Z(n237) );
  MUX2_X1 U849 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n238) );
  MUX2_X1 U850 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n239) );
  MUX2_X1 U851 ( .A(n239), .B(n238), .S(N11), .Z(n240) );
  MUX2_X1 U852 ( .A(n240), .B(n237), .S(N12), .Z(n241) );
  MUX2_X1 U853 ( .A(n241), .B(n234), .S(N13), .Z(n242) );
  MUX2_X1 U854 ( .A(n242), .B(n227), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_29 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  BUF_X1 U3 ( .A(n250), .Z(n248) );
  BUF_X1 U4 ( .A(N10), .Z(n249) );
  BUF_X1 U5 ( .A(n250), .Z(n245) );
  BUF_X1 U6 ( .A(n250), .Z(n246) );
  BUF_X1 U7 ( .A(n250), .Z(n247) );
  BUF_X1 U8 ( .A(N10), .Z(n250) );
  INV_X1 U9 ( .A(n1111), .ZN(n841) );
  INV_X1 U10 ( .A(n1100), .ZN(n840) );
  INV_X1 U11 ( .A(n1090), .ZN(n839) );
  INV_X1 U12 ( .A(n1080), .ZN(n838) );
  INV_X1 U13 ( .A(n1070), .ZN(n837) );
  INV_X1 U14 ( .A(n1060), .ZN(n836) );
  INV_X1 U15 ( .A(n1051), .ZN(n835) );
  INV_X1 U16 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U19 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U20 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U21 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U22 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U23 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U24 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U26 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U27 ( .A(n1131), .ZN(n816) );
  INV_X1 U28 ( .A(n1121), .ZN(n815) );
  INV_X1 U29 ( .A(n887), .ZN(n814) );
  INV_X1 U30 ( .A(n878), .ZN(n813) );
  INV_X1 U31 ( .A(n869), .ZN(n812) );
  INV_X1 U32 ( .A(n860), .ZN(n811) );
  INV_X1 U33 ( .A(n851), .ZN(n810) );
  INV_X1 U34 ( .A(n987), .ZN(n828) );
  INV_X1 U35 ( .A(n978), .ZN(n827) );
  INV_X1 U36 ( .A(n969), .ZN(n826) );
  INV_X1 U37 ( .A(n914), .ZN(n820) );
  INV_X1 U38 ( .A(n905), .ZN(n819) );
  INV_X1 U39 ( .A(n896), .ZN(n818) );
  INV_X1 U40 ( .A(n1033), .ZN(n833) );
  INV_X1 U41 ( .A(n1023), .ZN(n832) );
  INV_X1 U42 ( .A(n1014), .ZN(n831) );
  INV_X1 U43 ( .A(n1005), .ZN(n830) );
  INV_X1 U44 ( .A(n996), .ZN(n829) );
  INV_X1 U45 ( .A(n960), .ZN(n825) );
  INV_X1 U46 ( .A(n950), .ZN(n824) );
  INV_X1 U47 ( .A(n941), .ZN(n823) );
  INV_X1 U48 ( .A(n932), .ZN(n822) );
  INV_X1 U49 ( .A(n923), .ZN(n821) );
  INV_X1 U50 ( .A(n1142), .ZN(n817) );
  BUF_X1 U51 ( .A(N11), .Z(n242) );
  BUF_X1 U52 ( .A(N11), .Z(n243) );
  BUF_X1 U53 ( .A(N11), .Z(n244) );
  INV_X1 U54 ( .A(N10), .ZN(n251) );
  BUF_X1 U55 ( .A(N12), .Z(n241) );
  NOR3_X1 U56 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U57 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U58 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U60 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U62 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U63 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U64 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U65 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U67 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U69 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U70 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U71 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U72 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U73 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U74 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U75 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U76 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U77 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U79 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U81 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U82 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U83 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U84 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U85 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U86 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U88 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U89 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U90 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U92 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U94 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U95 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U96 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U97 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U98 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U99 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U100 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U101 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U102 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U103 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U104 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U105 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U106 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U107 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U108 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U109 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U110 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U111 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U112 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U113 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U114 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U115 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U116 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U117 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U118 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U119 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U120 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U121 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U122 ( .A(n988), .ZN(n705) );
  AOI22_X1 U123 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U124 ( .A(n986), .ZN(n704) );
  AOI22_X1 U125 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U126 ( .A(n985), .ZN(n703) );
  AOI22_X1 U127 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U128 ( .A(n984), .ZN(n702) );
  AOI22_X1 U129 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U130 ( .A(n983), .ZN(n701) );
  AOI22_X1 U131 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U132 ( .A(n982), .ZN(n700) );
  AOI22_X1 U133 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U134 ( .A(n981), .ZN(n699) );
  AOI22_X1 U135 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U136 ( .A(n980), .ZN(n698) );
  AOI22_X1 U137 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U138 ( .A(n951), .ZN(n673) );
  AOI22_X1 U139 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U140 ( .A(n949), .ZN(n672) );
  AOI22_X1 U141 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U142 ( .A(n948), .ZN(n671) );
  AOI22_X1 U143 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U144 ( .A(n947), .ZN(n670) );
  AOI22_X1 U145 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U146 ( .A(n946), .ZN(n669) );
  AOI22_X1 U147 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U148 ( .A(n945), .ZN(n668) );
  AOI22_X1 U149 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U150 ( .A(n944), .ZN(n667) );
  AOI22_X1 U151 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U152 ( .A(n943), .ZN(n666) );
  AOI22_X1 U153 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U154 ( .A(n915), .ZN(n641) );
  AOI22_X1 U155 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U156 ( .A(n913), .ZN(n640) );
  AOI22_X1 U157 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U158 ( .A(n912), .ZN(n639) );
  AOI22_X1 U159 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U160 ( .A(n911), .ZN(n638) );
  AOI22_X1 U161 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U162 ( .A(n910), .ZN(n637) );
  AOI22_X1 U163 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U164 ( .A(n909), .ZN(n636) );
  AOI22_X1 U165 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U166 ( .A(n908), .ZN(n635) );
  AOI22_X1 U167 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U168 ( .A(n907), .ZN(n634) );
  AOI22_X1 U169 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U170 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U171 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U172 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U173 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U174 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U175 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U176 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U177 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U178 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U179 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U180 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U181 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U182 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U183 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U184 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U185 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U186 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U187 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U188 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U189 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U190 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U191 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U192 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U193 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U194 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U195 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U196 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U197 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U198 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U199 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U200 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U201 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U202 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U203 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U204 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U205 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U206 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U207 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U208 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U209 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U210 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U211 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U212 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U213 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U214 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U215 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U216 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U217 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U218 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U219 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U220 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U221 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U222 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U223 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U224 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U225 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U226 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U227 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U228 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U229 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U230 ( .A(n999), .ZN(n715) );
  AOI22_X1 U231 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U232 ( .A(n998), .ZN(n714) );
  AOI22_X1 U233 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U234 ( .A(n942), .ZN(n665) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U236 ( .A(n940), .ZN(n664) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U238 ( .A(n939), .ZN(n663) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U240 ( .A(n938), .ZN(n662) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U242 ( .A(n937), .ZN(n661) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U244 ( .A(n936), .ZN(n660) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U246 ( .A(n935), .ZN(n659) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U248 ( .A(n934), .ZN(n658) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U250 ( .A(n933), .ZN(n657) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U252 ( .A(n931), .ZN(n656) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U254 ( .A(n930), .ZN(n655) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U256 ( .A(n929), .ZN(n654) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U258 ( .A(n928), .ZN(n653) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U260 ( .A(n927), .ZN(n652) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U262 ( .A(n926), .ZN(n651) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U264 ( .A(n925), .ZN(n650) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U266 ( .A(n979), .ZN(n697) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U268 ( .A(n977), .ZN(n696) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U270 ( .A(n976), .ZN(n695) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U272 ( .A(n975), .ZN(n694) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U274 ( .A(n974), .ZN(n693) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U276 ( .A(n973), .ZN(n692) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U278 ( .A(n972), .ZN(n691) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U280 ( .A(n971), .ZN(n690) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U282 ( .A(n970), .ZN(n689) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U284 ( .A(n968), .ZN(n688) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U286 ( .A(n967), .ZN(n687) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U288 ( .A(n966), .ZN(n686) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U290 ( .A(n965), .ZN(n685) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U292 ( .A(n964), .ZN(n684) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U294 ( .A(n963), .ZN(n683) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U296 ( .A(n962), .ZN(n682) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U298 ( .A(n906), .ZN(n633) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U300 ( .A(n904), .ZN(n632) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U302 ( .A(n903), .ZN(n631) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U304 ( .A(n902), .ZN(n630) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U306 ( .A(n901), .ZN(n629) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U308 ( .A(n900), .ZN(n628) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U310 ( .A(n899), .ZN(n627) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U312 ( .A(n898), .ZN(n626) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U314 ( .A(n897), .ZN(n625) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U316 ( .A(n895), .ZN(n624) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U318 ( .A(n894), .ZN(n623) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U320 ( .A(n893), .ZN(n622) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U322 ( .A(n892), .ZN(n621) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U324 ( .A(n891), .ZN(n620) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U326 ( .A(n890), .ZN(n619) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U328 ( .A(n889), .ZN(n618) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U330 ( .A(N12), .ZN(n253) );
  INV_X1 U331 ( .A(N11), .ZN(n252) );
  INV_X1 U332 ( .A(n997), .ZN(n713) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U334 ( .A(n995), .ZN(n712) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U336 ( .A(n994), .ZN(n711) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U338 ( .A(n993), .ZN(n710) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U340 ( .A(n992), .ZN(n709) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U342 ( .A(n991), .ZN(n708) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U344 ( .A(n990), .ZN(n707) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U346 ( .A(n989), .ZN(n706) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U348 ( .A(n924), .ZN(n649) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U350 ( .A(n922), .ZN(n648) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U352 ( .A(n921), .ZN(n647) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U354 ( .A(n920), .ZN(n646) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U356 ( .A(n919), .ZN(n645) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U358 ( .A(n918), .ZN(n644) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U360 ( .A(n917), .ZN(n643) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U362 ( .A(n916), .ZN(n642) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U364 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U366 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U368 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U370 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U372 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U374 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U376 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U378 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U380 ( .A(n961), .ZN(n681) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U382 ( .A(n959), .ZN(n680) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U384 ( .A(n958), .ZN(n679) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U386 ( .A(n957), .ZN(n678) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U388 ( .A(n956), .ZN(n677) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U390 ( .A(n955), .ZN(n676) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U392 ( .A(n954), .ZN(n675) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U394 ( .A(n953), .ZN(n674) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U396 ( .A(n888), .ZN(n617) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U398 ( .A(n886), .ZN(n616) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U400 ( .A(n885), .ZN(n615) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U402 ( .A(n884), .ZN(n614) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U404 ( .A(n883), .ZN(n613) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U406 ( .A(n882), .ZN(n612) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U408 ( .A(n881), .ZN(n611) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U410 ( .A(n880), .ZN(n610) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U412 ( .A(n879), .ZN(n609) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U414 ( .A(n877), .ZN(n608) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U416 ( .A(n876), .ZN(n607) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U418 ( .A(n875), .ZN(n606) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U420 ( .A(n874), .ZN(n605) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U422 ( .A(n873), .ZN(n604) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U424 ( .A(n872), .ZN(n603) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U426 ( .A(n871), .ZN(n602) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U428 ( .A(n870), .ZN(n601) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U430 ( .A(n868), .ZN(n600) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U432 ( .A(n867), .ZN(n599) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U434 ( .A(n866), .ZN(n598) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U436 ( .A(n865), .ZN(n597) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U438 ( .A(n864), .ZN(n596) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U440 ( .A(n863), .ZN(n595) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U442 ( .A(n862), .ZN(n594) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U444 ( .A(n861), .ZN(n293) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U446 ( .A(n859), .ZN(n292) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U448 ( .A(n858), .ZN(n291) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U450 ( .A(n857), .ZN(n290) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U452 ( .A(n856), .ZN(n289) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U454 ( .A(n855), .ZN(n288) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U456 ( .A(n854), .ZN(n287) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U458 ( .A(n853), .ZN(n286) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U460 ( .A(n852), .ZN(n285) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U462 ( .A(n850), .ZN(n284) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U464 ( .A(n849), .ZN(n283) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U466 ( .A(n848), .ZN(n282) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U468 ( .A(n847), .ZN(n281) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U470 ( .A(n846), .ZN(n280) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U472 ( .A(n845), .ZN(n279) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U474 ( .A(n844), .ZN(n278) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U476 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U477 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U478 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U479 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U480 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U481 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U482 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U483 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U484 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U485 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U486 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U487 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U488 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U489 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U490 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U491 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U492 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U494 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U496 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U498 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U500 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U502 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U504 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U506 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U508 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U510 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U512 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U514 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U516 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U518 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U520 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U522 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U524 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U526 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U528 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U530 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U532 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U534 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U536 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U538 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U540 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U542 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U544 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U546 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U548 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U550 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U552 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U554 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U556 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U558 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U560 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U562 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U564 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U566 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U568 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U570 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U572 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U574 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U576 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U578 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U580 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U582 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U584 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U586 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U588 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U590 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U592 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U594 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U596 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U598 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U600 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U602 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U604 ( .A(N13), .ZN(n842) );
  INV_X1 U605 ( .A(N14), .ZN(n843) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n249), .Z(n1) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n249), .Z(n2) );
  MUX2_X1 U608 ( .A(n2), .B(n1), .S(n242), .Z(n3) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n249), .Z(n4) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n248), .Z(n5) );
  MUX2_X1 U611 ( .A(n5), .B(n4), .S(n242), .Z(n6) );
  MUX2_X1 U612 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n249), .Z(n8) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n249), .Z(n9) );
  MUX2_X1 U615 ( .A(n9), .B(n8), .S(N11), .Z(n10) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n249), .Z(n11) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n248), .Z(n12) );
  MUX2_X1 U618 ( .A(n12), .B(n11), .S(n244), .Z(n13) );
  MUX2_X1 U619 ( .A(n13), .B(n10), .S(n241), .Z(n14) );
  MUX2_X1 U620 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n245), .Z(n16) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n245), .Z(n17) );
  MUX2_X1 U623 ( .A(n17), .B(n16), .S(n242), .Z(n18) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n245), .Z(n20) );
  MUX2_X1 U626 ( .A(n20), .B(n19), .S(n242), .Z(n21) );
  MUX2_X1 U627 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n245), .Z(n23) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n245), .Z(n24) );
  MUX2_X1 U630 ( .A(n24), .B(n23), .S(n242), .Z(n25) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n245), .Z(n26) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n245), .Z(n27) );
  MUX2_X1 U633 ( .A(n27), .B(n26), .S(n242), .Z(n28) );
  MUX2_X1 U634 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U635 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U636 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n245), .Z(n31) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n245), .Z(n32) );
  MUX2_X1 U639 ( .A(n32), .B(n31), .S(n242), .Z(n33) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U642 ( .A(n35), .B(n34), .S(n242), .Z(n36) );
  MUX2_X1 U643 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n246), .Z(n38) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n246), .Z(n39) );
  MUX2_X1 U646 ( .A(n39), .B(n38), .S(n242), .Z(n40) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n246), .Z(n41) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n246), .Z(n42) );
  MUX2_X1 U649 ( .A(n42), .B(n41), .S(n242), .Z(n43) );
  MUX2_X1 U650 ( .A(n43), .B(n40), .S(n241), .Z(n44) );
  MUX2_X1 U651 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n246), .Z(n46) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n246), .Z(n47) );
  MUX2_X1 U654 ( .A(n47), .B(n46), .S(n242), .Z(n48) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n246), .Z(n49) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n246), .Z(n50) );
  MUX2_X1 U657 ( .A(n50), .B(n49), .S(n242), .Z(n51) );
  MUX2_X1 U658 ( .A(n51), .B(n48), .S(n241), .Z(n52) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n246), .Z(n53) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n246), .Z(n54) );
  MUX2_X1 U661 ( .A(n54), .B(n53), .S(n242), .Z(n55) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n246), .Z(n56) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n246), .Z(n57) );
  MUX2_X1 U664 ( .A(n57), .B(n56), .S(n242), .Z(n58) );
  MUX2_X1 U665 ( .A(n58), .B(n55), .S(n241), .Z(n59) );
  MUX2_X1 U666 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U667 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n247), .Z(n61) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n247), .Z(n62) );
  MUX2_X1 U670 ( .A(n62), .B(n61), .S(n243), .Z(n63) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n247), .Z(n64) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n247), .Z(n65) );
  MUX2_X1 U673 ( .A(n65), .B(n64), .S(n243), .Z(n66) );
  MUX2_X1 U674 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n247), .Z(n68) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n247), .Z(n69) );
  MUX2_X1 U677 ( .A(n69), .B(n68), .S(n243), .Z(n70) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n247), .Z(n71) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n247), .Z(n72) );
  MUX2_X1 U680 ( .A(n72), .B(n71), .S(n243), .Z(n73) );
  MUX2_X1 U681 ( .A(n73), .B(n70), .S(N12), .Z(n74) );
  MUX2_X1 U682 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n247), .Z(n76) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n247), .Z(n77) );
  MUX2_X1 U685 ( .A(n77), .B(n76), .S(n243), .Z(n78) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n247), .Z(n79) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n247), .Z(n80) );
  MUX2_X1 U688 ( .A(n80), .B(n79), .S(n243), .Z(n81) );
  MUX2_X1 U689 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n248), .Z(n83) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n247), .Z(n84) );
  MUX2_X1 U692 ( .A(n84), .B(n83), .S(n243), .Z(n85) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n246), .Z(n86) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n245), .Z(n87) );
  MUX2_X1 U695 ( .A(n87), .B(n86), .S(n243), .Z(n88) );
  MUX2_X1 U696 ( .A(n88), .B(n85), .S(N12), .Z(n89) );
  MUX2_X1 U697 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U698 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n248), .Z(n91) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n247), .Z(n92) );
  MUX2_X1 U701 ( .A(n92), .B(n91), .S(n243), .Z(n93) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n248), .Z(n95) );
  MUX2_X1 U704 ( .A(n95), .B(n94), .S(n243), .Z(n96) );
  MUX2_X1 U705 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n245), .Z(n98) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n245), .Z(n99) );
  MUX2_X1 U708 ( .A(n99), .B(n98), .S(n243), .Z(n100) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n246), .Z(n101) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n246), .Z(n102) );
  MUX2_X1 U711 ( .A(n102), .B(n101), .S(n243), .Z(n103) );
  MUX2_X1 U712 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U713 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n249), .Z(n106) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(N10), .Z(n107) );
  MUX2_X1 U716 ( .A(n107), .B(n106), .S(n244), .Z(n108) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n249), .Z(n109) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n110) );
  MUX2_X1 U719 ( .A(n110), .B(n109), .S(n244), .Z(n111) );
  MUX2_X1 U720 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n249), .Z(n113) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n250), .Z(n114) );
  MUX2_X1 U723 ( .A(n114), .B(n113), .S(n244), .Z(n115) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n249), .Z(n116) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n117) );
  MUX2_X1 U726 ( .A(n117), .B(n116), .S(n244), .Z(n118) );
  MUX2_X1 U727 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U728 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U729 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(N10), .Z(n121) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(N10), .Z(n122) );
  MUX2_X1 U732 ( .A(n122), .B(n121), .S(n244), .Z(n123) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(N10), .Z(n124) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n125) );
  MUX2_X1 U735 ( .A(n125), .B(n124), .S(n244), .Z(n126) );
  MUX2_X1 U736 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n248), .Z(n128) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n248), .Z(n129) );
  MUX2_X1 U739 ( .A(n129), .B(n128), .S(n244), .Z(n130) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n248), .Z(n131) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n248), .Z(n132) );
  MUX2_X1 U742 ( .A(n132), .B(n131), .S(n244), .Z(n133) );
  MUX2_X1 U743 ( .A(n133), .B(n130), .S(N12), .Z(n134) );
  MUX2_X1 U744 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n248), .Z(n136) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n248), .Z(n137) );
  MUX2_X1 U747 ( .A(n137), .B(n136), .S(n244), .Z(n138) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n248), .Z(n139) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n248), .Z(n140) );
  MUX2_X1 U750 ( .A(n140), .B(n139), .S(n244), .Z(n141) );
  MUX2_X1 U751 ( .A(n141), .B(n138), .S(N12), .Z(n142) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n248), .Z(n143) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n248), .Z(n144) );
  MUX2_X1 U754 ( .A(n144), .B(n143), .S(n244), .Z(n145) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n248), .Z(n146) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n248), .Z(n147) );
  MUX2_X1 U757 ( .A(n147), .B(n146), .S(n244), .Z(n148) );
  MUX2_X1 U758 ( .A(n148), .B(n145), .S(N12), .Z(n149) );
  MUX2_X1 U759 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U760 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n249), .Z(n151) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n249), .Z(n152) );
  MUX2_X1 U763 ( .A(n152), .B(n151), .S(n242), .Z(n153) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n249), .Z(n154) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n249), .Z(n155) );
  MUX2_X1 U766 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U767 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n249), .Z(n158) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n249), .Z(n159) );
  MUX2_X1 U770 ( .A(n159), .B(n158), .S(N11), .Z(n160) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n249), .Z(n161) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n249), .Z(n162) );
  MUX2_X1 U773 ( .A(n162), .B(n161), .S(n242), .Z(n163) );
  MUX2_X1 U774 ( .A(n163), .B(n160), .S(n241), .Z(n164) );
  MUX2_X1 U775 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n249), .Z(n166) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n249), .Z(n167) );
  MUX2_X1 U778 ( .A(n167), .B(n166), .S(N11), .Z(n168) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n249), .Z(n169) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n249), .Z(n170) );
  MUX2_X1 U781 ( .A(n170), .B(n169), .S(n243), .Z(n171) );
  MUX2_X1 U782 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n245), .Z(n173) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n250), .Z(n174) );
  MUX2_X1 U785 ( .A(n174), .B(n173), .S(N11), .Z(n175) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n247), .Z(n176) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n246), .Z(n177) );
  MUX2_X1 U788 ( .A(n177), .B(n176), .S(n243), .Z(n178) );
  MUX2_X1 U789 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U790 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U791 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n250), .Z(n181) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n245), .Z(n182) );
  MUX2_X1 U794 ( .A(n182), .B(n181), .S(N11), .Z(n183) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n250), .Z(n184) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n246), .Z(n185) );
  MUX2_X1 U797 ( .A(n185), .B(n184), .S(N11), .Z(n186) );
  MUX2_X1 U798 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n247), .Z(n188) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n250), .Z(n189) );
  MUX2_X1 U801 ( .A(n189), .B(n188), .S(N11), .Z(n190) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n250), .Z(n191) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n250), .Z(n192) );
  MUX2_X1 U804 ( .A(n192), .B(n191), .S(n244), .Z(n193) );
  MUX2_X1 U805 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U806 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n250), .Z(n196) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n250), .Z(n197) );
  MUX2_X1 U809 ( .A(n197), .B(n196), .S(n242), .Z(n198) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n250), .Z(n199) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n250), .Z(n200) );
  MUX2_X1 U812 ( .A(n200), .B(n199), .S(n244), .Z(n201) );
  MUX2_X1 U813 ( .A(n201), .B(n198), .S(n241), .Z(n202) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n250), .Z(n203) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n250), .Z(n204) );
  MUX2_X1 U816 ( .A(n204), .B(n203), .S(n244), .Z(n205) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n250), .Z(n206) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n250), .Z(n207) );
  MUX2_X1 U819 ( .A(n207), .B(n206), .S(N11), .Z(n208) );
  MUX2_X1 U820 ( .A(n208), .B(n205), .S(n241), .Z(n209) );
  MUX2_X1 U821 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U822 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n250), .Z(n211) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n247), .Z(n212) );
  MUX2_X1 U825 ( .A(n212), .B(n211), .S(n243), .Z(n213) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n249), .Z(n214) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n250), .Z(n215) );
  MUX2_X1 U828 ( .A(n215), .B(n214), .S(n244), .Z(n216) );
  MUX2_X1 U829 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n245), .Z(n218) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(N10), .Z(n219) );
  MUX2_X1 U832 ( .A(n219), .B(n218), .S(n243), .Z(n220) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n250), .Z(n221) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n246), .Z(n222) );
  MUX2_X1 U835 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U836 ( .A(n223), .B(n220), .S(n241), .Z(n224) );
  MUX2_X1 U837 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n247), .Z(n226) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n227) );
  MUX2_X1 U840 ( .A(n227), .B(n226), .S(N11), .Z(n228) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n250), .Z(n229) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n230) );
  MUX2_X1 U843 ( .A(n230), .B(n229), .S(N11), .Z(n231) );
  MUX2_X1 U844 ( .A(n231), .B(n228), .S(N12), .Z(n232) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n233) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n234) );
  MUX2_X1 U847 ( .A(n234), .B(n233), .S(n243), .Z(n235) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n236) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n237) );
  MUX2_X1 U850 ( .A(n237), .B(n236), .S(N11), .Z(n238) );
  MUX2_X1 U851 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U852 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U853 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_28 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X2 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(n250), .Z(n247) );
  BUF_X1 U4 ( .A(N10), .Z(n248) );
  BUF_X1 U5 ( .A(n250), .Z(n249) );
  BUF_X1 U6 ( .A(n250), .Z(n246) );
  BUF_X1 U7 ( .A(n250), .Z(n245) );
  BUF_X1 U8 ( .A(N10), .Z(n250) );
  INV_X1 U9 ( .A(n1111), .ZN(n841) );
  INV_X1 U10 ( .A(n1100), .ZN(n840) );
  INV_X1 U11 ( .A(n1090), .ZN(n839) );
  INV_X1 U12 ( .A(n1080), .ZN(n838) );
  INV_X1 U13 ( .A(n1070), .ZN(n837) );
  INV_X1 U14 ( .A(n1060), .ZN(n836) );
  INV_X1 U15 ( .A(n1051), .ZN(n835) );
  INV_X1 U16 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U19 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U20 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U21 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U22 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U23 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U24 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U26 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U27 ( .A(n1131), .ZN(n816) );
  INV_X1 U28 ( .A(n1121), .ZN(n815) );
  INV_X1 U29 ( .A(n887), .ZN(n814) );
  INV_X1 U30 ( .A(n878), .ZN(n813) );
  INV_X1 U31 ( .A(n869), .ZN(n812) );
  INV_X1 U32 ( .A(n860), .ZN(n811) );
  INV_X1 U33 ( .A(n851), .ZN(n810) );
  INV_X1 U34 ( .A(n987), .ZN(n828) );
  INV_X1 U35 ( .A(n978), .ZN(n827) );
  INV_X1 U36 ( .A(n969), .ZN(n826) );
  INV_X1 U37 ( .A(n914), .ZN(n820) );
  INV_X1 U38 ( .A(n905), .ZN(n819) );
  INV_X1 U39 ( .A(n896), .ZN(n818) );
  INV_X1 U40 ( .A(n1033), .ZN(n833) );
  INV_X1 U41 ( .A(n1023), .ZN(n832) );
  INV_X1 U42 ( .A(n1014), .ZN(n831) );
  INV_X1 U43 ( .A(n1005), .ZN(n830) );
  INV_X1 U44 ( .A(n996), .ZN(n829) );
  INV_X1 U45 ( .A(n960), .ZN(n825) );
  INV_X1 U46 ( .A(n950), .ZN(n824) );
  INV_X1 U47 ( .A(n941), .ZN(n823) );
  INV_X1 U48 ( .A(n932), .ZN(n822) );
  INV_X1 U49 ( .A(n923), .ZN(n821) );
  INV_X1 U50 ( .A(n1142), .ZN(n817) );
  BUF_X1 U51 ( .A(N11), .Z(n242) );
  BUF_X1 U52 ( .A(N11), .Z(n243) );
  BUF_X1 U53 ( .A(N11), .Z(n244) );
  INV_X1 U54 ( .A(N10), .ZN(n251) );
  BUF_X1 U55 ( .A(N12), .Z(n241) );
  NOR3_X1 U56 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U57 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U58 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U60 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U62 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U63 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U64 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U65 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U67 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U69 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U70 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U71 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U72 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U73 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U74 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U75 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U76 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U77 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U79 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U81 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U82 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U83 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U84 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U85 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U86 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U88 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U89 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U90 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U92 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U94 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U95 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U96 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U97 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U98 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U99 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U100 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U101 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U102 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U103 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U104 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U105 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U106 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U107 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U108 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U109 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U110 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U111 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U112 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U113 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U114 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U115 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U116 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U117 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U118 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U119 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U120 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U121 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U122 ( .A(n988), .ZN(n705) );
  AOI22_X1 U123 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U124 ( .A(n986), .ZN(n704) );
  AOI22_X1 U125 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U126 ( .A(n985), .ZN(n703) );
  AOI22_X1 U127 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U128 ( .A(n984), .ZN(n702) );
  AOI22_X1 U129 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U130 ( .A(n983), .ZN(n701) );
  AOI22_X1 U131 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U132 ( .A(n982), .ZN(n700) );
  AOI22_X1 U133 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U134 ( .A(n981), .ZN(n699) );
  AOI22_X1 U135 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U136 ( .A(n980), .ZN(n698) );
  AOI22_X1 U137 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U138 ( .A(n948), .ZN(n671) );
  AOI22_X1 U139 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U140 ( .A(n947), .ZN(n670) );
  AOI22_X1 U141 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U142 ( .A(n946), .ZN(n669) );
  AOI22_X1 U143 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U144 ( .A(n945), .ZN(n668) );
  AOI22_X1 U145 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U146 ( .A(n944), .ZN(n667) );
  AOI22_X1 U147 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U148 ( .A(n943), .ZN(n666) );
  AOI22_X1 U149 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U150 ( .A(n915), .ZN(n641) );
  AOI22_X1 U151 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U152 ( .A(n913), .ZN(n640) );
  AOI22_X1 U153 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U154 ( .A(n912), .ZN(n639) );
  AOI22_X1 U155 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U156 ( .A(n911), .ZN(n638) );
  AOI22_X1 U157 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U158 ( .A(n910), .ZN(n637) );
  AOI22_X1 U159 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U160 ( .A(n909), .ZN(n636) );
  AOI22_X1 U161 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U162 ( .A(n908), .ZN(n635) );
  AOI22_X1 U163 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U164 ( .A(n907), .ZN(n634) );
  AOI22_X1 U165 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U166 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U167 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U168 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U169 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U170 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U171 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U172 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U173 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U174 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U175 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U176 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U177 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U178 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U179 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U180 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U181 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U182 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U183 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U184 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U185 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U186 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U187 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U188 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U189 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U190 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U191 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U192 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U193 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U194 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U195 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U196 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U197 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U198 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U199 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U200 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U201 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U202 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U203 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U204 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U205 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U206 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U207 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U208 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U209 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U210 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U211 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U212 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U213 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U214 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U215 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U216 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U217 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U218 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U219 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U220 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U221 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U222 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U223 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U224 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U225 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U226 ( .A(n999), .ZN(n715) );
  AOI22_X1 U227 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U228 ( .A(n998), .ZN(n714) );
  AOI22_X1 U229 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U230 ( .A(n951), .ZN(n673) );
  AOI22_X1 U231 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U232 ( .A(n949), .ZN(n672) );
  AOI22_X1 U233 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U234 ( .A(n979), .ZN(n697) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U236 ( .A(n977), .ZN(n696) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U238 ( .A(n976), .ZN(n695) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U240 ( .A(n975), .ZN(n694) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U242 ( .A(n974), .ZN(n693) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U244 ( .A(n973), .ZN(n692) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U246 ( .A(n972), .ZN(n691) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U248 ( .A(n971), .ZN(n690) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U250 ( .A(n970), .ZN(n689) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U252 ( .A(n968), .ZN(n688) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U254 ( .A(n967), .ZN(n687) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U256 ( .A(n966), .ZN(n686) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U258 ( .A(n965), .ZN(n685) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U260 ( .A(n964), .ZN(n684) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U262 ( .A(n963), .ZN(n683) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U264 ( .A(n962), .ZN(n682) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U266 ( .A(n942), .ZN(n665) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U268 ( .A(n940), .ZN(n664) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U270 ( .A(n939), .ZN(n663) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U272 ( .A(n938), .ZN(n662) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U274 ( .A(n937), .ZN(n661) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U276 ( .A(n936), .ZN(n660) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U278 ( .A(n935), .ZN(n659) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U280 ( .A(n934), .ZN(n658) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U282 ( .A(n933), .ZN(n657) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U284 ( .A(n931), .ZN(n656) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U286 ( .A(n930), .ZN(n655) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U288 ( .A(n929), .ZN(n654) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U290 ( .A(n928), .ZN(n653) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U292 ( .A(n927), .ZN(n652) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U294 ( .A(n926), .ZN(n651) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U296 ( .A(n925), .ZN(n650) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U298 ( .A(n906), .ZN(n633) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U300 ( .A(n904), .ZN(n632) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U302 ( .A(n903), .ZN(n631) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U304 ( .A(n902), .ZN(n630) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U306 ( .A(n901), .ZN(n629) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U308 ( .A(n900), .ZN(n628) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U310 ( .A(n899), .ZN(n627) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U312 ( .A(n898), .ZN(n626) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U314 ( .A(n897), .ZN(n625) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U316 ( .A(n895), .ZN(n624) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U318 ( .A(n894), .ZN(n623) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U320 ( .A(n893), .ZN(n622) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U322 ( .A(n892), .ZN(n621) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U324 ( .A(n891), .ZN(n620) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U326 ( .A(n890), .ZN(n619) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U328 ( .A(n889), .ZN(n618) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U330 ( .A(N12), .ZN(n253) );
  INV_X1 U331 ( .A(N11), .ZN(n252) );
  INV_X1 U332 ( .A(n997), .ZN(n713) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U334 ( .A(n995), .ZN(n712) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U336 ( .A(n994), .ZN(n711) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U338 ( .A(n993), .ZN(n710) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U340 ( .A(n992), .ZN(n709) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U342 ( .A(n991), .ZN(n708) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U344 ( .A(n990), .ZN(n707) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U346 ( .A(n989), .ZN(n706) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U348 ( .A(n924), .ZN(n649) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U350 ( .A(n922), .ZN(n648) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U352 ( .A(n921), .ZN(n647) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U354 ( .A(n920), .ZN(n646) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U356 ( .A(n919), .ZN(n645) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U358 ( .A(n918), .ZN(n644) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U360 ( .A(n917), .ZN(n643) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U362 ( .A(n916), .ZN(n642) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U364 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U366 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U368 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U370 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U372 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U374 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U376 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U378 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U380 ( .A(n961), .ZN(n681) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U382 ( .A(n959), .ZN(n680) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U384 ( .A(n958), .ZN(n679) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U386 ( .A(n957), .ZN(n678) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U388 ( .A(n956), .ZN(n677) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U390 ( .A(n955), .ZN(n676) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U392 ( .A(n954), .ZN(n675) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U394 ( .A(n953), .ZN(n674) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U396 ( .A(n888), .ZN(n617) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U398 ( .A(n886), .ZN(n616) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U400 ( .A(n885), .ZN(n615) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U402 ( .A(n884), .ZN(n614) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U404 ( .A(n883), .ZN(n613) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U406 ( .A(n882), .ZN(n612) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U408 ( .A(n881), .ZN(n611) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U410 ( .A(n880), .ZN(n610) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U412 ( .A(n879), .ZN(n609) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U414 ( .A(n877), .ZN(n608) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U416 ( .A(n876), .ZN(n607) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U418 ( .A(n875), .ZN(n606) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U420 ( .A(n874), .ZN(n605) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U422 ( .A(n873), .ZN(n604) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U424 ( .A(n872), .ZN(n603) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U426 ( .A(n871), .ZN(n602) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U428 ( .A(n870), .ZN(n601) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U430 ( .A(n868), .ZN(n600) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U432 ( .A(n867), .ZN(n599) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U434 ( .A(n866), .ZN(n598) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U436 ( .A(n865), .ZN(n597) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U438 ( .A(n864), .ZN(n596) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U440 ( .A(n863), .ZN(n595) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U442 ( .A(n862), .ZN(n594) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U444 ( .A(n861), .ZN(n293) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U446 ( .A(n859), .ZN(n292) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U448 ( .A(n858), .ZN(n291) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U450 ( .A(n857), .ZN(n290) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U452 ( .A(n856), .ZN(n289) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U454 ( .A(n855), .ZN(n288) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U456 ( .A(n854), .ZN(n287) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U458 ( .A(n853), .ZN(n286) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U460 ( .A(n852), .ZN(n285) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U462 ( .A(n850), .ZN(n284) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U464 ( .A(n849), .ZN(n283) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U466 ( .A(n848), .ZN(n282) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U468 ( .A(n847), .ZN(n281) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U470 ( .A(n846), .ZN(n280) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U472 ( .A(n845), .ZN(n279) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U474 ( .A(n844), .ZN(n278) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U476 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U477 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U478 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U479 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U480 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U481 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U482 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U483 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U484 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U485 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U486 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U487 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U488 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U489 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U490 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U491 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U492 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U494 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U496 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U498 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U500 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U502 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U504 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U506 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U508 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U510 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U512 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U514 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U516 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U518 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U520 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U522 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U524 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U526 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U528 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U530 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U532 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U534 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U536 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U538 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U540 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U542 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U544 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U546 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U548 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U550 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U552 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U554 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U556 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U558 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U560 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U562 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U564 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U566 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U568 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U570 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U572 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U574 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U576 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U578 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U580 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U582 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U584 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U586 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U588 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U590 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U592 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U594 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U596 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U598 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U600 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U602 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U604 ( .A(N13), .ZN(n842) );
  INV_X1 U605 ( .A(N14), .ZN(n843) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n248), .Z(n1) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n248), .Z(n2) );
  MUX2_X1 U608 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n248), .Z(n4) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n248), .Z(n5) );
  MUX2_X1 U611 ( .A(n5), .B(n4), .S(n244), .Z(n6) );
  MUX2_X1 U612 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n248), .Z(n8) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n249), .Z(n9) );
  MUX2_X1 U615 ( .A(n9), .B(n8), .S(n242), .Z(n10) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n248), .Z(n11) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n247), .Z(n12) );
  MUX2_X1 U618 ( .A(n12), .B(n11), .S(n242), .Z(n13) );
  MUX2_X1 U619 ( .A(n13), .B(n10), .S(N12), .Z(n14) );
  MUX2_X1 U620 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n245), .Z(n16) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n245), .Z(n17) );
  MUX2_X1 U623 ( .A(n17), .B(n16), .S(n242), .Z(n18) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n245), .Z(n20) );
  MUX2_X1 U626 ( .A(n20), .B(n19), .S(n242), .Z(n21) );
  MUX2_X1 U627 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n245), .Z(n23) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n245), .Z(n24) );
  MUX2_X1 U630 ( .A(n24), .B(n23), .S(n242), .Z(n25) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n245), .Z(n26) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n245), .Z(n27) );
  MUX2_X1 U633 ( .A(n27), .B(n26), .S(n242), .Z(n28) );
  MUX2_X1 U634 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U635 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U636 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n245), .Z(n31) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n245), .Z(n32) );
  MUX2_X1 U639 ( .A(n32), .B(n31), .S(n242), .Z(n33) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U642 ( .A(n35), .B(n34), .S(n242), .Z(n36) );
  MUX2_X1 U643 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n246), .Z(n38) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n246), .Z(n39) );
  MUX2_X1 U646 ( .A(n39), .B(n38), .S(n242), .Z(n40) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n246), .Z(n41) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n246), .Z(n42) );
  MUX2_X1 U649 ( .A(n42), .B(n41), .S(n242), .Z(n43) );
  MUX2_X1 U650 ( .A(n43), .B(n40), .S(n241), .Z(n44) );
  MUX2_X1 U651 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n246), .Z(n46) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n246), .Z(n47) );
  MUX2_X1 U654 ( .A(n47), .B(n46), .S(n242), .Z(n48) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n246), .Z(n49) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n246), .Z(n50) );
  MUX2_X1 U657 ( .A(n50), .B(n49), .S(n242), .Z(n51) );
  MUX2_X1 U658 ( .A(n51), .B(n48), .S(n241), .Z(n52) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n246), .Z(n53) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n246), .Z(n54) );
  MUX2_X1 U661 ( .A(n54), .B(n53), .S(n242), .Z(n55) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n246), .Z(n56) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n246), .Z(n57) );
  MUX2_X1 U664 ( .A(n57), .B(n56), .S(n242), .Z(n58) );
  MUX2_X1 U665 ( .A(n58), .B(n55), .S(n241), .Z(n59) );
  MUX2_X1 U666 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U667 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n250), .Z(n61) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n247), .Z(n62) );
  MUX2_X1 U670 ( .A(n62), .B(n61), .S(n243), .Z(n63) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n249), .Z(n64) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n245), .Z(n65) );
  MUX2_X1 U673 ( .A(n65), .B(n64), .S(n243), .Z(n66) );
  MUX2_X1 U674 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n250), .Z(n68) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n249), .Z(n69) );
  MUX2_X1 U677 ( .A(n69), .B(n68), .S(n243), .Z(n70) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n245), .Z(n71) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n249), .Z(n72) );
  MUX2_X1 U680 ( .A(n72), .B(n71), .S(n243), .Z(n73) );
  MUX2_X1 U681 ( .A(n73), .B(n70), .S(n241), .Z(n74) );
  MUX2_X1 U682 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n250), .Z(n76) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n247), .Z(n77) );
  MUX2_X1 U685 ( .A(n77), .B(n76), .S(n243), .Z(n78) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n246), .Z(n79) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n247), .Z(n80) );
  MUX2_X1 U688 ( .A(n80), .B(n79), .S(n243), .Z(n81) );
  MUX2_X1 U689 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n250), .Z(n83) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n250), .Z(n84) );
  MUX2_X1 U692 ( .A(n84), .B(n83), .S(n243), .Z(n85) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n250), .Z(n86) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n250), .Z(n87) );
  MUX2_X1 U695 ( .A(n87), .B(n86), .S(n243), .Z(n88) );
  MUX2_X1 U696 ( .A(n88), .B(n85), .S(n241), .Z(n89) );
  MUX2_X1 U697 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U698 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n247), .Z(n91) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n245), .Z(n92) );
  MUX2_X1 U701 ( .A(n92), .B(n91), .S(n243), .Z(n93) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n249), .Z(n94) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n250), .Z(n95) );
  MUX2_X1 U704 ( .A(n95), .B(n94), .S(n243), .Z(n96) );
  MUX2_X1 U705 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n249), .Z(n98) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n250), .Z(n99) );
  MUX2_X1 U708 ( .A(n99), .B(n98), .S(n243), .Z(n100) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n247), .Z(n101) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n250), .Z(n102) );
  MUX2_X1 U711 ( .A(n102), .B(n101), .S(n243), .Z(n103) );
  MUX2_X1 U712 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U713 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n247), .Z(n106) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n247), .Z(n107) );
  MUX2_X1 U716 ( .A(n107), .B(n106), .S(n244), .Z(n108) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n247), .Z(n109) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n247), .Z(n110) );
  MUX2_X1 U719 ( .A(n110), .B(n109), .S(n244), .Z(n111) );
  MUX2_X1 U720 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n247), .Z(n113) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n247), .Z(n114) );
  MUX2_X1 U723 ( .A(n114), .B(n113), .S(n244), .Z(n115) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n247), .Z(n116) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n247), .Z(n117) );
  MUX2_X1 U726 ( .A(n117), .B(n116), .S(n244), .Z(n118) );
  MUX2_X1 U727 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U728 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U729 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n247), .Z(n121) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n247), .Z(n122) );
  MUX2_X1 U732 ( .A(n122), .B(n121), .S(n244), .Z(n123) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n247), .Z(n124) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n247), .Z(n125) );
  MUX2_X1 U735 ( .A(n125), .B(n124), .S(n244), .Z(n126) );
  MUX2_X1 U736 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n248), .Z(n128) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n248), .Z(n129) );
  MUX2_X1 U739 ( .A(n129), .B(n128), .S(n244), .Z(n130) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n248), .Z(n131) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n248), .Z(n132) );
  MUX2_X1 U742 ( .A(n132), .B(n131), .S(n244), .Z(n133) );
  MUX2_X1 U743 ( .A(n133), .B(n130), .S(n241), .Z(n134) );
  MUX2_X1 U744 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n248), .Z(n136) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n248), .Z(n137) );
  MUX2_X1 U747 ( .A(n137), .B(n136), .S(n244), .Z(n138) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n248), .Z(n139) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n248), .Z(n140) );
  MUX2_X1 U750 ( .A(n140), .B(n139), .S(n244), .Z(n141) );
  MUX2_X1 U751 ( .A(n141), .B(n138), .S(n241), .Z(n142) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n248), .Z(n143) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n248), .Z(n144) );
  MUX2_X1 U754 ( .A(n144), .B(n143), .S(n244), .Z(n145) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n248), .Z(n146) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n248), .Z(n147) );
  MUX2_X1 U757 ( .A(n147), .B(n146), .S(n244), .Z(n148) );
  MUX2_X1 U758 ( .A(n148), .B(n145), .S(n241), .Z(n149) );
  MUX2_X1 U759 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U760 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n249), .Z(n151) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n249), .Z(n152) );
  MUX2_X1 U763 ( .A(n152), .B(n151), .S(N11), .Z(n153) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n249), .Z(n154) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n249), .Z(n155) );
  MUX2_X1 U766 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U767 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n249), .Z(n158) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n249), .Z(n159) );
  MUX2_X1 U770 ( .A(n159), .B(n158), .S(N11), .Z(n160) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n249), .Z(n161) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n249), .Z(n162) );
  MUX2_X1 U773 ( .A(n162), .B(n161), .S(n244), .Z(n163) );
  MUX2_X1 U774 ( .A(n163), .B(n160), .S(N12), .Z(n164) );
  MUX2_X1 U775 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n249), .Z(n166) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n249), .Z(n167) );
  MUX2_X1 U778 ( .A(n167), .B(n166), .S(N11), .Z(n168) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n249), .Z(n169) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n249), .Z(n170) );
  MUX2_X1 U781 ( .A(n170), .B(n169), .S(n243), .Z(n171) );
  MUX2_X1 U782 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(N10), .Z(n173) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n250), .Z(n174) );
  MUX2_X1 U785 ( .A(n174), .B(n173), .S(n242), .Z(n175) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n250), .Z(n176) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n250), .Z(n177) );
  MUX2_X1 U788 ( .A(n177), .B(n176), .S(n243), .Z(n178) );
  MUX2_X1 U789 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U790 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U791 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n246), .Z(n181) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n250), .Z(n182) );
  MUX2_X1 U794 ( .A(n182), .B(n181), .S(N11), .Z(n183) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n245), .Z(n184) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n248), .Z(n185) );
  MUX2_X1 U797 ( .A(n185), .B(n184), .S(N11), .Z(n186) );
  MUX2_X1 U798 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(N10), .Z(n188) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(N10), .Z(n189) );
  MUX2_X1 U801 ( .A(n189), .B(n188), .S(N11), .Z(n190) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n250), .Z(n191) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n250), .Z(n192) );
  MUX2_X1 U804 ( .A(n192), .B(n191), .S(n242), .Z(n193) );
  MUX2_X1 U805 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U806 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n246), .Z(n196) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n246), .Z(n197) );
  MUX2_X1 U809 ( .A(n197), .B(n196), .S(N11), .Z(n198) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(N10), .Z(n199) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n200) );
  MUX2_X1 U812 ( .A(n200), .B(n199), .S(n242), .Z(n201) );
  MUX2_X1 U813 ( .A(n201), .B(n198), .S(N12), .Z(n202) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n203) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n204) );
  MUX2_X1 U816 ( .A(n204), .B(n203), .S(n243), .Z(n205) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n250), .Z(n206) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n207) );
  MUX2_X1 U819 ( .A(n207), .B(n206), .S(N11), .Z(n208) );
  MUX2_X1 U820 ( .A(n208), .B(n205), .S(N12), .Z(n209) );
  MUX2_X1 U821 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U822 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n250), .Z(n211) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n245), .Z(n212) );
  MUX2_X1 U825 ( .A(n212), .B(n211), .S(n243), .Z(n213) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n246), .Z(n214) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n250), .Z(n215) );
  MUX2_X1 U828 ( .A(n215), .B(n214), .S(n244), .Z(n216) );
  MUX2_X1 U829 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(N10), .Z(n218) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(N10), .Z(n219) );
  MUX2_X1 U832 ( .A(n219), .B(n218), .S(n244), .Z(n220) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n248), .Z(n221) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n246), .Z(n222) );
  MUX2_X1 U835 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U836 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U837 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n248), .Z(n226) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n227) );
  MUX2_X1 U840 ( .A(n227), .B(n226), .S(n243), .Z(n228) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n248), .Z(n229) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n250), .Z(n230) );
  MUX2_X1 U843 ( .A(n230), .B(n229), .S(N11), .Z(n231) );
  MUX2_X1 U844 ( .A(n231), .B(n228), .S(N12), .Z(n232) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n233) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n234) );
  MUX2_X1 U847 ( .A(n234), .B(n233), .S(n244), .Z(n235) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n248), .Z(n236) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n237) );
  MUX2_X1 U850 ( .A(n237), .B(n236), .S(N11), .Z(n238) );
  MUX2_X1 U851 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U852 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U853 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_27 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  BUF_X1 U3 ( .A(N10), .Z(n247) );
  BUF_X1 U4 ( .A(n250), .Z(n248) );
  BUF_X1 U5 ( .A(n250), .Z(n249) );
  BUF_X1 U6 ( .A(n250), .Z(n246) );
  BUF_X1 U7 ( .A(n250), .Z(n245) );
  BUF_X1 U8 ( .A(N10), .Z(n250) );
  INV_X1 U9 ( .A(n1111), .ZN(n841) );
  INV_X1 U10 ( .A(n1100), .ZN(n840) );
  INV_X1 U11 ( .A(n1090), .ZN(n839) );
  INV_X1 U12 ( .A(n1080), .ZN(n838) );
  INV_X1 U13 ( .A(n1070), .ZN(n837) );
  INV_X1 U14 ( .A(n1060), .ZN(n836) );
  INV_X1 U15 ( .A(n1051), .ZN(n835) );
  INV_X1 U16 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U19 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U20 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U21 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U22 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U23 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U24 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U26 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U27 ( .A(n1131), .ZN(n816) );
  INV_X1 U28 ( .A(n1121), .ZN(n815) );
  INV_X1 U29 ( .A(n887), .ZN(n814) );
  INV_X1 U30 ( .A(n878), .ZN(n813) );
  INV_X1 U31 ( .A(n869), .ZN(n812) );
  INV_X1 U32 ( .A(n860), .ZN(n811) );
  INV_X1 U33 ( .A(n851), .ZN(n810) );
  INV_X1 U34 ( .A(n987), .ZN(n828) );
  INV_X1 U35 ( .A(n978), .ZN(n827) );
  INV_X1 U36 ( .A(n969), .ZN(n826) );
  INV_X1 U37 ( .A(n914), .ZN(n820) );
  INV_X1 U38 ( .A(n905), .ZN(n819) );
  INV_X1 U39 ( .A(n896), .ZN(n818) );
  INV_X1 U40 ( .A(n1033), .ZN(n833) );
  INV_X1 U41 ( .A(n1023), .ZN(n832) );
  INV_X1 U42 ( .A(n1014), .ZN(n831) );
  INV_X1 U43 ( .A(n1005), .ZN(n830) );
  INV_X1 U44 ( .A(n996), .ZN(n829) );
  INV_X1 U45 ( .A(n960), .ZN(n825) );
  INV_X1 U46 ( .A(n950), .ZN(n824) );
  INV_X1 U47 ( .A(n941), .ZN(n823) );
  INV_X1 U48 ( .A(n932), .ZN(n822) );
  INV_X1 U49 ( .A(n923), .ZN(n821) );
  INV_X1 U50 ( .A(n1142), .ZN(n817) );
  BUF_X1 U51 ( .A(N11), .Z(n243) );
  BUF_X1 U52 ( .A(N11), .Z(n244) );
  INV_X1 U53 ( .A(N10), .ZN(n251) );
  BUF_X1 U54 ( .A(N12), .Z(n241) );
  NOR3_X1 U55 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U56 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U57 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U58 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U59 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U60 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U61 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U62 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U63 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U64 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U65 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U67 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U69 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U70 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U71 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U72 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U73 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U74 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U75 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U76 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U77 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U79 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U81 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U82 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U83 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U84 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U85 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U86 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U87 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U88 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U89 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U90 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U91 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U92 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U93 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U94 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U95 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U96 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U97 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U98 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U99 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U100 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U101 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U102 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U103 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U104 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U105 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U106 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U107 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U108 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U109 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U110 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U111 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U112 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U113 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U114 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U115 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U116 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U117 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U118 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U119 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U120 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U121 ( .A(n988), .ZN(n705) );
  AOI22_X1 U122 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U123 ( .A(n986), .ZN(n704) );
  AOI22_X1 U124 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U125 ( .A(n985), .ZN(n703) );
  AOI22_X1 U126 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U127 ( .A(n984), .ZN(n702) );
  AOI22_X1 U128 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U129 ( .A(n983), .ZN(n701) );
  AOI22_X1 U130 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U131 ( .A(n982), .ZN(n700) );
  AOI22_X1 U132 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U133 ( .A(n981), .ZN(n699) );
  AOI22_X1 U134 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U135 ( .A(n980), .ZN(n698) );
  AOI22_X1 U136 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U137 ( .A(n949), .ZN(n672) );
  AOI22_X1 U138 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U139 ( .A(n948), .ZN(n671) );
  AOI22_X1 U140 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U141 ( .A(n947), .ZN(n670) );
  AOI22_X1 U142 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U143 ( .A(n946), .ZN(n669) );
  AOI22_X1 U144 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U145 ( .A(n945), .ZN(n668) );
  AOI22_X1 U146 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U147 ( .A(n944), .ZN(n667) );
  AOI22_X1 U148 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U149 ( .A(n943), .ZN(n666) );
  AOI22_X1 U150 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U151 ( .A(n915), .ZN(n641) );
  AOI22_X1 U152 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U153 ( .A(n913), .ZN(n640) );
  AOI22_X1 U154 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U155 ( .A(n912), .ZN(n639) );
  AOI22_X1 U156 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U157 ( .A(n911), .ZN(n638) );
  AOI22_X1 U158 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U159 ( .A(n910), .ZN(n637) );
  AOI22_X1 U160 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U161 ( .A(n909), .ZN(n636) );
  AOI22_X1 U162 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U163 ( .A(n908), .ZN(n635) );
  AOI22_X1 U164 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U165 ( .A(n907), .ZN(n634) );
  AOI22_X1 U166 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U167 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U168 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U169 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U170 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U171 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U172 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U173 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U174 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U175 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U176 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U177 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U178 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U179 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U180 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U181 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U182 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U183 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U184 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U185 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U186 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U187 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U188 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U189 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U190 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U191 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U192 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U193 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U194 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U195 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U196 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U197 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U198 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U199 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U200 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U201 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U202 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U203 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U204 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U205 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U206 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U207 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U208 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U209 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U210 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U211 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U212 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U213 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U214 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U215 ( .A(n998), .ZN(n714) );
  AOI22_X1 U216 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U217 ( .A(n951), .ZN(n673) );
  AOI22_X1 U218 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U219 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U220 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U221 ( .A(n999), .ZN(n715) );
  AOI22_X1 U222 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U223 ( .A(n979), .ZN(n697) );
  AOI22_X1 U224 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U225 ( .A(n977), .ZN(n696) );
  AOI22_X1 U226 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U227 ( .A(n976), .ZN(n695) );
  AOI22_X1 U228 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U229 ( .A(n975), .ZN(n694) );
  AOI22_X1 U230 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U231 ( .A(n974), .ZN(n693) );
  AOI22_X1 U232 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U233 ( .A(n973), .ZN(n692) );
  AOI22_X1 U234 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U235 ( .A(n972), .ZN(n691) );
  AOI22_X1 U236 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U237 ( .A(n971), .ZN(n690) );
  AOI22_X1 U238 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U239 ( .A(n970), .ZN(n689) );
  AOI22_X1 U240 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U241 ( .A(n968), .ZN(n688) );
  AOI22_X1 U242 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U243 ( .A(n967), .ZN(n687) );
  AOI22_X1 U244 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U245 ( .A(n966), .ZN(n686) );
  AOI22_X1 U246 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U247 ( .A(n965), .ZN(n685) );
  AOI22_X1 U248 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U249 ( .A(n964), .ZN(n684) );
  AOI22_X1 U250 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U251 ( .A(n963), .ZN(n683) );
  AOI22_X1 U252 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U253 ( .A(n962), .ZN(n682) );
  AOI22_X1 U254 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U255 ( .A(n942), .ZN(n665) );
  AOI22_X1 U256 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U257 ( .A(n940), .ZN(n664) );
  AOI22_X1 U258 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U259 ( .A(n939), .ZN(n663) );
  AOI22_X1 U260 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U261 ( .A(n938), .ZN(n662) );
  AOI22_X1 U262 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U263 ( .A(n937), .ZN(n661) );
  AOI22_X1 U264 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U265 ( .A(n936), .ZN(n660) );
  AOI22_X1 U266 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U267 ( .A(n935), .ZN(n659) );
  AOI22_X1 U268 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U269 ( .A(n934), .ZN(n658) );
  AOI22_X1 U270 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U271 ( .A(n933), .ZN(n657) );
  AOI22_X1 U272 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U273 ( .A(n931), .ZN(n656) );
  AOI22_X1 U274 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U275 ( .A(n930), .ZN(n655) );
  AOI22_X1 U276 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U277 ( .A(n929), .ZN(n654) );
  AOI22_X1 U278 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U279 ( .A(n928), .ZN(n653) );
  AOI22_X1 U280 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U281 ( .A(n927), .ZN(n652) );
  AOI22_X1 U282 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U283 ( .A(n926), .ZN(n651) );
  AOI22_X1 U284 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U285 ( .A(n925), .ZN(n650) );
  AOI22_X1 U286 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U287 ( .A(n906), .ZN(n633) );
  AOI22_X1 U288 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U289 ( .A(n904), .ZN(n632) );
  AOI22_X1 U290 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U291 ( .A(n903), .ZN(n631) );
  AOI22_X1 U292 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U293 ( .A(n902), .ZN(n630) );
  AOI22_X1 U294 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U295 ( .A(n901), .ZN(n629) );
  AOI22_X1 U296 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U297 ( .A(n900), .ZN(n628) );
  AOI22_X1 U298 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U299 ( .A(n899), .ZN(n627) );
  AOI22_X1 U300 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U301 ( .A(n898), .ZN(n626) );
  AOI22_X1 U302 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U303 ( .A(n897), .ZN(n625) );
  AOI22_X1 U304 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U305 ( .A(n895), .ZN(n624) );
  AOI22_X1 U306 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U307 ( .A(n894), .ZN(n623) );
  AOI22_X1 U308 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U309 ( .A(n893), .ZN(n622) );
  AOI22_X1 U310 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U311 ( .A(n892), .ZN(n621) );
  AOI22_X1 U312 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U313 ( .A(n891), .ZN(n620) );
  AOI22_X1 U314 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U315 ( .A(n890), .ZN(n619) );
  AOI22_X1 U316 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U317 ( .A(n889), .ZN(n618) );
  AOI22_X1 U318 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U319 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U320 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U321 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U322 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U323 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U324 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U325 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U326 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U327 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U328 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U329 ( .A(N12), .ZN(n253) );
  INV_X1 U330 ( .A(N11), .ZN(n252) );
  INV_X1 U331 ( .A(n997), .ZN(n713) );
  AOI22_X1 U332 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U333 ( .A(n995), .ZN(n712) );
  AOI22_X1 U334 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U335 ( .A(n994), .ZN(n711) );
  AOI22_X1 U336 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U337 ( .A(n993), .ZN(n710) );
  AOI22_X1 U338 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U339 ( .A(n992), .ZN(n709) );
  AOI22_X1 U340 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U341 ( .A(n991), .ZN(n708) );
  AOI22_X1 U342 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U343 ( .A(n990), .ZN(n707) );
  AOI22_X1 U344 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U345 ( .A(n989), .ZN(n706) );
  AOI22_X1 U346 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U347 ( .A(n924), .ZN(n649) );
  AOI22_X1 U348 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U349 ( .A(n922), .ZN(n648) );
  AOI22_X1 U350 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U351 ( .A(n921), .ZN(n647) );
  AOI22_X1 U352 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U353 ( .A(n920), .ZN(n646) );
  AOI22_X1 U354 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U355 ( .A(n919), .ZN(n645) );
  AOI22_X1 U356 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U357 ( .A(n918), .ZN(n644) );
  AOI22_X1 U358 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U359 ( .A(n917), .ZN(n643) );
  AOI22_X1 U360 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U361 ( .A(n916), .ZN(n642) );
  AOI22_X1 U362 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U363 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U364 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U365 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U366 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U367 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U368 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U369 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U370 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U371 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U372 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U373 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U374 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U375 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U376 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U377 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U378 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U379 ( .A(n961), .ZN(n681) );
  AOI22_X1 U380 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U381 ( .A(n959), .ZN(n680) );
  AOI22_X1 U382 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U383 ( .A(n958), .ZN(n679) );
  AOI22_X1 U384 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U385 ( .A(n957), .ZN(n678) );
  AOI22_X1 U386 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U387 ( .A(n956), .ZN(n677) );
  AOI22_X1 U388 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U389 ( .A(n955), .ZN(n676) );
  AOI22_X1 U390 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U391 ( .A(n954), .ZN(n675) );
  AOI22_X1 U392 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U393 ( .A(n953), .ZN(n674) );
  AOI22_X1 U394 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U395 ( .A(n888), .ZN(n617) );
  AOI22_X1 U396 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U397 ( .A(n886), .ZN(n616) );
  AOI22_X1 U398 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U399 ( .A(n885), .ZN(n615) );
  AOI22_X1 U400 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U401 ( .A(n884), .ZN(n614) );
  AOI22_X1 U402 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U403 ( .A(n883), .ZN(n613) );
  AOI22_X1 U404 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U405 ( .A(n882), .ZN(n612) );
  AOI22_X1 U406 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U407 ( .A(n881), .ZN(n611) );
  AOI22_X1 U408 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U409 ( .A(n880), .ZN(n610) );
  AOI22_X1 U410 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U411 ( .A(n879), .ZN(n609) );
  AOI22_X1 U412 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U413 ( .A(n877), .ZN(n608) );
  AOI22_X1 U414 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U415 ( .A(n876), .ZN(n607) );
  AOI22_X1 U416 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U417 ( .A(n875), .ZN(n606) );
  AOI22_X1 U418 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U419 ( .A(n874), .ZN(n605) );
  AOI22_X1 U420 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U421 ( .A(n873), .ZN(n604) );
  AOI22_X1 U422 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U423 ( .A(n872), .ZN(n603) );
  AOI22_X1 U424 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U425 ( .A(n871), .ZN(n602) );
  AOI22_X1 U426 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U427 ( .A(n870), .ZN(n601) );
  AOI22_X1 U428 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U429 ( .A(n868), .ZN(n600) );
  AOI22_X1 U430 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U431 ( .A(n867), .ZN(n599) );
  AOI22_X1 U432 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U433 ( .A(n866), .ZN(n598) );
  AOI22_X1 U434 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U435 ( .A(n865), .ZN(n597) );
  AOI22_X1 U436 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U437 ( .A(n864), .ZN(n596) );
  AOI22_X1 U438 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U439 ( .A(n863), .ZN(n595) );
  AOI22_X1 U440 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U441 ( .A(n862), .ZN(n594) );
  AOI22_X1 U442 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U443 ( .A(n861), .ZN(n293) );
  AOI22_X1 U444 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U445 ( .A(n859), .ZN(n292) );
  AOI22_X1 U446 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U447 ( .A(n858), .ZN(n291) );
  AOI22_X1 U448 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U449 ( .A(n857), .ZN(n290) );
  AOI22_X1 U450 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U451 ( .A(n856), .ZN(n289) );
  AOI22_X1 U452 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U453 ( .A(n855), .ZN(n288) );
  AOI22_X1 U454 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U455 ( .A(n854), .ZN(n287) );
  AOI22_X1 U456 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U457 ( .A(n853), .ZN(n286) );
  AOI22_X1 U458 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U459 ( .A(n852), .ZN(n285) );
  AOI22_X1 U460 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U461 ( .A(n850), .ZN(n284) );
  AOI22_X1 U462 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U463 ( .A(n849), .ZN(n283) );
  AOI22_X1 U464 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U465 ( .A(n848), .ZN(n282) );
  AOI22_X1 U466 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U467 ( .A(n847), .ZN(n281) );
  AOI22_X1 U468 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U469 ( .A(n846), .ZN(n280) );
  AOI22_X1 U470 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U471 ( .A(n845), .ZN(n279) );
  AOI22_X1 U472 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U473 ( .A(n844), .ZN(n278) );
  AOI22_X1 U474 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U475 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U476 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U477 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U478 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U479 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U480 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U481 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U482 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U483 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U484 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U485 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U486 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U487 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U488 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U489 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U490 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U491 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U492 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U493 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U494 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U495 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U496 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U497 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U498 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U499 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U500 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U501 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U502 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U503 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U504 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U505 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U506 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U507 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U508 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U509 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U510 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U511 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U512 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U513 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U514 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U515 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U516 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U517 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U518 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U519 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U520 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U521 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U522 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U523 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U524 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U525 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U526 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U527 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U528 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U529 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U530 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U531 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U532 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U533 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U534 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U535 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U536 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U537 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U538 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U539 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U540 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U541 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U542 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U543 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U544 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U545 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U546 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U547 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U548 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U549 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U550 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U551 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U552 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U553 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U554 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U555 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U556 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U557 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U558 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U559 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U560 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U561 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U562 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U563 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U564 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U565 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U566 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U567 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U568 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U569 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U570 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U571 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U572 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U573 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U574 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U575 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U576 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U577 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U578 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U579 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U580 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U581 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U582 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U583 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U584 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U585 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U586 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U587 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U588 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U589 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U590 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U591 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U592 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U593 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U594 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U595 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U596 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U597 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U598 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U599 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U600 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U601 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U602 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U603 ( .A(N13), .ZN(n842) );
  INV_X1 U604 ( .A(N14), .ZN(n843) );
  MUX2_X1 U605 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n247), .Z(n1) );
  MUX2_X1 U606 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n247), .Z(n2) );
  MUX2_X1 U607 ( .A(n2), .B(n1), .S(n242), .Z(n3) );
  MUX2_X1 U608 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n247), .Z(n4) );
  MUX2_X1 U609 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n247), .Z(n5) );
  MUX2_X1 U610 ( .A(n5), .B(n4), .S(n242), .Z(n6) );
  MUX2_X1 U611 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U612 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n247), .Z(n8) );
  MUX2_X1 U613 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n249), .Z(n9) );
  MUX2_X1 U614 ( .A(n9), .B(n8), .S(n242), .Z(n10) );
  MUX2_X1 U615 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n247), .Z(n11) );
  MUX2_X1 U616 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n248), .Z(n12) );
  MUX2_X1 U617 ( .A(n12), .B(n11), .S(n242), .Z(n13) );
  MUX2_X1 U618 ( .A(n13), .B(n10), .S(N12), .Z(n14) );
  MUX2_X1 U619 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U620 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n245), .Z(n16) );
  MUX2_X1 U621 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n245), .Z(n17) );
  MUX2_X1 U622 ( .A(n17), .B(n16), .S(n243), .Z(n18) );
  MUX2_X1 U623 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U624 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n245), .Z(n20) );
  MUX2_X1 U625 ( .A(n20), .B(n19), .S(n243), .Z(n21) );
  MUX2_X1 U626 ( .A(n21), .B(n18), .S(N12), .Z(n22) );
  MUX2_X1 U627 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n245), .Z(n23) );
  MUX2_X1 U628 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n245), .Z(n24) );
  MUX2_X1 U629 ( .A(n24), .B(n23), .S(n243), .Z(n25) );
  MUX2_X1 U630 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n245), .Z(n26) );
  MUX2_X1 U631 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n245), .Z(n27) );
  MUX2_X1 U632 ( .A(n27), .B(n26), .S(n243), .Z(n28) );
  MUX2_X1 U633 ( .A(n28), .B(n25), .S(N12), .Z(n29) );
  MUX2_X1 U634 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U635 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U636 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n245), .Z(n31) );
  MUX2_X1 U637 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n245), .Z(n32) );
  MUX2_X1 U638 ( .A(n32), .B(n31), .S(n243), .Z(n33) );
  MUX2_X1 U639 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U640 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U641 ( .A(n35), .B(n34), .S(n243), .Z(n36) );
  MUX2_X1 U642 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U643 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n246), .Z(n38) );
  MUX2_X1 U644 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n246), .Z(n39) );
  MUX2_X1 U645 ( .A(n39), .B(n38), .S(n243), .Z(n40) );
  MUX2_X1 U646 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n246), .Z(n41) );
  MUX2_X1 U647 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n246), .Z(n42) );
  MUX2_X1 U648 ( .A(n42), .B(n41), .S(n243), .Z(n43) );
  MUX2_X1 U649 ( .A(n43), .B(n40), .S(n241), .Z(n44) );
  MUX2_X1 U650 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U651 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n246), .Z(n46) );
  MUX2_X1 U652 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n246), .Z(n47) );
  MUX2_X1 U653 ( .A(n47), .B(n46), .S(n243), .Z(n48) );
  MUX2_X1 U654 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n246), .Z(n49) );
  MUX2_X1 U655 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n246), .Z(n50) );
  MUX2_X1 U656 ( .A(n50), .B(n49), .S(n243), .Z(n51) );
  MUX2_X1 U657 ( .A(n51), .B(n48), .S(n241), .Z(n52) );
  MUX2_X1 U658 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n246), .Z(n53) );
  MUX2_X1 U659 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n246), .Z(n54) );
  MUX2_X1 U660 ( .A(n54), .B(n53), .S(n243), .Z(n55) );
  MUX2_X1 U661 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n246), .Z(n56) );
  MUX2_X1 U662 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n246), .Z(n57) );
  MUX2_X1 U663 ( .A(n57), .B(n56), .S(n243), .Z(n58) );
  MUX2_X1 U664 ( .A(n58), .B(n55), .S(n241), .Z(n59) );
  MUX2_X1 U665 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U666 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U667 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n245), .Z(n61) );
  MUX2_X1 U668 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n245), .Z(n62) );
  MUX2_X1 U669 ( .A(n62), .B(n61), .S(n244), .Z(n63) );
  MUX2_X1 U670 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n246), .Z(n64) );
  MUX2_X1 U671 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n249), .Z(n65) );
  MUX2_X1 U672 ( .A(n65), .B(n64), .S(n244), .Z(n66) );
  MUX2_X1 U673 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U674 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n248), .Z(n68) );
  MUX2_X1 U675 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n246), .Z(n69) );
  MUX2_X1 U676 ( .A(n69), .B(n68), .S(n244), .Z(n70) );
  MUX2_X1 U677 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n246), .Z(n71) );
  MUX2_X1 U678 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n245), .Z(n72) );
  MUX2_X1 U679 ( .A(n72), .B(n71), .S(n244), .Z(n73) );
  MUX2_X1 U680 ( .A(n73), .B(n70), .S(n241), .Z(n74) );
  MUX2_X1 U681 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U682 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n248), .Z(n76) );
  MUX2_X1 U683 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n248), .Z(n77) );
  MUX2_X1 U684 ( .A(n77), .B(n76), .S(n244), .Z(n78) );
  MUX2_X1 U685 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n249), .Z(n79) );
  MUX2_X1 U686 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n248), .Z(n80) );
  MUX2_X1 U687 ( .A(n80), .B(n79), .S(n244), .Z(n81) );
  MUX2_X1 U688 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U689 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n250), .Z(n83) );
  MUX2_X1 U690 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n250), .Z(n84) );
  MUX2_X1 U691 ( .A(n84), .B(n83), .S(n244), .Z(n85) );
  MUX2_X1 U692 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n250), .Z(n86) );
  MUX2_X1 U693 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n246), .Z(n87) );
  MUX2_X1 U694 ( .A(n87), .B(n86), .S(n244), .Z(n88) );
  MUX2_X1 U695 ( .A(n88), .B(n85), .S(n241), .Z(n89) );
  MUX2_X1 U696 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U697 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U698 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n250), .Z(n91) );
  MUX2_X1 U699 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n92) );
  MUX2_X1 U700 ( .A(n92), .B(n91), .S(n244), .Z(n93) );
  MUX2_X1 U701 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U702 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n250), .Z(n95) );
  MUX2_X1 U703 ( .A(n95), .B(n94), .S(n244), .Z(n96) );
  MUX2_X1 U704 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U705 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n98) );
  MUX2_X1 U706 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n250), .Z(n99) );
  MUX2_X1 U707 ( .A(n99), .B(n98), .S(n244), .Z(n100) );
  MUX2_X1 U708 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n250), .Z(n101) );
  MUX2_X1 U709 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n250), .Z(n102) );
  MUX2_X1 U710 ( .A(n102), .B(n101), .S(n244), .Z(n103) );
  MUX2_X1 U711 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U712 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U713 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n247), .Z(n106) );
  MUX2_X1 U714 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n247), .Z(n107) );
  MUX2_X1 U715 ( .A(n107), .B(n106), .S(n243), .Z(n108) );
  MUX2_X1 U716 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n247), .Z(n109) );
  MUX2_X1 U717 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n247), .Z(n110) );
  MUX2_X1 U718 ( .A(n110), .B(n109), .S(N11), .Z(n111) );
  MUX2_X1 U719 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U720 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n247), .Z(n113) );
  MUX2_X1 U721 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n247), .Z(n114) );
  MUX2_X1 U722 ( .A(n114), .B(n113), .S(n244), .Z(n115) );
  MUX2_X1 U723 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n247), .Z(n116) );
  MUX2_X1 U724 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n247), .Z(n117) );
  MUX2_X1 U725 ( .A(n117), .B(n116), .S(N11), .Z(n118) );
  MUX2_X1 U726 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U727 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U728 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U729 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n247), .Z(n121) );
  MUX2_X1 U730 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n247), .Z(n122) );
  MUX2_X1 U731 ( .A(n122), .B(n121), .S(N11), .Z(n123) );
  MUX2_X1 U732 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n247), .Z(n124) );
  MUX2_X1 U733 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n247), .Z(n125) );
  MUX2_X1 U734 ( .A(n125), .B(n124), .S(N11), .Z(n126) );
  MUX2_X1 U735 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U736 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n248), .Z(n128) );
  MUX2_X1 U737 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n248), .Z(n129) );
  MUX2_X1 U738 ( .A(n129), .B(n128), .S(N11), .Z(n130) );
  MUX2_X1 U739 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n248), .Z(n131) );
  MUX2_X1 U740 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n248), .Z(n132) );
  MUX2_X1 U741 ( .A(n132), .B(n131), .S(n242), .Z(n133) );
  MUX2_X1 U742 ( .A(n133), .B(n130), .S(n241), .Z(n134) );
  MUX2_X1 U743 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U744 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n248), .Z(n136) );
  MUX2_X1 U745 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n248), .Z(n137) );
  MUX2_X1 U746 ( .A(n137), .B(n136), .S(N11), .Z(n138) );
  MUX2_X1 U747 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n248), .Z(n139) );
  MUX2_X1 U748 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n248), .Z(n140) );
  MUX2_X1 U749 ( .A(n140), .B(n139), .S(n244), .Z(n141) );
  MUX2_X1 U750 ( .A(n141), .B(n138), .S(n241), .Z(n142) );
  MUX2_X1 U751 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n248), .Z(n143) );
  MUX2_X1 U752 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n248), .Z(n144) );
  MUX2_X1 U753 ( .A(n144), .B(n143), .S(n243), .Z(n145) );
  MUX2_X1 U754 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n248), .Z(n146) );
  MUX2_X1 U755 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n248), .Z(n147) );
  MUX2_X1 U756 ( .A(n147), .B(n146), .S(n244), .Z(n148) );
  MUX2_X1 U757 ( .A(n148), .B(n145), .S(n241), .Z(n149) );
  MUX2_X1 U758 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U759 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U760 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n249), .Z(n151) );
  MUX2_X1 U761 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n249), .Z(n152) );
  MUX2_X1 U762 ( .A(n152), .B(n151), .S(n243), .Z(n153) );
  MUX2_X1 U763 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n249), .Z(n154) );
  MUX2_X1 U764 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n249), .Z(n155) );
  MUX2_X1 U765 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U766 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U767 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n249), .Z(n158) );
  MUX2_X1 U768 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n249), .Z(n159) );
  MUX2_X1 U769 ( .A(n159), .B(n158), .S(n242), .Z(n160) );
  MUX2_X1 U770 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n249), .Z(n161) );
  MUX2_X1 U771 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n249), .Z(n162) );
  MUX2_X1 U772 ( .A(n162), .B(n161), .S(N11), .Z(n163) );
  MUX2_X1 U773 ( .A(n163), .B(n160), .S(N12), .Z(n164) );
  MUX2_X1 U774 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U775 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n249), .Z(n166) );
  MUX2_X1 U776 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n249), .Z(n167) );
  MUX2_X1 U777 ( .A(n167), .B(n166), .S(n244), .Z(n168) );
  MUX2_X1 U778 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n249), .Z(n169) );
  MUX2_X1 U779 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n249), .Z(n170) );
  MUX2_X1 U780 ( .A(n170), .B(n169), .S(N11), .Z(n171) );
  MUX2_X1 U781 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U782 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n247), .Z(n173) );
  MUX2_X1 U783 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(N10), .Z(n174) );
  MUX2_X1 U784 ( .A(n174), .B(n173), .S(n242), .Z(n175) );
  MUX2_X1 U785 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n176) );
  MUX2_X1 U786 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n250), .Z(n177) );
  MUX2_X1 U787 ( .A(n177), .B(n176), .S(N11), .Z(n178) );
  MUX2_X1 U788 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U789 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U790 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U791 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n249), .Z(n181) );
  MUX2_X1 U792 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n250), .Z(n182) );
  MUX2_X1 U793 ( .A(n182), .B(n181), .S(N11), .Z(n183) );
  MUX2_X1 U794 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n248), .Z(n184) );
  MUX2_X1 U795 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n245), .Z(n185) );
  MUX2_X1 U796 ( .A(n185), .B(n184), .S(n244), .Z(n186) );
  MUX2_X1 U797 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U798 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n250), .Z(n188) );
  MUX2_X1 U799 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n245), .Z(n189) );
  MUX2_X1 U800 ( .A(n189), .B(n188), .S(n243), .Z(n190) );
  MUX2_X1 U801 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n246), .Z(n191) );
  MUX2_X1 U802 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(N10), .Z(n192) );
  MUX2_X1 U803 ( .A(n192), .B(n191), .S(N11), .Z(n193) );
  MUX2_X1 U804 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U805 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U806 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n245), .Z(n196) );
  MUX2_X1 U807 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n250), .Z(n197) );
  MUX2_X1 U808 ( .A(n197), .B(n196), .S(n242), .Z(n198) );
  MUX2_X1 U809 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n250), .Z(n199) );
  MUX2_X1 U810 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n200) );
  MUX2_X1 U811 ( .A(n200), .B(n199), .S(n243), .Z(n201) );
  MUX2_X1 U812 ( .A(n201), .B(n198), .S(n241), .Z(n202) );
  MUX2_X1 U813 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n250), .Z(n203) );
  MUX2_X1 U814 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n204) );
  MUX2_X1 U815 ( .A(n204), .B(n203), .S(n242), .Z(n205) );
  MUX2_X1 U816 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n206) );
  MUX2_X1 U817 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n207) );
  MUX2_X1 U818 ( .A(n207), .B(n206), .S(n244), .Z(n208) );
  MUX2_X1 U819 ( .A(n208), .B(n205), .S(N12), .Z(n209) );
  MUX2_X1 U820 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U821 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U822 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n250), .Z(n211) );
  MUX2_X1 U823 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n246), .Z(n212) );
  MUX2_X1 U824 ( .A(n212), .B(n211), .S(n242), .Z(n213) );
  MUX2_X1 U825 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n249), .Z(n214) );
  MUX2_X1 U826 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(N10), .Z(n215) );
  MUX2_X1 U827 ( .A(n215), .B(n214), .S(n242), .Z(n216) );
  MUX2_X1 U828 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U829 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n247), .Z(n218) );
  MUX2_X1 U830 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n250), .Z(n219) );
  MUX2_X1 U831 ( .A(n219), .B(n218), .S(n242), .Z(n220) );
  MUX2_X1 U832 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n247), .Z(n221) );
  MUX2_X1 U833 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n222) );
  MUX2_X1 U834 ( .A(n222), .B(n221), .S(n243), .Z(n223) );
  MUX2_X1 U835 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U836 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U837 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n247), .Z(n226) );
  MUX2_X1 U838 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n250), .Z(n227) );
  MUX2_X1 U839 ( .A(n227), .B(n226), .S(n242), .Z(n228) );
  MUX2_X1 U840 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n247), .Z(n229) );
  MUX2_X1 U841 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n230) );
  MUX2_X1 U842 ( .A(n230), .B(n229), .S(N11), .Z(n231) );
  MUX2_X1 U843 ( .A(n231), .B(n228), .S(n241), .Z(n232) );
  MUX2_X1 U844 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n233) );
  MUX2_X1 U845 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n234) );
  MUX2_X1 U846 ( .A(n234), .B(n233), .S(n242), .Z(n235) );
  MUX2_X1 U847 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n236) );
  MUX2_X1 U848 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n237) );
  MUX2_X1 U849 ( .A(n237), .B(n236), .S(n242), .Z(n238) );
  MUX2_X1 U850 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U851 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U852 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U853 ( .A(N11), .Z(n242) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_26 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X2 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(N10), .Z(n248) );
  BUF_X1 U4 ( .A(n250), .Z(n249) );
  BUF_X1 U5 ( .A(n250), .Z(n246) );
  BUF_X1 U6 ( .A(n250), .Z(n245) );
  BUF_X1 U7 ( .A(n250), .Z(n247) );
  BUF_X1 U8 ( .A(N10), .Z(n250) );
  INV_X1 U9 ( .A(n1111), .ZN(n841) );
  INV_X1 U10 ( .A(n1100), .ZN(n840) );
  INV_X1 U11 ( .A(n1090), .ZN(n839) );
  INV_X1 U12 ( .A(n1080), .ZN(n838) );
  INV_X1 U13 ( .A(n1070), .ZN(n837) );
  INV_X1 U14 ( .A(n1060), .ZN(n836) );
  INV_X1 U15 ( .A(n1051), .ZN(n835) );
  INV_X1 U16 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U19 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U20 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U21 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U22 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U23 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U24 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U26 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U27 ( .A(n1131), .ZN(n816) );
  INV_X1 U28 ( .A(n1121), .ZN(n815) );
  INV_X1 U29 ( .A(n887), .ZN(n814) );
  INV_X1 U30 ( .A(n878), .ZN(n813) );
  INV_X1 U31 ( .A(n869), .ZN(n812) );
  INV_X1 U32 ( .A(n860), .ZN(n811) );
  INV_X1 U33 ( .A(n851), .ZN(n810) );
  INV_X1 U34 ( .A(n987), .ZN(n828) );
  INV_X1 U35 ( .A(n978), .ZN(n827) );
  INV_X1 U36 ( .A(n969), .ZN(n826) );
  INV_X1 U37 ( .A(n914), .ZN(n820) );
  INV_X1 U38 ( .A(n905), .ZN(n819) );
  INV_X1 U39 ( .A(n896), .ZN(n818) );
  INV_X1 U40 ( .A(n1033), .ZN(n833) );
  INV_X1 U41 ( .A(n1023), .ZN(n832) );
  INV_X1 U42 ( .A(n1014), .ZN(n831) );
  INV_X1 U43 ( .A(n1005), .ZN(n830) );
  INV_X1 U44 ( .A(n996), .ZN(n829) );
  INV_X1 U45 ( .A(n960), .ZN(n825) );
  INV_X1 U46 ( .A(n950), .ZN(n824) );
  INV_X1 U47 ( .A(n941), .ZN(n823) );
  INV_X1 U48 ( .A(n932), .ZN(n822) );
  INV_X1 U49 ( .A(n923), .ZN(n821) );
  INV_X1 U50 ( .A(n1142), .ZN(n817) );
  BUF_X1 U51 ( .A(N11), .Z(n242) );
  BUF_X1 U52 ( .A(N11), .Z(n243) );
  BUF_X1 U53 ( .A(N11), .Z(n244) );
  INV_X1 U54 ( .A(N10), .ZN(n251) );
  BUF_X1 U55 ( .A(N12), .Z(n241) );
  NOR3_X1 U56 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U57 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U58 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U60 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U62 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U63 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U64 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U65 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U67 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U69 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U70 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U71 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U72 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U73 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U74 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U75 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U76 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U77 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U79 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U81 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U82 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U83 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U84 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U85 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U86 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U88 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U89 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U90 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U92 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U94 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U95 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U96 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U97 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U98 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U99 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U100 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U101 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U102 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U103 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U104 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U105 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U106 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U107 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U108 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U109 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U110 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U111 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U112 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U113 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U114 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U115 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U116 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U117 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U118 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U119 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U120 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U121 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U122 ( .A(n988), .ZN(n705) );
  AOI22_X1 U123 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U124 ( .A(n986), .ZN(n704) );
  AOI22_X1 U125 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U126 ( .A(n985), .ZN(n703) );
  AOI22_X1 U127 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U128 ( .A(n984), .ZN(n702) );
  AOI22_X1 U129 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U130 ( .A(n983), .ZN(n701) );
  AOI22_X1 U131 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U132 ( .A(n982), .ZN(n700) );
  AOI22_X1 U133 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U134 ( .A(n981), .ZN(n699) );
  AOI22_X1 U135 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U136 ( .A(n980), .ZN(n698) );
  AOI22_X1 U137 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U138 ( .A(n951), .ZN(n673) );
  AOI22_X1 U139 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U140 ( .A(n949), .ZN(n672) );
  AOI22_X1 U141 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U142 ( .A(n948), .ZN(n671) );
  AOI22_X1 U143 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U144 ( .A(n947), .ZN(n670) );
  AOI22_X1 U145 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U146 ( .A(n946), .ZN(n669) );
  AOI22_X1 U147 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U148 ( .A(n945), .ZN(n668) );
  AOI22_X1 U149 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U150 ( .A(n944), .ZN(n667) );
  AOI22_X1 U151 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U152 ( .A(n943), .ZN(n666) );
  AOI22_X1 U153 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U154 ( .A(n915), .ZN(n641) );
  AOI22_X1 U155 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U156 ( .A(n913), .ZN(n640) );
  AOI22_X1 U157 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U158 ( .A(n912), .ZN(n639) );
  AOI22_X1 U159 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U160 ( .A(n911), .ZN(n638) );
  AOI22_X1 U161 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U162 ( .A(n910), .ZN(n637) );
  AOI22_X1 U163 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U164 ( .A(n909), .ZN(n636) );
  AOI22_X1 U165 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U166 ( .A(n908), .ZN(n635) );
  AOI22_X1 U167 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U168 ( .A(n907), .ZN(n634) );
  AOI22_X1 U169 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U170 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U171 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U172 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U173 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U174 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U175 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U176 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U177 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U178 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U179 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U180 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U181 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U182 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U183 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U184 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U185 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U186 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U187 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U188 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U189 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U190 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U191 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U192 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U193 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U194 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U195 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U196 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U197 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U198 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U199 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U200 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U201 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U202 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U203 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U204 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U205 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U206 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U207 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U208 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U209 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U210 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U211 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U212 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U213 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U214 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U215 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U216 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U217 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U218 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U219 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U220 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U221 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U222 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U223 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U224 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U225 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U226 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U227 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U228 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U229 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U230 ( .A(n999), .ZN(n715) );
  AOI22_X1 U231 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U232 ( .A(n998), .ZN(n714) );
  AOI22_X1 U233 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U234 ( .A(n979), .ZN(n697) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U236 ( .A(n977), .ZN(n696) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U238 ( .A(n976), .ZN(n695) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U240 ( .A(n975), .ZN(n694) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U242 ( .A(n974), .ZN(n693) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U244 ( .A(n973), .ZN(n692) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U246 ( .A(n972), .ZN(n691) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U248 ( .A(n971), .ZN(n690) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U250 ( .A(n970), .ZN(n689) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U252 ( .A(n968), .ZN(n688) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U254 ( .A(n967), .ZN(n687) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U256 ( .A(n966), .ZN(n686) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U258 ( .A(n965), .ZN(n685) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U260 ( .A(n964), .ZN(n684) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U262 ( .A(n963), .ZN(n683) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U264 ( .A(n962), .ZN(n682) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U266 ( .A(n942), .ZN(n665) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U268 ( .A(n940), .ZN(n664) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U270 ( .A(n939), .ZN(n663) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U272 ( .A(n938), .ZN(n662) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U274 ( .A(n937), .ZN(n661) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U276 ( .A(n936), .ZN(n660) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U278 ( .A(n935), .ZN(n659) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U280 ( .A(n934), .ZN(n658) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U282 ( .A(n933), .ZN(n657) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U284 ( .A(n931), .ZN(n656) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U286 ( .A(n930), .ZN(n655) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U288 ( .A(n929), .ZN(n654) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U290 ( .A(n928), .ZN(n653) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U292 ( .A(n927), .ZN(n652) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U294 ( .A(n926), .ZN(n651) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U296 ( .A(n925), .ZN(n650) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U298 ( .A(n906), .ZN(n633) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U300 ( .A(n904), .ZN(n632) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U302 ( .A(n903), .ZN(n631) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U304 ( .A(n902), .ZN(n630) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U306 ( .A(n901), .ZN(n629) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U308 ( .A(n900), .ZN(n628) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U310 ( .A(n899), .ZN(n627) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U312 ( .A(n898), .ZN(n626) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U314 ( .A(n897), .ZN(n625) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U316 ( .A(n895), .ZN(n624) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U318 ( .A(n894), .ZN(n623) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U320 ( .A(n893), .ZN(n622) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U322 ( .A(n892), .ZN(n621) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U324 ( .A(n891), .ZN(n620) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U326 ( .A(n890), .ZN(n619) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U328 ( .A(n889), .ZN(n618) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U330 ( .A(N12), .ZN(n253) );
  INV_X1 U331 ( .A(N11), .ZN(n252) );
  INV_X1 U332 ( .A(n997), .ZN(n713) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U334 ( .A(n995), .ZN(n712) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U336 ( .A(n994), .ZN(n711) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U338 ( .A(n993), .ZN(n710) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U340 ( .A(n992), .ZN(n709) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U342 ( .A(n991), .ZN(n708) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U344 ( .A(n990), .ZN(n707) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U346 ( .A(n989), .ZN(n706) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U348 ( .A(n924), .ZN(n649) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U350 ( .A(n922), .ZN(n648) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U352 ( .A(n921), .ZN(n647) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U354 ( .A(n920), .ZN(n646) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U356 ( .A(n919), .ZN(n645) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U358 ( .A(n918), .ZN(n644) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U360 ( .A(n917), .ZN(n643) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U362 ( .A(n916), .ZN(n642) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U364 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U366 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U368 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U370 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U372 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U374 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U376 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U378 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U380 ( .A(n961), .ZN(n681) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U382 ( .A(n959), .ZN(n680) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U384 ( .A(n958), .ZN(n679) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U386 ( .A(n957), .ZN(n678) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U388 ( .A(n956), .ZN(n677) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U390 ( .A(n955), .ZN(n676) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U392 ( .A(n954), .ZN(n675) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U394 ( .A(n953), .ZN(n674) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U396 ( .A(n888), .ZN(n617) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U398 ( .A(n886), .ZN(n616) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U400 ( .A(n885), .ZN(n615) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U402 ( .A(n884), .ZN(n614) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U404 ( .A(n883), .ZN(n613) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U406 ( .A(n882), .ZN(n612) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U408 ( .A(n881), .ZN(n611) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U410 ( .A(n880), .ZN(n610) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U412 ( .A(n879), .ZN(n609) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U414 ( .A(n877), .ZN(n608) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U416 ( .A(n876), .ZN(n607) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U418 ( .A(n875), .ZN(n606) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U420 ( .A(n874), .ZN(n605) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U422 ( .A(n873), .ZN(n604) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U424 ( .A(n872), .ZN(n603) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U426 ( .A(n871), .ZN(n602) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U428 ( .A(n870), .ZN(n601) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U430 ( .A(n868), .ZN(n600) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U432 ( .A(n867), .ZN(n599) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U434 ( .A(n866), .ZN(n598) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U436 ( .A(n865), .ZN(n597) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U438 ( .A(n864), .ZN(n596) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U440 ( .A(n863), .ZN(n595) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U442 ( .A(n862), .ZN(n594) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U444 ( .A(n861), .ZN(n293) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U446 ( .A(n859), .ZN(n292) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U448 ( .A(n858), .ZN(n291) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U450 ( .A(n857), .ZN(n290) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U452 ( .A(n856), .ZN(n289) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U454 ( .A(n855), .ZN(n288) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U456 ( .A(n854), .ZN(n287) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U458 ( .A(n853), .ZN(n286) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U460 ( .A(n852), .ZN(n285) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U462 ( .A(n850), .ZN(n284) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U464 ( .A(n849), .ZN(n283) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U466 ( .A(n848), .ZN(n282) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U468 ( .A(n847), .ZN(n281) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U470 ( .A(n846), .ZN(n280) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U472 ( .A(n845), .ZN(n279) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U474 ( .A(n844), .ZN(n278) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U476 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U477 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U478 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U479 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U480 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U481 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U482 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U483 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U484 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U485 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U486 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U487 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U488 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U489 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U490 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U491 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U492 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U494 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U496 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U498 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U500 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U502 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U504 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U506 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U508 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U510 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U512 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U514 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U516 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U518 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U520 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U522 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U524 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U526 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U528 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U530 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U532 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U534 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U536 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U538 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U540 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U542 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U544 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U546 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U548 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U550 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U552 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U554 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U556 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U558 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U560 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U562 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U564 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U566 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U568 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U570 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U572 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U574 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U576 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U578 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U580 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U582 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U584 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U586 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U588 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U590 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U592 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U594 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U596 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U598 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U600 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U602 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U604 ( .A(N13), .ZN(n842) );
  INV_X1 U605 ( .A(N14), .ZN(n843) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n248), .Z(n1) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n248), .Z(n2) );
  MUX2_X1 U608 ( .A(n2), .B(n1), .S(n243), .Z(n3) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n248), .Z(n4) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n249), .Z(n5) );
  MUX2_X1 U611 ( .A(n5), .B(n4), .S(n244), .Z(n6) );
  MUX2_X1 U612 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n248), .Z(n8) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n249), .Z(n9) );
  MUX2_X1 U615 ( .A(n9), .B(n8), .S(n243), .Z(n10) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n248), .Z(n11) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n246), .Z(n12) );
  MUX2_X1 U618 ( .A(n12), .B(n11), .S(N11), .Z(n13) );
  MUX2_X1 U619 ( .A(n13), .B(n10), .S(n241), .Z(n14) );
  MUX2_X1 U620 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n245), .Z(n16) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n245), .Z(n17) );
  MUX2_X1 U623 ( .A(n17), .B(n16), .S(n242), .Z(n18) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n245), .Z(n20) );
  MUX2_X1 U626 ( .A(n20), .B(n19), .S(n243), .Z(n21) );
  MUX2_X1 U627 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n245), .Z(n23) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n245), .Z(n24) );
  MUX2_X1 U630 ( .A(n24), .B(n23), .S(N11), .Z(n25) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n245), .Z(n26) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n245), .Z(n27) );
  MUX2_X1 U633 ( .A(n27), .B(n26), .S(n244), .Z(n28) );
  MUX2_X1 U634 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U635 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U636 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n245), .Z(n31) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n245), .Z(n32) );
  MUX2_X1 U639 ( .A(n32), .B(n31), .S(N11), .Z(n33) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U642 ( .A(n35), .B(n34), .S(n242), .Z(n36) );
  MUX2_X1 U643 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n246), .Z(n38) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n246), .Z(n39) );
  MUX2_X1 U646 ( .A(n39), .B(n38), .S(N11), .Z(n40) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n246), .Z(n41) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n246), .Z(n42) );
  MUX2_X1 U649 ( .A(n42), .B(n41), .S(n242), .Z(n43) );
  MUX2_X1 U650 ( .A(n43), .B(n40), .S(n241), .Z(n44) );
  MUX2_X1 U651 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n246), .Z(n46) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n246), .Z(n47) );
  MUX2_X1 U654 ( .A(n47), .B(n46), .S(n244), .Z(n48) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n246), .Z(n49) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n246), .Z(n50) );
  MUX2_X1 U657 ( .A(n50), .B(n49), .S(n243), .Z(n51) );
  MUX2_X1 U658 ( .A(n51), .B(n48), .S(n241), .Z(n52) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n246), .Z(n53) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n246), .Z(n54) );
  MUX2_X1 U661 ( .A(n54), .B(n53), .S(N11), .Z(n55) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n246), .Z(n56) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n246), .Z(n57) );
  MUX2_X1 U664 ( .A(n57), .B(n56), .S(N11), .Z(n58) );
  MUX2_X1 U665 ( .A(n58), .B(n55), .S(n241), .Z(n59) );
  MUX2_X1 U666 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U667 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n247), .Z(n61) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n247), .Z(n62) );
  MUX2_X1 U670 ( .A(n62), .B(n61), .S(n242), .Z(n63) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n247), .Z(n64) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n247), .Z(n65) );
  MUX2_X1 U673 ( .A(n65), .B(n64), .S(n242), .Z(n66) );
  MUX2_X1 U674 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n247), .Z(n68) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n247), .Z(n69) );
  MUX2_X1 U677 ( .A(n69), .B(n68), .S(n242), .Z(n70) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n247), .Z(n71) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n247), .Z(n72) );
  MUX2_X1 U680 ( .A(n72), .B(n71), .S(n242), .Z(n73) );
  MUX2_X1 U681 ( .A(n73), .B(n70), .S(N12), .Z(n74) );
  MUX2_X1 U682 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n247), .Z(n76) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n247), .Z(n77) );
  MUX2_X1 U685 ( .A(n77), .B(n76), .S(n242), .Z(n78) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n247), .Z(n79) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n247), .Z(n80) );
  MUX2_X1 U688 ( .A(n80), .B(n79), .S(n242), .Z(n81) );
  MUX2_X1 U689 ( .A(n81), .B(n78), .S(N12), .Z(n82) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n249), .Z(n83) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n246), .Z(n84) );
  MUX2_X1 U692 ( .A(n84), .B(n83), .S(n242), .Z(n85) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n247), .Z(n86) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n245), .Z(n87) );
  MUX2_X1 U695 ( .A(n87), .B(n86), .S(n242), .Z(n88) );
  MUX2_X1 U696 ( .A(n88), .B(n85), .S(N12), .Z(n89) );
  MUX2_X1 U697 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U698 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n249), .Z(n91) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n246), .Z(n92) );
  MUX2_X1 U701 ( .A(n92), .B(n91), .S(n242), .Z(n93) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n245), .Z(n94) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n245), .Z(n95) );
  MUX2_X1 U704 ( .A(n95), .B(n94), .S(n242), .Z(n96) );
  MUX2_X1 U705 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n98) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n249), .Z(n99) );
  MUX2_X1 U708 ( .A(n99), .B(n98), .S(n242), .Z(n100) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n247), .Z(n101) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n247), .Z(n102) );
  MUX2_X1 U711 ( .A(n102), .B(n101), .S(n242), .Z(n103) );
  MUX2_X1 U712 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U713 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n248), .Z(n106) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(N10), .Z(n107) );
  MUX2_X1 U716 ( .A(n107), .B(n106), .S(n243), .Z(n108) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n248), .Z(n109) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n250), .Z(n110) );
  MUX2_X1 U719 ( .A(n110), .B(n109), .S(n243), .Z(n111) );
  MUX2_X1 U720 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n248), .Z(n113) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n114) );
  MUX2_X1 U723 ( .A(n114), .B(n113), .S(n243), .Z(n115) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n250), .Z(n116) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n117) );
  MUX2_X1 U726 ( .A(n117), .B(n116), .S(n243), .Z(n118) );
  MUX2_X1 U727 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U728 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U729 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(N10), .Z(n121) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(N10), .Z(n122) );
  MUX2_X1 U732 ( .A(n122), .B(n121), .S(n243), .Z(n123) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(N10), .Z(n124) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n125) );
  MUX2_X1 U735 ( .A(n125), .B(n124), .S(n243), .Z(n126) );
  MUX2_X1 U736 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n248), .Z(n128) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n248), .Z(n129) );
  MUX2_X1 U739 ( .A(n129), .B(n128), .S(n243), .Z(n130) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n248), .Z(n131) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n248), .Z(n132) );
  MUX2_X1 U742 ( .A(n132), .B(n131), .S(n243), .Z(n133) );
  MUX2_X1 U743 ( .A(n133), .B(n130), .S(N12), .Z(n134) );
  MUX2_X1 U744 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n248), .Z(n136) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n248), .Z(n137) );
  MUX2_X1 U747 ( .A(n137), .B(n136), .S(n243), .Z(n138) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n248), .Z(n139) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n248), .Z(n140) );
  MUX2_X1 U750 ( .A(n140), .B(n139), .S(n243), .Z(n141) );
  MUX2_X1 U751 ( .A(n141), .B(n138), .S(N12), .Z(n142) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n248), .Z(n143) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n248), .Z(n144) );
  MUX2_X1 U754 ( .A(n144), .B(n143), .S(n243), .Z(n145) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n248), .Z(n146) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n248), .Z(n147) );
  MUX2_X1 U757 ( .A(n147), .B(n146), .S(n243), .Z(n148) );
  MUX2_X1 U758 ( .A(n148), .B(n145), .S(N12), .Z(n149) );
  MUX2_X1 U759 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U760 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n249), .Z(n151) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n249), .Z(n152) );
  MUX2_X1 U763 ( .A(n152), .B(n151), .S(n244), .Z(n153) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n249), .Z(n154) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n249), .Z(n155) );
  MUX2_X1 U766 ( .A(n155), .B(n154), .S(n244), .Z(n156) );
  MUX2_X1 U767 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n249), .Z(n158) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n249), .Z(n159) );
  MUX2_X1 U770 ( .A(n159), .B(n158), .S(n244), .Z(n160) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n249), .Z(n161) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n249), .Z(n162) );
  MUX2_X1 U773 ( .A(n162), .B(n161), .S(n244), .Z(n163) );
  MUX2_X1 U774 ( .A(n163), .B(n160), .S(n241), .Z(n164) );
  MUX2_X1 U775 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n249), .Z(n166) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n249), .Z(n167) );
  MUX2_X1 U778 ( .A(n167), .B(n166), .S(n244), .Z(n168) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n249), .Z(n169) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n249), .Z(n170) );
  MUX2_X1 U781 ( .A(n170), .B(n169), .S(n244), .Z(n171) );
  MUX2_X1 U782 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n248), .Z(n173) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n245), .Z(n174) );
  MUX2_X1 U785 ( .A(n174), .B(n173), .S(n244), .Z(n175) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n250), .Z(n176) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n246), .Z(n177) );
  MUX2_X1 U788 ( .A(n177), .B(n176), .S(n244), .Z(n178) );
  MUX2_X1 U789 ( .A(n178), .B(n175), .S(n241), .Z(n179) );
  MUX2_X1 U790 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U791 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n247), .Z(n181) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n248), .Z(n182) );
  MUX2_X1 U794 ( .A(n182), .B(n181), .S(n244), .Z(n183) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n246), .Z(n184) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n250), .Z(n185) );
  MUX2_X1 U797 ( .A(n185), .B(n184), .S(n244), .Z(n186) );
  MUX2_X1 U798 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n250), .Z(n188) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n250), .Z(n189) );
  MUX2_X1 U801 ( .A(n189), .B(n188), .S(n244), .Z(n190) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n250), .Z(n191) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n250), .Z(n192) );
  MUX2_X1 U804 ( .A(n192), .B(n191), .S(n244), .Z(n193) );
  MUX2_X1 U805 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U806 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n250), .Z(n196) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n250), .Z(n197) );
  MUX2_X1 U809 ( .A(n197), .B(n196), .S(N11), .Z(n198) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n250), .Z(n199) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n250), .Z(n200) );
  MUX2_X1 U812 ( .A(n200), .B(n199), .S(n242), .Z(n201) );
  MUX2_X1 U813 ( .A(n201), .B(n198), .S(N12), .Z(n202) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n250), .Z(n203) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n247), .Z(n204) );
  MUX2_X1 U816 ( .A(n204), .B(n203), .S(N11), .Z(n205) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n250), .Z(n206) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n250), .Z(n207) );
  MUX2_X1 U819 ( .A(n207), .B(n206), .S(n242), .Z(n208) );
  MUX2_X1 U820 ( .A(n208), .B(n205), .S(N12), .Z(n209) );
  MUX2_X1 U821 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U822 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n250), .Z(n211) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n245), .Z(n212) );
  MUX2_X1 U825 ( .A(n212), .B(n211), .S(N11), .Z(n213) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n248), .Z(n214) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n250), .Z(n215) );
  MUX2_X1 U828 ( .A(n215), .B(n214), .S(N11), .Z(n216) );
  MUX2_X1 U829 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n245), .Z(n218) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(N10), .Z(n219) );
  MUX2_X1 U832 ( .A(n219), .B(n218), .S(N11), .Z(n220) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n250), .Z(n221) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n222) );
  MUX2_X1 U835 ( .A(n222), .B(n221), .S(n243), .Z(n223) );
  MUX2_X1 U836 ( .A(n223), .B(n220), .S(n241), .Z(n224) );
  MUX2_X1 U837 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n250), .Z(n226) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n227) );
  MUX2_X1 U840 ( .A(n227), .B(n226), .S(N11), .Z(n228) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n246), .Z(n229) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n230) );
  MUX2_X1 U843 ( .A(n230), .B(n229), .S(n244), .Z(n231) );
  MUX2_X1 U844 ( .A(n231), .B(n228), .S(n241), .Z(n232) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n247), .Z(n233) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n234) );
  MUX2_X1 U847 ( .A(n234), .B(n233), .S(N11), .Z(n235) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n236) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n237) );
  MUX2_X1 U850 ( .A(n237), .B(n236), .S(n244), .Z(n238) );
  MUX2_X1 U851 ( .A(n238), .B(n235), .S(n241), .Z(n239) );
  MUX2_X1 U852 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U853 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_25 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n256), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n257), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n258), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n259), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n260), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n261), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n262), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n263), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n264), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n265), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n266), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n267), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n268), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n269), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n270), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n271), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n272), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n273), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n274), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n275), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n276), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n277), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n278), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n279), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n280), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n281), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n282), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n283), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n284), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n285), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n286), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n287), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n288), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n289), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n290), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n291), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n292), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n293), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n594), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n595), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n596), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n597), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n598), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n599), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n600), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n601), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n602), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n603), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n604), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n605), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n606), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n607), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n608), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n609), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n610), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n611), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n612), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n613), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n614), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n615), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n616), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n617), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n618), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n619), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n620), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n621), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n622), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n623), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n624), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n625), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n626), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n627), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n628), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n629), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n630), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n631), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n632), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n633), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n634), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n635), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n636), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n637), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n638), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n639), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n640), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n641), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n642), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n643), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n644), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n645), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n646), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n647), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n648), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n649), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n650), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n651), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n652), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n653), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n654), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n655), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n656), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n657), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n658), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n659), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n660), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n661), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n662), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n663), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n664), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n665), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n666), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n667), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n668), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n669), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n670), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n671), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n672), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n673), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n674), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n675), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n676), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n677), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n678), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n679), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n680), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n681), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n682), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n683), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n684), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n685), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n686), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n687), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n688), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n689), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n690), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n691), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n692), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n693), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n694), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n695), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n696), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n697), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n698), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n699), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n700), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n701), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n702), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n703), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n704), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n705), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n706), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n707), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n708), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n709), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n710), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n711), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n712), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n713), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n714), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n715), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n716), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n717), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n718), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n719), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n720), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n721), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n722), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n723), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n724), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n725), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n726), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n727), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n728), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n729), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n730), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n731), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n732), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n733), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n734), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n735), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n736), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n737), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n738), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n739), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n740), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n741), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n742), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n743), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n744), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n745), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n746), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n747), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n748), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n749), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n750), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n751), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n752), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n753), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n754), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n755), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n756), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n757), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n758), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n759), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n760), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n761), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n762), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n763), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n764), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n765), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n766), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n767), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n768), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n769), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n770), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n771), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n772), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n773), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n774), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n775), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n776), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n777), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n778), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n779), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n780), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n781), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n782), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n783), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n784), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n785), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n786), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n787), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n788), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n789), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n790), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n791), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n792), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n793), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n794), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n795), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n796), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n797), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n798), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n799), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n800), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n801), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n802), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n803), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n804), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n805), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n806), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n807), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n808), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n809), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n810), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n811), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  DFF_X2 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(n252), .Z(n250) );
  BUF_X1 U5 ( .A(N10), .Z(n251) );
  BUF_X1 U6 ( .A(n252), .Z(n247) );
  BUF_X1 U7 ( .A(n252), .Z(n248) );
  BUF_X1 U8 ( .A(n252), .Z(n249) );
  BUF_X1 U9 ( .A(N10), .Z(n252) );
  INV_X1 U10 ( .A(n1113), .ZN(n843) );
  INV_X1 U11 ( .A(n1102), .ZN(n842) );
  INV_X1 U12 ( .A(n1092), .ZN(n841) );
  INV_X1 U13 ( .A(n1082), .ZN(n840) );
  INV_X1 U14 ( .A(n1072), .ZN(n839) );
  INV_X1 U15 ( .A(n1062), .ZN(n838) );
  INV_X1 U16 ( .A(n1053), .ZN(n837) );
  INV_X1 U17 ( .A(n1044), .ZN(n836) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1105) );
  NOR3_X1 U19 ( .A1(N11), .A2(N12), .A3(n253), .ZN(n1094) );
  NAND2_X1 U20 ( .A1(n1104), .A2(n1136), .ZN(n1062) );
  NAND2_X1 U21 ( .A1(n1105), .A2(n1104), .ZN(n1113) );
  NAND2_X1 U22 ( .A1(n1094), .A2(n1104), .ZN(n1102) );
  NAND2_X1 U23 ( .A1(n1084), .A2(n1104), .ZN(n1092) );
  NAND2_X1 U24 ( .A1(n1074), .A2(n1104), .ZN(n1082) );
  NAND2_X1 U25 ( .A1(n1064), .A2(n1104), .ZN(n1072) );
  NAND2_X1 U26 ( .A1(n1104), .A2(n1125), .ZN(n1053) );
  NAND2_X1 U27 ( .A1(n1104), .A2(n1115), .ZN(n1044) );
  INV_X1 U28 ( .A(n1133), .ZN(n818) );
  INV_X1 U29 ( .A(n1123), .ZN(n817) );
  INV_X1 U30 ( .A(n889), .ZN(n816) );
  INV_X1 U31 ( .A(n880), .ZN(n815) );
  INV_X1 U32 ( .A(n871), .ZN(n814) );
  INV_X1 U33 ( .A(n862), .ZN(n813) );
  INV_X1 U34 ( .A(n853), .ZN(n812) );
  INV_X1 U35 ( .A(n989), .ZN(n830) );
  INV_X1 U36 ( .A(n980), .ZN(n829) );
  INV_X1 U37 ( .A(n971), .ZN(n828) );
  INV_X1 U38 ( .A(n916), .ZN(n822) );
  INV_X1 U39 ( .A(n907), .ZN(n821) );
  INV_X1 U40 ( .A(n898), .ZN(n820) );
  INV_X1 U41 ( .A(n1035), .ZN(n835) );
  INV_X1 U42 ( .A(n1025), .ZN(n834) );
  INV_X1 U43 ( .A(n1016), .ZN(n833) );
  INV_X1 U44 ( .A(n1007), .ZN(n832) );
  INV_X1 U45 ( .A(n998), .ZN(n831) );
  INV_X1 U46 ( .A(n962), .ZN(n827) );
  INV_X1 U47 ( .A(n952), .ZN(n826) );
  INV_X1 U48 ( .A(n943), .ZN(n825) );
  INV_X1 U49 ( .A(n934), .ZN(n824) );
  INV_X1 U50 ( .A(n925), .ZN(n823) );
  INV_X1 U51 ( .A(n1144), .ZN(n819) );
  BUF_X1 U52 ( .A(N11), .Z(n245) );
  BUF_X1 U53 ( .A(N11), .Z(n246) );
  INV_X1 U54 ( .A(N10), .ZN(n253) );
  BUF_X1 U55 ( .A(N12), .Z(n243) );
  NOR3_X1 U56 ( .A1(n255), .A2(N10), .A3(n254), .ZN(n1125) );
  NOR3_X1 U57 ( .A1(n255), .A2(n253), .A3(n254), .ZN(n1115) );
  NOR3_X1 U58 ( .A1(n253), .A2(N11), .A3(n255), .ZN(n1136) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n254), .ZN(n1084) );
  NOR3_X1 U60 ( .A1(n253), .A2(N12), .A3(n254), .ZN(n1074) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n255), .ZN(n1064) );
  NAND2_X1 U62 ( .A1(n1027), .A2(n1136), .ZN(n989) );
  NAND2_X1 U63 ( .A1(n954), .A2(n1136), .ZN(n916) );
  NAND2_X1 U64 ( .A1(n1027), .A2(n1064), .ZN(n998) );
  NAND2_X1 U65 ( .A1(n954), .A2(n1064), .ZN(n925) );
  NAND2_X1 U66 ( .A1(n1027), .A2(n1105), .ZN(n1035) );
  NAND2_X1 U67 ( .A1(n1027), .A2(n1094), .ZN(n1025) );
  NAND2_X1 U68 ( .A1(n954), .A2(n1105), .ZN(n962) );
  NAND2_X1 U69 ( .A1(n954), .A2(n1094), .ZN(n952) );
  NAND2_X1 U70 ( .A1(n1105), .A2(n1135), .ZN(n889) );
  NAND2_X1 U71 ( .A1(n1094), .A2(n1135), .ZN(n880) );
  NAND2_X1 U72 ( .A1(n1084), .A2(n1135), .ZN(n871) );
  NAND2_X1 U73 ( .A1(n1074), .A2(n1135), .ZN(n862) );
  NAND2_X1 U74 ( .A1(n1064), .A2(n1135), .ZN(n853) );
  NAND2_X1 U75 ( .A1(n1136), .A2(n1135), .ZN(n1144) );
  NAND2_X1 U76 ( .A1(n1125), .A2(n1135), .ZN(n1133) );
  NAND2_X1 U77 ( .A1(n1115), .A2(n1135), .ZN(n1123) );
  NAND2_X1 U78 ( .A1(n1027), .A2(n1084), .ZN(n1016) );
  NAND2_X1 U79 ( .A1(n1027), .A2(n1074), .ZN(n1007) );
  NAND2_X1 U80 ( .A1(n954), .A2(n1084), .ZN(n943) );
  NAND2_X1 U81 ( .A1(n954), .A2(n1074), .ZN(n934) );
  NAND2_X1 U82 ( .A1(n1027), .A2(n1125), .ZN(n980) );
  NAND2_X1 U83 ( .A1(n954), .A2(n1125), .ZN(n907) );
  NAND2_X1 U84 ( .A1(n1027), .A2(n1115), .ZN(n971) );
  NAND2_X1 U85 ( .A1(n954), .A2(n1115), .ZN(n898) );
  AND3_X1 U86 ( .A1(n844), .A2(n845), .A3(wr_en), .ZN(n1104) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1135) );
  AND3_X1 U88 ( .A1(N13), .A2(n845), .A3(wr_en), .ZN(n1027) );
  AND3_X1 U89 ( .A1(N14), .A2(n844), .A3(wr_en), .ZN(n954) );
  INV_X1 U90 ( .A(n1063), .ZN(n771) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n838), .B1(n1062), .B2(\mem[5][0] ), 
        .ZN(n1063) );
  INV_X1 U92 ( .A(n1061), .ZN(n770) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n838), .B1(n1062), .B2(\mem[5][1] ), 
        .ZN(n1061) );
  INV_X1 U94 ( .A(n1060), .ZN(n769) );
  AOI22_X1 U95 ( .A1(data_in[2]), .A2(n838), .B1(n1062), .B2(\mem[5][2] ), 
        .ZN(n1060) );
  INV_X1 U96 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U97 ( .A1(data_in[3]), .A2(n838), .B1(n1062), .B2(\mem[5][3] ), 
        .ZN(n1059) );
  INV_X1 U98 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U99 ( .A1(data_in[4]), .A2(n838), .B1(n1062), .B2(\mem[5][4] ), 
        .ZN(n1058) );
  INV_X1 U100 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U101 ( .A1(data_in[5]), .A2(n838), .B1(n1062), .B2(\mem[5][5] ), 
        .ZN(n1057) );
  INV_X1 U102 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U103 ( .A1(data_in[6]), .A2(n838), .B1(n1062), .B2(\mem[5][6] ), 
        .ZN(n1056) );
  INV_X1 U104 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U105 ( .A1(data_in[7]), .A2(n838), .B1(n1062), .B2(\mem[5][7] ), 
        .ZN(n1055) );
  INV_X1 U106 ( .A(n1026), .ZN(n739) );
  AOI22_X1 U107 ( .A1(data_in[0]), .A2(n834), .B1(n1025), .B2(\mem[9][0] ), 
        .ZN(n1026) );
  INV_X1 U108 ( .A(n1024), .ZN(n738) );
  AOI22_X1 U109 ( .A1(data_in[1]), .A2(n834), .B1(n1025), .B2(\mem[9][1] ), 
        .ZN(n1024) );
  INV_X1 U110 ( .A(n1023), .ZN(n737) );
  AOI22_X1 U111 ( .A1(data_in[2]), .A2(n834), .B1(n1025), .B2(\mem[9][2] ), 
        .ZN(n1023) );
  INV_X1 U112 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U113 ( .A1(data_in[3]), .A2(n834), .B1(n1025), .B2(\mem[9][3] ), 
        .ZN(n1022) );
  INV_X1 U114 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U115 ( .A1(data_in[4]), .A2(n834), .B1(n1025), .B2(\mem[9][4] ), 
        .ZN(n1021) );
  INV_X1 U116 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U117 ( .A1(data_in[5]), .A2(n834), .B1(n1025), .B2(\mem[9][5] ), 
        .ZN(n1020) );
  INV_X1 U118 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U119 ( .A1(data_in[6]), .A2(n834), .B1(n1025), .B2(\mem[9][6] ), 
        .ZN(n1019) );
  INV_X1 U120 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U121 ( .A1(data_in[7]), .A2(n834), .B1(n1025), .B2(\mem[9][7] ), 
        .ZN(n1018) );
  INV_X1 U122 ( .A(n990), .ZN(n707) );
  AOI22_X1 U123 ( .A1(data_in[0]), .A2(n830), .B1(n989), .B2(\mem[13][0] ), 
        .ZN(n990) );
  INV_X1 U124 ( .A(n988), .ZN(n706) );
  AOI22_X1 U125 ( .A1(data_in[1]), .A2(n830), .B1(n989), .B2(\mem[13][1] ), 
        .ZN(n988) );
  INV_X1 U126 ( .A(n987), .ZN(n705) );
  AOI22_X1 U127 ( .A1(data_in[2]), .A2(n830), .B1(n989), .B2(\mem[13][2] ), 
        .ZN(n987) );
  INV_X1 U128 ( .A(n986), .ZN(n704) );
  AOI22_X1 U129 ( .A1(data_in[3]), .A2(n830), .B1(n989), .B2(\mem[13][3] ), 
        .ZN(n986) );
  INV_X1 U130 ( .A(n985), .ZN(n703) );
  AOI22_X1 U131 ( .A1(data_in[4]), .A2(n830), .B1(n989), .B2(\mem[13][4] ), 
        .ZN(n985) );
  INV_X1 U132 ( .A(n984), .ZN(n702) );
  AOI22_X1 U133 ( .A1(data_in[5]), .A2(n830), .B1(n989), .B2(\mem[13][5] ), 
        .ZN(n984) );
  INV_X1 U134 ( .A(n983), .ZN(n701) );
  AOI22_X1 U135 ( .A1(data_in[6]), .A2(n830), .B1(n989), .B2(\mem[13][6] ), 
        .ZN(n983) );
  INV_X1 U136 ( .A(n982), .ZN(n700) );
  AOI22_X1 U137 ( .A1(data_in[7]), .A2(n830), .B1(n989), .B2(\mem[13][7] ), 
        .ZN(n982) );
  INV_X1 U138 ( .A(n913), .ZN(n640) );
  AOI22_X1 U139 ( .A1(data_in[3]), .A2(n822), .B1(n916), .B2(\mem[21][3] ), 
        .ZN(n913) );
  INV_X1 U140 ( .A(n912), .ZN(n639) );
  AOI22_X1 U141 ( .A1(data_in[4]), .A2(n822), .B1(n916), .B2(\mem[21][4] ), 
        .ZN(n912) );
  INV_X1 U142 ( .A(n911), .ZN(n638) );
  AOI22_X1 U143 ( .A1(data_in[5]), .A2(n822), .B1(n916), .B2(\mem[21][5] ), 
        .ZN(n911) );
  INV_X1 U144 ( .A(n910), .ZN(n637) );
  AOI22_X1 U145 ( .A1(data_in[6]), .A2(n822), .B1(n916), .B2(\mem[21][6] ), 
        .ZN(n910) );
  INV_X1 U146 ( .A(n909), .ZN(n636) );
  AOI22_X1 U147 ( .A1(data_in[7]), .A2(n822), .B1(n916), .B2(\mem[21][7] ), 
        .ZN(n909) );
  INV_X1 U148 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U149 ( .A1(data_in[0]), .A2(n833), .B1(n1016), .B2(\mem[10][0] ), 
        .ZN(n1017) );
  INV_X1 U150 ( .A(n1015), .ZN(n730) );
  AOI22_X1 U151 ( .A1(data_in[1]), .A2(n833), .B1(n1016), .B2(\mem[10][1] ), 
        .ZN(n1015) );
  INV_X1 U152 ( .A(n1014), .ZN(n729) );
  AOI22_X1 U153 ( .A1(data_in[2]), .A2(n833), .B1(n1016), .B2(\mem[10][2] ), 
        .ZN(n1014) );
  INV_X1 U154 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U155 ( .A1(data_in[3]), .A2(n833), .B1(n1016), .B2(\mem[10][3] ), 
        .ZN(n1013) );
  INV_X1 U156 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U157 ( .A1(data_in[4]), .A2(n833), .B1(n1016), .B2(\mem[10][4] ), 
        .ZN(n1012) );
  INV_X1 U158 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U159 ( .A1(data_in[5]), .A2(n833), .B1(n1016), .B2(\mem[10][5] ), 
        .ZN(n1011) );
  INV_X1 U160 ( .A(n953), .ZN(n675) );
  AOI22_X1 U161 ( .A1(data_in[0]), .A2(n826), .B1(n952), .B2(\mem[17][0] ), 
        .ZN(n953) );
  INV_X1 U162 ( .A(n951), .ZN(n674) );
  AOI22_X1 U163 ( .A1(data_in[1]), .A2(n826), .B1(n952), .B2(\mem[17][1] ), 
        .ZN(n951) );
  INV_X1 U164 ( .A(n950), .ZN(n673) );
  AOI22_X1 U165 ( .A1(data_in[2]), .A2(n826), .B1(n952), .B2(\mem[17][2] ), 
        .ZN(n950) );
  INV_X1 U166 ( .A(n949), .ZN(n672) );
  AOI22_X1 U167 ( .A1(data_in[3]), .A2(n826), .B1(n952), .B2(\mem[17][3] ), 
        .ZN(n949) );
  INV_X1 U168 ( .A(n948), .ZN(n671) );
  AOI22_X1 U169 ( .A1(data_in[4]), .A2(n826), .B1(n952), .B2(\mem[17][4] ), 
        .ZN(n948) );
  INV_X1 U170 ( .A(n947), .ZN(n670) );
  AOI22_X1 U171 ( .A1(data_in[5]), .A2(n826), .B1(n952), .B2(\mem[17][5] ), 
        .ZN(n947) );
  INV_X1 U172 ( .A(n946), .ZN(n669) );
  AOI22_X1 U173 ( .A1(data_in[6]), .A2(n826), .B1(n952), .B2(\mem[17][6] ), 
        .ZN(n946) );
  INV_X1 U174 ( .A(n945), .ZN(n668) );
  AOI22_X1 U175 ( .A1(data_in[7]), .A2(n826), .B1(n952), .B2(\mem[17][7] ), 
        .ZN(n945) );
  INV_X1 U176 ( .A(n917), .ZN(n643) );
  AOI22_X1 U177 ( .A1(data_in[0]), .A2(n822), .B1(n916), .B2(\mem[21][0] ), 
        .ZN(n917) );
  INV_X1 U178 ( .A(n915), .ZN(n642) );
  AOI22_X1 U179 ( .A1(data_in[1]), .A2(n822), .B1(n916), .B2(\mem[21][1] ), 
        .ZN(n915) );
  INV_X1 U180 ( .A(n914), .ZN(n641) );
  AOI22_X1 U181 ( .A1(data_in[2]), .A2(n822), .B1(n916), .B2(\mem[21][2] ), 
        .ZN(n914) );
  INV_X1 U182 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U183 ( .A1(data_in[0]), .A2(n837), .B1(n1053), .B2(\mem[6][0] ), 
        .ZN(n1054) );
  INV_X1 U184 ( .A(n1052), .ZN(n762) );
  AOI22_X1 U185 ( .A1(data_in[1]), .A2(n837), .B1(n1053), .B2(\mem[6][1] ), 
        .ZN(n1052) );
  INV_X1 U186 ( .A(n1051), .ZN(n761) );
  AOI22_X1 U187 ( .A1(data_in[2]), .A2(n837), .B1(n1053), .B2(\mem[6][2] ), 
        .ZN(n1051) );
  INV_X1 U188 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U189 ( .A1(data_in[3]), .A2(n837), .B1(n1053), .B2(\mem[6][3] ), 
        .ZN(n1050) );
  INV_X1 U190 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U191 ( .A1(data_in[4]), .A2(n837), .B1(n1053), .B2(\mem[6][4] ), 
        .ZN(n1049) );
  INV_X1 U192 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U193 ( .A1(data_in[5]), .A2(n837), .B1(n1053), .B2(\mem[6][5] ), 
        .ZN(n1048) );
  INV_X1 U194 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U195 ( .A1(data_in[6]), .A2(n837), .B1(n1053), .B2(\mem[6][6] ), 
        .ZN(n1047) );
  INV_X1 U196 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U197 ( .A1(data_in[7]), .A2(n837), .B1(n1053), .B2(\mem[6][7] ), 
        .ZN(n1046) );
  INV_X1 U198 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U199 ( .A1(data_in[0]), .A2(n836), .B1(n1044), .B2(\mem[7][0] ), 
        .ZN(n1045) );
  INV_X1 U200 ( .A(n1043), .ZN(n754) );
  AOI22_X1 U201 ( .A1(data_in[1]), .A2(n836), .B1(n1044), .B2(\mem[7][1] ), 
        .ZN(n1043) );
  INV_X1 U202 ( .A(n1042), .ZN(n753) );
  AOI22_X1 U203 ( .A1(data_in[2]), .A2(n836), .B1(n1044), .B2(\mem[7][2] ), 
        .ZN(n1042) );
  INV_X1 U204 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U205 ( .A1(data_in[3]), .A2(n836), .B1(n1044), .B2(\mem[7][3] ), 
        .ZN(n1041) );
  INV_X1 U206 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U207 ( .A1(data_in[4]), .A2(n836), .B1(n1044), .B2(\mem[7][4] ), 
        .ZN(n1040) );
  INV_X1 U208 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U209 ( .A1(data_in[5]), .A2(n836), .B1(n1044), .B2(\mem[7][5] ), 
        .ZN(n1039) );
  INV_X1 U210 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U211 ( .A1(data_in[6]), .A2(n836), .B1(n1044), .B2(\mem[7][6] ), 
        .ZN(n1038) );
  INV_X1 U212 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U213 ( .A1(data_in[7]), .A2(n836), .B1(n1044), .B2(\mem[7][7] ), 
        .ZN(n1037) );
  INV_X1 U214 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U215 ( .A1(data_in[6]), .A2(n833), .B1(n1016), .B2(\mem[10][6] ), 
        .ZN(n1010) );
  INV_X1 U216 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U217 ( .A1(data_in[7]), .A2(n833), .B1(n1016), .B2(\mem[10][7] ), 
        .ZN(n1009) );
  INV_X1 U218 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U219 ( .A1(data_in[0]), .A2(n832), .B1(n1007), .B2(\mem[11][0] ), 
        .ZN(n1008) );
  INV_X1 U220 ( .A(n1006), .ZN(n722) );
  AOI22_X1 U221 ( .A1(data_in[1]), .A2(n832), .B1(n1007), .B2(\mem[11][1] ), 
        .ZN(n1006) );
  INV_X1 U222 ( .A(n1005), .ZN(n721) );
  AOI22_X1 U223 ( .A1(data_in[2]), .A2(n832), .B1(n1007), .B2(\mem[11][2] ), 
        .ZN(n1005) );
  INV_X1 U224 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U225 ( .A1(data_in[3]), .A2(n832), .B1(n1007), .B2(\mem[11][3] ), 
        .ZN(n1004) );
  INV_X1 U226 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U227 ( .A1(data_in[4]), .A2(n832), .B1(n1007), .B2(\mem[11][4] ), 
        .ZN(n1003) );
  INV_X1 U228 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U229 ( .A1(data_in[5]), .A2(n832), .B1(n1007), .B2(\mem[11][5] ), 
        .ZN(n1002) );
  INV_X1 U230 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U231 ( .A1(data_in[6]), .A2(n832), .B1(n1007), .B2(\mem[11][6] ), 
        .ZN(n1001) );
  INV_X1 U232 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U233 ( .A1(data_in[7]), .A2(n832), .B1(n1007), .B2(\mem[11][7] ), 
        .ZN(n1000) );
  INV_X1 U234 ( .A(n981), .ZN(n699) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n829), .B1(n980), .B2(\mem[14][0] ), 
        .ZN(n981) );
  INV_X1 U236 ( .A(n979), .ZN(n698) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n829), .B1(n980), .B2(\mem[14][1] ), 
        .ZN(n979) );
  INV_X1 U238 ( .A(n978), .ZN(n697) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n829), .B1(n980), .B2(\mem[14][2] ), 
        .ZN(n978) );
  INV_X1 U240 ( .A(n977), .ZN(n696) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n829), .B1(n980), .B2(\mem[14][3] ), 
        .ZN(n977) );
  INV_X1 U242 ( .A(n976), .ZN(n695) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n829), .B1(n980), .B2(\mem[14][4] ), 
        .ZN(n976) );
  INV_X1 U244 ( .A(n975), .ZN(n694) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n829), .B1(n980), .B2(\mem[14][5] ), 
        .ZN(n975) );
  INV_X1 U246 ( .A(n974), .ZN(n693) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n829), .B1(n980), .B2(\mem[14][6] ), 
        .ZN(n974) );
  INV_X1 U248 ( .A(n973), .ZN(n692) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n829), .B1(n980), .B2(\mem[14][7] ), 
        .ZN(n973) );
  INV_X1 U250 ( .A(n972), .ZN(n691) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n828), .B1(n971), .B2(\mem[15][0] ), 
        .ZN(n972) );
  INV_X1 U252 ( .A(n970), .ZN(n690) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n828), .B1(n971), .B2(\mem[15][1] ), 
        .ZN(n970) );
  INV_X1 U254 ( .A(n969), .ZN(n689) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n828), .B1(n971), .B2(\mem[15][2] ), 
        .ZN(n969) );
  INV_X1 U256 ( .A(n968), .ZN(n688) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n828), .B1(n971), .B2(\mem[15][3] ), 
        .ZN(n968) );
  INV_X1 U258 ( .A(n967), .ZN(n687) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n828), .B1(n971), .B2(\mem[15][4] ), 
        .ZN(n967) );
  INV_X1 U260 ( .A(n966), .ZN(n686) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n828), .B1(n971), .B2(\mem[15][5] ), 
        .ZN(n966) );
  INV_X1 U262 ( .A(n965), .ZN(n685) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n828), .B1(n971), .B2(\mem[15][6] ), 
        .ZN(n965) );
  INV_X1 U264 ( .A(n964), .ZN(n684) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n828), .B1(n971), .B2(\mem[15][7] ), 
        .ZN(n964) );
  INV_X1 U266 ( .A(n944), .ZN(n667) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n825), .B1(n943), .B2(\mem[18][0] ), 
        .ZN(n944) );
  INV_X1 U268 ( .A(n942), .ZN(n666) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n825), .B1(n943), .B2(\mem[18][1] ), 
        .ZN(n942) );
  INV_X1 U270 ( .A(n941), .ZN(n665) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n825), .B1(n943), .B2(\mem[18][2] ), 
        .ZN(n941) );
  INV_X1 U272 ( .A(n940), .ZN(n664) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n825), .B1(n943), .B2(\mem[18][3] ), 
        .ZN(n940) );
  INV_X1 U274 ( .A(n939), .ZN(n663) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n825), .B1(n943), .B2(\mem[18][4] ), 
        .ZN(n939) );
  INV_X1 U276 ( .A(n938), .ZN(n662) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n825), .B1(n943), .B2(\mem[18][5] ), 
        .ZN(n938) );
  INV_X1 U278 ( .A(n937), .ZN(n661) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n825), .B1(n943), .B2(\mem[18][6] ), 
        .ZN(n937) );
  INV_X1 U280 ( .A(n936), .ZN(n660) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n825), .B1(n943), .B2(\mem[18][7] ), 
        .ZN(n936) );
  INV_X1 U282 ( .A(n935), .ZN(n659) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n824), .B1(n934), .B2(\mem[19][0] ), 
        .ZN(n935) );
  INV_X1 U284 ( .A(n933), .ZN(n658) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n824), .B1(n934), .B2(\mem[19][1] ), 
        .ZN(n933) );
  INV_X1 U286 ( .A(n932), .ZN(n657) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n824), .B1(n934), .B2(\mem[19][2] ), 
        .ZN(n932) );
  INV_X1 U288 ( .A(n931), .ZN(n656) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n824), .B1(n934), .B2(\mem[19][3] ), 
        .ZN(n931) );
  INV_X1 U290 ( .A(n930), .ZN(n655) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n824), .B1(n934), .B2(\mem[19][4] ), 
        .ZN(n930) );
  INV_X1 U292 ( .A(n929), .ZN(n654) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n824), .B1(n934), .B2(\mem[19][5] ), 
        .ZN(n929) );
  INV_X1 U294 ( .A(n928), .ZN(n653) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n824), .B1(n934), .B2(\mem[19][6] ), 
        .ZN(n928) );
  INV_X1 U296 ( .A(n927), .ZN(n652) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n824), .B1(n934), .B2(\mem[19][7] ), 
        .ZN(n927) );
  INV_X1 U298 ( .A(n908), .ZN(n635) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n821), .B1(n907), .B2(\mem[22][0] ), 
        .ZN(n908) );
  INV_X1 U300 ( .A(n906), .ZN(n634) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n821), .B1(n907), .B2(\mem[22][1] ), 
        .ZN(n906) );
  INV_X1 U302 ( .A(n905), .ZN(n633) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n821), .B1(n907), .B2(\mem[22][2] ), 
        .ZN(n905) );
  INV_X1 U304 ( .A(n904), .ZN(n632) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n821), .B1(n907), .B2(\mem[22][3] ), 
        .ZN(n904) );
  INV_X1 U306 ( .A(n903), .ZN(n631) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n821), .B1(n907), .B2(\mem[22][4] ), 
        .ZN(n903) );
  INV_X1 U308 ( .A(n902), .ZN(n630) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n821), .B1(n907), .B2(\mem[22][5] ), 
        .ZN(n902) );
  INV_X1 U310 ( .A(n901), .ZN(n629) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n821), .B1(n907), .B2(\mem[22][6] ), 
        .ZN(n901) );
  INV_X1 U312 ( .A(n900), .ZN(n628) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n821), .B1(n907), .B2(\mem[22][7] ), 
        .ZN(n900) );
  INV_X1 U314 ( .A(n899), .ZN(n627) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n820), .B1(n898), .B2(\mem[23][0] ), 
        .ZN(n899) );
  INV_X1 U316 ( .A(n897), .ZN(n626) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n820), .B1(n898), .B2(\mem[23][1] ), 
        .ZN(n897) );
  INV_X1 U318 ( .A(n896), .ZN(n625) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n820), .B1(n898), .B2(\mem[23][2] ), 
        .ZN(n896) );
  INV_X1 U320 ( .A(n895), .ZN(n624) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n820), .B1(n898), .B2(\mem[23][3] ), 
        .ZN(n895) );
  INV_X1 U322 ( .A(n894), .ZN(n623) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n820), .B1(n898), .B2(\mem[23][4] ), 
        .ZN(n894) );
  INV_X1 U324 ( .A(n893), .ZN(n622) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n820), .B1(n898), .B2(\mem[23][5] ), 
        .ZN(n893) );
  INV_X1 U326 ( .A(n892), .ZN(n621) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n820), .B1(n898), .B2(\mem[23][6] ), 
        .ZN(n892) );
  INV_X1 U328 ( .A(n891), .ZN(n620) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n820), .B1(n898), .B2(\mem[23][7] ), 
        .ZN(n891) );
  INV_X1 U330 ( .A(N12), .ZN(n255) );
  INV_X1 U331 ( .A(N11), .ZN(n254) );
  INV_X1 U332 ( .A(n999), .ZN(n715) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n831), .B1(n998), .B2(\mem[12][0] ), 
        .ZN(n999) );
  INV_X1 U334 ( .A(n997), .ZN(n714) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n831), .B1(n998), .B2(\mem[12][1] ), 
        .ZN(n997) );
  INV_X1 U336 ( .A(n996), .ZN(n713) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n831), .B1(n998), .B2(\mem[12][2] ), 
        .ZN(n996) );
  INV_X1 U338 ( .A(n995), .ZN(n712) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n831), .B1(n998), .B2(\mem[12][3] ), 
        .ZN(n995) );
  INV_X1 U340 ( .A(n994), .ZN(n711) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n831), .B1(n998), .B2(\mem[12][4] ), 
        .ZN(n994) );
  INV_X1 U342 ( .A(n993), .ZN(n710) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n831), .B1(n998), .B2(\mem[12][5] ), 
        .ZN(n993) );
  INV_X1 U344 ( .A(n992), .ZN(n709) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n831), .B1(n998), .B2(\mem[12][6] ), 
        .ZN(n992) );
  INV_X1 U346 ( .A(n991), .ZN(n708) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n831), .B1(n998), .B2(\mem[12][7] ), 
        .ZN(n991) );
  INV_X1 U348 ( .A(n926), .ZN(n651) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n823), .B1(n925), .B2(\mem[20][0] ), 
        .ZN(n926) );
  INV_X1 U350 ( .A(n924), .ZN(n650) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n823), .B1(n925), .B2(\mem[20][1] ), 
        .ZN(n924) );
  INV_X1 U352 ( .A(n923), .ZN(n649) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n823), .B1(n925), .B2(\mem[20][2] ), 
        .ZN(n923) );
  INV_X1 U354 ( .A(n922), .ZN(n648) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n823), .B1(n925), .B2(\mem[20][3] ), 
        .ZN(n922) );
  INV_X1 U356 ( .A(n921), .ZN(n647) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n823), .B1(n925), .B2(\mem[20][4] ), 
        .ZN(n921) );
  INV_X1 U358 ( .A(n920), .ZN(n646) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n823), .B1(n925), .B2(\mem[20][5] ), 
        .ZN(n920) );
  INV_X1 U360 ( .A(n919), .ZN(n645) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n823), .B1(n925), .B2(\mem[20][6] ), 
        .ZN(n919) );
  INV_X1 U362 ( .A(n918), .ZN(n644) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n823), .B1(n925), .B2(\mem[20][7] ), 
        .ZN(n918) );
  INV_X1 U364 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n835), .B1(n1035), .B2(\mem[8][0] ), 
        .ZN(n1036) );
  INV_X1 U366 ( .A(n1034), .ZN(n746) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n835), .B1(n1035), .B2(\mem[8][1] ), 
        .ZN(n1034) );
  INV_X1 U368 ( .A(n1033), .ZN(n745) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n835), .B1(n1035), .B2(\mem[8][2] ), 
        .ZN(n1033) );
  INV_X1 U370 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n835), .B1(n1035), .B2(\mem[8][3] ), 
        .ZN(n1032) );
  INV_X1 U372 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n835), .B1(n1035), .B2(\mem[8][4] ), 
        .ZN(n1031) );
  INV_X1 U374 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n835), .B1(n1035), .B2(\mem[8][5] ), 
        .ZN(n1030) );
  INV_X1 U376 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n835), .B1(n1035), .B2(\mem[8][6] ), 
        .ZN(n1029) );
  INV_X1 U378 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n835), .B1(n1035), .B2(\mem[8][7] ), 
        .ZN(n1028) );
  INV_X1 U380 ( .A(n963), .ZN(n683) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n827), .B1(n962), .B2(\mem[16][0] ), 
        .ZN(n963) );
  INV_X1 U382 ( .A(n961), .ZN(n682) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n827), .B1(n962), .B2(\mem[16][1] ), 
        .ZN(n961) );
  INV_X1 U384 ( .A(n960), .ZN(n681) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n827), .B1(n962), .B2(\mem[16][2] ), 
        .ZN(n960) );
  INV_X1 U386 ( .A(n959), .ZN(n680) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n827), .B1(n962), .B2(\mem[16][3] ), 
        .ZN(n959) );
  INV_X1 U388 ( .A(n958), .ZN(n679) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n827), .B1(n962), .B2(\mem[16][4] ), 
        .ZN(n958) );
  INV_X1 U390 ( .A(n957), .ZN(n678) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n827), .B1(n962), .B2(\mem[16][5] ), 
        .ZN(n957) );
  INV_X1 U392 ( .A(n956), .ZN(n677) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n827), .B1(n962), .B2(\mem[16][6] ), 
        .ZN(n956) );
  INV_X1 U394 ( .A(n955), .ZN(n676) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n827), .B1(n962), .B2(\mem[16][7] ), 
        .ZN(n955) );
  INV_X1 U396 ( .A(n890), .ZN(n619) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n816), .B1(n889), .B2(\mem[24][0] ), 
        .ZN(n890) );
  INV_X1 U398 ( .A(n888), .ZN(n618) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n816), .B1(n889), .B2(\mem[24][1] ), 
        .ZN(n888) );
  INV_X1 U400 ( .A(n887), .ZN(n617) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n816), .B1(n889), .B2(\mem[24][2] ), 
        .ZN(n887) );
  INV_X1 U402 ( .A(n886), .ZN(n616) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n816), .B1(n889), .B2(\mem[24][3] ), 
        .ZN(n886) );
  INV_X1 U404 ( .A(n885), .ZN(n615) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n816), .B1(n889), .B2(\mem[24][4] ), 
        .ZN(n885) );
  INV_X1 U406 ( .A(n884), .ZN(n614) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n816), .B1(n889), .B2(\mem[24][5] ), 
        .ZN(n884) );
  INV_X1 U408 ( .A(n883), .ZN(n613) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n816), .B1(n889), .B2(\mem[24][6] ), 
        .ZN(n883) );
  INV_X1 U410 ( .A(n882), .ZN(n612) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n816), .B1(n889), .B2(\mem[24][7] ), 
        .ZN(n882) );
  INV_X1 U412 ( .A(n881), .ZN(n611) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n815), .B1(n880), .B2(\mem[25][0] ), 
        .ZN(n881) );
  INV_X1 U414 ( .A(n879), .ZN(n610) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n815), .B1(n880), .B2(\mem[25][1] ), 
        .ZN(n879) );
  INV_X1 U416 ( .A(n878), .ZN(n609) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n815), .B1(n880), .B2(\mem[25][2] ), 
        .ZN(n878) );
  INV_X1 U418 ( .A(n877), .ZN(n608) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n815), .B1(n880), .B2(\mem[25][3] ), 
        .ZN(n877) );
  INV_X1 U420 ( .A(n876), .ZN(n607) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n815), .B1(n880), .B2(\mem[25][4] ), 
        .ZN(n876) );
  INV_X1 U422 ( .A(n875), .ZN(n606) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n815), .B1(n880), .B2(\mem[25][5] ), 
        .ZN(n875) );
  INV_X1 U424 ( .A(n874), .ZN(n605) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n815), .B1(n880), .B2(\mem[25][6] ), 
        .ZN(n874) );
  INV_X1 U426 ( .A(n873), .ZN(n604) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n815), .B1(n880), .B2(\mem[25][7] ), 
        .ZN(n873) );
  INV_X1 U428 ( .A(n872), .ZN(n603) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n814), .B1(n871), .B2(\mem[26][0] ), 
        .ZN(n872) );
  INV_X1 U430 ( .A(n870), .ZN(n602) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n814), .B1(n871), .B2(\mem[26][1] ), 
        .ZN(n870) );
  INV_X1 U432 ( .A(n869), .ZN(n601) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n814), .B1(n871), .B2(\mem[26][2] ), 
        .ZN(n869) );
  INV_X1 U434 ( .A(n868), .ZN(n600) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n814), .B1(n871), .B2(\mem[26][3] ), 
        .ZN(n868) );
  INV_X1 U436 ( .A(n867), .ZN(n599) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n814), .B1(n871), .B2(\mem[26][4] ), 
        .ZN(n867) );
  INV_X1 U438 ( .A(n866), .ZN(n598) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n814), .B1(n871), .B2(\mem[26][5] ), 
        .ZN(n866) );
  INV_X1 U440 ( .A(n865), .ZN(n597) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n814), .B1(n871), .B2(\mem[26][6] ), 
        .ZN(n865) );
  INV_X1 U442 ( .A(n864), .ZN(n596) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n814), .B1(n871), .B2(\mem[26][7] ), 
        .ZN(n864) );
  INV_X1 U444 ( .A(n863), .ZN(n595) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n813), .B1(n862), .B2(\mem[27][0] ), 
        .ZN(n863) );
  INV_X1 U446 ( .A(n861), .ZN(n594) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n813), .B1(n862), .B2(\mem[27][1] ), 
        .ZN(n861) );
  INV_X1 U448 ( .A(n860), .ZN(n293) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n813), .B1(n862), .B2(\mem[27][2] ), 
        .ZN(n860) );
  INV_X1 U450 ( .A(n859), .ZN(n292) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n813), .B1(n862), .B2(\mem[27][3] ), 
        .ZN(n859) );
  INV_X1 U452 ( .A(n858), .ZN(n291) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n813), .B1(n862), .B2(\mem[27][4] ), 
        .ZN(n858) );
  INV_X1 U454 ( .A(n857), .ZN(n290) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n813), .B1(n862), .B2(\mem[27][5] ), 
        .ZN(n857) );
  INV_X1 U456 ( .A(n856), .ZN(n289) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n813), .B1(n862), .B2(\mem[27][6] ), 
        .ZN(n856) );
  INV_X1 U458 ( .A(n855), .ZN(n288) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n813), .B1(n862), .B2(\mem[27][7] ), 
        .ZN(n855) );
  INV_X1 U460 ( .A(n854), .ZN(n287) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n812), .B1(n853), .B2(\mem[28][0] ), 
        .ZN(n854) );
  INV_X1 U462 ( .A(n852), .ZN(n286) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n812), .B1(n853), .B2(\mem[28][1] ), 
        .ZN(n852) );
  INV_X1 U464 ( .A(n851), .ZN(n285) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n812), .B1(n853), .B2(\mem[28][2] ), 
        .ZN(n851) );
  INV_X1 U466 ( .A(n850), .ZN(n284) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n812), .B1(n853), .B2(\mem[28][3] ), 
        .ZN(n850) );
  INV_X1 U468 ( .A(n849), .ZN(n283) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n812), .B1(n853), .B2(\mem[28][4] ), 
        .ZN(n849) );
  INV_X1 U470 ( .A(n848), .ZN(n282) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n812), .B1(n853), .B2(\mem[28][5] ), 
        .ZN(n848) );
  INV_X1 U472 ( .A(n847), .ZN(n281) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n812), .B1(n853), .B2(\mem[28][6] ), 
        .ZN(n847) );
  INV_X1 U474 ( .A(n846), .ZN(n280) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n812), .B1(n853), .B2(\mem[28][7] ), 
        .ZN(n846) );
  INV_X1 U476 ( .A(n1145), .ZN(n279) );
  AOI22_X1 U477 ( .A1(n819), .A2(data_in[0]), .B1(n1144), .B2(\mem[29][0] ), 
        .ZN(n1145) );
  INV_X1 U478 ( .A(n1143), .ZN(n278) );
  AOI22_X1 U479 ( .A1(n819), .A2(data_in[1]), .B1(n1144), .B2(\mem[29][1] ), 
        .ZN(n1143) );
  INV_X1 U480 ( .A(n1142), .ZN(n277) );
  AOI22_X1 U481 ( .A1(n819), .A2(data_in[2]), .B1(n1144), .B2(\mem[29][2] ), 
        .ZN(n1142) );
  INV_X1 U482 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U483 ( .A1(n819), .A2(data_in[3]), .B1(n1144), .B2(\mem[29][3] ), 
        .ZN(n1141) );
  INV_X1 U484 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U485 ( .A1(n819), .A2(data_in[4]), .B1(n1144), .B2(\mem[29][4] ), 
        .ZN(n1140) );
  INV_X1 U486 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U487 ( .A1(n819), .A2(data_in[5]), .B1(n1144), .B2(\mem[29][5] ), 
        .ZN(n1139) );
  INV_X1 U488 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U489 ( .A1(n819), .A2(data_in[6]), .B1(n1144), .B2(\mem[29][6] ), 
        .ZN(n1138) );
  INV_X1 U490 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U491 ( .A1(n819), .A2(data_in[7]), .B1(n1144), .B2(\mem[29][7] ), 
        .ZN(n1137) );
  INV_X1 U492 ( .A(n1134), .ZN(n271) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n818), .B1(n1133), .B2(\mem[30][0] ), 
        .ZN(n1134) );
  INV_X1 U494 ( .A(n1132), .ZN(n270) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n818), .B1(n1133), .B2(\mem[30][1] ), 
        .ZN(n1132) );
  INV_X1 U496 ( .A(n1131), .ZN(n269) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n818), .B1(n1133), .B2(\mem[30][2] ), 
        .ZN(n1131) );
  INV_X1 U498 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n818), .B1(n1133), .B2(\mem[30][3] ), 
        .ZN(n1130) );
  INV_X1 U500 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n818), .B1(n1133), .B2(\mem[30][4] ), 
        .ZN(n1129) );
  INV_X1 U502 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n818), .B1(n1133), .B2(\mem[30][5] ), 
        .ZN(n1128) );
  INV_X1 U504 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n818), .B1(n1133), .B2(\mem[30][6] ), 
        .ZN(n1127) );
  INV_X1 U506 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n818), .B1(n1133), .B2(\mem[30][7] ), 
        .ZN(n1126) );
  INV_X1 U508 ( .A(n1124), .ZN(n263) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n817), .B1(n1123), .B2(\mem[31][0] ), 
        .ZN(n1124) );
  INV_X1 U510 ( .A(n1122), .ZN(n262) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n817), .B1(n1123), .B2(\mem[31][1] ), 
        .ZN(n1122) );
  INV_X1 U512 ( .A(n1121), .ZN(n261) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n817), .B1(n1123), .B2(\mem[31][2] ), 
        .ZN(n1121) );
  INV_X1 U514 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n817), .B1(n1123), .B2(\mem[31][3] ), 
        .ZN(n1120) );
  INV_X1 U516 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n817), .B1(n1123), .B2(\mem[31][4] ), 
        .ZN(n1119) );
  INV_X1 U518 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n817), .B1(n1123), .B2(\mem[31][5] ), 
        .ZN(n1118) );
  INV_X1 U520 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n817), .B1(n1123), .B2(\mem[31][6] ), 
        .ZN(n1117) );
  INV_X1 U522 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n817), .B1(n1123), .B2(\mem[31][7] ), 
        .ZN(n1116) );
  INV_X1 U524 ( .A(n1114), .ZN(n811) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n843), .B1(n1113), .B2(\mem[0][0] ), 
        .ZN(n1114) );
  INV_X1 U526 ( .A(n1112), .ZN(n810) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n843), .B1(n1113), .B2(\mem[0][1] ), 
        .ZN(n1112) );
  INV_X1 U528 ( .A(n1111), .ZN(n809) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n843), .B1(n1113), .B2(\mem[0][2] ), 
        .ZN(n1111) );
  INV_X1 U530 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n843), .B1(n1113), .B2(\mem[0][3] ), 
        .ZN(n1110) );
  INV_X1 U532 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n843), .B1(n1113), .B2(\mem[0][4] ), 
        .ZN(n1109) );
  INV_X1 U534 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n843), .B1(n1113), .B2(\mem[0][5] ), 
        .ZN(n1108) );
  INV_X1 U536 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n843), .B1(n1113), .B2(\mem[0][6] ), 
        .ZN(n1107) );
  INV_X1 U538 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n843), .B1(n1113), .B2(\mem[0][7] ), 
        .ZN(n1106) );
  INV_X1 U540 ( .A(n1103), .ZN(n803) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[1][0] ), 
        .ZN(n1103) );
  INV_X1 U542 ( .A(n1101), .ZN(n802) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[1][1] ), 
        .ZN(n1101) );
  INV_X1 U544 ( .A(n1100), .ZN(n801) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[1][2] ), 
        .ZN(n1100) );
  INV_X1 U546 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[1][3] ), 
        .ZN(n1099) );
  INV_X1 U548 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[1][4] ), 
        .ZN(n1098) );
  INV_X1 U550 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[1][5] ), 
        .ZN(n1097) );
  INV_X1 U552 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[1][6] ), 
        .ZN(n1096) );
  INV_X1 U554 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[1][7] ), 
        .ZN(n1095) );
  INV_X1 U556 ( .A(n1093), .ZN(n795) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n841), .B1(n1092), .B2(\mem[2][0] ), 
        .ZN(n1093) );
  INV_X1 U558 ( .A(n1091), .ZN(n794) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n841), .B1(n1092), .B2(\mem[2][1] ), 
        .ZN(n1091) );
  INV_X1 U560 ( .A(n1090), .ZN(n793) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n841), .B1(n1092), .B2(\mem[2][2] ), 
        .ZN(n1090) );
  INV_X1 U562 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n841), .B1(n1092), .B2(\mem[2][3] ), 
        .ZN(n1089) );
  INV_X1 U564 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n841), .B1(n1092), .B2(\mem[2][4] ), 
        .ZN(n1088) );
  INV_X1 U566 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n841), .B1(n1092), .B2(\mem[2][5] ), 
        .ZN(n1087) );
  INV_X1 U568 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n841), .B1(n1092), .B2(\mem[2][6] ), 
        .ZN(n1086) );
  INV_X1 U570 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n841), .B1(n1092), .B2(\mem[2][7] ), 
        .ZN(n1085) );
  INV_X1 U572 ( .A(n1083), .ZN(n787) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n840), .B1(n1082), .B2(\mem[3][0] ), 
        .ZN(n1083) );
  INV_X1 U574 ( .A(n1081), .ZN(n786) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n840), .B1(n1082), .B2(\mem[3][1] ), 
        .ZN(n1081) );
  INV_X1 U576 ( .A(n1080), .ZN(n785) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n840), .B1(n1082), .B2(\mem[3][2] ), 
        .ZN(n1080) );
  INV_X1 U578 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n840), .B1(n1082), .B2(\mem[3][3] ), 
        .ZN(n1079) );
  INV_X1 U580 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n840), .B1(n1082), .B2(\mem[3][4] ), 
        .ZN(n1078) );
  INV_X1 U582 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n840), .B1(n1082), .B2(\mem[3][5] ), 
        .ZN(n1077) );
  INV_X1 U584 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n840), .B1(n1082), .B2(\mem[3][6] ), 
        .ZN(n1076) );
  INV_X1 U586 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n840), .B1(n1082), .B2(\mem[3][7] ), 
        .ZN(n1075) );
  INV_X1 U588 ( .A(n1073), .ZN(n779) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n839), .B1(n1072), .B2(\mem[4][0] ), 
        .ZN(n1073) );
  INV_X1 U590 ( .A(n1071), .ZN(n778) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n839), .B1(n1072), .B2(\mem[4][1] ), 
        .ZN(n1071) );
  INV_X1 U592 ( .A(n1070), .ZN(n777) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n839), .B1(n1072), .B2(\mem[4][2] ), 
        .ZN(n1070) );
  INV_X1 U594 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n839), .B1(n1072), .B2(\mem[4][3] ), 
        .ZN(n1069) );
  INV_X1 U596 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n839), .B1(n1072), .B2(\mem[4][4] ), 
        .ZN(n1068) );
  INV_X1 U598 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n839), .B1(n1072), .B2(\mem[4][5] ), 
        .ZN(n1067) );
  INV_X1 U600 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n839), .B1(n1072), .B2(\mem[4][6] ), 
        .ZN(n1066) );
  INV_X1 U602 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n839), .B1(n1072), .B2(\mem[4][7] ), 
        .ZN(n1065) );
  INV_X1 U604 ( .A(N13), .ZN(n844) );
  INV_X1 U605 ( .A(N14), .ZN(n845) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n251), .Z(n3) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n251), .Z(n4) );
  MUX2_X1 U608 ( .A(n4), .B(n3), .S(n244), .Z(n5) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n251), .Z(n6) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n251), .Z(n7) );
  MUX2_X1 U611 ( .A(n7), .B(n6), .S(n244), .Z(n8) );
  MUX2_X1 U612 ( .A(n8), .B(n5), .S(n243), .Z(n9) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n251), .Z(n10) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n250), .Z(n11) );
  MUX2_X1 U615 ( .A(n11), .B(n10), .S(n244), .Z(n12) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n251), .Z(n13) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n250), .Z(n14) );
  MUX2_X1 U618 ( .A(n14), .B(n13), .S(n244), .Z(n15) );
  MUX2_X1 U619 ( .A(n15), .B(n12), .S(n243), .Z(n16) );
  MUX2_X1 U620 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n247), .Z(n18) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n247), .Z(n19) );
  MUX2_X1 U623 ( .A(n19), .B(n18), .S(N11), .Z(n20) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n247), .Z(n21) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n247), .Z(n22) );
  MUX2_X1 U626 ( .A(n22), .B(n21), .S(N11), .Z(n23) );
  MUX2_X1 U627 ( .A(n23), .B(n20), .S(n243), .Z(n24) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n247), .Z(n25) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n247), .Z(n26) );
  MUX2_X1 U630 ( .A(n26), .B(n25), .S(N11), .Z(n27) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n247), .Z(n28) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n247), .Z(n29) );
  MUX2_X1 U633 ( .A(n29), .B(n28), .S(n246), .Z(n30) );
  MUX2_X1 U634 ( .A(n30), .B(n27), .S(n243), .Z(n31) );
  MUX2_X1 U635 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U636 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n247), .Z(n33) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n247), .Z(n34) );
  MUX2_X1 U639 ( .A(n34), .B(n33), .S(n246), .Z(n35) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n247), .Z(n36) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n247), .Z(n37) );
  MUX2_X1 U642 ( .A(n37), .B(n36), .S(N11), .Z(n38) );
  MUX2_X1 U643 ( .A(n38), .B(n35), .S(n243), .Z(n39) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n248), .Z(n40) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n248), .Z(n41) );
  MUX2_X1 U646 ( .A(n41), .B(n40), .S(N11), .Z(n42) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n248), .Z(n43) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n248), .Z(n44) );
  MUX2_X1 U649 ( .A(n44), .B(n43), .S(n244), .Z(n45) );
  MUX2_X1 U650 ( .A(n45), .B(n42), .S(N12), .Z(n46) );
  MUX2_X1 U651 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n248), .Z(n48) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n248), .Z(n49) );
  MUX2_X1 U654 ( .A(n49), .B(n48), .S(N11), .Z(n50) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n248), .Z(n51) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n248), .Z(n52) );
  MUX2_X1 U657 ( .A(n52), .B(n51), .S(n246), .Z(n53) );
  MUX2_X1 U658 ( .A(n53), .B(n50), .S(N12), .Z(n54) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n248), .Z(n55) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n248), .Z(n56) );
  MUX2_X1 U661 ( .A(n56), .B(n55), .S(N11), .Z(n57) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n248), .Z(n58) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n248), .Z(n59) );
  MUX2_X1 U664 ( .A(n59), .B(n58), .S(n245), .Z(n60) );
  MUX2_X1 U665 ( .A(n60), .B(n57), .S(N12), .Z(n61) );
  MUX2_X1 U666 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U667 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n249), .Z(n63) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n249), .Z(n64) );
  MUX2_X1 U670 ( .A(n64), .B(n63), .S(n245), .Z(n65) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n249), .Z(n66) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n249), .Z(n67) );
  MUX2_X1 U673 ( .A(n67), .B(n66), .S(n246), .Z(n68) );
  MUX2_X1 U674 ( .A(n68), .B(n65), .S(n243), .Z(n69) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n249), .Z(n70) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n249), .Z(n71) );
  MUX2_X1 U677 ( .A(n71), .B(n70), .S(n244), .Z(n72) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n249), .Z(n73) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n249), .Z(n74) );
  MUX2_X1 U680 ( .A(n74), .B(n73), .S(N11), .Z(n75) );
  MUX2_X1 U681 ( .A(n75), .B(n72), .S(n243), .Z(n76) );
  MUX2_X1 U682 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n249), .Z(n78) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n249), .Z(n79) );
  MUX2_X1 U685 ( .A(n79), .B(n78), .S(n245), .Z(n80) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n249), .Z(n81) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n249), .Z(n82) );
  MUX2_X1 U688 ( .A(n82), .B(n81), .S(N11), .Z(n83) );
  MUX2_X1 U689 ( .A(n83), .B(n80), .S(n243), .Z(n84) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n249), .Z(n85) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n250), .Z(n86) );
  MUX2_X1 U692 ( .A(n86), .B(n85), .S(n244), .Z(n87) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n247), .Z(n88) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n250), .Z(n89) );
  MUX2_X1 U695 ( .A(n89), .B(n88), .S(N11), .Z(n90) );
  MUX2_X1 U696 ( .A(n90), .B(n87), .S(n243), .Z(n91) );
  MUX2_X1 U697 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U698 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n248), .Z(n93) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U701 ( .A(n94), .B(n93), .S(n246), .Z(n95) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n249), .Z(n96) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n248), .Z(n97) );
  MUX2_X1 U704 ( .A(n97), .B(n96), .S(n245), .Z(n98) );
  MUX2_X1 U705 ( .A(n98), .B(n95), .S(n243), .Z(n99) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n252), .Z(n100) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n248), .Z(n101) );
  MUX2_X1 U708 ( .A(n101), .B(n100), .S(N11), .Z(n102) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n247), .Z(n103) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n249), .Z(n104) );
  MUX2_X1 U711 ( .A(n104), .B(n103), .S(N11), .Z(n105) );
  MUX2_X1 U712 ( .A(n105), .B(n102), .S(n243), .Z(n106) );
  MUX2_X1 U713 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n251), .Z(n108) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(N10), .Z(n109) );
  MUX2_X1 U716 ( .A(n109), .B(n108), .S(n244), .Z(n110) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(N10), .Z(n111) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n112) );
  MUX2_X1 U719 ( .A(n112), .B(n111), .S(n246), .Z(n113) );
  MUX2_X1 U720 ( .A(n113), .B(n110), .S(n243), .Z(n114) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n252), .Z(n115) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n116) );
  MUX2_X1 U723 ( .A(n116), .B(n115), .S(n244), .Z(n117) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n118) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n119) );
  MUX2_X1 U726 ( .A(n119), .B(n118), .S(n245), .Z(n120) );
  MUX2_X1 U727 ( .A(n120), .B(n117), .S(n243), .Z(n121) );
  MUX2_X1 U728 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U729 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n251), .Z(n123) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(N10), .Z(n124) );
  MUX2_X1 U732 ( .A(n124), .B(n123), .S(n244), .Z(n125) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n251), .Z(n126) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n251), .Z(n127) );
  MUX2_X1 U735 ( .A(n127), .B(n126), .S(n244), .Z(n128) );
  MUX2_X1 U736 ( .A(n128), .B(n125), .S(n243), .Z(n129) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n250), .Z(n130) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n250), .Z(n131) );
  MUX2_X1 U739 ( .A(n131), .B(n130), .S(n244), .Z(n132) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n250), .Z(n133) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n250), .Z(n134) );
  MUX2_X1 U742 ( .A(n134), .B(n133), .S(N11), .Z(n135) );
  MUX2_X1 U743 ( .A(n135), .B(n132), .S(n243), .Z(n136) );
  MUX2_X1 U744 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n250), .Z(n138) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n250), .Z(n139) );
  MUX2_X1 U747 ( .A(n139), .B(n138), .S(n244), .Z(n140) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n250), .Z(n141) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n250), .Z(n142) );
  MUX2_X1 U750 ( .A(n142), .B(n141), .S(n245), .Z(n143) );
  MUX2_X1 U751 ( .A(n143), .B(n140), .S(n243), .Z(n144) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n250), .Z(n145) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n250), .Z(n146) );
  MUX2_X1 U754 ( .A(n146), .B(n145), .S(n244), .Z(n147) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n250), .Z(n148) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n250), .Z(n149) );
  MUX2_X1 U757 ( .A(n149), .B(n148), .S(n244), .Z(n150) );
  MUX2_X1 U758 ( .A(n150), .B(n147), .S(n243), .Z(n151) );
  MUX2_X1 U759 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U760 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n251), .Z(n153) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n251), .Z(n154) );
  MUX2_X1 U763 ( .A(n154), .B(n153), .S(n245), .Z(n155) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n251), .Z(n156) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n251), .Z(n157) );
  MUX2_X1 U766 ( .A(n157), .B(n156), .S(n245), .Z(n158) );
  MUX2_X1 U767 ( .A(n158), .B(n155), .S(n243), .Z(n159) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n251), .Z(n160) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n251), .Z(n161) );
  MUX2_X1 U770 ( .A(n161), .B(n160), .S(n245), .Z(n162) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n251), .Z(n163) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n251), .Z(n164) );
  MUX2_X1 U773 ( .A(n164), .B(n163), .S(n245), .Z(n165) );
  MUX2_X1 U774 ( .A(n165), .B(n162), .S(n243), .Z(n166) );
  MUX2_X1 U775 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n251), .Z(n168) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n251), .Z(n169) );
  MUX2_X1 U778 ( .A(n169), .B(n168), .S(n245), .Z(n170) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n251), .Z(n171) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n251), .Z(n172) );
  MUX2_X1 U781 ( .A(n172), .B(n171), .S(n245), .Z(n173) );
  MUX2_X1 U782 ( .A(n173), .B(n170), .S(n243), .Z(n174) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n251), .Z(n175) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n247), .Z(n176) );
  MUX2_X1 U785 ( .A(n176), .B(n175), .S(n245), .Z(n177) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n249), .Z(n178) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n247), .Z(n179) );
  MUX2_X1 U788 ( .A(n179), .B(n178), .S(n245), .Z(n180) );
  MUX2_X1 U789 ( .A(n180), .B(n177), .S(n243), .Z(n181) );
  MUX2_X1 U790 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U791 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n248), .Z(n183) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n252), .Z(n184) );
  MUX2_X1 U794 ( .A(n184), .B(n183), .S(n245), .Z(n185) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n252), .Z(n186) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n252), .Z(n187) );
  MUX2_X1 U797 ( .A(n187), .B(n186), .S(n245), .Z(n188) );
  MUX2_X1 U798 ( .A(n188), .B(n185), .S(n243), .Z(n189) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n252), .Z(n190) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n248), .Z(n191) );
  MUX2_X1 U801 ( .A(n191), .B(n190), .S(n245), .Z(n192) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n252), .Z(n193) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n252), .Z(n194) );
  MUX2_X1 U804 ( .A(n194), .B(n193), .S(n245), .Z(n195) );
  MUX2_X1 U805 ( .A(n195), .B(n192), .S(N12), .Z(n196) );
  MUX2_X1 U806 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n252), .Z(n198) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n252), .Z(n199) );
  MUX2_X1 U809 ( .A(n199), .B(n198), .S(n246), .Z(n200) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n252), .Z(n201) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n247), .Z(n202) );
  MUX2_X1 U812 ( .A(n202), .B(n201), .S(n246), .Z(n203) );
  MUX2_X1 U813 ( .A(n203), .B(n200), .S(N12), .Z(n204) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n252), .Z(n205) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n252), .Z(n206) );
  MUX2_X1 U816 ( .A(n206), .B(n205), .S(n246), .Z(n207) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n252), .Z(n208) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n249), .Z(n209) );
  MUX2_X1 U819 ( .A(n209), .B(n208), .S(n246), .Z(n210) );
  MUX2_X1 U820 ( .A(n210), .B(n207), .S(N12), .Z(n211) );
  MUX2_X1 U821 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U822 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n250), .Z(n213) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n252), .Z(n214) );
  MUX2_X1 U825 ( .A(n214), .B(n213), .S(n246), .Z(n215) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n252), .Z(n216) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n252), .Z(n217) );
  MUX2_X1 U828 ( .A(n217), .B(n216), .S(n246), .Z(n218) );
  MUX2_X1 U829 ( .A(n218), .B(n215), .S(n243), .Z(n219) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n252), .Z(n220) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(N10), .Z(n221) );
  MUX2_X1 U832 ( .A(n221), .B(n220), .S(n246), .Z(n222) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(N10), .Z(n223) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n252), .Z(n224) );
  MUX2_X1 U835 ( .A(n224), .B(n223), .S(n246), .Z(n225) );
  MUX2_X1 U836 ( .A(n225), .B(n222), .S(N12), .Z(n226) );
  MUX2_X1 U837 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n252), .Z(n228) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n229) );
  MUX2_X1 U840 ( .A(n229), .B(n228), .S(n246), .Z(n230) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(N10), .Z(n231) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n232) );
  MUX2_X1 U843 ( .A(n232), .B(n231), .S(n246), .Z(n233) );
  MUX2_X1 U844 ( .A(n233), .B(n230), .S(N12), .Z(n234) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n235) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n247), .Z(n236) );
  MUX2_X1 U847 ( .A(n236), .B(n235), .S(n246), .Z(n237) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n238) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n248), .Z(n239) );
  MUX2_X1 U850 ( .A(n239), .B(n238), .S(n246), .Z(n240) );
  MUX2_X1 U851 ( .A(n240), .B(n237), .S(N12), .Z(n241) );
  MUX2_X1 U852 ( .A(n241), .B(n234), .S(N13), .Z(n242) );
  MUX2_X1 U853 ( .A(n242), .B(n227), .S(N14), .Z(N15) );
  CLKBUF_X1 U854 ( .A(N11), .Z(n244) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_24 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  BUF_X1 U3 ( .A(n250), .Z(n248) );
  BUF_X1 U4 ( .A(N10), .Z(n249) );
  BUF_X1 U5 ( .A(n250), .Z(n246) );
  BUF_X1 U6 ( .A(n250), .Z(n245) );
  BUF_X1 U7 ( .A(n250), .Z(n247) );
  BUF_X1 U8 ( .A(N10), .Z(n250) );
  INV_X1 U9 ( .A(n1111), .ZN(n841) );
  INV_X1 U10 ( .A(n1100), .ZN(n840) );
  INV_X1 U11 ( .A(n1090), .ZN(n839) );
  INV_X1 U12 ( .A(n1080), .ZN(n838) );
  INV_X1 U13 ( .A(n1070), .ZN(n837) );
  INV_X1 U14 ( .A(n1060), .ZN(n836) );
  INV_X1 U15 ( .A(n1051), .ZN(n835) );
  INV_X1 U16 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U19 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U20 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U21 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U22 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U23 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U24 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U26 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U27 ( .A(n1131), .ZN(n816) );
  INV_X1 U28 ( .A(n1121), .ZN(n815) );
  INV_X1 U29 ( .A(n887), .ZN(n814) );
  INV_X1 U30 ( .A(n878), .ZN(n813) );
  INV_X1 U31 ( .A(n869), .ZN(n812) );
  INV_X1 U32 ( .A(n860), .ZN(n811) );
  INV_X1 U33 ( .A(n851), .ZN(n810) );
  INV_X1 U34 ( .A(n987), .ZN(n828) );
  INV_X1 U35 ( .A(n978), .ZN(n827) );
  INV_X1 U36 ( .A(n969), .ZN(n826) );
  INV_X1 U37 ( .A(n914), .ZN(n820) );
  INV_X1 U38 ( .A(n905), .ZN(n819) );
  INV_X1 U39 ( .A(n896), .ZN(n818) );
  INV_X1 U40 ( .A(n1033), .ZN(n833) );
  INV_X1 U41 ( .A(n1023), .ZN(n832) );
  INV_X1 U42 ( .A(n1014), .ZN(n831) );
  INV_X1 U43 ( .A(n1005), .ZN(n830) );
  INV_X1 U44 ( .A(n996), .ZN(n829) );
  INV_X1 U45 ( .A(n960), .ZN(n825) );
  INV_X1 U46 ( .A(n950), .ZN(n824) );
  INV_X1 U47 ( .A(n941), .ZN(n823) );
  INV_X1 U48 ( .A(n932), .ZN(n822) );
  INV_X1 U49 ( .A(n923), .ZN(n821) );
  INV_X1 U50 ( .A(n1142), .ZN(n817) );
  BUF_X1 U51 ( .A(N11), .Z(n242) );
  BUF_X1 U52 ( .A(N11), .Z(n243) );
  BUF_X1 U53 ( .A(N11), .Z(n244) );
  INV_X1 U54 ( .A(N10), .ZN(n251) );
  BUF_X1 U55 ( .A(N12), .Z(n241) );
  NOR3_X1 U56 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U57 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U58 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U60 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U62 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U63 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U64 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U65 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U67 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U69 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U70 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U71 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U72 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U73 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U74 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U75 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U76 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U77 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U79 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U81 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U82 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U83 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U84 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U85 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U86 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U88 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U89 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U90 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U92 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U94 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U95 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U96 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U97 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U98 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U99 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U100 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U101 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U102 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U103 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U104 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U105 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U106 ( .A(n912), .ZN(n639) );
  AOI22_X1 U107 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U108 ( .A(n911), .ZN(n638) );
  AOI22_X1 U109 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U110 ( .A(n910), .ZN(n637) );
  AOI22_X1 U111 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U112 ( .A(n909), .ZN(n636) );
  AOI22_X1 U113 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U114 ( .A(n908), .ZN(n635) );
  AOI22_X1 U115 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U116 ( .A(n907), .ZN(n634) );
  AOI22_X1 U117 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U118 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U119 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U120 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U121 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U122 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U123 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U124 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U125 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U126 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U127 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U128 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U129 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U130 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U131 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U132 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U133 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U134 ( .A(n988), .ZN(n705) );
  AOI22_X1 U135 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U136 ( .A(n986), .ZN(n704) );
  AOI22_X1 U137 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U138 ( .A(n985), .ZN(n703) );
  AOI22_X1 U139 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U140 ( .A(n984), .ZN(n702) );
  AOI22_X1 U141 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U142 ( .A(n983), .ZN(n701) );
  AOI22_X1 U143 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U144 ( .A(n982), .ZN(n700) );
  AOI22_X1 U145 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U146 ( .A(n981), .ZN(n699) );
  AOI22_X1 U147 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U148 ( .A(n980), .ZN(n698) );
  AOI22_X1 U149 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U150 ( .A(n926), .ZN(n651) );
  AOI22_X1 U151 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U152 ( .A(n925), .ZN(n650) );
  AOI22_X1 U153 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U154 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U155 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U156 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U157 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U158 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U159 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U160 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U161 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U162 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U163 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U164 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U165 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U166 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U167 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U168 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U169 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U170 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U171 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U172 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U173 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U174 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U175 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U176 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U177 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U178 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U179 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U180 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U181 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U182 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U183 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U184 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U185 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U186 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U187 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U188 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U189 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U190 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U191 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U192 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U193 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U194 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U195 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U196 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U197 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U198 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U199 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U200 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U201 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U202 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U203 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U204 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U205 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U206 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U207 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U208 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U209 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U210 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U211 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U212 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U213 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U214 ( .A(n999), .ZN(n715) );
  AOI22_X1 U215 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U216 ( .A(n998), .ZN(n714) );
  AOI22_X1 U217 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U218 ( .A(n951), .ZN(n673) );
  AOI22_X1 U219 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U220 ( .A(n949), .ZN(n672) );
  AOI22_X1 U221 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U222 ( .A(n948), .ZN(n671) );
  AOI22_X1 U223 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U224 ( .A(n947), .ZN(n670) );
  AOI22_X1 U225 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U226 ( .A(n946), .ZN(n669) );
  AOI22_X1 U227 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U228 ( .A(n945), .ZN(n668) );
  AOI22_X1 U229 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U230 ( .A(n944), .ZN(n667) );
  AOI22_X1 U231 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U232 ( .A(n943), .ZN(n666) );
  AOI22_X1 U233 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U234 ( .A(n915), .ZN(n641) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U236 ( .A(n913), .ZN(n640) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U238 ( .A(n979), .ZN(n697) );
  AOI22_X1 U239 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U240 ( .A(n977), .ZN(n696) );
  AOI22_X1 U241 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U242 ( .A(n976), .ZN(n695) );
  AOI22_X1 U243 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U244 ( .A(n975), .ZN(n694) );
  AOI22_X1 U245 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U246 ( .A(n974), .ZN(n693) );
  AOI22_X1 U247 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U248 ( .A(n973), .ZN(n692) );
  AOI22_X1 U249 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U250 ( .A(n972), .ZN(n691) );
  AOI22_X1 U251 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U252 ( .A(n971), .ZN(n690) );
  AOI22_X1 U253 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U254 ( .A(n970), .ZN(n689) );
  AOI22_X1 U255 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U256 ( .A(n968), .ZN(n688) );
  AOI22_X1 U257 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U258 ( .A(n967), .ZN(n687) );
  AOI22_X1 U259 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U260 ( .A(n966), .ZN(n686) );
  AOI22_X1 U261 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U262 ( .A(n965), .ZN(n685) );
  AOI22_X1 U263 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U264 ( .A(n964), .ZN(n684) );
  AOI22_X1 U265 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U266 ( .A(n963), .ZN(n683) );
  AOI22_X1 U267 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U268 ( .A(n962), .ZN(n682) );
  AOI22_X1 U269 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U270 ( .A(n942), .ZN(n665) );
  AOI22_X1 U271 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U272 ( .A(n940), .ZN(n664) );
  AOI22_X1 U273 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U274 ( .A(n939), .ZN(n663) );
  AOI22_X1 U275 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U276 ( .A(n938), .ZN(n662) );
  AOI22_X1 U277 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U278 ( .A(n937), .ZN(n661) );
  AOI22_X1 U279 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U280 ( .A(n936), .ZN(n660) );
  AOI22_X1 U281 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U282 ( .A(n935), .ZN(n659) );
  AOI22_X1 U283 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U284 ( .A(n934), .ZN(n658) );
  AOI22_X1 U285 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U286 ( .A(n933), .ZN(n657) );
  AOI22_X1 U287 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U288 ( .A(n931), .ZN(n656) );
  AOI22_X1 U289 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U290 ( .A(n930), .ZN(n655) );
  AOI22_X1 U291 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U292 ( .A(n929), .ZN(n654) );
  AOI22_X1 U293 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U294 ( .A(n928), .ZN(n653) );
  AOI22_X1 U295 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U296 ( .A(n927), .ZN(n652) );
  AOI22_X1 U297 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U298 ( .A(n906), .ZN(n633) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U300 ( .A(n904), .ZN(n632) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U302 ( .A(n903), .ZN(n631) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U304 ( .A(n902), .ZN(n630) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U306 ( .A(n901), .ZN(n629) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U308 ( .A(n900), .ZN(n628) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U310 ( .A(n899), .ZN(n627) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U312 ( .A(n898), .ZN(n626) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U314 ( .A(n897), .ZN(n625) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U316 ( .A(n895), .ZN(n624) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U318 ( .A(n894), .ZN(n623) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U320 ( .A(n893), .ZN(n622) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U322 ( .A(n892), .ZN(n621) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U324 ( .A(n891), .ZN(n620) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U326 ( .A(n890), .ZN(n619) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U328 ( .A(n889), .ZN(n618) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U330 ( .A(N12), .ZN(n253) );
  INV_X1 U331 ( .A(N11), .ZN(n252) );
  INV_X1 U332 ( .A(n997), .ZN(n713) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U334 ( .A(n995), .ZN(n712) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U336 ( .A(n994), .ZN(n711) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U338 ( .A(n993), .ZN(n710) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U340 ( .A(n992), .ZN(n709) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U342 ( .A(n991), .ZN(n708) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U344 ( .A(n990), .ZN(n707) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U346 ( .A(n989), .ZN(n706) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U348 ( .A(n924), .ZN(n649) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U350 ( .A(n922), .ZN(n648) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U352 ( .A(n921), .ZN(n647) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U354 ( .A(n920), .ZN(n646) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U356 ( .A(n919), .ZN(n645) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U358 ( .A(n918), .ZN(n644) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U360 ( .A(n917), .ZN(n643) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U362 ( .A(n916), .ZN(n642) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U364 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U366 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U368 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U370 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U372 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U374 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U376 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U378 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U380 ( .A(n961), .ZN(n681) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U382 ( .A(n959), .ZN(n680) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U384 ( .A(n958), .ZN(n679) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U386 ( .A(n957), .ZN(n678) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U388 ( .A(n956), .ZN(n677) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U390 ( .A(n955), .ZN(n676) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U392 ( .A(n954), .ZN(n675) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U394 ( .A(n953), .ZN(n674) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U396 ( .A(n888), .ZN(n617) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U398 ( .A(n886), .ZN(n616) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U400 ( .A(n885), .ZN(n615) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U402 ( .A(n884), .ZN(n614) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U404 ( .A(n883), .ZN(n613) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U406 ( .A(n882), .ZN(n612) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U408 ( .A(n881), .ZN(n611) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U410 ( .A(n880), .ZN(n610) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U412 ( .A(n879), .ZN(n609) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U414 ( .A(n877), .ZN(n608) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U416 ( .A(n876), .ZN(n607) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U418 ( .A(n875), .ZN(n606) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U420 ( .A(n874), .ZN(n605) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U422 ( .A(n873), .ZN(n604) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U424 ( .A(n872), .ZN(n603) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U426 ( .A(n871), .ZN(n602) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U428 ( .A(n870), .ZN(n601) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U430 ( .A(n868), .ZN(n600) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U432 ( .A(n867), .ZN(n599) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U434 ( .A(n866), .ZN(n598) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U436 ( .A(n865), .ZN(n597) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U438 ( .A(n864), .ZN(n596) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U440 ( .A(n863), .ZN(n595) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U442 ( .A(n862), .ZN(n594) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U444 ( .A(n861), .ZN(n293) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U446 ( .A(n859), .ZN(n292) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U448 ( .A(n858), .ZN(n291) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U450 ( .A(n857), .ZN(n290) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U452 ( .A(n856), .ZN(n289) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U454 ( .A(n855), .ZN(n288) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U456 ( .A(n854), .ZN(n287) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U458 ( .A(n853), .ZN(n286) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U460 ( .A(n852), .ZN(n285) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U462 ( .A(n850), .ZN(n284) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U464 ( .A(n849), .ZN(n283) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U466 ( .A(n848), .ZN(n282) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U468 ( .A(n847), .ZN(n281) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U470 ( .A(n846), .ZN(n280) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U472 ( .A(n845), .ZN(n279) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U474 ( .A(n844), .ZN(n278) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U476 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U477 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U478 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U479 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U480 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U481 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U482 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U483 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U484 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U485 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U486 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U487 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U488 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U489 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U490 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U491 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U492 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U494 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U496 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U498 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U500 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U502 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U504 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U506 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U508 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U510 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U512 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U514 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U516 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U518 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U520 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U522 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U524 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U526 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U528 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U530 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U532 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U534 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U536 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U538 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U540 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U542 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U544 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U546 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U548 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U550 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U552 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U554 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U556 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U558 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U560 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U562 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U564 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U566 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U568 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U570 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U572 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U574 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U576 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U578 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U580 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U582 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U584 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U586 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U588 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U590 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U592 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U594 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U596 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U598 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U600 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U602 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U604 ( .A(N13), .ZN(n842) );
  INV_X1 U605 ( .A(N14), .ZN(n843) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n249), .Z(n1) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n249), .Z(n2) );
  MUX2_X1 U608 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n249), .Z(n4) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n248), .Z(n5) );
  MUX2_X1 U611 ( .A(n5), .B(n4), .S(n243), .Z(n6) );
  MUX2_X1 U612 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n249), .Z(n8) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n248), .Z(n9) );
  MUX2_X1 U615 ( .A(n9), .B(n8), .S(n243), .Z(n10) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n249), .Z(n11) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n248), .Z(n12) );
  MUX2_X1 U618 ( .A(n12), .B(n11), .S(n244), .Z(n13) );
  MUX2_X1 U619 ( .A(n13), .B(n10), .S(N12), .Z(n14) );
  MUX2_X1 U620 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n245), .Z(n16) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n245), .Z(n17) );
  MUX2_X1 U623 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n245), .Z(n20) );
  MUX2_X1 U626 ( .A(n20), .B(n19), .S(N11), .Z(n21) );
  MUX2_X1 U627 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n245), .Z(n23) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n245), .Z(n24) );
  MUX2_X1 U630 ( .A(n24), .B(n23), .S(N11), .Z(n25) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n245), .Z(n26) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n245), .Z(n27) );
  MUX2_X1 U633 ( .A(n27), .B(n26), .S(N11), .Z(n28) );
  MUX2_X1 U634 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U635 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U636 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n245), .Z(n31) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n245), .Z(n32) );
  MUX2_X1 U639 ( .A(n32), .B(n31), .S(n242), .Z(n33) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U642 ( .A(n35), .B(n34), .S(N11), .Z(n36) );
  MUX2_X1 U643 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n246), .Z(n38) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n246), .Z(n39) );
  MUX2_X1 U646 ( .A(n39), .B(n38), .S(n244), .Z(n40) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n246), .Z(n41) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n246), .Z(n42) );
  MUX2_X1 U649 ( .A(n42), .B(n41), .S(n242), .Z(n43) );
  MUX2_X1 U650 ( .A(n43), .B(n40), .S(n241), .Z(n44) );
  MUX2_X1 U651 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n246), .Z(n46) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n246), .Z(n47) );
  MUX2_X1 U654 ( .A(n47), .B(n46), .S(n243), .Z(n48) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n246), .Z(n49) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n246), .Z(n50) );
  MUX2_X1 U657 ( .A(n50), .B(n49), .S(n244), .Z(n51) );
  MUX2_X1 U658 ( .A(n51), .B(n48), .S(n241), .Z(n52) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n246), .Z(n53) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n246), .Z(n54) );
  MUX2_X1 U661 ( .A(n54), .B(n53), .S(n243), .Z(n55) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n246), .Z(n56) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n246), .Z(n57) );
  MUX2_X1 U664 ( .A(n57), .B(n56), .S(N11), .Z(n58) );
  MUX2_X1 U665 ( .A(n58), .B(n55), .S(n241), .Z(n59) );
  MUX2_X1 U666 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U667 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n247), .Z(n61) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n247), .Z(n62) );
  MUX2_X1 U670 ( .A(n62), .B(n61), .S(N11), .Z(n63) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n247), .Z(n64) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n247), .Z(n65) );
  MUX2_X1 U673 ( .A(n65), .B(n64), .S(n244), .Z(n66) );
  MUX2_X1 U674 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n247), .Z(n68) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n247), .Z(n69) );
  MUX2_X1 U677 ( .A(n69), .B(n68), .S(N11), .Z(n70) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n247), .Z(n71) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n247), .Z(n72) );
  MUX2_X1 U680 ( .A(n72), .B(n71), .S(n244), .Z(n73) );
  MUX2_X1 U681 ( .A(n73), .B(n70), .S(n241), .Z(n74) );
  MUX2_X1 U682 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n247), .Z(n76) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n247), .Z(n77) );
  MUX2_X1 U685 ( .A(n77), .B(n76), .S(N11), .Z(n78) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n247), .Z(n79) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n247), .Z(n80) );
  MUX2_X1 U688 ( .A(n80), .B(n79), .S(n243), .Z(n81) );
  MUX2_X1 U689 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n246), .Z(n83) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n247), .Z(n84) );
  MUX2_X1 U692 ( .A(n84), .B(n83), .S(n242), .Z(n85) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n246), .Z(n86) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n246), .Z(n87) );
  MUX2_X1 U695 ( .A(n87), .B(n86), .S(n242), .Z(n88) );
  MUX2_X1 U696 ( .A(n88), .B(n85), .S(n241), .Z(n89) );
  MUX2_X1 U697 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U698 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n247), .Z(n91) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n92) );
  MUX2_X1 U701 ( .A(n92), .B(n91), .S(N11), .Z(n93) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n247), .Z(n95) );
  MUX2_X1 U704 ( .A(n95), .B(n94), .S(n242), .Z(n96) );
  MUX2_X1 U705 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n98) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n248), .Z(n99) );
  MUX2_X1 U708 ( .A(n99), .B(n98), .S(N11), .Z(n100) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n245), .Z(n101) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n248), .Z(n102) );
  MUX2_X1 U711 ( .A(n102), .B(n101), .S(N11), .Z(n103) );
  MUX2_X1 U712 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U713 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n249), .Z(n106) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n250), .Z(n107) );
  MUX2_X1 U716 ( .A(n107), .B(n106), .S(n242), .Z(n108) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n249), .Z(n109) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n110) );
  MUX2_X1 U719 ( .A(n110), .B(n109), .S(n242), .Z(n111) );
  MUX2_X1 U720 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n250), .Z(n113) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n114) );
  MUX2_X1 U723 ( .A(n114), .B(n113), .S(n242), .Z(n115) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n116) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n117) );
  MUX2_X1 U726 ( .A(n117), .B(n116), .S(n242), .Z(n118) );
  MUX2_X1 U727 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U728 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U729 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n249), .Z(n121) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(N10), .Z(n122) );
  MUX2_X1 U732 ( .A(n122), .B(n121), .S(n242), .Z(n123) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n249), .Z(n124) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n125) );
  MUX2_X1 U735 ( .A(n125), .B(n124), .S(n242), .Z(n126) );
  MUX2_X1 U736 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n248), .Z(n128) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n248), .Z(n129) );
  MUX2_X1 U739 ( .A(n129), .B(n128), .S(n242), .Z(n130) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n248), .Z(n131) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n248), .Z(n132) );
  MUX2_X1 U742 ( .A(n132), .B(n131), .S(n242), .Z(n133) );
  MUX2_X1 U743 ( .A(n133), .B(n130), .S(n241), .Z(n134) );
  MUX2_X1 U744 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n248), .Z(n136) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n248), .Z(n137) );
  MUX2_X1 U747 ( .A(n137), .B(n136), .S(n242), .Z(n138) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n248), .Z(n139) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n248), .Z(n140) );
  MUX2_X1 U750 ( .A(n140), .B(n139), .S(n242), .Z(n141) );
  MUX2_X1 U751 ( .A(n141), .B(n138), .S(n241), .Z(n142) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n248), .Z(n143) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n248), .Z(n144) );
  MUX2_X1 U754 ( .A(n144), .B(n143), .S(n242), .Z(n145) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n248), .Z(n146) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n248), .Z(n147) );
  MUX2_X1 U757 ( .A(n147), .B(n146), .S(n242), .Z(n148) );
  MUX2_X1 U758 ( .A(n148), .B(n145), .S(n241), .Z(n149) );
  MUX2_X1 U759 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U760 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n249), .Z(n151) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n249), .Z(n152) );
  MUX2_X1 U763 ( .A(n152), .B(n151), .S(n243), .Z(n153) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n249), .Z(n154) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n249), .Z(n155) );
  MUX2_X1 U766 ( .A(n155), .B(n154), .S(n243), .Z(n156) );
  MUX2_X1 U767 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n249), .Z(n158) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n249), .Z(n159) );
  MUX2_X1 U770 ( .A(n159), .B(n158), .S(n243), .Z(n160) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n249), .Z(n161) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n249), .Z(n162) );
  MUX2_X1 U773 ( .A(n162), .B(n161), .S(n243), .Z(n163) );
  MUX2_X1 U774 ( .A(n163), .B(n160), .S(N12), .Z(n164) );
  MUX2_X1 U775 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n249), .Z(n166) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n249), .Z(n167) );
  MUX2_X1 U778 ( .A(n167), .B(n166), .S(n243), .Z(n168) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n249), .Z(n169) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n249), .Z(n170) );
  MUX2_X1 U781 ( .A(n170), .B(n169), .S(n243), .Z(n171) );
  MUX2_X1 U782 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n250), .Z(n173) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n245), .Z(n174) );
  MUX2_X1 U785 ( .A(n174), .B(n173), .S(n243), .Z(n175) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n247), .Z(n176) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n250), .Z(n177) );
  MUX2_X1 U788 ( .A(n177), .B(n176), .S(n243), .Z(n178) );
  MUX2_X1 U789 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U790 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U791 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n246), .Z(n181) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n245), .Z(n182) );
  MUX2_X1 U794 ( .A(n182), .B(n181), .S(n243), .Z(n183) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n250), .Z(n184) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n250), .Z(n185) );
  MUX2_X1 U797 ( .A(n185), .B(n184), .S(n243), .Z(n186) );
  MUX2_X1 U798 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n246), .Z(n188) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n250), .Z(n189) );
  MUX2_X1 U801 ( .A(n189), .B(n188), .S(n243), .Z(n190) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n250), .Z(n191) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n250), .Z(n192) );
  MUX2_X1 U804 ( .A(n192), .B(n191), .S(n243), .Z(n193) );
  MUX2_X1 U805 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U806 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n249), .Z(n196) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(N10), .Z(n197) );
  MUX2_X1 U809 ( .A(n197), .B(n196), .S(n244), .Z(n198) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n249), .Z(n199) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n250), .Z(n200) );
  MUX2_X1 U812 ( .A(n200), .B(n199), .S(n244), .Z(n201) );
  MUX2_X1 U813 ( .A(n201), .B(n198), .S(N12), .Z(n202) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n203) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n250), .Z(n204) );
  MUX2_X1 U816 ( .A(n204), .B(n203), .S(n244), .Z(n205) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n250), .Z(n206) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n250), .Z(n207) );
  MUX2_X1 U819 ( .A(n207), .B(n206), .S(n244), .Z(n208) );
  MUX2_X1 U820 ( .A(n208), .B(n205), .S(N12), .Z(n209) );
  MUX2_X1 U821 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U822 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n245), .Z(n211) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n247), .Z(n212) );
  MUX2_X1 U825 ( .A(n212), .B(n211), .S(n244), .Z(n213) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n248), .Z(n214) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(N10), .Z(n215) );
  MUX2_X1 U828 ( .A(n215), .B(n214), .S(n244), .Z(n216) );
  MUX2_X1 U829 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n247), .Z(n218) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n250), .Z(n219) );
  MUX2_X1 U832 ( .A(n219), .B(n218), .S(n244), .Z(n220) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n246), .Z(n221) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n222) );
  MUX2_X1 U835 ( .A(n222), .B(n221), .S(n244), .Z(n223) );
  MUX2_X1 U836 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U837 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n250), .Z(n226) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n245), .Z(n227) );
  MUX2_X1 U840 ( .A(n227), .B(n226), .S(n244), .Z(n228) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n250), .Z(n229) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n230) );
  MUX2_X1 U843 ( .A(n230), .B(n229), .S(n244), .Z(n231) );
  MUX2_X1 U844 ( .A(n231), .B(n228), .S(N12), .Z(n232) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n250), .Z(n233) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n234) );
  MUX2_X1 U847 ( .A(n234), .B(n233), .S(n244), .Z(n235) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n236) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n237) );
  MUX2_X1 U850 ( .A(n237), .B(n236), .S(n244), .Z(n238) );
  MUX2_X1 U851 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U852 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U853 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_23 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  BUF_X1 U3 ( .A(n250), .Z(n248) );
  BUF_X1 U4 ( .A(N10), .Z(n249) );
  BUF_X1 U5 ( .A(n250), .Z(n246) );
  BUF_X1 U6 ( .A(n250), .Z(n245) );
  BUF_X1 U7 ( .A(n250), .Z(n247) );
  BUF_X1 U8 ( .A(N10), .Z(n250) );
  INV_X1 U9 ( .A(n1111), .ZN(n841) );
  INV_X1 U10 ( .A(n1100), .ZN(n840) );
  INV_X1 U11 ( .A(n1090), .ZN(n839) );
  INV_X1 U12 ( .A(n1080), .ZN(n838) );
  INV_X1 U13 ( .A(n1070), .ZN(n837) );
  INV_X1 U14 ( .A(n1060), .ZN(n836) );
  INV_X1 U15 ( .A(n1051), .ZN(n835) );
  INV_X1 U16 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U19 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U20 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U21 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U22 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U23 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U24 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U26 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U27 ( .A(n1131), .ZN(n816) );
  INV_X1 U28 ( .A(n1121), .ZN(n815) );
  INV_X1 U29 ( .A(n887), .ZN(n814) );
  INV_X1 U30 ( .A(n878), .ZN(n813) );
  INV_X1 U31 ( .A(n869), .ZN(n812) );
  INV_X1 U32 ( .A(n860), .ZN(n811) );
  INV_X1 U33 ( .A(n851), .ZN(n810) );
  INV_X1 U34 ( .A(n987), .ZN(n828) );
  INV_X1 U35 ( .A(n978), .ZN(n827) );
  INV_X1 U36 ( .A(n969), .ZN(n826) );
  INV_X1 U37 ( .A(n914), .ZN(n820) );
  INV_X1 U38 ( .A(n905), .ZN(n819) );
  INV_X1 U39 ( .A(n896), .ZN(n818) );
  INV_X1 U40 ( .A(n1033), .ZN(n833) );
  INV_X1 U41 ( .A(n1023), .ZN(n832) );
  INV_X1 U42 ( .A(n1014), .ZN(n831) );
  INV_X1 U43 ( .A(n1005), .ZN(n830) );
  INV_X1 U44 ( .A(n996), .ZN(n829) );
  INV_X1 U45 ( .A(n960), .ZN(n825) );
  INV_X1 U46 ( .A(n950), .ZN(n824) );
  INV_X1 U47 ( .A(n941), .ZN(n823) );
  INV_X1 U48 ( .A(n932), .ZN(n822) );
  INV_X1 U49 ( .A(n923), .ZN(n821) );
  INV_X1 U50 ( .A(n1142), .ZN(n817) );
  BUF_X1 U51 ( .A(N11), .Z(n243) );
  BUF_X1 U52 ( .A(N11), .Z(n244) );
  INV_X1 U53 ( .A(N10), .ZN(n251) );
  BUF_X1 U54 ( .A(N12), .Z(n241) );
  NOR3_X1 U55 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U56 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U57 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U58 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U59 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U60 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U61 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U62 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U63 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U64 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U65 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U67 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U69 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U70 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U71 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U72 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U73 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U74 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U75 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U76 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U77 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U79 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U81 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U82 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U83 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U84 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U85 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U86 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U87 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U88 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U89 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U90 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U91 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U92 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U93 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U94 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U95 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U96 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U97 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U98 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U99 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U100 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U101 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U102 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U103 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U104 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U105 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U106 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U107 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U108 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U109 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U110 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U111 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U112 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U113 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U114 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U115 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U116 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U117 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U118 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U119 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U120 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U121 ( .A(n988), .ZN(n705) );
  AOI22_X1 U122 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U123 ( .A(n986), .ZN(n704) );
  AOI22_X1 U124 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U125 ( .A(n985), .ZN(n703) );
  AOI22_X1 U126 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U127 ( .A(n984), .ZN(n702) );
  AOI22_X1 U128 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U129 ( .A(n983), .ZN(n701) );
  AOI22_X1 U130 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U131 ( .A(n982), .ZN(n700) );
  AOI22_X1 U132 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U133 ( .A(n981), .ZN(n699) );
  AOI22_X1 U134 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U135 ( .A(n980), .ZN(n698) );
  AOI22_X1 U136 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U137 ( .A(n951), .ZN(n673) );
  AOI22_X1 U138 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U139 ( .A(n949), .ZN(n672) );
  AOI22_X1 U140 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U141 ( .A(n948), .ZN(n671) );
  AOI22_X1 U142 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U143 ( .A(n947), .ZN(n670) );
  AOI22_X1 U144 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U145 ( .A(n946), .ZN(n669) );
  AOI22_X1 U146 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U147 ( .A(n945), .ZN(n668) );
  AOI22_X1 U148 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U149 ( .A(n944), .ZN(n667) );
  AOI22_X1 U150 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U151 ( .A(n943), .ZN(n666) );
  AOI22_X1 U152 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U153 ( .A(n915), .ZN(n641) );
  AOI22_X1 U154 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U155 ( .A(n913), .ZN(n640) );
  AOI22_X1 U156 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U157 ( .A(n912), .ZN(n639) );
  AOI22_X1 U158 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U159 ( .A(n911), .ZN(n638) );
  AOI22_X1 U160 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U161 ( .A(n910), .ZN(n637) );
  AOI22_X1 U162 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U163 ( .A(n909), .ZN(n636) );
  AOI22_X1 U164 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U165 ( .A(n908), .ZN(n635) );
  AOI22_X1 U166 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U167 ( .A(n907), .ZN(n634) );
  AOI22_X1 U168 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U169 ( .A(n935), .ZN(n659) );
  AOI22_X1 U170 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U171 ( .A(n934), .ZN(n658) );
  AOI22_X1 U172 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U173 ( .A(n933), .ZN(n657) );
  AOI22_X1 U174 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U175 ( .A(n931), .ZN(n656) );
  AOI22_X1 U176 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U177 ( .A(n930), .ZN(n655) );
  AOI22_X1 U178 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U179 ( .A(n929), .ZN(n654) );
  AOI22_X1 U180 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U181 ( .A(n928), .ZN(n653) );
  AOI22_X1 U182 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U183 ( .A(n927), .ZN(n652) );
  AOI22_X1 U184 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U185 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U186 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U187 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U188 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U189 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U190 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U191 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U192 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U193 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U194 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U195 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U196 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U197 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U198 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U199 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U200 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U201 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U202 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U203 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U204 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U205 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U206 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U207 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U208 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U209 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U210 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U211 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U212 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U213 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U214 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U215 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U216 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U217 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U218 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U219 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U220 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U221 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U222 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U223 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U224 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U225 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U226 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U227 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U228 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U229 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U230 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U231 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U232 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U233 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U234 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U235 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U236 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U237 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U238 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U239 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U240 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U241 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U242 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U243 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U244 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U245 ( .A(n972), .ZN(n691) );
  AOI22_X1 U246 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U247 ( .A(n971), .ZN(n690) );
  AOI22_X1 U248 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U249 ( .A(n970), .ZN(n689) );
  AOI22_X1 U250 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U251 ( .A(n968), .ZN(n688) );
  AOI22_X1 U252 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U253 ( .A(n967), .ZN(n687) );
  AOI22_X1 U254 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U255 ( .A(n966), .ZN(n686) );
  AOI22_X1 U256 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U257 ( .A(n965), .ZN(n685) );
  AOI22_X1 U258 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U259 ( .A(n964), .ZN(n684) );
  AOI22_X1 U260 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U261 ( .A(n963), .ZN(n683) );
  AOI22_X1 U262 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U263 ( .A(n962), .ZN(n682) );
  AOI22_X1 U264 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U265 ( .A(n942), .ZN(n665) );
  AOI22_X1 U266 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U267 ( .A(n940), .ZN(n664) );
  AOI22_X1 U268 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U269 ( .A(n939), .ZN(n663) );
  AOI22_X1 U270 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U271 ( .A(n938), .ZN(n662) );
  AOI22_X1 U272 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U273 ( .A(n937), .ZN(n661) );
  AOI22_X1 U274 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U275 ( .A(n936), .ZN(n660) );
  AOI22_X1 U276 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U277 ( .A(n926), .ZN(n651) );
  AOI22_X1 U278 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U279 ( .A(n925), .ZN(n650) );
  AOI22_X1 U280 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U281 ( .A(n906), .ZN(n633) );
  AOI22_X1 U282 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U283 ( .A(n904), .ZN(n632) );
  AOI22_X1 U284 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U285 ( .A(n903), .ZN(n631) );
  AOI22_X1 U286 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U287 ( .A(n902), .ZN(n630) );
  AOI22_X1 U288 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U289 ( .A(n901), .ZN(n629) );
  AOI22_X1 U290 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U291 ( .A(n900), .ZN(n628) );
  AOI22_X1 U292 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U293 ( .A(n899), .ZN(n627) );
  AOI22_X1 U294 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U295 ( .A(n898), .ZN(n626) );
  AOI22_X1 U296 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U297 ( .A(n897), .ZN(n625) );
  AOI22_X1 U298 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U299 ( .A(n895), .ZN(n624) );
  AOI22_X1 U300 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U301 ( .A(n894), .ZN(n623) );
  AOI22_X1 U302 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U303 ( .A(n893), .ZN(n622) );
  AOI22_X1 U304 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U305 ( .A(n892), .ZN(n621) );
  AOI22_X1 U306 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U307 ( .A(n891), .ZN(n620) );
  AOI22_X1 U308 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U309 ( .A(n890), .ZN(n619) );
  AOI22_X1 U310 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U311 ( .A(n889), .ZN(n618) );
  AOI22_X1 U312 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U313 ( .A(n999), .ZN(n715) );
  AOI22_X1 U314 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U315 ( .A(n998), .ZN(n714) );
  AOI22_X1 U316 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U317 ( .A(n979), .ZN(n697) );
  AOI22_X1 U318 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U319 ( .A(n977), .ZN(n696) );
  AOI22_X1 U320 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U321 ( .A(n976), .ZN(n695) );
  AOI22_X1 U322 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U323 ( .A(n975), .ZN(n694) );
  AOI22_X1 U324 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U325 ( .A(n974), .ZN(n693) );
  AOI22_X1 U326 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U327 ( .A(n973), .ZN(n692) );
  AOI22_X1 U328 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U329 ( .A(N12), .ZN(n253) );
  INV_X1 U330 ( .A(N11), .ZN(n252) );
  INV_X1 U331 ( .A(n997), .ZN(n713) );
  AOI22_X1 U332 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U333 ( .A(n995), .ZN(n712) );
  AOI22_X1 U334 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U335 ( .A(n994), .ZN(n711) );
  AOI22_X1 U336 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U337 ( .A(n993), .ZN(n710) );
  AOI22_X1 U338 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U339 ( .A(n992), .ZN(n709) );
  AOI22_X1 U340 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U341 ( .A(n991), .ZN(n708) );
  AOI22_X1 U342 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U343 ( .A(n990), .ZN(n707) );
  AOI22_X1 U344 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U345 ( .A(n989), .ZN(n706) );
  AOI22_X1 U346 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U347 ( .A(n924), .ZN(n649) );
  AOI22_X1 U348 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U349 ( .A(n922), .ZN(n648) );
  AOI22_X1 U350 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U351 ( .A(n921), .ZN(n647) );
  AOI22_X1 U352 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U353 ( .A(n920), .ZN(n646) );
  AOI22_X1 U354 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U355 ( .A(n919), .ZN(n645) );
  AOI22_X1 U356 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U357 ( .A(n918), .ZN(n644) );
  AOI22_X1 U358 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U359 ( .A(n917), .ZN(n643) );
  AOI22_X1 U360 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U361 ( .A(n916), .ZN(n642) );
  AOI22_X1 U362 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U363 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U364 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U365 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U366 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U367 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U368 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U369 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U370 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U371 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U372 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U373 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U374 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U375 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U376 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U377 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U378 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U379 ( .A(n961), .ZN(n681) );
  AOI22_X1 U380 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U381 ( .A(n959), .ZN(n680) );
  AOI22_X1 U382 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U383 ( .A(n958), .ZN(n679) );
  AOI22_X1 U384 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U385 ( .A(n957), .ZN(n678) );
  AOI22_X1 U386 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U387 ( .A(n956), .ZN(n677) );
  AOI22_X1 U388 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U389 ( .A(n955), .ZN(n676) );
  AOI22_X1 U390 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U391 ( .A(n954), .ZN(n675) );
  AOI22_X1 U392 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U393 ( .A(n953), .ZN(n674) );
  AOI22_X1 U394 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U395 ( .A(n888), .ZN(n617) );
  AOI22_X1 U396 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U397 ( .A(n886), .ZN(n616) );
  AOI22_X1 U398 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U399 ( .A(n885), .ZN(n615) );
  AOI22_X1 U400 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U401 ( .A(n884), .ZN(n614) );
  AOI22_X1 U402 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U403 ( .A(n883), .ZN(n613) );
  AOI22_X1 U404 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U405 ( .A(n882), .ZN(n612) );
  AOI22_X1 U406 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U407 ( .A(n881), .ZN(n611) );
  AOI22_X1 U408 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U409 ( .A(n880), .ZN(n610) );
  AOI22_X1 U410 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U411 ( .A(n879), .ZN(n609) );
  AOI22_X1 U412 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U413 ( .A(n877), .ZN(n608) );
  AOI22_X1 U414 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U415 ( .A(n876), .ZN(n607) );
  AOI22_X1 U416 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U417 ( .A(n875), .ZN(n606) );
  AOI22_X1 U418 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U419 ( .A(n874), .ZN(n605) );
  AOI22_X1 U420 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U421 ( .A(n873), .ZN(n604) );
  AOI22_X1 U422 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U423 ( .A(n872), .ZN(n603) );
  AOI22_X1 U424 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U425 ( .A(n871), .ZN(n602) );
  AOI22_X1 U426 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U427 ( .A(n870), .ZN(n601) );
  AOI22_X1 U428 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U429 ( .A(n868), .ZN(n600) );
  AOI22_X1 U430 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U431 ( .A(n867), .ZN(n599) );
  AOI22_X1 U432 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U433 ( .A(n866), .ZN(n598) );
  AOI22_X1 U434 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U435 ( .A(n865), .ZN(n597) );
  AOI22_X1 U436 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U437 ( .A(n864), .ZN(n596) );
  AOI22_X1 U438 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U439 ( .A(n863), .ZN(n595) );
  AOI22_X1 U440 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U441 ( .A(n862), .ZN(n594) );
  AOI22_X1 U442 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U443 ( .A(n861), .ZN(n293) );
  AOI22_X1 U444 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U445 ( .A(n859), .ZN(n292) );
  AOI22_X1 U446 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U447 ( .A(n858), .ZN(n291) );
  AOI22_X1 U448 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U449 ( .A(n857), .ZN(n290) );
  AOI22_X1 U450 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U451 ( .A(n856), .ZN(n289) );
  AOI22_X1 U452 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U453 ( .A(n855), .ZN(n288) );
  AOI22_X1 U454 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U455 ( .A(n854), .ZN(n287) );
  AOI22_X1 U456 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U457 ( .A(n853), .ZN(n286) );
  AOI22_X1 U458 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U459 ( .A(n852), .ZN(n285) );
  AOI22_X1 U460 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U461 ( .A(n850), .ZN(n284) );
  AOI22_X1 U462 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U463 ( .A(n849), .ZN(n283) );
  AOI22_X1 U464 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U465 ( .A(n848), .ZN(n282) );
  AOI22_X1 U466 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U467 ( .A(n847), .ZN(n281) );
  AOI22_X1 U468 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U469 ( .A(n846), .ZN(n280) );
  AOI22_X1 U470 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U471 ( .A(n845), .ZN(n279) );
  AOI22_X1 U472 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U473 ( .A(n844), .ZN(n278) );
  AOI22_X1 U474 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U475 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U476 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U477 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U478 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U479 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U480 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U481 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U482 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U483 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U484 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U485 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U486 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U487 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U488 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U489 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U490 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U491 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U492 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U493 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U494 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U495 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U496 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U497 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U498 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U499 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U500 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U501 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U502 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U503 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U504 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U505 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U506 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U507 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U508 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U509 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U510 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U511 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U512 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U513 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U514 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U515 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U516 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U517 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U518 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U519 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U520 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U521 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U522 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U523 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U524 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U525 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U526 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U527 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U528 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U529 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U530 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U531 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U532 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U533 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U534 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U535 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U536 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U537 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U538 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U539 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U540 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U541 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U542 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U543 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U544 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U545 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U546 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U547 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U548 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U549 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U550 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U551 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U552 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U553 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U554 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U555 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U556 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U557 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U558 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U559 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U560 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U561 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U562 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U563 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U564 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U565 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U566 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U567 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U568 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U569 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U570 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U571 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U572 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U573 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U574 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U575 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U576 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U577 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U578 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U579 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U580 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U581 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U582 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U583 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U584 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U585 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U586 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U587 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U588 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U589 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U590 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U591 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U592 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U593 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U594 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U595 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U596 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U597 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U598 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U599 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U600 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U601 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U602 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U603 ( .A(N13), .ZN(n842) );
  INV_X1 U604 ( .A(N14), .ZN(n843) );
  MUX2_X1 U605 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n249), .Z(n1) );
  MUX2_X1 U606 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n249), .Z(n2) );
  MUX2_X1 U607 ( .A(n2), .B(n1), .S(n242), .Z(n3) );
  MUX2_X1 U608 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n249), .Z(n4) );
  MUX2_X1 U609 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n248), .Z(n5) );
  MUX2_X1 U610 ( .A(n5), .B(n4), .S(n242), .Z(n6) );
  MUX2_X1 U611 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U612 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n249), .Z(n8) );
  MUX2_X1 U613 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n248), .Z(n9) );
  MUX2_X1 U614 ( .A(n9), .B(n8), .S(n242), .Z(n10) );
  MUX2_X1 U615 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n249), .Z(n11) );
  MUX2_X1 U616 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n248), .Z(n12) );
  MUX2_X1 U617 ( .A(n12), .B(n11), .S(n242), .Z(n13) );
  MUX2_X1 U618 ( .A(n13), .B(n10), .S(N12), .Z(n14) );
  MUX2_X1 U619 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U620 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n245), .Z(n16) );
  MUX2_X1 U621 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n245), .Z(n17) );
  MUX2_X1 U622 ( .A(n17), .B(n16), .S(n243), .Z(n18) );
  MUX2_X1 U623 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U624 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n245), .Z(n20) );
  MUX2_X1 U625 ( .A(n20), .B(n19), .S(n243), .Z(n21) );
  MUX2_X1 U626 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U627 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n245), .Z(n23) );
  MUX2_X1 U628 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n245), .Z(n24) );
  MUX2_X1 U629 ( .A(n24), .B(n23), .S(n243), .Z(n25) );
  MUX2_X1 U630 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n245), .Z(n26) );
  MUX2_X1 U631 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n245), .Z(n27) );
  MUX2_X1 U632 ( .A(n27), .B(n26), .S(n243), .Z(n28) );
  MUX2_X1 U633 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U634 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U635 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U636 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n245), .Z(n31) );
  MUX2_X1 U637 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n245), .Z(n32) );
  MUX2_X1 U638 ( .A(n32), .B(n31), .S(n243), .Z(n33) );
  MUX2_X1 U639 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U640 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U641 ( .A(n35), .B(n34), .S(n243), .Z(n36) );
  MUX2_X1 U642 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U643 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n246), .Z(n38) );
  MUX2_X1 U644 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n246), .Z(n39) );
  MUX2_X1 U645 ( .A(n39), .B(n38), .S(n243), .Z(n40) );
  MUX2_X1 U646 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n246), .Z(n41) );
  MUX2_X1 U647 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n246), .Z(n42) );
  MUX2_X1 U648 ( .A(n42), .B(n41), .S(n243), .Z(n43) );
  MUX2_X1 U649 ( .A(n43), .B(n40), .S(n241), .Z(n44) );
  MUX2_X1 U650 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U651 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n246), .Z(n46) );
  MUX2_X1 U652 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n246), .Z(n47) );
  MUX2_X1 U653 ( .A(n47), .B(n46), .S(n243), .Z(n48) );
  MUX2_X1 U654 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n246), .Z(n49) );
  MUX2_X1 U655 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n246), .Z(n50) );
  MUX2_X1 U656 ( .A(n50), .B(n49), .S(n243), .Z(n51) );
  MUX2_X1 U657 ( .A(n51), .B(n48), .S(n241), .Z(n52) );
  MUX2_X1 U658 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n246), .Z(n53) );
  MUX2_X1 U659 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n246), .Z(n54) );
  MUX2_X1 U660 ( .A(n54), .B(n53), .S(n243), .Z(n55) );
  MUX2_X1 U661 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n246), .Z(n56) );
  MUX2_X1 U662 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n246), .Z(n57) );
  MUX2_X1 U663 ( .A(n57), .B(n56), .S(n243), .Z(n58) );
  MUX2_X1 U664 ( .A(n58), .B(n55), .S(n241), .Z(n59) );
  MUX2_X1 U665 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U666 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U667 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n247), .Z(n61) );
  MUX2_X1 U668 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n247), .Z(n62) );
  MUX2_X1 U669 ( .A(n62), .B(n61), .S(n244), .Z(n63) );
  MUX2_X1 U670 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n247), .Z(n64) );
  MUX2_X1 U671 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n247), .Z(n65) );
  MUX2_X1 U672 ( .A(n65), .B(n64), .S(n244), .Z(n66) );
  MUX2_X1 U673 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U674 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n247), .Z(n68) );
  MUX2_X1 U675 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n247), .Z(n69) );
  MUX2_X1 U676 ( .A(n69), .B(n68), .S(n244), .Z(n70) );
  MUX2_X1 U677 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n247), .Z(n71) );
  MUX2_X1 U678 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n247), .Z(n72) );
  MUX2_X1 U679 ( .A(n72), .B(n71), .S(n244), .Z(n73) );
  MUX2_X1 U680 ( .A(n73), .B(n70), .S(n241), .Z(n74) );
  MUX2_X1 U681 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U682 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n247), .Z(n76) );
  MUX2_X1 U683 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n247), .Z(n77) );
  MUX2_X1 U684 ( .A(n77), .B(n76), .S(n244), .Z(n78) );
  MUX2_X1 U685 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n247), .Z(n79) );
  MUX2_X1 U686 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n247), .Z(n80) );
  MUX2_X1 U687 ( .A(n80), .B(n79), .S(n244), .Z(n81) );
  MUX2_X1 U688 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U689 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n246), .Z(n83) );
  MUX2_X1 U690 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n247), .Z(n84) );
  MUX2_X1 U691 ( .A(n84), .B(n83), .S(n244), .Z(n85) );
  MUX2_X1 U692 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n246), .Z(n86) );
  MUX2_X1 U693 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n246), .Z(n87) );
  MUX2_X1 U694 ( .A(n87), .B(n86), .S(n244), .Z(n88) );
  MUX2_X1 U695 ( .A(n88), .B(n85), .S(n241), .Z(n89) );
  MUX2_X1 U696 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U697 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U698 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n247), .Z(n91) );
  MUX2_X1 U699 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n92) );
  MUX2_X1 U700 ( .A(n92), .B(n91), .S(n244), .Z(n93) );
  MUX2_X1 U701 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U702 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n247), .Z(n95) );
  MUX2_X1 U703 ( .A(n95), .B(n94), .S(n244), .Z(n96) );
  MUX2_X1 U704 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U705 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n98) );
  MUX2_X1 U706 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n248), .Z(n99) );
  MUX2_X1 U707 ( .A(n99), .B(n98), .S(n244), .Z(n100) );
  MUX2_X1 U708 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n245), .Z(n101) );
  MUX2_X1 U709 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n248), .Z(n102) );
  MUX2_X1 U710 ( .A(n102), .B(n101), .S(n244), .Z(n103) );
  MUX2_X1 U711 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U712 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U713 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n249), .Z(n106) );
  MUX2_X1 U714 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n250), .Z(n107) );
  MUX2_X1 U715 ( .A(n107), .B(n106), .S(N11), .Z(n108) );
  MUX2_X1 U716 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n249), .Z(n109) );
  MUX2_X1 U717 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n110) );
  MUX2_X1 U718 ( .A(n110), .B(n109), .S(N11), .Z(n111) );
  MUX2_X1 U719 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U720 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n250), .Z(n113) );
  MUX2_X1 U721 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n114) );
  MUX2_X1 U722 ( .A(n114), .B(n113), .S(N11), .Z(n115) );
  MUX2_X1 U723 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n116) );
  MUX2_X1 U724 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n117) );
  MUX2_X1 U725 ( .A(n117), .B(n116), .S(n244), .Z(n118) );
  MUX2_X1 U726 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U727 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U728 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U729 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n249), .Z(n121) );
  MUX2_X1 U730 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(N10), .Z(n122) );
  MUX2_X1 U731 ( .A(n122), .B(n121), .S(n244), .Z(n123) );
  MUX2_X1 U732 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n249), .Z(n124) );
  MUX2_X1 U733 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n125) );
  MUX2_X1 U734 ( .A(n125), .B(n124), .S(N11), .Z(n126) );
  MUX2_X1 U735 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U736 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n248), .Z(n128) );
  MUX2_X1 U737 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n248), .Z(n129) );
  MUX2_X1 U738 ( .A(n129), .B(n128), .S(N11), .Z(n130) );
  MUX2_X1 U739 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n248), .Z(n131) );
  MUX2_X1 U740 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n248), .Z(n132) );
  MUX2_X1 U741 ( .A(n132), .B(n131), .S(n242), .Z(n133) );
  MUX2_X1 U742 ( .A(n133), .B(n130), .S(n241), .Z(n134) );
  MUX2_X1 U743 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U744 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n248), .Z(n136) );
  MUX2_X1 U745 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n248), .Z(n137) );
  MUX2_X1 U746 ( .A(n137), .B(n136), .S(N11), .Z(n138) );
  MUX2_X1 U747 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n248), .Z(n139) );
  MUX2_X1 U748 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n248), .Z(n140) );
  MUX2_X1 U749 ( .A(n140), .B(n139), .S(n244), .Z(n141) );
  MUX2_X1 U750 ( .A(n141), .B(n138), .S(n241), .Z(n142) );
  MUX2_X1 U751 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n248), .Z(n143) );
  MUX2_X1 U752 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n248), .Z(n144) );
  MUX2_X1 U753 ( .A(n144), .B(n143), .S(N11), .Z(n145) );
  MUX2_X1 U754 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n248), .Z(n146) );
  MUX2_X1 U755 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n248), .Z(n147) );
  MUX2_X1 U756 ( .A(n147), .B(n146), .S(n243), .Z(n148) );
  MUX2_X1 U757 ( .A(n148), .B(n145), .S(n241), .Z(n149) );
  MUX2_X1 U758 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U759 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U760 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n249), .Z(n151) );
  MUX2_X1 U761 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n249), .Z(n152) );
  MUX2_X1 U762 ( .A(n152), .B(n151), .S(n244), .Z(n153) );
  MUX2_X1 U763 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n249), .Z(n154) );
  MUX2_X1 U764 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n249), .Z(n155) );
  MUX2_X1 U765 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U766 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U767 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n249), .Z(n158) );
  MUX2_X1 U768 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n249), .Z(n159) );
  MUX2_X1 U769 ( .A(n159), .B(n158), .S(n242), .Z(n160) );
  MUX2_X1 U770 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n249), .Z(n161) );
  MUX2_X1 U771 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n249), .Z(n162) );
  MUX2_X1 U772 ( .A(n162), .B(n161), .S(N11), .Z(n163) );
  MUX2_X1 U773 ( .A(n163), .B(n160), .S(N12), .Z(n164) );
  MUX2_X1 U774 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U775 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n249), .Z(n166) );
  MUX2_X1 U776 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n249), .Z(n167) );
  MUX2_X1 U777 ( .A(n167), .B(n166), .S(n243), .Z(n168) );
  MUX2_X1 U778 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n249), .Z(n169) );
  MUX2_X1 U779 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n249), .Z(n170) );
  MUX2_X1 U780 ( .A(n170), .B(n169), .S(N11), .Z(n171) );
  MUX2_X1 U781 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U782 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n250), .Z(n173) );
  MUX2_X1 U783 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n245), .Z(n174) );
  MUX2_X1 U784 ( .A(n174), .B(n173), .S(n242), .Z(n175) );
  MUX2_X1 U785 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n247), .Z(n176) );
  MUX2_X1 U786 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n250), .Z(n177) );
  MUX2_X1 U787 ( .A(n177), .B(n176), .S(N11), .Z(n178) );
  MUX2_X1 U788 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U789 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U790 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U791 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n246), .Z(n181) );
  MUX2_X1 U792 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n245), .Z(n182) );
  MUX2_X1 U793 ( .A(n182), .B(n181), .S(n243), .Z(n183) );
  MUX2_X1 U794 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n250), .Z(n184) );
  MUX2_X1 U795 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n250), .Z(n185) );
  MUX2_X1 U796 ( .A(n185), .B(n184), .S(n243), .Z(n186) );
  MUX2_X1 U797 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U798 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n246), .Z(n188) );
  MUX2_X1 U799 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n250), .Z(n189) );
  MUX2_X1 U800 ( .A(n189), .B(n188), .S(n244), .Z(n190) );
  MUX2_X1 U801 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n250), .Z(n191) );
  MUX2_X1 U802 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n250), .Z(n192) );
  MUX2_X1 U803 ( .A(n192), .B(n191), .S(N11), .Z(n193) );
  MUX2_X1 U804 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U805 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U806 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n249), .Z(n196) );
  MUX2_X1 U807 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(N10), .Z(n197) );
  MUX2_X1 U808 ( .A(n197), .B(n196), .S(n242), .Z(n198) );
  MUX2_X1 U809 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n249), .Z(n199) );
  MUX2_X1 U810 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n250), .Z(n200) );
  MUX2_X1 U811 ( .A(n200), .B(n199), .S(n244), .Z(n201) );
  MUX2_X1 U812 ( .A(n201), .B(n198), .S(N12), .Z(n202) );
  MUX2_X1 U813 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n203) );
  MUX2_X1 U814 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n250), .Z(n204) );
  MUX2_X1 U815 ( .A(n204), .B(n203), .S(n242), .Z(n205) );
  MUX2_X1 U816 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n250), .Z(n206) );
  MUX2_X1 U817 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n250), .Z(n207) );
  MUX2_X1 U818 ( .A(n207), .B(n206), .S(n243), .Z(n208) );
  MUX2_X1 U819 ( .A(n208), .B(n205), .S(N12), .Z(n209) );
  MUX2_X1 U820 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U821 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U822 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n245), .Z(n211) );
  MUX2_X1 U823 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n247), .Z(n212) );
  MUX2_X1 U824 ( .A(n212), .B(n211), .S(n242), .Z(n213) );
  MUX2_X1 U825 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n248), .Z(n214) );
  MUX2_X1 U826 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(N10), .Z(n215) );
  MUX2_X1 U827 ( .A(n215), .B(n214), .S(n242), .Z(n216) );
  MUX2_X1 U828 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U829 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n247), .Z(n218) );
  MUX2_X1 U830 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n250), .Z(n219) );
  MUX2_X1 U831 ( .A(n219), .B(n218), .S(n242), .Z(n220) );
  MUX2_X1 U832 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n246), .Z(n221) );
  MUX2_X1 U833 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n222) );
  MUX2_X1 U834 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U835 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U836 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U837 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n250), .Z(n226) );
  MUX2_X1 U838 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n245), .Z(n227) );
  MUX2_X1 U839 ( .A(n227), .B(n226), .S(n242), .Z(n228) );
  MUX2_X1 U840 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n250), .Z(n229) );
  MUX2_X1 U841 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n230) );
  MUX2_X1 U842 ( .A(n230), .B(n229), .S(n243), .Z(n231) );
  MUX2_X1 U843 ( .A(n231), .B(n228), .S(N12), .Z(n232) );
  MUX2_X1 U844 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n250), .Z(n233) );
  MUX2_X1 U845 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n234) );
  MUX2_X1 U846 ( .A(n234), .B(n233), .S(n242), .Z(n235) );
  MUX2_X1 U847 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n236) );
  MUX2_X1 U848 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n237) );
  MUX2_X1 U849 ( .A(n237), .B(n236), .S(n242), .Z(n238) );
  MUX2_X1 U850 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U851 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U852 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U853 ( .A(N11), .Z(n242) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_22 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(N10), .Z(n247) );
  BUF_X1 U4 ( .A(n250), .Z(n248) );
  BUF_X1 U5 ( .A(n250), .Z(n249) );
  BUF_X1 U6 ( .A(n250), .Z(n246) );
  BUF_X1 U7 ( .A(n250), .Z(n245) );
  BUF_X1 U8 ( .A(N10), .Z(n250) );
  INV_X1 U9 ( .A(n1111), .ZN(n841) );
  INV_X1 U10 ( .A(n1100), .ZN(n840) );
  INV_X1 U11 ( .A(n1090), .ZN(n839) );
  INV_X1 U12 ( .A(n1080), .ZN(n838) );
  INV_X1 U13 ( .A(n1070), .ZN(n837) );
  INV_X1 U14 ( .A(n1060), .ZN(n836) );
  INV_X1 U15 ( .A(n1051), .ZN(n835) );
  INV_X1 U16 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U19 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U20 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U21 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U22 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U23 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U24 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U26 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U27 ( .A(n1131), .ZN(n816) );
  INV_X1 U28 ( .A(n1121), .ZN(n815) );
  INV_X1 U29 ( .A(n887), .ZN(n814) );
  INV_X1 U30 ( .A(n878), .ZN(n813) );
  INV_X1 U31 ( .A(n869), .ZN(n812) );
  INV_X1 U32 ( .A(n860), .ZN(n811) );
  INV_X1 U33 ( .A(n851), .ZN(n810) );
  INV_X1 U34 ( .A(n987), .ZN(n828) );
  INV_X1 U35 ( .A(n978), .ZN(n827) );
  INV_X1 U36 ( .A(n969), .ZN(n826) );
  INV_X1 U37 ( .A(n914), .ZN(n820) );
  INV_X1 U38 ( .A(n905), .ZN(n819) );
  INV_X1 U39 ( .A(n896), .ZN(n818) );
  INV_X1 U40 ( .A(n1033), .ZN(n833) );
  INV_X1 U41 ( .A(n1023), .ZN(n832) );
  INV_X1 U42 ( .A(n1014), .ZN(n831) );
  INV_X1 U43 ( .A(n1005), .ZN(n830) );
  INV_X1 U44 ( .A(n996), .ZN(n829) );
  INV_X1 U45 ( .A(n960), .ZN(n825) );
  INV_X1 U46 ( .A(n950), .ZN(n824) );
  INV_X1 U47 ( .A(n941), .ZN(n823) );
  INV_X1 U48 ( .A(n932), .ZN(n822) );
  INV_X1 U49 ( .A(n923), .ZN(n821) );
  INV_X1 U50 ( .A(n1142), .ZN(n817) );
  BUF_X1 U51 ( .A(N11), .Z(n243) );
  BUF_X1 U52 ( .A(N11), .Z(n244) );
  INV_X1 U53 ( .A(N10), .ZN(n251) );
  BUF_X1 U54 ( .A(N12), .Z(n241) );
  NOR3_X1 U55 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U56 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U57 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U58 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U59 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U60 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U61 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U62 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U63 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U64 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U65 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U67 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U69 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U70 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U71 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U72 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U73 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U74 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U75 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U76 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U77 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U79 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U81 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U82 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U83 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U84 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U85 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U86 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U87 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U88 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U89 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U90 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U91 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U92 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U93 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U94 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U95 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U96 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U97 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U98 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U99 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U100 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U101 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U102 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U103 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U104 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U105 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U106 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U107 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U108 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U109 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U110 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U111 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U112 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U113 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U114 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U115 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U116 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U117 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U118 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U119 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U120 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U121 ( .A(n988), .ZN(n705) );
  AOI22_X1 U122 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U123 ( .A(n986), .ZN(n704) );
  AOI22_X1 U124 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U125 ( .A(n985), .ZN(n703) );
  AOI22_X1 U126 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U127 ( .A(n984), .ZN(n702) );
  AOI22_X1 U128 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U129 ( .A(n983), .ZN(n701) );
  AOI22_X1 U130 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U131 ( .A(n982), .ZN(n700) );
  AOI22_X1 U132 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U133 ( .A(n981), .ZN(n699) );
  AOI22_X1 U134 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U135 ( .A(n980), .ZN(n698) );
  AOI22_X1 U136 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U137 ( .A(n943), .ZN(n666) );
  AOI22_X1 U138 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U139 ( .A(n915), .ZN(n641) );
  AOI22_X1 U140 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U141 ( .A(n913), .ZN(n640) );
  AOI22_X1 U142 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U143 ( .A(n912), .ZN(n639) );
  AOI22_X1 U144 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U145 ( .A(n911), .ZN(n638) );
  AOI22_X1 U146 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U147 ( .A(n910), .ZN(n637) );
  AOI22_X1 U148 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U149 ( .A(n909), .ZN(n636) );
  AOI22_X1 U150 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U151 ( .A(n908), .ZN(n635) );
  AOI22_X1 U152 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U153 ( .A(n907), .ZN(n634) );
  AOI22_X1 U154 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U155 ( .A(n942), .ZN(n665) );
  AOI22_X1 U156 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U157 ( .A(n940), .ZN(n664) );
  AOI22_X1 U158 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U159 ( .A(n939), .ZN(n663) );
  AOI22_X1 U160 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U161 ( .A(n938), .ZN(n662) );
  AOI22_X1 U162 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U163 ( .A(n937), .ZN(n661) );
  AOI22_X1 U164 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U165 ( .A(n936), .ZN(n660) );
  AOI22_X1 U166 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U167 ( .A(n935), .ZN(n659) );
  AOI22_X1 U168 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U169 ( .A(n934), .ZN(n658) );
  AOI22_X1 U170 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U171 ( .A(n933), .ZN(n657) );
  AOI22_X1 U172 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U173 ( .A(n931), .ZN(n656) );
  AOI22_X1 U174 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U175 ( .A(n930), .ZN(n655) );
  AOI22_X1 U176 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U177 ( .A(n929), .ZN(n654) );
  AOI22_X1 U178 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U179 ( .A(n928), .ZN(n653) );
  AOI22_X1 U180 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U181 ( .A(n927), .ZN(n652) );
  AOI22_X1 U182 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U183 ( .A(n926), .ZN(n651) );
  AOI22_X1 U184 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U185 ( .A(n925), .ZN(n650) );
  AOI22_X1 U186 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U187 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U188 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U189 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U190 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U191 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U192 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U193 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U194 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U195 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U196 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U197 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U198 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U199 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U200 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U201 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U202 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U203 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U204 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U205 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U206 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U207 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U208 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U209 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U210 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U211 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U212 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U213 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U214 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U215 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U216 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U217 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U218 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U219 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U220 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U221 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U222 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U223 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U224 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U225 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U226 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U227 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U228 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U229 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U230 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U231 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U232 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U233 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U234 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U235 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U236 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U237 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U238 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U239 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U240 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U241 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U242 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U243 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U244 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U245 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U246 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U247 ( .A(n999), .ZN(n715) );
  AOI22_X1 U248 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U249 ( .A(n998), .ZN(n714) );
  AOI22_X1 U250 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U251 ( .A(n951), .ZN(n673) );
  AOI22_X1 U252 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U253 ( .A(n949), .ZN(n672) );
  AOI22_X1 U254 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U255 ( .A(n948), .ZN(n671) );
  AOI22_X1 U256 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U257 ( .A(n947), .ZN(n670) );
  AOI22_X1 U258 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U259 ( .A(n946), .ZN(n669) );
  AOI22_X1 U260 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U261 ( .A(n945), .ZN(n668) );
  AOI22_X1 U262 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U263 ( .A(n944), .ZN(n667) );
  AOI22_X1 U264 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U265 ( .A(n979), .ZN(n697) );
  AOI22_X1 U266 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U267 ( .A(n977), .ZN(n696) );
  AOI22_X1 U268 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U269 ( .A(n976), .ZN(n695) );
  AOI22_X1 U270 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U271 ( .A(n975), .ZN(n694) );
  AOI22_X1 U272 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U273 ( .A(n974), .ZN(n693) );
  AOI22_X1 U274 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U275 ( .A(n973), .ZN(n692) );
  AOI22_X1 U276 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U277 ( .A(n972), .ZN(n691) );
  AOI22_X1 U278 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U279 ( .A(n971), .ZN(n690) );
  AOI22_X1 U280 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U281 ( .A(n970), .ZN(n689) );
  AOI22_X1 U282 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U283 ( .A(n968), .ZN(n688) );
  AOI22_X1 U284 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U285 ( .A(n967), .ZN(n687) );
  AOI22_X1 U286 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U287 ( .A(n966), .ZN(n686) );
  AOI22_X1 U288 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U289 ( .A(n965), .ZN(n685) );
  AOI22_X1 U290 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U291 ( .A(n964), .ZN(n684) );
  AOI22_X1 U292 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U293 ( .A(n963), .ZN(n683) );
  AOI22_X1 U294 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U295 ( .A(n962), .ZN(n682) );
  AOI22_X1 U296 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U297 ( .A(n906), .ZN(n633) );
  AOI22_X1 U298 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U299 ( .A(n904), .ZN(n632) );
  AOI22_X1 U300 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U301 ( .A(n903), .ZN(n631) );
  AOI22_X1 U302 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U303 ( .A(n902), .ZN(n630) );
  AOI22_X1 U304 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U305 ( .A(n901), .ZN(n629) );
  AOI22_X1 U306 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U307 ( .A(n900), .ZN(n628) );
  AOI22_X1 U308 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U309 ( .A(n899), .ZN(n627) );
  AOI22_X1 U310 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U311 ( .A(n898), .ZN(n626) );
  AOI22_X1 U312 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U313 ( .A(n897), .ZN(n625) );
  AOI22_X1 U314 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U315 ( .A(n895), .ZN(n624) );
  AOI22_X1 U316 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U317 ( .A(n894), .ZN(n623) );
  AOI22_X1 U318 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U319 ( .A(n893), .ZN(n622) );
  AOI22_X1 U320 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U321 ( .A(n892), .ZN(n621) );
  AOI22_X1 U322 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U323 ( .A(n891), .ZN(n620) );
  AOI22_X1 U324 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U325 ( .A(n890), .ZN(n619) );
  AOI22_X1 U326 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U327 ( .A(n889), .ZN(n618) );
  AOI22_X1 U328 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U329 ( .A(N12), .ZN(n253) );
  INV_X1 U330 ( .A(N11), .ZN(n252) );
  INV_X1 U331 ( .A(n997), .ZN(n713) );
  AOI22_X1 U332 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U333 ( .A(n995), .ZN(n712) );
  AOI22_X1 U334 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U335 ( .A(n994), .ZN(n711) );
  AOI22_X1 U336 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U337 ( .A(n993), .ZN(n710) );
  AOI22_X1 U338 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U339 ( .A(n992), .ZN(n709) );
  AOI22_X1 U340 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U341 ( .A(n991), .ZN(n708) );
  AOI22_X1 U342 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U343 ( .A(n990), .ZN(n707) );
  AOI22_X1 U344 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U345 ( .A(n989), .ZN(n706) );
  AOI22_X1 U346 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U347 ( .A(n924), .ZN(n649) );
  AOI22_X1 U348 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U349 ( .A(n922), .ZN(n648) );
  AOI22_X1 U350 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U351 ( .A(n921), .ZN(n647) );
  AOI22_X1 U352 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U353 ( .A(n920), .ZN(n646) );
  AOI22_X1 U354 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U355 ( .A(n919), .ZN(n645) );
  AOI22_X1 U356 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U357 ( .A(n918), .ZN(n644) );
  AOI22_X1 U358 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U359 ( .A(n917), .ZN(n643) );
  AOI22_X1 U360 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U361 ( .A(n916), .ZN(n642) );
  AOI22_X1 U362 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U363 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U364 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U365 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U366 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U367 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U368 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U369 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U370 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U371 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U372 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U373 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U374 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U375 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U376 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U377 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U378 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U379 ( .A(n961), .ZN(n681) );
  AOI22_X1 U380 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U381 ( .A(n959), .ZN(n680) );
  AOI22_X1 U382 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U383 ( .A(n958), .ZN(n679) );
  AOI22_X1 U384 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U385 ( .A(n957), .ZN(n678) );
  AOI22_X1 U386 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U387 ( .A(n956), .ZN(n677) );
  AOI22_X1 U388 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U389 ( .A(n955), .ZN(n676) );
  AOI22_X1 U390 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U391 ( .A(n954), .ZN(n675) );
  AOI22_X1 U392 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U393 ( .A(n953), .ZN(n674) );
  AOI22_X1 U394 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U395 ( .A(n888), .ZN(n617) );
  AOI22_X1 U396 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U397 ( .A(n886), .ZN(n616) );
  AOI22_X1 U398 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U399 ( .A(n885), .ZN(n615) );
  AOI22_X1 U400 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U401 ( .A(n884), .ZN(n614) );
  AOI22_X1 U402 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U403 ( .A(n883), .ZN(n613) );
  AOI22_X1 U404 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U405 ( .A(n882), .ZN(n612) );
  AOI22_X1 U406 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U407 ( .A(n881), .ZN(n611) );
  AOI22_X1 U408 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U409 ( .A(n880), .ZN(n610) );
  AOI22_X1 U410 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U411 ( .A(n879), .ZN(n609) );
  AOI22_X1 U412 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U413 ( .A(n877), .ZN(n608) );
  AOI22_X1 U414 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U415 ( .A(n876), .ZN(n607) );
  AOI22_X1 U416 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U417 ( .A(n875), .ZN(n606) );
  AOI22_X1 U418 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U419 ( .A(n874), .ZN(n605) );
  AOI22_X1 U420 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U421 ( .A(n873), .ZN(n604) );
  AOI22_X1 U422 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U423 ( .A(n872), .ZN(n603) );
  AOI22_X1 U424 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U425 ( .A(n871), .ZN(n602) );
  AOI22_X1 U426 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U427 ( .A(n870), .ZN(n601) );
  AOI22_X1 U428 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U429 ( .A(n868), .ZN(n600) );
  AOI22_X1 U430 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U431 ( .A(n867), .ZN(n599) );
  AOI22_X1 U432 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U433 ( .A(n866), .ZN(n598) );
  AOI22_X1 U434 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U435 ( .A(n865), .ZN(n597) );
  AOI22_X1 U436 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U437 ( .A(n864), .ZN(n596) );
  AOI22_X1 U438 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U439 ( .A(n863), .ZN(n595) );
  AOI22_X1 U440 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U441 ( .A(n862), .ZN(n594) );
  AOI22_X1 U442 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U443 ( .A(n861), .ZN(n293) );
  AOI22_X1 U444 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U445 ( .A(n859), .ZN(n292) );
  AOI22_X1 U446 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U447 ( .A(n858), .ZN(n291) );
  AOI22_X1 U448 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U449 ( .A(n857), .ZN(n290) );
  AOI22_X1 U450 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U451 ( .A(n856), .ZN(n289) );
  AOI22_X1 U452 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U453 ( .A(n855), .ZN(n288) );
  AOI22_X1 U454 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U455 ( .A(n854), .ZN(n287) );
  AOI22_X1 U456 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U457 ( .A(n853), .ZN(n286) );
  AOI22_X1 U458 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U459 ( .A(n852), .ZN(n285) );
  AOI22_X1 U460 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U461 ( .A(n850), .ZN(n284) );
  AOI22_X1 U462 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U463 ( .A(n849), .ZN(n283) );
  AOI22_X1 U464 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U465 ( .A(n848), .ZN(n282) );
  AOI22_X1 U466 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U467 ( .A(n847), .ZN(n281) );
  AOI22_X1 U468 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U469 ( .A(n846), .ZN(n280) );
  AOI22_X1 U470 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U471 ( .A(n845), .ZN(n279) );
  AOI22_X1 U472 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U473 ( .A(n844), .ZN(n278) );
  AOI22_X1 U474 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U475 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U476 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U477 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U478 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U479 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U480 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U481 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U482 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U483 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U484 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U485 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U486 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U487 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U488 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U489 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U490 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U491 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U492 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U493 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U494 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U495 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U496 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U497 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U498 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U499 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U500 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U501 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U502 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U503 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U504 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U505 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U506 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U507 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U508 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U509 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U510 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U511 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U512 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U513 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U514 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U515 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U516 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U517 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U518 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U519 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U520 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U521 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U522 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U523 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U524 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U525 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U526 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U527 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U528 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U529 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U530 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U531 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U532 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U533 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U534 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U535 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U536 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U537 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U538 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U539 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U540 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U541 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U542 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U543 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U544 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U545 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U546 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U547 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U548 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U549 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U550 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U551 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U552 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U553 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U554 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U555 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U556 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U557 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U558 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U559 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U560 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U561 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U562 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U563 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U564 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U565 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U566 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U567 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U568 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U569 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U570 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U571 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U572 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U573 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U574 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U575 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U576 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U577 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U578 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U579 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U580 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U581 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U582 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U583 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U584 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U585 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U586 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U587 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U588 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U589 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U590 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U591 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U592 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U593 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U594 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U595 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U596 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U597 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U598 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U599 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U600 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U601 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U602 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U603 ( .A(N13), .ZN(n842) );
  INV_X1 U604 ( .A(N14), .ZN(n843) );
  MUX2_X1 U605 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n247), .Z(n1) );
  MUX2_X1 U606 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n247), .Z(n2) );
  MUX2_X1 U607 ( .A(n2), .B(n1), .S(n242), .Z(n3) );
  MUX2_X1 U608 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n247), .Z(n4) );
  MUX2_X1 U609 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n247), .Z(n5) );
  MUX2_X1 U610 ( .A(n5), .B(n4), .S(n242), .Z(n6) );
  MUX2_X1 U611 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U612 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n247), .Z(n8) );
  MUX2_X1 U613 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n247), .Z(n9) );
  MUX2_X1 U614 ( .A(n9), .B(n8), .S(n242), .Z(n10) );
  MUX2_X1 U615 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n247), .Z(n11) );
  MUX2_X1 U616 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n247), .Z(n12) );
  MUX2_X1 U617 ( .A(n12), .B(n11), .S(n242), .Z(n13) );
  MUX2_X1 U618 ( .A(n13), .B(n10), .S(n241), .Z(n14) );
  MUX2_X1 U619 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U620 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n245), .Z(n16) );
  MUX2_X1 U621 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n245), .Z(n17) );
  MUX2_X1 U622 ( .A(n17), .B(n16), .S(n243), .Z(n18) );
  MUX2_X1 U623 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U624 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n245), .Z(n20) );
  MUX2_X1 U625 ( .A(n20), .B(n19), .S(n243), .Z(n21) );
  MUX2_X1 U626 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U627 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n245), .Z(n23) );
  MUX2_X1 U628 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n245), .Z(n24) );
  MUX2_X1 U629 ( .A(n24), .B(n23), .S(n243), .Z(n25) );
  MUX2_X1 U630 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n245), .Z(n26) );
  MUX2_X1 U631 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n245), .Z(n27) );
  MUX2_X1 U632 ( .A(n27), .B(n26), .S(n243), .Z(n28) );
  MUX2_X1 U633 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U634 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U635 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U636 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n245), .Z(n31) );
  MUX2_X1 U637 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n245), .Z(n32) );
  MUX2_X1 U638 ( .A(n32), .B(n31), .S(n243), .Z(n33) );
  MUX2_X1 U639 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U640 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U641 ( .A(n35), .B(n34), .S(n243), .Z(n36) );
  MUX2_X1 U642 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U643 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n246), .Z(n38) );
  MUX2_X1 U644 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n246), .Z(n39) );
  MUX2_X1 U645 ( .A(n39), .B(n38), .S(n243), .Z(n40) );
  MUX2_X1 U646 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n246), .Z(n41) );
  MUX2_X1 U647 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n246), .Z(n42) );
  MUX2_X1 U648 ( .A(n42), .B(n41), .S(n243), .Z(n43) );
  MUX2_X1 U649 ( .A(n43), .B(n40), .S(N12), .Z(n44) );
  MUX2_X1 U650 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U651 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n246), .Z(n46) );
  MUX2_X1 U652 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n246), .Z(n47) );
  MUX2_X1 U653 ( .A(n47), .B(n46), .S(n243), .Z(n48) );
  MUX2_X1 U654 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n246), .Z(n49) );
  MUX2_X1 U655 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n246), .Z(n50) );
  MUX2_X1 U656 ( .A(n50), .B(n49), .S(n243), .Z(n51) );
  MUX2_X1 U657 ( .A(n51), .B(n48), .S(N12), .Z(n52) );
  MUX2_X1 U658 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n246), .Z(n53) );
  MUX2_X1 U659 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n246), .Z(n54) );
  MUX2_X1 U660 ( .A(n54), .B(n53), .S(n243), .Z(n55) );
  MUX2_X1 U661 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n246), .Z(n56) );
  MUX2_X1 U662 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n246), .Z(n57) );
  MUX2_X1 U663 ( .A(n57), .B(n56), .S(n243), .Z(n58) );
  MUX2_X1 U664 ( .A(n58), .B(n55), .S(N12), .Z(n59) );
  MUX2_X1 U665 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U666 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U667 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n245), .Z(n61) );
  MUX2_X1 U668 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n249), .Z(n62) );
  MUX2_X1 U669 ( .A(n62), .B(n61), .S(n243), .Z(n63) );
  MUX2_X1 U670 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n248), .Z(n64) );
  MUX2_X1 U671 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n249), .Z(n65) );
  MUX2_X1 U672 ( .A(n65), .B(n64), .S(N11), .Z(n66) );
  MUX2_X1 U673 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U674 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n246), .Z(n68) );
  MUX2_X1 U675 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n245), .Z(n69) );
  MUX2_X1 U676 ( .A(n69), .B(n68), .S(N11), .Z(n70) );
  MUX2_X1 U677 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n248), .Z(n71) );
  MUX2_X1 U678 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n249), .Z(n72) );
  MUX2_X1 U679 ( .A(n72), .B(n71), .S(n244), .Z(n73) );
  MUX2_X1 U680 ( .A(n73), .B(n70), .S(n241), .Z(n74) );
  MUX2_X1 U681 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U682 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n248), .Z(n76) );
  MUX2_X1 U683 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n246), .Z(n77) );
  MUX2_X1 U684 ( .A(n77), .B(n76), .S(N11), .Z(n78) );
  MUX2_X1 U685 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n245), .Z(n79) );
  MUX2_X1 U686 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n248), .Z(n80) );
  MUX2_X1 U687 ( .A(n80), .B(n79), .S(n243), .Z(n81) );
  MUX2_X1 U688 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U689 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n250), .Z(n83) );
  MUX2_X1 U690 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n246), .Z(n84) );
  MUX2_X1 U691 ( .A(n84), .B(n83), .S(N11), .Z(n85) );
  MUX2_X1 U692 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n245), .Z(n86) );
  MUX2_X1 U693 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n246), .Z(n87) );
  MUX2_X1 U694 ( .A(n87), .B(n86), .S(n244), .Z(n88) );
  MUX2_X1 U695 ( .A(n88), .B(n85), .S(n241), .Z(n89) );
  MUX2_X1 U696 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U697 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U698 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n249), .Z(n91) );
  MUX2_X1 U699 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n92) );
  MUX2_X1 U700 ( .A(n92), .B(n91), .S(n244), .Z(n93) );
  MUX2_X1 U701 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n248), .Z(n94) );
  MUX2_X1 U702 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n246), .Z(n95) );
  MUX2_X1 U703 ( .A(n95), .B(n94), .S(N11), .Z(n96) );
  MUX2_X1 U704 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U705 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n98) );
  MUX2_X1 U706 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n248), .Z(n99) );
  MUX2_X1 U707 ( .A(n99), .B(n98), .S(N11), .Z(n100) );
  MUX2_X1 U708 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n250), .Z(n101) );
  MUX2_X1 U709 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n249), .Z(n102) );
  MUX2_X1 U710 ( .A(n102), .B(n101), .S(n242), .Z(n103) );
  MUX2_X1 U711 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U712 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U713 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n247), .Z(n106) );
  MUX2_X1 U714 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n247), .Z(n107) );
  MUX2_X1 U715 ( .A(n107), .B(n106), .S(n244), .Z(n108) );
  MUX2_X1 U716 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n247), .Z(n109) );
  MUX2_X1 U717 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n247), .Z(n110) );
  MUX2_X1 U718 ( .A(n110), .B(n109), .S(n242), .Z(n111) );
  MUX2_X1 U719 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U720 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n247), .Z(n113) );
  MUX2_X1 U721 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n247), .Z(n114) );
  MUX2_X1 U722 ( .A(n114), .B(n113), .S(n243), .Z(n115) );
  MUX2_X1 U723 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n247), .Z(n116) );
  MUX2_X1 U724 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n247), .Z(n117) );
  MUX2_X1 U725 ( .A(n117), .B(n116), .S(N11), .Z(n118) );
  MUX2_X1 U726 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U727 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U728 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U729 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n247), .Z(n121) );
  MUX2_X1 U730 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n247), .Z(n122) );
  MUX2_X1 U731 ( .A(n122), .B(n121), .S(n243), .Z(n123) );
  MUX2_X1 U732 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n247), .Z(n124) );
  MUX2_X1 U733 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n247), .Z(n125) );
  MUX2_X1 U734 ( .A(n125), .B(n124), .S(n244), .Z(n126) );
  MUX2_X1 U735 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U736 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n248), .Z(n128) );
  MUX2_X1 U737 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n248), .Z(n129) );
  MUX2_X1 U738 ( .A(n129), .B(n128), .S(n242), .Z(n130) );
  MUX2_X1 U739 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n248), .Z(n131) );
  MUX2_X1 U740 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n248), .Z(n132) );
  MUX2_X1 U741 ( .A(n132), .B(n131), .S(N11), .Z(n133) );
  MUX2_X1 U742 ( .A(n133), .B(n130), .S(n241), .Z(n134) );
  MUX2_X1 U743 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U744 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n248), .Z(n136) );
  MUX2_X1 U745 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n248), .Z(n137) );
  MUX2_X1 U746 ( .A(n137), .B(n136), .S(N11), .Z(n138) );
  MUX2_X1 U747 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n248), .Z(n139) );
  MUX2_X1 U748 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n248), .Z(n140) );
  MUX2_X1 U749 ( .A(n140), .B(n139), .S(N11), .Z(n141) );
  MUX2_X1 U750 ( .A(n141), .B(n138), .S(n241), .Z(n142) );
  MUX2_X1 U751 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n248), .Z(n143) );
  MUX2_X1 U752 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n248), .Z(n144) );
  MUX2_X1 U753 ( .A(n144), .B(n143), .S(N11), .Z(n145) );
  MUX2_X1 U754 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n248), .Z(n146) );
  MUX2_X1 U755 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n248), .Z(n147) );
  MUX2_X1 U756 ( .A(n147), .B(n146), .S(N11), .Z(n148) );
  MUX2_X1 U757 ( .A(n148), .B(n145), .S(n241), .Z(n149) );
  MUX2_X1 U758 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U759 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U760 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n249), .Z(n151) );
  MUX2_X1 U761 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n249), .Z(n152) );
  MUX2_X1 U762 ( .A(n152), .B(n151), .S(n242), .Z(n153) );
  MUX2_X1 U763 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n249), .Z(n154) );
  MUX2_X1 U764 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n249), .Z(n155) );
  MUX2_X1 U765 ( .A(n155), .B(n154), .S(n242), .Z(n156) );
  MUX2_X1 U766 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U767 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n249), .Z(n158) );
  MUX2_X1 U768 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n249), .Z(n159) );
  MUX2_X1 U769 ( .A(n159), .B(n158), .S(n242), .Z(n160) );
  MUX2_X1 U770 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n249), .Z(n161) );
  MUX2_X1 U771 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n249), .Z(n162) );
  MUX2_X1 U772 ( .A(n162), .B(n161), .S(n243), .Z(n163) );
  MUX2_X1 U773 ( .A(n163), .B(n160), .S(N12), .Z(n164) );
  MUX2_X1 U774 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U775 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n249), .Z(n166) );
  MUX2_X1 U776 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n249), .Z(n167) );
  MUX2_X1 U777 ( .A(n167), .B(n166), .S(n242), .Z(n168) );
  MUX2_X1 U778 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n249), .Z(n169) );
  MUX2_X1 U779 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n249), .Z(n170) );
  MUX2_X1 U780 ( .A(n170), .B(n169), .S(n243), .Z(n171) );
  MUX2_X1 U781 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U782 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n250), .Z(n173) );
  MUX2_X1 U783 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n250), .Z(n174) );
  MUX2_X1 U784 ( .A(n174), .B(n173), .S(n244), .Z(n175) );
  MUX2_X1 U785 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n250), .Z(n176) );
  MUX2_X1 U786 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n250), .Z(n177) );
  MUX2_X1 U787 ( .A(n177), .B(n176), .S(n242), .Z(n178) );
  MUX2_X1 U788 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U789 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U790 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U791 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n245), .Z(n181) );
  MUX2_X1 U792 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n250), .Z(n182) );
  MUX2_X1 U793 ( .A(n182), .B(n181), .S(n242), .Z(n183) );
  MUX2_X1 U794 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n250), .Z(n184) );
  MUX2_X1 U795 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n250), .Z(n185) );
  MUX2_X1 U796 ( .A(n185), .B(n184), .S(n242), .Z(n186) );
  MUX2_X1 U797 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U798 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n250), .Z(n188) );
  MUX2_X1 U799 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n250), .Z(n189) );
  MUX2_X1 U800 ( .A(n189), .B(n188), .S(n242), .Z(n190) );
  MUX2_X1 U801 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n246), .Z(n191) );
  MUX2_X1 U802 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n250), .Z(n192) );
  MUX2_X1 U803 ( .A(n192), .B(n191), .S(N11), .Z(n193) );
  MUX2_X1 U804 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U805 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U806 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n250), .Z(n196) );
  MUX2_X1 U807 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(N10), .Z(n197) );
  MUX2_X1 U808 ( .A(n197), .B(n196), .S(n244), .Z(n198) );
  MUX2_X1 U809 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(N10), .Z(n199) );
  MUX2_X1 U810 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n250), .Z(n200) );
  MUX2_X1 U811 ( .A(n200), .B(n199), .S(n244), .Z(n201) );
  MUX2_X1 U812 ( .A(n201), .B(n198), .S(n241), .Z(n202) );
  MUX2_X1 U813 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n203) );
  MUX2_X1 U814 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n250), .Z(n204) );
  MUX2_X1 U815 ( .A(n204), .B(n203), .S(n244), .Z(n205) );
  MUX2_X1 U816 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n206) );
  MUX2_X1 U817 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n250), .Z(n207) );
  MUX2_X1 U818 ( .A(n207), .B(n206), .S(n244), .Z(n208) );
  MUX2_X1 U819 ( .A(n208), .B(n205), .S(N12), .Z(n209) );
  MUX2_X1 U820 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U821 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U822 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n249), .Z(n211) );
  MUX2_X1 U823 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(N10), .Z(n212) );
  MUX2_X1 U824 ( .A(n212), .B(n211), .S(n244), .Z(n213) );
  MUX2_X1 U825 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(N10), .Z(n214) );
  MUX2_X1 U826 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(N10), .Z(n215) );
  MUX2_X1 U827 ( .A(n215), .B(n214), .S(n244), .Z(n216) );
  MUX2_X1 U828 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U829 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n247), .Z(n218) );
  MUX2_X1 U830 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(N10), .Z(n219) );
  MUX2_X1 U831 ( .A(n219), .B(n218), .S(n244), .Z(n220) );
  MUX2_X1 U832 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n250), .Z(n221) );
  MUX2_X1 U833 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n222) );
  MUX2_X1 U834 ( .A(n222), .B(n221), .S(n244), .Z(n223) );
  MUX2_X1 U835 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U836 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U837 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n247), .Z(n226) );
  MUX2_X1 U838 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n250), .Z(n227) );
  MUX2_X1 U839 ( .A(n227), .B(n226), .S(n244), .Z(n228) );
  MUX2_X1 U840 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n247), .Z(n229) );
  MUX2_X1 U841 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n230) );
  MUX2_X1 U842 ( .A(n230), .B(n229), .S(n244), .Z(n231) );
  MUX2_X1 U843 ( .A(n231), .B(n228), .S(n241), .Z(n232) );
  MUX2_X1 U844 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n233) );
  MUX2_X1 U845 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n234) );
  MUX2_X1 U846 ( .A(n234), .B(n233), .S(n244), .Z(n235) );
  MUX2_X1 U847 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n236) );
  MUX2_X1 U848 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n237) );
  MUX2_X1 U849 ( .A(n237), .B(n236), .S(n244), .Z(n238) );
  MUX2_X1 U850 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U851 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U852 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U853 ( .A(N11), .Z(n242) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_21 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(n250), .Z(n249) );
  BUF_X1 U4 ( .A(n250), .Z(n245) );
  BUF_X1 U5 ( .A(n250), .Z(n246) );
  BUF_X1 U6 ( .A(n250), .Z(n247) );
  BUF_X1 U7 ( .A(n250), .Z(n248) );
  BUF_X1 U8 ( .A(N10), .Z(n250) );
  INV_X1 U9 ( .A(n1111), .ZN(n841) );
  INV_X1 U10 ( .A(n1100), .ZN(n840) );
  INV_X1 U11 ( .A(n1090), .ZN(n839) );
  INV_X1 U12 ( .A(n1080), .ZN(n838) );
  INV_X1 U13 ( .A(n1070), .ZN(n837) );
  INV_X1 U14 ( .A(n1060), .ZN(n836) );
  INV_X1 U15 ( .A(n1051), .ZN(n835) );
  INV_X1 U16 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U19 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U20 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U21 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U22 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U23 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U24 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U26 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U27 ( .A(n1131), .ZN(n816) );
  INV_X1 U28 ( .A(n1121), .ZN(n815) );
  INV_X1 U29 ( .A(n887), .ZN(n814) );
  INV_X1 U30 ( .A(n878), .ZN(n813) );
  INV_X1 U31 ( .A(n869), .ZN(n812) );
  INV_X1 U32 ( .A(n860), .ZN(n811) );
  INV_X1 U33 ( .A(n851), .ZN(n810) );
  INV_X1 U34 ( .A(n987), .ZN(n828) );
  INV_X1 U35 ( .A(n978), .ZN(n827) );
  INV_X1 U36 ( .A(n969), .ZN(n826) );
  INV_X1 U37 ( .A(n914), .ZN(n820) );
  INV_X1 U38 ( .A(n905), .ZN(n819) );
  INV_X1 U39 ( .A(n896), .ZN(n818) );
  INV_X1 U40 ( .A(n1033), .ZN(n833) );
  INV_X1 U41 ( .A(n1023), .ZN(n832) );
  INV_X1 U42 ( .A(n1014), .ZN(n831) );
  INV_X1 U43 ( .A(n1005), .ZN(n830) );
  INV_X1 U44 ( .A(n996), .ZN(n829) );
  INV_X1 U45 ( .A(n960), .ZN(n825) );
  INV_X1 U46 ( .A(n950), .ZN(n824) );
  INV_X1 U47 ( .A(n941), .ZN(n823) );
  INV_X1 U48 ( .A(n932), .ZN(n822) );
  INV_X1 U49 ( .A(n923), .ZN(n821) );
  INV_X1 U50 ( .A(n1142), .ZN(n817) );
  BUF_X1 U51 ( .A(N11), .Z(n242) );
  BUF_X1 U52 ( .A(N11), .Z(n243) );
  BUF_X1 U53 ( .A(N11), .Z(n244) );
  INV_X1 U54 ( .A(N10), .ZN(n251) );
  BUF_X1 U55 ( .A(N12), .Z(n241) );
  NOR3_X1 U56 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U57 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U58 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U60 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U62 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U63 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U64 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U65 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U67 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U69 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U70 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U71 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U72 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U73 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U74 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U75 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U76 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U77 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U79 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U81 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U82 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U83 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U84 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U85 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U86 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U88 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U89 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U90 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U92 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U94 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U95 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U96 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U97 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U98 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U99 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U100 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U101 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U102 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U103 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U104 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U105 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U106 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U107 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U108 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U109 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U110 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U111 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U112 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U113 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U114 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U115 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U116 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U117 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U118 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U119 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U120 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U121 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U122 ( .A(n988), .ZN(n705) );
  AOI22_X1 U123 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U124 ( .A(n986), .ZN(n704) );
  AOI22_X1 U125 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U126 ( .A(n985), .ZN(n703) );
  AOI22_X1 U127 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U128 ( .A(n984), .ZN(n702) );
  AOI22_X1 U129 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U130 ( .A(n983), .ZN(n701) );
  AOI22_X1 U131 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U132 ( .A(n982), .ZN(n700) );
  AOI22_X1 U133 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U134 ( .A(n981), .ZN(n699) );
  AOI22_X1 U135 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U136 ( .A(n980), .ZN(n698) );
  AOI22_X1 U137 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U138 ( .A(n951), .ZN(n673) );
  AOI22_X1 U139 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U140 ( .A(n949), .ZN(n672) );
  AOI22_X1 U141 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U142 ( .A(n948), .ZN(n671) );
  AOI22_X1 U143 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U144 ( .A(n947), .ZN(n670) );
  AOI22_X1 U145 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U146 ( .A(n946), .ZN(n669) );
  AOI22_X1 U147 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U148 ( .A(n945), .ZN(n668) );
  AOI22_X1 U149 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U150 ( .A(n944), .ZN(n667) );
  AOI22_X1 U151 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U152 ( .A(n943), .ZN(n666) );
  AOI22_X1 U153 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U154 ( .A(n915), .ZN(n641) );
  AOI22_X1 U155 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U156 ( .A(n913), .ZN(n640) );
  AOI22_X1 U157 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U158 ( .A(n912), .ZN(n639) );
  AOI22_X1 U159 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U160 ( .A(n911), .ZN(n638) );
  AOI22_X1 U161 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U162 ( .A(n910), .ZN(n637) );
  AOI22_X1 U163 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U164 ( .A(n909), .ZN(n636) );
  AOI22_X1 U165 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U166 ( .A(n908), .ZN(n635) );
  AOI22_X1 U167 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U168 ( .A(n907), .ZN(n634) );
  AOI22_X1 U169 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U170 ( .A(n942), .ZN(n665) );
  AOI22_X1 U171 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U172 ( .A(n940), .ZN(n664) );
  AOI22_X1 U173 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U174 ( .A(n939), .ZN(n663) );
  AOI22_X1 U175 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U176 ( .A(n938), .ZN(n662) );
  AOI22_X1 U177 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U178 ( .A(n937), .ZN(n661) );
  AOI22_X1 U179 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U180 ( .A(n936), .ZN(n660) );
  AOI22_X1 U181 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U182 ( .A(n935), .ZN(n659) );
  AOI22_X1 U183 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U184 ( .A(n934), .ZN(n658) );
  AOI22_X1 U185 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U186 ( .A(n933), .ZN(n657) );
  AOI22_X1 U187 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U188 ( .A(n931), .ZN(n656) );
  AOI22_X1 U189 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U190 ( .A(n930), .ZN(n655) );
  AOI22_X1 U191 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U192 ( .A(n929), .ZN(n654) );
  AOI22_X1 U193 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U194 ( .A(n928), .ZN(n653) );
  AOI22_X1 U195 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U196 ( .A(n927), .ZN(n652) );
  AOI22_X1 U197 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U198 ( .A(n926), .ZN(n651) );
  AOI22_X1 U199 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U200 ( .A(n925), .ZN(n650) );
  AOI22_X1 U201 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U202 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U203 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U204 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U205 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U206 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U207 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U208 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U209 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U210 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U211 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U212 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U213 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U214 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U215 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U216 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U217 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U218 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U219 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U220 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U221 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U222 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U223 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U224 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U225 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U226 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U227 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U228 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U229 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U230 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U231 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U232 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U233 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U234 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U236 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U238 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U240 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U242 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U244 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U246 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U248 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U250 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U252 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U254 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U256 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U258 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U260 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U262 ( .A(n999), .ZN(n715) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U264 ( .A(n998), .ZN(n714) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U266 ( .A(n979), .ZN(n697) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U268 ( .A(n977), .ZN(n696) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U270 ( .A(n976), .ZN(n695) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U272 ( .A(n975), .ZN(n694) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U274 ( .A(n974), .ZN(n693) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U276 ( .A(n973), .ZN(n692) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U278 ( .A(n972), .ZN(n691) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U280 ( .A(n971), .ZN(n690) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U282 ( .A(n970), .ZN(n689) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U284 ( .A(n968), .ZN(n688) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U286 ( .A(n967), .ZN(n687) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U288 ( .A(n966), .ZN(n686) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U290 ( .A(n965), .ZN(n685) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U292 ( .A(n964), .ZN(n684) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U294 ( .A(n906), .ZN(n633) );
  AOI22_X1 U295 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U296 ( .A(n904), .ZN(n632) );
  AOI22_X1 U297 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U298 ( .A(n903), .ZN(n631) );
  AOI22_X1 U299 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U300 ( .A(n902), .ZN(n630) );
  AOI22_X1 U301 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U302 ( .A(n901), .ZN(n629) );
  AOI22_X1 U303 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U304 ( .A(n900), .ZN(n628) );
  AOI22_X1 U305 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U306 ( .A(n899), .ZN(n627) );
  AOI22_X1 U307 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U308 ( .A(n898), .ZN(n626) );
  AOI22_X1 U309 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U310 ( .A(n897), .ZN(n625) );
  AOI22_X1 U311 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U312 ( .A(n895), .ZN(n624) );
  AOI22_X1 U313 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U314 ( .A(n894), .ZN(n623) );
  AOI22_X1 U315 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U316 ( .A(n893), .ZN(n622) );
  AOI22_X1 U317 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U318 ( .A(n892), .ZN(n621) );
  AOI22_X1 U319 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U320 ( .A(n891), .ZN(n620) );
  AOI22_X1 U321 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U322 ( .A(n890), .ZN(n619) );
  AOI22_X1 U323 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U324 ( .A(n889), .ZN(n618) );
  AOI22_X1 U325 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U326 ( .A(n963), .ZN(n683) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U328 ( .A(n962), .ZN(n682) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U330 ( .A(N12), .ZN(n253) );
  INV_X1 U331 ( .A(N11), .ZN(n252) );
  INV_X1 U332 ( .A(n997), .ZN(n713) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U334 ( .A(n995), .ZN(n712) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U336 ( .A(n994), .ZN(n711) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U338 ( .A(n993), .ZN(n710) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U340 ( .A(n992), .ZN(n709) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U342 ( .A(n991), .ZN(n708) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U344 ( .A(n990), .ZN(n707) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U346 ( .A(n989), .ZN(n706) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U348 ( .A(n924), .ZN(n649) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U350 ( .A(n922), .ZN(n648) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U352 ( .A(n921), .ZN(n647) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U354 ( .A(n920), .ZN(n646) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U356 ( .A(n919), .ZN(n645) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U358 ( .A(n918), .ZN(n644) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U360 ( .A(n917), .ZN(n643) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U362 ( .A(n916), .ZN(n642) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U364 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U366 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U368 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U370 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U372 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U374 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U376 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U378 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U380 ( .A(n961), .ZN(n681) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U382 ( .A(n959), .ZN(n680) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U384 ( .A(n958), .ZN(n679) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U386 ( .A(n957), .ZN(n678) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U388 ( .A(n956), .ZN(n677) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U390 ( .A(n955), .ZN(n676) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U392 ( .A(n954), .ZN(n675) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U394 ( .A(n953), .ZN(n674) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U396 ( .A(n888), .ZN(n617) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U398 ( .A(n886), .ZN(n616) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U400 ( .A(n885), .ZN(n615) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U402 ( .A(n884), .ZN(n614) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U404 ( .A(n883), .ZN(n613) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U406 ( .A(n882), .ZN(n612) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U408 ( .A(n881), .ZN(n611) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U410 ( .A(n880), .ZN(n610) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U412 ( .A(n879), .ZN(n609) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U414 ( .A(n877), .ZN(n608) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U416 ( .A(n876), .ZN(n607) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U418 ( .A(n875), .ZN(n606) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U420 ( .A(n874), .ZN(n605) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U422 ( .A(n873), .ZN(n604) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U424 ( .A(n872), .ZN(n603) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U426 ( .A(n871), .ZN(n602) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U428 ( .A(n870), .ZN(n601) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U430 ( .A(n868), .ZN(n600) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U432 ( .A(n867), .ZN(n599) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U434 ( .A(n866), .ZN(n598) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U436 ( .A(n865), .ZN(n597) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U438 ( .A(n864), .ZN(n596) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U440 ( .A(n863), .ZN(n595) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U442 ( .A(n862), .ZN(n594) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U444 ( .A(n861), .ZN(n293) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U446 ( .A(n859), .ZN(n292) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U448 ( .A(n858), .ZN(n291) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U450 ( .A(n857), .ZN(n290) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U452 ( .A(n856), .ZN(n289) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U454 ( .A(n855), .ZN(n288) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U456 ( .A(n854), .ZN(n287) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U458 ( .A(n853), .ZN(n286) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U460 ( .A(n852), .ZN(n285) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U462 ( .A(n850), .ZN(n284) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U464 ( .A(n849), .ZN(n283) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U466 ( .A(n848), .ZN(n282) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U468 ( .A(n847), .ZN(n281) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U470 ( .A(n846), .ZN(n280) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U472 ( .A(n845), .ZN(n279) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U474 ( .A(n844), .ZN(n278) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U476 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U477 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U478 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U479 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U480 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U481 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U482 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U483 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U484 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U485 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U486 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U487 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U488 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U489 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U490 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U491 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U492 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U494 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U496 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U498 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U500 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U502 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U504 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U506 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U508 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U510 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U512 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U514 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U516 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U518 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U520 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U522 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U524 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U526 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U528 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U530 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U532 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U534 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U536 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U538 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U540 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U542 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U544 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U546 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U548 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U550 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U552 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U554 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U556 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U558 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U560 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U562 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U564 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U566 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U568 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U570 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U572 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U574 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U576 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U578 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U580 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U582 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U584 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U586 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U588 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U590 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U592 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U594 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U596 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U598 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U600 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U602 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U604 ( .A(N13), .ZN(n842) );
  INV_X1 U605 ( .A(N14), .ZN(n843) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n249), .Z(n1) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n245), .Z(n2) );
  MUX2_X1 U608 ( .A(n2), .B(n1), .S(n242), .Z(n3) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n249), .Z(n4) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n249), .Z(n5) );
  MUX2_X1 U611 ( .A(n5), .B(n4), .S(n244), .Z(n6) );
  MUX2_X1 U612 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n250), .Z(n8) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n248), .Z(n9) );
  MUX2_X1 U615 ( .A(n9), .B(n8), .S(n243), .Z(n10) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n247), .Z(n11) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n247), .Z(n12) );
  MUX2_X1 U618 ( .A(n12), .B(n11), .S(n243), .Z(n13) );
  MUX2_X1 U619 ( .A(n13), .B(n10), .S(n241), .Z(n14) );
  MUX2_X1 U620 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n245), .Z(n16) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n245), .Z(n17) );
  MUX2_X1 U623 ( .A(n17), .B(n16), .S(n242), .Z(n18) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n245), .Z(n20) );
  MUX2_X1 U626 ( .A(n20), .B(n19), .S(n242), .Z(n21) );
  MUX2_X1 U627 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n245), .Z(n23) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n245), .Z(n24) );
  MUX2_X1 U630 ( .A(n24), .B(n23), .S(n242), .Z(n25) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n245), .Z(n26) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n245), .Z(n27) );
  MUX2_X1 U633 ( .A(n27), .B(n26), .S(n242), .Z(n28) );
  MUX2_X1 U634 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U635 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U636 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n245), .Z(n31) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n245), .Z(n32) );
  MUX2_X1 U639 ( .A(n32), .B(n31), .S(n242), .Z(n33) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U642 ( .A(n35), .B(n34), .S(n242), .Z(n36) );
  MUX2_X1 U643 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n246), .Z(n38) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n246), .Z(n39) );
  MUX2_X1 U646 ( .A(n39), .B(n38), .S(n242), .Z(n40) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n246), .Z(n41) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n246), .Z(n42) );
  MUX2_X1 U649 ( .A(n42), .B(n41), .S(n242), .Z(n43) );
  MUX2_X1 U650 ( .A(n43), .B(n40), .S(N12), .Z(n44) );
  MUX2_X1 U651 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n246), .Z(n46) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n246), .Z(n47) );
  MUX2_X1 U654 ( .A(n47), .B(n46), .S(n242), .Z(n48) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n246), .Z(n49) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n246), .Z(n50) );
  MUX2_X1 U657 ( .A(n50), .B(n49), .S(n242), .Z(n51) );
  MUX2_X1 U658 ( .A(n51), .B(n48), .S(N12), .Z(n52) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n246), .Z(n53) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n246), .Z(n54) );
  MUX2_X1 U661 ( .A(n54), .B(n53), .S(n242), .Z(n55) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n246), .Z(n56) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n246), .Z(n57) );
  MUX2_X1 U664 ( .A(n57), .B(n56), .S(n242), .Z(n58) );
  MUX2_X1 U665 ( .A(n58), .B(n55), .S(N12), .Z(n59) );
  MUX2_X1 U666 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U667 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n247), .Z(n61) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n247), .Z(n62) );
  MUX2_X1 U670 ( .A(n62), .B(n61), .S(n243), .Z(n63) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n247), .Z(n64) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n247), .Z(n65) );
  MUX2_X1 U673 ( .A(n65), .B(n64), .S(n243), .Z(n66) );
  MUX2_X1 U674 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n247), .Z(n68) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n247), .Z(n69) );
  MUX2_X1 U677 ( .A(n69), .B(n68), .S(n243), .Z(n70) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n247), .Z(n71) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n247), .Z(n72) );
  MUX2_X1 U680 ( .A(n72), .B(n71), .S(n243), .Z(n73) );
  MUX2_X1 U681 ( .A(n73), .B(n70), .S(n241), .Z(n74) );
  MUX2_X1 U682 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n247), .Z(n76) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n247), .Z(n77) );
  MUX2_X1 U685 ( .A(n77), .B(n76), .S(n243), .Z(n78) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n247), .Z(n79) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n247), .Z(n80) );
  MUX2_X1 U688 ( .A(n80), .B(n79), .S(n243), .Z(n81) );
  MUX2_X1 U689 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n248), .Z(n83) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n248), .Z(n84) );
  MUX2_X1 U692 ( .A(n84), .B(n83), .S(n243), .Z(n85) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n248), .Z(n86) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n248), .Z(n87) );
  MUX2_X1 U695 ( .A(n87), .B(n86), .S(n243), .Z(n88) );
  MUX2_X1 U696 ( .A(n88), .B(n85), .S(n241), .Z(n89) );
  MUX2_X1 U697 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U698 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n248), .Z(n91) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n248), .Z(n92) );
  MUX2_X1 U701 ( .A(n92), .B(n91), .S(n243), .Z(n93) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n248), .Z(n94) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n248), .Z(n95) );
  MUX2_X1 U704 ( .A(n95), .B(n94), .S(n243), .Z(n96) );
  MUX2_X1 U705 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n248), .Z(n98) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n248), .Z(n99) );
  MUX2_X1 U708 ( .A(n99), .B(n98), .S(n243), .Z(n100) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n248), .Z(n101) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n248), .Z(n102) );
  MUX2_X1 U711 ( .A(n102), .B(n101), .S(n243), .Z(n103) );
  MUX2_X1 U712 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U713 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n250), .Z(n106) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(N10), .Z(n107) );
  MUX2_X1 U716 ( .A(n107), .B(n106), .S(n244), .Z(n108) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(N10), .Z(n109) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n246), .Z(n110) );
  MUX2_X1 U719 ( .A(n110), .B(n109), .S(n244), .Z(n111) );
  MUX2_X1 U720 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(N10), .Z(n113) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n250), .Z(n114) );
  MUX2_X1 U723 ( .A(n114), .B(n113), .S(n244), .Z(n115) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n116) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n246), .Z(n117) );
  MUX2_X1 U726 ( .A(n117), .B(n116), .S(n244), .Z(n118) );
  MUX2_X1 U727 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U728 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U729 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n246), .Z(n121) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(N10), .Z(n122) );
  MUX2_X1 U732 ( .A(n122), .B(n121), .S(n244), .Z(n123) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(N10), .Z(n124) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n125) );
  MUX2_X1 U735 ( .A(n125), .B(n124), .S(n244), .Z(n126) );
  MUX2_X1 U736 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n249), .Z(n128) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(N10), .Z(n129) );
  MUX2_X1 U739 ( .A(n129), .B(n128), .S(n244), .Z(n130) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n250), .Z(n131) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(N10), .Z(n132) );
  MUX2_X1 U742 ( .A(n132), .B(n131), .S(n244), .Z(n133) );
  MUX2_X1 U743 ( .A(n133), .B(n130), .S(n241), .Z(n134) );
  MUX2_X1 U744 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n249), .Z(n136) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n250), .Z(n137) );
  MUX2_X1 U747 ( .A(n137), .B(n136), .S(n244), .Z(n138) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n246), .Z(n139) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(N10), .Z(n140) );
  MUX2_X1 U750 ( .A(n140), .B(n139), .S(n244), .Z(n141) );
  MUX2_X1 U751 ( .A(n141), .B(n138), .S(n241), .Z(n142) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(N10), .Z(n143) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(N10), .Z(n144) );
  MUX2_X1 U754 ( .A(n144), .B(n143), .S(n244), .Z(n145) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(N10), .Z(n146) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n147) );
  MUX2_X1 U757 ( .A(n147), .B(n146), .S(n244), .Z(n148) );
  MUX2_X1 U758 ( .A(n148), .B(n145), .S(n241), .Z(n149) );
  MUX2_X1 U759 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U760 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n249), .Z(n151) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n249), .Z(n152) );
  MUX2_X1 U763 ( .A(n152), .B(n151), .S(n242), .Z(n153) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n249), .Z(n154) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n249), .Z(n155) );
  MUX2_X1 U766 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U767 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n249), .Z(n158) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n249), .Z(n159) );
  MUX2_X1 U770 ( .A(n159), .B(n158), .S(N11), .Z(n160) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n249), .Z(n161) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n249), .Z(n162) );
  MUX2_X1 U773 ( .A(n162), .B(n161), .S(N11), .Z(n163) );
  MUX2_X1 U774 ( .A(n163), .B(n160), .S(N12), .Z(n164) );
  MUX2_X1 U775 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n249), .Z(n166) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n249), .Z(n167) );
  MUX2_X1 U778 ( .A(n167), .B(n166), .S(n244), .Z(n168) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n249), .Z(n169) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n249), .Z(n170) );
  MUX2_X1 U781 ( .A(n170), .B(n169), .S(N11), .Z(n171) );
  MUX2_X1 U782 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n250), .Z(n173) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n245), .Z(n174) );
  MUX2_X1 U785 ( .A(n174), .B(n173), .S(N11), .Z(n175) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n250), .Z(n176) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n245), .Z(n177) );
  MUX2_X1 U788 ( .A(n177), .B(n176), .S(n244), .Z(n178) );
  MUX2_X1 U789 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U790 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U791 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n245), .Z(n181) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n248), .Z(n182) );
  MUX2_X1 U794 ( .A(n182), .B(n181), .S(n243), .Z(n183) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n249), .Z(n184) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n250), .Z(n185) );
  MUX2_X1 U797 ( .A(n185), .B(n184), .S(N11), .Z(n186) );
  MUX2_X1 U798 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n250), .Z(n188) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n250), .Z(n189) );
  MUX2_X1 U801 ( .A(n189), .B(n188), .S(N11), .Z(n190) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n247), .Z(n191) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n250), .Z(n192) );
  MUX2_X1 U804 ( .A(n192), .B(n191), .S(n242), .Z(n193) );
  MUX2_X1 U805 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U806 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n248), .Z(n196) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n250), .Z(n197) );
  MUX2_X1 U809 ( .A(n197), .B(n196), .S(n243), .Z(n198) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n246), .Z(n199) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n247), .Z(n200) );
  MUX2_X1 U812 ( .A(n200), .B(n199), .S(N11), .Z(n201) );
  MUX2_X1 U813 ( .A(n201), .B(n198), .S(n241), .Z(n202) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n248), .Z(n203) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n250), .Z(n204) );
  MUX2_X1 U816 ( .A(n204), .B(n203), .S(n243), .Z(n205) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n250), .Z(n206) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n247), .Z(n207) );
  MUX2_X1 U819 ( .A(n207), .B(n206), .S(N11), .Z(n208) );
  MUX2_X1 U820 ( .A(n208), .B(n205), .S(N12), .Z(n209) );
  MUX2_X1 U821 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U822 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n247), .Z(n211) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n247), .Z(n212) );
  MUX2_X1 U825 ( .A(n212), .B(n211), .S(n242), .Z(n213) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n245), .Z(n214) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n248), .Z(n215) );
  MUX2_X1 U828 ( .A(n215), .B(n214), .S(n242), .Z(n216) );
  MUX2_X1 U829 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n250), .Z(n218) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n248), .Z(n219) );
  MUX2_X1 U832 ( .A(n219), .B(n218), .S(N11), .Z(n220) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n250), .Z(n221) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n248), .Z(n222) );
  MUX2_X1 U835 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U836 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U837 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(N10), .Z(n226) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n246), .Z(n227) );
  MUX2_X1 U840 ( .A(n227), .B(n226), .S(n244), .Z(n228) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n250), .Z(n229) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n246), .Z(n230) );
  MUX2_X1 U843 ( .A(n230), .B(n229), .S(N11), .Z(n231) );
  MUX2_X1 U844 ( .A(n231), .B(n228), .S(n241), .Z(n232) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n245), .Z(n233) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n250), .Z(n234) );
  MUX2_X1 U847 ( .A(n234), .B(n233), .S(n244), .Z(n235) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n250), .Z(n236) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n250), .Z(n237) );
  MUX2_X1 U850 ( .A(n237), .B(n236), .S(N11), .Z(n238) );
  MUX2_X1 U851 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U852 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U853 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_20 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n256), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n257), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n258), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n259), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n260), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n261), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n262), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n263), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n264), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n265), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n266), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n267), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n268), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n269), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n270), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n271), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n272), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n273), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n274), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n275), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n276), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n277), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n278), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n279), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n280), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n281), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n282), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n283), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n284), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n285), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n286), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n287), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n288), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n289), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n290), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n291), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n292), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n293), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n594), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n595), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n596), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n597), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n598), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n599), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n600), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n601), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n602), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n603), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n604), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n605), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n606), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n607), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n608), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n609), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n610), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n611), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n612), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n613), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n614), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n615), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n616), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n617), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n618), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n619), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n620), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n621), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n622), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n623), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n624), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n625), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n626), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n627), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n628), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n629), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n630), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n631), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n632), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n633), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n634), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n635), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n636), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n637), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n638), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n639), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n640), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n641), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n642), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n643), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n644), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n645), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n646), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n647), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n648), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n649), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n650), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n651), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n652), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n653), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n654), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n655), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n656), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n657), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n658), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n659), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n660), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n661), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n662), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n663), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n664), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n665), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n666), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n667), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n668), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n669), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n670), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n671), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n672), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n673), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n674), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n675), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n676), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n677), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n678), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n679), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n680), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n681), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n682), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n683), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n684), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n685), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n686), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n687), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n688), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n689), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n690), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n691), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n692), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n693), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n694), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n695), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n696), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n697), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n698), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n699), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n700), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n701), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n702), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n703), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n704), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n705), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n706), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n707), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n708), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n709), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n710), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n711), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n712), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n713), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n714), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n715), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n716), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n717), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n718), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n719), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n720), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n721), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n722), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n723), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n724), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n725), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n726), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n727), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n728), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n729), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n730), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n731), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n732), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n733), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n734), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n735), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n736), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n737), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n738), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n739), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n740), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n741), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n742), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n743), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n744), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n745), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n746), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n747), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n748), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n749), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n750), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n751), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n752), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n753), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n754), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n755), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n756), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n757), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n758), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n759), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n760), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n761), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n762), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n763), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n764), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n765), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n766), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n767), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n768), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n769), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n770), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n771), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n772), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n773), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n774), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n775), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n776), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n777), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n778), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n779), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n780), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n781), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n782), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n783), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n784), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n785), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n786), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n787), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n788), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n789), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n790), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n791), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n792), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n793), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n794), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n795), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n796), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n797), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n798), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n799), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n800), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n801), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n802), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n803), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n804), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n805), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n806), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n807), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n808), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n809), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n810), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n811), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(n252), .Z(n249) );
  BUF_X1 U5 ( .A(N10), .Z(n250) );
  BUF_X1 U6 ( .A(n252), .Z(n251) );
  BUF_X1 U7 ( .A(n252), .Z(n248) );
  BUF_X1 U8 ( .A(n252), .Z(n247) );
  BUF_X1 U9 ( .A(N10), .Z(n252) );
  INV_X1 U10 ( .A(n1113), .ZN(n843) );
  INV_X1 U11 ( .A(n1102), .ZN(n842) );
  INV_X1 U12 ( .A(n1092), .ZN(n841) );
  INV_X1 U13 ( .A(n1082), .ZN(n840) );
  INV_X1 U14 ( .A(n1072), .ZN(n839) );
  INV_X1 U15 ( .A(n1062), .ZN(n838) );
  INV_X1 U16 ( .A(n1053), .ZN(n837) );
  INV_X1 U17 ( .A(n1044), .ZN(n836) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1105) );
  NOR3_X1 U19 ( .A1(N11), .A2(N12), .A3(n253), .ZN(n1094) );
  NAND2_X1 U20 ( .A1(n1104), .A2(n1136), .ZN(n1062) );
  NAND2_X1 U21 ( .A1(n1105), .A2(n1104), .ZN(n1113) );
  NAND2_X1 U22 ( .A1(n1094), .A2(n1104), .ZN(n1102) );
  NAND2_X1 U23 ( .A1(n1084), .A2(n1104), .ZN(n1092) );
  NAND2_X1 U24 ( .A1(n1074), .A2(n1104), .ZN(n1082) );
  NAND2_X1 U25 ( .A1(n1064), .A2(n1104), .ZN(n1072) );
  NAND2_X1 U26 ( .A1(n1104), .A2(n1125), .ZN(n1053) );
  NAND2_X1 U27 ( .A1(n1104), .A2(n1115), .ZN(n1044) );
  INV_X1 U28 ( .A(n1133), .ZN(n818) );
  INV_X1 U29 ( .A(n1123), .ZN(n817) );
  INV_X1 U30 ( .A(n889), .ZN(n816) );
  INV_X1 U31 ( .A(n880), .ZN(n815) );
  INV_X1 U32 ( .A(n871), .ZN(n814) );
  INV_X1 U33 ( .A(n862), .ZN(n813) );
  INV_X1 U34 ( .A(n853), .ZN(n812) );
  INV_X1 U35 ( .A(n989), .ZN(n830) );
  INV_X1 U36 ( .A(n980), .ZN(n829) );
  INV_X1 U37 ( .A(n971), .ZN(n828) );
  INV_X1 U38 ( .A(n916), .ZN(n822) );
  INV_X1 U39 ( .A(n907), .ZN(n821) );
  INV_X1 U40 ( .A(n898), .ZN(n820) );
  INV_X1 U41 ( .A(n1035), .ZN(n835) );
  INV_X1 U42 ( .A(n1025), .ZN(n834) );
  INV_X1 U43 ( .A(n1016), .ZN(n833) );
  INV_X1 U44 ( .A(n1007), .ZN(n832) );
  INV_X1 U45 ( .A(n998), .ZN(n831) );
  INV_X1 U46 ( .A(n962), .ZN(n827) );
  INV_X1 U47 ( .A(n952), .ZN(n826) );
  INV_X1 U48 ( .A(n943), .ZN(n825) );
  INV_X1 U49 ( .A(n934), .ZN(n824) );
  INV_X1 U50 ( .A(n925), .ZN(n823) );
  INV_X1 U51 ( .A(n1144), .ZN(n819) );
  BUF_X1 U52 ( .A(N11), .Z(n244) );
  BUF_X1 U53 ( .A(N11), .Z(n245) );
  BUF_X1 U54 ( .A(N11), .Z(n246) );
  INV_X1 U55 ( .A(N10), .ZN(n253) );
  BUF_X1 U56 ( .A(N12), .Z(n243) );
  NOR3_X1 U57 ( .A1(n255), .A2(N10), .A3(n254), .ZN(n1125) );
  NOR3_X1 U58 ( .A1(n255), .A2(n253), .A3(n254), .ZN(n1115) );
  NOR3_X1 U59 ( .A1(n253), .A2(N11), .A3(n255), .ZN(n1136) );
  NOR3_X1 U60 ( .A1(N10), .A2(N12), .A3(n254), .ZN(n1084) );
  NOR3_X1 U61 ( .A1(n253), .A2(N12), .A3(n254), .ZN(n1074) );
  NOR3_X1 U62 ( .A1(N10), .A2(N11), .A3(n255), .ZN(n1064) );
  NAND2_X1 U63 ( .A1(n1027), .A2(n1136), .ZN(n989) );
  NAND2_X1 U64 ( .A1(n954), .A2(n1136), .ZN(n916) );
  NAND2_X1 U65 ( .A1(n1027), .A2(n1064), .ZN(n998) );
  NAND2_X1 U66 ( .A1(n954), .A2(n1064), .ZN(n925) );
  NAND2_X1 U67 ( .A1(n1027), .A2(n1105), .ZN(n1035) );
  NAND2_X1 U68 ( .A1(n1027), .A2(n1094), .ZN(n1025) );
  NAND2_X1 U69 ( .A1(n954), .A2(n1105), .ZN(n962) );
  NAND2_X1 U70 ( .A1(n954), .A2(n1094), .ZN(n952) );
  NAND2_X1 U71 ( .A1(n1105), .A2(n1135), .ZN(n889) );
  NAND2_X1 U72 ( .A1(n1094), .A2(n1135), .ZN(n880) );
  NAND2_X1 U73 ( .A1(n1084), .A2(n1135), .ZN(n871) );
  NAND2_X1 U74 ( .A1(n1074), .A2(n1135), .ZN(n862) );
  NAND2_X1 U75 ( .A1(n1064), .A2(n1135), .ZN(n853) );
  NAND2_X1 U76 ( .A1(n1136), .A2(n1135), .ZN(n1144) );
  NAND2_X1 U77 ( .A1(n1125), .A2(n1135), .ZN(n1133) );
  NAND2_X1 U78 ( .A1(n1115), .A2(n1135), .ZN(n1123) );
  NAND2_X1 U79 ( .A1(n1027), .A2(n1084), .ZN(n1016) );
  NAND2_X1 U80 ( .A1(n1027), .A2(n1074), .ZN(n1007) );
  NAND2_X1 U81 ( .A1(n954), .A2(n1084), .ZN(n943) );
  NAND2_X1 U82 ( .A1(n954), .A2(n1074), .ZN(n934) );
  NAND2_X1 U83 ( .A1(n1027), .A2(n1125), .ZN(n980) );
  NAND2_X1 U84 ( .A1(n954), .A2(n1125), .ZN(n907) );
  NAND2_X1 U85 ( .A1(n1027), .A2(n1115), .ZN(n971) );
  NAND2_X1 U86 ( .A1(n954), .A2(n1115), .ZN(n898) );
  AND3_X1 U87 ( .A1(n844), .A2(n845), .A3(wr_en), .ZN(n1104) );
  AND3_X1 U88 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1135) );
  AND3_X1 U89 ( .A1(N13), .A2(n845), .A3(wr_en), .ZN(n1027) );
  AND3_X1 U90 ( .A1(N14), .A2(n844), .A3(wr_en), .ZN(n954) );
  INV_X1 U91 ( .A(n1063), .ZN(n771) );
  AOI22_X1 U92 ( .A1(data_in[0]), .A2(n838), .B1(n1062), .B2(\mem[5][0] ), 
        .ZN(n1063) );
  INV_X1 U93 ( .A(n1061), .ZN(n770) );
  AOI22_X1 U94 ( .A1(data_in[1]), .A2(n838), .B1(n1062), .B2(\mem[5][1] ), 
        .ZN(n1061) );
  INV_X1 U95 ( .A(n1060), .ZN(n769) );
  AOI22_X1 U96 ( .A1(data_in[2]), .A2(n838), .B1(n1062), .B2(\mem[5][2] ), 
        .ZN(n1060) );
  INV_X1 U97 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U98 ( .A1(data_in[3]), .A2(n838), .B1(n1062), .B2(\mem[5][3] ), 
        .ZN(n1059) );
  INV_X1 U99 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U100 ( .A1(data_in[4]), .A2(n838), .B1(n1062), .B2(\mem[5][4] ), 
        .ZN(n1058) );
  INV_X1 U101 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U102 ( .A1(data_in[5]), .A2(n838), .B1(n1062), .B2(\mem[5][5] ), 
        .ZN(n1057) );
  INV_X1 U103 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U104 ( .A1(data_in[6]), .A2(n838), .B1(n1062), .B2(\mem[5][6] ), 
        .ZN(n1056) );
  INV_X1 U105 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U106 ( .A1(data_in[7]), .A2(n838), .B1(n1062), .B2(\mem[5][7] ), 
        .ZN(n1055) );
  INV_X1 U107 ( .A(n1026), .ZN(n739) );
  AOI22_X1 U108 ( .A1(data_in[0]), .A2(n834), .B1(n1025), .B2(\mem[9][0] ), 
        .ZN(n1026) );
  INV_X1 U109 ( .A(n1024), .ZN(n738) );
  AOI22_X1 U110 ( .A1(data_in[1]), .A2(n834), .B1(n1025), .B2(\mem[9][1] ), 
        .ZN(n1024) );
  INV_X1 U111 ( .A(n1023), .ZN(n737) );
  AOI22_X1 U112 ( .A1(data_in[2]), .A2(n834), .B1(n1025), .B2(\mem[9][2] ), 
        .ZN(n1023) );
  INV_X1 U113 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U114 ( .A1(data_in[3]), .A2(n834), .B1(n1025), .B2(\mem[9][3] ), 
        .ZN(n1022) );
  INV_X1 U115 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U116 ( .A1(data_in[4]), .A2(n834), .B1(n1025), .B2(\mem[9][4] ), 
        .ZN(n1021) );
  INV_X1 U117 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U118 ( .A1(data_in[5]), .A2(n834), .B1(n1025), .B2(\mem[9][5] ), 
        .ZN(n1020) );
  INV_X1 U119 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U120 ( .A1(data_in[6]), .A2(n834), .B1(n1025), .B2(\mem[9][6] ), 
        .ZN(n1019) );
  INV_X1 U121 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U122 ( .A1(data_in[7]), .A2(n834), .B1(n1025), .B2(\mem[9][7] ), 
        .ZN(n1018) );
  INV_X1 U123 ( .A(n990), .ZN(n707) );
  AOI22_X1 U124 ( .A1(data_in[0]), .A2(n830), .B1(n989), .B2(\mem[13][0] ), 
        .ZN(n990) );
  INV_X1 U125 ( .A(n988), .ZN(n706) );
  AOI22_X1 U126 ( .A1(data_in[1]), .A2(n830), .B1(n989), .B2(\mem[13][1] ), 
        .ZN(n988) );
  INV_X1 U127 ( .A(n987), .ZN(n705) );
  AOI22_X1 U128 ( .A1(data_in[2]), .A2(n830), .B1(n989), .B2(\mem[13][2] ), 
        .ZN(n987) );
  INV_X1 U129 ( .A(n986), .ZN(n704) );
  AOI22_X1 U130 ( .A1(data_in[3]), .A2(n830), .B1(n989), .B2(\mem[13][3] ), 
        .ZN(n986) );
  INV_X1 U131 ( .A(n985), .ZN(n703) );
  AOI22_X1 U132 ( .A1(data_in[4]), .A2(n830), .B1(n989), .B2(\mem[13][4] ), 
        .ZN(n985) );
  INV_X1 U133 ( .A(n984), .ZN(n702) );
  AOI22_X1 U134 ( .A1(data_in[5]), .A2(n830), .B1(n989), .B2(\mem[13][5] ), 
        .ZN(n984) );
  INV_X1 U135 ( .A(n983), .ZN(n701) );
  AOI22_X1 U136 ( .A1(data_in[6]), .A2(n830), .B1(n989), .B2(\mem[13][6] ), 
        .ZN(n983) );
  INV_X1 U137 ( .A(n982), .ZN(n700) );
  AOI22_X1 U138 ( .A1(data_in[7]), .A2(n830), .B1(n989), .B2(\mem[13][7] ), 
        .ZN(n982) );
  INV_X1 U139 ( .A(n950), .ZN(n673) );
  AOI22_X1 U140 ( .A1(data_in[2]), .A2(n826), .B1(n952), .B2(\mem[17][2] ), 
        .ZN(n950) );
  INV_X1 U141 ( .A(n949), .ZN(n672) );
  AOI22_X1 U142 ( .A1(data_in[3]), .A2(n826), .B1(n952), .B2(\mem[17][3] ), 
        .ZN(n949) );
  INV_X1 U143 ( .A(n948), .ZN(n671) );
  AOI22_X1 U144 ( .A1(data_in[4]), .A2(n826), .B1(n952), .B2(\mem[17][4] ), 
        .ZN(n948) );
  INV_X1 U145 ( .A(n947), .ZN(n670) );
  AOI22_X1 U146 ( .A1(data_in[5]), .A2(n826), .B1(n952), .B2(\mem[17][5] ), 
        .ZN(n947) );
  INV_X1 U147 ( .A(n946), .ZN(n669) );
  AOI22_X1 U148 ( .A1(data_in[6]), .A2(n826), .B1(n952), .B2(\mem[17][6] ), 
        .ZN(n946) );
  INV_X1 U149 ( .A(n945), .ZN(n668) );
  AOI22_X1 U150 ( .A1(data_in[7]), .A2(n826), .B1(n952), .B2(\mem[17][7] ), 
        .ZN(n945) );
  INV_X1 U151 ( .A(n917), .ZN(n643) );
  AOI22_X1 U152 ( .A1(data_in[0]), .A2(n822), .B1(n916), .B2(\mem[21][0] ), 
        .ZN(n917) );
  INV_X1 U153 ( .A(n915), .ZN(n642) );
  AOI22_X1 U154 ( .A1(data_in[1]), .A2(n822), .B1(n916), .B2(\mem[21][1] ), 
        .ZN(n915) );
  INV_X1 U155 ( .A(n914), .ZN(n641) );
  AOI22_X1 U156 ( .A1(data_in[2]), .A2(n822), .B1(n916), .B2(\mem[21][2] ), 
        .ZN(n914) );
  INV_X1 U157 ( .A(n913), .ZN(n640) );
  AOI22_X1 U158 ( .A1(data_in[3]), .A2(n822), .B1(n916), .B2(\mem[21][3] ), 
        .ZN(n913) );
  INV_X1 U159 ( .A(n912), .ZN(n639) );
  AOI22_X1 U160 ( .A1(data_in[4]), .A2(n822), .B1(n916), .B2(\mem[21][4] ), 
        .ZN(n912) );
  INV_X1 U161 ( .A(n911), .ZN(n638) );
  AOI22_X1 U162 ( .A1(data_in[5]), .A2(n822), .B1(n916), .B2(\mem[21][5] ), 
        .ZN(n911) );
  INV_X1 U163 ( .A(n910), .ZN(n637) );
  AOI22_X1 U164 ( .A1(data_in[6]), .A2(n822), .B1(n916), .B2(\mem[21][6] ), 
        .ZN(n910) );
  INV_X1 U165 ( .A(n909), .ZN(n636) );
  AOI22_X1 U166 ( .A1(data_in[7]), .A2(n822), .B1(n916), .B2(\mem[21][7] ), 
        .ZN(n909) );
  INV_X1 U167 ( .A(n966), .ZN(n686) );
  AOI22_X1 U168 ( .A1(data_in[5]), .A2(n828), .B1(n971), .B2(\mem[15][5] ), 
        .ZN(n966) );
  INV_X1 U169 ( .A(n965), .ZN(n685) );
  AOI22_X1 U170 ( .A1(data_in[6]), .A2(n828), .B1(n971), .B2(\mem[15][6] ), 
        .ZN(n965) );
  INV_X1 U171 ( .A(n964), .ZN(n684) );
  AOI22_X1 U172 ( .A1(data_in[7]), .A2(n828), .B1(n971), .B2(\mem[15][7] ), 
        .ZN(n964) );
  INV_X1 U173 ( .A(n944), .ZN(n667) );
  AOI22_X1 U174 ( .A1(data_in[0]), .A2(n825), .B1(n943), .B2(\mem[18][0] ), 
        .ZN(n944) );
  INV_X1 U175 ( .A(n942), .ZN(n666) );
  AOI22_X1 U176 ( .A1(data_in[1]), .A2(n825), .B1(n943), .B2(\mem[18][1] ), 
        .ZN(n942) );
  INV_X1 U177 ( .A(n941), .ZN(n665) );
  AOI22_X1 U178 ( .A1(data_in[2]), .A2(n825), .B1(n943), .B2(\mem[18][2] ), 
        .ZN(n941) );
  INV_X1 U179 ( .A(n940), .ZN(n664) );
  AOI22_X1 U180 ( .A1(data_in[3]), .A2(n825), .B1(n943), .B2(\mem[18][3] ), 
        .ZN(n940) );
  INV_X1 U181 ( .A(n939), .ZN(n663) );
  AOI22_X1 U182 ( .A1(data_in[4]), .A2(n825), .B1(n943), .B2(\mem[18][4] ), 
        .ZN(n939) );
  INV_X1 U183 ( .A(n938), .ZN(n662) );
  AOI22_X1 U184 ( .A1(data_in[5]), .A2(n825), .B1(n943), .B2(\mem[18][5] ), 
        .ZN(n938) );
  INV_X1 U185 ( .A(n937), .ZN(n661) );
  AOI22_X1 U186 ( .A1(data_in[6]), .A2(n825), .B1(n943), .B2(\mem[18][6] ), 
        .ZN(n937) );
  INV_X1 U187 ( .A(n936), .ZN(n660) );
  AOI22_X1 U188 ( .A1(data_in[7]), .A2(n825), .B1(n943), .B2(\mem[18][7] ), 
        .ZN(n936) );
  INV_X1 U189 ( .A(n935), .ZN(n659) );
  AOI22_X1 U190 ( .A1(data_in[0]), .A2(n824), .B1(n934), .B2(\mem[19][0] ), 
        .ZN(n935) );
  INV_X1 U191 ( .A(n933), .ZN(n658) );
  AOI22_X1 U192 ( .A1(data_in[1]), .A2(n824), .B1(n934), .B2(\mem[19][1] ), 
        .ZN(n933) );
  INV_X1 U193 ( .A(n932), .ZN(n657) );
  AOI22_X1 U194 ( .A1(data_in[2]), .A2(n824), .B1(n934), .B2(\mem[19][2] ), 
        .ZN(n932) );
  INV_X1 U195 ( .A(n931), .ZN(n656) );
  AOI22_X1 U196 ( .A1(data_in[3]), .A2(n824), .B1(n934), .B2(\mem[19][3] ), 
        .ZN(n931) );
  INV_X1 U197 ( .A(n930), .ZN(n655) );
  AOI22_X1 U198 ( .A1(data_in[4]), .A2(n824), .B1(n934), .B2(\mem[19][4] ), 
        .ZN(n930) );
  INV_X1 U199 ( .A(n929), .ZN(n654) );
  AOI22_X1 U200 ( .A1(data_in[5]), .A2(n824), .B1(n934), .B2(\mem[19][5] ), 
        .ZN(n929) );
  INV_X1 U201 ( .A(n928), .ZN(n653) );
  AOI22_X1 U202 ( .A1(data_in[6]), .A2(n824), .B1(n934), .B2(\mem[19][6] ), 
        .ZN(n928) );
  INV_X1 U203 ( .A(n927), .ZN(n652) );
  AOI22_X1 U204 ( .A1(data_in[7]), .A2(n824), .B1(n934), .B2(\mem[19][7] ), 
        .ZN(n927) );
  INV_X1 U205 ( .A(n908), .ZN(n635) );
  AOI22_X1 U206 ( .A1(data_in[0]), .A2(n821), .B1(n907), .B2(\mem[22][0] ), 
        .ZN(n908) );
  INV_X1 U207 ( .A(n906), .ZN(n634) );
  AOI22_X1 U208 ( .A1(data_in[1]), .A2(n821), .B1(n907), .B2(\mem[22][1] ), 
        .ZN(n906) );
  INV_X1 U209 ( .A(n905), .ZN(n633) );
  AOI22_X1 U210 ( .A1(data_in[2]), .A2(n821), .B1(n907), .B2(\mem[22][2] ), 
        .ZN(n905) );
  INV_X1 U211 ( .A(n904), .ZN(n632) );
  AOI22_X1 U212 ( .A1(data_in[3]), .A2(n821), .B1(n907), .B2(\mem[22][3] ), 
        .ZN(n904) );
  INV_X1 U213 ( .A(n903), .ZN(n631) );
  AOI22_X1 U214 ( .A1(data_in[4]), .A2(n821), .B1(n907), .B2(\mem[22][4] ), 
        .ZN(n903) );
  INV_X1 U215 ( .A(n902), .ZN(n630) );
  AOI22_X1 U216 ( .A1(data_in[5]), .A2(n821), .B1(n907), .B2(\mem[22][5] ), 
        .ZN(n902) );
  INV_X1 U217 ( .A(n901), .ZN(n629) );
  AOI22_X1 U218 ( .A1(data_in[6]), .A2(n821), .B1(n907), .B2(\mem[22][6] ), 
        .ZN(n901) );
  INV_X1 U219 ( .A(n900), .ZN(n628) );
  AOI22_X1 U220 ( .A1(data_in[7]), .A2(n821), .B1(n907), .B2(\mem[22][7] ), 
        .ZN(n900) );
  INV_X1 U221 ( .A(n899), .ZN(n627) );
  AOI22_X1 U222 ( .A1(data_in[0]), .A2(n820), .B1(n898), .B2(\mem[23][0] ), 
        .ZN(n899) );
  INV_X1 U223 ( .A(n897), .ZN(n626) );
  AOI22_X1 U224 ( .A1(data_in[1]), .A2(n820), .B1(n898), .B2(\mem[23][1] ), 
        .ZN(n897) );
  INV_X1 U225 ( .A(n896), .ZN(n625) );
  AOI22_X1 U226 ( .A1(data_in[2]), .A2(n820), .B1(n898), .B2(\mem[23][2] ), 
        .ZN(n896) );
  INV_X1 U227 ( .A(n895), .ZN(n624) );
  AOI22_X1 U228 ( .A1(data_in[3]), .A2(n820), .B1(n898), .B2(\mem[23][3] ), 
        .ZN(n895) );
  INV_X1 U229 ( .A(n894), .ZN(n623) );
  AOI22_X1 U230 ( .A1(data_in[4]), .A2(n820), .B1(n898), .B2(\mem[23][4] ), 
        .ZN(n894) );
  INV_X1 U231 ( .A(n893), .ZN(n622) );
  AOI22_X1 U232 ( .A1(data_in[5]), .A2(n820), .B1(n898), .B2(\mem[23][5] ), 
        .ZN(n893) );
  INV_X1 U233 ( .A(n892), .ZN(n621) );
  AOI22_X1 U234 ( .A1(data_in[6]), .A2(n820), .B1(n898), .B2(\mem[23][6] ), 
        .ZN(n892) );
  INV_X1 U235 ( .A(n891), .ZN(n620) );
  AOI22_X1 U236 ( .A1(data_in[7]), .A2(n820), .B1(n898), .B2(\mem[23][7] ), 
        .ZN(n891) );
  INV_X1 U237 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U238 ( .A1(data_in[0]), .A2(n837), .B1(n1053), .B2(\mem[6][0] ), 
        .ZN(n1054) );
  INV_X1 U239 ( .A(n1052), .ZN(n762) );
  AOI22_X1 U240 ( .A1(data_in[1]), .A2(n837), .B1(n1053), .B2(\mem[6][1] ), 
        .ZN(n1052) );
  INV_X1 U241 ( .A(n1051), .ZN(n761) );
  AOI22_X1 U242 ( .A1(data_in[2]), .A2(n837), .B1(n1053), .B2(\mem[6][2] ), 
        .ZN(n1051) );
  INV_X1 U243 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U244 ( .A1(data_in[3]), .A2(n837), .B1(n1053), .B2(\mem[6][3] ), 
        .ZN(n1050) );
  INV_X1 U245 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U246 ( .A1(data_in[4]), .A2(n837), .B1(n1053), .B2(\mem[6][4] ), 
        .ZN(n1049) );
  INV_X1 U247 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U248 ( .A1(data_in[5]), .A2(n837), .B1(n1053), .B2(\mem[6][5] ), 
        .ZN(n1048) );
  INV_X1 U249 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U250 ( .A1(data_in[6]), .A2(n837), .B1(n1053), .B2(\mem[6][6] ), 
        .ZN(n1047) );
  INV_X1 U251 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U252 ( .A1(data_in[7]), .A2(n837), .B1(n1053), .B2(\mem[6][7] ), 
        .ZN(n1046) );
  INV_X1 U253 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U254 ( .A1(data_in[0]), .A2(n836), .B1(n1044), .B2(\mem[7][0] ), 
        .ZN(n1045) );
  INV_X1 U255 ( .A(n1043), .ZN(n754) );
  AOI22_X1 U256 ( .A1(data_in[1]), .A2(n836), .B1(n1044), .B2(\mem[7][1] ), 
        .ZN(n1043) );
  INV_X1 U257 ( .A(n1042), .ZN(n753) );
  AOI22_X1 U258 ( .A1(data_in[2]), .A2(n836), .B1(n1044), .B2(\mem[7][2] ), 
        .ZN(n1042) );
  INV_X1 U259 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U260 ( .A1(data_in[3]), .A2(n836), .B1(n1044), .B2(\mem[7][3] ), 
        .ZN(n1041) );
  INV_X1 U261 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U262 ( .A1(data_in[4]), .A2(n836), .B1(n1044), .B2(\mem[7][4] ), 
        .ZN(n1040) );
  INV_X1 U263 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U264 ( .A1(data_in[5]), .A2(n836), .B1(n1044), .B2(\mem[7][5] ), 
        .ZN(n1039) );
  INV_X1 U265 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U266 ( .A1(data_in[6]), .A2(n836), .B1(n1044), .B2(\mem[7][6] ), 
        .ZN(n1038) );
  INV_X1 U267 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U268 ( .A1(data_in[7]), .A2(n836), .B1(n1044), .B2(\mem[7][7] ), 
        .ZN(n1037) );
  INV_X1 U269 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U270 ( .A1(data_in[0]), .A2(n833), .B1(n1016), .B2(\mem[10][0] ), 
        .ZN(n1017) );
  INV_X1 U271 ( .A(n1014), .ZN(n729) );
  AOI22_X1 U272 ( .A1(data_in[2]), .A2(n833), .B1(n1016), .B2(\mem[10][2] ), 
        .ZN(n1014) );
  INV_X1 U273 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U274 ( .A1(data_in[3]), .A2(n833), .B1(n1016), .B2(\mem[10][3] ), 
        .ZN(n1013) );
  INV_X1 U275 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U276 ( .A1(data_in[4]), .A2(n833), .B1(n1016), .B2(\mem[10][4] ), 
        .ZN(n1012) );
  INV_X1 U277 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U278 ( .A1(data_in[5]), .A2(n833), .B1(n1016), .B2(\mem[10][5] ), 
        .ZN(n1011) );
  INV_X1 U279 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U280 ( .A1(data_in[6]), .A2(n833), .B1(n1016), .B2(\mem[10][6] ), 
        .ZN(n1010) );
  INV_X1 U281 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U282 ( .A1(data_in[7]), .A2(n833), .B1(n1016), .B2(\mem[10][7] ), 
        .ZN(n1009) );
  INV_X1 U283 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U284 ( .A1(data_in[0]), .A2(n832), .B1(n1007), .B2(\mem[11][0] ), 
        .ZN(n1008) );
  INV_X1 U285 ( .A(n1006), .ZN(n722) );
  AOI22_X1 U286 ( .A1(data_in[1]), .A2(n832), .B1(n1007), .B2(\mem[11][1] ), 
        .ZN(n1006) );
  INV_X1 U287 ( .A(n1005), .ZN(n721) );
  AOI22_X1 U288 ( .A1(data_in[2]), .A2(n832), .B1(n1007), .B2(\mem[11][2] ), 
        .ZN(n1005) );
  INV_X1 U289 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U290 ( .A1(data_in[3]), .A2(n832), .B1(n1007), .B2(\mem[11][3] ), 
        .ZN(n1004) );
  INV_X1 U291 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U292 ( .A1(data_in[4]), .A2(n832), .B1(n1007), .B2(\mem[11][4] ), 
        .ZN(n1003) );
  INV_X1 U293 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U294 ( .A1(data_in[5]), .A2(n832), .B1(n1007), .B2(\mem[11][5] ), 
        .ZN(n1002) );
  INV_X1 U295 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U296 ( .A1(data_in[6]), .A2(n832), .B1(n1007), .B2(\mem[11][6] ), 
        .ZN(n1001) );
  INV_X1 U297 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U298 ( .A1(data_in[7]), .A2(n832), .B1(n1007), .B2(\mem[11][7] ), 
        .ZN(n1000) );
  INV_X1 U299 ( .A(n953), .ZN(n675) );
  AOI22_X1 U300 ( .A1(data_in[0]), .A2(n826), .B1(n952), .B2(\mem[17][0] ), 
        .ZN(n953) );
  INV_X1 U301 ( .A(n951), .ZN(n674) );
  AOI22_X1 U302 ( .A1(data_in[1]), .A2(n826), .B1(n952), .B2(\mem[17][1] ), 
        .ZN(n951) );
  INV_X1 U303 ( .A(n981), .ZN(n699) );
  AOI22_X1 U304 ( .A1(data_in[0]), .A2(n829), .B1(n980), .B2(\mem[14][0] ), 
        .ZN(n981) );
  INV_X1 U305 ( .A(n979), .ZN(n698) );
  AOI22_X1 U306 ( .A1(data_in[1]), .A2(n829), .B1(n980), .B2(\mem[14][1] ), 
        .ZN(n979) );
  INV_X1 U307 ( .A(n978), .ZN(n697) );
  AOI22_X1 U308 ( .A1(data_in[2]), .A2(n829), .B1(n980), .B2(\mem[14][2] ), 
        .ZN(n978) );
  INV_X1 U309 ( .A(n977), .ZN(n696) );
  AOI22_X1 U310 ( .A1(data_in[3]), .A2(n829), .B1(n980), .B2(\mem[14][3] ), 
        .ZN(n977) );
  INV_X1 U311 ( .A(n976), .ZN(n695) );
  AOI22_X1 U312 ( .A1(data_in[4]), .A2(n829), .B1(n980), .B2(\mem[14][4] ), 
        .ZN(n976) );
  INV_X1 U313 ( .A(n975), .ZN(n694) );
  AOI22_X1 U314 ( .A1(data_in[5]), .A2(n829), .B1(n980), .B2(\mem[14][5] ), 
        .ZN(n975) );
  INV_X1 U315 ( .A(n974), .ZN(n693) );
  AOI22_X1 U316 ( .A1(data_in[6]), .A2(n829), .B1(n980), .B2(\mem[14][6] ), 
        .ZN(n974) );
  INV_X1 U317 ( .A(n973), .ZN(n692) );
  AOI22_X1 U318 ( .A1(data_in[7]), .A2(n829), .B1(n980), .B2(\mem[14][7] ), 
        .ZN(n973) );
  INV_X1 U319 ( .A(n972), .ZN(n691) );
  AOI22_X1 U320 ( .A1(data_in[0]), .A2(n828), .B1(n971), .B2(\mem[15][0] ), 
        .ZN(n972) );
  INV_X1 U321 ( .A(n970), .ZN(n690) );
  AOI22_X1 U322 ( .A1(data_in[1]), .A2(n828), .B1(n971), .B2(\mem[15][1] ), 
        .ZN(n970) );
  INV_X1 U323 ( .A(n969), .ZN(n689) );
  AOI22_X1 U324 ( .A1(data_in[2]), .A2(n828), .B1(n971), .B2(\mem[15][2] ), 
        .ZN(n969) );
  INV_X1 U325 ( .A(n968), .ZN(n688) );
  AOI22_X1 U326 ( .A1(data_in[3]), .A2(n828), .B1(n971), .B2(\mem[15][3] ), 
        .ZN(n968) );
  INV_X1 U327 ( .A(n967), .ZN(n687) );
  AOI22_X1 U328 ( .A1(data_in[4]), .A2(n828), .B1(n971), .B2(\mem[15][4] ), 
        .ZN(n967) );
  INV_X1 U329 ( .A(n1015), .ZN(n730) );
  AOI22_X1 U330 ( .A1(data_in[1]), .A2(n833), .B1(n1016), .B2(\mem[10][1] ), 
        .ZN(n1015) );
  INV_X1 U331 ( .A(N12), .ZN(n255) );
  INV_X1 U332 ( .A(N11), .ZN(n254) );
  INV_X1 U333 ( .A(n999), .ZN(n715) );
  AOI22_X1 U334 ( .A1(data_in[0]), .A2(n831), .B1(n998), .B2(\mem[12][0] ), 
        .ZN(n999) );
  INV_X1 U335 ( .A(n997), .ZN(n714) );
  AOI22_X1 U336 ( .A1(data_in[1]), .A2(n831), .B1(n998), .B2(\mem[12][1] ), 
        .ZN(n997) );
  INV_X1 U337 ( .A(n996), .ZN(n713) );
  AOI22_X1 U338 ( .A1(data_in[2]), .A2(n831), .B1(n998), .B2(\mem[12][2] ), 
        .ZN(n996) );
  INV_X1 U339 ( .A(n995), .ZN(n712) );
  AOI22_X1 U340 ( .A1(data_in[3]), .A2(n831), .B1(n998), .B2(\mem[12][3] ), 
        .ZN(n995) );
  INV_X1 U341 ( .A(n994), .ZN(n711) );
  AOI22_X1 U342 ( .A1(data_in[4]), .A2(n831), .B1(n998), .B2(\mem[12][4] ), 
        .ZN(n994) );
  INV_X1 U343 ( .A(n993), .ZN(n710) );
  AOI22_X1 U344 ( .A1(data_in[5]), .A2(n831), .B1(n998), .B2(\mem[12][5] ), 
        .ZN(n993) );
  INV_X1 U345 ( .A(n992), .ZN(n709) );
  AOI22_X1 U346 ( .A1(data_in[6]), .A2(n831), .B1(n998), .B2(\mem[12][6] ), 
        .ZN(n992) );
  INV_X1 U347 ( .A(n991), .ZN(n708) );
  AOI22_X1 U348 ( .A1(data_in[7]), .A2(n831), .B1(n998), .B2(\mem[12][7] ), 
        .ZN(n991) );
  INV_X1 U349 ( .A(n926), .ZN(n651) );
  AOI22_X1 U350 ( .A1(data_in[0]), .A2(n823), .B1(n925), .B2(\mem[20][0] ), 
        .ZN(n926) );
  INV_X1 U351 ( .A(n924), .ZN(n650) );
  AOI22_X1 U352 ( .A1(data_in[1]), .A2(n823), .B1(n925), .B2(\mem[20][1] ), 
        .ZN(n924) );
  INV_X1 U353 ( .A(n923), .ZN(n649) );
  AOI22_X1 U354 ( .A1(data_in[2]), .A2(n823), .B1(n925), .B2(\mem[20][2] ), 
        .ZN(n923) );
  INV_X1 U355 ( .A(n922), .ZN(n648) );
  AOI22_X1 U356 ( .A1(data_in[3]), .A2(n823), .B1(n925), .B2(\mem[20][3] ), 
        .ZN(n922) );
  INV_X1 U357 ( .A(n921), .ZN(n647) );
  AOI22_X1 U358 ( .A1(data_in[4]), .A2(n823), .B1(n925), .B2(\mem[20][4] ), 
        .ZN(n921) );
  INV_X1 U359 ( .A(n920), .ZN(n646) );
  AOI22_X1 U360 ( .A1(data_in[5]), .A2(n823), .B1(n925), .B2(\mem[20][5] ), 
        .ZN(n920) );
  INV_X1 U361 ( .A(n919), .ZN(n645) );
  AOI22_X1 U362 ( .A1(data_in[6]), .A2(n823), .B1(n925), .B2(\mem[20][6] ), 
        .ZN(n919) );
  INV_X1 U363 ( .A(n918), .ZN(n644) );
  AOI22_X1 U364 ( .A1(data_in[7]), .A2(n823), .B1(n925), .B2(\mem[20][7] ), 
        .ZN(n918) );
  INV_X1 U365 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U366 ( .A1(data_in[0]), .A2(n835), .B1(n1035), .B2(\mem[8][0] ), 
        .ZN(n1036) );
  INV_X1 U367 ( .A(n1034), .ZN(n746) );
  AOI22_X1 U368 ( .A1(data_in[1]), .A2(n835), .B1(n1035), .B2(\mem[8][1] ), 
        .ZN(n1034) );
  INV_X1 U369 ( .A(n1033), .ZN(n745) );
  AOI22_X1 U370 ( .A1(data_in[2]), .A2(n835), .B1(n1035), .B2(\mem[8][2] ), 
        .ZN(n1033) );
  INV_X1 U371 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U372 ( .A1(data_in[3]), .A2(n835), .B1(n1035), .B2(\mem[8][3] ), 
        .ZN(n1032) );
  INV_X1 U373 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U374 ( .A1(data_in[4]), .A2(n835), .B1(n1035), .B2(\mem[8][4] ), 
        .ZN(n1031) );
  INV_X1 U375 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U376 ( .A1(data_in[5]), .A2(n835), .B1(n1035), .B2(\mem[8][5] ), 
        .ZN(n1030) );
  INV_X1 U377 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U378 ( .A1(data_in[6]), .A2(n835), .B1(n1035), .B2(\mem[8][6] ), 
        .ZN(n1029) );
  INV_X1 U379 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U380 ( .A1(data_in[7]), .A2(n835), .B1(n1035), .B2(\mem[8][7] ), 
        .ZN(n1028) );
  INV_X1 U381 ( .A(n963), .ZN(n683) );
  AOI22_X1 U382 ( .A1(data_in[0]), .A2(n827), .B1(n962), .B2(\mem[16][0] ), 
        .ZN(n963) );
  INV_X1 U383 ( .A(n961), .ZN(n682) );
  AOI22_X1 U384 ( .A1(data_in[1]), .A2(n827), .B1(n962), .B2(\mem[16][1] ), 
        .ZN(n961) );
  INV_X1 U385 ( .A(n960), .ZN(n681) );
  AOI22_X1 U386 ( .A1(data_in[2]), .A2(n827), .B1(n962), .B2(\mem[16][2] ), 
        .ZN(n960) );
  INV_X1 U387 ( .A(n959), .ZN(n680) );
  AOI22_X1 U388 ( .A1(data_in[3]), .A2(n827), .B1(n962), .B2(\mem[16][3] ), 
        .ZN(n959) );
  INV_X1 U389 ( .A(n958), .ZN(n679) );
  AOI22_X1 U390 ( .A1(data_in[4]), .A2(n827), .B1(n962), .B2(\mem[16][4] ), 
        .ZN(n958) );
  INV_X1 U391 ( .A(n957), .ZN(n678) );
  AOI22_X1 U392 ( .A1(data_in[5]), .A2(n827), .B1(n962), .B2(\mem[16][5] ), 
        .ZN(n957) );
  INV_X1 U393 ( .A(n956), .ZN(n677) );
  AOI22_X1 U394 ( .A1(data_in[6]), .A2(n827), .B1(n962), .B2(\mem[16][6] ), 
        .ZN(n956) );
  INV_X1 U395 ( .A(n955), .ZN(n676) );
  AOI22_X1 U396 ( .A1(data_in[7]), .A2(n827), .B1(n962), .B2(\mem[16][7] ), 
        .ZN(n955) );
  INV_X1 U397 ( .A(n890), .ZN(n619) );
  AOI22_X1 U398 ( .A1(data_in[0]), .A2(n816), .B1(n889), .B2(\mem[24][0] ), 
        .ZN(n890) );
  INV_X1 U399 ( .A(n888), .ZN(n618) );
  AOI22_X1 U400 ( .A1(data_in[1]), .A2(n816), .B1(n889), .B2(\mem[24][1] ), 
        .ZN(n888) );
  INV_X1 U401 ( .A(n887), .ZN(n617) );
  AOI22_X1 U402 ( .A1(data_in[2]), .A2(n816), .B1(n889), .B2(\mem[24][2] ), 
        .ZN(n887) );
  INV_X1 U403 ( .A(n886), .ZN(n616) );
  AOI22_X1 U404 ( .A1(data_in[3]), .A2(n816), .B1(n889), .B2(\mem[24][3] ), 
        .ZN(n886) );
  INV_X1 U405 ( .A(n885), .ZN(n615) );
  AOI22_X1 U406 ( .A1(data_in[4]), .A2(n816), .B1(n889), .B2(\mem[24][4] ), 
        .ZN(n885) );
  INV_X1 U407 ( .A(n884), .ZN(n614) );
  AOI22_X1 U408 ( .A1(data_in[5]), .A2(n816), .B1(n889), .B2(\mem[24][5] ), 
        .ZN(n884) );
  INV_X1 U409 ( .A(n883), .ZN(n613) );
  AOI22_X1 U410 ( .A1(data_in[6]), .A2(n816), .B1(n889), .B2(\mem[24][6] ), 
        .ZN(n883) );
  INV_X1 U411 ( .A(n882), .ZN(n612) );
  AOI22_X1 U412 ( .A1(data_in[7]), .A2(n816), .B1(n889), .B2(\mem[24][7] ), 
        .ZN(n882) );
  INV_X1 U413 ( .A(n881), .ZN(n611) );
  AOI22_X1 U414 ( .A1(data_in[0]), .A2(n815), .B1(n880), .B2(\mem[25][0] ), 
        .ZN(n881) );
  INV_X1 U415 ( .A(n879), .ZN(n610) );
  AOI22_X1 U416 ( .A1(data_in[1]), .A2(n815), .B1(n880), .B2(\mem[25][1] ), 
        .ZN(n879) );
  INV_X1 U417 ( .A(n878), .ZN(n609) );
  AOI22_X1 U418 ( .A1(data_in[2]), .A2(n815), .B1(n880), .B2(\mem[25][2] ), 
        .ZN(n878) );
  INV_X1 U419 ( .A(n877), .ZN(n608) );
  AOI22_X1 U420 ( .A1(data_in[3]), .A2(n815), .B1(n880), .B2(\mem[25][3] ), 
        .ZN(n877) );
  INV_X1 U421 ( .A(n876), .ZN(n607) );
  AOI22_X1 U422 ( .A1(data_in[4]), .A2(n815), .B1(n880), .B2(\mem[25][4] ), 
        .ZN(n876) );
  INV_X1 U423 ( .A(n875), .ZN(n606) );
  AOI22_X1 U424 ( .A1(data_in[5]), .A2(n815), .B1(n880), .B2(\mem[25][5] ), 
        .ZN(n875) );
  INV_X1 U425 ( .A(n874), .ZN(n605) );
  AOI22_X1 U426 ( .A1(data_in[6]), .A2(n815), .B1(n880), .B2(\mem[25][6] ), 
        .ZN(n874) );
  INV_X1 U427 ( .A(n873), .ZN(n604) );
  AOI22_X1 U428 ( .A1(data_in[7]), .A2(n815), .B1(n880), .B2(\mem[25][7] ), 
        .ZN(n873) );
  INV_X1 U429 ( .A(n872), .ZN(n603) );
  AOI22_X1 U430 ( .A1(data_in[0]), .A2(n814), .B1(n871), .B2(\mem[26][0] ), 
        .ZN(n872) );
  INV_X1 U431 ( .A(n870), .ZN(n602) );
  AOI22_X1 U432 ( .A1(data_in[1]), .A2(n814), .B1(n871), .B2(\mem[26][1] ), 
        .ZN(n870) );
  INV_X1 U433 ( .A(n869), .ZN(n601) );
  AOI22_X1 U434 ( .A1(data_in[2]), .A2(n814), .B1(n871), .B2(\mem[26][2] ), 
        .ZN(n869) );
  INV_X1 U435 ( .A(n868), .ZN(n600) );
  AOI22_X1 U436 ( .A1(data_in[3]), .A2(n814), .B1(n871), .B2(\mem[26][3] ), 
        .ZN(n868) );
  INV_X1 U437 ( .A(n867), .ZN(n599) );
  AOI22_X1 U438 ( .A1(data_in[4]), .A2(n814), .B1(n871), .B2(\mem[26][4] ), 
        .ZN(n867) );
  INV_X1 U439 ( .A(n866), .ZN(n598) );
  AOI22_X1 U440 ( .A1(data_in[5]), .A2(n814), .B1(n871), .B2(\mem[26][5] ), 
        .ZN(n866) );
  INV_X1 U441 ( .A(n865), .ZN(n597) );
  AOI22_X1 U442 ( .A1(data_in[6]), .A2(n814), .B1(n871), .B2(\mem[26][6] ), 
        .ZN(n865) );
  INV_X1 U443 ( .A(n864), .ZN(n596) );
  AOI22_X1 U444 ( .A1(data_in[7]), .A2(n814), .B1(n871), .B2(\mem[26][7] ), 
        .ZN(n864) );
  INV_X1 U445 ( .A(n863), .ZN(n595) );
  AOI22_X1 U446 ( .A1(data_in[0]), .A2(n813), .B1(n862), .B2(\mem[27][0] ), 
        .ZN(n863) );
  INV_X1 U447 ( .A(n861), .ZN(n594) );
  AOI22_X1 U448 ( .A1(data_in[1]), .A2(n813), .B1(n862), .B2(\mem[27][1] ), 
        .ZN(n861) );
  INV_X1 U449 ( .A(n860), .ZN(n293) );
  AOI22_X1 U450 ( .A1(data_in[2]), .A2(n813), .B1(n862), .B2(\mem[27][2] ), 
        .ZN(n860) );
  INV_X1 U451 ( .A(n859), .ZN(n292) );
  AOI22_X1 U452 ( .A1(data_in[3]), .A2(n813), .B1(n862), .B2(\mem[27][3] ), 
        .ZN(n859) );
  INV_X1 U453 ( .A(n858), .ZN(n291) );
  AOI22_X1 U454 ( .A1(data_in[4]), .A2(n813), .B1(n862), .B2(\mem[27][4] ), 
        .ZN(n858) );
  INV_X1 U455 ( .A(n857), .ZN(n290) );
  AOI22_X1 U456 ( .A1(data_in[5]), .A2(n813), .B1(n862), .B2(\mem[27][5] ), 
        .ZN(n857) );
  INV_X1 U457 ( .A(n856), .ZN(n289) );
  AOI22_X1 U458 ( .A1(data_in[6]), .A2(n813), .B1(n862), .B2(\mem[27][6] ), 
        .ZN(n856) );
  INV_X1 U459 ( .A(n855), .ZN(n288) );
  AOI22_X1 U460 ( .A1(data_in[7]), .A2(n813), .B1(n862), .B2(\mem[27][7] ), 
        .ZN(n855) );
  INV_X1 U461 ( .A(n854), .ZN(n287) );
  AOI22_X1 U462 ( .A1(data_in[0]), .A2(n812), .B1(n853), .B2(\mem[28][0] ), 
        .ZN(n854) );
  INV_X1 U463 ( .A(n852), .ZN(n286) );
  AOI22_X1 U464 ( .A1(data_in[1]), .A2(n812), .B1(n853), .B2(\mem[28][1] ), 
        .ZN(n852) );
  INV_X1 U465 ( .A(n851), .ZN(n285) );
  AOI22_X1 U466 ( .A1(data_in[2]), .A2(n812), .B1(n853), .B2(\mem[28][2] ), 
        .ZN(n851) );
  INV_X1 U467 ( .A(n850), .ZN(n284) );
  AOI22_X1 U468 ( .A1(data_in[3]), .A2(n812), .B1(n853), .B2(\mem[28][3] ), 
        .ZN(n850) );
  INV_X1 U469 ( .A(n849), .ZN(n283) );
  AOI22_X1 U470 ( .A1(data_in[4]), .A2(n812), .B1(n853), .B2(\mem[28][4] ), 
        .ZN(n849) );
  INV_X1 U471 ( .A(n848), .ZN(n282) );
  AOI22_X1 U472 ( .A1(data_in[5]), .A2(n812), .B1(n853), .B2(\mem[28][5] ), 
        .ZN(n848) );
  INV_X1 U473 ( .A(n847), .ZN(n281) );
  AOI22_X1 U474 ( .A1(data_in[6]), .A2(n812), .B1(n853), .B2(\mem[28][6] ), 
        .ZN(n847) );
  INV_X1 U475 ( .A(n846), .ZN(n280) );
  AOI22_X1 U476 ( .A1(data_in[7]), .A2(n812), .B1(n853), .B2(\mem[28][7] ), 
        .ZN(n846) );
  INV_X1 U477 ( .A(n1145), .ZN(n279) );
  AOI22_X1 U478 ( .A1(n819), .A2(data_in[0]), .B1(n1144), .B2(\mem[29][0] ), 
        .ZN(n1145) );
  INV_X1 U479 ( .A(n1143), .ZN(n278) );
  AOI22_X1 U480 ( .A1(n819), .A2(data_in[1]), .B1(n1144), .B2(\mem[29][1] ), 
        .ZN(n1143) );
  INV_X1 U481 ( .A(n1142), .ZN(n277) );
  AOI22_X1 U482 ( .A1(n819), .A2(data_in[2]), .B1(n1144), .B2(\mem[29][2] ), 
        .ZN(n1142) );
  INV_X1 U483 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U484 ( .A1(n819), .A2(data_in[3]), .B1(n1144), .B2(\mem[29][3] ), 
        .ZN(n1141) );
  INV_X1 U485 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U486 ( .A1(n819), .A2(data_in[4]), .B1(n1144), .B2(\mem[29][4] ), 
        .ZN(n1140) );
  INV_X1 U487 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U488 ( .A1(n819), .A2(data_in[5]), .B1(n1144), .B2(\mem[29][5] ), 
        .ZN(n1139) );
  INV_X1 U489 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U490 ( .A1(n819), .A2(data_in[6]), .B1(n1144), .B2(\mem[29][6] ), 
        .ZN(n1138) );
  INV_X1 U491 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U492 ( .A1(n819), .A2(data_in[7]), .B1(n1144), .B2(\mem[29][7] ), 
        .ZN(n1137) );
  INV_X1 U493 ( .A(n1134), .ZN(n271) );
  AOI22_X1 U494 ( .A1(data_in[0]), .A2(n818), .B1(n1133), .B2(\mem[30][0] ), 
        .ZN(n1134) );
  INV_X1 U495 ( .A(n1132), .ZN(n270) );
  AOI22_X1 U496 ( .A1(data_in[1]), .A2(n818), .B1(n1133), .B2(\mem[30][1] ), 
        .ZN(n1132) );
  INV_X1 U497 ( .A(n1131), .ZN(n269) );
  AOI22_X1 U498 ( .A1(data_in[2]), .A2(n818), .B1(n1133), .B2(\mem[30][2] ), 
        .ZN(n1131) );
  INV_X1 U499 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U500 ( .A1(data_in[3]), .A2(n818), .B1(n1133), .B2(\mem[30][3] ), 
        .ZN(n1130) );
  INV_X1 U501 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U502 ( .A1(data_in[4]), .A2(n818), .B1(n1133), .B2(\mem[30][4] ), 
        .ZN(n1129) );
  INV_X1 U503 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U504 ( .A1(data_in[5]), .A2(n818), .B1(n1133), .B2(\mem[30][5] ), 
        .ZN(n1128) );
  INV_X1 U505 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U506 ( .A1(data_in[6]), .A2(n818), .B1(n1133), .B2(\mem[30][6] ), 
        .ZN(n1127) );
  INV_X1 U507 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U508 ( .A1(data_in[7]), .A2(n818), .B1(n1133), .B2(\mem[30][7] ), 
        .ZN(n1126) );
  INV_X1 U509 ( .A(n1124), .ZN(n263) );
  AOI22_X1 U510 ( .A1(data_in[0]), .A2(n817), .B1(n1123), .B2(\mem[31][0] ), 
        .ZN(n1124) );
  INV_X1 U511 ( .A(n1122), .ZN(n262) );
  AOI22_X1 U512 ( .A1(data_in[1]), .A2(n817), .B1(n1123), .B2(\mem[31][1] ), 
        .ZN(n1122) );
  INV_X1 U513 ( .A(n1121), .ZN(n261) );
  AOI22_X1 U514 ( .A1(data_in[2]), .A2(n817), .B1(n1123), .B2(\mem[31][2] ), 
        .ZN(n1121) );
  INV_X1 U515 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U516 ( .A1(data_in[3]), .A2(n817), .B1(n1123), .B2(\mem[31][3] ), 
        .ZN(n1120) );
  INV_X1 U517 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U518 ( .A1(data_in[4]), .A2(n817), .B1(n1123), .B2(\mem[31][4] ), 
        .ZN(n1119) );
  INV_X1 U519 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U520 ( .A1(data_in[5]), .A2(n817), .B1(n1123), .B2(\mem[31][5] ), 
        .ZN(n1118) );
  INV_X1 U521 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U522 ( .A1(data_in[6]), .A2(n817), .B1(n1123), .B2(\mem[31][6] ), 
        .ZN(n1117) );
  INV_X1 U523 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U524 ( .A1(data_in[7]), .A2(n817), .B1(n1123), .B2(\mem[31][7] ), 
        .ZN(n1116) );
  INV_X1 U525 ( .A(n1114), .ZN(n811) );
  AOI22_X1 U526 ( .A1(data_in[0]), .A2(n843), .B1(n1113), .B2(\mem[0][0] ), 
        .ZN(n1114) );
  INV_X1 U527 ( .A(n1112), .ZN(n810) );
  AOI22_X1 U528 ( .A1(data_in[1]), .A2(n843), .B1(n1113), .B2(\mem[0][1] ), 
        .ZN(n1112) );
  INV_X1 U529 ( .A(n1111), .ZN(n809) );
  AOI22_X1 U530 ( .A1(data_in[2]), .A2(n843), .B1(n1113), .B2(\mem[0][2] ), 
        .ZN(n1111) );
  INV_X1 U531 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U532 ( .A1(data_in[3]), .A2(n843), .B1(n1113), .B2(\mem[0][3] ), 
        .ZN(n1110) );
  INV_X1 U533 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U534 ( .A1(data_in[4]), .A2(n843), .B1(n1113), .B2(\mem[0][4] ), 
        .ZN(n1109) );
  INV_X1 U535 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U536 ( .A1(data_in[5]), .A2(n843), .B1(n1113), .B2(\mem[0][5] ), 
        .ZN(n1108) );
  INV_X1 U537 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U538 ( .A1(data_in[6]), .A2(n843), .B1(n1113), .B2(\mem[0][6] ), 
        .ZN(n1107) );
  INV_X1 U539 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U540 ( .A1(data_in[7]), .A2(n843), .B1(n1113), .B2(\mem[0][7] ), 
        .ZN(n1106) );
  INV_X1 U541 ( .A(n1103), .ZN(n803) );
  AOI22_X1 U542 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[1][0] ), 
        .ZN(n1103) );
  INV_X1 U543 ( .A(n1101), .ZN(n802) );
  AOI22_X1 U544 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[1][1] ), 
        .ZN(n1101) );
  INV_X1 U545 ( .A(n1100), .ZN(n801) );
  AOI22_X1 U546 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[1][2] ), 
        .ZN(n1100) );
  INV_X1 U547 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U548 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[1][3] ), 
        .ZN(n1099) );
  INV_X1 U549 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U550 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[1][4] ), 
        .ZN(n1098) );
  INV_X1 U551 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U552 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[1][5] ), 
        .ZN(n1097) );
  INV_X1 U553 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U554 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[1][6] ), 
        .ZN(n1096) );
  INV_X1 U555 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U556 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[1][7] ), 
        .ZN(n1095) );
  INV_X1 U557 ( .A(n1093), .ZN(n795) );
  AOI22_X1 U558 ( .A1(data_in[0]), .A2(n841), .B1(n1092), .B2(\mem[2][0] ), 
        .ZN(n1093) );
  INV_X1 U559 ( .A(n1091), .ZN(n794) );
  AOI22_X1 U560 ( .A1(data_in[1]), .A2(n841), .B1(n1092), .B2(\mem[2][1] ), 
        .ZN(n1091) );
  INV_X1 U561 ( .A(n1090), .ZN(n793) );
  AOI22_X1 U562 ( .A1(data_in[2]), .A2(n841), .B1(n1092), .B2(\mem[2][2] ), 
        .ZN(n1090) );
  INV_X1 U563 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U564 ( .A1(data_in[3]), .A2(n841), .B1(n1092), .B2(\mem[2][3] ), 
        .ZN(n1089) );
  INV_X1 U565 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U566 ( .A1(data_in[4]), .A2(n841), .B1(n1092), .B2(\mem[2][4] ), 
        .ZN(n1088) );
  INV_X1 U567 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U568 ( .A1(data_in[5]), .A2(n841), .B1(n1092), .B2(\mem[2][5] ), 
        .ZN(n1087) );
  INV_X1 U569 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U570 ( .A1(data_in[6]), .A2(n841), .B1(n1092), .B2(\mem[2][6] ), 
        .ZN(n1086) );
  INV_X1 U571 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U572 ( .A1(data_in[7]), .A2(n841), .B1(n1092), .B2(\mem[2][7] ), 
        .ZN(n1085) );
  INV_X1 U573 ( .A(n1083), .ZN(n787) );
  AOI22_X1 U574 ( .A1(data_in[0]), .A2(n840), .B1(n1082), .B2(\mem[3][0] ), 
        .ZN(n1083) );
  INV_X1 U575 ( .A(n1081), .ZN(n786) );
  AOI22_X1 U576 ( .A1(data_in[1]), .A2(n840), .B1(n1082), .B2(\mem[3][1] ), 
        .ZN(n1081) );
  INV_X1 U577 ( .A(n1080), .ZN(n785) );
  AOI22_X1 U578 ( .A1(data_in[2]), .A2(n840), .B1(n1082), .B2(\mem[3][2] ), 
        .ZN(n1080) );
  INV_X1 U579 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U580 ( .A1(data_in[3]), .A2(n840), .B1(n1082), .B2(\mem[3][3] ), 
        .ZN(n1079) );
  INV_X1 U581 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U582 ( .A1(data_in[4]), .A2(n840), .B1(n1082), .B2(\mem[3][4] ), 
        .ZN(n1078) );
  INV_X1 U583 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U584 ( .A1(data_in[5]), .A2(n840), .B1(n1082), .B2(\mem[3][5] ), 
        .ZN(n1077) );
  INV_X1 U585 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U586 ( .A1(data_in[6]), .A2(n840), .B1(n1082), .B2(\mem[3][6] ), 
        .ZN(n1076) );
  INV_X1 U587 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U588 ( .A1(data_in[7]), .A2(n840), .B1(n1082), .B2(\mem[3][7] ), 
        .ZN(n1075) );
  INV_X1 U589 ( .A(n1073), .ZN(n779) );
  AOI22_X1 U590 ( .A1(data_in[0]), .A2(n839), .B1(n1072), .B2(\mem[4][0] ), 
        .ZN(n1073) );
  INV_X1 U591 ( .A(n1071), .ZN(n778) );
  AOI22_X1 U592 ( .A1(data_in[1]), .A2(n839), .B1(n1072), .B2(\mem[4][1] ), 
        .ZN(n1071) );
  INV_X1 U593 ( .A(n1070), .ZN(n777) );
  AOI22_X1 U594 ( .A1(data_in[2]), .A2(n839), .B1(n1072), .B2(\mem[4][2] ), 
        .ZN(n1070) );
  INV_X1 U595 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U596 ( .A1(data_in[3]), .A2(n839), .B1(n1072), .B2(\mem[4][3] ), 
        .ZN(n1069) );
  INV_X1 U597 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U598 ( .A1(data_in[4]), .A2(n839), .B1(n1072), .B2(\mem[4][4] ), 
        .ZN(n1068) );
  INV_X1 U599 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U600 ( .A1(data_in[5]), .A2(n839), .B1(n1072), .B2(\mem[4][5] ), 
        .ZN(n1067) );
  INV_X1 U601 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U602 ( .A1(data_in[6]), .A2(n839), .B1(n1072), .B2(\mem[4][6] ), 
        .ZN(n1066) );
  INV_X1 U603 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U604 ( .A1(data_in[7]), .A2(n839), .B1(n1072), .B2(\mem[4][7] ), 
        .ZN(n1065) );
  INV_X1 U605 ( .A(N13), .ZN(n844) );
  INV_X1 U606 ( .A(N14), .ZN(n845) );
  MUX2_X1 U607 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n250), .Z(n3) );
  MUX2_X1 U608 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n250), .Z(n4) );
  MUX2_X1 U609 ( .A(n4), .B(n3), .S(n245), .Z(n5) );
  MUX2_X1 U610 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n250), .Z(n6) );
  MUX2_X1 U611 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n250), .Z(n7) );
  MUX2_X1 U612 ( .A(n7), .B(n6), .S(N11), .Z(n8) );
  MUX2_X1 U613 ( .A(n8), .B(n5), .S(n243), .Z(n9) );
  MUX2_X1 U614 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n250), .Z(n10) );
  MUX2_X1 U615 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n249), .Z(n11) );
  MUX2_X1 U616 ( .A(n11), .B(n10), .S(n246), .Z(n12) );
  MUX2_X1 U617 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n250), .Z(n13) );
  MUX2_X1 U618 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n251), .Z(n14) );
  MUX2_X1 U619 ( .A(n14), .B(n13), .S(N11), .Z(n15) );
  MUX2_X1 U620 ( .A(n15), .B(n12), .S(N12), .Z(n16) );
  MUX2_X1 U621 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U622 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n247), .Z(n18) );
  MUX2_X1 U623 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n247), .Z(n19) );
  MUX2_X1 U624 ( .A(n19), .B(n18), .S(n244), .Z(n20) );
  MUX2_X1 U625 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n247), .Z(n21) );
  MUX2_X1 U626 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n247), .Z(n22) );
  MUX2_X1 U627 ( .A(n22), .B(n21), .S(n244), .Z(n23) );
  MUX2_X1 U628 ( .A(n23), .B(n20), .S(n243), .Z(n24) );
  MUX2_X1 U629 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n247), .Z(n25) );
  MUX2_X1 U630 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n247), .Z(n26) );
  MUX2_X1 U631 ( .A(n26), .B(n25), .S(n244), .Z(n27) );
  MUX2_X1 U632 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n247), .Z(n28) );
  MUX2_X1 U633 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n247), .Z(n29) );
  MUX2_X1 U634 ( .A(n29), .B(n28), .S(n244), .Z(n30) );
  MUX2_X1 U635 ( .A(n30), .B(n27), .S(n243), .Z(n31) );
  MUX2_X1 U636 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U637 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U638 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n247), .Z(n33) );
  MUX2_X1 U639 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n247), .Z(n34) );
  MUX2_X1 U640 ( .A(n34), .B(n33), .S(n244), .Z(n35) );
  MUX2_X1 U641 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n247), .Z(n36) );
  MUX2_X1 U642 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n247), .Z(n37) );
  MUX2_X1 U643 ( .A(n37), .B(n36), .S(n244), .Z(n38) );
  MUX2_X1 U644 ( .A(n38), .B(n35), .S(n243), .Z(n39) );
  MUX2_X1 U645 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n248), .Z(n40) );
  MUX2_X1 U646 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n248), .Z(n41) );
  MUX2_X1 U647 ( .A(n41), .B(n40), .S(n244), .Z(n42) );
  MUX2_X1 U648 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n248), .Z(n43) );
  MUX2_X1 U649 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n248), .Z(n44) );
  MUX2_X1 U650 ( .A(n44), .B(n43), .S(n244), .Z(n45) );
  MUX2_X1 U651 ( .A(n45), .B(n42), .S(n243), .Z(n46) );
  MUX2_X1 U652 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U653 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n248), .Z(n48) );
  MUX2_X1 U654 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n248), .Z(n49) );
  MUX2_X1 U655 ( .A(n49), .B(n48), .S(n244), .Z(n50) );
  MUX2_X1 U656 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n248), .Z(n51) );
  MUX2_X1 U657 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n248), .Z(n52) );
  MUX2_X1 U658 ( .A(n52), .B(n51), .S(n244), .Z(n53) );
  MUX2_X1 U659 ( .A(n53), .B(n50), .S(n243), .Z(n54) );
  MUX2_X1 U660 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n248), .Z(n55) );
  MUX2_X1 U661 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n248), .Z(n56) );
  MUX2_X1 U662 ( .A(n56), .B(n55), .S(n244), .Z(n57) );
  MUX2_X1 U663 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n248), .Z(n58) );
  MUX2_X1 U664 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n248), .Z(n59) );
  MUX2_X1 U665 ( .A(n59), .B(n58), .S(n244), .Z(n60) );
  MUX2_X1 U666 ( .A(n60), .B(n57), .S(n243), .Z(n61) );
  MUX2_X1 U667 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U668 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U669 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n247), .Z(n63) );
  MUX2_X1 U670 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n252), .Z(n64) );
  MUX2_X1 U671 ( .A(n64), .B(n63), .S(n245), .Z(n65) );
  MUX2_X1 U672 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n252), .Z(n66) );
  MUX2_X1 U673 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n247), .Z(n67) );
  MUX2_X1 U674 ( .A(n67), .B(n66), .S(n245), .Z(n68) );
  MUX2_X1 U675 ( .A(n68), .B(n65), .S(n243), .Z(n69) );
  MUX2_X1 U676 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n252), .Z(n70) );
  MUX2_X1 U677 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n251), .Z(n71) );
  MUX2_X1 U678 ( .A(n71), .B(n70), .S(n245), .Z(n72) );
  MUX2_X1 U679 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n252), .Z(n73) );
  MUX2_X1 U680 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n248), .Z(n74) );
  MUX2_X1 U681 ( .A(n74), .B(n73), .S(n245), .Z(n75) );
  MUX2_X1 U682 ( .A(n75), .B(n72), .S(n243), .Z(n76) );
  MUX2_X1 U683 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U684 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n249), .Z(n78) );
  MUX2_X1 U685 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n248), .Z(n79) );
  MUX2_X1 U686 ( .A(n79), .B(n78), .S(n245), .Z(n80) );
  MUX2_X1 U687 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n252), .Z(n81) );
  MUX2_X1 U688 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n249), .Z(n82) );
  MUX2_X1 U689 ( .A(n82), .B(n81), .S(n245), .Z(n83) );
  MUX2_X1 U690 ( .A(n83), .B(n80), .S(n243), .Z(n84) );
  MUX2_X1 U691 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n249), .Z(n85) );
  MUX2_X1 U692 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n252), .Z(n86) );
  MUX2_X1 U693 ( .A(n86), .B(n85), .S(n245), .Z(n87) );
  MUX2_X1 U694 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n252), .Z(n88) );
  MUX2_X1 U695 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n252), .Z(n89) );
  MUX2_X1 U696 ( .A(n89), .B(n88), .S(n245), .Z(n90) );
  MUX2_X1 U697 ( .A(n90), .B(n87), .S(n243), .Z(n91) );
  MUX2_X1 U698 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U699 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U700 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n249), .Z(n93) );
  MUX2_X1 U701 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n251), .Z(n94) );
  MUX2_X1 U702 ( .A(n94), .B(n93), .S(n245), .Z(n95) );
  MUX2_X1 U703 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n251), .Z(n96) );
  MUX2_X1 U704 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n252), .Z(n97) );
  MUX2_X1 U705 ( .A(n97), .B(n96), .S(n245), .Z(n98) );
  MUX2_X1 U706 ( .A(n98), .B(n95), .S(n243), .Z(n99) );
  MUX2_X1 U707 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n249), .Z(n100) );
  MUX2_X1 U708 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n252), .Z(n101) );
  MUX2_X1 U709 ( .A(n101), .B(n100), .S(n245), .Z(n102) );
  MUX2_X1 U710 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n248), .Z(n103) );
  MUX2_X1 U711 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n252), .Z(n104) );
  MUX2_X1 U712 ( .A(n104), .B(n103), .S(n245), .Z(n105) );
  MUX2_X1 U713 ( .A(n105), .B(n102), .S(n243), .Z(n106) );
  MUX2_X1 U714 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U715 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n249), .Z(n108) );
  MUX2_X1 U716 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n249), .Z(n109) );
  MUX2_X1 U717 ( .A(n109), .B(n108), .S(n246), .Z(n110) );
  MUX2_X1 U718 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n249), .Z(n111) );
  MUX2_X1 U719 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n249), .Z(n112) );
  MUX2_X1 U720 ( .A(n112), .B(n111), .S(n246), .Z(n113) );
  MUX2_X1 U721 ( .A(n113), .B(n110), .S(n243), .Z(n114) );
  MUX2_X1 U722 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n249), .Z(n115) );
  MUX2_X1 U723 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n249), .Z(n116) );
  MUX2_X1 U724 ( .A(n116), .B(n115), .S(n246), .Z(n117) );
  MUX2_X1 U725 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n249), .Z(n118) );
  MUX2_X1 U726 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n249), .Z(n119) );
  MUX2_X1 U727 ( .A(n119), .B(n118), .S(n246), .Z(n120) );
  MUX2_X1 U728 ( .A(n120), .B(n117), .S(n243), .Z(n121) );
  MUX2_X1 U729 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U730 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U731 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n249), .Z(n123) );
  MUX2_X1 U732 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n249), .Z(n124) );
  MUX2_X1 U733 ( .A(n124), .B(n123), .S(n246), .Z(n125) );
  MUX2_X1 U734 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n249), .Z(n126) );
  MUX2_X1 U735 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n249), .Z(n127) );
  MUX2_X1 U736 ( .A(n127), .B(n126), .S(n246), .Z(n128) );
  MUX2_X1 U737 ( .A(n128), .B(n125), .S(n243), .Z(n129) );
  MUX2_X1 U738 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n250), .Z(n130) );
  MUX2_X1 U739 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n250), .Z(n131) );
  MUX2_X1 U740 ( .A(n131), .B(n130), .S(n246), .Z(n132) );
  MUX2_X1 U741 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n250), .Z(n133) );
  MUX2_X1 U742 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n250), .Z(n134) );
  MUX2_X1 U743 ( .A(n134), .B(n133), .S(n246), .Z(n135) );
  MUX2_X1 U744 ( .A(n135), .B(n132), .S(n243), .Z(n136) );
  MUX2_X1 U745 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U746 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n250), .Z(n138) );
  MUX2_X1 U747 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n250), .Z(n139) );
  MUX2_X1 U748 ( .A(n139), .B(n138), .S(n246), .Z(n140) );
  MUX2_X1 U749 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n250), .Z(n141) );
  MUX2_X1 U750 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n250), .Z(n142) );
  MUX2_X1 U751 ( .A(n142), .B(n141), .S(n246), .Z(n143) );
  MUX2_X1 U752 ( .A(n143), .B(n140), .S(n243), .Z(n144) );
  MUX2_X1 U753 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n250), .Z(n145) );
  MUX2_X1 U754 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n250), .Z(n146) );
  MUX2_X1 U755 ( .A(n146), .B(n145), .S(n246), .Z(n147) );
  MUX2_X1 U756 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n250), .Z(n148) );
  MUX2_X1 U757 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n250), .Z(n149) );
  MUX2_X1 U758 ( .A(n149), .B(n148), .S(n246), .Z(n150) );
  MUX2_X1 U759 ( .A(n150), .B(n147), .S(n243), .Z(n151) );
  MUX2_X1 U760 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U761 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U762 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n251), .Z(n153) );
  MUX2_X1 U763 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n251), .Z(n154) );
  MUX2_X1 U764 ( .A(n154), .B(n153), .S(n245), .Z(n155) );
  MUX2_X1 U765 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n251), .Z(n156) );
  MUX2_X1 U766 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n251), .Z(n157) );
  MUX2_X1 U767 ( .A(n157), .B(n156), .S(N11), .Z(n158) );
  MUX2_X1 U768 ( .A(n158), .B(n155), .S(n243), .Z(n159) );
  MUX2_X1 U769 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n251), .Z(n160) );
  MUX2_X1 U770 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n251), .Z(n161) );
  MUX2_X1 U771 ( .A(n161), .B(n160), .S(N11), .Z(n162) );
  MUX2_X1 U772 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n251), .Z(n163) );
  MUX2_X1 U773 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n251), .Z(n164) );
  MUX2_X1 U774 ( .A(n164), .B(n163), .S(n245), .Z(n165) );
  MUX2_X1 U775 ( .A(n165), .B(n162), .S(N12), .Z(n166) );
  MUX2_X1 U776 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U777 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n251), .Z(n168) );
  MUX2_X1 U778 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n251), .Z(n169) );
  MUX2_X1 U779 ( .A(n169), .B(n168), .S(N11), .Z(n170) );
  MUX2_X1 U780 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n251), .Z(n171) );
  MUX2_X1 U781 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n251), .Z(n172) );
  MUX2_X1 U782 ( .A(n172), .B(n171), .S(N11), .Z(n173) );
  MUX2_X1 U783 ( .A(n173), .B(n170), .S(n243), .Z(n174) );
  MUX2_X1 U784 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n252), .Z(n175) );
  MUX2_X1 U785 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n252), .Z(n176) );
  MUX2_X1 U786 ( .A(n176), .B(n175), .S(N11), .Z(n177) );
  MUX2_X1 U787 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n252), .Z(n178) );
  MUX2_X1 U788 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n252), .Z(n179) );
  MUX2_X1 U789 ( .A(n179), .B(n178), .S(n244), .Z(n180) );
  MUX2_X1 U790 ( .A(n180), .B(n177), .S(N12), .Z(n181) );
  MUX2_X1 U791 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U792 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U793 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n248), .Z(n183) );
  MUX2_X1 U794 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n252), .Z(n184) );
  MUX2_X1 U795 ( .A(n184), .B(n183), .S(n246), .Z(n185) );
  MUX2_X1 U796 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n252), .Z(n186) );
  MUX2_X1 U797 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(N10), .Z(n187) );
  MUX2_X1 U798 ( .A(n187), .B(n186), .S(N11), .Z(n188) );
  MUX2_X1 U799 ( .A(n188), .B(n185), .S(n243), .Z(n189) );
  MUX2_X1 U800 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n250), .Z(n190) );
  MUX2_X1 U801 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(N10), .Z(n191) );
  MUX2_X1 U802 ( .A(n191), .B(n190), .S(N11), .Z(n192) );
  MUX2_X1 U803 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(N10), .Z(n193) );
  MUX2_X1 U804 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n252), .Z(n194) );
  MUX2_X1 U805 ( .A(n194), .B(n193), .S(n246), .Z(n195) );
  MUX2_X1 U806 ( .A(n195), .B(n192), .S(N12), .Z(n196) );
  MUX2_X1 U807 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U808 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n251), .Z(n198) );
  MUX2_X1 U809 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n252), .Z(n199) );
  MUX2_X1 U810 ( .A(n199), .B(n198), .S(n245), .Z(n200) );
  MUX2_X1 U811 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n248), .Z(n201) );
  MUX2_X1 U812 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n202) );
  MUX2_X1 U813 ( .A(n202), .B(n201), .S(n244), .Z(n203) );
  MUX2_X1 U814 ( .A(n203), .B(n200), .S(N12), .Z(n204) );
  MUX2_X1 U815 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n247), .Z(n205) );
  MUX2_X1 U816 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n206) );
  MUX2_X1 U817 ( .A(n206), .B(n205), .S(n245), .Z(n207) );
  MUX2_X1 U818 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n208) );
  MUX2_X1 U819 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n209) );
  MUX2_X1 U820 ( .A(n209), .B(n208), .S(N11), .Z(n210) );
  MUX2_X1 U821 ( .A(n210), .B(n207), .S(N12), .Z(n211) );
  MUX2_X1 U822 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U823 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U824 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n247), .Z(n213) );
  MUX2_X1 U825 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n247), .Z(n214) );
  MUX2_X1 U826 ( .A(n214), .B(n213), .S(n244), .Z(n215) );
  MUX2_X1 U827 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n251), .Z(n216) );
  MUX2_X1 U828 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(N10), .Z(n217) );
  MUX2_X1 U829 ( .A(n217), .B(n216), .S(n244), .Z(n218) );
  MUX2_X1 U830 ( .A(n218), .B(n215), .S(n243), .Z(n219) );
  MUX2_X1 U831 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n250), .Z(n220) );
  MUX2_X1 U832 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n252), .Z(n221) );
  MUX2_X1 U833 ( .A(n221), .B(n220), .S(N11), .Z(n222) );
  MUX2_X1 U834 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n250), .Z(n223) );
  MUX2_X1 U835 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n224) );
  MUX2_X1 U836 ( .A(n224), .B(n223), .S(N11), .Z(n225) );
  MUX2_X1 U837 ( .A(n225), .B(n222), .S(N12), .Z(n226) );
  MUX2_X1 U838 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U839 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n250), .Z(n228) );
  MUX2_X1 U840 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n248), .Z(n229) );
  MUX2_X1 U841 ( .A(n229), .B(n228), .S(n246), .Z(n230) );
  MUX2_X1 U842 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n250), .Z(n231) );
  MUX2_X1 U843 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n232) );
  MUX2_X1 U844 ( .A(n232), .B(n231), .S(n244), .Z(n233) );
  MUX2_X1 U845 ( .A(n233), .B(n230), .S(N12), .Z(n234) );
  MUX2_X1 U846 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n235) );
  MUX2_X1 U847 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n236) );
  MUX2_X1 U848 ( .A(n236), .B(n235), .S(n246), .Z(n237) );
  MUX2_X1 U849 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n238) );
  MUX2_X1 U850 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n239) );
  MUX2_X1 U851 ( .A(n239), .B(n238), .S(N11), .Z(n240) );
  MUX2_X1 U852 ( .A(n240), .B(n237), .S(N12), .Z(n241) );
  MUX2_X1 U853 ( .A(n241), .B(n234), .S(N13), .Z(n242) );
  MUX2_X1 U854 ( .A(n242), .B(n227), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_19 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n256), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n257), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n258), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n259), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n260), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n261), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n262), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n263), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n264), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n265), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n266), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n267), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n268), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n269), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n270), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n271), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n272), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n273), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n274), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n275), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n276), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n277), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n278), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n279), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n280), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n281), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n282), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n283), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n284), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n285), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n286), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n287), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n288), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n289), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n290), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n291), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n292), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n293), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n594), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n595), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n596), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n597), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n598), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n599), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n600), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n601), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n602), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n603), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n604), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n605), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n606), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n607), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n608), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n609), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n610), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n611), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n612), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n613), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n614), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n615), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n616), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n617), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n618), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n619), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n620), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n621), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n622), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n623), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n624), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n625), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n626), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n627), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n628), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n629), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n630), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n631), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n632), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n633), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n634), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n635), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n636), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n637), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n638), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n639), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n640), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n641), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n642), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n643), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n644), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n645), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n646), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n647), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n648), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n649), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n650), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n651), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n652), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n653), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n654), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n655), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n656), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n657), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n658), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n659), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n660), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n661), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n662), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n663), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n664), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n665), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n666), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n667), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n668), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n669), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n670), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n671), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n672), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n673), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n674), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n675), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n676), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n677), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n678), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n679), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n680), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n681), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n682), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n683), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n684), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n685), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n686), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n687), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n688), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n689), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n690), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n691), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n692), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n693), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n694), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n695), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n696), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n697), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n698), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n699), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n700), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n701), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n702), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n703), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n704), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n705), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n706), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n707), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n708), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n709), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n710), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n711), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n712), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n713), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n714), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n715), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n716), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n717), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n718), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n719), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n720), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n721), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n722), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n723), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n724), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n725), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n726), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n727), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n728), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n729), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n730), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n731), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n732), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n733), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n734), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n735), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n736), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n737), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n738), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n739), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n740), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n741), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n742), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n743), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n744), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n745), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n746), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n747), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n748), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n749), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n750), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n751), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n752), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n753), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n754), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n755), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n756), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n757), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n758), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n759), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n760), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n761), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n762), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n763), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n764), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n765), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n766), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n767), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n768), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n769), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n770), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n771), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n772), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n773), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n774), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n775), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n776), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n777), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n778), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n779), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n780), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n781), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n782), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n783), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n784), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n785), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n786), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n787), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n788), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n789), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n790), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n791), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n792), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n793), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n794), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n795), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n796), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n797), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n798), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n799), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n800), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n801), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n802), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n803), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n804), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n805), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n806), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n807), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n808), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n809), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n810), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n811), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X2 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(n252), .Z(n249) );
  BUF_X1 U5 ( .A(n252), .Z(n250) );
  BUF_X1 U6 ( .A(N10), .Z(n251) );
  BUF_X1 U7 ( .A(n252), .Z(n248) );
  BUF_X1 U8 ( .A(n252), .Z(n247) );
  BUF_X1 U9 ( .A(N10), .Z(n252) );
  INV_X1 U10 ( .A(n1113), .ZN(n843) );
  INV_X1 U11 ( .A(n1102), .ZN(n842) );
  INV_X1 U12 ( .A(n1092), .ZN(n841) );
  INV_X1 U13 ( .A(n1082), .ZN(n840) );
  INV_X1 U14 ( .A(n1072), .ZN(n839) );
  INV_X1 U15 ( .A(n1062), .ZN(n838) );
  INV_X1 U16 ( .A(n1053), .ZN(n837) );
  INV_X1 U17 ( .A(n1044), .ZN(n836) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1105) );
  NOR3_X1 U19 ( .A1(N11), .A2(N12), .A3(n253), .ZN(n1094) );
  NAND2_X1 U20 ( .A1(n1104), .A2(n1136), .ZN(n1062) );
  NAND2_X1 U21 ( .A1(n1105), .A2(n1104), .ZN(n1113) );
  NAND2_X1 U22 ( .A1(n1094), .A2(n1104), .ZN(n1102) );
  NAND2_X1 U23 ( .A1(n1084), .A2(n1104), .ZN(n1092) );
  NAND2_X1 U24 ( .A1(n1074), .A2(n1104), .ZN(n1082) );
  NAND2_X1 U25 ( .A1(n1064), .A2(n1104), .ZN(n1072) );
  NAND2_X1 U26 ( .A1(n1104), .A2(n1125), .ZN(n1053) );
  NAND2_X1 U27 ( .A1(n1104), .A2(n1115), .ZN(n1044) );
  INV_X1 U28 ( .A(n1133), .ZN(n818) );
  INV_X1 U29 ( .A(n1123), .ZN(n817) );
  INV_X1 U30 ( .A(n889), .ZN(n816) );
  INV_X1 U31 ( .A(n880), .ZN(n815) );
  INV_X1 U32 ( .A(n871), .ZN(n814) );
  INV_X1 U33 ( .A(n862), .ZN(n813) );
  INV_X1 U34 ( .A(n853), .ZN(n812) );
  INV_X1 U35 ( .A(n989), .ZN(n830) );
  INV_X1 U36 ( .A(n980), .ZN(n829) );
  INV_X1 U37 ( .A(n971), .ZN(n828) );
  INV_X1 U38 ( .A(n916), .ZN(n822) );
  INV_X1 U39 ( .A(n907), .ZN(n821) );
  INV_X1 U40 ( .A(n898), .ZN(n820) );
  INV_X1 U41 ( .A(n1035), .ZN(n835) );
  INV_X1 U42 ( .A(n1025), .ZN(n834) );
  INV_X1 U43 ( .A(n1016), .ZN(n833) );
  INV_X1 U44 ( .A(n1007), .ZN(n832) );
  INV_X1 U45 ( .A(n998), .ZN(n831) );
  INV_X1 U46 ( .A(n962), .ZN(n827) );
  INV_X1 U47 ( .A(n952), .ZN(n826) );
  INV_X1 U48 ( .A(n943), .ZN(n825) );
  INV_X1 U49 ( .A(n934), .ZN(n824) );
  INV_X1 U50 ( .A(n925), .ZN(n823) );
  INV_X1 U51 ( .A(n1144), .ZN(n819) );
  BUF_X1 U52 ( .A(N11), .Z(n244) );
  BUF_X1 U53 ( .A(N11), .Z(n245) );
  BUF_X1 U54 ( .A(N11), .Z(n246) );
  INV_X1 U55 ( .A(N10), .ZN(n253) );
  BUF_X1 U56 ( .A(N12), .Z(n243) );
  NOR3_X1 U57 ( .A1(n255), .A2(N10), .A3(n254), .ZN(n1125) );
  NOR3_X1 U58 ( .A1(n255), .A2(n253), .A3(n254), .ZN(n1115) );
  NOR3_X1 U59 ( .A1(n253), .A2(N11), .A3(n255), .ZN(n1136) );
  NOR3_X1 U60 ( .A1(N10), .A2(N12), .A3(n254), .ZN(n1084) );
  NOR3_X1 U61 ( .A1(n253), .A2(N12), .A3(n254), .ZN(n1074) );
  NOR3_X1 U62 ( .A1(N10), .A2(N11), .A3(n255), .ZN(n1064) );
  NAND2_X1 U63 ( .A1(n1027), .A2(n1136), .ZN(n989) );
  NAND2_X1 U64 ( .A1(n954), .A2(n1136), .ZN(n916) );
  NAND2_X1 U65 ( .A1(n1027), .A2(n1064), .ZN(n998) );
  NAND2_X1 U66 ( .A1(n954), .A2(n1064), .ZN(n925) );
  NAND2_X1 U67 ( .A1(n1027), .A2(n1105), .ZN(n1035) );
  NAND2_X1 U68 ( .A1(n1027), .A2(n1094), .ZN(n1025) );
  NAND2_X1 U69 ( .A1(n954), .A2(n1105), .ZN(n962) );
  NAND2_X1 U70 ( .A1(n954), .A2(n1094), .ZN(n952) );
  NAND2_X1 U71 ( .A1(n1105), .A2(n1135), .ZN(n889) );
  NAND2_X1 U72 ( .A1(n1094), .A2(n1135), .ZN(n880) );
  NAND2_X1 U73 ( .A1(n1084), .A2(n1135), .ZN(n871) );
  NAND2_X1 U74 ( .A1(n1074), .A2(n1135), .ZN(n862) );
  NAND2_X1 U75 ( .A1(n1064), .A2(n1135), .ZN(n853) );
  NAND2_X1 U76 ( .A1(n1136), .A2(n1135), .ZN(n1144) );
  NAND2_X1 U77 ( .A1(n1125), .A2(n1135), .ZN(n1133) );
  NAND2_X1 U78 ( .A1(n1115), .A2(n1135), .ZN(n1123) );
  NAND2_X1 U79 ( .A1(n1027), .A2(n1084), .ZN(n1016) );
  NAND2_X1 U80 ( .A1(n1027), .A2(n1074), .ZN(n1007) );
  NAND2_X1 U81 ( .A1(n954), .A2(n1084), .ZN(n943) );
  NAND2_X1 U82 ( .A1(n954), .A2(n1074), .ZN(n934) );
  NAND2_X1 U83 ( .A1(n1027), .A2(n1125), .ZN(n980) );
  NAND2_X1 U84 ( .A1(n954), .A2(n1125), .ZN(n907) );
  NAND2_X1 U85 ( .A1(n1027), .A2(n1115), .ZN(n971) );
  NAND2_X1 U86 ( .A1(n954), .A2(n1115), .ZN(n898) );
  AND3_X1 U87 ( .A1(n844), .A2(n845), .A3(wr_en), .ZN(n1104) );
  AND3_X1 U88 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1135) );
  AND3_X1 U89 ( .A1(N13), .A2(n845), .A3(wr_en), .ZN(n1027) );
  AND3_X1 U90 ( .A1(N14), .A2(n844), .A3(wr_en), .ZN(n954) );
  INV_X1 U91 ( .A(n1063), .ZN(n771) );
  AOI22_X1 U92 ( .A1(data_in[0]), .A2(n838), .B1(n1062), .B2(\mem[5][0] ), 
        .ZN(n1063) );
  INV_X1 U93 ( .A(n1061), .ZN(n770) );
  AOI22_X1 U94 ( .A1(data_in[1]), .A2(n838), .B1(n1062), .B2(\mem[5][1] ), 
        .ZN(n1061) );
  INV_X1 U95 ( .A(n1060), .ZN(n769) );
  AOI22_X1 U96 ( .A1(data_in[2]), .A2(n838), .B1(n1062), .B2(\mem[5][2] ), 
        .ZN(n1060) );
  INV_X1 U97 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U98 ( .A1(data_in[3]), .A2(n838), .B1(n1062), .B2(\mem[5][3] ), 
        .ZN(n1059) );
  INV_X1 U99 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U100 ( .A1(data_in[4]), .A2(n838), .B1(n1062), .B2(\mem[5][4] ), 
        .ZN(n1058) );
  INV_X1 U101 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U102 ( .A1(data_in[5]), .A2(n838), .B1(n1062), .B2(\mem[5][5] ), 
        .ZN(n1057) );
  INV_X1 U103 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U104 ( .A1(data_in[6]), .A2(n838), .B1(n1062), .B2(\mem[5][6] ), 
        .ZN(n1056) );
  INV_X1 U105 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U106 ( .A1(data_in[7]), .A2(n838), .B1(n1062), .B2(\mem[5][7] ), 
        .ZN(n1055) );
  INV_X1 U107 ( .A(n1026), .ZN(n739) );
  AOI22_X1 U108 ( .A1(data_in[0]), .A2(n834), .B1(n1025), .B2(\mem[9][0] ), 
        .ZN(n1026) );
  INV_X1 U109 ( .A(n1024), .ZN(n738) );
  AOI22_X1 U110 ( .A1(data_in[1]), .A2(n834), .B1(n1025), .B2(\mem[9][1] ), 
        .ZN(n1024) );
  INV_X1 U111 ( .A(n1023), .ZN(n737) );
  AOI22_X1 U112 ( .A1(data_in[2]), .A2(n834), .B1(n1025), .B2(\mem[9][2] ), 
        .ZN(n1023) );
  INV_X1 U113 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U114 ( .A1(data_in[3]), .A2(n834), .B1(n1025), .B2(\mem[9][3] ), 
        .ZN(n1022) );
  INV_X1 U115 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U116 ( .A1(data_in[4]), .A2(n834), .B1(n1025), .B2(\mem[9][4] ), 
        .ZN(n1021) );
  INV_X1 U117 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U118 ( .A1(data_in[5]), .A2(n834), .B1(n1025), .B2(\mem[9][5] ), 
        .ZN(n1020) );
  INV_X1 U119 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U120 ( .A1(data_in[6]), .A2(n834), .B1(n1025), .B2(\mem[9][6] ), 
        .ZN(n1019) );
  INV_X1 U121 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U122 ( .A1(data_in[7]), .A2(n834), .B1(n1025), .B2(\mem[9][7] ), 
        .ZN(n1018) );
  INV_X1 U123 ( .A(n990), .ZN(n707) );
  AOI22_X1 U124 ( .A1(data_in[0]), .A2(n830), .B1(n989), .B2(\mem[13][0] ), 
        .ZN(n990) );
  INV_X1 U125 ( .A(n988), .ZN(n706) );
  AOI22_X1 U126 ( .A1(data_in[1]), .A2(n830), .B1(n989), .B2(\mem[13][1] ), 
        .ZN(n988) );
  INV_X1 U127 ( .A(n987), .ZN(n705) );
  AOI22_X1 U128 ( .A1(data_in[2]), .A2(n830), .B1(n989), .B2(\mem[13][2] ), 
        .ZN(n987) );
  INV_X1 U129 ( .A(n986), .ZN(n704) );
  AOI22_X1 U130 ( .A1(data_in[3]), .A2(n830), .B1(n989), .B2(\mem[13][3] ), 
        .ZN(n986) );
  INV_X1 U131 ( .A(n985), .ZN(n703) );
  AOI22_X1 U132 ( .A1(data_in[4]), .A2(n830), .B1(n989), .B2(\mem[13][4] ), 
        .ZN(n985) );
  INV_X1 U133 ( .A(n984), .ZN(n702) );
  AOI22_X1 U134 ( .A1(data_in[5]), .A2(n830), .B1(n989), .B2(\mem[13][5] ), 
        .ZN(n984) );
  INV_X1 U135 ( .A(n983), .ZN(n701) );
  AOI22_X1 U136 ( .A1(data_in[6]), .A2(n830), .B1(n989), .B2(\mem[13][6] ), 
        .ZN(n983) );
  INV_X1 U137 ( .A(n982), .ZN(n700) );
  AOI22_X1 U138 ( .A1(data_in[7]), .A2(n830), .B1(n989), .B2(\mem[13][7] ), 
        .ZN(n982) );
  INV_X1 U139 ( .A(n953), .ZN(n675) );
  AOI22_X1 U140 ( .A1(data_in[0]), .A2(n826), .B1(n952), .B2(\mem[17][0] ), 
        .ZN(n953) );
  INV_X1 U141 ( .A(n951), .ZN(n674) );
  AOI22_X1 U142 ( .A1(data_in[1]), .A2(n826), .B1(n952), .B2(\mem[17][1] ), 
        .ZN(n951) );
  INV_X1 U143 ( .A(n950), .ZN(n673) );
  AOI22_X1 U144 ( .A1(data_in[2]), .A2(n826), .B1(n952), .B2(\mem[17][2] ), 
        .ZN(n950) );
  INV_X1 U145 ( .A(n949), .ZN(n672) );
  AOI22_X1 U146 ( .A1(data_in[3]), .A2(n826), .B1(n952), .B2(\mem[17][3] ), 
        .ZN(n949) );
  INV_X1 U147 ( .A(n948), .ZN(n671) );
  AOI22_X1 U148 ( .A1(data_in[4]), .A2(n826), .B1(n952), .B2(\mem[17][4] ), 
        .ZN(n948) );
  INV_X1 U149 ( .A(n947), .ZN(n670) );
  AOI22_X1 U150 ( .A1(data_in[5]), .A2(n826), .B1(n952), .B2(\mem[17][5] ), 
        .ZN(n947) );
  INV_X1 U151 ( .A(n946), .ZN(n669) );
  AOI22_X1 U152 ( .A1(data_in[6]), .A2(n826), .B1(n952), .B2(\mem[17][6] ), 
        .ZN(n946) );
  INV_X1 U153 ( .A(n945), .ZN(n668) );
  AOI22_X1 U154 ( .A1(data_in[7]), .A2(n826), .B1(n952), .B2(\mem[17][7] ), 
        .ZN(n945) );
  INV_X1 U155 ( .A(n917), .ZN(n643) );
  AOI22_X1 U156 ( .A1(data_in[0]), .A2(n822), .B1(n916), .B2(\mem[21][0] ), 
        .ZN(n917) );
  INV_X1 U157 ( .A(n915), .ZN(n642) );
  AOI22_X1 U158 ( .A1(data_in[1]), .A2(n822), .B1(n916), .B2(\mem[21][1] ), 
        .ZN(n915) );
  INV_X1 U159 ( .A(n914), .ZN(n641) );
  AOI22_X1 U160 ( .A1(data_in[2]), .A2(n822), .B1(n916), .B2(\mem[21][2] ), 
        .ZN(n914) );
  INV_X1 U161 ( .A(n913), .ZN(n640) );
  AOI22_X1 U162 ( .A1(data_in[3]), .A2(n822), .B1(n916), .B2(\mem[21][3] ), 
        .ZN(n913) );
  INV_X1 U163 ( .A(n912), .ZN(n639) );
  AOI22_X1 U164 ( .A1(data_in[4]), .A2(n822), .B1(n916), .B2(\mem[21][4] ), 
        .ZN(n912) );
  INV_X1 U165 ( .A(n911), .ZN(n638) );
  AOI22_X1 U166 ( .A1(data_in[5]), .A2(n822), .B1(n916), .B2(\mem[21][5] ), 
        .ZN(n911) );
  INV_X1 U167 ( .A(n910), .ZN(n637) );
  AOI22_X1 U168 ( .A1(data_in[6]), .A2(n822), .B1(n916), .B2(\mem[21][6] ), 
        .ZN(n910) );
  INV_X1 U169 ( .A(n909), .ZN(n636) );
  AOI22_X1 U170 ( .A1(data_in[7]), .A2(n822), .B1(n916), .B2(\mem[21][7] ), 
        .ZN(n909) );
  INV_X1 U171 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U172 ( .A1(data_in[0]), .A2(n837), .B1(n1053), .B2(\mem[6][0] ), 
        .ZN(n1054) );
  INV_X1 U173 ( .A(n1052), .ZN(n762) );
  AOI22_X1 U174 ( .A1(data_in[1]), .A2(n837), .B1(n1053), .B2(\mem[6][1] ), 
        .ZN(n1052) );
  INV_X1 U175 ( .A(n1051), .ZN(n761) );
  AOI22_X1 U176 ( .A1(data_in[2]), .A2(n837), .B1(n1053), .B2(\mem[6][2] ), 
        .ZN(n1051) );
  INV_X1 U177 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U178 ( .A1(data_in[3]), .A2(n837), .B1(n1053), .B2(\mem[6][3] ), 
        .ZN(n1050) );
  INV_X1 U179 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U180 ( .A1(data_in[4]), .A2(n837), .B1(n1053), .B2(\mem[6][4] ), 
        .ZN(n1049) );
  INV_X1 U181 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U182 ( .A1(data_in[5]), .A2(n837), .B1(n1053), .B2(\mem[6][5] ), 
        .ZN(n1048) );
  INV_X1 U183 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U184 ( .A1(data_in[6]), .A2(n837), .B1(n1053), .B2(\mem[6][6] ), 
        .ZN(n1047) );
  INV_X1 U185 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U186 ( .A1(data_in[7]), .A2(n837), .B1(n1053), .B2(\mem[6][7] ), 
        .ZN(n1046) );
  INV_X1 U187 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U188 ( .A1(data_in[0]), .A2(n836), .B1(n1044), .B2(\mem[7][0] ), 
        .ZN(n1045) );
  INV_X1 U189 ( .A(n1043), .ZN(n754) );
  AOI22_X1 U190 ( .A1(data_in[1]), .A2(n836), .B1(n1044), .B2(\mem[7][1] ), 
        .ZN(n1043) );
  INV_X1 U191 ( .A(n1042), .ZN(n753) );
  AOI22_X1 U192 ( .A1(data_in[2]), .A2(n836), .B1(n1044), .B2(\mem[7][2] ), 
        .ZN(n1042) );
  INV_X1 U193 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U194 ( .A1(data_in[3]), .A2(n836), .B1(n1044), .B2(\mem[7][3] ), 
        .ZN(n1041) );
  INV_X1 U195 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U196 ( .A1(data_in[4]), .A2(n836), .B1(n1044), .B2(\mem[7][4] ), 
        .ZN(n1040) );
  INV_X1 U197 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U198 ( .A1(data_in[5]), .A2(n836), .B1(n1044), .B2(\mem[7][5] ), 
        .ZN(n1039) );
  INV_X1 U199 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U200 ( .A1(data_in[6]), .A2(n836), .B1(n1044), .B2(\mem[7][6] ), 
        .ZN(n1038) );
  INV_X1 U201 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U202 ( .A1(data_in[7]), .A2(n836), .B1(n1044), .B2(\mem[7][7] ), 
        .ZN(n1037) );
  INV_X1 U203 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U204 ( .A1(data_in[0]), .A2(n833), .B1(n1016), .B2(\mem[10][0] ), 
        .ZN(n1017) );
  INV_X1 U205 ( .A(n1015), .ZN(n730) );
  AOI22_X1 U206 ( .A1(data_in[1]), .A2(n833), .B1(n1016), .B2(\mem[10][1] ), 
        .ZN(n1015) );
  INV_X1 U207 ( .A(n1014), .ZN(n729) );
  AOI22_X1 U208 ( .A1(data_in[2]), .A2(n833), .B1(n1016), .B2(\mem[10][2] ), 
        .ZN(n1014) );
  INV_X1 U209 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U210 ( .A1(data_in[3]), .A2(n833), .B1(n1016), .B2(\mem[10][3] ), 
        .ZN(n1013) );
  INV_X1 U211 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U212 ( .A1(data_in[4]), .A2(n833), .B1(n1016), .B2(\mem[10][4] ), 
        .ZN(n1012) );
  INV_X1 U213 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U214 ( .A1(data_in[6]), .A2(n833), .B1(n1016), .B2(\mem[10][6] ), 
        .ZN(n1010) );
  INV_X1 U215 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U216 ( .A1(data_in[7]), .A2(n833), .B1(n1016), .B2(\mem[10][7] ), 
        .ZN(n1009) );
  INV_X1 U217 ( .A(n1006), .ZN(n722) );
  AOI22_X1 U218 ( .A1(data_in[1]), .A2(n832), .B1(n1007), .B2(\mem[11][1] ), 
        .ZN(n1006) );
  INV_X1 U219 ( .A(n1005), .ZN(n721) );
  AOI22_X1 U220 ( .A1(data_in[2]), .A2(n832), .B1(n1007), .B2(\mem[11][2] ), 
        .ZN(n1005) );
  INV_X1 U221 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U222 ( .A1(data_in[3]), .A2(n832), .B1(n1007), .B2(\mem[11][3] ), 
        .ZN(n1004) );
  INV_X1 U223 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U224 ( .A1(data_in[4]), .A2(n832), .B1(n1007), .B2(\mem[11][4] ), 
        .ZN(n1003) );
  INV_X1 U225 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U226 ( .A1(data_in[5]), .A2(n832), .B1(n1007), .B2(\mem[11][5] ), 
        .ZN(n1002) );
  INV_X1 U227 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U228 ( .A1(data_in[6]), .A2(n832), .B1(n1007), .B2(\mem[11][6] ), 
        .ZN(n1001) );
  INV_X1 U229 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U230 ( .A1(data_in[7]), .A2(n832), .B1(n1007), .B2(\mem[11][7] ), 
        .ZN(n1000) );
  INV_X1 U231 ( .A(n975), .ZN(n694) );
  AOI22_X1 U232 ( .A1(data_in[5]), .A2(n829), .B1(n980), .B2(\mem[14][5] ), 
        .ZN(n975) );
  INV_X1 U233 ( .A(n974), .ZN(n693) );
  AOI22_X1 U234 ( .A1(data_in[6]), .A2(n829), .B1(n980), .B2(\mem[14][6] ), 
        .ZN(n974) );
  INV_X1 U235 ( .A(n973), .ZN(n692) );
  AOI22_X1 U236 ( .A1(data_in[7]), .A2(n829), .B1(n980), .B2(\mem[14][7] ), 
        .ZN(n973) );
  INV_X1 U237 ( .A(n972), .ZN(n691) );
  AOI22_X1 U238 ( .A1(data_in[0]), .A2(n828), .B1(n971), .B2(\mem[15][0] ), 
        .ZN(n972) );
  INV_X1 U239 ( .A(n970), .ZN(n690) );
  AOI22_X1 U240 ( .A1(data_in[1]), .A2(n828), .B1(n971), .B2(\mem[15][1] ), 
        .ZN(n970) );
  INV_X1 U241 ( .A(n969), .ZN(n689) );
  AOI22_X1 U242 ( .A1(data_in[2]), .A2(n828), .B1(n971), .B2(\mem[15][2] ), 
        .ZN(n969) );
  INV_X1 U243 ( .A(n968), .ZN(n688) );
  AOI22_X1 U244 ( .A1(data_in[3]), .A2(n828), .B1(n971), .B2(\mem[15][3] ), 
        .ZN(n968) );
  INV_X1 U245 ( .A(n967), .ZN(n687) );
  AOI22_X1 U246 ( .A1(data_in[4]), .A2(n828), .B1(n971), .B2(\mem[15][4] ), 
        .ZN(n967) );
  INV_X1 U247 ( .A(n966), .ZN(n686) );
  AOI22_X1 U248 ( .A1(data_in[5]), .A2(n828), .B1(n971), .B2(\mem[15][5] ), 
        .ZN(n966) );
  INV_X1 U249 ( .A(n965), .ZN(n685) );
  AOI22_X1 U250 ( .A1(data_in[6]), .A2(n828), .B1(n971), .B2(\mem[15][6] ), 
        .ZN(n965) );
  INV_X1 U251 ( .A(n964), .ZN(n684) );
  AOI22_X1 U252 ( .A1(data_in[7]), .A2(n828), .B1(n971), .B2(\mem[15][7] ), 
        .ZN(n964) );
  INV_X1 U253 ( .A(n944), .ZN(n667) );
  AOI22_X1 U254 ( .A1(data_in[0]), .A2(n825), .B1(n943), .B2(\mem[18][0] ), 
        .ZN(n944) );
  INV_X1 U255 ( .A(n942), .ZN(n666) );
  AOI22_X1 U256 ( .A1(data_in[1]), .A2(n825), .B1(n943), .B2(\mem[18][1] ), 
        .ZN(n942) );
  INV_X1 U257 ( .A(n941), .ZN(n665) );
  AOI22_X1 U258 ( .A1(data_in[2]), .A2(n825), .B1(n943), .B2(\mem[18][2] ), 
        .ZN(n941) );
  INV_X1 U259 ( .A(n940), .ZN(n664) );
  AOI22_X1 U260 ( .A1(data_in[3]), .A2(n825), .B1(n943), .B2(\mem[18][3] ), 
        .ZN(n940) );
  INV_X1 U261 ( .A(n939), .ZN(n663) );
  AOI22_X1 U262 ( .A1(data_in[4]), .A2(n825), .B1(n943), .B2(\mem[18][4] ), 
        .ZN(n939) );
  INV_X1 U263 ( .A(n938), .ZN(n662) );
  AOI22_X1 U264 ( .A1(data_in[5]), .A2(n825), .B1(n943), .B2(\mem[18][5] ), 
        .ZN(n938) );
  INV_X1 U265 ( .A(n937), .ZN(n661) );
  AOI22_X1 U266 ( .A1(data_in[6]), .A2(n825), .B1(n943), .B2(\mem[18][6] ), 
        .ZN(n937) );
  INV_X1 U267 ( .A(n936), .ZN(n660) );
  AOI22_X1 U268 ( .A1(data_in[7]), .A2(n825), .B1(n943), .B2(\mem[18][7] ), 
        .ZN(n936) );
  INV_X1 U269 ( .A(n935), .ZN(n659) );
  AOI22_X1 U270 ( .A1(data_in[0]), .A2(n824), .B1(n934), .B2(\mem[19][0] ), 
        .ZN(n935) );
  INV_X1 U271 ( .A(n933), .ZN(n658) );
  AOI22_X1 U272 ( .A1(data_in[1]), .A2(n824), .B1(n934), .B2(\mem[19][1] ), 
        .ZN(n933) );
  INV_X1 U273 ( .A(n932), .ZN(n657) );
  AOI22_X1 U274 ( .A1(data_in[2]), .A2(n824), .B1(n934), .B2(\mem[19][2] ), 
        .ZN(n932) );
  INV_X1 U275 ( .A(n931), .ZN(n656) );
  AOI22_X1 U276 ( .A1(data_in[3]), .A2(n824), .B1(n934), .B2(\mem[19][3] ), 
        .ZN(n931) );
  INV_X1 U277 ( .A(n930), .ZN(n655) );
  AOI22_X1 U278 ( .A1(data_in[4]), .A2(n824), .B1(n934), .B2(\mem[19][4] ), 
        .ZN(n930) );
  INV_X1 U279 ( .A(n929), .ZN(n654) );
  AOI22_X1 U280 ( .A1(data_in[5]), .A2(n824), .B1(n934), .B2(\mem[19][5] ), 
        .ZN(n929) );
  INV_X1 U281 ( .A(n928), .ZN(n653) );
  AOI22_X1 U282 ( .A1(data_in[6]), .A2(n824), .B1(n934), .B2(\mem[19][6] ), 
        .ZN(n928) );
  INV_X1 U283 ( .A(n927), .ZN(n652) );
  AOI22_X1 U284 ( .A1(data_in[7]), .A2(n824), .B1(n934), .B2(\mem[19][7] ), 
        .ZN(n927) );
  INV_X1 U285 ( .A(n908), .ZN(n635) );
  AOI22_X1 U286 ( .A1(data_in[0]), .A2(n821), .B1(n907), .B2(\mem[22][0] ), 
        .ZN(n908) );
  INV_X1 U287 ( .A(n906), .ZN(n634) );
  AOI22_X1 U288 ( .A1(data_in[1]), .A2(n821), .B1(n907), .B2(\mem[22][1] ), 
        .ZN(n906) );
  INV_X1 U289 ( .A(n905), .ZN(n633) );
  AOI22_X1 U290 ( .A1(data_in[2]), .A2(n821), .B1(n907), .B2(\mem[22][2] ), 
        .ZN(n905) );
  INV_X1 U291 ( .A(n904), .ZN(n632) );
  AOI22_X1 U292 ( .A1(data_in[3]), .A2(n821), .B1(n907), .B2(\mem[22][3] ), 
        .ZN(n904) );
  INV_X1 U293 ( .A(n903), .ZN(n631) );
  AOI22_X1 U294 ( .A1(data_in[4]), .A2(n821), .B1(n907), .B2(\mem[22][4] ), 
        .ZN(n903) );
  INV_X1 U295 ( .A(n902), .ZN(n630) );
  AOI22_X1 U296 ( .A1(data_in[5]), .A2(n821), .B1(n907), .B2(\mem[22][5] ), 
        .ZN(n902) );
  INV_X1 U297 ( .A(n901), .ZN(n629) );
  AOI22_X1 U298 ( .A1(data_in[6]), .A2(n821), .B1(n907), .B2(\mem[22][6] ), 
        .ZN(n901) );
  INV_X1 U299 ( .A(n900), .ZN(n628) );
  AOI22_X1 U300 ( .A1(data_in[7]), .A2(n821), .B1(n907), .B2(\mem[22][7] ), 
        .ZN(n900) );
  INV_X1 U301 ( .A(n899), .ZN(n627) );
  AOI22_X1 U302 ( .A1(data_in[0]), .A2(n820), .B1(n898), .B2(\mem[23][0] ), 
        .ZN(n899) );
  INV_X1 U303 ( .A(n897), .ZN(n626) );
  AOI22_X1 U304 ( .A1(data_in[1]), .A2(n820), .B1(n898), .B2(\mem[23][1] ), 
        .ZN(n897) );
  INV_X1 U305 ( .A(n896), .ZN(n625) );
  AOI22_X1 U306 ( .A1(data_in[2]), .A2(n820), .B1(n898), .B2(\mem[23][2] ), 
        .ZN(n896) );
  INV_X1 U307 ( .A(n895), .ZN(n624) );
  AOI22_X1 U308 ( .A1(data_in[3]), .A2(n820), .B1(n898), .B2(\mem[23][3] ), 
        .ZN(n895) );
  INV_X1 U309 ( .A(n894), .ZN(n623) );
  AOI22_X1 U310 ( .A1(data_in[4]), .A2(n820), .B1(n898), .B2(\mem[23][4] ), 
        .ZN(n894) );
  INV_X1 U311 ( .A(n893), .ZN(n622) );
  AOI22_X1 U312 ( .A1(data_in[5]), .A2(n820), .B1(n898), .B2(\mem[23][5] ), 
        .ZN(n893) );
  INV_X1 U313 ( .A(n892), .ZN(n621) );
  AOI22_X1 U314 ( .A1(data_in[6]), .A2(n820), .B1(n898), .B2(\mem[23][6] ), 
        .ZN(n892) );
  INV_X1 U315 ( .A(n891), .ZN(n620) );
  AOI22_X1 U316 ( .A1(data_in[7]), .A2(n820), .B1(n898), .B2(\mem[23][7] ), 
        .ZN(n891) );
  INV_X1 U317 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U318 ( .A1(data_in[5]), .A2(n833), .B1(n1016), .B2(\mem[10][5] ), 
        .ZN(n1011) );
  INV_X1 U319 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U320 ( .A1(data_in[0]), .A2(n832), .B1(n1007), .B2(\mem[11][0] ), 
        .ZN(n1008) );
  INV_X1 U321 ( .A(n981), .ZN(n699) );
  AOI22_X1 U322 ( .A1(data_in[0]), .A2(n829), .B1(n980), .B2(\mem[14][0] ), 
        .ZN(n981) );
  INV_X1 U323 ( .A(n979), .ZN(n698) );
  AOI22_X1 U324 ( .A1(data_in[1]), .A2(n829), .B1(n980), .B2(\mem[14][1] ), 
        .ZN(n979) );
  INV_X1 U325 ( .A(n978), .ZN(n697) );
  AOI22_X1 U326 ( .A1(data_in[2]), .A2(n829), .B1(n980), .B2(\mem[14][2] ), 
        .ZN(n978) );
  INV_X1 U327 ( .A(n977), .ZN(n696) );
  AOI22_X1 U328 ( .A1(data_in[3]), .A2(n829), .B1(n980), .B2(\mem[14][3] ), 
        .ZN(n977) );
  INV_X1 U329 ( .A(n976), .ZN(n695) );
  AOI22_X1 U330 ( .A1(data_in[4]), .A2(n829), .B1(n980), .B2(\mem[14][4] ), 
        .ZN(n976) );
  INV_X1 U331 ( .A(N12), .ZN(n255) );
  INV_X1 U332 ( .A(N11), .ZN(n254) );
  INV_X1 U333 ( .A(n999), .ZN(n715) );
  AOI22_X1 U334 ( .A1(data_in[0]), .A2(n831), .B1(n998), .B2(\mem[12][0] ), 
        .ZN(n999) );
  INV_X1 U335 ( .A(n997), .ZN(n714) );
  AOI22_X1 U336 ( .A1(data_in[1]), .A2(n831), .B1(n998), .B2(\mem[12][1] ), 
        .ZN(n997) );
  INV_X1 U337 ( .A(n996), .ZN(n713) );
  AOI22_X1 U338 ( .A1(data_in[2]), .A2(n831), .B1(n998), .B2(\mem[12][2] ), 
        .ZN(n996) );
  INV_X1 U339 ( .A(n995), .ZN(n712) );
  AOI22_X1 U340 ( .A1(data_in[3]), .A2(n831), .B1(n998), .B2(\mem[12][3] ), 
        .ZN(n995) );
  INV_X1 U341 ( .A(n994), .ZN(n711) );
  AOI22_X1 U342 ( .A1(data_in[4]), .A2(n831), .B1(n998), .B2(\mem[12][4] ), 
        .ZN(n994) );
  INV_X1 U343 ( .A(n993), .ZN(n710) );
  AOI22_X1 U344 ( .A1(data_in[5]), .A2(n831), .B1(n998), .B2(\mem[12][5] ), 
        .ZN(n993) );
  INV_X1 U345 ( .A(n992), .ZN(n709) );
  AOI22_X1 U346 ( .A1(data_in[6]), .A2(n831), .B1(n998), .B2(\mem[12][6] ), 
        .ZN(n992) );
  INV_X1 U347 ( .A(n991), .ZN(n708) );
  AOI22_X1 U348 ( .A1(data_in[7]), .A2(n831), .B1(n998), .B2(\mem[12][7] ), 
        .ZN(n991) );
  INV_X1 U349 ( .A(n926), .ZN(n651) );
  AOI22_X1 U350 ( .A1(data_in[0]), .A2(n823), .B1(n925), .B2(\mem[20][0] ), 
        .ZN(n926) );
  INV_X1 U351 ( .A(n924), .ZN(n650) );
  AOI22_X1 U352 ( .A1(data_in[1]), .A2(n823), .B1(n925), .B2(\mem[20][1] ), 
        .ZN(n924) );
  INV_X1 U353 ( .A(n923), .ZN(n649) );
  AOI22_X1 U354 ( .A1(data_in[2]), .A2(n823), .B1(n925), .B2(\mem[20][2] ), 
        .ZN(n923) );
  INV_X1 U355 ( .A(n922), .ZN(n648) );
  AOI22_X1 U356 ( .A1(data_in[3]), .A2(n823), .B1(n925), .B2(\mem[20][3] ), 
        .ZN(n922) );
  INV_X1 U357 ( .A(n921), .ZN(n647) );
  AOI22_X1 U358 ( .A1(data_in[4]), .A2(n823), .B1(n925), .B2(\mem[20][4] ), 
        .ZN(n921) );
  INV_X1 U359 ( .A(n920), .ZN(n646) );
  AOI22_X1 U360 ( .A1(data_in[5]), .A2(n823), .B1(n925), .B2(\mem[20][5] ), 
        .ZN(n920) );
  INV_X1 U361 ( .A(n919), .ZN(n645) );
  AOI22_X1 U362 ( .A1(data_in[6]), .A2(n823), .B1(n925), .B2(\mem[20][6] ), 
        .ZN(n919) );
  INV_X1 U363 ( .A(n918), .ZN(n644) );
  AOI22_X1 U364 ( .A1(data_in[7]), .A2(n823), .B1(n925), .B2(\mem[20][7] ), 
        .ZN(n918) );
  INV_X1 U365 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U366 ( .A1(data_in[0]), .A2(n835), .B1(n1035), .B2(\mem[8][0] ), 
        .ZN(n1036) );
  INV_X1 U367 ( .A(n1034), .ZN(n746) );
  AOI22_X1 U368 ( .A1(data_in[1]), .A2(n835), .B1(n1035), .B2(\mem[8][1] ), 
        .ZN(n1034) );
  INV_X1 U369 ( .A(n1033), .ZN(n745) );
  AOI22_X1 U370 ( .A1(data_in[2]), .A2(n835), .B1(n1035), .B2(\mem[8][2] ), 
        .ZN(n1033) );
  INV_X1 U371 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U372 ( .A1(data_in[3]), .A2(n835), .B1(n1035), .B2(\mem[8][3] ), 
        .ZN(n1032) );
  INV_X1 U373 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U374 ( .A1(data_in[4]), .A2(n835), .B1(n1035), .B2(\mem[8][4] ), 
        .ZN(n1031) );
  INV_X1 U375 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U376 ( .A1(data_in[5]), .A2(n835), .B1(n1035), .B2(\mem[8][5] ), 
        .ZN(n1030) );
  INV_X1 U377 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U378 ( .A1(data_in[6]), .A2(n835), .B1(n1035), .B2(\mem[8][6] ), 
        .ZN(n1029) );
  INV_X1 U379 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U380 ( .A1(data_in[7]), .A2(n835), .B1(n1035), .B2(\mem[8][7] ), 
        .ZN(n1028) );
  INV_X1 U381 ( .A(n963), .ZN(n683) );
  AOI22_X1 U382 ( .A1(data_in[0]), .A2(n827), .B1(n962), .B2(\mem[16][0] ), 
        .ZN(n963) );
  INV_X1 U383 ( .A(n961), .ZN(n682) );
  AOI22_X1 U384 ( .A1(data_in[1]), .A2(n827), .B1(n962), .B2(\mem[16][1] ), 
        .ZN(n961) );
  INV_X1 U385 ( .A(n960), .ZN(n681) );
  AOI22_X1 U386 ( .A1(data_in[2]), .A2(n827), .B1(n962), .B2(\mem[16][2] ), 
        .ZN(n960) );
  INV_X1 U387 ( .A(n959), .ZN(n680) );
  AOI22_X1 U388 ( .A1(data_in[3]), .A2(n827), .B1(n962), .B2(\mem[16][3] ), 
        .ZN(n959) );
  INV_X1 U389 ( .A(n958), .ZN(n679) );
  AOI22_X1 U390 ( .A1(data_in[4]), .A2(n827), .B1(n962), .B2(\mem[16][4] ), 
        .ZN(n958) );
  INV_X1 U391 ( .A(n957), .ZN(n678) );
  AOI22_X1 U392 ( .A1(data_in[5]), .A2(n827), .B1(n962), .B2(\mem[16][5] ), 
        .ZN(n957) );
  INV_X1 U393 ( .A(n956), .ZN(n677) );
  AOI22_X1 U394 ( .A1(data_in[6]), .A2(n827), .B1(n962), .B2(\mem[16][6] ), 
        .ZN(n956) );
  INV_X1 U395 ( .A(n955), .ZN(n676) );
  AOI22_X1 U396 ( .A1(data_in[7]), .A2(n827), .B1(n962), .B2(\mem[16][7] ), 
        .ZN(n955) );
  INV_X1 U397 ( .A(n890), .ZN(n619) );
  AOI22_X1 U398 ( .A1(data_in[0]), .A2(n816), .B1(n889), .B2(\mem[24][0] ), 
        .ZN(n890) );
  INV_X1 U399 ( .A(n888), .ZN(n618) );
  AOI22_X1 U400 ( .A1(data_in[1]), .A2(n816), .B1(n889), .B2(\mem[24][1] ), 
        .ZN(n888) );
  INV_X1 U401 ( .A(n887), .ZN(n617) );
  AOI22_X1 U402 ( .A1(data_in[2]), .A2(n816), .B1(n889), .B2(\mem[24][2] ), 
        .ZN(n887) );
  INV_X1 U403 ( .A(n886), .ZN(n616) );
  AOI22_X1 U404 ( .A1(data_in[3]), .A2(n816), .B1(n889), .B2(\mem[24][3] ), 
        .ZN(n886) );
  INV_X1 U405 ( .A(n885), .ZN(n615) );
  AOI22_X1 U406 ( .A1(data_in[4]), .A2(n816), .B1(n889), .B2(\mem[24][4] ), 
        .ZN(n885) );
  INV_X1 U407 ( .A(n884), .ZN(n614) );
  AOI22_X1 U408 ( .A1(data_in[5]), .A2(n816), .B1(n889), .B2(\mem[24][5] ), 
        .ZN(n884) );
  INV_X1 U409 ( .A(n883), .ZN(n613) );
  AOI22_X1 U410 ( .A1(data_in[6]), .A2(n816), .B1(n889), .B2(\mem[24][6] ), 
        .ZN(n883) );
  INV_X1 U411 ( .A(n882), .ZN(n612) );
  AOI22_X1 U412 ( .A1(data_in[7]), .A2(n816), .B1(n889), .B2(\mem[24][7] ), 
        .ZN(n882) );
  INV_X1 U413 ( .A(n881), .ZN(n611) );
  AOI22_X1 U414 ( .A1(data_in[0]), .A2(n815), .B1(n880), .B2(\mem[25][0] ), 
        .ZN(n881) );
  INV_X1 U415 ( .A(n879), .ZN(n610) );
  AOI22_X1 U416 ( .A1(data_in[1]), .A2(n815), .B1(n880), .B2(\mem[25][1] ), 
        .ZN(n879) );
  INV_X1 U417 ( .A(n878), .ZN(n609) );
  AOI22_X1 U418 ( .A1(data_in[2]), .A2(n815), .B1(n880), .B2(\mem[25][2] ), 
        .ZN(n878) );
  INV_X1 U419 ( .A(n877), .ZN(n608) );
  AOI22_X1 U420 ( .A1(data_in[3]), .A2(n815), .B1(n880), .B2(\mem[25][3] ), 
        .ZN(n877) );
  INV_X1 U421 ( .A(n876), .ZN(n607) );
  AOI22_X1 U422 ( .A1(data_in[4]), .A2(n815), .B1(n880), .B2(\mem[25][4] ), 
        .ZN(n876) );
  INV_X1 U423 ( .A(n875), .ZN(n606) );
  AOI22_X1 U424 ( .A1(data_in[5]), .A2(n815), .B1(n880), .B2(\mem[25][5] ), 
        .ZN(n875) );
  INV_X1 U425 ( .A(n874), .ZN(n605) );
  AOI22_X1 U426 ( .A1(data_in[6]), .A2(n815), .B1(n880), .B2(\mem[25][6] ), 
        .ZN(n874) );
  INV_X1 U427 ( .A(n873), .ZN(n604) );
  AOI22_X1 U428 ( .A1(data_in[7]), .A2(n815), .B1(n880), .B2(\mem[25][7] ), 
        .ZN(n873) );
  INV_X1 U429 ( .A(n872), .ZN(n603) );
  AOI22_X1 U430 ( .A1(data_in[0]), .A2(n814), .B1(n871), .B2(\mem[26][0] ), 
        .ZN(n872) );
  INV_X1 U431 ( .A(n870), .ZN(n602) );
  AOI22_X1 U432 ( .A1(data_in[1]), .A2(n814), .B1(n871), .B2(\mem[26][1] ), 
        .ZN(n870) );
  INV_X1 U433 ( .A(n869), .ZN(n601) );
  AOI22_X1 U434 ( .A1(data_in[2]), .A2(n814), .B1(n871), .B2(\mem[26][2] ), 
        .ZN(n869) );
  INV_X1 U435 ( .A(n868), .ZN(n600) );
  AOI22_X1 U436 ( .A1(data_in[3]), .A2(n814), .B1(n871), .B2(\mem[26][3] ), 
        .ZN(n868) );
  INV_X1 U437 ( .A(n867), .ZN(n599) );
  AOI22_X1 U438 ( .A1(data_in[4]), .A2(n814), .B1(n871), .B2(\mem[26][4] ), 
        .ZN(n867) );
  INV_X1 U439 ( .A(n866), .ZN(n598) );
  AOI22_X1 U440 ( .A1(data_in[5]), .A2(n814), .B1(n871), .B2(\mem[26][5] ), 
        .ZN(n866) );
  INV_X1 U441 ( .A(n865), .ZN(n597) );
  AOI22_X1 U442 ( .A1(data_in[6]), .A2(n814), .B1(n871), .B2(\mem[26][6] ), 
        .ZN(n865) );
  INV_X1 U443 ( .A(n864), .ZN(n596) );
  AOI22_X1 U444 ( .A1(data_in[7]), .A2(n814), .B1(n871), .B2(\mem[26][7] ), 
        .ZN(n864) );
  INV_X1 U445 ( .A(n863), .ZN(n595) );
  AOI22_X1 U446 ( .A1(data_in[0]), .A2(n813), .B1(n862), .B2(\mem[27][0] ), 
        .ZN(n863) );
  INV_X1 U447 ( .A(n861), .ZN(n594) );
  AOI22_X1 U448 ( .A1(data_in[1]), .A2(n813), .B1(n862), .B2(\mem[27][1] ), 
        .ZN(n861) );
  INV_X1 U449 ( .A(n860), .ZN(n293) );
  AOI22_X1 U450 ( .A1(data_in[2]), .A2(n813), .B1(n862), .B2(\mem[27][2] ), 
        .ZN(n860) );
  INV_X1 U451 ( .A(n859), .ZN(n292) );
  AOI22_X1 U452 ( .A1(data_in[3]), .A2(n813), .B1(n862), .B2(\mem[27][3] ), 
        .ZN(n859) );
  INV_X1 U453 ( .A(n858), .ZN(n291) );
  AOI22_X1 U454 ( .A1(data_in[4]), .A2(n813), .B1(n862), .B2(\mem[27][4] ), 
        .ZN(n858) );
  INV_X1 U455 ( .A(n857), .ZN(n290) );
  AOI22_X1 U456 ( .A1(data_in[5]), .A2(n813), .B1(n862), .B2(\mem[27][5] ), 
        .ZN(n857) );
  INV_X1 U457 ( .A(n856), .ZN(n289) );
  AOI22_X1 U458 ( .A1(data_in[6]), .A2(n813), .B1(n862), .B2(\mem[27][6] ), 
        .ZN(n856) );
  INV_X1 U459 ( .A(n855), .ZN(n288) );
  AOI22_X1 U460 ( .A1(data_in[7]), .A2(n813), .B1(n862), .B2(\mem[27][7] ), 
        .ZN(n855) );
  INV_X1 U461 ( .A(n854), .ZN(n287) );
  AOI22_X1 U462 ( .A1(data_in[0]), .A2(n812), .B1(n853), .B2(\mem[28][0] ), 
        .ZN(n854) );
  INV_X1 U463 ( .A(n852), .ZN(n286) );
  AOI22_X1 U464 ( .A1(data_in[1]), .A2(n812), .B1(n853), .B2(\mem[28][1] ), 
        .ZN(n852) );
  INV_X1 U465 ( .A(n851), .ZN(n285) );
  AOI22_X1 U466 ( .A1(data_in[2]), .A2(n812), .B1(n853), .B2(\mem[28][2] ), 
        .ZN(n851) );
  INV_X1 U467 ( .A(n850), .ZN(n284) );
  AOI22_X1 U468 ( .A1(data_in[3]), .A2(n812), .B1(n853), .B2(\mem[28][3] ), 
        .ZN(n850) );
  INV_X1 U469 ( .A(n849), .ZN(n283) );
  AOI22_X1 U470 ( .A1(data_in[4]), .A2(n812), .B1(n853), .B2(\mem[28][4] ), 
        .ZN(n849) );
  INV_X1 U471 ( .A(n848), .ZN(n282) );
  AOI22_X1 U472 ( .A1(data_in[5]), .A2(n812), .B1(n853), .B2(\mem[28][5] ), 
        .ZN(n848) );
  INV_X1 U473 ( .A(n847), .ZN(n281) );
  AOI22_X1 U474 ( .A1(data_in[6]), .A2(n812), .B1(n853), .B2(\mem[28][6] ), 
        .ZN(n847) );
  INV_X1 U475 ( .A(n846), .ZN(n280) );
  AOI22_X1 U476 ( .A1(data_in[7]), .A2(n812), .B1(n853), .B2(\mem[28][7] ), 
        .ZN(n846) );
  INV_X1 U477 ( .A(n1145), .ZN(n279) );
  AOI22_X1 U478 ( .A1(n819), .A2(data_in[0]), .B1(n1144), .B2(\mem[29][0] ), 
        .ZN(n1145) );
  INV_X1 U479 ( .A(n1143), .ZN(n278) );
  AOI22_X1 U480 ( .A1(n819), .A2(data_in[1]), .B1(n1144), .B2(\mem[29][1] ), 
        .ZN(n1143) );
  INV_X1 U481 ( .A(n1142), .ZN(n277) );
  AOI22_X1 U482 ( .A1(n819), .A2(data_in[2]), .B1(n1144), .B2(\mem[29][2] ), 
        .ZN(n1142) );
  INV_X1 U483 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U484 ( .A1(n819), .A2(data_in[3]), .B1(n1144), .B2(\mem[29][3] ), 
        .ZN(n1141) );
  INV_X1 U485 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U486 ( .A1(n819), .A2(data_in[4]), .B1(n1144), .B2(\mem[29][4] ), 
        .ZN(n1140) );
  INV_X1 U487 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U488 ( .A1(n819), .A2(data_in[5]), .B1(n1144), .B2(\mem[29][5] ), 
        .ZN(n1139) );
  INV_X1 U489 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U490 ( .A1(n819), .A2(data_in[6]), .B1(n1144), .B2(\mem[29][6] ), 
        .ZN(n1138) );
  INV_X1 U491 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U492 ( .A1(n819), .A2(data_in[7]), .B1(n1144), .B2(\mem[29][7] ), 
        .ZN(n1137) );
  INV_X1 U493 ( .A(n1134), .ZN(n271) );
  AOI22_X1 U494 ( .A1(data_in[0]), .A2(n818), .B1(n1133), .B2(\mem[30][0] ), 
        .ZN(n1134) );
  INV_X1 U495 ( .A(n1132), .ZN(n270) );
  AOI22_X1 U496 ( .A1(data_in[1]), .A2(n818), .B1(n1133), .B2(\mem[30][1] ), 
        .ZN(n1132) );
  INV_X1 U497 ( .A(n1131), .ZN(n269) );
  AOI22_X1 U498 ( .A1(data_in[2]), .A2(n818), .B1(n1133), .B2(\mem[30][2] ), 
        .ZN(n1131) );
  INV_X1 U499 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U500 ( .A1(data_in[3]), .A2(n818), .B1(n1133), .B2(\mem[30][3] ), 
        .ZN(n1130) );
  INV_X1 U501 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U502 ( .A1(data_in[4]), .A2(n818), .B1(n1133), .B2(\mem[30][4] ), 
        .ZN(n1129) );
  INV_X1 U503 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U504 ( .A1(data_in[5]), .A2(n818), .B1(n1133), .B2(\mem[30][5] ), 
        .ZN(n1128) );
  INV_X1 U505 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U506 ( .A1(data_in[6]), .A2(n818), .B1(n1133), .B2(\mem[30][6] ), 
        .ZN(n1127) );
  INV_X1 U507 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U508 ( .A1(data_in[7]), .A2(n818), .B1(n1133), .B2(\mem[30][7] ), 
        .ZN(n1126) );
  INV_X1 U509 ( .A(n1124), .ZN(n263) );
  AOI22_X1 U510 ( .A1(data_in[0]), .A2(n817), .B1(n1123), .B2(\mem[31][0] ), 
        .ZN(n1124) );
  INV_X1 U511 ( .A(n1122), .ZN(n262) );
  AOI22_X1 U512 ( .A1(data_in[1]), .A2(n817), .B1(n1123), .B2(\mem[31][1] ), 
        .ZN(n1122) );
  INV_X1 U513 ( .A(n1121), .ZN(n261) );
  AOI22_X1 U514 ( .A1(data_in[2]), .A2(n817), .B1(n1123), .B2(\mem[31][2] ), 
        .ZN(n1121) );
  INV_X1 U515 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U516 ( .A1(data_in[3]), .A2(n817), .B1(n1123), .B2(\mem[31][3] ), 
        .ZN(n1120) );
  INV_X1 U517 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U518 ( .A1(data_in[4]), .A2(n817), .B1(n1123), .B2(\mem[31][4] ), 
        .ZN(n1119) );
  INV_X1 U519 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U520 ( .A1(data_in[5]), .A2(n817), .B1(n1123), .B2(\mem[31][5] ), 
        .ZN(n1118) );
  INV_X1 U521 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U522 ( .A1(data_in[6]), .A2(n817), .B1(n1123), .B2(\mem[31][6] ), 
        .ZN(n1117) );
  INV_X1 U523 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U524 ( .A1(data_in[7]), .A2(n817), .B1(n1123), .B2(\mem[31][7] ), 
        .ZN(n1116) );
  INV_X1 U525 ( .A(n1114), .ZN(n811) );
  AOI22_X1 U526 ( .A1(data_in[0]), .A2(n843), .B1(n1113), .B2(\mem[0][0] ), 
        .ZN(n1114) );
  INV_X1 U527 ( .A(n1112), .ZN(n810) );
  AOI22_X1 U528 ( .A1(data_in[1]), .A2(n843), .B1(n1113), .B2(\mem[0][1] ), 
        .ZN(n1112) );
  INV_X1 U529 ( .A(n1111), .ZN(n809) );
  AOI22_X1 U530 ( .A1(data_in[2]), .A2(n843), .B1(n1113), .B2(\mem[0][2] ), 
        .ZN(n1111) );
  INV_X1 U531 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U532 ( .A1(data_in[3]), .A2(n843), .B1(n1113), .B2(\mem[0][3] ), 
        .ZN(n1110) );
  INV_X1 U533 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U534 ( .A1(data_in[4]), .A2(n843), .B1(n1113), .B2(\mem[0][4] ), 
        .ZN(n1109) );
  INV_X1 U535 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U536 ( .A1(data_in[5]), .A2(n843), .B1(n1113), .B2(\mem[0][5] ), 
        .ZN(n1108) );
  INV_X1 U537 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U538 ( .A1(data_in[6]), .A2(n843), .B1(n1113), .B2(\mem[0][6] ), 
        .ZN(n1107) );
  INV_X1 U539 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U540 ( .A1(data_in[7]), .A2(n843), .B1(n1113), .B2(\mem[0][7] ), 
        .ZN(n1106) );
  INV_X1 U541 ( .A(n1103), .ZN(n803) );
  AOI22_X1 U542 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[1][0] ), 
        .ZN(n1103) );
  INV_X1 U543 ( .A(n1101), .ZN(n802) );
  AOI22_X1 U544 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[1][1] ), 
        .ZN(n1101) );
  INV_X1 U545 ( .A(n1100), .ZN(n801) );
  AOI22_X1 U546 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[1][2] ), 
        .ZN(n1100) );
  INV_X1 U547 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U548 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[1][3] ), 
        .ZN(n1099) );
  INV_X1 U549 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U550 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[1][4] ), 
        .ZN(n1098) );
  INV_X1 U551 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U552 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[1][5] ), 
        .ZN(n1097) );
  INV_X1 U553 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U554 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[1][6] ), 
        .ZN(n1096) );
  INV_X1 U555 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U556 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[1][7] ), 
        .ZN(n1095) );
  INV_X1 U557 ( .A(n1093), .ZN(n795) );
  AOI22_X1 U558 ( .A1(data_in[0]), .A2(n841), .B1(n1092), .B2(\mem[2][0] ), 
        .ZN(n1093) );
  INV_X1 U559 ( .A(n1091), .ZN(n794) );
  AOI22_X1 U560 ( .A1(data_in[1]), .A2(n841), .B1(n1092), .B2(\mem[2][1] ), 
        .ZN(n1091) );
  INV_X1 U561 ( .A(n1090), .ZN(n793) );
  AOI22_X1 U562 ( .A1(data_in[2]), .A2(n841), .B1(n1092), .B2(\mem[2][2] ), 
        .ZN(n1090) );
  INV_X1 U563 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U564 ( .A1(data_in[3]), .A2(n841), .B1(n1092), .B2(\mem[2][3] ), 
        .ZN(n1089) );
  INV_X1 U565 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U566 ( .A1(data_in[4]), .A2(n841), .B1(n1092), .B2(\mem[2][4] ), 
        .ZN(n1088) );
  INV_X1 U567 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U568 ( .A1(data_in[5]), .A2(n841), .B1(n1092), .B2(\mem[2][5] ), 
        .ZN(n1087) );
  INV_X1 U569 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U570 ( .A1(data_in[6]), .A2(n841), .B1(n1092), .B2(\mem[2][6] ), 
        .ZN(n1086) );
  INV_X1 U571 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U572 ( .A1(data_in[7]), .A2(n841), .B1(n1092), .B2(\mem[2][7] ), 
        .ZN(n1085) );
  INV_X1 U573 ( .A(n1083), .ZN(n787) );
  AOI22_X1 U574 ( .A1(data_in[0]), .A2(n840), .B1(n1082), .B2(\mem[3][0] ), 
        .ZN(n1083) );
  INV_X1 U575 ( .A(n1081), .ZN(n786) );
  AOI22_X1 U576 ( .A1(data_in[1]), .A2(n840), .B1(n1082), .B2(\mem[3][1] ), 
        .ZN(n1081) );
  INV_X1 U577 ( .A(n1080), .ZN(n785) );
  AOI22_X1 U578 ( .A1(data_in[2]), .A2(n840), .B1(n1082), .B2(\mem[3][2] ), 
        .ZN(n1080) );
  INV_X1 U579 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U580 ( .A1(data_in[3]), .A2(n840), .B1(n1082), .B2(\mem[3][3] ), 
        .ZN(n1079) );
  INV_X1 U581 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U582 ( .A1(data_in[4]), .A2(n840), .B1(n1082), .B2(\mem[3][4] ), 
        .ZN(n1078) );
  INV_X1 U583 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U584 ( .A1(data_in[5]), .A2(n840), .B1(n1082), .B2(\mem[3][5] ), 
        .ZN(n1077) );
  INV_X1 U585 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U586 ( .A1(data_in[6]), .A2(n840), .B1(n1082), .B2(\mem[3][6] ), 
        .ZN(n1076) );
  INV_X1 U587 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U588 ( .A1(data_in[7]), .A2(n840), .B1(n1082), .B2(\mem[3][7] ), 
        .ZN(n1075) );
  INV_X1 U589 ( .A(n1073), .ZN(n779) );
  AOI22_X1 U590 ( .A1(data_in[0]), .A2(n839), .B1(n1072), .B2(\mem[4][0] ), 
        .ZN(n1073) );
  INV_X1 U591 ( .A(n1071), .ZN(n778) );
  AOI22_X1 U592 ( .A1(data_in[1]), .A2(n839), .B1(n1072), .B2(\mem[4][1] ), 
        .ZN(n1071) );
  INV_X1 U593 ( .A(n1070), .ZN(n777) );
  AOI22_X1 U594 ( .A1(data_in[2]), .A2(n839), .B1(n1072), .B2(\mem[4][2] ), 
        .ZN(n1070) );
  INV_X1 U595 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U596 ( .A1(data_in[3]), .A2(n839), .B1(n1072), .B2(\mem[4][3] ), 
        .ZN(n1069) );
  INV_X1 U597 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U598 ( .A1(data_in[4]), .A2(n839), .B1(n1072), .B2(\mem[4][4] ), 
        .ZN(n1068) );
  INV_X1 U599 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U600 ( .A1(data_in[5]), .A2(n839), .B1(n1072), .B2(\mem[4][5] ), 
        .ZN(n1067) );
  INV_X1 U601 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U602 ( .A1(data_in[6]), .A2(n839), .B1(n1072), .B2(\mem[4][6] ), 
        .ZN(n1066) );
  INV_X1 U603 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U604 ( .A1(data_in[7]), .A2(n839), .B1(n1072), .B2(\mem[4][7] ), 
        .ZN(n1065) );
  INV_X1 U605 ( .A(N13), .ZN(n844) );
  INV_X1 U606 ( .A(N14), .ZN(n845) );
  MUX2_X1 U607 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n251), .Z(n3) );
  MUX2_X1 U608 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n251), .Z(n4) );
  MUX2_X1 U609 ( .A(n4), .B(n3), .S(n244), .Z(n5) );
  MUX2_X1 U610 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n251), .Z(n6) );
  MUX2_X1 U611 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n251), .Z(n7) );
  MUX2_X1 U612 ( .A(n7), .B(n6), .S(n246), .Z(n8) );
  MUX2_X1 U613 ( .A(n8), .B(n5), .S(n243), .Z(n9) );
  MUX2_X1 U614 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n251), .Z(n10) );
  MUX2_X1 U615 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n251), .Z(n11) );
  MUX2_X1 U616 ( .A(n11), .B(n10), .S(n245), .Z(n12) );
  MUX2_X1 U617 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n251), .Z(n13) );
  MUX2_X1 U618 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n251), .Z(n14) );
  MUX2_X1 U619 ( .A(n14), .B(n13), .S(N11), .Z(n15) );
  MUX2_X1 U620 ( .A(n15), .B(n12), .S(n243), .Z(n16) );
  MUX2_X1 U621 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U622 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n247), .Z(n18) );
  MUX2_X1 U623 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n247), .Z(n19) );
  MUX2_X1 U624 ( .A(n19), .B(n18), .S(n244), .Z(n20) );
  MUX2_X1 U625 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n247), .Z(n21) );
  MUX2_X1 U626 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n247), .Z(n22) );
  MUX2_X1 U627 ( .A(n22), .B(n21), .S(n244), .Z(n23) );
  MUX2_X1 U628 ( .A(n23), .B(n20), .S(n243), .Z(n24) );
  MUX2_X1 U629 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n247), .Z(n25) );
  MUX2_X1 U630 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n247), .Z(n26) );
  MUX2_X1 U631 ( .A(n26), .B(n25), .S(n244), .Z(n27) );
  MUX2_X1 U632 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n247), .Z(n28) );
  MUX2_X1 U633 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n247), .Z(n29) );
  MUX2_X1 U634 ( .A(n29), .B(n28), .S(n244), .Z(n30) );
  MUX2_X1 U635 ( .A(n30), .B(n27), .S(n243), .Z(n31) );
  MUX2_X1 U636 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U637 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U638 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n247), .Z(n33) );
  MUX2_X1 U639 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n247), .Z(n34) );
  MUX2_X1 U640 ( .A(n34), .B(n33), .S(n244), .Z(n35) );
  MUX2_X1 U641 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n247), .Z(n36) );
  MUX2_X1 U642 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n247), .Z(n37) );
  MUX2_X1 U643 ( .A(n37), .B(n36), .S(n244), .Z(n38) );
  MUX2_X1 U644 ( .A(n38), .B(n35), .S(n243), .Z(n39) );
  MUX2_X1 U645 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n248), .Z(n40) );
  MUX2_X1 U646 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n248), .Z(n41) );
  MUX2_X1 U647 ( .A(n41), .B(n40), .S(n244), .Z(n42) );
  MUX2_X1 U648 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n248), .Z(n43) );
  MUX2_X1 U649 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n248), .Z(n44) );
  MUX2_X1 U650 ( .A(n44), .B(n43), .S(n244), .Z(n45) );
  MUX2_X1 U651 ( .A(n45), .B(n42), .S(n243), .Z(n46) );
  MUX2_X1 U652 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U653 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n248), .Z(n48) );
  MUX2_X1 U654 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n248), .Z(n49) );
  MUX2_X1 U655 ( .A(n49), .B(n48), .S(n244), .Z(n50) );
  MUX2_X1 U656 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n248), .Z(n51) );
  MUX2_X1 U657 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n248), .Z(n52) );
  MUX2_X1 U658 ( .A(n52), .B(n51), .S(n244), .Z(n53) );
  MUX2_X1 U659 ( .A(n53), .B(n50), .S(n243), .Z(n54) );
  MUX2_X1 U660 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n248), .Z(n55) );
  MUX2_X1 U661 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n248), .Z(n56) );
  MUX2_X1 U662 ( .A(n56), .B(n55), .S(n244), .Z(n57) );
  MUX2_X1 U663 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n248), .Z(n58) );
  MUX2_X1 U664 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n248), .Z(n59) );
  MUX2_X1 U665 ( .A(n59), .B(n58), .S(n244), .Z(n60) );
  MUX2_X1 U666 ( .A(n60), .B(n57), .S(n243), .Z(n61) );
  MUX2_X1 U667 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U668 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U669 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n250), .Z(n63) );
  MUX2_X1 U670 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n249), .Z(n64) );
  MUX2_X1 U671 ( .A(n64), .B(n63), .S(n245), .Z(n65) );
  MUX2_X1 U672 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n248), .Z(n66) );
  MUX2_X1 U673 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n249), .Z(n67) );
  MUX2_X1 U674 ( .A(n67), .B(n66), .S(n245), .Z(n68) );
  MUX2_X1 U675 ( .A(n68), .B(n65), .S(n243), .Z(n69) );
  MUX2_X1 U676 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n250), .Z(n70) );
  MUX2_X1 U677 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n247), .Z(n71) );
  MUX2_X1 U678 ( .A(n71), .B(n70), .S(n245), .Z(n72) );
  MUX2_X1 U679 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n248), .Z(n73) );
  MUX2_X1 U680 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n249), .Z(n74) );
  MUX2_X1 U681 ( .A(n74), .B(n73), .S(n245), .Z(n75) );
  MUX2_X1 U682 ( .A(n75), .B(n72), .S(N12), .Z(n76) );
  MUX2_X1 U683 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U684 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n247), .Z(n78) );
  MUX2_X1 U685 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n250), .Z(n79) );
  MUX2_X1 U686 ( .A(n79), .B(n78), .S(n245), .Z(n80) );
  MUX2_X1 U687 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n247), .Z(n81) );
  MUX2_X1 U688 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n248), .Z(n82) );
  MUX2_X1 U689 ( .A(n82), .B(n81), .S(n245), .Z(n83) );
  MUX2_X1 U690 ( .A(n83), .B(n80), .S(n243), .Z(n84) );
  MUX2_X1 U691 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n252), .Z(n85) );
  MUX2_X1 U692 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n250), .Z(n86) );
  MUX2_X1 U693 ( .A(n86), .B(n85), .S(n245), .Z(n87) );
  MUX2_X1 U694 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n252), .Z(n88) );
  MUX2_X1 U695 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n248), .Z(n89) );
  MUX2_X1 U696 ( .A(n89), .B(n88), .S(n245), .Z(n90) );
  MUX2_X1 U697 ( .A(n90), .B(n87), .S(N12), .Z(n91) );
  MUX2_X1 U698 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U699 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U700 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n250), .Z(n93) );
  MUX2_X1 U701 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U702 ( .A(n94), .B(n93), .S(n245), .Z(n95) );
  MUX2_X1 U703 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n248), .Z(n96) );
  MUX2_X1 U704 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n252), .Z(n97) );
  MUX2_X1 U705 ( .A(n97), .B(n96), .S(n245), .Z(n98) );
  MUX2_X1 U706 ( .A(n98), .B(n95), .S(n243), .Z(n99) );
  MUX2_X1 U707 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n249), .Z(n100) );
  MUX2_X1 U708 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n252), .Z(n101) );
  MUX2_X1 U709 ( .A(n101), .B(n100), .S(n245), .Z(n102) );
  MUX2_X1 U710 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n252), .Z(n103) );
  MUX2_X1 U711 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n247), .Z(n104) );
  MUX2_X1 U712 ( .A(n104), .B(n103), .S(n245), .Z(n105) );
  MUX2_X1 U713 ( .A(n105), .B(n102), .S(N12), .Z(n106) );
  MUX2_X1 U714 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U715 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n249), .Z(n108) );
  MUX2_X1 U716 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n249), .Z(n109) );
  MUX2_X1 U717 ( .A(n109), .B(n108), .S(n246), .Z(n110) );
  MUX2_X1 U718 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n249), .Z(n111) );
  MUX2_X1 U719 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n249), .Z(n112) );
  MUX2_X1 U720 ( .A(n112), .B(n111), .S(n246), .Z(n113) );
  MUX2_X1 U721 ( .A(n113), .B(n110), .S(n243), .Z(n114) );
  MUX2_X1 U722 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n249), .Z(n115) );
  MUX2_X1 U723 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n249), .Z(n116) );
  MUX2_X1 U724 ( .A(n116), .B(n115), .S(n246), .Z(n117) );
  MUX2_X1 U725 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n249), .Z(n118) );
  MUX2_X1 U726 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n249), .Z(n119) );
  MUX2_X1 U727 ( .A(n119), .B(n118), .S(n246), .Z(n120) );
  MUX2_X1 U728 ( .A(n120), .B(n117), .S(N12), .Z(n121) );
  MUX2_X1 U729 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U730 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U731 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n249), .Z(n123) );
  MUX2_X1 U732 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n249), .Z(n124) );
  MUX2_X1 U733 ( .A(n124), .B(n123), .S(n246), .Z(n125) );
  MUX2_X1 U734 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n249), .Z(n126) );
  MUX2_X1 U735 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n249), .Z(n127) );
  MUX2_X1 U736 ( .A(n127), .B(n126), .S(n246), .Z(n128) );
  MUX2_X1 U737 ( .A(n128), .B(n125), .S(n243), .Z(n129) );
  MUX2_X1 U738 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n250), .Z(n130) );
  MUX2_X1 U739 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n250), .Z(n131) );
  MUX2_X1 U740 ( .A(n131), .B(n130), .S(n246), .Z(n132) );
  MUX2_X1 U741 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n250), .Z(n133) );
  MUX2_X1 U742 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n250), .Z(n134) );
  MUX2_X1 U743 ( .A(n134), .B(n133), .S(n246), .Z(n135) );
  MUX2_X1 U744 ( .A(n135), .B(n132), .S(N12), .Z(n136) );
  MUX2_X1 U745 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U746 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n250), .Z(n138) );
  MUX2_X1 U747 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n250), .Z(n139) );
  MUX2_X1 U748 ( .A(n139), .B(n138), .S(n246), .Z(n140) );
  MUX2_X1 U749 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n250), .Z(n141) );
  MUX2_X1 U750 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n250), .Z(n142) );
  MUX2_X1 U751 ( .A(n142), .B(n141), .S(n246), .Z(n143) );
  MUX2_X1 U752 ( .A(n143), .B(n140), .S(n243), .Z(n144) );
  MUX2_X1 U753 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n250), .Z(n145) );
  MUX2_X1 U754 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n250), .Z(n146) );
  MUX2_X1 U755 ( .A(n146), .B(n145), .S(n246), .Z(n147) );
  MUX2_X1 U756 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n250), .Z(n148) );
  MUX2_X1 U757 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n250), .Z(n149) );
  MUX2_X1 U758 ( .A(n149), .B(n148), .S(n246), .Z(n150) );
  MUX2_X1 U759 ( .A(n150), .B(n147), .S(N12), .Z(n151) );
  MUX2_X1 U760 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U761 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U762 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n251), .Z(n153) );
  MUX2_X1 U763 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n251), .Z(n154) );
  MUX2_X1 U764 ( .A(n154), .B(n153), .S(N11), .Z(n155) );
  MUX2_X1 U765 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n251), .Z(n156) );
  MUX2_X1 U766 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n251), .Z(n157) );
  MUX2_X1 U767 ( .A(n157), .B(n156), .S(N11), .Z(n158) );
  MUX2_X1 U768 ( .A(n158), .B(n155), .S(n243), .Z(n159) );
  MUX2_X1 U769 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n251), .Z(n160) );
  MUX2_X1 U770 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n251), .Z(n161) );
  MUX2_X1 U771 ( .A(n161), .B(n160), .S(N11), .Z(n162) );
  MUX2_X1 U772 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n251), .Z(n163) );
  MUX2_X1 U773 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n251), .Z(n164) );
  MUX2_X1 U774 ( .A(n164), .B(n163), .S(N11), .Z(n165) );
  MUX2_X1 U775 ( .A(n165), .B(n162), .S(n243), .Z(n166) );
  MUX2_X1 U776 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U777 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n251), .Z(n168) );
  MUX2_X1 U778 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n251), .Z(n169) );
  MUX2_X1 U779 ( .A(n169), .B(n168), .S(N11), .Z(n170) );
  MUX2_X1 U780 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n251), .Z(n171) );
  MUX2_X1 U781 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n251), .Z(n172) );
  MUX2_X1 U782 ( .A(n172), .B(n171), .S(N11), .Z(n173) );
  MUX2_X1 U783 ( .A(n173), .B(n170), .S(n243), .Z(n174) );
  MUX2_X1 U784 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n252), .Z(n175) );
  MUX2_X1 U785 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n252), .Z(n176) );
  MUX2_X1 U786 ( .A(n176), .B(n175), .S(N11), .Z(n177) );
  MUX2_X1 U787 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n247), .Z(n178) );
  MUX2_X1 U788 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n249), .Z(n179) );
  MUX2_X1 U789 ( .A(n179), .B(n178), .S(N11), .Z(n180) );
  MUX2_X1 U790 ( .A(n180), .B(n177), .S(n243), .Z(n181) );
  MUX2_X1 U791 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U792 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U793 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n252), .Z(n183) );
  MUX2_X1 U794 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n252), .Z(n184) );
  MUX2_X1 U795 ( .A(n184), .B(n183), .S(N11), .Z(n185) );
  MUX2_X1 U796 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n248), .Z(n186) );
  MUX2_X1 U797 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n252), .Z(n187) );
  MUX2_X1 U798 ( .A(n187), .B(n186), .S(n246), .Z(n188) );
  MUX2_X1 U799 ( .A(n188), .B(n185), .S(n243), .Z(n189) );
  MUX2_X1 U800 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n252), .Z(n190) );
  MUX2_X1 U801 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n252), .Z(n191) );
  MUX2_X1 U802 ( .A(n191), .B(n190), .S(n245), .Z(n192) );
  MUX2_X1 U803 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n252), .Z(n193) );
  MUX2_X1 U804 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n252), .Z(n194) );
  MUX2_X1 U805 ( .A(n194), .B(n193), .S(n246), .Z(n195) );
  MUX2_X1 U806 ( .A(n195), .B(n192), .S(N12), .Z(n196) );
  MUX2_X1 U807 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U808 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n252), .Z(n198) );
  MUX2_X1 U809 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(N10), .Z(n199) );
  MUX2_X1 U810 ( .A(n199), .B(n198), .S(n244), .Z(n200) );
  MUX2_X1 U811 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(N10), .Z(n201) );
  MUX2_X1 U812 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n252), .Z(n202) );
  MUX2_X1 U813 ( .A(n202), .B(n201), .S(n246), .Z(n203) );
  MUX2_X1 U814 ( .A(n203), .B(n200), .S(N12), .Z(n204) );
  MUX2_X1 U815 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n205) );
  MUX2_X1 U816 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n252), .Z(n206) );
  MUX2_X1 U817 ( .A(n206), .B(n205), .S(n244), .Z(n207) );
  MUX2_X1 U818 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n208) );
  MUX2_X1 U819 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n252), .Z(n209) );
  MUX2_X1 U820 ( .A(n209), .B(n208), .S(N11), .Z(n210) );
  MUX2_X1 U821 ( .A(n210), .B(n207), .S(N12), .Z(n211) );
  MUX2_X1 U822 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U823 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U824 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n249), .Z(n213) );
  MUX2_X1 U825 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(N10), .Z(n214) );
  MUX2_X1 U826 ( .A(n214), .B(n213), .S(n244), .Z(n215) );
  MUX2_X1 U827 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(N10), .Z(n216) );
  MUX2_X1 U828 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(N10), .Z(n217) );
  MUX2_X1 U829 ( .A(n217), .B(n216), .S(n244), .Z(n218) );
  MUX2_X1 U830 ( .A(n218), .B(n215), .S(n243), .Z(n219) );
  MUX2_X1 U831 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n251), .Z(n220) );
  MUX2_X1 U832 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(N10), .Z(n221) );
  MUX2_X1 U833 ( .A(n221), .B(n220), .S(n246), .Z(n222) );
  MUX2_X1 U834 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n252), .Z(n223) );
  MUX2_X1 U835 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n224) );
  MUX2_X1 U836 ( .A(n224), .B(n223), .S(N11), .Z(n225) );
  MUX2_X1 U837 ( .A(n225), .B(n222), .S(n243), .Z(n226) );
  MUX2_X1 U838 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U839 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n251), .Z(n228) );
  MUX2_X1 U840 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n252), .Z(n229) );
  MUX2_X1 U841 ( .A(n229), .B(n228), .S(n245), .Z(n230) );
  MUX2_X1 U842 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n251), .Z(n231) );
  MUX2_X1 U843 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n232) );
  MUX2_X1 U844 ( .A(n232), .B(n231), .S(n245), .Z(n233) );
  MUX2_X1 U845 ( .A(n233), .B(n230), .S(n243), .Z(n234) );
  MUX2_X1 U846 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n235) );
  MUX2_X1 U847 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n236) );
  MUX2_X1 U848 ( .A(n236), .B(n235), .S(n245), .Z(n237) );
  MUX2_X1 U849 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n238) );
  MUX2_X1 U850 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n239) );
  MUX2_X1 U851 ( .A(n239), .B(n238), .S(N11), .Z(n240) );
  MUX2_X1 U852 ( .A(n240), .B(n237), .S(n243), .Z(n241) );
  MUX2_X1 U853 ( .A(n241), .B(n234), .S(N13), .Z(n242) );
  MUX2_X1 U854 ( .A(n242), .B(n227), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_18 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n256), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n257), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n258), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n259), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n260), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n261), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n262), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n263), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n264), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n265), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n266), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n267), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n268), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n269), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n270), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n271), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n272), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n273), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n274), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n275), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n276), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n277), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n278), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n279), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n280), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n281), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n282), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n283), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n284), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n285), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n286), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n287), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n288), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n289), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n290), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n291), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n292), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n293), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n594), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n595), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n596), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n597), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n598), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n599), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n600), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n601), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n602), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n603), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n604), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n605), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n606), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n607), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n608), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n609), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n610), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n611), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n612), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n613), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n614), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n615), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n616), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n617), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n618), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n619), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n620), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n621), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n622), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n623), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n624), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n625), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n626), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n627), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n628), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n629), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n630), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n631), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n632), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n633), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n634), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n635), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n636), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n637), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n638), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n639), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n640), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n641), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n642), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n643), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n644), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n645), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n646), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n647), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n648), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n649), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n650), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n651), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n652), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n653), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n654), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n655), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n656), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n657), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n658), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n659), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n660), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n661), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n662), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n663), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n664), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n665), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n666), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n667), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n668), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n669), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n670), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n671), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n672), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n673), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n674), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n675), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n676), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n677), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n678), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n679), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n680), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n681), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n682), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n683), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n684), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n685), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n686), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n687), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n688), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n689), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n690), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n691), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n692), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n693), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n694), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n695), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n696), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n697), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n698), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n699), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n700), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n701), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n702), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n703), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n704), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n705), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n706), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n707), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n708), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n709), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n710), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n711), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n712), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n713), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n714), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n715), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n716), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n717), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n718), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n719), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n720), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n721), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n722), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n723), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n724), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n725), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n726), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n727), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n728), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n729), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n730), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n731), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n732), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n733), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n734), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n735), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n736), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n737), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n738), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n739), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n740), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n741), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n742), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n743), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n744), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n745), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n746), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n747), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n748), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n749), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n750), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n751), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n752), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n753), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n754), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n755), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n756), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n757), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n758), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n759), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n760), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n761), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n762), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n763), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n764), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n765), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n766), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n767), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n768), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n769), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n770), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n771), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n772), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n773), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n774), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n775), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n776), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n777), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n778), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n779), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n780), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n781), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n782), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n783), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n784), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n785), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n786), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n787), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n788), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n789), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n790), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n791), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n792), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n793), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n794), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n795), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n796), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n797), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n798), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n799), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n800), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n801), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n802), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n803), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n804), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n805), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n806), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n807), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n808), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n809), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n810), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n811), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .QN(n1) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[1]) );
  BUF_X1 U4 ( .A(N10), .Z(n251) );
  BUF_X1 U5 ( .A(n252), .Z(n248) );
  BUF_X1 U6 ( .A(n252), .Z(n247) );
  BUF_X1 U7 ( .A(n252), .Z(n249) );
  BUF_X1 U8 ( .A(n252), .Z(n250) );
  BUF_X1 U9 ( .A(N10), .Z(n252) );
  INV_X1 U10 ( .A(n1113), .ZN(n843) );
  INV_X1 U11 ( .A(n1102), .ZN(n842) );
  INV_X1 U12 ( .A(n1092), .ZN(n841) );
  INV_X1 U13 ( .A(n1082), .ZN(n840) );
  INV_X1 U14 ( .A(n1072), .ZN(n839) );
  INV_X1 U15 ( .A(n1062), .ZN(n838) );
  INV_X1 U16 ( .A(n1053), .ZN(n837) );
  INV_X1 U17 ( .A(n1044), .ZN(n836) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1105) );
  NOR3_X1 U19 ( .A1(N11), .A2(N12), .A3(n253), .ZN(n1094) );
  NAND2_X1 U20 ( .A1(n1104), .A2(n1136), .ZN(n1062) );
  NAND2_X1 U21 ( .A1(n1105), .A2(n1104), .ZN(n1113) );
  NAND2_X1 U22 ( .A1(n1094), .A2(n1104), .ZN(n1102) );
  NAND2_X1 U23 ( .A1(n1084), .A2(n1104), .ZN(n1092) );
  NAND2_X1 U24 ( .A1(n1074), .A2(n1104), .ZN(n1082) );
  NAND2_X1 U25 ( .A1(n1064), .A2(n1104), .ZN(n1072) );
  NAND2_X1 U26 ( .A1(n1104), .A2(n1125), .ZN(n1053) );
  NAND2_X1 U27 ( .A1(n1104), .A2(n1115), .ZN(n1044) );
  INV_X1 U28 ( .A(n1133), .ZN(n818) );
  INV_X1 U29 ( .A(n1123), .ZN(n817) );
  INV_X1 U30 ( .A(n889), .ZN(n816) );
  INV_X1 U31 ( .A(n880), .ZN(n815) );
  INV_X1 U32 ( .A(n871), .ZN(n814) );
  INV_X1 U33 ( .A(n862), .ZN(n813) );
  INV_X1 U34 ( .A(n853), .ZN(n812) );
  INV_X1 U35 ( .A(n989), .ZN(n830) );
  INV_X1 U36 ( .A(n980), .ZN(n829) );
  INV_X1 U37 ( .A(n971), .ZN(n828) );
  INV_X1 U38 ( .A(n916), .ZN(n822) );
  INV_X1 U39 ( .A(n907), .ZN(n821) );
  INV_X1 U40 ( .A(n898), .ZN(n820) );
  INV_X1 U41 ( .A(n1035), .ZN(n835) );
  INV_X1 U42 ( .A(n1025), .ZN(n834) );
  INV_X1 U43 ( .A(n1016), .ZN(n833) );
  INV_X1 U44 ( .A(n1007), .ZN(n832) );
  INV_X1 U45 ( .A(n998), .ZN(n831) );
  INV_X1 U46 ( .A(n962), .ZN(n827) );
  INV_X1 U47 ( .A(n952), .ZN(n826) );
  INV_X1 U48 ( .A(n943), .ZN(n825) );
  INV_X1 U49 ( .A(n934), .ZN(n824) );
  INV_X1 U50 ( .A(n925), .ZN(n823) );
  INV_X1 U51 ( .A(n1144), .ZN(n819) );
  BUF_X1 U52 ( .A(N11), .Z(n245) );
  BUF_X1 U53 ( .A(N11), .Z(n246) );
  INV_X1 U54 ( .A(N10), .ZN(n253) );
  BUF_X1 U55 ( .A(N12), .Z(n243) );
  NOR3_X1 U56 ( .A1(n255), .A2(N10), .A3(n254), .ZN(n1125) );
  NOR3_X1 U57 ( .A1(n255), .A2(n253), .A3(n254), .ZN(n1115) );
  NOR3_X1 U58 ( .A1(n253), .A2(N11), .A3(n255), .ZN(n1136) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n254), .ZN(n1084) );
  NOR3_X1 U60 ( .A1(n253), .A2(N12), .A3(n254), .ZN(n1074) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n255), .ZN(n1064) );
  NAND2_X1 U62 ( .A1(n1027), .A2(n1136), .ZN(n989) );
  NAND2_X1 U63 ( .A1(n954), .A2(n1136), .ZN(n916) );
  NAND2_X1 U64 ( .A1(n1027), .A2(n1064), .ZN(n998) );
  NAND2_X1 U65 ( .A1(n954), .A2(n1064), .ZN(n925) );
  NAND2_X1 U66 ( .A1(n1027), .A2(n1105), .ZN(n1035) );
  NAND2_X1 U67 ( .A1(n1027), .A2(n1094), .ZN(n1025) );
  NAND2_X1 U68 ( .A1(n954), .A2(n1105), .ZN(n962) );
  NAND2_X1 U69 ( .A1(n954), .A2(n1094), .ZN(n952) );
  NAND2_X1 U70 ( .A1(n1105), .A2(n1135), .ZN(n889) );
  NAND2_X1 U71 ( .A1(n1094), .A2(n1135), .ZN(n880) );
  NAND2_X1 U72 ( .A1(n1084), .A2(n1135), .ZN(n871) );
  NAND2_X1 U73 ( .A1(n1074), .A2(n1135), .ZN(n862) );
  NAND2_X1 U74 ( .A1(n1064), .A2(n1135), .ZN(n853) );
  NAND2_X1 U75 ( .A1(n1136), .A2(n1135), .ZN(n1144) );
  NAND2_X1 U76 ( .A1(n1125), .A2(n1135), .ZN(n1133) );
  NAND2_X1 U77 ( .A1(n1115), .A2(n1135), .ZN(n1123) );
  NAND2_X1 U78 ( .A1(n1027), .A2(n1084), .ZN(n1016) );
  NAND2_X1 U79 ( .A1(n1027), .A2(n1074), .ZN(n1007) );
  NAND2_X1 U80 ( .A1(n954), .A2(n1084), .ZN(n943) );
  NAND2_X1 U81 ( .A1(n954), .A2(n1074), .ZN(n934) );
  NAND2_X1 U82 ( .A1(n1027), .A2(n1125), .ZN(n980) );
  NAND2_X1 U83 ( .A1(n954), .A2(n1125), .ZN(n907) );
  NAND2_X1 U84 ( .A1(n1027), .A2(n1115), .ZN(n971) );
  NAND2_X1 U85 ( .A1(n954), .A2(n1115), .ZN(n898) );
  AND3_X1 U86 ( .A1(n844), .A2(n845), .A3(wr_en), .ZN(n1104) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1135) );
  AND3_X1 U88 ( .A1(N13), .A2(n845), .A3(wr_en), .ZN(n1027) );
  AND3_X1 U89 ( .A1(N14), .A2(n844), .A3(wr_en), .ZN(n954) );
  INV_X1 U90 ( .A(n984), .ZN(n702) );
  AOI22_X1 U91 ( .A1(data_in[5]), .A2(n830), .B1(n989), .B2(\mem[13][5] ), 
        .ZN(n984) );
  INV_X1 U92 ( .A(n983), .ZN(n701) );
  AOI22_X1 U93 ( .A1(data_in[6]), .A2(n830), .B1(n989), .B2(\mem[13][6] ), 
        .ZN(n983) );
  INV_X1 U94 ( .A(n982), .ZN(n700) );
  AOI22_X1 U95 ( .A1(data_in[7]), .A2(n830), .B1(n989), .B2(\mem[13][7] ), 
        .ZN(n982) );
  INV_X1 U96 ( .A(n1063), .ZN(n771) );
  AOI22_X1 U97 ( .A1(data_in[0]), .A2(n838), .B1(n1062), .B2(\mem[5][0] ), 
        .ZN(n1063) );
  INV_X1 U98 ( .A(n1061), .ZN(n770) );
  AOI22_X1 U99 ( .A1(data_in[1]), .A2(n838), .B1(n1062), .B2(\mem[5][1] ), 
        .ZN(n1061) );
  INV_X1 U100 ( .A(n1060), .ZN(n769) );
  AOI22_X1 U101 ( .A1(data_in[2]), .A2(n838), .B1(n1062), .B2(\mem[5][2] ), 
        .ZN(n1060) );
  INV_X1 U102 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U103 ( .A1(data_in[3]), .A2(n838), .B1(n1062), .B2(\mem[5][3] ), 
        .ZN(n1059) );
  INV_X1 U104 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U105 ( .A1(data_in[4]), .A2(n838), .B1(n1062), .B2(\mem[5][4] ), 
        .ZN(n1058) );
  INV_X1 U106 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U107 ( .A1(data_in[5]), .A2(n838), .B1(n1062), .B2(\mem[5][5] ), 
        .ZN(n1057) );
  INV_X1 U108 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U109 ( .A1(data_in[6]), .A2(n838), .B1(n1062), .B2(\mem[5][6] ), 
        .ZN(n1056) );
  INV_X1 U110 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U111 ( .A1(data_in[7]), .A2(n838), .B1(n1062), .B2(\mem[5][7] ), 
        .ZN(n1055) );
  INV_X1 U112 ( .A(n1026), .ZN(n739) );
  AOI22_X1 U113 ( .A1(data_in[0]), .A2(n834), .B1(n1025), .B2(\mem[9][0] ), 
        .ZN(n1026) );
  INV_X1 U114 ( .A(n1024), .ZN(n738) );
  AOI22_X1 U115 ( .A1(data_in[1]), .A2(n834), .B1(n1025), .B2(\mem[9][1] ), 
        .ZN(n1024) );
  INV_X1 U116 ( .A(n1023), .ZN(n737) );
  AOI22_X1 U117 ( .A1(data_in[2]), .A2(n834), .B1(n1025), .B2(\mem[9][2] ), 
        .ZN(n1023) );
  INV_X1 U118 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U119 ( .A1(data_in[3]), .A2(n834), .B1(n1025), .B2(\mem[9][3] ), 
        .ZN(n1022) );
  INV_X1 U120 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U121 ( .A1(data_in[4]), .A2(n834), .B1(n1025), .B2(\mem[9][4] ), 
        .ZN(n1021) );
  INV_X1 U122 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U123 ( .A1(data_in[5]), .A2(n834), .B1(n1025), .B2(\mem[9][5] ), 
        .ZN(n1020) );
  INV_X1 U124 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U125 ( .A1(data_in[6]), .A2(n834), .B1(n1025), .B2(\mem[9][6] ), 
        .ZN(n1019) );
  INV_X1 U126 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U127 ( .A1(data_in[7]), .A2(n834), .B1(n1025), .B2(\mem[9][7] ), 
        .ZN(n1018) );
  INV_X1 U128 ( .A(n990), .ZN(n707) );
  AOI22_X1 U129 ( .A1(data_in[0]), .A2(n830), .B1(n989), .B2(\mem[13][0] ), 
        .ZN(n990) );
  INV_X1 U130 ( .A(n988), .ZN(n706) );
  AOI22_X1 U131 ( .A1(data_in[1]), .A2(n830), .B1(n989), .B2(\mem[13][1] ), 
        .ZN(n988) );
  INV_X1 U132 ( .A(n987), .ZN(n705) );
  AOI22_X1 U133 ( .A1(data_in[2]), .A2(n830), .B1(n989), .B2(\mem[13][2] ), 
        .ZN(n987) );
  INV_X1 U134 ( .A(n986), .ZN(n704) );
  AOI22_X1 U135 ( .A1(data_in[3]), .A2(n830), .B1(n989), .B2(\mem[13][3] ), 
        .ZN(n986) );
  INV_X1 U136 ( .A(n985), .ZN(n703) );
  AOI22_X1 U137 ( .A1(data_in[4]), .A2(n830), .B1(n989), .B2(\mem[13][4] ), 
        .ZN(n985) );
  INV_X1 U138 ( .A(n953), .ZN(n675) );
  AOI22_X1 U139 ( .A1(data_in[0]), .A2(n826), .B1(n952), .B2(\mem[17][0] ), 
        .ZN(n953) );
  INV_X1 U140 ( .A(n951), .ZN(n674) );
  AOI22_X1 U141 ( .A1(data_in[1]), .A2(n826), .B1(n952), .B2(\mem[17][1] ), 
        .ZN(n951) );
  INV_X1 U142 ( .A(n950), .ZN(n673) );
  AOI22_X1 U143 ( .A1(data_in[2]), .A2(n826), .B1(n952), .B2(\mem[17][2] ), 
        .ZN(n950) );
  INV_X1 U144 ( .A(n949), .ZN(n672) );
  AOI22_X1 U145 ( .A1(data_in[3]), .A2(n826), .B1(n952), .B2(\mem[17][3] ), 
        .ZN(n949) );
  INV_X1 U146 ( .A(n948), .ZN(n671) );
  AOI22_X1 U147 ( .A1(data_in[4]), .A2(n826), .B1(n952), .B2(\mem[17][4] ), 
        .ZN(n948) );
  INV_X1 U148 ( .A(n947), .ZN(n670) );
  AOI22_X1 U149 ( .A1(data_in[5]), .A2(n826), .B1(n952), .B2(\mem[17][5] ), 
        .ZN(n947) );
  INV_X1 U150 ( .A(n946), .ZN(n669) );
  AOI22_X1 U151 ( .A1(data_in[6]), .A2(n826), .B1(n952), .B2(\mem[17][6] ), 
        .ZN(n946) );
  INV_X1 U152 ( .A(n945), .ZN(n668) );
  AOI22_X1 U153 ( .A1(data_in[7]), .A2(n826), .B1(n952), .B2(\mem[17][7] ), 
        .ZN(n945) );
  INV_X1 U154 ( .A(n917), .ZN(n643) );
  AOI22_X1 U155 ( .A1(data_in[0]), .A2(n822), .B1(n916), .B2(\mem[21][0] ), 
        .ZN(n917) );
  INV_X1 U156 ( .A(n915), .ZN(n642) );
  AOI22_X1 U157 ( .A1(data_in[1]), .A2(n822), .B1(n916), .B2(\mem[21][1] ), 
        .ZN(n915) );
  INV_X1 U158 ( .A(n914), .ZN(n641) );
  AOI22_X1 U159 ( .A1(data_in[2]), .A2(n822), .B1(n916), .B2(\mem[21][2] ), 
        .ZN(n914) );
  INV_X1 U160 ( .A(n913), .ZN(n640) );
  AOI22_X1 U161 ( .A1(data_in[3]), .A2(n822), .B1(n916), .B2(\mem[21][3] ), 
        .ZN(n913) );
  INV_X1 U162 ( .A(n912), .ZN(n639) );
  AOI22_X1 U163 ( .A1(data_in[4]), .A2(n822), .B1(n916), .B2(\mem[21][4] ), 
        .ZN(n912) );
  INV_X1 U164 ( .A(n911), .ZN(n638) );
  AOI22_X1 U165 ( .A1(data_in[5]), .A2(n822), .B1(n916), .B2(\mem[21][5] ), 
        .ZN(n911) );
  INV_X1 U166 ( .A(n910), .ZN(n637) );
  AOI22_X1 U167 ( .A1(data_in[6]), .A2(n822), .B1(n916), .B2(\mem[21][6] ), 
        .ZN(n910) );
  INV_X1 U168 ( .A(n909), .ZN(n636) );
  AOI22_X1 U169 ( .A1(data_in[7]), .A2(n822), .B1(n916), .B2(\mem[21][7] ), 
        .ZN(n909) );
  INV_X1 U170 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U171 ( .A1(data_in[0]), .A2(n837), .B1(n1053), .B2(\mem[6][0] ), 
        .ZN(n1054) );
  INV_X1 U172 ( .A(n1052), .ZN(n762) );
  AOI22_X1 U173 ( .A1(data_in[1]), .A2(n837), .B1(n1053), .B2(\mem[6][1] ), 
        .ZN(n1052) );
  INV_X1 U174 ( .A(n1051), .ZN(n761) );
  AOI22_X1 U175 ( .A1(data_in[2]), .A2(n837), .B1(n1053), .B2(\mem[6][2] ), 
        .ZN(n1051) );
  INV_X1 U176 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U177 ( .A1(data_in[3]), .A2(n837), .B1(n1053), .B2(\mem[6][3] ), 
        .ZN(n1050) );
  INV_X1 U178 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U179 ( .A1(data_in[4]), .A2(n837), .B1(n1053), .B2(\mem[6][4] ), 
        .ZN(n1049) );
  INV_X1 U180 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U181 ( .A1(data_in[5]), .A2(n837), .B1(n1053), .B2(\mem[6][5] ), 
        .ZN(n1048) );
  INV_X1 U182 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U183 ( .A1(data_in[6]), .A2(n837), .B1(n1053), .B2(\mem[6][6] ), 
        .ZN(n1047) );
  INV_X1 U184 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U185 ( .A1(data_in[7]), .A2(n837), .B1(n1053), .B2(\mem[6][7] ), 
        .ZN(n1046) );
  INV_X1 U186 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U187 ( .A1(data_in[0]), .A2(n836), .B1(n1044), .B2(\mem[7][0] ), 
        .ZN(n1045) );
  INV_X1 U188 ( .A(n1043), .ZN(n754) );
  AOI22_X1 U189 ( .A1(data_in[1]), .A2(n836), .B1(n1044), .B2(\mem[7][1] ), 
        .ZN(n1043) );
  INV_X1 U190 ( .A(n1042), .ZN(n753) );
  AOI22_X1 U191 ( .A1(data_in[2]), .A2(n836), .B1(n1044), .B2(\mem[7][2] ), 
        .ZN(n1042) );
  INV_X1 U192 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U193 ( .A1(data_in[3]), .A2(n836), .B1(n1044), .B2(\mem[7][3] ), 
        .ZN(n1041) );
  INV_X1 U194 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U195 ( .A1(data_in[4]), .A2(n836), .B1(n1044), .B2(\mem[7][4] ), 
        .ZN(n1040) );
  INV_X1 U196 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U197 ( .A1(data_in[5]), .A2(n836), .B1(n1044), .B2(\mem[7][5] ), 
        .ZN(n1039) );
  INV_X1 U198 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U199 ( .A1(data_in[6]), .A2(n836), .B1(n1044), .B2(\mem[7][6] ), 
        .ZN(n1038) );
  INV_X1 U200 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U201 ( .A1(data_in[7]), .A2(n836), .B1(n1044), .B2(\mem[7][7] ), 
        .ZN(n1037) );
  INV_X1 U202 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U203 ( .A1(data_in[0]), .A2(n833), .B1(n1016), .B2(\mem[10][0] ), 
        .ZN(n1017) );
  INV_X1 U204 ( .A(n1015), .ZN(n730) );
  AOI22_X1 U205 ( .A1(data_in[1]), .A2(n833), .B1(n1016), .B2(\mem[10][1] ), 
        .ZN(n1015) );
  INV_X1 U206 ( .A(n1014), .ZN(n729) );
  AOI22_X1 U207 ( .A1(data_in[2]), .A2(n833), .B1(n1016), .B2(\mem[10][2] ), 
        .ZN(n1014) );
  INV_X1 U208 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U209 ( .A1(data_in[3]), .A2(n833), .B1(n1016), .B2(\mem[10][3] ), 
        .ZN(n1013) );
  INV_X1 U210 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U211 ( .A1(data_in[4]), .A2(n833), .B1(n1016), .B2(\mem[10][4] ), 
        .ZN(n1012) );
  INV_X1 U212 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U213 ( .A1(data_in[5]), .A2(n833), .B1(n1016), .B2(\mem[10][5] ), 
        .ZN(n1011) );
  INV_X1 U214 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U215 ( .A1(data_in[6]), .A2(n833), .B1(n1016), .B2(\mem[10][6] ), 
        .ZN(n1010) );
  INV_X1 U216 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U217 ( .A1(data_in[7]), .A2(n833), .B1(n1016), .B2(\mem[10][7] ), 
        .ZN(n1009) );
  INV_X1 U218 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U219 ( .A1(data_in[0]), .A2(n832), .B1(n1007), .B2(\mem[11][0] ), 
        .ZN(n1008) );
  INV_X1 U220 ( .A(n1006), .ZN(n722) );
  AOI22_X1 U221 ( .A1(data_in[1]), .A2(n832), .B1(n1007), .B2(\mem[11][1] ), 
        .ZN(n1006) );
  INV_X1 U222 ( .A(n1005), .ZN(n721) );
  AOI22_X1 U223 ( .A1(data_in[2]), .A2(n832), .B1(n1007), .B2(\mem[11][2] ), 
        .ZN(n1005) );
  INV_X1 U224 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U225 ( .A1(data_in[3]), .A2(n832), .B1(n1007), .B2(\mem[11][3] ), 
        .ZN(n1004) );
  INV_X1 U226 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U227 ( .A1(data_in[4]), .A2(n832), .B1(n1007), .B2(\mem[11][4] ), 
        .ZN(n1003) );
  INV_X1 U228 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U229 ( .A1(data_in[5]), .A2(n832), .B1(n1007), .B2(\mem[11][5] ), 
        .ZN(n1002) );
  INV_X1 U230 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U231 ( .A1(data_in[6]), .A2(n832), .B1(n1007), .B2(\mem[11][6] ), 
        .ZN(n1001) );
  INV_X1 U232 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U233 ( .A1(data_in[7]), .A2(n832), .B1(n1007), .B2(\mem[11][7] ), 
        .ZN(n1000) );
  INV_X1 U234 ( .A(n981), .ZN(n699) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n829), .B1(n980), .B2(\mem[14][0] ), 
        .ZN(n981) );
  INV_X1 U236 ( .A(n979), .ZN(n698) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n829), .B1(n980), .B2(\mem[14][1] ), 
        .ZN(n979) );
  INV_X1 U238 ( .A(n978), .ZN(n697) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n829), .B1(n980), .B2(\mem[14][2] ), 
        .ZN(n978) );
  INV_X1 U240 ( .A(n977), .ZN(n696) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n829), .B1(n980), .B2(\mem[14][3] ), 
        .ZN(n977) );
  INV_X1 U242 ( .A(n976), .ZN(n695) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n829), .B1(n980), .B2(\mem[14][4] ), 
        .ZN(n976) );
  INV_X1 U244 ( .A(n975), .ZN(n694) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n829), .B1(n980), .B2(\mem[14][5] ), 
        .ZN(n975) );
  INV_X1 U246 ( .A(n974), .ZN(n693) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n829), .B1(n980), .B2(\mem[14][6] ), 
        .ZN(n974) );
  INV_X1 U248 ( .A(n973), .ZN(n692) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n829), .B1(n980), .B2(\mem[14][7] ), 
        .ZN(n973) );
  INV_X1 U250 ( .A(n972), .ZN(n691) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n828), .B1(n971), .B2(\mem[15][0] ), 
        .ZN(n972) );
  INV_X1 U252 ( .A(n970), .ZN(n690) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n828), .B1(n971), .B2(\mem[15][1] ), 
        .ZN(n970) );
  INV_X1 U254 ( .A(n969), .ZN(n689) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n828), .B1(n971), .B2(\mem[15][2] ), 
        .ZN(n969) );
  INV_X1 U256 ( .A(n968), .ZN(n688) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n828), .B1(n971), .B2(\mem[15][3] ), 
        .ZN(n968) );
  INV_X1 U258 ( .A(n967), .ZN(n687) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n828), .B1(n971), .B2(\mem[15][4] ), 
        .ZN(n967) );
  INV_X1 U260 ( .A(n966), .ZN(n686) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n828), .B1(n971), .B2(\mem[15][5] ), 
        .ZN(n966) );
  INV_X1 U262 ( .A(n965), .ZN(n685) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n828), .B1(n971), .B2(\mem[15][6] ), 
        .ZN(n965) );
  INV_X1 U264 ( .A(n964), .ZN(n684) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n828), .B1(n971), .B2(\mem[15][7] ), 
        .ZN(n964) );
  INV_X1 U266 ( .A(n944), .ZN(n667) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n825), .B1(n943), .B2(\mem[18][0] ), 
        .ZN(n944) );
  INV_X1 U268 ( .A(n942), .ZN(n666) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n825), .B1(n943), .B2(\mem[18][1] ), 
        .ZN(n942) );
  INV_X1 U270 ( .A(n941), .ZN(n665) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n825), .B1(n943), .B2(\mem[18][2] ), 
        .ZN(n941) );
  INV_X1 U272 ( .A(n940), .ZN(n664) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n825), .B1(n943), .B2(\mem[18][3] ), 
        .ZN(n940) );
  INV_X1 U274 ( .A(n939), .ZN(n663) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n825), .B1(n943), .B2(\mem[18][4] ), 
        .ZN(n939) );
  INV_X1 U276 ( .A(n938), .ZN(n662) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n825), .B1(n943), .B2(\mem[18][5] ), 
        .ZN(n938) );
  INV_X1 U278 ( .A(n937), .ZN(n661) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n825), .B1(n943), .B2(\mem[18][6] ), 
        .ZN(n937) );
  INV_X1 U280 ( .A(n936), .ZN(n660) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n825), .B1(n943), .B2(\mem[18][7] ), 
        .ZN(n936) );
  INV_X1 U282 ( .A(n935), .ZN(n659) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n824), .B1(n934), .B2(\mem[19][0] ), 
        .ZN(n935) );
  INV_X1 U284 ( .A(n933), .ZN(n658) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n824), .B1(n934), .B2(\mem[19][1] ), 
        .ZN(n933) );
  INV_X1 U286 ( .A(n932), .ZN(n657) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n824), .B1(n934), .B2(\mem[19][2] ), 
        .ZN(n932) );
  INV_X1 U288 ( .A(n931), .ZN(n656) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n824), .B1(n934), .B2(\mem[19][3] ), 
        .ZN(n931) );
  INV_X1 U290 ( .A(n930), .ZN(n655) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n824), .B1(n934), .B2(\mem[19][4] ), 
        .ZN(n930) );
  INV_X1 U292 ( .A(n929), .ZN(n654) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n824), .B1(n934), .B2(\mem[19][5] ), 
        .ZN(n929) );
  INV_X1 U294 ( .A(n928), .ZN(n653) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n824), .B1(n934), .B2(\mem[19][6] ), 
        .ZN(n928) );
  INV_X1 U296 ( .A(n927), .ZN(n652) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n824), .B1(n934), .B2(\mem[19][7] ), 
        .ZN(n927) );
  INV_X1 U298 ( .A(n908), .ZN(n635) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n821), .B1(n907), .B2(\mem[22][0] ), 
        .ZN(n908) );
  INV_X1 U300 ( .A(n906), .ZN(n634) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n821), .B1(n907), .B2(\mem[22][1] ), 
        .ZN(n906) );
  INV_X1 U302 ( .A(n905), .ZN(n633) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n821), .B1(n907), .B2(\mem[22][2] ), 
        .ZN(n905) );
  INV_X1 U304 ( .A(n904), .ZN(n632) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n821), .B1(n907), .B2(\mem[22][3] ), 
        .ZN(n904) );
  INV_X1 U306 ( .A(n903), .ZN(n631) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n821), .B1(n907), .B2(\mem[22][4] ), 
        .ZN(n903) );
  INV_X1 U308 ( .A(n902), .ZN(n630) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n821), .B1(n907), .B2(\mem[22][5] ), 
        .ZN(n902) );
  INV_X1 U310 ( .A(n901), .ZN(n629) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n821), .B1(n907), .B2(\mem[22][6] ), 
        .ZN(n901) );
  INV_X1 U312 ( .A(n900), .ZN(n628) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n821), .B1(n907), .B2(\mem[22][7] ), 
        .ZN(n900) );
  INV_X1 U314 ( .A(n899), .ZN(n627) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n820), .B1(n898), .B2(\mem[23][0] ), 
        .ZN(n899) );
  INV_X1 U316 ( .A(n897), .ZN(n626) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n820), .B1(n898), .B2(\mem[23][1] ), 
        .ZN(n897) );
  INV_X1 U318 ( .A(n896), .ZN(n625) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n820), .B1(n898), .B2(\mem[23][2] ), 
        .ZN(n896) );
  INV_X1 U320 ( .A(n895), .ZN(n624) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n820), .B1(n898), .B2(\mem[23][3] ), 
        .ZN(n895) );
  INV_X1 U322 ( .A(n894), .ZN(n623) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n820), .B1(n898), .B2(\mem[23][4] ), 
        .ZN(n894) );
  INV_X1 U324 ( .A(n893), .ZN(n622) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n820), .B1(n898), .B2(\mem[23][5] ), 
        .ZN(n893) );
  INV_X1 U326 ( .A(n892), .ZN(n621) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n820), .B1(n898), .B2(\mem[23][6] ), 
        .ZN(n892) );
  INV_X1 U328 ( .A(n891), .ZN(n620) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n820), .B1(n898), .B2(\mem[23][7] ), 
        .ZN(n891) );
  INV_X1 U330 ( .A(N12), .ZN(n255) );
  INV_X1 U331 ( .A(N11), .ZN(n254) );
  INV_X1 U332 ( .A(n999), .ZN(n715) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n831), .B1(n998), .B2(\mem[12][0] ), 
        .ZN(n999) );
  INV_X1 U334 ( .A(n997), .ZN(n714) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n831), .B1(n998), .B2(\mem[12][1] ), 
        .ZN(n997) );
  INV_X1 U336 ( .A(n996), .ZN(n713) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n831), .B1(n998), .B2(\mem[12][2] ), 
        .ZN(n996) );
  INV_X1 U338 ( .A(n995), .ZN(n712) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n831), .B1(n998), .B2(\mem[12][3] ), 
        .ZN(n995) );
  INV_X1 U340 ( .A(n994), .ZN(n711) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n831), .B1(n998), .B2(\mem[12][4] ), 
        .ZN(n994) );
  INV_X1 U342 ( .A(n993), .ZN(n710) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n831), .B1(n998), .B2(\mem[12][5] ), 
        .ZN(n993) );
  INV_X1 U344 ( .A(n992), .ZN(n709) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n831), .B1(n998), .B2(\mem[12][6] ), 
        .ZN(n992) );
  INV_X1 U346 ( .A(n991), .ZN(n708) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n831), .B1(n998), .B2(\mem[12][7] ), 
        .ZN(n991) );
  INV_X1 U348 ( .A(n926), .ZN(n651) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n823), .B1(n925), .B2(\mem[20][0] ), 
        .ZN(n926) );
  INV_X1 U350 ( .A(n924), .ZN(n650) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n823), .B1(n925), .B2(\mem[20][1] ), 
        .ZN(n924) );
  INV_X1 U352 ( .A(n923), .ZN(n649) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n823), .B1(n925), .B2(\mem[20][2] ), 
        .ZN(n923) );
  INV_X1 U354 ( .A(n922), .ZN(n648) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n823), .B1(n925), .B2(\mem[20][3] ), 
        .ZN(n922) );
  INV_X1 U356 ( .A(n921), .ZN(n647) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n823), .B1(n925), .B2(\mem[20][4] ), 
        .ZN(n921) );
  INV_X1 U358 ( .A(n920), .ZN(n646) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n823), .B1(n925), .B2(\mem[20][5] ), 
        .ZN(n920) );
  INV_X1 U360 ( .A(n919), .ZN(n645) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n823), .B1(n925), .B2(\mem[20][6] ), 
        .ZN(n919) );
  INV_X1 U362 ( .A(n918), .ZN(n644) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n823), .B1(n925), .B2(\mem[20][7] ), 
        .ZN(n918) );
  INV_X1 U364 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n835), .B1(n1035), .B2(\mem[8][0] ), 
        .ZN(n1036) );
  INV_X1 U366 ( .A(n1034), .ZN(n746) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n835), .B1(n1035), .B2(\mem[8][1] ), 
        .ZN(n1034) );
  INV_X1 U368 ( .A(n1033), .ZN(n745) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n835), .B1(n1035), .B2(\mem[8][2] ), 
        .ZN(n1033) );
  INV_X1 U370 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n835), .B1(n1035), .B2(\mem[8][3] ), 
        .ZN(n1032) );
  INV_X1 U372 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n835), .B1(n1035), .B2(\mem[8][4] ), 
        .ZN(n1031) );
  INV_X1 U374 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n835), .B1(n1035), .B2(\mem[8][5] ), 
        .ZN(n1030) );
  INV_X1 U376 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n835), .B1(n1035), .B2(\mem[8][6] ), 
        .ZN(n1029) );
  INV_X1 U378 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n835), .B1(n1035), .B2(\mem[8][7] ), 
        .ZN(n1028) );
  INV_X1 U380 ( .A(n963), .ZN(n683) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n827), .B1(n962), .B2(\mem[16][0] ), 
        .ZN(n963) );
  INV_X1 U382 ( .A(n961), .ZN(n682) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n827), .B1(n962), .B2(\mem[16][1] ), 
        .ZN(n961) );
  INV_X1 U384 ( .A(n960), .ZN(n681) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n827), .B1(n962), .B2(\mem[16][2] ), 
        .ZN(n960) );
  INV_X1 U386 ( .A(n959), .ZN(n680) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n827), .B1(n962), .B2(\mem[16][3] ), 
        .ZN(n959) );
  INV_X1 U388 ( .A(n958), .ZN(n679) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n827), .B1(n962), .B2(\mem[16][4] ), 
        .ZN(n958) );
  INV_X1 U390 ( .A(n957), .ZN(n678) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n827), .B1(n962), .B2(\mem[16][5] ), 
        .ZN(n957) );
  INV_X1 U392 ( .A(n956), .ZN(n677) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n827), .B1(n962), .B2(\mem[16][6] ), 
        .ZN(n956) );
  INV_X1 U394 ( .A(n955), .ZN(n676) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n827), .B1(n962), .B2(\mem[16][7] ), 
        .ZN(n955) );
  INV_X1 U396 ( .A(n890), .ZN(n619) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n816), .B1(n889), .B2(\mem[24][0] ), 
        .ZN(n890) );
  INV_X1 U398 ( .A(n888), .ZN(n618) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n816), .B1(n889), .B2(\mem[24][1] ), 
        .ZN(n888) );
  INV_X1 U400 ( .A(n887), .ZN(n617) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n816), .B1(n889), .B2(\mem[24][2] ), 
        .ZN(n887) );
  INV_X1 U402 ( .A(n886), .ZN(n616) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n816), .B1(n889), .B2(\mem[24][3] ), 
        .ZN(n886) );
  INV_X1 U404 ( .A(n885), .ZN(n615) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n816), .B1(n889), .B2(\mem[24][4] ), 
        .ZN(n885) );
  INV_X1 U406 ( .A(n884), .ZN(n614) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n816), .B1(n889), .B2(\mem[24][5] ), 
        .ZN(n884) );
  INV_X1 U408 ( .A(n883), .ZN(n613) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n816), .B1(n889), .B2(\mem[24][6] ), 
        .ZN(n883) );
  INV_X1 U410 ( .A(n882), .ZN(n612) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n816), .B1(n889), .B2(\mem[24][7] ), 
        .ZN(n882) );
  INV_X1 U412 ( .A(n881), .ZN(n611) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n815), .B1(n880), .B2(\mem[25][0] ), 
        .ZN(n881) );
  INV_X1 U414 ( .A(n879), .ZN(n610) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n815), .B1(n880), .B2(\mem[25][1] ), 
        .ZN(n879) );
  INV_X1 U416 ( .A(n878), .ZN(n609) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n815), .B1(n880), .B2(\mem[25][2] ), 
        .ZN(n878) );
  INV_X1 U418 ( .A(n877), .ZN(n608) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n815), .B1(n880), .B2(\mem[25][3] ), 
        .ZN(n877) );
  INV_X1 U420 ( .A(n876), .ZN(n607) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n815), .B1(n880), .B2(\mem[25][4] ), 
        .ZN(n876) );
  INV_X1 U422 ( .A(n875), .ZN(n606) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n815), .B1(n880), .B2(\mem[25][5] ), 
        .ZN(n875) );
  INV_X1 U424 ( .A(n874), .ZN(n605) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n815), .B1(n880), .B2(\mem[25][6] ), 
        .ZN(n874) );
  INV_X1 U426 ( .A(n873), .ZN(n604) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n815), .B1(n880), .B2(\mem[25][7] ), 
        .ZN(n873) );
  INV_X1 U428 ( .A(n872), .ZN(n603) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n814), .B1(n871), .B2(\mem[26][0] ), 
        .ZN(n872) );
  INV_X1 U430 ( .A(n870), .ZN(n602) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n814), .B1(n871), .B2(\mem[26][1] ), 
        .ZN(n870) );
  INV_X1 U432 ( .A(n869), .ZN(n601) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n814), .B1(n871), .B2(\mem[26][2] ), 
        .ZN(n869) );
  INV_X1 U434 ( .A(n868), .ZN(n600) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n814), .B1(n871), .B2(\mem[26][3] ), 
        .ZN(n868) );
  INV_X1 U436 ( .A(n867), .ZN(n599) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n814), .B1(n871), .B2(\mem[26][4] ), 
        .ZN(n867) );
  INV_X1 U438 ( .A(n866), .ZN(n598) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n814), .B1(n871), .B2(\mem[26][5] ), 
        .ZN(n866) );
  INV_X1 U440 ( .A(n865), .ZN(n597) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n814), .B1(n871), .B2(\mem[26][6] ), 
        .ZN(n865) );
  INV_X1 U442 ( .A(n864), .ZN(n596) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n814), .B1(n871), .B2(\mem[26][7] ), 
        .ZN(n864) );
  INV_X1 U444 ( .A(n863), .ZN(n595) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n813), .B1(n862), .B2(\mem[27][0] ), 
        .ZN(n863) );
  INV_X1 U446 ( .A(n861), .ZN(n594) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n813), .B1(n862), .B2(\mem[27][1] ), 
        .ZN(n861) );
  INV_X1 U448 ( .A(n860), .ZN(n293) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n813), .B1(n862), .B2(\mem[27][2] ), 
        .ZN(n860) );
  INV_X1 U450 ( .A(n859), .ZN(n292) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n813), .B1(n862), .B2(\mem[27][3] ), 
        .ZN(n859) );
  INV_X1 U452 ( .A(n858), .ZN(n291) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n813), .B1(n862), .B2(\mem[27][4] ), 
        .ZN(n858) );
  INV_X1 U454 ( .A(n857), .ZN(n290) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n813), .B1(n862), .B2(\mem[27][5] ), 
        .ZN(n857) );
  INV_X1 U456 ( .A(n856), .ZN(n289) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n813), .B1(n862), .B2(\mem[27][6] ), 
        .ZN(n856) );
  INV_X1 U458 ( .A(n855), .ZN(n288) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n813), .B1(n862), .B2(\mem[27][7] ), 
        .ZN(n855) );
  INV_X1 U460 ( .A(n854), .ZN(n287) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n812), .B1(n853), .B2(\mem[28][0] ), 
        .ZN(n854) );
  INV_X1 U462 ( .A(n852), .ZN(n286) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n812), .B1(n853), .B2(\mem[28][1] ), 
        .ZN(n852) );
  INV_X1 U464 ( .A(n851), .ZN(n285) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n812), .B1(n853), .B2(\mem[28][2] ), 
        .ZN(n851) );
  INV_X1 U466 ( .A(n850), .ZN(n284) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n812), .B1(n853), .B2(\mem[28][3] ), 
        .ZN(n850) );
  INV_X1 U468 ( .A(n849), .ZN(n283) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n812), .B1(n853), .B2(\mem[28][4] ), 
        .ZN(n849) );
  INV_X1 U470 ( .A(n848), .ZN(n282) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n812), .B1(n853), .B2(\mem[28][5] ), 
        .ZN(n848) );
  INV_X1 U472 ( .A(n847), .ZN(n281) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n812), .B1(n853), .B2(\mem[28][6] ), 
        .ZN(n847) );
  INV_X1 U474 ( .A(n846), .ZN(n280) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n812), .B1(n853), .B2(\mem[28][7] ), 
        .ZN(n846) );
  INV_X1 U476 ( .A(n1145), .ZN(n279) );
  AOI22_X1 U477 ( .A1(n819), .A2(data_in[0]), .B1(n1144), .B2(\mem[29][0] ), 
        .ZN(n1145) );
  INV_X1 U478 ( .A(n1143), .ZN(n278) );
  AOI22_X1 U479 ( .A1(n819), .A2(data_in[1]), .B1(n1144), .B2(\mem[29][1] ), 
        .ZN(n1143) );
  INV_X1 U480 ( .A(n1142), .ZN(n277) );
  AOI22_X1 U481 ( .A1(n819), .A2(data_in[2]), .B1(n1144), .B2(\mem[29][2] ), 
        .ZN(n1142) );
  INV_X1 U482 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U483 ( .A1(n819), .A2(data_in[3]), .B1(n1144), .B2(\mem[29][3] ), 
        .ZN(n1141) );
  INV_X1 U484 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U485 ( .A1(n819), .A2(data_in[4]), .B1(n1144), .B2(\mem[29][4] ), 
        .ZN(n1140) );
  INV_X1 U486 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U487 ( .A1(n819), .A2(data_in[5]), .B1(n1144), .B2(\mem[29][5] ), 
        .ZN(n1139) );
  INV_X1 U488 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U489 ( .A1(n819), .A2(data_in[6]), .B1(n1144), .B2(\mem[29][6] ), 
        .ZN(n1138) );
  INV_X1 U490 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U491 ( .A1(n819), .A2(data_in[7]), .B1(n1144), .B2(\mem[29][7] ), 
        .ZN(n1137) );
  INV_X1 U492 ( .A(n1134), .ZN(n271) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n818), .B1(n1133), .B2(\mem[30][0] ), 
        .ZN(n1134) );
  INV_X1 U494 ( .A(n1132), .ZN(n270) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n818), .B1(n1133), .B2(\mem[30][1] ), 
        .ZN(n1132) );
  INV_X1 U496 ( .A(n1131), .ZN(n269) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n818), .B1(n1133), .B2(\mem[30][2] ), 
        .ZN(n1131) );
  INV_X1 U498 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n818), .B1(n1133), .B2(\mem[30][3] ), 
        .ZN(n1130) );
  INV_X1 U500 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n818), .B1(n1133), .B2(\mem[30][4] ), 
        .ZN(n1129) );
  INV_X1 U502 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n818), .B1(n1133), .B2(\mem[30][5] ), 
        .ZN(n1128) );
  INV_X1 U504 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n818), .B1(n1133), .B2(\mem[30][6] ), 
        .ZN(n1127) );
  INV_X1 U506 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n818), .B1(n1133), .B2(\mem[30][7] ), 
        .ZN(n1126) );
  INV_X1 U508 ( .A(n1124), .ZN(n263) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n817), .B1(n1123), .B2(\mem[31][0] ), 
        .ZN(n1124) );
  INV_X1 U510 ( .A(n1122), .ZN(n262) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n817), .B1(n1123), .B2(\mem[31][1] ), 
        .ZN(n1122) );
  INV_X1 U512 ( .A(n1121), .ZN(n261) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n817), .B1(n1123), .B2(\mem[31][2] ), 
        .ZN(n1121) );
  INV_X1 U514 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n817), .B1(n1123), .B2(\mem[31][3] ), 
        .ZN(n1120) );
  INV_X1 U516 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n817), .B1(n1123), .B2(\mem[31][4] ), 
        .ZN(n1119) );
  INV_X1 U518 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n817), .B1(n1123), .B2(\mem[31][5] ), 
        .ZN(n1118) );
  INV_X1 U520 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n817), .B1(n1123), .B2(\mem[31][6] ), 
        .ZN(n1117) );
  INV_X1 U522 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n817), .B1(n1123), .B2(\mem[31][7] ), 
        .ZN(n1116) );
  INV_X1 U524 ( .A(n1114), .ZN(n811) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n843), .B1(n1113), .B2(\mem[0][0] ), 
        .ZN(n1114) );
  INV_X1 U526 ( .A(n1112), .ZN(n810) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n843), .B1(n1113), .B2(\mem[0][1] ), 
        .ZN(n1112) );
  INV_X1 U528 ( .A(n1111), .ZN(n809) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n843), .B1(n1113), .B2(\mem[0][2] ), 
        .ZN(n1111) );
  INV_X1 U530 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n843), .B1(n1113), .B2(\mem[0][3] ), 
        .ZN(n1110) );
  INV_X1 U532 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n843), .B1(n1113), .B2(\mem[0][4] ), 
        .ZN(n1109) );
  INV_X1 U534 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n843), .B1(n1113), .B2(\mem[0][5] ), 
        .ZN(n1108) );
  INV_X1 U536 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n843), .B1(n1113), .B2(\mem[0][6] ), 
        .ZN(n1107) );
  INV_X1 U538 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n843), .B1(n1113), .B2(\mem[0][7] ), 
        .ZN(n1106) );
  INV_X1 U540 ( .A(n1103), .ZN(n803) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[1][0] ), 
        .ZN(n1103) );
  INV_X1 U542 ( .A(n1101), .ZN(n802) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[1][1] ), 
        .ZN(n1101) );
  INV_X1 U544 ( .A(n1100), .ZN(n801) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[1][2] ), 
        .ZN(n1100) );
  INV_X1 U546 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[1][3] ), 
        .ZN(n1099) );
  INV_X1 U548 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[1][4] ), 
        .ZN(n1098) );
  INV_X1 U550 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[1][5] ), 
        .ZN(n1097) );
  INV_X1 U552 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[1][6] ), 
        .ZN(n1096) );
  INV_X1 U554 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[1][7] ), 
        .ZN(n1095) );
  INV_X1 U556 ( .A(n1093), .ZN(n795) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n841), .B1(n1092), .B2(\mem[2][0] ), 
        .ZN(n1093) );
  INV_X1 U558 ( .A(n1091), .ZN(n794) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n841), .B1(n1092), .B2(\mem[2][1] ), 
        .ZN(n1091) );
  INV_X1 U560 ( .A(n1090), .ZN(n793) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n841), .B1(n1092), .B2(\mem[2][2] ), 
        .ZN(n1090) );
  INV_X1 U562 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n841), .B1(n1092), .B2(\mem[2][3] ), 
        .ZN(n1089) );
  INV_X1 U564 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n841), .B1(n1092), .B2(\mem[2][4] ), 
        .ZN(n1088) );
  INV_X1 U566 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n841), .B1(n1092), .B2(\mem[2][5] ), 
        .ZN(n1087) );
  INV_X1 U568 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n841), .B1(n1092), .B2(\mem[2][6] ), 
        .ZN(n1086) );
  INV_X1 U570 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n841), .B1(n1092), .B2(\mem[2][7] ), 
        .ZN(n1085) );
  INV_X1 U572 ( .A(n1083), .ZN(n787) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n840), .B1(n1082), .B2(\mem[3][0] ), 
        .ZN(n1083) );
  INV_X1 U574 ( .A(n1081), .ZN(n786) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n840), .B1(n1082), .B2(\mem[3][1] ), 
        .ZN(n1081) );
  INV_X1 U576 ( .A(n1080), .ZN(n785) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n840), .B1(n1082), .B2(\mem[3][2] ), 
        .ZN(n1080) );
  INV_X1 U578 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n840), .B1(n1082), .B2(\mem[3][3] ), 
        .ZN(n1079) );
  INV_X1 U580 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n840), .B1(n1082), .B2(\mem[3][4] ), 
        .ZN(n1078) );
  INV_X1 U582 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n840), .B1(n1082), .B2(\mem[3][5] ), 
        .ZN(n1077) );
  INV_X1 U584 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n840), .B1(n1082), .B2(\mem[3][6] ), 
        .ZN(n1076) );
  INV_X1 U586 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n840), .B1(n1082), .B2(\mem[3][7] ), 
        .ZN(n1075) );
  INV_X1 U588 ( .A(n1073), .ZN(n779) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n839), .B1(n1072), .B2(\mem[4][0] ), 
        .ZN(n1073) );
  INV_X1 U590 ( .A(n1071), .ZN(n778) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n839), .B1(n1072), .B2(\mem[4][1] ), 
        .ZN(n1071) );
  INV_X1 U592 ( .A(n1070), .ZN(n777) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n839), .B1(n1072), .B2(\mem[4][2] ), 
        .ZN(n1070) );
  INV_X1 U594 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n839), .B1(n1072), .B2(\mem[4][3] ), 
        .ZN(n1069) );
  INV_X1 U596 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n839), .B1(n1072), .B2(\mem[4][4] ), 
        .ZN(n1068) );
  INV_X1 U598 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n839), .B1(n1072), .B2(\mem[4][5] ), 
        .ZN(n1067) );
  INV_X1 U600 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n839), .B1(n1072), .B2(\mem[4][6] ), 
        .ZN(n1066) );
  INV_X1 U602 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n839), .B1(n1072), .B2(\mem[4][7] ), 
        .ZN(n1065) );
  INV_X1 U604 ( .A(N13), .ZN(n844) );
  INV_X1 U605 ( .A(N14), .ZN(n845) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n251), .Z(n3) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n251), .Z(n4) );
  MUX2_X1 U608 ( .A(n4), .B(n3), .S(n244), .Z(n5) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n251), .Z(n6) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n248), .Z(n7) );
  MUX2_X1 U611 ( .A(n7), .B(n6), .S(n244), .Z(n8) );
  MUX2_X1 U612 ( .A(n8), .B(n5), .S(n243), .Z(n9) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n251), .Z(n10) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n247), .Z(n11) );
  MUX2_X1 U615 ( .A(n11), .B(n10), .S(n244), .Z(n12) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n247), .Z(n13) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n249), .Z(n14) );
  MUX2_X1 U618 ( .A(n14), .B(n13), .S(n244), .Z(n15) );
  MUX2_X1 U619 ( .A(n15), .B(n12), .S(N12), .Z(n16) );
  MUX2_X1 U620 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n247), .Z(n18) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n247), .Z(n19) );
  MUX2_X1 U623 ( .A(n19), .B(n18), .S(N11), .Z(n20) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n247), .Z(n21) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n247), .Z(n22) );
  MUX2_X1 U626 ( .A(n22), .B(n21), .S(n244), .Z(n23) );
  MUX2_X1 U627 ( .A(n23), .B(n20), .S(N12), .Z(n24) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n247), .Z(n25) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n247), .Z(n26) );
  MUX2_X1 U630 ( .A(n26), .B(n25), .S(n246), .Z(n27) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n247), .Z(n28) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n247), .Z(n29) );
  MUX2_X1 U633 ( .A(n29), .B(n28), .S(n246), .Z(n30) );
  MUX2_X1 U634 ( .A(n30), .B(n27), .S(N12), .Z(n31) );
  MUX2_X1 U635 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U636 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n247), .Z(n33) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n247), .Z(n34) );
  MUX2_X1 U639 ( .A(n34), .B(n33), .S(N11), .Z(n35) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n247), .Z(n36) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n247), .Z(n37) );
  MUX2_X1 U642 ( .A(n37), .B(n36), .S(N11), .Z(n38) );
  MUX2_X1 U643 ( .A(n38), .B(n35), .S(n243), .Z(n39) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n248), .Z(n40) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n248), .Z(n41) );
  MUX2_X1 U646 ( .A(n41), .B(n40), .S(N11), .Z(n42) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n248), .Z(n43) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n248), .Z(n44) );
  MUX2_X1 U649 ( .A(n44), .B(n43), .S(n244), .Z(n45) );
  MUX2_X1 U650 ( .A(n45), .B(n42), .S(n243), .Z(n46) );
  MUX2_X1 U651 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n248), .Z(n48) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n248), .Z(n49) );
  MUX2_X1 U654 ( .A(n49), .B(n48), .S(N11), .Z(n50) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n248), .Z(n51) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n248), .Z(n52) );
  MUX2_X1 U657 ( .A(n52), .B(n51), .S(n246), .Z(n53) );
  MUX2_X1 U658 ( .A(n53), .B(n50), .S(n243), .Z(n54) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n248), .Z(n55) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n248), .Z(n56) );
  MUX2_X1 U661 ( .A(n56), .B(n55), .S(n245), .Z(n57) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n248), .Z(n58) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n248), .Z(n59) );
  MUX2_X1 U664 ( .A(n59), .B(n58), .S(n245), .Z(n60) );
  MUX2_X1 U665 ( .A(n60), .B(n57), .S(n243), .Z(n61) );
  MUX2_X1 U666 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U667 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n249), .Z(n63) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n249), .Z(n64) );
  MUX2_X1 U670 ( .A(n64), .B(n63), .S(n246), .Z(n65) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n249), .Z(n66) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n249), .Z(n67) );
  MUX2_X1 U673 ( .A(n67), .B(n66), .S(N11), .Z(n68) );
  MUX2_X1 U674 ( .A(n68), .B(n65), .S(n243), .Z(n69) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n249), .Z(n70) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n249), .Z(n71) );
  MUX2_X1 U677 ( .A(n71), .B(n70), .S(N11), .Z(n72) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n249), .Z(n73) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n249), .Z(n74) );
  MUX2_X1 U680 ( .A(n74), .B(n73), .S(N11), .Z(n75) );
  MUX2_X1 U681 ( .A(n75), .B(n72), .S(n243), .Z(n76) );
  MUX2_X1 U682 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n249), .Z(n78) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n249), .Z(n79) );
  MUX2_X1 U685 ( .A(n79), .B(n78), .S(n245), .Z(n80) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n249), .Z(n81) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n249), .Z(n82) );
  MUX2_X1 U688 ( .A(n82), .B(n81), .S(N11), .Z(n83) );
  MUX2_X1 U689 ( .A(n83), .B(n80), .S(n243), .Z(n84) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n250), .Z(n85) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n250), .Z(n86) );
  MUX2_X1 U692 ( .A(n86), .B(n85), .S(N11), .Z(n87) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n250), .Z(n88) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n250), .Z(n89) );
  MUX2_X1 U695 ( .A(n89), .B(n88), .S(N11), .Z(n90) );
  MUX2_X1 U696 ( .A(n90), .B(n87), .S(n243), .Z(n91) );
  MUX2_X1 U697 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U698 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n250), .Z(n93) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U701 ( .A(n94), .B(n93), .S(N11), .Z(n95) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n250), .Z(n96) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n250), .Z(n97) );
  MUX2_X1 U704 ( .A(n97), .B(n96), .S(n246), .Z(n98) );
  MUX2_X1 U705 ( .A(n98), .B(n95), .S(n243), .Z(n99) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n100) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n250), .Z(n101) );
  MUX2_X1 U708 ( .A(n101), .B(n100), .S(n245), .Z(n102) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n250), .Z(n103) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n250), .Z(n104) );
  MUX2_X1 U711 ( .A(n104), .B(n103), .S(n244), .Z(n105) );
  MUX2_X1 U712 ( .A(n105), .B(n102), .S(n243), .Z(n106) );
  MUX2_X1 U713 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n251), .Z(n108) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n249), .Z(n109) );
  MUX2_X1 U716 ( .A(n109), .B(n108), .S(n244), .Z(n110) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n252), .Z(n111) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n250), .Z(n112) );
  MUX2_X1 U719 ( .A(n112), .B(n111), .S(n244), .Z(n113) );
  MUX2_X1 U720 ( .A(n113), .B(n110), .S(n243), .Z(n114) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n247), .Z(n115) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n252), .Z(n116) );
  MUX2_X1 U723 ( .A(n116), .B(n115), .S(n244), .Z(n117) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n248), .Z(n118) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n119) );
  MUX2_X1 U726 ( .A(n119), .B(n118), .S(n244), .Z(n120) );
  MUX2_X1 U727 ( .A(n120), .B(n117), .S(n243), .Z(n121) );
  MUX2_X1 U728 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U729 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(N10), .Z(n123) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(N10), .Z(n124) );
  MUX2_X1 U732 ( .A(n124), .B(n123), .S(n244), .Z(n125) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(N10), .Z(n126) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n127) );
  MUX2_X1 U735 ( .A(n127), .B(n126), .S(n245), .Z(n128) );
  MUX2_X1 U736 ( .A(n128), .B(n125), .S(n243), .Z(n129) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n251), .Z(n130) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n252), .Z(n131) );
  MUX2_X1 U739 ( .A(n131), .B(n130), .S(n244), .Z(n132) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n251), .Z(n133) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(N10), .Z(n134) );
  MUX2_X1 U742 ( .A(n134), .B(n133), .S(N11), .Z(n135) );
  MUX2_X1 U743 ( .A(n135), .B(n132), .S(n243), .Z(n136) );
  MUX2_X1 U744 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n251), .Z(n138) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n252), .Z(n139) );
  MUX2_X1 U747 ( .A(n139), .B(n138), .S(n244), .Z(n140) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n251), .Z(n141) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(N10), .Z(n142) );
  MUX2_X1 U750 ( .A(n142), .B(n141), .S(n245), .Z(n143) );
  MUX2_X1 U751 ( .A(n143), .B(n140), .S(n243), .Z(n144) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(N10), .Z(n145) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(N10), .Z(n146) );
  MUX2_X1 U754 ( .A(n146), .B(n145), .S(n246), .Z(n147) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(N10), .Z(n148) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n149) );
  MUX2_X1 U757 ( .A(n149), .B(n148), .S(n244), .Z(n150) );
  MUX2_X1 U758 ( .A(n150), .B(n147), .S(n243), .Z(n151) );
  MUX2_X1 U759 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U760 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n251), .Z(n153) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n251), .Z(n154) );
  MUX2_X1 U763 ( .A(n154), .B(n153), .S(n245), .Z(n155) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n251), .Z(n156) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n251), .Z(n157) );
  MUX2_X1 U766 ( .A(n157), .B(n156), .S(n245), .Z(n158) );
  MUX2_X1 U767 ( .A(n158), .B(n155), .S(n243), .Z(n159) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n251), .Z(n160) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n251), .Z(n161) );
  MUX2_X1 U770 ( .A(n161), .B(n160), .S(n245), .Z(n162) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n251), .Z(n163) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n251), .Z(n164) );
  MUX2_X1 U773 ( .A(n164), .B(n163), .S(n245), .Z(n165) );
  MUX2_X1 U774 ( .A(n165), .B(n162), .S(N12), .Z(n166) );
  MUX2_X1 U775 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n251), .Z(n168) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n251), .Z(n169) );
  MUX2_X1 U778 ( .A(n169), .B(n168), .S(n245), .Z(n170) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n251), .Z(n171) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n251), .Z(n172) );
  MUX2_X1 U781 ( .A(n172), .B(n171), .S(n245), .Z(n173) );
  MUX2_X1 U782 ( .A(n173), .B(n170), .S(n243), .Z(n174) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n248), .Z(n175) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n252), .Z(n176) );
  MUX2_X1 U785 ( .A(n176), .B(n175), .S(n245), .Z(n177) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n252), .Z(n178) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n252), .Z(n179) );
  MUX2_X1 U788 ( .A(n179), .B(n178), .S(n245), .Z(n180) );
  MUX2_X1 U789 ( .A(n180), .B(n177), .S(N12), .Z(n181) );
  MUX2_X1 U790 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U791 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n252), .Z(n183) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n250), .Z(n184) );
  MUX2_X1 U794 ( .A(n184), .B(n183), .S(n245), .Z(n185) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n251), .Z(n186) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n247), .Z(n187) );
  MUX2_X1 U797 ( .A(n187), .B(n186), .S(n245), .Z(n188) );
  MUX2_X1 U798 ( .A(n188), .B(n185), .S(n243), .Z(n189) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n252), .Z(n190) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n252), .Z(n191) );
  MUX2_X1 U801 ( .A(n191), .B(n190), .S(n245), .Z(n192) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n249), .Z(n193) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n248), .Z(n194) );
  MUX2_X1 U804 ( .A(n194), .B(n193), .S(n245), .Z(n195) );
  MUX2_X1 U805 ( .A(n195), .B(n192), .S(N12), .Z(n196) );
  MUX2_X1 U806 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n248), .Z(n198) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n252), .Z(n199) );
  MUX2_X1 U809 ( .A(n199), .B(n198), .S(n246), .Z(n200) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n247), .Z(n201) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n250), .Z(n202) );
  MUX2_X1 U812 ( .A(n202), .B(n201), .S(n246), .Z(n203) );
  MUX2_X1 U813 ( .A(n203), .B(n200), .S(n243), .Z(n204) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n252), .Z(n205) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n249), .Z(n206) );
  MUX2_X1 U816 ( .A(n206), .B(n205), .S(n246), .Z(n207) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n248), .Z(n208) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n247), .Z(n209) );
  MUX2_X1 U819 ( .A(n209), .B(n208), .S(n246), .Z(n210) );
  MUX2_X1 U820 ( .A(n210), .B(n207), .S(N12), .Z(n211) );
  MUX2_X1 U821 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U822 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n252), .Z(n213) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n249), .Z(n214) );
  MUX2_X1 U825 ( .A(n214), .B(n213), .S(n246), .Z(n215) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n250), .Z(n216) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n252), .Z(n217) );
  MUX2_X1 U828 ( .A(n217), .B(n216), .S(n246), .Z(n218) );
  MUX2_X1 U829 ( .A(n218), .B(n215), .S(n243), .Z(n219) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n252), .Z(n220) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n252), .Z(n221) );
  MUX2_X1 U832 ( .A(n221), .B(n220), .S(n246), .Z(n222) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(N10), .Z(n223) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n249), .Z(n224) );
  MUX2_X1 U835 ( .A(n224), .B(n223), .S(n246), .Z(n225) );
  MUX2_X1 U836 ( .A(n225), .B(n222), .S(N12), .Z(n226) );
  MUX2_X1 U837 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n252), .Z(n228) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n229) );
  MUX2_X1 U840 ( .A(n229), .B(n228), .S(n246), .Z(n230) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n251), .Z(n231) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n250), .Z(n232) );
  MUX2_X1 U843 ( .A(n232), .B(n231), .S(n246), .Z(n233) );
  MUX2_X1 U844 ( .A(n233), .B(n230), .S(n243), .Z(n234) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n235) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n252), .Z(n236) );
  MUX2_X1 U847 ( .A(n236), .B(n235), .S(n246), .Z(n237) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n252), .Z(n238) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n252), .Z(n239) );
  MUX2_X1 U850 ( .A(n239), .B(n238), .S(n246), .Z(n240) );
  MUX2_X1 U851 ( .A(n240), .B(n237), .S(N12), .Z(n241) );
  MUX2_X1 U852 ( .A(n241), .B(n234), .S(N13), .Z(n242) );
  MUX2_X1 U853 ( .A(n242), .B(n227), .S(N14), .Z(N15) );
  CLKBUF_X1 U854 ( .A(N11), .Z(n244) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_17 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n256), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n257), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n258), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n259), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n260), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n261), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n262), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n263), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n264), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n265), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n266), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n267), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n268), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n269), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n270), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n271), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n272), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n273), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n274), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n275), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n276), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n277), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n278), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n279), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n280), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n281), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n282), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n283), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n284), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n285), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n286), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n287), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n288), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n289), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n290), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n291), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n292), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n293), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n594), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n595), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n596), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n597), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n598), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n599), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n600), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n601), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n602), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n603), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n604), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n605), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n606), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n607), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n608), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n609), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n610), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n611), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n612), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n613), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n614), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n615), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n616), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n617), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n618), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n619), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n620), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n621), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n622), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n623), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n624), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n625), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n626), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n627), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n628), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n629), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n630), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n631), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n632), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n633), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n634), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n635), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n636), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n637), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n638), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n639), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n640), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n641), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n642), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n643), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n644), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n645), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n646), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n647), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n648), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n649), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n650), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n651), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n652), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n653), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n654), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n655), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n656), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n657), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n658), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n659), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n660), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n661), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n662), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n663), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n664), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n665), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n666), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n667), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n668), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n669), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n670), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n671), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n672), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n673), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n674), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n675), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n676), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n677), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n678), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n679), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n680), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n681), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n682), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n683), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n684), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n685), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n686), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n687), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n688), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n689), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n690), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n691), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n692), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n693), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n694), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n695), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n696), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n697), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n698), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n699), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n700), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n701), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n702), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n703), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n704), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n705), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n706), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n707), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n708), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n709), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n710), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n711), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n712), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n713), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n714), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n715), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n716), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n717), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n718), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n719), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n720), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n721), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n722), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n723), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n724), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n725), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n726), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n727), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n728), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n729), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n730), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n731), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n732), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n733), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n734), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n735), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n736), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n737), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n738), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n739), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n740), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n741), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n742), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n743), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n744), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n745), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n746), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n747), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n748), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n749), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n750), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n751), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n752), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n753), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n754), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n755), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n756), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n757), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n758), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n759), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n760), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n761), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n762), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n763), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n764), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n765), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n766), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n767), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n768), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n769), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n770), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n771), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n772), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n773), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n774), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n775), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n776), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n777), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n778), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n779), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n780), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n781), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n782), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n783), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n784), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n785), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n786), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n787), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n788), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n789), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n790), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n791), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n792), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n793), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n794), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n795), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n796), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n797), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n798), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n799), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n800), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n801), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n802), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n803), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n804), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n805), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n806), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n807), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n808), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n809), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n810), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n811), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(n252), .Z(n250) );
  BUF_X1 U5 ( .A(N10), .Z(n251) );
  BUF_X1 U6 ( .A(n252), .Z(n247) );
  BUF_X1 U7 ( .A(n252), .Z(n248) );
  BUF_X1 U8 ( .A(n252), .Z(n249) );
  BUF_X1 U9 ( .A(N10), .Z(n252) );
  INV_X1 U10 ( .A(n1113), .ZN(n843) );
  INV_X1 U11 ( .A(n1102), .ZN(n842) );
  INV_X1 U12 ( .A(n1092), .ZN(n841) );
  INV_X1 U13 ( .A(n1082), .ZN(n840) );
  INV_X1 U14 ( .A(n1072), .ZN(n839) );
  INV_X1 U15 ( .A(n1062), .ZN(n838) );
  INV_X1 U16 ( .A(n1053), .ZN(n837) );
  INV_X1 U17 ( .A(n1044), .ZN(n836) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1105) );
  NOR3_X1 U19 ( .A1(N11), .A2(N12), .A3(n253), .ZN(n1094) );
  NAND2_X1 U20 ( .A1(n1104), .A2(n1136), .ZN(n1062) );
  NAND2_X1 U21 ( .A1(n1105), .A2(n1104), .ZN(n1113) );
  NAND2_X1 U22 ( .A1(n1094), .A2(n1104), .ZN(n1102) );
  NAND2_X1 U23 ( .A1(n1084), .A2(n1104), .ZN(n1092) );
  NAND2_X1 U24 ( .A1(n1074), .A2(n1104), .ZN(n1082) );
  NAND2_X1 U25 ( .A1(n1064), .A2(n1104), .ZN(n1072) );
  NAND2_X1 U26 ( .A1(n1104), .A2(n1125), .ZN(n1053) );
  NAND2_X1 U27 ( .A1(n1104), .A2(n1115), .ZN(n1044) );
  INV_X1 U28 ( .A(n1133), .ZN(n818) );
  INV_X1 U29 ( .A(n1123), .ZN(n817) );
  INV_X1 U30 ( .A(n889), .ZN(n816) );
  INV_X1 U31 ( .A(n880), .ZN(n815) );
  INV_X1 U32 ( .A(n871), .ZN(n814) );
  INV_X1 U33 ( .A(n862), .ZN(n813) );
  INV_X1 U34 ( .A(n853), .ZN(n812) );
  INV_X1 U35 ( .A(n989), .ZN(n830) );
  INV_X1 U36 ( .A(n980), .ZN(n829) );
  INV_X1 U37 ( .A(n971), .ZN(n828) );
  INV_X1 U38 ( .A(n916), .ZN(n822) );
  INV_X1 U39 ( .A(n907), .ZN(n821) );
  INV_X1 U40 ( .A(n898), .ZN(n820) );
  INV_X1 U41 ( .A(n1035), .ZN(n835) );
  INV_X1 U42 ( .A(n1025), .ZN(n834) );
  INV_X1 U43 ( .A(n1016), .ZN(n833) );
  INV_X1 U44 ( .A(n1007), .ZN(n832) );
  INV_X1 U45 ( .A(n998), .ZN(n831) );
  INV_X1 U46 ( .A(n962), .ZN(n827) );
  INV_X1 U47 ( .A(n952), .ZN(n826) );
  INV_X1 U48 ( .A(n943), .ZN(n825) );
  INV_X1 U49 ( .A(n934), .ZN(n824) );
  INV_X1 U50 ( .A(n925), .ZN(n823) );
  INV_X1 U51 ( .A(n1144), .ZN(n819) );
  BUF_X1 U52 ( .A(N11), .Z(n244) );
  BUF_X1 U53 ( .A(N11), .Z(n245) );
  BUF_X1 U54 ( .A(N11), .Z(n246) );
  INV_X1 U55 ( .A(N10), .ZN(n253) );
  BUF_X1 U56 ( .A(N12), .Z(n243) );
  NOR3_X1 U57 ( .A1(n255), .A2(N10), .A3(n254), .ZN(n1125) );
  NOR3_X1 U58 ( .A1(n255), .A2(n253), .A3(n254), .ZN(n1115) );
  NOR3_X1 U59 ( .A1(n253), .A2(N11), .A3(n255), .ZN(n1136) );
  NOR3_X1 U60 ( .A1(N10), .A2(N12), .A3(n254), .ZN(n1084) );
  NOR3_X1 U61 ( .A1(n253), .A2(N12), .A3(n254), .ZN(n1074) );
  NOR3_X1 U62 ( .A1(N10), .A2(N11), .A3(n255), .ZN(n1064) );
  NAND2_X1 U63 ( .A1(n1027), .A2(n1136), .ZN(n989) );
  NAND2_X1 U64 ( .A1(n954), .A2(n1136), .ZN(n916) );
  NAND2_X1 U65 ( .A1(n1027), .A2(n1064), .ZN(n998) );
  NAND2_X1 U66 ( .A1(n954), .A2(n1064), .ZN(n925) );
  NAND2_X1 U67 ( .A1(n1027), .A2(n1105), .ZN(n1035) );
  NAND2_X1 U68 ( .A1(n1027), .A2(n1094), .ZN(n1025) );
  NAND2_X1 U69 ( .A1(n954), .A2(n1105), .ZN(n962) );
  NAND2_X1 U70 ( .A1(n954), .A2(n1094), .ZN(n952) );
  NAND2_X1 U71 ( .A1(n1105), .A2(n1135), .ZN(n889) );
  NAND2_X1 U72 ( .A1(n1094), .A2(n1135), .ZN(n880) );
  NAND2_X1 U73 ( .A1(n1084), .A2(n1135), .ZN(n871) );
  NAND2_X1 U74 ( .A1(n1074), .A2(n1135), .ZN(n862) );
  NAND2_X1 U75 ( .A1(n1064), .A2(n1135), .ZN(n853) );
  NAND2_X1 U76 ( .A1(n1136), .A2(n1135), .ZN(n1144) );
  NAND2_X1 U77 ( .A1(n1125), .A2(n1135), .ZN(n1133) );
  NAND2_X1 U78 ( .A1(n1115), .A2(n1135), .ZN(n1123) );
  NAND2_X1 U79 ( .A1(n1027), .A2(n1084), .ZN(n1016) );
  NAND2_X1 U80 ( .A1(n1027), .A2(n1074), .ZN(n1007) );
  NAND2_X1 U81 ( .A1(n954), .A2(n1084), .ZN(n943) );
  NAND2_X1 U82 ( .A1(n954), .A2(n1074), .ZN(n934) );
  NAND2_X1 U83 ( .A1(n1027), .A2(n1125), .ZN(n980) );
  NAND2_X1 U84 ( .A1(n954), .A2(n1125), .ZN(n907) );
  NAND2_X1 U85 ( .A1(n1027), .A2(n1115), .ZN(n971) );
  NAND2_X1 U86 ( .A1(n954), .A2(n1115), .ZN(n898) );
  AND3_X1 U87 ( .A1(n844), .A2(n845), .A3(wr_en), .ZN(n1104) );
  AND3_X1 U88 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1135) );
  AND3_X1 U89 ( .A1(N13), .A2(n845), .A3(wr_en), .ZN(n1027) );
  AND3_X1 U90 ( .A1(N14), .A2(n844), .A3(wr_en), .ZN(n954) );
  INV_X1 U91 ( .A(n1063), .ZN(n771) );
  AOI22_X1 U92 ( .A1(data_in[0]), .A2(n838), .B1(n1062), .B2(\mem[5][0] ), 
        .ZN(n1063) );
  INV_X1 U93 ( .A(n1061), .ZN(n770) );
  AOI22_X1 U94 ( .A1(data_in[1]), .A2(n838), .B1(n1062), .B2(\mem[5][1] ), 
        .ZN(n1061) );
  INV_X1 U95 ( .A(n1060), .ZN(n769) );
  AOI22_X1 U96 ( .A1(data_in[2]), .A2(n838), .B1(n1062), .B2(\mem[5][2] ), 
        .ZN(n1060) );
  INV_X1 U97 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U98 ( .A1(data_in[3]), .A2(n838), .B1(n1062), .B2(\mem[5][3] ), 
        .ZN(n1059) );
  INV_X1 U99 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U100 ( .A1(data_in[4]), .A2(n838), .B1(n1062), .B2(\mem[5][4] ), 
        .ZN(n1058) );
  INV_X1 U101 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U102 ( .A1(data_in[5]), .A2(n838), .B1(n1062), .B2(\mem[5][5] ), 
        .ZN(n1057) );
  INV_X1 U103 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U104 ( .A1(data_in[6]), .A2(n838), .B1(n1062), .B2(\mem[5][6] ), 
        .ZN(n1056) );
  INV_X1 U105 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U106 ( .A1(data_in[7]), .A2(n838), .B1(n1062), .B2(\mem[5][7] ), 
        .ZN(n1055) );
  INV_X1 U107 ( .A(n1026), .ZN(n739) );
  AOI22_X1 U108 ( .A1(data_in[0]), .A2(n834), .B1(n1025), .B2(\mem[9][0] ), 
        .ZN(n1026) );
  INV_X1 U109 ( .A(n1024), .ZN(n738) );
  AOI22_X1 U110 ( .A1(data_in[1]), .A2(n834), .B1(n1025), .B2(\mem[9][1] ), 
        .ZN(n1024) );
  INV_X1 U111 ( .A(n1023), .ZN(n737) );
  AOI22_X1 U112 ( .A1(data_in[2]), .A2(n834), .B1(n1025), .B2(\mem[9][2] ), 
        .ZN(n1023) );
  INV_X1 U113 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U114 ( .A1(data_in[3]), .A2(n834), .B1(n1025), .B2(\mem[9][3] ), 
        .ZN(n1022) );
  INV_X1 U115 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U116 ( .A1(data_in[4]), .A2(n834), .B1(n1025), .B2(\mem[9][4] ), 
        .ZN(n1021) );
  INV_X1 U117 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U118 ( .A1(data_in[5]), .A2(n834), .B1(n1025), .B2(\mem[9][5] ), 
        .ZN(n1020) );
  INV_X1 U119 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U120 ( .A1(data_in[6]), .A2(n834), .B1(n1025), .B2(\mem[9][6] ), 
        .ZN(n1019) );
  INV_X1 U121 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U122 ( .A1(data_in[7]), .A2(n834), .B1(n1025), .B2(\mem[9][7] ), 
        .ZN(n1018) );
  INV_X1 U123 ( .A(n990), .ZN(n707) );
  AOI22_X1 U124 ( .A1(data_in[0]), .A2(n830), .B1(n989), .B2(\mem[13][0] ), 
        .ZN(n990) );
  INV_X1 U125 ( .A(n988), .ZN(n706) );
  AOI22_X1 U126 ( .A1(data_in[1]), .A2(n830), .B1(n989), .B2(\mem[13][1] ), 
        .ZN(n988) );
  INV_X1 U127 ( .A(n987), .ZN(n705) );
  AOI22_X1 U128 ( .A1(data_in[2]), .A2(n830), .B1(n989), .B2(\mem[13][2] ), 
        .ZN(n987) );
  INV_X1 U129 ( .A(n986), .ZN(n704) );
  AOI22_X1 U130 ( .A1(data_in[3]), .A2(n830), .B1(n989), .B2(\mem[13][3] ), 
        .ZN(n986) );
  INV_X1 U131 ( .A(n985), .ZN(n703) );
  AOI22_X1 U132 ( .A1(data_in[4]), .A2(n830), .B1(n989), .B2(\mem[13][4] ), 
        .ZN(n985) );
  INV_X1 U133 ( .A(n984), .ZN(n702) );
  AOI22_X1 U134 ( .A1(data_in[5]), .A2(n830), .B1(n989), .B2(\mem[13][5] ), 
        .ZN(n984) );
  INV_X1 U135 ( .A(n983), .ZN(n701) );
  AOI22_X1 U136 ( .A1(data_in[6]), .A2(n830), .B1(n989), .B2(\mem[13][6] ), 
        .ZN(n983) );
  INV_X1 U137 ( .A(n982), .ZN(n700) );
  AOI22_X1 U138 ( .A1(data_in[7]), .A2(n830), .B1(n989), .B2(\mem[13][7] ), 
        .ZN(n982) );
  INV_X1 U139 ( .A(n953), .ZN(n675) );
  AOI22_X1 U140 ( .A1(data_in[0]), .A2(n826), .B1(n952), .B2(\mem[17][0] ), 
        .ZN(n953) );
  INV_X1 U141 ( .A(n951), .ZN(n674) );
  AOI22_X1 U142 ( .A1(data_in[1]), .A2(n826), .B1(n952), .B2(\mem[17][1] ), 
        .ZN(n951) );
  INV_X1 U143 ( .A(n950), .ZN(n673) );
  AOI22_X1 U144 ( .A1(data_in[2]), .A2(n826), .B1(n952), .B2(\mem[17][2] ), 
        .ZN(n950) );
  INV_X1 U145 ( .A(n949), .ZN(n672) );
  AOI22_X1 U146 ( .A1(data_in[3]), .A2(n826), .B1(n952), .B2(\mem[17][3] ), 
        .ZN(n949) );
  INV_X1 U147 ( .A(n948), .ZN(n671) );
  AOI22_X1 U148 ( .A1(data_in[4]), .A2(n826), .B1(n952), .B2(\mem[17][4] ), 
        .ZN(n948) );
  INV_X1 U149 ( .A(n947), .ZN(n670) );
  AOI22_X1 U150 ( .A1(data_in[5]), .A2(n826), .B1(n952), .B2(\mem[17][5] ), 
        .ZN(n947) );
  INV_X1 U151 ( .A(n946), .ZN(n669) );
  AOI22_X1 U152 ( .A1(data_in[6]), .A2(n826), .B1(n952), .B2(\mem[17][6] ), 
        .ZN(n946) );
  INV_X1 U153 ( .A(n945), .ZN(n668) );
  AOI22_X1 U154 ( .A1(data_in[7]), .A2(n826), .B1(n952), .B2(\mem[17][7] ), 
        .ZN(n945) );
  INV_X1 U155 ( .A(n917), .ZN(n643) );
  AOI22_X1 U156 ( .A1(data_in[0]), .A2(n822), .B1(n916), .B2(\mem[21][0] ), 
        .ZN(n917) );
  INV_X1 U157 ( .A(n915), .ZN(n642) );
  AOI22_X1 U158 ( .A1(data_in[1]), .A2(n822), .B1(n916), .B2(\mem[21][1] ), 
        .ZN(n915) );
  INV_X1 U159 ( .A(n914), .ZN(n641) );
  AOI22_X1 U160 ( .A1(data_in[2]), .A2(n822), .B1(n916), .B2(\mem[21][2] ), 
        .ZN(n914) );
  INV_X1 U161 ( .A(n913), .ZN(n640) );
  AOI22_X1 U162 ( .A1(data_in[3]), .A2(n822), .B1(n916), .B2(\mem[21][3] ), 
        .ZN(n913) );
  INV_X1 U163 ( .A(n912), .ZN(n639) );
  AOI22_X1 U164 ( .A1(data_in[4]), .A2(n822), .B1(n916), .B2(\mem[21][4] ), 
        .ZN(n912) );
  INV_X1 U165 ( .A(n911), .ZN(n638) );
  AOI22_X1 U166 ( .A1(data_in[5]), .A2(n822), .B1(n916), .B2(\mem[21][5] ), 
        .ZN(n911) );
  INV_X1 U167 ( .A(n910), .ZN(n637) );
  AOI22_X1 U168 ( .A1(data_in[6]), .A2(n822), .B1(n916), .B2(\mem[21][6] ), 
        .ZN(n910) );
  INV_X1 U169 ( .A(n909), .ZN(n636) );
  AOI22_X1 U170 ( .A1(data_in[7]), .A2(n822), .B1(n916), .B2(\mem[21][7] ), 
        .ZN(n909) );
  INV_X1 U171 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U172 ( .A1(data_in[0]), .A2(n833), .B1(n1016), .B2(\mem[10][0] ), 
        .ZN(n1017) );
  INV_X1 U173 ( .A(n1015), .ZN(n730) );
  AOI22_X1 U174 ( .A1(data_in[1]), .A2(n833), .B1(n1016), .B2(\mem[10][1] ), 
        .ZN(n1015) );
  INV_X1 U175 ( .A(n1014), .ZN(n729) );
  AOI22_X1 U176 ( .A1(data_in[2]), .A2(n833), .B1(n1016), .B2(\mem[10][2] ), 
        .ZN(n1014) );
  INV_X1 U177 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U178 ( .A1(data_in[3]), .A2(n833), .B1(n1016), .B2(\mem[10][3] ), 
        .ZN(n1013) );
  INV_X1 U179 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U180 ( .A1(data_in[4]), .A2(n833), .B1(n1016), .B2(\mem[10][4] ), 
        .ZN(n1012) );
  INV_X1 U181 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U182 ( .A1(data_in[5]), .A2(n833), .B1(n1016), .B2(\mem[10][5] ), 
        .ZN(n1011) );
  INV_X1 U183 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U184 ( .A1(data_in[6]), .A2(n833), .B1(n1016), .B2(\mem[10][6] ), 
        .ZN(n1010) );
  INV_X1 U185 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U186 ( .A1(data_in[7]), .A2(n833), .B1(n1016), .B2(\mem[10][7] ), 
        .ZN(n1009) );
  INV_X1 U187 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U188 ( .A1(data_in[0]), .A2(n832), .B1(n1007), .B2(\mem[11][0] ), 
        .ZN(n1008) );
  INV_X1 U189 ( .A(n1006), .ZN(n722) );
  AOI22_X1 U190 ( .A1(data_in[1]), .A2(n832), .B1(n1007), .B2(\mem[11][1] ), 
        .ZN(n1006) );
  INV_X1 U191 ( .A(n1005), .ZN(n721) );
  AOI22_X1 U192 ( .A1(data_in[2]), .A2(n832), .B1(n1007), .B2(\mem[11][2] ), 
        .ZN(n1005) );
  INV_X1 U193 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U194 ( .A1(data_in[3]), .A2(n832), .B1(n1007), .B2(\mem[11][3] ), 
        .ZN(n1004) );
  INV_X1 U195 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U196 ( .A1(data_in[4]), .A2(n832), .B1(n1007), .B2(\mem[11][4] ), 
        .ZN(n1003) );
  INV_X1 U197 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U198 ( .A1(data_in[5]), .A2(n832), .B1(n1007), .B2(\mem[11][5] ), 
        .ZN(n1002) );
  INV_X1 U199 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U200 ( .A1(data_in[6]), .A2(n832), .B1(n1007), .B2(\mem[11][6] ), 
        .ZN(n1001) );
  INV_X1 U201 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U202 ( .A1(data_in[7]), .A2(n832), .B1(n1007), .B2(\mem[11][7] ), 
        .ZN(n1000) );
  INV_X1 U203 ( .A(n981), .ZN(n699) );
  AOI22_X1 U204 ( .A1(data_in[0]), .A2(n829), .B1(n980), .B2(\mem[14][0] ), 
        .ZN(n981) );
  INV_X1 U205 ( .A(n979), .ZN(n698) );
  AOI22_X1 U206 ( .A1(data_in[1]), .A2(n829), .B1(n980), .B2(\mem[14][1] ), 
        .ZN(n979) );
  INV_X1 U207 ( .A(n978), .ZN(n697) );
  AOI22_X1 U208 ( .A1(data_in[2]), .A2(n829), .B1(n980), .B2(\mem[14][2] ), 
        .ZN(n978) );
  INV_X1 U209 ( .A(n977), .ZN(n696) );
  AOI22_X1 U210 ( .A1(data_in[3]), .A2(n829), .B1(n980), .B2(\mem[14][3] ), 
        .ZN(n977) );
  INV_X1 U211 ( .A(n976), .ZN(n695) );
  AOI22_X1 U212 ( .A1(data_in[4]), .A2(n829), .B1(n980), .B2(\mem[14][4] ), 
        .ZN(n976) );
  INV_X1 U213 ( .A(n975), .ZN(n694) );
  AOI22_X1 U214 ( .A1(data_in[5]), .A2(n829), .B1(n980), .B2(\mem[14][5] ), 
        .ZN(n975) );
  INV_X1 U215 ( .A(n974), .ZN(n693) );
  AOI22_X1 U216 ( .A1(data_in[6]), .A2(n829), .B1(n980), .B2(\mem[14][6] ), 
        .ZN(n974) );
  INV_X1 U217 ( .A(n973), .ZN(n692) );
  AOI22_X1 U218 ( .A1(data_in[7]), .A2(n829), .B1(n980), .B2(\mem[14][7] ), 
        .ZN(n973) );
  INV_X1 U219 ( .A(n972), .ZN(n691) );
  AOI22_X1 U220 ( .A1(data_in[0]), .A2(n828), .B1(n971), .B2(\mem[15][0] ), 
        .ZN(n972) );
  INV_X1 U221 ( .A(n970), .ZN(n690) );
  AOI22_X1 U222 ( .A1(data_in[1]), .A2(n828), .B1(n971), .B2(\mem[15][1] ), 
        .ZN(n970) );
  INV_X1 U223 ( .A(n969), .ZN(n689) );
  AOI22_X1 U224 ( .A1(data_in[2]), .A2(n828), .B1(n971), .B2(\mem[15][2] ), 
        .ZN(n969) );
  INV_X1 U225 ( .A(n968), .ZN(n688) );
  AOI22_X1 U226 ( .A1(data_in[3]), .A2(n828), .B1(n971), .B2(\mem[15][3] ), 
        .ZN(n968) );
  INV_X1 U227 ( .A(n967), .ZN(n687) );
  AOI22_X1 U228 ( .A1(data_in[4]), .A2(n828), .B1(n971), .B2(\mem[15][4] ), 
        .ZN(n967) );
  INV_X1 U229 ( .A(n966), .ZN(n686) );
  AOI22_X1 U230 ( .A1(data_in[5]), .A2(n828), .B1(n971), .B2(\mem[15][5] ), 
        .ZN(n966) );
  INV_X1 U231 ( .A(n965), .ZN(n685) );
  AOI22_X1 U232 ( .A1(data_in[6]), .A2(n828), .B1(n971), .B2(\mem[15][6] ), 
        .ZN(n965) );
  INV_X1 U233 ( .A(n964), .ZN(n684) );
  AOI22_X1 U234 ( .A1(data_in[7]), .A2(n828), .B1(n971), .B2(\mem[15][7] ), 
        .ZN(n964) );
  INV_X1 U235 ( .A(n944), .ZN(n667) );
  AOI22_X1 U236 ( .A1(data_in[0]), .A2(n825), .B1(n943), .B2(\mem[18][0] ), 
        .ZN(n944) );
  INV_X1 U237 ( .A(n942), .ZN(n666) );
  AOI22_X1 U238 ( .A1(data_in[1]), .A2(n825), .B1(n943), .B2(\mem[18][1] ), 
        .ZN(n942) );
  INV_X1 U239 ( .A(n941), .ZN(n665) );
  AOI22_X1 U240 ( .A1(data_in[2]), .A2(n825), .B1(n943), .B2(\mem[18][2] ), 
        .ZN(n941) );
  INV_X1 U241 ( .A(n940), .ZN(n664) );
  AOI22_X1 U242 ( .A1(data_in[3]), .A2(n825), .B1(n943), .B2(\mem[18][3] ), 
        .ZN(n940) );
  INV_X1 U243 ( .A(n939), .ZN(n663) );
  AOI22_X1 U244 ( .A1(data_in[4]), .A2(n825), .B1(n943), .B2(\mem[18][4] ), 
        .ZN(n939) );
  INV_X1 U245 ( .A(n938), .ZN(n662) );
  AOI22_X1 U246 ( .A1(data_in[5]), .A2(n825), .B1(n943), .B2(\mem[18][5] ), 
        .ZN(n938) );
  INV_X1 U247 ( .A(n937), .ZN(n661) );
  AOI22_X1 U248 ( .A1(data_in[6]), .A2(n825), .B1(n943), .B2(\mem[18][6] ), 
        .ZN(n937) );
  INV_X1 U249 ( .A(n936), .ZN(n660) );
  AOI22_X1 U250 ( .A1(data_in[7]), .A2(n825), .B1(n943), .B2(\mem[18][7] ), 
        .ZN(n936) );
  INV_X1 U251 ( .A(n935), .ZN(n659) );
  AOI22_X1 U252 ( .A1(data_in[0]), .A2(n824), .B1(n934), .B2(\mem[19][0] ), 
        .ZN(n935) );
  INV_X1 U253 ( .A(n933), .ZN(n658) );
  AOI22_X1 U254 ( .A1(data_in[1]), .A2(n824), .B1(n934), .B2(\mem[19][1] ), 
        .ZN(n933) );
  INV_X1 U255 ( .A(n932), .ZN(n657) );
  AOI22_X1 U256 ( .A1(data_in[2]), .A2(n824), .B1(n934), .B2(\mem[19][2] ), 
        .ZN(n932) );
  INV_X1 U257 ( .A(n931), .ZN(n656) );
  AOI22_X1 U258 ( .A1(data_in[3]), .A2(n824), .B1(n934), .B2(\mem[19][3] ), 
        .ZN(n931) );
  INV_X1 U259 ( .A(n930), .ZN(n655) );
  AOI22_X1 U260 ( .A1(data_in[4]), .A2(n824), .B1(n934), .B2(\mem[19][4] ), 
        .ZN(n930) );
  INV_X1 U261 ( .A(n929), .ZN(n654) );
  AOI22_X1 U262 ( .A1(data_in[5]), .A2(n824), .B1(n934), .B2(\mem[19][5] ), 
        .ZN(n929) );
  INV_X1 U263 ( .A(n928), .ZN(n653) );
  AOI22_X1 U264 ( .A1(data_in[6]), .A2(n824), .B1(n934), .B2(\mem[19][6] ), 
        .ZN(n928) );
  INV_X1 U265 ( .A(n927), .ZN(n652) );
  AOI22_X1 U266 ( .A1(data_in[7]), .A2(n824), .B1(n934), .B2(\mem[19][7] ), 
        .ZN(n927) );
  INV_X1 U267 ( .A(n908), .ZN(n635) );
  AOI22_X1 U268 ( .A1(data_in[0]), .A2(n821), .B1(n907), .B2(\mem[22][0] ), 
        .ZN(n908) );
  INV_X1 U269 ( .A(n906), .ZN(n634) );
  AOI22_X1 U270 ( .A1(data_in[1]), .A2(n821), .B1(n907), .B2(\mem[22][1] ), 
        .ZN(n906) );
  INV_X1 U271 ( .A(n905), .ZN(n633) );
  AOI22_X1 U272 ( .A1(data_in[2]), .A2(n821), .B1(n907), .B2(\mem[22][2] ), 
        .ZN(n905) );
  INV_X1 U273 ( .A(n904), .ZN(n632) );
  AOI22_X1 U274 ( .A1(data_in[3]), .A2(n821), .B1(n907), .B2(\mem[22][3] ), 
        .ZN(n904) );
  INV_X1 U275 ( .A(n903), .ZN(n631) );
  AOI22_X1 U276 ( .A1(data_in[4]), .A2(n821), .B1(n907), .B2(\mem[22][4] ), 
        .ZN(n903) );
  INV_X1 U277 ( .A(n902), .ZN(n630) );
  AOI22_X1 U278 ( .A1(data_in[5]), .A2(n821), .B1(n907), .B2(\mem[22][5] ), 
        .ZN(n902) );
  INV_X1 U279 ( .A(n901), .ZN(n629) );
  AOI22_X1 U280 ( .A1(data_in[6]), .A2(n821), .B1(n907), .B2(\mem[22][6] ), 
        .ZN(n901) );
  INV_X1 U281 ( .A(n900), .ZN(n628) );
  AOI22_X1 U282 ( .A1(data_in[7]), .A2(n821), .B1(n907), .B2(\mem[22][7] ), 
        .ZN(n900) );
  INV_X1 U283 ( .A(n899), .ZN(n627) );
  AOI22_X1 U284 ( .A1(data_in[0]), .A2(n820), .B1(n898), .B2(\mem[23][0] ), 
        .ZN(n899) );
  INV_X1 U285 ( .A(n897), .ZN(n626) );
  AOI22_X1 U286 ( .A1(data_in[1]), .A2(n820), .B1(n898), .B2(\mem[23][1] ), 
        .ZN(n897) );
  INV_X1 U287 ( .A(n896), .ZN(n625) );
  AOI22_X1 U288 ( .A1(data_in[2]), .A2(n820), .B1(n898), .B2(\mem[23][2] ), 
        .ZN(n896) );
  INV_X1 U289 ( .A(n895), .ZN(n624) );
  AOI22_X1 U290 ( .A1(data_in[3]), .A2(n820), .B1(n898), .B2(\mem[23][3] ), 
        .ZN(n895) );
  INV_X1 U291 ( .A(n894), .ZN(n623) );
  AOI22_X1 U292 ( .A1(data_in[4]), .A2(n820), .B1(n898), .B2(\mem[23][4] ), 
        .ZN(n894) );
  INV_X1 U293 ( .A(n893), .ZN(n622) );
  AOI22_X1 U294 ( .A1(data_in[5]), .A2(n820), .B1(n898), .B2(\mem[23][5] ), 
        .ZN(n893) );
  INV_X1 U295 ( .A(n892), .ZN(n621) );
  AOI22_X1 U296 ( .A1(data_in[6]), .A2(n820), .B1(n898), .B2(\mem[23][6] ), 
        .ZN(n892) );
  INV_X1 U297 ( .A(n891), .ZN(n620) );
  AOI22_X1 U298 ( .A1(data_in[7]), .A2(n820), .B1(n898), .B2(\mem[23][7] ), 
        .ZN(n891) );
  INV_X1 U299 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U300 ( .A1(data_in[0]), .A2(n837), .B1(n1053), .B2(\mem[6][0] ), 
        .ZN(n1054) );
  INV_X1 U301 ( .A(n1052), .ZN(n762) );
  AOI22_X1 U302 ( .A1(data_in[1]), .A2(n837), .B1(n1053), .B2(\mem[6][1] ), 
        .ZN(n1052) );
  INV_X1 U303 ( .A(n1051), .ZN(n761) );
  AOI22_X1 U304 ( .A1(data_in[2]), .A2(n837), .B1(n1053), .B2(\mem[6][2] ), 
        .ZN(n1051) );
  INV_X1 U305 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U306 ( .A1(data_in[3]), .A2(n837), .B1(n1053), .B2(\mem[6][3] ), 
        .ZN(n1050) );
  INV_X1 U307 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U308 ( .A1(data_in[4]), .A2(n837), .B1(n1053), .B2(\mem[6][4] ), 
        .ZN(n1049) );
  INV_X1 U309 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U310 ( .A1(data_in[5]), .A2(n837), .B1(n1053), .B2(\mem[6][5] ), 
        .ZN(n1048) );
  INV_X1 U311 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U312 ( .A1(data_in[6]), .A2(n837), .B1(n1053), .B2(\mem[6][6] ), 
        .ZN(n1047) );
  INV_X1 U313 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U314 ( .A1(data_in[7]), .A2(n837), .B1(n1053), .B2(\mem[6][7] ), 
        .ZN(n1046) );
  INV_X1 U315 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U316 ( .A1(data_in[0]), .A2(n836), .B1(n1044), .B2(\mem[7][0] ), 
        .ZN(n1045) );
  INV_X1 U317 ( .A(n1043), .ZN(n754) );
  AOI22_X1 U318 ( .A1(data_in[1]), .A2(n836), .B1(n1044), .B2(\mem[7][1] ), 
        .ZN(n1043) );
  INV_X1 U319 ( .A(n1042), .ZN(n753) );
  AOI22_X1 U320 ( .A1(data_in[2]), .A2(n836), .B1(n1044), .B2(\mem[7][2] ), 
        .ZN(n1042) );
  INV_X1 U321 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U322 ( .A1(data_in[3]), .A2(n836), .B1(n1044), .B2(\mem[7][3] ), 
        .ZN(n1041) );
  INV_X1 U323 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U324 ( .A1(data_in[4]), .A2(n836), .B1(n1044), .B2(\mem[7][4] ), 
        .ZN(n1040) );
  INV_X1 U325 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U326 ( .A1(data_in[5]), .A2(n836), .B1(n1044), .B2(\mem[7][5] ), 
        .ZN(n1039) );
  INV_X1 U327 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U328 ( .A1(data_in[6]), .A2(n836), .B1(n1044), .B2(\mem[7][6] ), 
        .ZN(n1038) );
  INV_X1 U329 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U330 ( .A1(data_in[7]), .A2(n836), .B1(n1044), .B2(\mem[7][7] ), 
        .ZN(n1037) );
  INV_X1 U331 ( .A(N12), .ZN(n255) );
  INV_X1 U332 ( .A(N11), .ZN(n254) );
  INV_X1 U333 ( .A(n999), .ZN(n715) );
  AOI22_X1 U334 ( .A1(data_in[0]), .A2(n831), .B1(n998), .B2(\mem[12][0] ), 
        .ZN(n999) );
  INV_X1 U335 ( .A(n997), .ZN(n714) );
  AOI22_X1 U336 ( .A1(data_in[1]), .A2(n831), .B1(n998), .B2(\mem[12][1] ), 
        .ZN(n997) );
  INV_X1 U337 ( .A(n996), .ZN(n713) );
  AOI22_X1 U338 ( .A1(data_in[2]), .A2(n831), .B1(n998), .B2(\mem[12][2] ), 
        .ZN(n996) );
  INV_X1 U339 ( .A(n995), .ZN(n712) );
  AOI22_X1 U340 ( .A1(data_in[3]), .A2(n831), .B1(n998), .B2(\mem[12][3] ), 
        .ZN(n995) );
  INV_X1 U341 ( .A(n994), .ZN(n711) );
  AOI22_X1 U342 ( .A1(data_in[4]), .A2(n831), .B1(n998), .B2(\mem[12][4] ), 
        .ZN(n994) );
  INV_X1 U343 ( .A(n993), .ZN(n710) );
  AOI22_X1 U344 ( .A1(data_in[5]), .A2(n831), .B1(n998), .B2(\mem[12][5] ), 
        .ZN(n993) );
  INV_X1 U345 ( .A(n992), .ZN(n709) );
  AOI22_X1 U346 ( .A1(data_in[6]), .A2(n831), .B1(n998), .B2(\mem[12][6] ), 
        .ZN(n992) );
  INV_X1 U347 ( .A(n991), .ZN(n708) );
  AOI22_X1 U348 ( .A1(data_in[7]), .A2(n831), .B1(n998), .B2(\mem[12][7] ), 
        .ZN(n991) );
  INV_X1 U349 ( .A(n926), .ZN(n651) );
  AOI22_X1 U350 ( .A1(data_in[0]), .A2(n823), .B1(n925), .B2(\mem[20][0] ), 
        .ZN(n926) );
  INV_X1 U351 ( .A(n924), .ZN(n650) );
  AOI22_X1 U352 ( .A1(data_in[1]), .A2(n823), .B1(n925), .B2(\mem[20][1] ), 
        .ZN(n924) );
  INV_X1 U353 ( .A(n923), .ZN(n649) );
  AOI22_X1 U354 ( .A1(data_in[2]), .A2(n823), .B1(n925), .B2(\mem[20][2] ), 
        .ZN(n923) );
  INV_X1 U355 ( .A(n922), .ZN(n648) );
  AOI22_X1 U356 ( .A1(data_in[3]), .A2(n823), .B1(n925), .B2(\mem[20][3] ), 
        .ZN(n922) );
  INV_X1 U357 ( .A(n921), .ZN(n647) );
  AOI22_X1 U358 ( .A1(data_in[4]), .A2(n823), .B1(n925), .B2(\mem[20][4] ), 
        .ZN(n921) );
  INV_X1 U359 ( .A(n920), .ZN(n646) );
  AOI22_X1 U360 ( .A1(data_in[5]), .A2(n823), .B1(n925), .B2(\mem[20][5] ), 
        .ZN(n920) );
  INV_X1 U361 ( .A(n919), .ZN(n645) );
  AOI22_X1 U362 ( .A1(data_in[6]), .A2(n823), .B1(n925), .B2(\mem[20][6] ), 
        .ZN(n919) );
  INV_X1 U363 ( .A(n918), .ZN(n644) );
  AOI22_X1 U364 ( .A1(data_in[7]), .A2(n823), .B1(n925), .B2(\mem[20][7] ), 
        .ZN(n918) );
  INV_X1 U365 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U366 ( .A1(data_in[0]), .A2(n835), .B1(n1035), .B2(\mem[8][0] ), 
        .ZN(n1036) );
  INV_X1 U367 ( .A(n1034), .ZN(n746) );
  AOI22_X1 U368 ( .A1(data_in[1]), .A2(n835), .B1(n1035), .B2(\mem[8][1] ), 
        .ZN(n1034) );
  INV_X1 U369 ( .A(n1033), .ZN(n745) );
  AOI22_X1 U370 ( .A1(data_in[2]), .A2(n835), .B1(n1035), .B2(\mem[8][2] ), 
        .ZN(n1033) );
  INV_X1 U371 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U372 ( .A1(data_in[3]), .A2(n835), .B1(n1035), .B2(\mem[8][3] ), 
        .ZN(n1032) );
  INV_X1 U373 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U374 ( .A1(data_in[4]), .A2(n835), .B1(n1035), .B2(\mem[8][4] ), 
        .ZN(n1031) );
  INV_X1 U375 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U376 ( .A1(data_in[5]), .A2(n835), .B1(n1035), .B2(\mem[8][5] ), 
        .ZN(n1030) );
  INV_X1 U377 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U378 ( .A1(data_in[6]), .A2(n835), .B1(n1035), .B2(\mem[8][6] ), 
        .ZN(n1029) );
  INV_X1 U379 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U380 ( .A1(data_in[7]), .A2(n835), .B1(n1035), .B2(\mem[8][7] ), 
        .ZN(n1028) );
  INV_X1 U381 ( .A(n963), .ZN(n683) );
  AOI22_X1 U382 ( .A1(data_in[0]), .A2(n827), .B1(n962), .B2(\mem[16][0] ), 
        .ZN(n963) );
  INV_X1 U383 ( .A(n961), .ZN(n682) );
  AOI22_X1 U384 ( .A1(data_in[1]), .A2(n827), .B1(n962), .B2(\mem[16][1] ), 
        .ZN(n961) );
  INV_X1 U385 ( .A(n960), .ZN(n681) );
  AOI22_X1 U386 ( .A1(data_in[2]), .A2(n827), .B1(n962), .B2(\mem[16][2] ), 
        .ZN(n960) );
  INV_X1 U387 ( .A(n959), .ZN(n680) );
  AOI22_X1 U388 ( .A1(data_in[3]), .A2(n827), .B1(n962), .B2(\mem[16][3] ), 
        .ZN(n959) );
  INV_X1 U389 ( .A(n958), .ZN(n679) );
  AOI22_X1 U390 ( .A1(data_in[4]), .A2(n827), .B1(n962), .B2(\mem[16][4] ), 
        .ZN(n958) );
  INV_X1 U391 ( .A(n957), .ZN(n678) );
  AOI22_X1 U392 ( .A1(data_in[5]), .A2(n827), .B1(n962), .B2(\mem[16][5] ), 
        .ZN(n957) );
  INV_X1 U393 ( .A(n956), .ZN(n677) );
  AOI22_X1 U394 ( .A1(data_in[6]), .A2(n827), .B1(n962), .B2(\mem[16][6] ), 
        .ZN(n956) );
  INV_X1 U395 ( .A(n955), .ZN(n676) );
  AOI22_X1 U396 ( .A1(data_in[7]), .A2(n827), .B1(n962), .B2(\mem[16][7] ), 
        .ZN(n955) );
  INV_X1 U397 ( .A(n890), .ZN(n619) );
  AOI22_X1 U398 ( .A1(data_in[0]), .A2(n816), .B1(n889), .B2(\mem[24][0] ), 
        .ZN(n890) );
  INV_X1 U399 ( .A(n888), .ZN(n618) );
  AOI22_X1 U400 ( .A1(data_in[1]), .A2(n816), .B1(n889), .B2(\mem[24][1] ), 
        .ZN(n888) );
  INV_X1 U401 ( .A(n887), .ZN(n617) );
  AOI22_X1 U402 ( .A1(data_in[2]), .A2(n816), .B1(n889), .B2(\mem[24][2] ), 
        .ZN(n887) );
  INV_X1 U403 ( .A(n886), .ZN(n616) );
  AOI22_X1 U404 ( .A1(data_in[3]), .A2(n816), .B1(n889), .B2(\mem[24][3] ), 
        .ZN(n886) );
  INV_X1 U405 ( .A(n885), .ZN(n615) );
  AOI22_X1 U406 ( .A1(data_in[4]), .A2(n816), .B1(n889), .B2(\mem[24][4] ), 
        .ZN(n885) );
  INV_X1 U407 ( .A(n884), .ZN(n614) );
  AOI22_X1 U408 ( .A1(data_in[5]), .A2(n816), .B1(n889), .B2(\mem[24][5] ), 
        .ZN(n884) );
  INV_X1 U409 ( .A(n883), .ZN(n613) );
  AOI22_X1 U410 ( .A1(data_in[6]), .A2(n816), .B1(n889), .B2(\mem[24][6] ), 
        .ZN(n883) );
  INV_X1 U411 ( .A(n882), .ZN(n612) );
  AOI22_X1 U412 ( .A1(data_in[7]), .A2(n816), .B1(n889), .B2(\mem[24][7] ), 
        .ZN(n882) );
  INV_X1 U413 ( .A(n881), .ZN(n611) );
  AOI22_X1 U414 ( .A1(data_in[0]), .A2(n815), .B1(n880), .B2(\mem[25][0] ), 
        .ZN(n881) );
  INV_X1 U415 ( .A(n879), .ZN(n610) );
  AOI22_X1 U416 ( .A1(data_in[1]), .A2(n815), .B1(n880), .B2(\mem[25][1] ), 
        .ZN(n879) );
  INV_X1 U417 ( .A(n878), .ZN(n609) );
  AOI22_X1 U418 ( .A1(data_in[2]), .A2(n815), .B1(n880), .B2(\mem[25][2] ), 
        .ZN(n878) );
  INV_X1 U419 ( .A(n877), .ZN(n608) );
  AOI22_X1 U420 ( .A1(data_in[3]), .A2(n815), .B1(n880), .B2(\mem[25][3] ), 
        .ZN(n877) );
  INV_X1 U421 ( .A(n876), .ZN(n607) );
  AOI22_X1 U422 ( .A1(data_in[4]), .A2(n815), .B1(n880), .B2(\mem[25][4] ), 
        .ZN(n876) );
  INV_X1 U423 ( .A(n875), .ZN(n606) );
  AOI22_X1 U424 ( .A1(data_in[5]), .A2(n815), .B1(n880), .B2(\mem[25][5] ), 
        .ZN(n875) );
  INV_X1 U425 ( .A(n874), .ZN(n605) );
  AOI22_X1 U426 ( .A1(data_in[6]), .A2(n815), .B1(n880), .B2(\mem[25][6] ), 
        .ZN(n874) );
  INV_X1 U427 ( .A(n873), .ZN(n604) );
  AOI22_X1 U428 ( .A1(data_in[7]), .A2(n815), .B1(n880), .B2(\mem[25][7] ), 
        .ZN(n873) );
  INV_X1 U429 ( .A(n872), .ZN(n603) );
  AOI22_X1 U430 ( .A1(data_in[0]), .A2(n814), .B1(n871), .B2(\mem[26][0] ), 
        .ZN(n872) );
  INV_X1 U431 ( .A(n870), .ZN(n602) );
  AOI22_X1 U432 ( .A1(data_in[1]), .A2(n814), .B1(n871), .B2(\mem[26][1] ), 
        .ZN(n870) );
  INV_X1 U433 ( .A(n869), .ZN(n601) );
  AOI22_X1 U434 ( .A1(data_in[2]), .A2(n814), .B1(n871), .B2(\mem[26][2] ), 
        .ZN(n869) );
  INV_X1 U435 ( .A(n868), .ZN(n600) );
  AOI22_X1 U436 ( .A1(data_in[3]), .A2(n814), .B1(n871), .B2(\mem[26][3] ), 
        .ZN(n868) );
  INV_X1 U437 ( .A(n867), .ZN(n599) );
  AOI22_X1 U438 ( .A1(data_in[4]), .A2(n814), .B1(n871), .B2(\mem[26][4] ), 
        .ZN(n867) );
  INV_X1 U439 ( .A(n866), .ZN(n598) );
  AOI22_X1 U440 ( .A1(data_in[5]), .A2(n814), .B1(n871), .B2(\mem[26][5] ), 
        .ZN(n866) );
  INV_X1 U441 ( .A(n865), .ZN(n597) );
  AOI22_X1 U442 ( .A1(data_in[6]), .A2(n814), .B1(n871), .B2(\mem[26][6] ), 
        .ZN(n865) );
  INV_X1 U443 ( .A(n864), .ZN(n596) );
  AOI22_X1 U444 ( .A1(data_in[7]), .A2(n814), .B1(n871), .B2(\mem[26][7] ), 
        .ZN(n864) );
  INV_X1 U445 ( .A(n863), .ZN(n595) );
  AOI22_X1 U446 ( .A1(data_in[0]), .A2(n813), .B1(n862), .B2(\mem[27][0] ), 
        .ZN(n863) );
  INV_X1 U447 ( .A(n861), .ZN(n594) );
  AOI22_X1 U448 ( .A1(data_in[1]), .A2(n813), .B1(n862), .B2(\mem[27][1] ), 
        .ZN(n861) );
  INV_X1 U449 ( .A(n860), .ZN(n293) );
  AOI22_X1 U450 ( .A1(data_in[2]), .A2(n813), .B1(n862), .B2(\mem[27][2] ), 
        .ZN(n860) );
  INV_X1 U451 ( .A(n859), .ZN(n292) );
  AOI22_X1 U452 ( .A1(data_in[3]), .A2(n813), .B1(n862), .B2(\mem[27][3] ), 
        .ZN(n859) );
  INV_X1 U453 ( .A(n858), .ZN(n291) );
  AOI22_X1 U454 ( .A1(data_in[4]), .A2(n813), .B1(n862), .B2(\mem[27][4] ), 
        .ZN(n858) );
  INV_X1 U455 ( .A(n857), .ZN(n290) );
  AOI22_X1 U456 ( .A1(data_in[5]), .A2(n813), .B1(n862), .B2(\mem[27][5] ), 
        .ZN(n857) );
  INV_X1 U457 ( .A(n856), .ZN(n289) );
  AOI22_X1 U458 ( .A1(data_in[6]), .A2(n813), .B1(n862), .B2(\mem[27][6] ), 
        .ZN(n856) );
  INV_X1 U459 ( .A(n855), .ZN(n288) );
  AOI22_X1 U460 ( .A1(data_in[7]), .A2(n813), .B1(n862), .B2(\mem[27][7] ), 
        .ZN(n855) );
  INV_X1 U461 ( .A(n854), .ZN(n287) );
  AOI22_X1 U462 ( .A1(data_in[0]), .A2(n812), .B1(n853), .B2(\mem[28][0] ), 
        .ZN(n854) );
  INV_X1 U463 ( .A(n852), .ZN(n286) );
  AOI22_X1 U464 ( .A1(data_in[1]), .A2(n812), .B1(n853), .B2(\mem[28][1] ), 
        .ZN(n852) );
  INV_X1 U465 ( .A(n851), .ZN(n285) );
  AOI22_X1 U466 ( .A1(data_in[2]), .A2(n812), .B1(n853), .B2(\mem[28][2] ), 
        .ZN(n851) );
  INV_X1 U467 ( .A(n850), .ZN(n284) );
  AOI22_X1 U468 ( .A1(data_in[3]), .A2(n812), .B1(n853), .B2(\mem[28][3] ), 
        .ZN(n850) );
  INV_X1 U469 ( .A(n849), .ZN(n283) );
  AOI22_X1 U470 ( .A1(data_in[4]), .A2(n812), .B1(n853), .B2(\mem[28][4] ), 
        .ZN(n849) );
  INV_X1 U471 ( .A(n848), .ZN(n282) );
  AOI22_X1 U472 ( .A1(data_in[5]), .A2(n812), .B1(n853), .B2(\mem[28][5] ), 
        .ZN(n848) );
  INV_X1 U473 ( .A(n847), .ZN(n281) );
  AOI22_X1 U474 ( .A1(data_in[6]), .A2(n812), .B1(n853), .B2(\mem[28][6] ), 
        .ZN(n847) );
  INV_X1 U475 ( .A(n846), .ZN(n280) );
  AOI22_X1 U476 ( .A1(data_in[7]), .A2(n812), .B1(n853), .B2(\mem[28][7] ), 
        .ZN(n846) );
  INV_X1 U477 ( .A(n1145), .ZN(n279) );
  AOI22_X1 U478 ( .A1(n819), .A2(data_in[0]), .B1(n1144), .B2(\mem[29][0] ), 
        .ZN(n1145) );
  INV_X1 U479 ( .A(n1143), .ZN(n278) );
  AOI22_X1 U480 ( .A1(n819), .A2(data_in[1]), .B1(n1144), .B2(\mem[29][1] ), 
        .ZN(n1143) );
  INV_X1 U481 ( .A(n1142), .ZN(n277) );
  AOI22_X1 U482 ( .A1(n819), .A2(data_in[2]), .B1(n1144), .B2(\mem[29][2] ), 
        .ZN(n1142) );
  INV_X1 U483 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U484 ( .A1(n819), .A2(data_in[3]), .B1(n1144), .B2(\mem[29][3] ), 
        .ZN(n1141) );
  INV_X1 U485 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U486 ( .A1(n819), .A2(data_in[4]), .B1(n1144), .B2(\mem[29][4] ), 
        .ZN(n1140) );
  INV_X1 U487 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U488 ( .A1(n819), .A2(data_in[5]), .B1(n1144), .B2(\mem[29][5] ), 
        .ZN(n1139) );
  INV_X1 U489 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U490 ( .A1(n819), .A2(data_in[6]), .B1(n1144), .B2(\mem[29][6] ), 
        .ZN(n1138) );
  INV_X1 U491 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U492 ( .A1(n819), .A2(data_in[7]), .B1(n1144), .B2(\mem[29][7] ), 
        .ZN(n1137) );
  INV_X1 U493 ( .A(n1134), .ZN(n271) );
  AOI22_X1 U494 ( .A1(data_in[0]), .A2(n818), .B1(n1133), .B2(\mem[30][0] ), 
        .ZN(n1134) );
  INV_X1 U495 ( .A(n1132), .ZN(n270) );
  AOI22_X1 U496 ( .A1(data_in[1]), .A2(n818), .B1(n1133), .B2(\mem[30][1] ), 
        .ZN(n1132) );
  INV_X1 U497 ( .A(n1131), .ZN(n269) );
  AOI22_X1 U498 ( .A1(data_in[2]), .A2(n818), .B1(n1133), .B2(\mem[30][2] ), 
        .ZN(n1131) );
  INV_X1 U499 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U500 ( .A1(data_in[3]), .A2(n818), .B1(n1133), .B2(\mem[30][3] ), 
        .ZN(n1130) );
  INV_X1 U501 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U502 ( .A1(data_in[4]), .A2(n818), .B1(n1133), .B2(\mem[30][4] ), 
        .ZN(n1129) );
  INV_X1 U503 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U504 ( .A1(data_in[5]), .A2(n818), .B1(n1133), .B2(\mem[30][5] ), 
        .ZN(n1128) );
  INV_X1 U505 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U506 ( .A1(data_in[6]), .A2(n818), .B1(n1133), .B2(\mem[30][6] ), 
        .ZN(n1127) );
  INV_X1 U507 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U508 ( .A1(data_in[7]), .A2(n818), .B1(n1133), .B2(\mem[30][7] ), 
        .ZN(n1126) );
  INV_X1 U509 ( .A(n1124), .ZN(n263) );
  AOI22_X1 U510 ( .A1(data_in[0]), .A2(n817), .B1(n1123), .B2(\mem[31][0] ), 
        .ZN(n1124) );
  INV_X1 U511 ( .A(n1122), .ZN(n262) );
  AOI22_X1 U512 ( .A1(data_in[1]), .A2(n817), .B1(n1123), .B2(\mem[31][1] ), 
        .ZN(n1122) );
  INV_X1 U513 ( .A(n1121), .ZN(n261) );
  AOI22_X1 U514 ( .A1(data_in[2]), .A2(n817), .B1(n1123), .B2(\mem[31][2] ), 
        .ZN(n1121) );
  INV_X1 U515 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U516 ( .A1(data_in[3]), .A2(n817), .B1(n1123), .B2(\mem[31][3] ), 
        .ZN(n1120) );
  INV_X1 U517 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U518 ( .A1(data_in[4]), .A2(n817), .B1(n1123), .B2(\mem[31][4] ), 
        .ZN(n1119) );
  INV_X1 U519 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U520 ( .A1(data_in[5]), .A2(n817), .B1(n1123), .B2(\mem[31][5] ), 
        .ZN(n1118) );
  INV_X1 U521 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U522 ( .A1(data_in[6]), .A2(n817), .B1(n1123), .B2(\mem[31][6] ), 
        .ZN(n1117) );
  INV_X1 U523 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U524 ( .A1(data_in[7]), .A2(n817), .B1(n1123), .B2(\mem[31][7] ), 
        .ZN(n1116) );
  INV_X1 U525 ( .A(n1114), .ZN(n811) );
  AOI22_X1 U526 ( .A1(data_in[0]), .A2(n843), .B1(n1113), .B2(\mem[0][0] ), 
        .ZN(n1114) );
  INV_X1 U527 ( .A(n1112), .ZN(n810) );
  AOI22_X1 U528 ( .A1(data_in[1]), .A2(n843), .B1(n1113), .B2(\mem[0][1] ), 
        .ZN(n1112) );
  INV_X1 U529 ( .A(n1111), .ZN(n809) );
  AOI22_X1 U530 ( .A1(data_in[2]), .A2(n843), .B1(n1113), .B2(\mem[0][2] ), 
        .ZN(n1111) );
  INV_X1 U531 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U532 ( .A1(data_in[3]), .A2(n843), .B1(n1113), .B2(\mem[0][3] ), 
        .ZN(n1110) );
  INV_X1 U533 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U534 ( .A1(data_in[4]), .A2(n843), .B1(n1113), .B2(\mem[0][4] ), 
        .ZN(n1109) );
  INV_X1 U535 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U536 ( .A1(data_in[5]), .A2(n843), .B1(n1113), .B2(\mem[0][5] ), 
        .ZN(n1108) );
  INV_X1 U537 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U538 ( .A1(data_in[6]), .A2(n843), .B1(n1113), .B2(\mem[0][6] ), 
        .ZN(n1107) );
  INV_X1 U539 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U540 ( .A1(data_in[7]), .A2(n843), .B1(n1113), .B2(\mem[0][7] ), 
        .ZN(n1106) );
  INV_X1 U541 ( .A(n1103), .ZN(n803) );
  AOI22_X1 U542 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[1][0] ), 
        .ZN(n1103) );
  INV_X1 U543 ( .A(n1101), .ZN(n802) );
  AOI22_X1 U544 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[1][1] ), 
        .ZN(n1101) );
  INV_X1 U545 ( .A(n1100), .ZN(n801) );
  AOI22_X1 U546 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[1][2] ), 
        .ZN(n1100) );
  INV_X1 U547 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U548 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[1][3] ), 
        .ZN(n1099) );
  INV_X1 U549 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U550 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[1][4] ), 
        .ZN(n1098) );
  INV_X1 U551 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U552 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[1][5] ), 
        .ZN(n1097) );
  INV_X1 U553 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U554 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[1][6] ), 
        .ZN(n1096) );
  INV_X1 U555 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U556 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[1][7] ), 
        .ZN(n1095) );
  INV_X1 U557 ( .A(n1093), .ZN(n795) );
  AOI22_X1 U558 ( .A1(data_in[0]), .A2(n841), .B1(n1092), .B2(\mem[2][0] ), 
        .ZN(n1093) );
  INV_X1 U559 ( .A(n1091), .ZN(n794) );
  AOI22_X1 U560 ( .A1(data_in[1]), .A2(n841), .B1(n1092), .B2(\mem[2][1] ), 
        .ZN(n1091) );
  INV_X1 U561 ( .A(n1090), .ZN(n793) );
  AOI22_X1 U562 ( .A1(data_in[2]), .A2(n841), .B1(n1092), .B2(\mem[2][2] ), 
        .ZN(n1090) );
  INV_X1 U563 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U564 ( .A1(data_in[3]), .A2(n841), .B1(n1092), .B2(\mem[2][3] ), 
        .ZN(n1089) );
  INV_X1 U565 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U566 ( .A1(data_in[4]), .A2(n841), .B1(n1092), .B2(\mem[2][4] ), 
        .ZN(n1088) );
  INV_X1 U567 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U568 ( .A1(data_in[5]), .A2(n841), .B1(n1092), .B2(\mem[2][5] ), 
        .ZN(n1087) );
  INV_X1 U569 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U570 ( .A1(data_in[6]), .A2(n841), .B1(n1092), .B2(\mem[2][6] ), 
        .ZN(n1086) );
  INV_X1 U571 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U572 ( .A1(data_in[7]), .A2(n841), .B1(n1092), .B2(\mem[2][7] ), 
        .ZN(n1085) );
  INV_X1 U573 ( .A(n1083), .ZN(n787) );
  AOI22_X1 U574 ( .A1(data_in[0]), .A2(n840), .B1(n1082), .B2(\mem[3][0] ), 
        .ZN(n1083) );
  INV_X1 U575 ( .A(n1081), .ZN(n786) );
  AOI22_X1 U576 ( .A1(data_in[1]), .A2(n840), .B1(n1082), .B2(\mem[3][1] ), 
        .ZN(n1081) );
  INV_X1 U577 ( .A(n1080), .ZN(n785) );
  AOI22_X1 U578 ( .A1(data_in[2]), .A2(n840), .B1(n1082), .B2(\mem[3][2] ), 
        .ZN(n1080) );
  INV_X1 U579 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U580 ( .A1(data_in[3]), .A2(n840), .B1(n1082), .B2(\mem[3][3] ), 
        .ZN(n1079) );
  INV_X1 U581 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U582 ( .A1(data_in[4]), .A2(n840), .B1(n1082), .B2(\mem[3][4] ), 
        .ZN(n1078) );
  INV_X1 U583 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U584 ( .A1(data_in[5]), .A2(n840), .B1(n1082), .B2(\mem[3][5] ), 
        .ZN(n1077) );
  INV_X1 U585 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U586 ( .A1(data_in[6]), .A2(n840), .B1(n1082), .B2(\mem[3][6] ), 
        .ZN(n1076) );
  INV_X1 U587 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U588 ( .A1(data_in[7]), .A2(n840), .B1(n1082), .B2(\mem[3][7] ), 
        .ZN(n1075) );
  INV_X1 U589 ( .A(n1073), .ZN(n779) );
  AOI22_X1 U590 ( .A1(data_in[0]), .A2(n839), .B1(n1072), .B2(\mem[4][0] ), 
        .ZN(n1073) );
  INV_X1 U591 ( .A(n1071), .ZN(n778) );
  AOI22_X1 U592 ( .A1(data_in[1]), .A2(n839), .B1(n1072), .B2(\mem[4][1] ), 
        .ZN(n1071) );
  INV_X1 U593 ( .A(n1070), .ZN(n777) );
  AOI22_X1 U594 ( .A1(data_in[2]), .A2(n839), .B1(n1072), .B2(\mem[4][2] ), 
        .ZN(n1070) );
  INV_X1 U595 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U596 ( .A1(data_in[3]), .A2(n839), .B1(n1072), .B2(\mem[4][3] ), 
        .ZN(n1069) );
  INV_X1 U597 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U598 ( .A1(data_in[4]), .A2(n839), .B1(n1072), .B2(\mem[4][4] ), 
        .ZN(n1068) );
  INV_X1 U599 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U600 ( .A1(data_in[5]), .A2(n839), .B1(n1072), .B2(\mem[4][5] ), 
        .ZN(n1067) );
  INV_X1 U601 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U602 ( .A1(data_in[6]), .A2(n839), .B1(n1072), .B2(\mem[4][6] ), 
        .ZN(n1066) );
  INV_X1 U603 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U604 ( .A1(data_in[7]), .A2(n839), .B1(n1072), .B2(\mem[4][7] ), 
        .ZN(n1065) );
  INV_X1 U605 ( .A(N13), .ZN(n844) );
  INV_X1 U606 ( .A(N14), .ZN(n845) );
  MUX2_X1 U607 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n251), .Z(n3) );
  MUX2_X1 U608 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n251), .Z(n4) );
  MUX2_X1 U609 ( .A(n4), .B(n3), .S(n244), .Z(n5) );
  MUX2_X1 U610 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n251), .Z(n6) );
  MUX2_X1 U611 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n251), .Z(n7) );
  MUX2_X1 U612 ( .A(n7), .B(n6), .S(n246), .Z(n8) );
  MUX2_X1 U613 ( .A(n8), .B(n5), .S(n243), .Z(n9) );
  MUX2_X1 U614 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n251), .Z(n10) );
  MUX2_X1 U615 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n251), .Z(n11) );
  MUX2_X1 U616 ( .A(n11), .B(n10), .S(n245), .Z(n12) );
  MUX2_X1 U617 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n251), .Z(n13) );
  MUX2_X1 U618 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n250), .Z(n14) );
  MUX2_X1 U619 ( .A(n14), .B(n13), .S(n245), .Z(n15) );
  MUX2_X1 U620 ( .A(n15), .B(n12), .S(n243), .Z(n16) );
  MUX2_X1 U621 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U622 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n247), .Z(n18) );
  MUX2_X1 U623 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n247), .Z(n19) );
  MUX2_X1 U624 ( .A(n19), .B(n18), .S(n244), .Z(n20) );
  MUX2_X1 U625 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n247), .Z(n21) );
  MUX2_X1 U626 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n247), .Z(n22) );
  MUX2_X1 U627 ( .A(n22), .B(n21), .S(n244), .Z(n23) );
  MUX2_X1 U628 ( .A(n23), .B(n20), .S(n243), .Z(n24) );
  MUX2_X1 U629 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n247), .Z(n25) );
  MUX2_X1 U630 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n247), .Z(n26) );
  MUX2_X1 U631 ( .A(n26), .B(n25), .S(n244), .Z(n27) );
  MUX2_X1 U632 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n247), .Z(n28) );
  MUX2_X1 U633 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n247), .Z(n29) );
  MUX2_X1 U634 ( .A(n29), .B(n28), .S(n244), .Z(n30) );
  MUX2_X1 U635 ( .A(n30), .B(n27), .S(n243), .Z(n31) );
  MUX2_X1 U636 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U637 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U638 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n247), .Z(n33) );
  MUX2_X1 U639 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n247), .Z(n34) );
  MUX2_X1 U640 ( .A(n34), .B(n33), .S(n244), .Z(n35) );
  MUX2_X1 U641 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n247), .Z(n36) );
  MUX2_X1 U642 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n247), .Z(n37) );
  MUX2_X1 U643 ( .A(n37), .B(n36), .S(n244), .Z(n38) );
  MUX2_X1 U644 ( .A(n38), .B(n35), .S(n243), .Z(n39) );
  MUX2_X1 U645 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n248), .Z(n40) );
  MUX2_X1 U646 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n248), .Z(n41) );
  MUX2_X1 U647 ( .A(n41), .B(n40), .S(n244), .Z(n42) );
  MUX2_X1 U648 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n248), .Z(n43) );
  MUX2_X1 U649 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n248), .Z(n44) );
  MUX2_X1 U650 ( .A(n44), .B(n43), .S(n244), .Z(n45) );
  MUX2_X1 U651 ( .A(n45), .B(n42), .S(N12), .Z(n46) );
  MUX2_X1 U652 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U653 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n248), .Z(n48) );
  MUX2_X1 U654 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n248), .Z(n49) );
  MUX2_X1 U655 ( .A(n49), .B(n48), .S(n244), .Z(n50) );
  MUX2_X1 U656 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n248), .Z(n51) );
  MUX2_X1 U657 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n248), .Z(n52) );
  MUX2_X1 U658 ( .A(n52), .B(n51), .S(n244), .Z(n53) );
  MUX2_X1 U659 ( .A(n53), .B(n50), .S(N12), .Z(n54) );
  MUX2_X1 U660 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n248), .Z(n55) );
  MUX2_X1 U661 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n248), .Z(n56) );
  MUX2_X1 U662 ( .A(n56), .B(n55), .S(n244), .Z(n57) );
  MUX2_X1 U663 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n248), .Z(n58) );
  MUX2_X1 U664 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n248), .Z(n59) );
  MUX2_X1 U665 ( .A(n59), .B(n58), .S(n244), .Z(n60) );
  MUX2_X1 U666 ( .A(n60), .B(n57), .S(N12), .Z(n61) );
  MUX2_X1 U667 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U668 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U669 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n249), .Z(n63) );
  MUX2_X1 U670 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n249), .Z(n64) );
  MUX2_X1 U671 ( .A(n64), .B(n63), .S(n245), .Z(n65) );
  MUX2_X1 U672 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n249), .Z(n66) );
  MUX2_X1 U673 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n249), .Z(n67) );
  MUX2_X1 U674 ( .A(n67), .B(n66), .S(n245), .Z(n68) );
  MUX2_X1 U675 ( .A(n68), .B(n65), .S(n243), .Z(n69) );
  MUX2_X1 U676 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n249), .Z(n70) );
  MUX2_X1 U677 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n249), .Z(n71) );
  MUX2_X1 U678 ( .A(n71), .B(n70), .S(n245), .Z(n72) );
  MUX2_X1 U679 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n249), .Z(n73) );
  MUX2_X1 U680 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n249), .Z(n74) );
  MUX2_X1 U681 ( .A(n74), .B(n73), .S(n245), .Z(n75) );
  MUX2_X1 U682 ( .A(n75), .B(n72), .S(n243), .Z(n76) );
  MUX2_X1 U683 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U684 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n249), .Z(n78) );
  MUX2_X1 U685 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n249), .Z(n79) );
  MUX2_X1 U686 ( .A(n79), .B(n78), .S(n245), .Z(n80) );
  MUX2_X1 U687 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n249), .Z(n81) );
  MUX2_X1 U688 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n249), .Z(n82) );
  MUX2_X1 U689 ( .A(n82), .B(n81), .S(n245), .Z(n83) );
  MUX2_X1 U690 ( .A(n83), .B(n80), .S(n243), .Z(n84) );
  MUX2_X1 U691 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n248), .Z(n85) );
  MUX2_X1 U692 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n250), .Z(n86) );
  MUX2_X1 U693 ( .A(n86), .B(n85), .S(n245), .Z(n87) );
  MUX2_X1 U694 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n249), .Z(n88) );
  MUX2_X1 U695 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n249), .Z(n89) );
  MUX2_X1 U696 ( .A(n89), .B(n88), .S(n245), .Z(n90) );
  MUX2_X1 U697 ( .A(n90), .B(n87), .S(n243), .Z(n91) );
  MUX2_X1 U698 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U699 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U700 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n250), .Z(n93) );
  MUX2_X1 U701 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n252), .Z(n94) );
  MUX2_X1 U702 ( .A(n94), .B(n93), .S(n245), .Z(n95) );
  MUX2_X1 U703 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n247), .Z(n96) );
  MUX2_X1 U704 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n248), .Z(n97) );
  MUX2_X1 U705 ( .A(n97), .B(n96), .S(n245), .Z(n98) );
  MUX2_X1 U706 ( .A(n98), .B(n95), .S(n243), .Z(n99) );
  MUX2_X1 U707 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n100) );
  MUX2_X1 U708 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n247), .Z(n101) );
  MUX2_X1 U709 ( .A(n101), .B(n100), .S(n245), .Z(n102) );
  MUX2_X1 U710 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n249), .Z(n103) );
  MUX2_X1 U711 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n248), .Z(n104) );
  MUX2_X1 U712 ( .A(n104), .B(n103), .S(n245), .Z(n105) );
  MUX2_X1 U713 ( .A(n105), .B(n102), .S(n243), .Z(n106) );
  MUX2_X1 U714 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U715 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n251), .Z(n108) );
  MUX2_X1 U716 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(N10), .Z(n109) );
  MUX2_X1 U717 ( .A(n109), .B(n108), .S(n246), .Z(n110) );
  MUX2_X1 U718 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n252), .Z(n111) );
  MUX2_X1 U719 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n112) );
  MUX2_X1 U720 ( .A(n112), .B(n111), .S(n246), .Z(n113) );
  MUX2_X1 U721 ( .A(n113), .B(n110), .S(n243), .Z(n114) );
  MUX2_X1 U722 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n252), .Z(n115) );
  MUX2_X1 U723 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n116) );
  MUX2_X1 U724 ( .A(n116), .B(n115), .S(n246), .Z(n117) );
  MUX2_X1 U725 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n118) );
  MUX2_X1 U726 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n119) );
  MUX2_X1 U727 ( .A(n119), .B(n118), .S(n246), .Z(n120) );
  MUX2_X1 U728 ( .A(n120), .B(n117), .S(n243), .Z(n121) );
  MUX2_X1 U729 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U730 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U731 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n251), .Z(n123) );
  MUX2_X1 U732 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(N10), .Z(n124) );
  MUX2_X1 U733 ( .A(n124), .B(n123), .S(n246), .Z(n125) );
  MUX2_X1 U734 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n251), .Z(n126) );
  MUX2_X1 U735 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n127) );
  MUX2_X1 U736 ( .A(n127), .B(n126), .S(n246), .Z(n128) );
  MUX2_X1 U737 ( .A(n128), .B(n125), .S(n243), .Z(n129) );
  MUX2_X1 U738 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n250), .Z(n130) );
  MUX2_X1 U739 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n250), .Z(n131) );
  MUX2_X1 U740 ( .A(n131), .B(n130), .S(n246), .Z(n132) );
  MUX2_X1 U741 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n250), .Z(n133) );
  MUX2_X1 U742 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n250), .Z(n134) );
  MUX2_X1 U743 ( .A(n134), .B(n133), .S(n246), .Z(n135) );
  MUX2_X1 U744 ( .A(n135), .B(n132), .S(n243), .Z(n136) );
  MUX2_X1 U745 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U746 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n250), .Z(n138) );
  MUX2_X1 U747 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n250), .Z(n139) );
  MUX2_X1 U748 ( .A(n139), .B(n138), .S(n246), .Z(n140) );
  MUX2_X1 U749 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n250), .Z(n141) );
  MUX2_X1 U750 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n250), .Z(n142) );
  MUX2_X1 U751 ( .A(n142), .B(n141), .S(n246), .Z(n143) );
  MUX2_X1 U752 ( .A(n143), .B(n140), .S(n243), .Z(n144) );
  MUX2_X1 U753 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n250), .Z(n145) );
  MUX2_X1 U754 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n250), .Z(n146) );
  MUX2_X1 U755 ( .A(n146), .B(n145), .S(n246), .Z(n147) );
  MUX2_X1 U756 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n250), .Z(n148) );
  MUX2_X1 U757 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n250), .Z(n149) );
  MUX2_X1 U758 ( .A(n149), .B(n148), .S(n246), .Z(n150) );
  MUX2_X1 U759 ( .A(n150), .B(n147), .S(n243), .Z(n151) );
  MUX2_X1 U760 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U761 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U762 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n251), .Z(n153) );
  MUX2_X1 U763 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n251), .Z(n154) );
  MUX2_X1 U764 ( .A(n154), .B(n153), .S(N11), .Z(n155) );
  MUX2_X1 U765 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n251), .Z(n156) );
  MUX2_X1 U766 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n251), .Z(n157) );
  MUX2_X1 U767 ( .A(n157), .B(n156), .S(N11), .Z(n158) );
  MUX2_X1 U768 ( .A(n158), .B(n155), .S(n243), .Z(n159) );
  MUX2_X1 U769 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n251), .Z(n160) );
  MUX2_X1 U770 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n251), .Z(n161) );
  MUX2_X1 U771 ( .A(n161), .B(n160), .S(N11), .Z(n162) );
  MUX2_X1 U772 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n251), .Z(n163) );
  MUX2_X1 U773 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n251), .Z(n164) );
  MUX2_X1 U774 ( .A(n164), .B(n163), .S(n246), .Z(n165) );
  MUX2_X1 U775 ( .A(n165), .B(n162), .S(N12), .Z(n166) );
  MUX2_X1 U776 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U777 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n251), .Z(n168) );
  MUX2_X1 U778 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n251), .Z(n169) );
  MUX2_X1 U779 ( .A(n169), .B(n168), .S(N11), .Z(n170) );
  MUX2_X1 U780 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n251), .Z(n171) );
  MUX2_X1 U781 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n251), .Z(n172) );
  MUX2_X1 U782 ( .A(n172), .B(n171), .S(n244), .Z(n173) );
  MUX2_X1 U783 ( .A(n173), .B(n170), .S(n243), .Z(n174) );
  MUX2_X1 U784 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n248), .Z(n175) );
  MUX2_X1 U785 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n247), .Z(n176) );
  MUX2_X1 U786 ( .A(n176), .B(n175), .S(N11), .Z(n177) );
  MUX2_X1 U787 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n252), .Z(n178) );
  MUX2_X1 U788 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n247), .Z(n179) );
  MUX2_X1 U789 ( .A(n179), .B(n178), .S(n246), .Z(n180) );
  MUX2_X1 U790 ( .A(n180), .B(n177), .S(N12), .Z(n181) );
  MUX2_X1 U791 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U792 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U793 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n252), .Z(n183) );
  MUX2_X1 U794 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n249), .Z(n184) );
  MUX2_X1 U795 ( .A(n184), .B(n183), .S(N11), .Z(n185) );
  MUX2_X1 U796 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n252), .Z(n186) );
  MUX2_X1 U797 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n252), .Z(n187) );
  MUX2_X1 U798 ( .A(n187), .B(n186), .S(N11), .Z(n188) );
  MUX2_X1 U799 ( .A(n188), .B(n185), .S(n243), .Z(n189) );
  MUX2_X1 U800 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n247), .Z(n190) );
  MUX2_X1 U801 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n250), .Z(n191) );
  MUX2_X1 U802 ( .A(n191), .B(n190), .S(N11), .Z(n192) );
  MUX2_X1 U803 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n247), .Z(n193) );
  MUX2_X1 U804 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n252), .Z(n194) );
  MUX2_X1 U805 ( .A(n194), .B(n193), .S(n244), .Z(n195) );
  MUX2_X1 U806 ( .A(n195), .B(n192), .S(N12), .Z(n196) );
  MUX2_X1 U807 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U808 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n252), .Z(n198) );
  MUX2_X1 U809 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n248), .Z(n199) );
  MUX2_X1 U810 ( .A(n199), .B(n198), .S(n245), .Z(n200) );
  MUX2_X1 U811 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n252), .Z(n201) );
  MUX2_X1 U812 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n252), .Z(n202) );
  MUX2_X1 U813 ( .A(n202), .B(n201), .S(n245), .Z(n203) );
  MUX2_X1 U814 ( .A(n203), .B(n200), .S(n243), .Z(n204) );
  MUX2_X1 U815 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n252), .Z(n205) );
  MUX2_X1 U816 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n251), .Z(n206) );
  MUX2_X1 U817 ( .A(n206), .B(n205), .S(n245), .Z(n207) );
  MUX2_X1 U818 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n249), .Z(n208) );
  MUX2_X1 U819 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n252), .Z(n209) );
  MUX2_X1 U820 ( .A(n209), .B(n208), .S(N11), .Z(n210) );
  MUX2_X1 U821 ( .A(n210), .B(n207), .S(N12), .Z(n211) );
  MUX2_X1 U822 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U823 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U824 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n252), .Z(n213) );
  MUX2_X1 U825 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n252), .Z(n214) );
  MUX2_X1 U826 ( .A(n214), .B(n213), .S(n244), .Z(n215) );
  MUX2_X1 U827 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n252), .Z(n216) );
  MUX2_X1 U828 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n252), .Z(n217) );
  MUX2_X1 U829 ( .A(n217), .B(n216), .S(n244), .Z(n218) );
  MUX2_X1 U830 ( .A(n218), .B(n215), .S(n243), .Z(n219) );
  MUX2_X1 U831 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n252), .Z(n220) );
  MUX2_X1 U832 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(N10), .Z(n221) );
  MUX2_X1 U833 ( .A(n221), .B(n220), .S(N11), .Z(n222) );
  MUX2_X1 U834 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(N10), .Z(n223) );
  MUX2_X1 U835 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n252), .Z(n224) );
  MUX2_X1 U836 ( .A(n224), .B(n223), .S(N11), .Z(n225) );
  MUX2_X1 U837 ( .A(n225), .B(n222), .S(N12), .Z(n226) );
  MUX2_X1 U838 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U839 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n252), .Z(n228) );
  MUX2_X1 U840 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n229) );
  MUX2_X1 U841 ( .A(n229), .B(n228), .S(n246), .Z(n230) );
  MUX2_X1 U842 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(N10), .Z(n231) );
  MUX2_X1 U843 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n232) );
  MUX2_X1 U844 ( .A(n232), .B(n231), .S(N11), .Z(n233) );
  MUX2_X1 U845 ( .A(n233), .B(n230), .S(n243), .Z(n234) );
  MUX2_X1 U846 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n235) );
  MUX2_X1 U847 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n248), .Z(n236) );
  MUX2_X1 U848 ( .A(n236), .B(n235), .S(n246), .Z(n237) );
  MUX2_X1 U849 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n238) );
  MUX2_X1 U850 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n249), .Z(n239) );
  MUX2_X1 U851 ( .A(n239), .B(n238), .S(N11), .Z(n240) );
  MUX2_X1 U852 ( .A(n240), .B(n237), .S(N12), .Z(n241) );
  MUX2_X1 U853 ( .A(n241), .B(n234), .S(N13), .Z(n242) );
  MUX2_X1 U854 ( .A(n242), .B(n227), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_16 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n256), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n257), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n258), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n259), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n260), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n261), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n262), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n263), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n264), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n265), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n266), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n267), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n268), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n269), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n270), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n271), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n272), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n273), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n274), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n275), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n276), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n277), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n278), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n279), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n280), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n281), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n282), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n283), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n284), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n285), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n286), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n287), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n288), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n289), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n290), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n291), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n292), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n293), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n594), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n595), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n596), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n597), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n598), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n599), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n600), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n601), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n602), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n603), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n604), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n605), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n606), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n607), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n608), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n609), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n610), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n611), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n612), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n613), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n614), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n615), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n616), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n617), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n618), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n619), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n620), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n621), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n622), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n623), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n624), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n625), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n626), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n627), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n628), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n629), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n630), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n631), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n632), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n633), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n634), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n635), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n636), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n637), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n638), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n639), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n640), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n641), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n642), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n643), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n644), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n645), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n646), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n647), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n648), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n649), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n650), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n651), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n652), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n653), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n654), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n655), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n656), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n657), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n658), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n659), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n660), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n661), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n662), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n663), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n664), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n665), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n666), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n667), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n668), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n669), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n670), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n671), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n672), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n673), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n674), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n675), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n676), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n677), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n678), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n679), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n680), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n681), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n682), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n683), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n684), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n685), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n686), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n687), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n688), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n689), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n690), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n691), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n692), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n693), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n694), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n695), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n696), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n697), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n698), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n699), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n700), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n701), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n702), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n703), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n704), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n705), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n706), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n707), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n708), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n709), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n710), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n711), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n712), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n713), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n714), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n715), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n716), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n717), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n718), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n719), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n720), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n721), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n722), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n723), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n724), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n725), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n726), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n727), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n728), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n729), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n730), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n731), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n732), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n733), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n734), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n735), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n736), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n737), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n738), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n739), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n740), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n741), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n742), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n743), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n744), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n745), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n746), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n747), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n748), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n749), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n750), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n751), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n752), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n753), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n754), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n755), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n756), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n757), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n758), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n759), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n760), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n761), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n762), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n763), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n764), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n765), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n766), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n767), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n768), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n769), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n770), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n771), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n772), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n773), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n774), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n775), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n776), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n777), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n778), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n779), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n780), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n781), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n782), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n783), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n784), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n785), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n786), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n787), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n788), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n789), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n790), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n791), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n792), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n793), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n794), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n795), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n796), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n797), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n798), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n799), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n800), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n801), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n802), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n803), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n804), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n805), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n806), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n807), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n808), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n809), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n810), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n811), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(n252), .Z(n248) );
  BUF_X1 U5 ( .A(n252), .Z(n249) );
  BUF_X1 U6 ( .A(n252), .Z(n250) );
  BUF_X1 U7 ( .A(n252), .Z(n251) );
  BUF_X1 U8 ( .A(N10), .Z(n252) );
  INV_X1 U9 ( .A(n1113), .ZN(n843) );
  INV_X1 U10 ( .A(n1102), .ZN(n842) );
  INV_X1 U11 ( .A(n1092), .ZN(n841) );
  INV_X1 U12 ( .A(n1082), .ZN(n840) );
  INV_X1 U13 ( .A(n1072), .ZN(n839) );
  INV_X1 U14 ( .A(n1062), .ZN(n838) );
  INV_X1 U15 ( .A(n1053), .ZN(n837) );
  INV_X1 U16 ( .A(n1044), .ZN(n836) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1105) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n253), .ZN(n1094) );
  NAND2_X1 U19 ( .A1(n1104), .A2(n1136), .ZN(n1062) );
  NAND2_X1 U20 ( .A1(n1105), .A2(n1104), .ZN(n1113) );
  NAND2_X1 U21 ( .A1(n1094), .A2(n1104), .ZN(n1102) );
  NAND2_X1 U22 ( .A1(n1084), .A2(n1104), .ZN(n1092) );
  NAND2_X1 U23 ( .A1(n1074), .A2(n1104), .ZN(n1082) );
  NAND2_X1 U24 ( .A1(n1064), .A2(n1104), .ZN(n1072) );
  NAND2_X1 U25 ( .A1(n1104), .A2(n1125), .ZN(n1053) );
  NAND2_X1 U26 ( .A1(n1104), .A2(n1115), .ZN(n1044) );
  INV_X1 U27 ( .A(n1133), .ZN(n818) );
  INV_X1 U28 ( .A(n1123), .ZN(n817) );
  INV_X1 U29 ( .A(n889), .ZN(n816) );
  INV_X1 U30 ( .A(n880), .ZN(n815) );
  INV_X1 U31 ( .A(n871), .ZN(n814) );
  INV_X1 U32 ( .A(n862), .ZN(n813) );
  INV_X1 U33 ( .A(n853), .ZN(n812) );
  INV_X1 U34 ( .A(n989), .ZN(n830) );
  INV_X1 U35 ( .A(n980), .ZN(n829) );
  INV_X1 U36 ( .A(n971), .ZN(n828) );
  INV_X1 U37 ( .A(n916), .ZN(n822) );
  INV_X1 U38 ( .A(n907), .ZN(n821) );
  INV_X1 U39 ( .A(n898), .ZN(n820) );
  INV_X1 U40 ( .A(n1035), .ZN(n835) );
  INV_X1 U41 ( .A(n1025), .ZN(n834) );
  INV_X1 U42 ( .A(n1016), .ZN(n833) );
  INV_X1 U43 ( .A(n1007), .ZN(n832) );
  INV_X1 U44 ( .A(n998), .ZN(n831) );
  INV_X1 U45 ( .A(n962), .ZN(n827) );
  INV_X1 U46 ( .A(n952), .ZN(n826) );
  INV_X1 U47 ( .A(n943), .ZN(n825) );
  INV_X1 U48 ( .A(n934), .ZN(n824) );
  INV_X1 U49 ( .A(n925), .ZN(n823) );
  INV_X1 U50 ( .A(n1144), .ZN(n819) );
  BUF_X1 U51 ( .A(N11), .Z(n244) );
  BUF_X1 U52 ( .A(N11), .Z(n245) );
  BUF_X1 U53 ( .A(N11), .Z(n246) );
  INV_X1 U54 ( .A(N10), .ZN(n253) );
  BUF_X1 U55 ( .A(N12), .Z(n243) );
  NOR3_X1 U56 ( .A1(n255), .A2(N10), .A3(n254), .ZN(n1125) );
  NOR3_X1 U57 ( .A1(n255), .A2(n253), .A3(n254), .ZN(n1115) );
  NOR3_X1 U58 ( .A1(n253), .A2(N11), .A3(n255), .ZN(n1136) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n254), .ZN(n1084) );
  NOR3_X1 U60 ( .A1(n253), .A2(N12), .A3(n254), .ZN(n1074) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n255), .ZN(n1064) );
  NAND2_X1 U62 ( .A1(n1027), .A2(n1136), .ZN(n989) );
  NAND2_X1 U63 ( .A1(n954), .A2(n1136), .ZN(n916) );
  NAND2_X1 U64 ( .A1(n1027), .A2(n1064), .ZN(n998) );
  NAND2_X1 U65 ( .A1(n954), .A2(n1064), .ZN(n925) );
  NAND2_X1 U66 ( .A1(n1027), .A2(n1105), .ZN(n1035) );
  NAND2_X1 U67 ( .A1(n1027), .A2(n1094), .ZN(n1025) );
  NAND2_X1 U68 ( .A1(n954), .A2(n1105), .ZN(n962) );
  NAND2_X1 U69 ( .A1(n954), .A2(n1094), .ZN(n952) );
  NAND2_X1 U70 ( .A1(n1105), .A2(n1135), .ZN(n889) );
  NAND2_X1 U71 ( .A1(n1094), .A2(n1135), .ZN(n880) );
  NAND2_X1 U72 ( .A1(n1084), .A2(n1135), .ZN(n871) );
  NAND2_X1 U73 ( .A1(n1074), .A2(n1135), .ZN(n862) );
  NAND2_X1 U74 ( .A1(n1064), .A2(n1135), .ZN(n853) );
  NAND2_X1 U75 ( .A1(n1136), .A2(n1135), .ZN(n1144) );
  NAND2_X1 U76 ( .A1(n1125), .A2(n1135), .ZN(n1133) );
  NAND2_X1 U77 ( .A1(n1115), .A2(n1135), .ZN(n1123) );
  NAND2_X1 U78 ( .A1(n1027), .A2(n1084), .ZN(n1016) );
  NAND2_X1 U79 ( .A1(n1027), .A2(n1074), .ZN(n1007) );
  NAND2_X1 U80 ( .A1(n954), .A2(n1084), .ZN(n943) );
  NAND2_X1 U81 ( .A1(n954), .A2(n1074), .ZN(n934) );
  NAND2_X1 U82 ( .A1(n1027), .A2(n1125), .ZN(n980) );
  NAND2_X1 U83 ( .A1(n954), .A2(n1125), .ZN(n907) );
  NAND2_X1 U84 ( .A1(n1027), .A2(n1115), .ZN(n971) );
  NAND2_X1 U85 ( .A1(n954), .A2(n1115), .ZN(n898) );
  AND3_X1 U86 ( .A1(n844), .A2(n845), .A3(wr_en), .ZN(n1104) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1135) );
  AND3_X1 U88 ( .A1(N13), .A2(n845), .A3(wr_en), .ZN(n1027) );
  AND3_X1 U89 ( .A1(N14), .A2(n844), .A3(wr_en), .ZN(n954) );
  INV_X1 U90 ( .A(n1063), .ZN(n771) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n838), .B1(n1062), .B2(\mem[5][0] ), 
        .ZN(n1063) );
  INV_X1 U92 ( .A(n1061), .ZN(n770) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n838), .B1(n1062), .B2(\mem[5][1] ), 
        .ZN(n1061) );
  INV_X1 U94 ( .A(n1060), .ZN(n769) );
  AOI22_X1 U95 ( .A1(data_in[2]), .A2(n838), .B1(n1062), .B2(\mem[5][2] ), 
        .ZN(n1060) );
  INV_X1 U96 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U97 ( .A1(data_in[3]), .A2(n838), .B1(n1062), .B2(\mem[5][3] ), 
        .ZN(n1059) );
  INV_X1 U98 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U99 ( .A1(data_in[4]), .A2(n838), .B1(n1062), .B2(\mem[5][4] ), 
        .ZN(n1058) );
  INV_X1 U100 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U101 ( .A1(data_in[5]), .A2(n838), .B1(n1062), .B2(\mem[5][5] ), 
        .ZN(n1057) );
  INV_X1 U102 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U103 ( .A1(data_in[6]), .A2(n838), .B1(n1062), .B2(\mem[5][6] ), 
        .ZN(n1056) );
  INV_X1 U104 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U105 ( .A1(data_in[7]), .A2(n838), .B1(n1062), .B2(\mem[5][7] ), 
        .ZN(n1055) );
  INV_X1 U106 ( .A(n1026), .ZN(n739) );
  AOI22_X1 U107 ( .A1(data_in[0]), .A2(n834), .B1(n1025), .B2(\mem[9][0] ), 
        .ZN(n1026) );
  INV_X1 U108 ( .A(n1024), .ZN(n738) );
  AOI22_X1 U109 ( .A1(data_in[1]), .A2(n834), .B1(n1025), .B2(\mem[9][1] ), 
        .ZN(n1024) );
  INV_X1 U110 ( .A(n1023), .ZN(n737) );
  AOI22_X1 U111 ( .A1(data_in[2]), .A2(n834), .B1(n1025), .B2(\mem[9][2] ), 
        .ZN(n1023) );
  INV_X1 U112 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U113 ( .A1(data_in[3]), .A2(n834), .B1(n1025), .B2(\mem[9][3] ), 
        .ZN(n1022) );
  INV_X1 U114 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U115 ( .A1(data_in[4]), .A2(n834), .B1(n1025), .B2(\mem[9][4] ), 
        .ZN(n1021) );
  INV_X1 U116 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U117 ( .A1(data_in[5]), .A2(n834), .B1(n1025), .B2(\mem[9][5] ), 
        .ZN(n1020) );
  INV_X1 U118 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U119 ( .A1(data_in[6]), .A2(n834), .B1(n1025), .B2(\mem[9][6] ), 
        .ZN(n1019) );
  INV_X1 U120 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U121 ( .A1(data_in[7]), .A2(n834), .B1(n1025), .B2(\mem[9][7] ), 
        .ZN(n1018) );
  INV_X1 U122 ( .A(n990), .ZN(n707) );
  AOI22_X1 U123 ( .A1(data_in[0]), .A2(n830), .B1(n989), .B2(\mem[13][0] ), 
        .ZN(n990) );
  INV_X1 U124 ( .A(n988), .ZN(n706) );
  AOI22_X1 U125 ( .A1(data_in[1]), .A2(n830), .B1(n989), .B2(\mem[13][1] ), 
        .ZN(n988) );
  INV_X1 U126 ( .A(n987), .ZN(n705) );
  AOI22_X1 U127 ( .A1(data_in[2]), .A2(n830), .B1(n989), .B2(\mem[13][2] ), 
        .ZN(n987) );
  INV_X1 U128 ( .A(n986), .ZN(n704) );
  AOI22_X1 U129 ( .A1(data_in[3]), .A2(n830), .B1(n989), .B2(\mem[13][3] ), 
        .ZN(n986) );
  INV_X1 U130 ( .A(n985), .ZN(n703) );
  AOI22_X1 U131 ( .A1(data_in[4]), .A2(n830), .B1(n989), .B2(\mem[13][4] ), 
        .ZN(n985) );
  INV_X1 U132 ( .A(n984), .ZN(n702) );
  AOI22_X1 U133 ( .A1(data_in[5]), .A2(n830), .B1(n989), .B2(\mem[13][5] ), 
        .ZN(n984) );
  INV_X1 U134 ( .A(n983), .ZN(n701) );
  AOI22_X1 U135 ( .A1(data_in[6]), .A2(n830), .B1(n989), .B2(\mem[13][6] ), 
        .ZN(n983) );
  INV_X1 U136 ( .A(n982), .ZN(n700) );
  AOI22_X1 U137 ( .A1(data_in[7]), .A2(n830), .B1(n989), .B2(\mem[13][7] ), 
        .ZN(n982) );
  INV_X1 U138 ( .A(n914), .ZN(n641) );
  AOI22_X1 U139 ( .A1(data_in[2]), .A2(n822), .B1(n916), .B2(\mem[21][2] ), 
        .ZN(n914) );
  INV_X1 U140 ( .A(n913), .ZN(n640) );
  AOI22_X1 U141 ( .A1(data_in[3]), .A2(n822), .B1(n916), .B2(\mem[21][3] ), 
        .ZN(n913) );
  INV_X1 U142 ( .A(n912), .ZN(n639) );
  AOI22_X1 U143 ( .A1(data_in[4]), .A2(n822), .B1(n916), .B2(\mem[21][4] ), 
        .ZN(n912) );
  INV_X1 U144 ( .A(n911), .ZN(n638) );
  AOI22_X1 U145 ( .A1(data_in[5]), .A2(n822), .B1(n916), .B2(\mem[21][5] ), 
        .ZN(n911) );
  INV_X1 U146 ( .A(n910), .ZN(n637) );
  AOI22_X1 U147 ( .A1(data_in[6]), .A2(n822), .B1(n916), .B2(\mem[21][6] ), 
        .ZN(n910) );
  INV_X1 U148 ( .A(n909), .ZN(n636) );
  AOI22_X1 U149 ( .A1(data_in[7]), .A2(n822), .B1(n916), .B2(\mem[21][7] ), 
        .ZN(n909) );
  INV_X1 U150 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U151 ( .A1(data_in[6]), .A2(n832), .B1(n1007), .B2(\mem[11][6] ), 
        .ZN(n1001) );
  INV_X1 U152 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U153 ( .A1(data_in[7]), .A2(n832), .B1(n1007), .B2(\mem[11][7] ), 
        .ZN(n1000) );
  INV_X1 U154 ( .A(n953), .ZN(n675) );
  AOI22_X1 U155 ( .A1(data_in[0]), .A2(n826), .B1(n952), .B2(\mem[17][0] ), 
        .ZN(n953) );
  INV_X1 U156 ( .A(n951), .ZN(n674) );
  AOI22_X1 U157 ( .A1(data_in[1]), .A2(n826), .B1(n952), .B2(\mem[17][1] ), 
        .ZN(n951) );
  INV_X1 U158 ( .A(n950), .ZN(n673) );
  AOI22_X1 U159 ( .A1(data_in[2]), .A2(n826), .B1(n952), .B2(\mem[17][2] ), 
        .ZN(n950) );
  INV_X1 U160 ( .A(n949), .ZN(n672) );
  AOI22_X1 U161 ( .A1(data_in[3]), .A2(n826), .B1(n952), .B2(\mem[17][3] ), 
        .ZN(n949) );
  INV_X1 U162 ( .A(n948), .ZN(n671) );
  AOI22_X1 U163 ( .A1(data_in[4]), .A2(n826), .B1(n952), .B2(\mem[17][4] ), 
        .ZN(n948) );
  INV_X1 U164 ( .A(n947), .ZN(n670) );
  AOI22_X1 U165 ( .A1(data_in[5]), .A2(n826), .B1(n952), .B2(\mem[17][5] ), 
        .ZN(n947) );
  INV_X1 U166 ( .A(n946), .ZN(n669) );
  AOI22_X1 U167 ( .A1(data_in[6]), .A2(n826), .B1(n952), .B2(\mem[17][6] ), 
        .ZN(n946) );
  INV_X1 U168 ( .A(n945), .ZN(n668) );
  AOI22_X1 U169 ( .A1(data_in[7]), .A2(n826), .B1(n952), .B2(\mem[17][7] ), 
        .ZN(n945) );
  INV_X1 U170 ( .A(n917), .ZN(n643) );
  AOI22_X1 U171 ( .A1(data_in[0]), .A2(n822), .B1(n916), .B2(\mem[21][0] ), 
        .ZN(n917) );
  INV_X1 U172 ( .A(n915), .ZN(n642) );
  AOI22_X1 U173 ( .A1(data_in[1]), .A2(n822), .B1(n916), .B2(\mem[21][1] ), 
        .ZN(n915) );
  INV_X1 U174 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U175 ( .A1(data_in[0]), .A2(n837), .B1(n1053), .B2(\mem[6][0] ), 
        .ZN(n1054) );
  INV_X1 U176 ( .A(n1052), .ZN(n762) );
  AOI22_X1 U177 ( .A1(data_in[1]), .A2(n837), .B1(n1053), .B2(\mem[6][1] ), 
        .ZN(n1052) );
  INV_X1 U178 ( .A(n1051), .ZN(n761) );
  AOI22_X1 U179 ( .A1(data_in[2]), .A2(n837), .B1(n1053), .B2(\mem[6][2] ), 
        .ZN(n1051) );
  INV_X1 U180 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U181 ( .A1(data_in[3]), .A2(n837), .B1(n1053), .B2(\mem[6][3] ), 
        .ZN(n1050) );
  INV_X1 U182 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U183 ( .A1(data_in[4]), .A2(n837), .B1(n1053), .B2(\mem[6][4] ), 
        .ZN(n1049) );
  INV_X1 U184 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U185 ( .A1(data_in[5]), .A2(n837), .B1(n1053), .B2(\mem[6][5] ), 
        .ZN(n1048) );
  INV_X1 U186 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U187 ( .A1(data_in[6]), .A2(n837), .B1(n1053), .B2(\mem[6][6] ), 
        .ZN(n1047) );
  INV_X1 U188 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U189 ( .A1(data_in[7]), .A2(n837), .B1(n1053), .B2(\mem[6][7] ), 
        .ZN(n1046) );
  INV_X1 U190 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U191 ( .A1(data_in[0]), .A2(n836), .B1(n1044), .B2(\mem[7][0] ), 
        .ZN(n1045) );
  INV_X1 U192 ( .A(n1043), .ZN(n754) );
  AOI22_X1 U193 ( .A1(data_in[1]), .A2(n836), .B1(n1044), .B2(\mem[7][1] ), 
        .ZN(n1043) );
  INV_X1 U194 ( .A(n1042), .ZN(n753) );
  AOI22_X1 U195 ( .A1(data_in[2]), .A2(n836), .B1(n1044), .B2(\mem[7][2] ), 
        .ZN(n1042) );
  INV_X1 U196 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U197 ( .A1(data_in[3]), .A2(n836), .B1(n1044), .B2(\mem[7][3] ), 
        .ZN(n1041) );
  INV_X1 U198 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U199 ( .A1(data_in[4]), .A2(n836), .B1(n1044), .B2(\mem[7][4] ), 
        .ZN(n1040) );
  INV_X1 U200 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U201 ( .A1(data_in[5]), .A2(n836), .B1(n1044), .B2(\mem[7][5] ), 
        .ZN(n1039) );
  INV_X1 U202 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U203 ( .A1(data_in[6]), .A2(n836), .B1(n1044), .B2(\mem[7][6] ), 
        .ZN(n1038) );
  INV_X1 U204 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U205 ( .A1(data_in[7]), .A2(n836), .B1(n1044), .B2(\mem[7][7] ), 
        .ZN(n1037) );
  INV_X1 U206 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U207 ( .A1(data_in[0]), .A2(n833), .B1(n1016), .B2(\mem[10][0] ), 
        .ZN(n1017) );
  INV_X1 U208 ( .A(n1015), .ZN(n730) );
  AOI22_X1 U209 ( .A1(data_in[1]), .A2(n833), .B1(n1016), .B2(\mem[10][1] ), 
        .ZN(n1015) );
  INV_X1 U210 ( .A(n1014), .ZN(n729) );
  AOI22_X1 U211 ( .A1(data_in[2]), .A2(n833), .B1(n1016), .B2(\mem[10][2] ), 
        .ZN(n1014) );
  INV_X1 U212 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U213 ( .A1(data_in[3]), .A2(n833), .B1(n1016), .B2(\mem[10][3] ), 
        .ZN(n1013) );
  INV_X1 U214 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U215 ( .A1(data_in[4]), .A2(n833), .B1(n1016), .B2(\mem[10][4] ), 
        .ZN(n1012) );
  INV_X1 U216 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U217 ( .A1(data_in[5]), .A2(n833), .B1(n1016), .B2(\mem[10][5] ), 
        .ZN(n1011) );
  INV_X1 U218 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U219 ( .A1(data_in[6]), .A2(n833), .B1(n1016), .B2(\mem[10][6] ), 
        .ZN(n1010) );
  INV_X1 U220 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U221 ( .A1(data_in[7]), .A2(n833), .B1(n1016), .B2(\mem[10][7] ), 
        .ZN(n1009) );
  INV_X1 U222 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U223 ( .A1(data_in[0]), .A2(n832), .B1(n1007), .B2(\mem[11][0] ), 
        .ZN(n1008) );
  INV_X1 U224 ( .A(n1006), .ZN(n722) );
  AOI22_X1 U225 ( .A1(data_in[1]), .A2(n832), .B1(n1007), .B2(\mem[11][1] ), 
        .ZN(n1006) );
  INV_X1 U226 ( .A(n1005), .ZN(n721) );
  AOI22_X1 U227 ( .A1(data_in[2]), .A2(n832), .B1(n1007), .B2(\mem[11][2] ), 
        .ZN(n1005) );
  INV_X1 U228 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U229 ( .A1(data_in[3]), .A2(n832), .B1(n1007), .B2(\mem[11][3] ), 
        .ZN(n1004) );
  INV_X1 U230 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U231 ( .A1(data_in[4]), .A2(n832), .B1(n1007), .B2(\mem[11][4] ), 
        .ZN(n1003) );
  INV_X1 U232 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U233 ( .A1(data_in[5]), .A2(n832), .B1(n1007), .B2(\mem[11][5] ), 
        .ZN(n1002) );
  INV_X1 U234 ( .A(n981), .ZN(n699) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n829), .B1(n980), .B2(\mem[14][0] ), 
        .ZN(n981) );
  INV_X1 U236 ( .A(n979), .ZN(n698) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n829), .B1(n980), .B2(\mem[14][1] ), 
        .ZN(n979) );
  INV_X1 U238 ( .A(n978), .ZN(n697) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n829), .B1(n980), .B2(\mem[14][2] ), 
        .ZN(n978) );
  INV_X1 U240 ( .A(n977), .ZN(n696) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n829), .B1(n980), .B2(\mem[14][3] ), 
        .ZN(n977) );
  INV_X1 U242 ( .A(n976), .ZN(n695) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n829), .B1(n980), .B2(\mem[14][4] ), 
        .ZN(n976) );
  INV_X1 U244 ( .A(n975), .ZN(n694) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n829), .B1(n980), .B2(\mem[14][5] ), 
        .ZN(n975) );
  INV_X1 U246 ( .A(n974), .ZN(n693) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n829), .B1(n980), .B2(\mem[14][6] ), 
        .ZN(n974) );
  INV_X1 U248 ( .A(n973), .ZN(n692) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n829), .B1(n980), .B2(\mem[14][7] ), 
        .ZN(n973) );
  INV_X1 U250 ( .A(n972), .ZN(n691) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n828), .B1(n971), .B2(\mem[15][0] ), 
        .ZN(n972) );
  INV_X1 U252 ( .A(n970), .ZN(n690) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n828), .B1(n971), .B2(\mem[15][1] ), 
        .ZN(n970) );
  INV_X1 U254 ( .A(n969), .ZN(n689) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n828), .B1(n971), .B2(\mem[15][2] ), 
        .ZN(n969) );
  INV_X1 U256 ( .A(n968), .ZN(n688) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n828), .B1(n971), .B2(\mem[15][3] ), 
        .ZN(n968) );
  INV_X1 U258 ( .A(n967), .ZN(n687) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n828), .B1(n971), .B2(\mem[15][4] ), 
        .ZN(n967) );
  INV_X1 U260 ( .A(n966), .ZN(n686) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n828), .B1(n971), .B2(\mem[15][5] ), 
        .ZN(n966) );
  INV_X1 U262 ( .A(n965), .ZN(n685) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n828), .B1(n971), .B2(\mem[15][6] ), 
        .ZN(n965) );
  INV_X1 U264 ( .A(n964), .ZN(n684) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n828), .B1(n971), .B2(\mem[15][7] ), 
        .ZN(n964) );
  INV_X1 U266 ( .A(n944), .ZN(n667) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n825), .B1(n943), .B2(\mem[18][0] ), 
        .ZN(n944) );
  INV_X1 U268 ( .A(n942), .ZN(n666) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n825), .B1(n943), .B2(\mem[18][1] ), 
        .ZN(n942) );
  INV_X1 U270 ( .A(n941), .ZN(n665) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n825), .B1(n943), .B2(\mem[18][2] ), 
        .ZN(n941) );
  INV_X1 U272 ( .A(n940), .ZN(n664) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n825), .B1(n943), .B2(\mem[18][3] ), 
        .ZN(n940) );
  INV_X1 U274 ( .A(n939), .ZN(n663) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n825), .B1(n943), .B2(\mem[18][4] ), 
        .ZN(n939) );
  INV_X1 U276 ( .A(n938), .ZN(n662) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n825), .B1(n943), .B2(\mem[18][5] ), 
        .ZN(n938) );
  INV_X1 U278 ( .A(n937), .ZN(n661) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n825), .B1(n943), .B2(\mem[18][6] ), 
        .ZN(n937) );
  INV_X1 U280 ( .A(n936), .ZN(n660) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n825), .B1(n943), .B2(\mem[18][7] ), 
        .ZN(n936) );
  INV_X1 U282 ( .A(n935), .ZN(n659) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n824), .B1(n934), .B2(\mem[19][0] ), 
        .ZN(n935) );
  INV_X1 U284 ( .A(n933), .ZN(n658) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n824), .B1(n934), .B2(\mem[19][1] ), 
        .ZN(n933) );
  INV_X1 U286 ( .A(n932), .ZN(n657) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n824), .B1(n934), .B2(\mem[19][2] ), 
        .ZN(n932) );
  INV_X1 U288 ( .A(n931), .ZN(n656) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n824), .B1(n934), .B2(\mem[19][3] ), 
        .ZN(n931) );
  INV_X1 U290 ( .A(n930), .ZN(n655) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n824), .B1(n934), .B2(\mem[19][4] ), 
        .ZN(n930) );
  INV_X1 U292 ( .A(n929), .ZN(n654) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n824), .B1(n934), .B2(\mem[19][5] ), 
        .ZN(n929) );
  INV_X1 U294 ( .A(n928), .ZN(n653) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n824), .B1(n934), .B2(\mem[19][6] ), 
        .ZN(n928) );
  INV_X1 U296 ( .A(n927), .ZN(n652) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n824), .B1(n934), .B2(\mem[19][7] ), 
        .ZN(n927) );
  INV_X1 U298 ( .A(n908), .ZN(n635) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n821), .B1(n907), .B2(\mem[22][0] ), 
        .ZN(n908) );
  INV_X1 U300 ( .A(n906), .ZN(n634) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n821), .B1(n907), .B2(\mem[22][1] ), 
        .ZN(n906) );
  INV_X1 U302 ( .A(n905), .ZN(n633) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n821), .B1(n907), .B2(\mem[22][2] ), 
        .ZN(n905) );
  INV_X1 U304 ( .A(n904), .ZN(n632) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n821), .B1(n907), .B2(\mem[22][3] ), 
        .ZN(n904) );
  INV_X1 U306 ( .A(n903), .ZN(n631) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n821), .B1(n907), .B2(\mem[22][4] ), 
        .ZN(n903) );
  INV_X1 U308 ( .A(n902), .ZN(n630) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n821), .B1(n907), .B2(\mem[22][5] ), 
        .ZN(n902) );
  INV_X1 U310 ( .A(n901), .ZN(n629) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n821), .B1(n907), .B2(\mem[22][6] ), 
        .ZN(n901) );
  INV_X1 U312 ( .A(n900), .ZN(n628) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n821), .B1(n907), .B2(\mem[22][7] ), 
        .ZN(n900) );
  INV_X1 U314 ( .A(n899), .ZN(n627) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n820), .B1(n898), .B2(\mem[23][0] ), 
        .ZN(n899) );
  INV_X1 U316 ( .A(n897), .ZN(n626) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n820), .B1(n898), .B2(\mem[23][1] ), 
        .ZN(n897) );
  INV_X1 U318 ( .A(n896), .ZN(n625) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n820), .B1(n898), .B2(\mem[23][2] ), 
        .ZN(n896) );
  INV_X1 U320 ( .A(n895), .ZN(n624) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n820), .B1(n898), .B2(\mem[23][3] ), 
        .ZN(n895) );
  INV_X1 U322 ( .A(n894), .ZN(n623) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n820), .B1(n898), .B2(\mem[23][4] ), 
        .ZN(n894) );
  INV_X1 U324 ( .A(n893), .ZN(n622) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n820), .B1(n898), .B2(\mem[23][5] ), 
        .ZN(n893) );
  INV_X1 U326 ( .A(n892), .ZN(n621) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n820), .B1(n898), .B2(\mem[23][6] ), 
        .ZN(n892) );
  INV_X1 U328 ( .A(n891), .ZN(n620) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n820), .B1(n898), .B2(\mem[23][7] ), 
        .ZN(n891) );
  INV_X1 U330 ( .A(N12), .ZN(n255) );
  INV_X1 U331 ( .A(N11), .ZN(n254) );
  INV_X1 U332 ( .A(n999), .ZN(n715) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n831), .B1(n998), .B2(\mem[12][0] ), 
        .ZN(n999) );
  INV_X1 U334 ( .A(n997), .ZN(n714) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n831), .B1(n998), .B2(\mem[12][1] ), 
        .ZN(n997) );
  INV_X1 U336 ( .A(n996), .ZN(n713) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n831), .B1(n998), .B2(\mem[12][2] ), 
        .ZN(n996) );
  INV_X1 U338 ( .A(n995), .ZN(n712) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n831), .B1(n998), .B2(\mem[12][3] ), 
        .ZN(n995) );
  INV_X1 U340 ( .A(n994), .ZN(n711) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n831), .B1(n998), .B2(\mem[12][4] ), 
        .ZN(n994) );
  INV_X1 U342 ( .A(n993), .ZN(n710) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n831), .B1(n998), .B2(\mem[12][5] ), 
        .ZN(n993) );
  INV_X1 U344 ( .A(n992), .ZN(n709) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n831), .B1(n998), .B2(\mem[12][6] ), 
        .ZN(n992) );
  INV_X1 U346 ( .A(n991), .ZN(n708) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n831), .B1(n998), .B2(\mem[12][7] ), 
        .ZN(n991) );
  INV_X1 U348 ( .A(n926), .ZN(n651) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n823), .B1(n925), .B2(\mem[20][0] ), 
        .ZN(n926) );
  INV_X1 U350 ( .A(n924), .ZN(n650) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n823), .B1(n925), .B2(\mem[20][1] ), 
        .ZN(n924) );
  INV_X1 U352 ( .A(n923), .ZN(n649) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n823), .B1(n925), .B2(\mem[20][2] ), 
        .ZN(n923) );
  INV_X1 U354 ( .A(n922), .ZN(n648) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n823), .B1(n925), .B2(\mem[20][3] ), 
        .ZN(n922) );
  INV_X1 U356 ( .A(n921), .ZN(n647) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n823), .B1(n925), .B2(\mem[20][4] ), 
        .ZN(n921) );
  INV_X1 U358 ( .A(n920), .ZN(n646) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n823), .B1(n925), .B2(\mem[20][5] ), 
        .ZN(n920) );
  INV_X1 U360 ( .A(n919), .ZN(n645) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n823), .B1(n925), .B2(\mem[20][6] ), 
        .ZN(n919) );
  INV_X1 U362 ( .A(n918), .ZN(n644) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n823), .B1(n925), .B2(\mem[20][7] ), 
        .ZN(n918) );
  INV_X1 U364 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n835), .B1(n1035), .B2(\mem[8][0] ), 
        .ZN(n1036) );
  INV_X1 U366 ( .A(n1034), .ZN(n746) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n835), .B1(n1035), .B2(\mem[8][1] ), 
        .ZN(n1034) );
  INV_X1 U368 ( .A(n1033), .ZN(n745) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n835), .B1(n1035), .B2(\mem[8][2] ), 
        .ZN(n1033) );
  INV_X1 U370 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n835), .B1(n1035), .B2(\mem[8][3] ), 
        .ZN(n1032) );
  INV_X1 U372 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n835), .B1(n1035), .B2(\mem[8][4] ), 
        .ZN(n1031) );
  INV_X1 U374 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n835), .B1(n1035), .B2(\mem[8][5] ), 
        .ZN(n1030) );
  INV_X1 U376 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n835), .B1(n1035), .B2(\mem[8][6] ), 
        .ZN(n1029) );
  INV_X1 U378 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n835), .B1(n1035), .B2(\mem[8][7] ), 
        .ZN(n1028) );
  INV_X1 U380 ( .A(n963), .ZN(n683) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n827), .B1(n962), .B2(\mem[16][0] ), 
        .ZN(n963) );
  INV_X1 U382 ( .A(n961), .ZN(n682) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n827), .B1(n962), .B2(\mem[16][1] ), 
        .ZN(n961) );
  INV_X1 U384 ( .A(n960), .ZN(n681) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n827), .B1(n962), .B2(\mem[16][2] ), 
        .ZN(n960) );
  INV_X1 U386 ( .A(n959), .ZN(n680) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n827), .B1(n962), .B2(\mem[16][3] ), 
        .ZN(n959) );
  INV_X1 U388 ( .A(n958), .ZN(n679) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n827), .B1(n962), .B2(\mem[16][4] ), 
        .ZN(n958) );
  INV_X1 U390 ( .A(n957), .ZN(n678) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n827), .B1(n962), .B2(\mem[16][5] ), 
        .ZN(n957) );
  INV_X1 U392 ( .A(n956), .ZN(n677) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n827), .B1(n962), .B2(\mem[16][6] ), 
        .ZN(n956) );
  INV_X1 U394 ( .A(n955), .ZN(n676) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n827), .B1(n962), .B2(\mem[16][7] ), 
        .ZN(n955) );
  INV_X1 U396 ( .A(n890), .ZN(n619) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n816), .B1(n889), .B2(\mem[24][0] ), 
        .ZN(n890) );
  INV_X1 U398 ( .A(n888), .ZN(n618) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n816), .B1(n889), .B2(\mem[24][1] ), 
        .ZN(n888) );
  INV_X1 U400 ( .A(n887), .ZN(n617) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n816), .B1(n889), .B2(\mem[24][2] ), 
        .ZN(n887) );
  INV_X1 U402 ( .A(n886), .ZN(n616) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n816), .B1(n889), .B2(\mem[24][3] ), 
        .ZN(n886) );
  INV_X1 U404 ( .A(n885), .ZN(n615) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n816), .B1(n889), .B2(\mem[24][4] ), 
        .ZN(n885) );
  INV_X1 U406 ( .A(n884), .ZN(n614) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n816), .B1(n889), .B2(\mem[24][5] ), 
        .ZN(n884) );
  INV_X1 U408 ( .A(n883), .ZN(n613) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n816), .B1(n889), .B2(\mem[24][6] ), 
        .ZN(n883) );
  INV_X1 U410 ( .A(n882), .ZN(n612) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n816), .B1(n889), .B2(\mem[24][7] ), 
        .ZN(n882) );
  INV_X1 U412 ( .A(n881), .ZN(n611) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n815), .B1(n880), .B2(\mem[25][0] ), 
        .ZN(n881) );
  INV_X1 U414 ( .A(n879), .ZN(n610) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n815), .B1(n880), .B2(\mem[25][1] ), 
        .ZN(n879) );
  INV_X1 U416 ( .A(n878), .ZN(n609) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n815), .B1(n880), .B2(\mem[25][2] ), 
        .ZN(n878) );
  INV_X1 U418 ( .A(n877), .ZN(n608) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n815), .B1(n880), .B2(\mem[25][3] ), 
        .ZN(n877) );
  INV_X1 U420 ( .A(n876), .ZN(n607) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n815), .B1(n880), .B2(\mem[25][4] ), 
        .ZN(n876) );
  INV_X1 U422 ( .A(n875), .ZN(n606) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n815), .B1(n880), .B2(\mem[25][5] ), 
        .ZN(n875) );
  INV_X1 U424 ( .A(n874), .ZN(n605) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n815), .B1(n880), .B2(\mem[25][6] ), 
        .ZN(n874) );
  INV_X1 U426 ( .A(n873), .ZN(n604) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n815), .B1(n880), .B2(\mem[25][7] ), 
        .ZN(n873) );
  INV_X1 U428 ( .A(n872), .ZN(n603) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n814), .B1(n871), .B2(\mem[26][0] ), 
        .ZN(n872) );
  INV_X1 U430 ( .A(n870), .ZN(n602) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n814), .B1(n871), .B2(\mem[26][1] ), 
        .ZN(n870) );
  INV_X1 U432 ( .A(n869), .ZN(n601) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n814), .B1(n871), .B2(\mem[26][2] ), 
        .ZN(n869) );
  INV_X1 U434 ( .A(n868), .ZN(n600) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n814), .B1(n871), .B2(\mem[26][3] ), 
        .ZN(n868) );
  INV_X1 U436 ( .A(n867), .ZN(n599) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n814), .B1(n871), .B2(\mem[26][4] ), 
        .ZN(n867) );
  INV_X1 U438 ( .A(n866), .ZN(n598) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n814), .B1(n871), .B2(\mem[26][5] ), 
        .ZN(n866) );
  INV_X1 U440 ( .A(n865), .ZN(n597) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n814), .B1(n871), .B2(\mem[26][6] ), 
        .ZN(n865) );
  INV_X1 U442 ( .A(n864), .ZN(n596) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n814), .B1(n871), .B2(\mem[26][7] ), 
        .ZN(n864) );
  INV_X1 U444 ( .A(n863), .ZN(n595) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n813), .B1(n862), .B2(\mem[27][0] ), 
        .ZN(n863) );
  INV_X1 U446 ( .A(n861), .ZN(n594) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n813), .B1(n862), .B2(\mem[27][1] ), 
        .ZN(n861) );
  INV_X1 U448 ( .A(n860), .ZN(n293) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n813), .B1(n862), .B2(\mem[27][2] ), 
        .ZN(n860) );
  INV_X1 U450 ( .A(n859), .ZN(n292) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n813), .B1(n862), .B2(\mem[27][3] ), 
        .ZN(n859) );
  INV_X1 U452 ( .A(n858), .ZN(n291) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n813), .B1(n862), .B2(\mem[27][4] ), 
        .ZN(n858) );
  INV_X1 U454 ( .A(n857), .ZN(n290) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n813), .B1(n862), .B2(\mem[27][5] ), 
        .ZN(n857) );
  INV_X1 U456 ( .A(n856), .ZN(n289) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n813), .B1(n862), .B2(\mem[27][6] ), 
        .ZN(n856) );
  INV_X1 U458 ( .A(n855), .ZN(n288) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n813), .B1(n862), .B2(\mem[27][7] ), 
        .ZN(n855) );
  INV_X1 U460 ( .A(n854), .ZN(n287) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n812), .B1(n853), .B2(\mem[28][0] ), 
        .ZN(n854) );
  INV_X1 U462 ( .A(n852), .ZN(n286) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n812), .B1(n853), .B2(\mem[28][1] ), 
        .ZN(n852) );
  INV_X1 U464 ( .A(n851), .ZN(n285) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n812), .B1(n853), .B2(\mem[28][2] ), 
        .ZN(n851) );
  INV_X1 U466 ( .A(n850), .ZN(n284) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n812), .B1(n853), .B2(\mem[28][3] ), 
        .ZN(n850) );
  INV_X1 U468 ( .A(n849), .ZN(n283) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n812), .B1(n853), .B2(\mem[28][4] ), 
        .ZN(n849) );
  INV_X1 U470 ( .A(n848), .ZN(n282) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n812), .B1(n853), .B2(\mem[28][5] ), 
        .ZN(n848) );
  INV_X1 U472 ( .A(n847), .ZN(n281) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n812), .B1(n853), .B2(\mem[28][6] ), 
        .ZN(n847) );
  INV_X1 U474 ( .A(n846), .ZN(n280) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n812), .B1(n853), .B2(\mem[28][7] ), 
        .ZN(n846) );
  INV_X1 U476 ( .A(n1145), .ZN(n279) );
  AOI22_X1 U477 ( .A1(n819), .A2(data_in[0]), .B1(n1144), .B2(\mem[29][0] ), 
        .ZN(n1145) );
  INV_X1 U478 ( .A(n1143), .ZN(n278) );
  AOI22_X1 U479 ( .A1(n819), .A2(data_in[1]), .B1(n1144), .B2(\mem[29][1] ), 
        .ZN(n1143) );
  INV_X1 U480 ( .A(n1142), .ZN(n277) );
  AOI22_X1 U481 ( .A1(n819), .A2(data_in[2]), .B1(n1144), .B2(\mem[29][2] ), 
        .ZN(n1142) );
  INV_X1 U482 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U483 ( .A1(n819), .A2(data_in[3]), .B1(n1144), .B2(\mem[29][3] ), 
        .ZN(n1141) );
  INV_X1 U484 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U485 ( .A1(n819), .A2(data_in[4]), .B1(n1144), .B2(\mem[29][4] ), 
        .ZN(n1140) );
  INV_X1 U486 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U487 ( .A1(n819), .A2(data_in[5]), .B1(n1144), .B2(\mem[29][5] ), 
        .ZN(n1139) );
  INV_X1 U488 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U489 ( .A1(n819), .A2(data_in[6]), .B1(n1144), .B2(\mem[29][6] ), 
        .ZN(n1138) );
  INV_X1 U490 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U491 ( .A1(n819), .A2(data_in[7]), .B1(n1144), .B2(\mem[29][7] ), 
        .ZN(n1137) );
  INV_X1 U492 ( .A(n1134), .ZN(n271) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n818), .B1(n1133), .B2(\mem[30][0] ), 
        .ZN(n1134) );
  INV_X1 U494 ( .A(n1132), .ZN(n270) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n818), .B1(n1133), .B2(\mem[30][1] ), 
        .ZN(n1132) );
  INV_X1 U496 ( .A(n1131), .ZN(n269) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n818), .B1(n1133), .B2(\mem[30][2] ), 
        .ZN(n1131) );
  INV_X1 U498 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n818), .B1(n1133), .B2(\mem[30][3] ), 
        .ZN(n1130) );
  INV_X1 U500 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n818), .B1(n1133), .B2(\mem[30][4] ), 
        .ZN(n1129) );
  INV_X1 U502 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n818), .B1(n1133), .B2(\mem[30][5] ), 
        .ZN(n1128) );
  INV_X1 U504 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n818), .B1(n1133), .B2(\mem[30][6] ), 
        .ZN(n1127) );
  INV_X1 U506 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n818), .B1(n1133), .B2(\mem[30][7] ), 
        .ZN(n1126) );
  INV_X1 U508 ( .A(n1124), .ZN(n263) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n817), .B1(n1123), .B2(\mem[31][0] ), 
        .ZN(n1124) );
  INV_X1 U510 ( .A(n1122), .ZN(n262) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n817), .B1(n1123), .B2(\mem[31][1] ), 
        .ZN(n1122) );
  INV_X1 U512 ( .A(n1121), .ZN(n261) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n817), .B1(n1123), .B2(\mem[31][2] ), 
        .ZN(n1121) );
  INV_X1 U514 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n817), .B1(n1123), .B2(\mem[31][3] ), 
        .ZN(n1120) );
  INV_X1 U516 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n817), .B1(n1123), .B2(\mem[31][4] ), 
        .ZN(n1119) );
  INV_X1 U518 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n817), .B1(n1123), .B2(\mem[31][5] ), 
        .ZN(n1118) );
  INV_X1 U520 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n817), .B1(n1123), .B2(\mem[31][6] ), 
        .ZN(n1117) );
  INV_X1 U522 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n817), .B1(n1123), .B2(\mem[31][7] ), 
        .ZN(n1116) );
  INV_X1 U524 ( .A(n1114), .ZN(n811) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n843), .B1(n1113), .B2(\mem[0][0] ), 
        .ZN(n1114) );
  INV_X1 U526 ( .A(n1112), .ZN(n810) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n843), .B1(n1113), .B2(\mem[0][1] ), 
        .ZN(n1112) );
  INV_X1 U528 ( .A(n1111), .ZN(n809) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n843), .B1(n1113), .B2(\mem[0][2] ), 
        .ZN(n1111) );
  INV_X1 U530 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n843), .B1(n1113), .B2(\mem[0][3] ), 
        .ZN(n1110) );
  INV_X1 U532 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n843), .B1(n1113), .B2(\mem[0][4] ), 
        .ZN(n1109) );
  INV_X1 U534 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n843), .B1(n1113), .B2(\mem[0][5] ), 
        .ZN(n1108) );
  INV_X1 U536 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n843), .B1(n1113), .B2(\mem[0][6] ), 
        .ZN(n1107) );
  INV_X1 U538 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n843), .B1(n1113), .B2(\mem[0][7] ), 
        .ZN(n1106) );
  INV_X1 U540 ( .A(n1103), .ZN(n803) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[1][0] ), 
        .ZN(n1103) );
  INV_X1 U542 ( .A(n1101), .ZN(n802) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[1][1] ), 
        .ZN(n1101) );
  INV_X1 U544 ( .A(n1100), .ZN(n801) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[1][2] ), 
        .ZN(n1100) );
  INV_X1 U546 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[1][3] ), 
        .ZN(n1099) );
  INV_X1 U548 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[1][4] ), 
        .ZN(n1098) );
  INV_X1 U550 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[1][5] ), 
        .ZN(n1097) );
  INV_X1 U552 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[1][6] ), 
        .ZN(n1096) );
  INV_X1 U554 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[1][7] ), 
        .ZN(n1095) );
  INV_X1 U556 ( .A(n1093), .ZN(n795) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n841), .B1(n1092), .B2(\mem[2][0] ), 
        .ZN(n1093) );
  INV_X1 U558 ( .A(n1091), .ZN(n794) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n841), .B1(n1092), .B2(\mem[2][1] ), 
        .ZN(n1091) );
  INV_X1 U560 ( .A(n1090), .ZN(n793) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n841), .B1(n1092), .B2(\mem[2][2] ), 
        .ZN(n1090) );
  INV_X1 U562 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n841), .B1(n1092), .B2(\mem[2][3] ), 
        .ZN(n1089) );
  INV_X1 U564 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n841), .B1(n1092), .B2(\mem[2][4] ), 
        .ZN(n1088) );
  INV_X1 U566 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n841), .B1(n1092), .B2(\mem[2][5] ), 
        .ZN(n1087) );
  INV_X1 U568 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n841), .B1(n1092), .B2(\mem[2][6] ), 
        .ZN(n1086) );
  INV_X1 U570 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n841), .B1(n1092), .B2(\mem[2][7] ), 
        .ZN(n1085) );
  INV_X1 U572 ( .A(n1083), .ZN(n787) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n840), .B1(n1082), .B2(\mem[3][0] ), 
        .ZN(n1083) );
  INV_X1 U574 ( .A(n1081), .ZN(n786) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n840), .B1(n1082), .B2(\mem[3][1] ), 
        .ZN(n1081) );
  INV_X1 U576 ( .A(n1080), .ZN(n785) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n840), .B1(n1082), .B2(\mem[3][2] ), 
        .ZN(n1080) );
  INV_X1 U578 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n840), .B1(n1082), .B2(\mem[3][3] ), 
        .ZN(n1079) );
  INV_X1 U580 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n840), .B1(n1082), .B2(\mem[3][4] ), 
        .ZN(n1078) );
  INV_X1 U582 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n840), .B1(n1082), .B2(\mem[3][5] ), 
        .ZN(n1077) );
  INV_X1 U584 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n840), .B1(n1082), .B2(\mem[3][6] ), 
        .ZN(n1076) );
  INV_X1 U586 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n840), .B1(n1082), .B2(\mem[3][7] ), 
        .ZN(n1075) );
  INV_X1 U588 ( .A(n1073), .ZN(n779) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n839), .B1(n1072), .B2(\mem[4][0] ), 
        .ZN(n1073) );
  INV_X1 U590 ( .A(n1071), .ZN(n778) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n839), .B1(n1072), .B2(\mem[4][1] ), 
        .ZN(n1071) );
  INV_X1 U592 ( .A(n1070), .ZN(n777) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n839), .B1(n1072), .B2(\mem[4][2] ), 
        .ZN(n1070) );
  INV_X1 U594 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n839), .B1(n1072), .B2(\mem[4][3] ), 
        .ZN(n1069) );
  INV_X1 U596 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n839), .B1(n1072), .B2(\mem[4][4] ), 
        .ZN(n1068) );
  INV_X1 U598 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n839), .B1(n1072), .B2(\mem[4][5] ), 
        .ZN(n1067) );
  INV_X1 U600 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n839), .B1(n1072), .B2(\mem[4][6] ), 
        .ZN(n1066) );
  INV_X1 U602 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n839), .B1(n1072), .B2(\mem[4][7] ), 
        .ZN(n1065) );
  INV_X1 U604 ( .A(N13), .ZN(n844) );
  INV_X1 U605 ( .A(N14), .ZN(n845) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n247), .Z(n3) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n247), .Z(n4) );
  MUX2_X1 U608 ( .A(n4), .B(n3), .S(n245), .Z(n5) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n247), .Z(n6) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n247), .Z(n7) );
  MUX2_X1 U611 ( .A(n7), .B(n6), .S(n245), .Z(n8) );
  MUX2_X1 U612 ( .A(n8), .B(n5), .S(n243), .Z(n9) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n247), .Z(n10) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n247), .Z(n11) );
  MUX2_X1 U615 ( .A(n11), .B(n10), .S(N11), .Z(n12) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n247), .Z(n13) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n247), .Z(n14) );
  MUX2_X1 U618 ( .A(n14), .B(n13), .S(N11), .Z(n15) );
  MUX2_X1 U619 ( .A(n15), .B(n12), .S(n243), .Z(n16) );
  MUX2_X1 U620 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n248), .Z(n18) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n248), .Z(n19) );
  MUX2_X1 U623 ( .A(n19), .B(n18), .S(n246), .Z(n20) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n248), .Z(n21) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n248), .Z(n22) );
  MUX2_X1 U626 ( .A(n22), .B(n21), .S(n244), .Z(n23) );
  MUX2_X1 U627 ( .A(n23), .B(n20), .S(n243), .Z(n24) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n248), .Z(n25) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n248), .Z(n26) );
  MUX2_X1 U630 ( .A(n26), .B(n25), .S(N11), .Z(n27) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n248), .Z(n28) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n248), .Z(n29) );
  MUX2_X1 U633 ( .A(n29), .B(n28), .S(n246), .Z(n30) );
  MUX2_X1 U634 ( .A(n30), .B(n27), .S(n243), .Z(n31) );
  MUX2_X1 U635 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U636 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n248), .Z(n33) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n248), .Z(n34) );
  MUX2_X1 U639 ( .A(n34), .B(n33), .S(n244), .Z(n35) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n248), .Z(n36) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n248), .Z(n37) );
  MUX2_X1 U642 ( .A(n37), .B(n36), .S(n244), .Z(n38) );
  MUX2_X1 U643 ( .A(n38), .B(n35), .S(n243), .Z(n39) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n249), .Z(n40) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n249), .Z(n41) );
  MUX2_X1 U646 ( .A(n41), .B(n40), .S(n246), .Z(n42) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n249), .Z(n43) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n249), .Z(n44) );
  MUX2_X1 U649 ( .A(n44), .B(n43), .S(n246), .Z(n45) );
  MUX2_X1 U650 ( .A(n45), .B(n42), .S(N12), .Z(n46) );
  MUX2_X1 U651 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n249), .Z(n48) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n249), .Z(n49) );
  MUX2_X1 U654 ( .A(n49), .B(n48), .S(N11), .Z(n50) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n249), .Z(n51) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n249), .Z(n52) );
  MUX2_X1 U657 ( .A(n52), .B(n51), .S(n245), .Z(n53) );
  MUX2_X1 U658 ( .A(n53), .B(n50), .S(N12), .Z(n54) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n249), .Z(n55) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n249), .Z(n56) );
  MUX2_X1 U661 ( .A(n56), .B(n55), .S(N11), .Z(n57) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n249), .Z(n58) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n249), .Z(n59) );
  MUX2_X1 U664 ( .A(n59), .B(n58), .S(N11), .Z(n60) );
  MUX2_X1 U665 ( .A(n60), .B(n57), .S(N12), .Z(n61) );
  MUX2_X1 U666 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U667 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n250), .Z(n63) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n250), .Z(n64) );
  MUX2_X1 U670 ( .A(n64), .B(n63), .S(n244), .Z(n65) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n250), .Z(n66) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n250), .Z(n67) );
  MUX2_X1 U673 ( .A(n67), .B(n66), .S(n244), .Z(n68) );
  MUX2_X1 U674 ( .A(n68), .B(n65), .S(n243), .Z(n69) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n250), .Z(n70) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n250), .Z(n71) );
  MUX2_X1 U677 ( .A(n71), .B(n70), .S(n244), .Z(n72) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n250), .Z(n73) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n250), .Z(n74) );
  MUX2_X1 U680 ( .A(n74), .B(n73), .S(n244), .Z(n75) );
  MUX2_X1 U681 ( .A(n75), .B(n72), .S(n243), .Z(n76) );
  MUX2_X1 U682 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n250), .Z(n78) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n250), .Z(n79) );
  MUX2_X1 U685 ( .A(n79), .B(n78), .S(n244), .Z(n80) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n250), .Z(n81) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n250), .Z(n82) );
  MUX2_X1 U688 ( .A(n82), .B(n81), .S(n244), .Z(n83) );
  MUX2_X1 U689 ( .A(n83), .B(n80), .S(n243), .Z(n84) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n251), .Z(n85) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n251), .Z(n86) );
  MUX2_X1 U692 ( .A(n86), .B(n85), .S(n244), .Z(n87) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n251), .Z(n88) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n251), .Z(n89) );
  MUX2_X1 U695 ( .A(n89), .B(n88), .S(n244), .Z(n90) );
  MUX2_X1 U696 ( .A(n90), .B(n87), .S(n243), .Z(n91) );
  MUX2_X1 U697 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U698 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n251), .Z(n93) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n251), .Z(n94) );
  MUX2_X1 U701 ( .A(n94), .B(n93), .S(n244), .Z(n95) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n251), .Z(n96) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n251), .Z(n97) );
  MUX2_X1 U704 ( .A(n97), .B(n96), .S(n244), .Z(n98) );
  MUX2_X1 U705 ( .A(n98), .B(n95), .S(n243), .Z(n99) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n251), .Z(n100) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n251), .Z(n101) );
  MUX2_X1 U708 ( .A(n101), .B(n100), .S(n244), .Z(n102) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n251), .Z(n103) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n251), .Z(n104) );
  MUX2_X1 U711 ( .A(n104), .B(n103), .S(n244), .Z(n105) );
  MUX2_X1 U712 ( .A(n105), .B(n102), .S(n243), .Z(n106) );
  MUX2_X1 U713 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n252), .Z(n108) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n247), .Z(n109) );
  MUX2_X1 U716 ( .A(n109), .B(n108), .S(n245), .Z(n110) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n252), .Z(n111) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n252), .Z(n112) );
  MUX2_X1 U719 ( .A(n112), .B(n111), .S(n245), .Z(n113) );
  MUX2_X1 U720 ( .A(n113), .B(n110), .S(n243), .Z(n114) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n249), .Z(n115) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n251), .Z(n116) );
  MUX2_X1 U723 ( .A(n116), .B(n115), .S(n245), .Z(n117) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n249), .Z(n118) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n252), .Z(n119) );
  MUX2_X1 U726 ( .A(n119), .B(n118), .S(n245), .Z(n120) );
  MUX2_X1 U727 ( .A(n120), .B(n117), .S(n243), .Z(n121) );
  MUX2_X1 U728 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U729 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(N10), .Z(n123) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n251), .Z(n124) );
  MUX2_X1 U732 ( .A(n124), .B(n123), .S(n245), .Z(n125) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n252), .Z(n126) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n252), .Z(n127) );
  MUX2_X1 U735 ( .A(n127), .B(n126), .S(n245), .Z(n128) );
  MUX2_X1 U736 ( .A(n128), .B(n125), .S(n243), .Z(n129) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n252), .Z(n130) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(N10), .Z(n131) );
  MUX2_X1 U739 ( .A(n131), .B(n130), .S(n245), .Z(n132) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(N10), .Z(n133) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n252), .Z(n134) );
  MUX2_X1 U742 ( .A(n134), .B(n133), .S(n245), .Z(n135) );
  MUX2_X1 U743 ( .A(n135), .B(n132), .S(n243), .Z(n136) );
  MUX2_X1 U744 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n248), .Z(n138) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(N10), .Z(n139) );
  MUX2_X1 U747 ( .A(n139), .B(n138), .S(n245), .Z(n140) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(N10), .Z(n141) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(N10), .Z(n142) );
  MUX2_X1 U750 ( .A(n142), .B(n141), .S(n245), .Z(n143) );
  MUX2_X1 U751 ( .A(n143), .B(n140), .S(n243), .Z(n144) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(N10), .Z(n145) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n248), .Z(n146) );
  MUX2_X1 U754 ( .A(n146), .B(n145), .S(n245), .Z(n147) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(N10), .Z(n148) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n247), .Z(n149) );
  MUX2_X1 U757 ( .A(n149), .B(n148), .S(n245), .Z(n150) );
  MUX2_X1 U758 ( .A(n150), .B(n147), .S(n243), .Z(n151) );
  MUX2_X1 U759 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U760 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n247), .Z(n153) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n252), .Z(n154) );
  MUX2_X1 U763 ( .A(n154), .B(n153), .S(n246), .Z(n155) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n247), .Z(n156) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(N10), .Z(n157) );
  MUX2_X1 U766 ( .A(n157), .B(n156), .S(n246), .Z(n158) );
  MUX2_X1 U767 ( .A(n158), .B(n155), .S(n243), .Z(n159) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(N10), .Z(n160) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(N10), .Z(n161) );
  MUX2_X1 U770 ( .A(n161), .B(n160), .S(n246), .Z(n162) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(N10), .Z(n163) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(N10), .Z(n164) );
  MUX2_X1 U773 ( .A(n164), .B(n163), .S(n246), .Z(n165) );
  MUX2_X1 U774 ( .A(n165), .B(n162), .S(N12), .Z(n166) );
  MUX2_X1 U775 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n247), .Z(n168) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(N10), .Z(n169) );
  MUX2_X1 U778 ( .A(n169), .B(n168), .S(n246), .Z(n170) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n250), .Z(n171) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(N10), .Z(n172) );
  MUX2_X1 U781 ( .A(n172), .B(n171), .S(n246), .Z(n173) );
  MUX2_X1 U782 ( .A(n173), .B(n170), .S(n243), .Z(n174) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n249), .Z(n175) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n250), .Z(n176) );
  MUX2_X1 U785 ( .A(n176), .B(n175), .S(n246), .Z(n177) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n249), .Z(n178) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n252), .Z(n179) );
  MUX2_X1 U788 ( .A(n179), .B(n178), .S(n246), .Z(n180) );
  MUX2_X1 U789 ( .A(n180), .B(n177), .S(N12), .Z(n181) );
  MUX2_X1 U790 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U791 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n247), .Z(n183) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n248), .Z(n184) );
  MUX2_X1 U794 ( .A(n184), .B(n183), .S(n246), .Z(n185) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n249), .Z(n186) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n251), .Z(n187) );
  MUX2_X1 U797 ( .A(n187), .B(n186), .S(n246), .Z(n188) );
  MUX2_X1 U798 ( .A(n188), .B(n185), .S(n243), .Z(n189) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n251), .Z(n190) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n248), .Z(n191) );
  MUX2_X1 U801 ( .A(n191), .B(n190), .S(n246), .Z(n192) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n250), .Z(n193) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n252), .Z(n194) );
  MUX2_X1 U804 ( .A(n194), .B(n193), .S(n246), .Z(n195) );
  MUX2_X1 U805 ( .A(n195), .B(n192), .S(N12), .Z(n196) );
  MUX2_X1 U806 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n247), .Z(n198) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n252), .Z(n199) );
  MUX2_X1 U809 ( .A(n199), .B(n198), .S(N11), .Z(n200) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n252), .Z(n201) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n250), .Z(n202) );
  MUX2_X1 U812 ( .A(n202), .B(n201), .S(n246), .Z(n203) );
  MUX2_X1 U813 ( .A(n203), .B(n200), .S(n243), .Z(n204) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n248), .Z(n205) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n252), .Z(n206) );
  MUX2_X1 U816 ( .A(n206), .B(n205), .S(N11), .Z(n207) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n252), .Z(n208) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n249), .Z(n209) );
  MUX2_X1 U819 ( .A(n209), .B(n208), .S(n244), .Z(n210) );
  MUX2_X1 U820 ( .A(n210), .B(n207), .S(N12), .Z(n211) );
  MUX2_X1 U821 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U822 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n252), .Z(n213) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n247), .Z(n214) );
  MUX2_X1 U825 ( .A(n214), .B(n213), .S(N11), .Z(n215) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n252), .Z(n216) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n251), .Z(n217) );
  MUX2_X1 U828 ( .A(n217), .B(n216), .S(N11), .Z(n218) );
  MUX2_X1 U829 ( .A(n218), .B(n215), .S(n243), .Z(n219) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n250), .Z(n220) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n252), .Z(n221) );
  MUX2_X1 U832 ( .A(n221), .B(n220), .S(N11), .Z(n222) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n250), .Z(n223) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n252), .Z(n224) );
  MUX2_X1 U835 ( .A(n224), .B(n223), .S(n245), .Z(n225) );
  MUX2_X1 U836 ( .A(n225), .B(n222), .S(N12), .Z(n226) );
  MUX2_X1 U837 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n251), .Z(n228) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n251), .Z(n229) );
  MUX2_X1 U840 ( .A(n229), .B(n228), .S(N11), .Z(n230) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n249), .Z(n231) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n252), .Z(n232) );
  MUX2_X1 U843 ( .A(n232), .B(n231), .S(n244), .Z(n233) );
  MUX2_X1 U844 ( .A(n233), .B(n230), .S(n243), .Z(n234) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n248), .Z(n235) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n247), .Z(n236) );
  MUX2_X1 U847 ( .A(n236), .B(n235), .S(N11), .Z(n237) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n248), .Z(n238) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n250), .Z(n239) );
  MUX2_X1 U850 ( .A(n239), .B(n238), .S(n245), .Z(n240) );
  MUX2_X1 U851 ( .A(n240), .B(n237), .S(N12), .Z(n241) );
  MUX2_X1 U852 ( .A(n241), .B(n234), .S(N13), .Z(n242) );
  MUX2_X1 U853 ( .A(n242), .B(n227), .S(N14), .Z(N15) );
  CLKBUF_X1 U854 ( .A(n252), .Z(n247) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_15 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n255), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n256), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n257), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n258), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n259), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n260), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n261), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n262), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n263), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n264), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n265), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n266), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n267), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n268), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n269), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n270), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n271), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n272), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n273), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n274), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n275), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n276), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n277), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n278), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n279), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n280), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n281), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n282), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n283), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n284), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n285), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n286), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n287), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n288), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n289), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n290), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n291), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n292), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n293), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n594), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n595), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n596), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n597), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n598), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n599), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n600), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n601), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n602), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n603), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n604), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n605), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n606), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n607), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n608), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n609), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n610), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n611), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n612), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n613), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n614), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n615), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n616), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n617), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n618), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n619), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n620), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n621), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n622), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n623), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n624), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n625), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n626), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n627), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n628), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n629), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n630), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n631), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n632), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n633), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n634), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n635), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n636), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n637), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n638), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n639), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n640), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n641), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n642), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n643), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n644), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n645), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n646), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n647), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n648), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n649), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n650), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n651), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n652), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n653), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n654), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n655), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n656), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n657), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n658), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n659), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n660), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n661), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n662), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n663), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n664), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n665), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n666), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n667), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n668), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n669), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n670), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n671), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n672), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n673), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n674), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n675), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n676), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n677), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n678), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n679), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n680), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n681), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n682), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n683), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n684), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n685), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n686), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n687), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n688), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n689), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n690), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n691), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n692), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n693), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n694), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n695), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n696), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n697), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n698), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n699), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n700), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n701), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n702), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n703), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n704), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n705), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n706), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n707), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n708), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n709), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n710), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n711), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n712), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n713), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n714), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n715), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n716), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n717), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n718), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n719), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n720), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n721), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n722), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n723), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n724), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n725), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n726), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n727), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n728), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n729), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n730), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n731), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n732), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n733), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n734), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n735), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n736), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n737), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n738), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n739), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n740), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n741), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n742), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n743), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n744), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n745), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n746), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n747), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n748), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n749), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n750), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n751), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n752), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n753), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n754), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n755), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n756), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n757), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n758), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n759), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n760), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n761), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n762), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n763), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n764), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n765), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n766), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n767), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n768), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n769), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n770), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n771), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n772), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n773), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n774), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n775), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n776), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n777), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n778), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n779), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n780), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n781), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n782), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n783), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n784), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n785), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n786), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n787), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n788), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n789), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n790), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n791), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n792), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n793), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n794), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n795), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n796), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n797), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n798), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n799), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n800), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n801), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n802), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n803), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n804), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n805), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n806), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n807), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n808), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n809), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n810), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  BUF_X1 U3 ( .A(n251), .Z(n248) );
  BUF_X1 U4 ( .A(n251), .Z(n247) );
  BUF_X1 U5 ( .A(n251), .Z(n249) );
  BUF_X1 U6 ( .A(n251), .Z(n250) );
  BUF_X1 U7 ( .A(N10), .Z(n251) );
  INV_X1 U8 ( .A(n1112), .ZN(n842) );
  INV_X1 U9 ( .A(n1101), .ZN(n841) );
  INV_X1 U10 ( .A(n1091), .ZN(n840) );
  INV_X1 U11 ( .A(n1081), .ZN(n839) );
  INV_X1 U12 ( .A(n1071), .ZN(n838) );
  INV_X1 U13 ( .A(n1061), .ZN(n837) );
  INV_X1 U14 ( .A(n1052), .ZN(n836) );
  INV_X1 U15 ( .A(n1043), .ZN(n835) );
  NOR3_X1 U16 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1104) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(n252), .ZN(n1093) );
  NAND2_X1 U18 ( .A1(n1103), .A2(n1135), .ZN(n1061) );
  NAND2_X1 U19 ( .A1(n1104), .A2(n1103), .ZN(n1112) );
  NAND2_X1 U20 ( .A1(n1093), .A2(n1103), .ZN(n1101) );
  NAND2_X1 U21 ( .A1(n1083), .A2(n1103), .ZN(n1091) );
  NAND2_X1 U22 ( .A1(n1073), .A2(n1103), .ZN(n1081) );
  NAND2_X1 U23 ( .A1(n1063), .A2(n1103), .ZN(n1071) );
  NAND2_X1 U24 ( .A1(n1103), .A2(n1124), .ZN(n1052) );
  NAND2_X1 U25 ( .A1(n1103), .A2(n1114), .ZN(n1043) );
  INV_X1 U26 ( .A(n1132), .ZN(n817) );
  INV_X1 U27 ( .A(n1122), .ZN(n816) );
  INV_X1 U28 ( .A(n888), .ZN(n815) );
  INV_X1 U29 ( .A(n879), .ZN(n814) );
  INV_X1 U30 ( .A(n870), .ZN(n813) );
  INV_X1 U31 ( .A(n861), .ZN(n812) );
  INV_X1 U32 ( .A(n852), .ZN(n811) );
  INV_X1 U33 ( .A(n988), .ZN(n829) );
  INV_X1 U34 ( .A(n979), .ZN(n828) );
  INV_X1 U35 ( .A(n970), .ZN(n827) );
  INV_X1 U36 ( .A(n915), .ZN(n821) );
  INV_X1 U37 ( .A(n906), .ZN(n820) );
  INV_X1 U38 ( .A(n897), .ZN(n819) );
  INV_X1 U39 ( .A(n1034), .ZN(n834) );
  INV_X1 U40 ( .A(n1024), .ZN(n833) );
  INV_X1 U41 ( .A(n1015), .ZN(n832) );
  INV_X1 U42 ( .A(n1006), .ZN(n831) );
  INV_X1 U43 ( .A(n997), .ZN(n830) );
  INV_X1 U44 ( .A(n961), .ZN(n826) );
  INV_X1 U45 ( .A(n951), .ZN(n825) );
  INV_X1 U46 ( .A(n942), .ZN(n824) );
  INV_X1 U47 ( .A(n933), .ZN(n823) );
  INV_X1 U48 ( .A(n924), .ZN(n822) );
  INV_X1 U49 ( .A(n1143), .ZN(n818) );
  BUF_X1 U50 ( .A(N11), .Z(n243) );
  BUF_X1 U51 ( .A(N11), .Z(n244) );
  BUF_X1 U52 ( .A(N11), .Z(n245) );
  INV_X1 U53 ( .A(N10), .ZN(n252) );
  BUF_X1 U54 ( .A(N12), .Z(n242) );
  NOR3_X1 U55 ( .A1(n254), .A2(N10), .A3(n253), .ZN(n1124) );
  NOR3_X1 U56 ( .A1(n254), .A2(n252), .A3(n253), .ZN(n1114) );
  NOR3_X1 U57 ( .A1(n252), .A2(N11), .A3(n254), .ZN(n1135) );
  NOR3_X1 U58 ( .A1(N10), .A2(N12), .A3(n253), .ZN(n1083) );
  NOR3_X1 U59 ( .A1(n252), .A2(N12), .A3(n253), .ZN(n1073) );
  NOR3_X1 U60 ( .A1(N10), .A2(N11), .A3(n254), .ZN(n1063) );
  NAND2_X1 U61 ( .A1(n1026), .A2(n1135), .ZN(n988) );
  NAND2_X1 U62 ( .A1(n953), .A2(n1135), .ZN(n915) );
  NAND2_X1 U63 ( .A1(n1026), .A2(n1063), .ZN(n997) );
  NAND2_X1 U64 ( .A1(n953), .A2(n1063), .ZN(n924) );
  NAND2_X1 U65 ( .A1(n1026), .A2(n1104), .ZN(n1034) );
  NAND2_X1 U66 ( .A1(n1026), .A2(n1093), .ZN(n1024) );
  NAND2_X1 U67 ( .A1(n953), .A2(n1104), .ZN(n961) );
  NAND2_X1 U68 ( .A1(n953), .A2(n1093), .ZN(n951) );
  NAND2_X1 U69 ( .A1(n1104), .A2(n1134), .ZN(n888) );
  NAND2_X1 U70 ( .A1(n1093), .A2(n1134), .ZN(n879) );
  NAND2_X1 U71 ( .A1(n1083), .A2(n1134), .ZN(n870) );
  NAND2_X1 U72 ( .A1(n1073), .A2(n1134), .ZN(n861) );
  NAND2_X1 U73 ( .A1(n1063), .A2(n1134), .ZN(n852) );
  NAND2_X1 U74 ( .A1(n1135), .A2(n1134), .ZN(n1143) );
  NAND2_X1 U75 ( .A1(n1124), .A2(n1134), .ZN(n1132) );
  NAND2_X1 U76 ( .A1(n1114), .A2(n1134), .ZN(n1122) );
  NAND2_X1 U77 ( .A1(n1026), .A2(n1083), .ZN(n1015) );
  NAND2_X1 U78 ( .A1(n1026), .A2(n1073), .ZN(n1006) );
  NAND2_X1 U79 ( .A1(n953), .A2(n1083), .ZN(n942) );
  NAND2_X1 U80 ( .A1(n953), .A2(n1073), .ZN(n933) );
  NAND2_X1 U81 ( .A1(n1026), .A2(n1124), .ZN(n979) );
  NAND2_X1 U82 ( .A1(n953), .A2(n1124), .ZN(n906) );
  NAND2_X1 U83 ( .A1(n1026), .A2(n1114), .ZN(n970) );
  NAND2_X1 U84 ( .A1(n953), .A2(n1114), .ZN(n897) );
  AND3_X1 U85 ( .A1(n843), .A2(n844), .A3(wr_en), .ZN(n1103) );
  AND3_X1 U86 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1134) );
  AND3_X1 U87 ( .A1(N13), .A2(n844), .A3(wr_en), .ZN(n1026) );
  AND3_X1 U88 ( .A1(N14), .A2(n843), .A3(wr_en), .ZN(n953) );
  INV_X1 U89 ( .A(n1062), .ZN(n770) );
  AOI22_X1 U90 ( .A1(data_in[0]), .A2(n837), .B1(n1061), .B2(\mem[5][0] ), 
        .ZN(n1062) );
  INV_X1 U91 ( .A(n1060), .ZN(n769) );
  AOI22_X1 U92 ( .A1(data_in[1]), .A2(n837), .B1(n1061), .B2(\mem[5][1] ), 
        .ZN(n1060) );
  INV_X1 U93 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U94 ( .A1(data_in[2]), .A2(n837), .B1(n1061), .B2(\mem[5][2] ), 
        .ZN(n1059) );
  INV_X1 U95 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U96 ( .A1(data_in[3]), .A2(n837), .B1(n1061), .B2(\mem[5][3] ), 
        .ZN(n1058) );
  INV_X1 U97 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U98 ( .A1(data_in[4]), .A2(n837), .B1(n1061), .B2(\mem[5][4] ), 
        .ZN(n1057) );
  INV_X1 U99 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U100 ( .A1(data_in[5]), .A2(n837), .B1(n1061), .B2(\mem[5][5] ), 
        .ZN(n1056) );
  INV_X1 U101 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U102 ( .A1(data_in[6]), .A2(n837), .B1(n1061), .B2(\mem[5][6] ), 
        .ZN(n1055) );
  INV_X1 U103 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U104 ( .A1(data_in[7]), .A2(n837), .B1(n1061), .B2(\mem[5][7] ), 
        .ZN(n1054) );
  INV_X1 U105 ( .A(n1025), .ZN(n738) );
  AOI22_X1 U106 ( .A1(data_in[0]), .A2(n833), .B1(n1024), .B2(\mem[9][0] ), 
        .ZN(n1025) );
  INV_X1 U107 ( .A(n1023), .ZN(n737) );
  AOI22_X1 U108 ( .A1(data_in[1]), .A2(n833), .B1(n1024), .B2(\mem[9][1] ), 
        .ZN(n1023) );
  INV_X1 U109 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U110 ( .A1(data_in[2]), .A2(n833), .B1(n1024), .B2(\mem[9][2] ), 
        .ZN(n1022) );
  INV_X1 U111 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U112 ( .A1(data_in[3]), .A2(n833), .B1(n1024), .B2(\mem[9][3] ), 
        .ZN(n1021) );
  INV_X1 U113 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U114 ( .A1(data_in[4]), .A2(n833), .B1(n1024), .B2(\mem[9][4] ), 
        .ZN(n1020) );
  INV_X1 U115 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U116 ( .A1(data_in[5]), .A2(n833), .B1(n1024), .B2(\mem[9][5] ), 
        .ZN(n1019) );
  INV_X1 U117 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U118 ( .A1(data_in[6]), .A2(n833), .B1(n1024), .B2(\mem[9][6] ), 
        .ZN(n1018) );
  INV_X1 U119 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U120 ( .A1(data_in[7]), .A2(n833), .B1(n1024), .B2(\mem[9][7] ), 
        .ZN(n1017) );
  INV_X1 U121 ( .A(n989), .ZN(n706) );
  AOI22_X1 U122 ( .A1(data_in[0]), .A2(n829), .B1(n988), .B2(\mem[13][0] ), 
        .ZN(n989) );
  INV_X1 U123 ( .A(n987), .ZN(n705) );
  AOI22_X1 U124 ( .A1(data_in[1]), .A2(n829), .B1(n988), .B2(\mem[13][1] ), 
        .ZN(n987) );
  INV_X1 U125 ( .A(n986), .ZN(n704) );
  AOI22_X1 U126 ( .A1(data_in[2]), .A2(n829), .B1(n988), .B2(\mem[13][2] ), 
        .ZN(n986) );
  INV_X1 U127 ( .A(n985), .ZN(n703) );
  AOI22_X1 U128 ( .A1(data_in[3]), .A2(n829), .B1(n988), .B2(\mem[13][3] ), 
        .ZN(n985) );
  INV_X1 U129 ( .A(n984), .ZN(n702) );
  AOI22_X1 U130 ( .A1(data_in[4]), .A2(n829), .B1(n988), .B2(\mem[13][4] ), 
        .ZN(n984) );
  INV_X1 U131 ( .A(n983), .ZN(n701) );
  AOI22_X1 U132 ( .A1(data_in[5]), .A2(n829), .B1(n988), .B2(\mem[13][5] ), 
        .ZN(n983) );
  INV_X1 U133 ( .A(n982), .ZN(n700) );
  AOI22_X1 U134 ( .A1(data_in[6]), .A2(n829), .B1(n988), .B2(\mem[13][6] ), 
        .ZN(n982) );
  INV_X1 U135 ( .A(n981), .ZN(n699) );
  AOI22_X1 U136 ( .A1(data_in[7]), .A2(n829), .B1(n988), .B2(\mem[13][7] ), 
        .ZN(n981) );
  INV_X1 U137 ( .A(n914), .ZN(n641) );
  AOI22_X1 U138 ( .A1(data_in[1]), .A2(n821), .B1(n915), .B2(\mem[21][1] ), 
        .ZN(n914) );
  INV_X1 U139 ( .A(n913), .ZN(n640) );
  AOI22_X1 U140 ( .A1(data_in[2]), .A2(n821), .B1(n915), .B2(\mem[21][2] ), 
        .ZN(n913) );
  INV_X1 U141 ( .A(n912), .ZN(n639) );
  AOI22_X1 U142 ( .A1(data_in[3]), .A2(n821), .B1(n915), .B2(\mem[21][3] ), 
        .ZN(n912) );
  INV_X1 U143 ( .A(n911), .ZN(n638) );
  AOI22_X1 U144 ( .A1(data_in[4]), .A2(n821), .B1(n915), .B2(\mem[21][4] ), 
        .ZN(n911) );
  INV_X1 U145 ( .A(n910), .ZN(n637) );
  AOI22_X1 U146 ( .A1(data_in[5]), .A2(n821), .B1(n915), .B2(\mem[21][5] ), 
        .ZN(n910) );
  INV_X1 U147 ( .A(n909), .ZN(n636) );
  AOI22_X1 U148 ( .A1(data_in[6]), .A2(n821), .B1(n915), .B2(\mem[21][6] ), 
        .ZN(n909) );
  INV_X1 U149 ( .A(n908), .ZN(n635) );
  AOI22_X1 U150 ( .A1(data_in[7]), .A2(n821), .B1(n915), .B2(\mem[21][7] ), 
        .ZN(n908) );
  INV_X1 U151 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U152 ( .A1(data_in[6]), .A2(n832), .B1(n1015), .B2(\mem[10][6] ), 
        .ZN(n1009) );
  INV_X1 U153 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U154 ( .A1(data_in[7]), .A2(n832), .B1(n1015), .B2(\mem[10][7] ), 
        .ZN(n1008) );
  INV_X1 U155 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U156 ( .A1(data_in[0]), .A2(n831), .B1(n1006), .B2(\mem[11][0] ), 
        .ZN(n1007) );
  INV_X1 U157 ( .A(n1005), .ZN(n721) );
  AOI22_X1 U158 ( .A1(data_in[1]), .A2(n831), .B1(n1006), .B2(\mem[11][1] ), 
        .ZN(n1005) );
  INV_X1 U159 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U160 ( .A1(data_in[2]), .A2(n831), .B1(n1006), .B2(\mem[11][2] ), 
        .ZN(n1004) );
  INV_X1 U161 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U162 ( .A1(data_in[3]), .A2(n831), .B1(n1006), .B2(\mem[11][3] ), 
        .ZN(n1003) );
  INV_X1 U163 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U164 ( .A1(data_in[4]), .A2(n831), .B1(n1006), .B2(\mem[11][4] ), 
        .ZN(n1002) );
  INV_X1 U165 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U166 ( .A1(data_in[5]), .A2(n831), .B1(n1006), .B2(\mem[11][5] ), 
        .ZN(n1001) );
  INV_X1 U167 ( .A(n952), .ZN(n674) );
  AOI22_X1 U168 ( .A1(data_in[0]), .A2(n825), .B1(n951), .B2(\mem[17][0] ), 
        .ZN(n952) );
  INV_X1 U169 ( .A(n950), .ZN(n673) );
  AOI22_X1 U170 ( .A1(data_in[1]), .A2(n825), .B1(n951), .B2(\mem[17][1] ), 
        .ZN(n950) );
  INV_X1 U171 ( .A(n949), .ZN(n672) );
  AOI22_X1 U172 ( .A1(data_in[2]), .A2(n825), .B1(n951), .B2(\mem[17][2] ), 
        .ZN(n949) );
  INV_X1 U173 ( .A(n948), .ZN(n671) );
  AOI22_X1 U174 ( .A1(data_in[3]), .A2(n825), .B1(n951), .B2(\mem[17][3] ), 
        .ZN(n948) );
  INV_X1 U175 ( .A(n947), .ZN(n670) );
  AOI22_X1 U176 ( .A1(data_in[4]), .A2(n825), .B1(n951), .B2(\mem[17][4] ), 
        .ZN(n947) );
  INV_X1 U177 ( .A(n946), .ZN(n669) );
  AOI22_X1 U178 ( .A1(data_in[5]), .A2(n825), .B1(n951), .B2(\mem[17][5] ), 
        .ZN(n946) );
  INV_X1 U179 ( .A(n945), .ZN(n668) );
  AOI22_X1 U180 ( .A1(data_in[6]), .A2(n825), .B1(n951), .B2(\mem[17][6] ), 
        .ZN(n945) );
  INV_X1 U181 ( .A(n944), .ZN(n667) );
  AOI22_X1 U182 ( .A1(data_in[7]), .A2(n825), .B1(n951), .B2(\mem[17][7] ), 
        .ZN(n944) );
  INV_X1 U183 ( .A(n916), .ZN(n642) );
  AOI22_X1 U184 ( .A1(data_in[0]), .A2(n821), .B1(n915), .B2(\mem[21][0] ), 
        .ZN(n916) );
  INV_X1 U185 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U186 ( .A1(data_in[6]), .A2(n831), .B1(n1006), .B2(\mem[11][6] ), 
        .ZN(n1000) );
  INV_X1 U187 ( .A(n999), .ZN(n715) );
  AOI22_X1 U188 ( .A1(data_in[7]), .A2(n831), .B1(n1006), .B2(\mem[11][7] ), 
        .ZN(n999) );
  INV_X1 U189 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U190 ( .A1(data_in[0]), .A2(n836), .B1(n1052), .B2(\mem[6][0] ), 
        .ZN(n1053) );
  INV_X1 U191 ( .A(n1051), .ZN(n761) );
  AOI22_X1 U192 ( .A1(data_in[1]), .A2(n836), .B1(n1052), .B2(\mem[6][1] ), 
        .ZN(n1051) );
  INV_X1 U193 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U194 ( .A1(data_in[2]), .A2(n836), .B1(n1052), .B2(\mem[6][2] ), 
        .ZN(n1050) );
  INV_X1 U195 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U196 ( .A1(data_in[3]), .A2(n836), .B1(n1052), .B2(\mem[6][3] ), 
        .ZN(n1049) );
  INV_X1 U197 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U198 ( .A1(data_in[4]), .A2(n836), .B1(n1052), .B2(\mem[6][4] ), 
        .ZN(n1048) );
  INV_X1 U199 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U200 ( .A1(data_in[5]), .A2(n836), .B1(n1052), .B2(\mem[6][5] ), 
        .ZN(n1047) );
  INV_X1 U201 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U202 ( .A1(data_in[6]), .A2(n836), .B1(n1052), .B2(\mem[6][6] ), 
        .ZN(n1046) );
  INV_X1 U203 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U204 ( .A1(data_in[7]), .A2(n836), .B1(n1052), .B2(\mem[6][7] ), 
        .ZN(n1045) );
  INV_X1 U205 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U206 ( .A1(data_in[0]), .A2(n835), .B1(n1043), .B2(\mem[7][0] ), 
        .ZN(n1044) );
  INV_X1 U207 ( .A(n1042), .ZN(n753) );
  AOI22_X1 U208 ( .A1(data_in[1]), .A2(n835), .B1(n1043), .B2(\mem[7][1] ), 
        .ZN(n1042) );
  INV_X1 U209 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U210 ( .A1(data_in[2]), .A2(n835), .B1(n1043), .B2(\mem[7][2] ), 
        .ZN(n1041) );
  INV_X1 U211 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U212 ( .A1(data_in[3]), .A2(n835), .B1(n1043), .B2(\mem[7][3] ), 
        .ZN(n1040) );
  INV_X1 U213 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U214 ( .A1(data_in[4]), .A2(n835), .B1(n1043), .B2(\mem[7][4] ), 
        .ZN(n1039) );
  INV_X1 U215 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U216 ( .A1(data_in[5]), .A2(n835), .B1(n1043), .B2(\mem[7][5] ), 
        .ZN(n1038) );
  INV_X1 U217 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U218 ( .A1(data_in[6]), .A2(n835), .B1(n1043), .B2(\mem[7][6] ), 
        .ZN(n1037) );
  INV_X1 U219 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U220 ( .A1(data_in[7]), .A2(n835), .B1(n1043), .B2(\mem[7][7] ), 
        .ZN(n1036) );
  INV_X1 U221 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U222 ( .A1(data_in[0]), .A2(n832), .B1(n1015), .B2(\mem[10][0] ), 
        .ZN(n1016) );
  INV_X1 U223 ( .A(n1014), .ZN(n729) );
  AOI22_X1 U224 ( .A1(data_in[1]), .A2(n832), .B1(n1015), .B2(\mem[10][1] ), 
        .ZN(n1014) );
  INV_X1 U225 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U226 ( .A1(data_in[2]), .A2(n832), .B1(n1015), .B2(\mem[10][2] ), 
        .ZN(n1013) );
  INV_X1 U227 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U228 ( .A1(data_in[3]), .A2(n832), .B1(n1015), .B2(\mem[10][3] ), 
        .ZN(n1012) );
  INV_X1 U229 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U230 ( .A1(data_in[4]), .A2(n832), .B1(n1015), .B2(\mem[10][4] ), 
        .ZN(n1011) );
  INV_X1 U231 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U232 ( .A1(data_in[5]), .A2(n832), .B1(n1015), .B2(\mem[10][5] ), 
        .ZN(n1010) );
  INV_X1 U233 ( .A(n980), .ZN(n698) );
  AOI22_X1 U234 ( .A1(data_in[0]), .A2(n828), .B1(n979), .B2(\mem[14][0] ), 
        .ZN(n980) );
  INV_X1 U235 ( .A(n978), .ZN(n697) );
  AOI22_X1 U236 ( .A1(data_in[1]), .A2(n828), .B1(n979), .B2(\mem[14][1] ), 
        .ZN(n978) );
  INV_X1 U237 ( .A(n977), .ZN(n696) );
  AOI22_X1 U238 ( .A1(data_in[2]), .A2(n828), .B1(n979), .B2(\mem[14][2] ), 
        .ZN(n977) );
  INV_X1 U239 ( .A(n976), .ZN(n695) );
  AOI22_X1 U240 ( .A1(data_in[3]), .A2(n828), .B1(n979), .B2(\mem[14][3] ), 
        .ZN(n976) );
  INV_X1 U241 ( .A(n975), .ZN(n694) );
  AOI22_X1 U242 ( .A1(data_in[4]), .A2(n828), .B1(n979), .B2(\mem[14][4] ), 
        .ZN(n975) );
  INV_X1 U243 ( .A(n974), .ZN(n693) );
  AOI22_X1 U244 ( .A1(data_in[5]), .A2(n828), .B1(n979), .B2(\mem[14][5] ), 
        .ZN(n974) );
  INV_X1 U245 ( .A(n973), .ZN(n692) );
  AOI22_X1 U246 ( .A1(data_in[6]), .A2(n828), .B1(n979), .B2(\mem[14][6] ), 
        .ZN(n973) );
  INV_X1 U247 ( .A(n972), .ZN(n691) );
  AOI22_X1 U248 ( .A1(data_in[7]), .A2(n828), .B1(n979), .B2(\mem[14][7] ), 
        .ZN(n972) );
  INV_X1 U249 ( .A(n971), .ZN(n690) );
  AOI22_X1 U250 ( .A1(data_in[0]), .A2(n827), .B1(n970), .B2(\mem[15][0] ), 
        .ZN(n971) );
  INV_X1 U251 ( .A(n969), .ZN(n689) );
  AOI22_X1 U252 ( .A1(data_in[1]), .A2(n827), .B1(n970), .B2(\mem[15][1] ), 
        .ZN(n969) );
  INV_X1 U253 ( .A(n968), .ZN(n688) );
  AOI22_X1 U254 ( .A1(data_in[2]), .A2(n827), .B1(n970), .B2(\mem[15][2] ), 
        .ZN(n968) );
  INV_X1 U255 ( .A(n967), .ZN(n687) );
  AOI22_X1 U256 ( .A1(data_in[3]), .A2(n827), .B1(n970), .B2(\mem[15][3] ), 
        .ZN(n967) );
  INV_X1 U257 ( .A(n966), .ZN(n686) );
  AOI22_X1 U258 ( .A1(data_in[4]), .A2(n827), .B1(n970), .B2(\mem[15][4] ), 
        .ZN(n966) );
  INV_X1 U259 ( .A(n965), .ZN(n685) );
  AOI22_X1 U260 ( .A1(data_in[5]), .A2(n827), .B1(n970), .B2(\mem[15][5] ), 
        .ZN(n965) );
  INV_X1 U261 ( .A(n964), .ZN(n684) );
  AOI22_X1 U262 ( .A1(data_in[6]), .A2(n827), .B1(n970), .B2(\mem[15][6] ), 
        .ZN(n964) );
  INV_X1 U263 ( .A(n963), .ZN(n683) );
  AOI22_X1 U264 ( .A1(data_in[7]), .A2(n827), .B1(n970), .B2(\mem[15][7] ), 
        .ZN(n963) );
  INV_X1 U265 ( .A(n943), .ZN(n666) );
  AOI22_X1 U266 ( .A1(data_in[0]), .A2(n824), .B1(n942), .B2(\mem[18][0] ), 
        .ZN(n943) );
  INV_X1 U267 ( .A(n941), .ZN(n665) );
  AOI22_X1 U268 ( .A1(data_in[1]), .A2(n824), .B1(n942), .B2(\mem[18][1] ), 
        .ZN(n941) );
  INV_X1 U269 ( .A(n940), .ZN(n664) );
  AOI22_X1 U270 ( .A1(data_in[2]), .A2(n824), .B1(n942), .B2(\mem[18][2] ), 
        .ZN(n940) );
  INV_X1 U271 ( .A(n939), .ZN(n663) );
  AOI22_X1 U272 ( .A1(data_in[3]), .A2(n824), .B1(n942), .B2(\mem[18][3] ), 
        .ZN(n939) );
  INV_X1 U273 ( .A(n938), .ZN(n662) );
  AOI22_X1 U274 ( .A1(data_in[4]), .A2(n824), .B1(n942), .B2(\mem[18][4] ), 
        .ZN(n938) );
  INV_X1 U275 ( .A(n937), .ZN(n661) );
  AOI22_X1 U276 ( .A1(data_in[5]), .A2(n824), .B1(n942), .B2(\mem[18][5] ), 
        .ZN(n937) );
  INV_X1 U277 ( .A(n936), .ZN(n660) );
  AOI22_X1 U278 ( .A1(data_in[6]), .A2(n824), .B1(n942), .B2(\mem[18][6] ), 
        .ZN(n936) );
  INV_X1 U279 ( .A(n935), .ZN(n659) );
  AOI22_X1 U280 ( .A1(data_in[7]), .A2(n824), .B1(n942), .B2(\mem[18][7] ), 
        .ZN(n935) );
  INV_X1 U281 ( .A(n934), .ZN(n658) );
  AOI22_X1 U282 ( .A1(data_in[0]), .A2(n823), .B1(n933), .B2(\mem[19][0] ), 
        .ZN(n934) );
  INV_X1 U283 ( .A(n932), .ZN(n657) );
  AOI22_X1 U284 ( .A1(data_in[1]), .A2(n823), .B1(n933), .B2(\mem[19][1] ), 
        .ZN(n932) );
  INV_X1 U285 ( .A(n931), .ZN(n656) );
  AOI22_X1 U286 ( .A1(data_in[2]), .A2(n823), .B1(n933), .B2(\mem[19][2] ), 
        .ZN(n931) );
  INV_X1 U287 ( .A(n930), .ZN(n655) );
  AOI22_X1 U288 ( .A1(data_in[3]), .A2(n823), .B1(n933), .B2(\mem[19][3] ), 
        .ZN(n930) );
  INV_X1 U289 ( .A(n929), .ZN(n654) );
  AOI22_X1 U290 ( .A1(data_in[4]), .A2(n823), .B1(n933), .B2(\mem[19][4] ), 
        .ZN(n929) );
  INV_X1 U291 ( .A(n928), .ZN(n653) );
  AOI22_X1 U292 ( .A1(data_in[5]), .A2(n823), .B1(n933), .B2(\mem[19][5] ), 
        .ZN(n928) );
  INV_X1 U293 ( .A(n927), .ZN(n652) );
  AOI22_X1 U294 ( .A1(data_in[6]), .A2(n823), .B1(n933), .B2(\mem[19][6] ), 
        .ZN(n927) );
  INV_X1 U295 ( .A(n926), .ZN(n651) );
  AOI22_X1 U296 ( .A1(data_in[7]), .A2(n823), .B1(n933), .B2(\mem[19][7] ), 
        .ZN(n926) );
  INV_X1 U297 ( .A(n907), .ZN(n634) );
  AOI22_X1 U298 ( .A1(data_in[0]), .A2(n820), .B1(n906), .B2(\mem[22][0] ), 
        .ZN(n907) );
  INV_X1 U299 ( .A(n905), .ZN(n633) );
  AOI22_X1 U300 ( .A1(data_in[1]), .A2(n820), .B1(n906), .B2(\mem[22][1] ), 
        .ZN(n905) );
  INV_X1 U301 ( .A(n904), .ZN(n632) );
  AOI22_X1 U302 ( .A1(data_in[2]), .A2(n820), .B1(n906), .B2(\mem[22][2] ), 
        .ZN(n904) );
  INV_X1 U303 ( .A(n903), .ZN(n631) );
  AOI22_X1 U304 ( .A1(data_in[3]), .A2(n820), .B1(n906), .B2(\mem[22][3] ), 
        .ZN(n903) );
  INV_X1 U305 ( .A(n902), .ZN(n630) );
  AOI22_X1 U306 ( .A1(data_in[4]), .A2(n820), .B1(n906), .B2(\mem[22][4] ), 
        .ZN(n902) );
  INV_X1 U307 ( .A(n901), .ZN(n629) );
  AOI22_X1 U308 ( .A1(data_in[5]), .A2(n820), .B1(n906), .B2(\mem[22][5] ), 
        .ZN(n901) );
  INV_X1 U309 ( .A(n900), .ZN(n628) );
  AOI22_X1 U310 ( .A1(data_in[6]), .A2(n820), .B1(n906), .B2(\mem[22][6] ), 
        .ZN(n900) );
  INV_X1 U311 ( .A(n899), .ZN(n627) );
  AOI22_X1 U312 ( .A1(data_in[7]), .A2(n820), .B1(n906), .B2(\mem[22][7] ), 
        .ZN(n899) );
  INV_X1 U313 ( .A(n898), .ZN(n626) );
  AOI22_X1 U314 ( .A1(data_in[0]), .A2(n819), .B1(n897), .B2(\mem[23][0] ), 
        .ZN(n898) );
  INV_X1 U315 ( .A(n896), .ZN(n625) );
  AOI22_X1 U316 ( .A1(data_in[1]), .A2(n819), .B1(n897), .B2(\mem[23][1] ), 
        .ZN(n896) );
  INV_X1 U317 ( .A(n895), .ZN(n624) );
  AOI22_X1 U318 ( .A1(data_in[2]), .A2(n819), .B1(n897), .B2(\mem[23][2] ), 
        .ZN(n895) );
  INV_X1 U319 ( .A(n894), .ZN(n623) );
  AOI22_X1 U320 ( .A1(data_in[3]), .A2(n819), .B1(n897), .B2(\mem[23][3] ), 
        .ZN(n894) );
  INV_X1 U321 ( .A(n893), .ZN(n622) );
  AOI22_X1 U322 ( .A1(data_in[4]), .A2(n819), .B1(n897), .B2(\mem[23][4] ), 
        .ZN(n893) );
  INV_X1 U323 ( .A(n892), .ZN(n621) );
  AOI22_X1 U324 ( .A1(data_in[5]), .A2(n819), .B1(n897), .B2(\mem[23][5] ), 
        .ZN(n892) );
  INV_X1 U325 ( .A(n891), .ZN(n620) );
  AOI22_X1 U326 ( .A1(data_in[6]), .A2(n819), .B1(n897), .B2(\mem[23][6] ), 
        .ZN(n891) );
  INV_X1 U327 ( .A(n890), .ZN(n619) );
  AOI22_X1 U328 ( .A1(data_in[7]), .A2(n819), .B1(n897), .B2(\mem[23][7] ), 
        .ZN(n890) );
  INV_X1 U329 ( .A(N12), .ZN(n254) );
  INV_X1 U330 ( .A(N11), .ZN(n253) );
  INV_X1 U331 ( .A(n998), .ZN(n714) );
  AOI22_X1 U332 ( .A1(data_in[0]), .A2(n830), .B1(n997), .B2(\mem[12][0] ), 
        .ZN(n998) );
  INV_X1 U333 ( .A(n996), .ZN(n713) );
  AOI22_X1 U334 ( .A1(data_in[1]), .A2(n830), .B1(n997), .B2(\mem[12][1] ), 
        .ZN(n996) );
  INV_X1 U335 ( .A(n995), .ZN(n712) );
  AOI22_X1 U336 ( .A1(data_in[2]), .A2(n830), .B1(n997), .B2(\mem[12][2] ), 
        .ZN(n995) );
  INV_X1 U337 ( .A(n994), .ZN(n711) );
  AOI22_X1 U338 ( .A1(data_in[3]), .A2(n830), .B1(n997), .B2(\mem[12][3] ), 
        .ZN(n994) );
  INV_X1 U339 ( .A(n993), .ZN(n710) );
  AOI22_X1 U340 ( .A1(data_in[4]), .A2(n830), .B1(n997), .B2(\mem[12][4] ), 
        .ZN(n993) );
  INV_X1 U341 ( .A(n992), .ZN(n709) );
  AOI22_X1 U342 ( .A1(data_in[5]), .A2(n830), .B1(n997), .B2(\mem[12][5] ), 
        .ZN(n992) );
  INV_X1 U343 ( .A(n991), .ZN(n708) );
  AOI22_X1 U344 ( .A1(data_in[6]), .A2(n830), .B1(n997), .B2(\mem[12][6] ), 
        .ZN(n991) );
  INV_X1 U345 ( .A(n990), .ZN(n707) );
  AOI22_X1 U346 ( .A1(data_in[7]), .A2(n830), .B1(n997), .B2(\mem[12][7] ), 
        .ZN(n990) );
  INV_X1 U347 ( .A(n925), .ZN(n650) );
  AOI22_X1 U348 ( .A1(data_in[0]), .A2(n822), .B1(n924), .B2(\mem[20][0] ), 
        .ZN(n925) );
  INV_X1 U349 ( .A(n923), .ZN(n649) );
  AOI22_X1 U350 ( .A1(data_in[1]), .A2(n822), .B1(n924), .B2(\mem[20][1] ), 
        .ZN(n923) );
  INV_X1 U351 ( .A(n922), .ZN(n648) );
  AOI22_X1 U352 ( .A1(data_in[2]), .A2(n822), .B1(n924), .B2(\mem[20][2] ), 
        .ZN(n922) );
  INV_X1 U353 ( .A(n921), .ZN(n647) );
  AOI22_X1 U354 ( .A1(data_in[3]), .A2(n822), .B1(n924), .B2(\mem[20][3] ), 
        .ZN(n921) );
  INV_X1 U355 ( .A(n920), .ZN(n646) );
  AOI22_X1 U356 ( .A1(data_in[4]), .A2(n822), .B1(n924), .B2(\mem[20][4] ), 
        .ZN(n920) );
  INV_X1 U357 ( .A(n919), .ZN(n645) );
  AOI22_X1 U358 ( .A1(data_in[5]), .A2(n822), .B1(n924), .B2(\mem[20][5] ), 
        .ZN(n919) );
  INV_X1 U359 ( .A(n918), .ZN(n644) );
  AOI22_X1 U360 ( .A1(data_in[6]), .A2(n822), .B1(n924), .B2(\mem[20][6] ), 
        .ZN(n918) );
  INV_X1 U361 ( .A(n917), .ZN(n643) );
  AOI22_X1 U362 ( .A1(data_in[7]), .A2(n822), .B1(n924), .B2(\mem[20][7] ), 
        .ZN(n917) );
  INV_X1 U363 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U364 ( .A1(data_in[0]), .A2(n834), .B1(n1034), .B2(\mem[8][0] ), 
        .ZN(n1035) );
  INV_X1 U365 ( .A(n1033), .ZN(n745) );
  AOI22_X1 U366 ( .A1(data_in[1]), .A2(n834), .B1(n1034), .B2(\mem[8][1] ), 
        .ZN(n1033) );
  INV_X1 U367 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U368 ( .A1(data_in[2]), .A2(n834), .B1(n1034), .B2(\mem[8][2] ), 
        .ZN(n1032) );
  INV_X1 U369 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U370 ( .A1(data_in[3]), .A2(n834), .B1(n1034), .B2(\mem[8][3] ), 
        .ZN(n1031) );
  INV_X1 U371 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U372 ( .A1(data_in[4]), .A2(n834), .B1(n1034), .B2(\mem[8][4] ), 
        .ZN(n1030) );
  INV_X1 U373 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U374 ( .A1(data_in[5]), .A2(n834), .B1(n1034), .B2(\mem[8][5] ), 
        .ZN(n1029) );
  INV_X1 U375 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U376 ( .A1(data_in[6]), .A2(n834), .B1(n1034), .B2(\mem[8][6] ), 
        .ZN(n1028) );
  INV_X1 U377 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U378 ( .A1(data_in[7]), .A2(n834), .B1(n1034), .B2(\mem[8][7] ), 
        .ZN(n1027) );
  INV_X1 U379 ( .A(n962), .ZN(n682) );
  AOI22_X1 U380 ( .A1(data_in[0]), .A2(n826), .B1(n961), .B2(\mem[16][0] ), 
        .ZN(n962) );
  INV_X1 U381 ( .A(n960), .ZN(n681) );
  AOI22_X1 U382 ( .A1(data_in[1]), .A2(n826), .B1(n961), .B2(\mem[16][1] ), 
        .ZN(n960) );
  INV_X1 U383 ( .A(n959), .ZN(n680) );
  AOI22_X1 U384 ( .A1(data_in[2]), .A2(n826), .B1(n961), .B2(\mem[16][2] ), 
        .ZN(n959) );
  INV_X1 U385 ( .A(n958), .ZN(n679) );
  AOI22_X1 U386 ( .A1(data_in[3]), .A2(n826), .B1(n961), .B2(\mem[16][3] ), 
        .ZN(n958) );
  INV_X1 U387 ( .A(n957), .ZN(n678) );
  AOI22_X1 U388 ( .A1(data_in[4]), .A2(n826), .B1(n961), .B2(\mem[16][4] ), 
        .ZN(n957) );
  INV_X1 U389 ( .A(n956), .ZN(n677) );
  AOI22_X1 U390 ( .A1(data_in[5]), .A2(n826), .B1(n961), .B2(\mem[16][5] ), 
        .ZN(n956) );
  INV_X1 U391 ( .A(n955), .ZN(n676) );
  AOI22_X1 U392 ( .A1(data_in[6]), .A2(n826), .B1(n961), .B2(\mem[16][6] ), 
        .ZN(n955) );
  INV_X1 U393 ( .A(n954), .ZN(n675) );
  AOI22_X1 U394 ( .A1(data_in[7]), .A2(n826), .B1(n961), .B2(\mem[16][7] ), 
        .ZN(n954) );
  INV_X1 U395 ( .A(n889), .ZN(n618) );
  AOI22_X1 U396 ( .A1(data_in[0]), .A2(n815), .B1(n888), .B2(\mem[24][0] ), 
        .ZN(n889) );
  INV_X1 U397 ( .A(n887), .ZN(n617) );
  AOI22_X1 U398 ( .A1(data_in[1]), .A2(n815), .B1(n888), .B2(\mem[24][1] ), 
        .ZN(n887) );
  INV_X1 U399 ( .A(n886), .ZN(n616) );
  AOI22_X1 U400 ( .A1(data_in[2]), .A2(n815), .B1(n888), .B2(\mem[24][2] ), 
        .ZN(n886) );
  INV_X1 U401 ( .A(n885), .ZN(n615) );
  AOI22_X1 U402 ( .A1(data_in[3]), .A2(n815), .B1(n888), .B2(\mem[24][3] ), 
        .ZN(n885) );
  INV_X1 U403 ( .A(n884), .ZN(n614) );
  AOI22_X1 U404 ( .A1(data_in[4]), .A2(n815), .B1(n888), .B2(\mem[24][4] ), 
        .ZN(n884) );
  INV_X1 U405 ( .A(n883), .ZN(n613) );
  AOI22_X1 U406 ( .A1(data_in[5]), .A2(n815), .B1(n888), .B2(\mem[24][5] ), 
        .ZN(n883) );
  INV_X1 U407 ( .A(n882), .ZN(n612) );
  AOI22_X1 U408 ( .A1(data_in[6]), .A2(n815), .B1(n888), .B2(\mem[24][6] ), 
        .ZN(n882) );
  INV_X1 U409 ( .A(n881), .ZN(n611) );
  AOI22_X1 U410 ( .A1(data_in[7]), .A2(n815), .B1(n888), .B2(\mem[24][7] ), 
        .ZN(n881) );
  INV_X1 U411 ( .A(n880), .ZN(n610) );
  AOI22_X1 U412 ( .A1(data_in[0]), .A2(n814), .B1(n879), .B2(\mem[25][0] ), 
        .ZN(n880) );
  INV_X1 U413 ( .A(n878), .ZN(n609) );
  AOI22_X1 U414 ( .A1(data_in[1]), .A2(n814), .B1(n879), .B2(\mem[25][1] ), 
        .ZN(n878) );
  INV_X1 U415 ( .A(n877), .ZN(n608) );
  AOI22_X1 U416 ( .A1(data_in[2]), .A2(n814), .B1(n879), .B2(\mem[25][2] ), 
        .ZN(n877) );
  INV_X1 U417 ( .A(n876), .ZN(n607) );
  AOI22_X1 U418 ( .A1(data_in[3]), .A2(n814), .B1(n879), .B2(\mem[25][3] ), 
        .ZN(n876) );
  INV_X1 U419 ( .A(n875), .ZN(n606) );
  AOI22_X1 U420 ( .A1(data_in[4]), .A2(n814), .B1(n879), .B2(\mem[25][4] ), 
        .ZN(n875) );
  INV_X1 U421 ( .A(n874), .ZN(n605) );
  AOI22_X1 U422 ( .A1(data_in[5]), .A2(n814), .B1(n879), .B2(\mem[25][5] ), 
        .ZN(n874) );
  INV_X1 U423 ( .A(n873), .ZN(n604) );
  AOI22_X1 U424 ( .A1(data_in[6]), .A2(n814), .B1(n879), .B2(\mem[25][6] ), 
        .ZN(n873) );
  INV_X1 U425 ( .A(n872), .ZN(n603) );
  AOI22_X1 U426 ( .A1(data_in[7]), .A2(n814), .B1(n879), .B2(\mem[25][7] ), 
        .ZN(n872) );
  INV_X1 U427 ( .A(n871), .ZN(n602) );
  AOI22_X1 U428 ( .A1(data_in[0]), .A2(n813), .B1(n870), .B2(\mem[26][0] ), 
        .ZN(n871) );
  INV_X1 U429 ( .A(n869), .ZN(n601) );
  AOI22_X1 U430 ( .A1(data_in[1]), .A2(n813), .B1(n870), .B2(\mem[26][1] ), 
        .ZN(n869) );
  INV_X1 U431 ( .A(n868), .ZN(n600) );
  AOI22_X1 U432 ( .A1(data_in[2]), .A2(n813), .B1(n870), .B2(\mem[26][2] ), 
        .ZN(n868) );
  INV_X1 U433 ( .A(n867), .ZN(n599) );
  AOI22_X1 U434 ( .A1(data_in[3]), .A2(n813), .B1(n870), .B2(\mem[26][3] ), 
        .ZN(n867) );
  INV_X1 U435 ( .A(n866), .ZN(n598) );
  AOI22_X1 U436 ( .A1(data_in[4]), .A2(n813), .B1(n870), .B2(\mem[26][4] ), 
        .ZN(n866) );
  INV_X1 U437 ( .A(n865), .ZN(n597) );
  AOI22_X1 U438 ( .A1(data_in[5]), .A2(n813), .B1(n870), .B2(\mem[26][5] ), 
        .ZN(n865) );
  INV_X1 U439 ( .A(n864), .ZN(n596) );
  AOI22_X1 U440 ( .A1(data_in[6]), .A2(n813), .B1(n870), .B2(\mem[26][6] ), 
        .ZN(n864) );
  INV_X1 U441 ( .A(n863), .ZN(n595) );
  AOI22_X1 U442 ( .A1(data_in[7]), .A2(n813), .B1(n870), .B2(\mem[26][7] ), 
        .ZN(n863) );
  INV_X1 U443 ( .A(n862), .ZN(n594) );
  AOI22_X1 U444 ( .A1(data_in[0]), .A2(n812), .B1(n861), .B2(\mem[27][0] ), 
        .ZN(n862) );
  INV_X1 U445 ( .A(n860), .ZN(n293) );
  AOI22_X1 U446 ( .A1(data_in[1]), .A2(n812), .B1(n861), .B2(\mem[27][1] ), 
        .ZN(n860) );
  INV_X1 U447 ( .A(n859), .ZN(n292) );
  AOI22_X1 U448 ( .A1(data_in[2]), .A2(n812), .B1(n861), .B2(\mem[27][2] ), 
        .ZN(n859) );
  INV_X1 U449 ( .A(n858), .ZN(n291) );
  AOI22_X1 U450 ( .A1(data_in[3]), .A2(n812), .B1(n861), .B2(\mem[27][3] ), 
        .ZN(n858) );
  INV_X1 U451 ( .A(n857), .ZN(n290) );
  AOI22_X1 U452 ( .A1(data_in[4]), .A2(n812), .B1(n861), .B2(\mem[27][4] ), 
        .ZN(n857) );
  INV_X1 U453 ( .A(n856), .ZN(n289) );
  AOI22_X1 U454 ( .A1(data_in[5]), .A2(n812), .B1(n861), .B2(\mem[27][5] ), 
        .ZN(n856) );
  INV_X1 U455 ( .A(n855), .ZN(n288) );
  AOI22_X1 U456 ( .A1(data_in[6]), .A2(n812), .B1(n861), .B2(\mem[27][6] ), 
        .ZN(n855) );
  INV_X1 U457 ( .A(n854), .ZN(n287) );
  AOI22_X1 U458 ( .A1(data_in[7]), .A2(n812), .B1(n861), .B2(\mem[27][7] ), 
        .ZN(n854) );
  INV_X1 U459 ( .A(n853), .ZN(n286) );
  AOI22_X1 U460 ( .A1(data_in[0]), .A2(n811), .B1(n852), .B2(\mem[28][0] ), 
        .ZN(n853) );
  INV_X1 U461 ( .A(n851), .ZN(n285) );
  AOI22_X1 U462 ( .A1(data_in[1]), .A2(n811), .B1(n852), .B2(\mem[28][1] ), 
        .ZN(n851) );
  INV_X1 U463 ( .A(n850), .ZN(n284) );
  AOI22_X1 U464 ( .A1(data_in[2]), .A2(n811), .B1(n852), .B2(\mem[28][2] ), 
        .ZN(n850) );
  INV_X1 U465 ( .A(n849), .ZN(n283) );
  AOI22_X1 U466 ( .A1(data_in[3]), .A2(n811), .B1(n852), .B2(\mem[28][3] ), 
        .ZN(n849) );
  INV_X1 U467 ( .A(n848), .ZN(n282) );
  AOI22_X1 U468 ( .A1(data_in[4]), .A2(n811), .B1(n852), .B2(\mem[28][4] ), 
        .ZN(n848) );
  INV_X1 U469 ( .A(n847), .ZN(n281) );
  AOI22_X1 U470 ( .A1(data_in[5]), .A2(n811), .B1(n852), .B2(\mem[28][5] ), 
        .ZN(n847) );
  INV_X1 U471 ( .A(n846), .ZN(n280) );
  AOI22_X1 U472 ( .A1(data_in[6]), .A2(n811), .B1(n852), .B2(\mem[28][6] ), 
        .ZN(n846) );
  INV_X1 U473 ( .A(n845), .ZN(n279) );
  AOI22_X1 U474 ( .A1(data_in[7]), .A2(n811), .B1(n852), .B2(\mem[28][7] ), 
        .ZN(n845) );
  INV_X1 U475 ( .A(n1144), .ZN(n278) );
  AOI22_X1 U476 ( .A1(n818), .A2(data_in[0]), .B1(n1143), .B2(\mem[29][0] ), 
        .ZN(n1144) );
  INV_X1 U477 ( .A(n1142), .ZN(n277) );
  AOI22_X1 U478 ( .A1(n818), .A2(data_in[1]), .B1(n1143), .B2(\mem[29][1] ), 
        .ZN(n1142) );
  INV_X1 U479 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U480 ( .A1(n818), .A2(data_in[2]), .B1(n1143), .B2(\mem[29][2] ), 
        .ZN(n1141) );
  INV_X1 U481 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U482 ( .A1(n818), .A2(data_in[3]), .B1(n1143), .B2(\mem[29][3] ), 
        .ZN(n1140) );
  INV_X1 U483 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U484 ( .A1(n818), .A2(data_in[4]), .B1(n1143), .B2(\mem[29][4] ), 
        .ZN(n1139) );
  INV_X1 U485 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U486 ( .A1(n818), .A2(data_in[5]), .B1(n1143), .B2(\mem[29][5] ), 
        .ZN(n1138) );
  INV_X1 U487 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U488 ( .A1(n818), .A2(data_in[6]), .B1(n1143), .B2(\mem[29][6] ), 
        .ZN(n1137) );
  INV_X1 U489 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U490 ( .A1(n818), .A2(data_in[7]), .B1(n1143), .B2(\mem[29][7] ), 
        .ZN(n1136) );
  INV_X1 U491 ( .A(n1133), .ZN(n270) );
  AOI22_X1 U492 ( .A1(data_in[0]), .A2(n817), .B1(n1132), .B2(\mem[30][0] ), 
        .ZN(n1133) );
  INV_X1 U493 ( .A(n1131), .ZN(n269) );
  AOI22_X1 U494 ( .A1(data_in[1]), .A2(n817), .B1(n1132), .B2(\mem[30][1] ), 
        .ZN(n1131) );
  INV_X1 U495 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U496 ( .A1(data_in[2]), .A2(n817), .B1(n1132), .B2(\mem[30][2] ), 
        .ZN(n1130) );
  INV_X1 U497 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U498 ( .A1(data_in[3]), .A2(n817), .B1(n1132), .B2(\mem[30][3] ), 
        .ZN(n1129) );
  INV_X1 U499 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U500 ( .A1(data_in[4]), .A2(n817), .B1(n1132), .B2(\mem[30][4] ), 
        .ZN(n1128) );
  INV_X1 U501 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U502 ( .A1(data_in[5]), .A2(n817), .B1(n1132), .B2(\mem[30][5] ), 
        .ZN(n1127) );
  INV_X1 U503 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U504 ( .A1(data_in[6]), .A2(n817), .B1(n1132), .B2(\mem[30][6] ), 
        .ZN(n1126) );
  INV_X1 U505 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U506 ( .A1(data_in[7]), .A2(n817), .B1(n1132), .B2(\mem[30][7] ), 
        .ZN(n1125) );
  INV_X1 U507 ( .A(n1123), .ZN(n262) );
  AOI22_X1 U508 ( .A1(data_in[0]), .A2(n816), .B1(n1122), .B2(\mem[31][0] ), 
        .ZN(n1123) );
  INV_X1 U509 ( .A(n1121), .ZN(n261) );
  AOI22_X1 U510 ( .A1(data_in[1]), .A2(n816), .B1(n1122), .B2(\mem[31][1] ), 
        .ZN(n1121) );
  INV_X1 U511 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U512 ( .A1(data_in[2]), .A2(n816), .B1(n1122), .B2(\mem[31][2] ), 
        .ZN(n1120) );
  INV_X1 U513 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U514 ( .A1(data_in[3]), .A2(n816), .B1(n1122), .B2(\mem[31][3] ), 
        .ZN(n1119) );
  INV_X1 U515 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U516 ( .A1(data_in[4]), .A2(n816), .B1(n1122), .B2(\mem[31][4] ), 
        .ZN(n1118) );
  INV_X1 U517 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U518 ( .A1(data_in[5]), .A2(n816), .B1(n1122), .B2(\mem[31][5] ), 
        .ZN(n1117) );
  INV_X1 U519 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U520 ( .A1(data_in[6]), .A2(n816), .B1(n1122), .B2(\mem[31][6] ), 
        .ZN(n1116) );
  INV_X1 U521 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U522 ( .A1(data_in[7]), .A2(n816), .B1(n1122), .B2(\mem[31][7] ), 
        .ZN(n1115) );
  INV_X1 U523 ( .A(n1113), .ZN(n810) );
  AOI22_X1 U524 ( .A1(data_in[0]), .A2(n842), .B1(n1112), .B2(\mem[0][0] ), 
        .ZN(n1113) );
  INV_X1 U525 ( .A(n1111), .ZN(n809) );
  AOI22_X1 U526 ( .A1(data_in[1]), .A2(n842), .B1(n1112), .B2(\mem[0][1] ), 
        .ZN(n1111) );
  INV_X1 U527 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U528 ( .A1(data_in[2]), .A2(n842), .B1(n1112), .B2(\mem[0][2] ), 
        .ZN(n1110) );
  INV_X1 U529 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U530 ( .A1(data_in[3]), .A2(n842), .B1(n1112), .B2(\mem[0][3] ), 
        .ZN(n1109) );
  INV_X1 U531 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U532 ( .A1(data_in[4]), .A2(n842), .B1(n1112), .B2(\mem[0][4] ), 
        .ZN(n1108) );
  INV_X1 U533 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U534 ( .A1(data_in[5]), .A2(n842), .B1(n1112), .B2(\mem[0][5] ), 
        .ZN(n1107) );
  INV_X1 U535 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U536 ( .A1(data_in[6]), .A2(n842), .B1(n1112), .B2(\mem[0][6] ), 
        .ZN(n1106) );
  INV_X1 U537 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U538 ( .A1(data_in[7]), .A2(n842), .B1(n1112), .B2(\mem[0][7] ), 
        .ZN(n1105) );
  INV_X1 U539 ( .A(n1102), .ZN(n802) );
  AOI22_X1 U540 ( .A1(data_in[0]), .A2(n841), .B1(n1101), .B2(\mem[1][0] ), 
        .ZN(n1102) );
  INV_X1 U541 ( .A(n1100), .ZN(n801) );
  AOI22_X1 U542 ( .A1(data_in[1]), .A2(n841), .B1(n1101), .B2(\mem[1][1] ), 
        .ZN(n1100) );
  INV_X1 U543 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U544 ( .A1(data_in[2]), .A2(n841), .B1(n1101), .B2(\mem[1][2] ), 
        .ZN(n1099) );
  INV_X1 U545 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U546 ( .A1(data_in[3]), .A2(n841), .B1(n1101), .B2(\mem[1][3] ), 
        .ZN(n1098) );
  INV_X1 U547 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U548 ( .A1(data_in[4]), .A2(n841), .B1(n1101), .B2(\mem[1][4] ), 
        .ZN(n1097) );
  INV_X1 U549 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U550 ( .A1(data_in[5]), .A2(n841), .B1(n1101), .B2(\mem[1][5] ), 
        .ZN(n1096) );
  INV_X1 U551 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U552 ( .A1(data_in[6]), .A2(n841), .B1(n1101), .B2(\mem[1][6] ), 
        .ZN(n1095) );
  INV_X1 U553 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U554 ( .A1(data_in[7]), .A2(n841), .B1(n1101), .B2(\mem[1][7] ), 
        .ZN(n1094) );
  INV_X1 U555 ( .A(n1092), .ZN(n794) );
  AOI22_X1 U556 ( .A1(data_in[0]), .A2(n840), .B1(n1091), .B2(\mem[2][0] ), 
        .ZN(n1092) );
  INV_X1 U557 ( .A(n1090), .ZN(n793) );
  AOI22_X1 U558 ( .A1(data_in[1]), .A2(n840), .B1(n1091), .B2(\mem[2][1] ), 
        .ZN(n1090) );
  INV_X1 U559 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U560 ( .A1(data_in[2]), .A2(n840), .B1(n1091), .B2(\mem[2][2] ), 
        .ZN(n1089) );
  INV_X1 U561 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U562 ( .A1(data_in[3]), .A2(n840), .B1(n1091), .B2(\mem[2][3] ), 
        .ZN(n1088) );
  INV_X1 U563 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U564 ( .A1(data_in[4]), .A2(n840), .B1(n1091), .B2(\mem[2][4] ), 
        .ZN(n1087) );
  INV_X1 U565 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U566 ( .A1(data_in[5]), .A2(n840), .B1(n1091), .B2(\mem[2][5] ), 
        .ZN(n1086) );
  INV_X1 U567 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U568 ( .A1(data_in[6]), .A2(n840), .B1(n1091), .B2(\mem[2][6] ), 
        .ZN(n1085) );
  INV_X1 U569 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U570 ( .A1(data_in[7]), .A2(n840), .B1(n1091), .B2(\mem[2][7] ), 
        .ZN(n1084) );
  INV_X1 U571 ( .A(n1082), .ZN(n786) );
  AOI22_X1 U572 ( .A1(data_in[0]), .A2(n839), .B1(n1081), .B2(\mem[3][0] ), 
        .ZN(n1082) );
  INV_X1 U573 ( .A(n1080), .ZN(n785) );
  AOI22_X1 U574 ( .A1(data_in[1]), .A2(n839), .B1(n1081), .B2(\mem[3][1] ), 
        .ZN(n1080) );
  INV_X1 U575 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U576 ( .A1(data_in[2]), .A2(n839), .B1(n1081), .B2(\mem[3][2] ), 
        .ZN(n1079) );
  INV_X1 U577 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U578 ( .A1(data_in[3]), .A2(n839), .B1(n1081), .B2(\mem[3][3] ), 
        .ZN(n1078) );
  INV_X1 U579 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U580 ( .A1(data_in[4]), .A2(n839), .B1(n1081), .B2(\mem[3][4] ), 
        .ZN(n1077) );
  INV_X1 U581 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U582 ( .A1(data_in[5]), .A2(n839), .B1(n1081), .B2(\mem[3][5] ), 
        .ZN(n1076) );
  INV_X1 U583 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U584 ( .A1(data_in[6]), .A2(n839), .B1(n1081), .B2(\mem[3][6] ), 
        .ZN(n1075) );
  INV_X1 U585 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U586 ( .A1(data_in[7]), .A2(n839), .B1(n1081), .B2(\mem[3][7] ), 
        .ZN(n1074) );
  INV_X1 U587 ( .A(n1072), .ZN(n778) );
  AOI22_X1 U588 ( .A1(data_in[0]), .A2(n838), .B1(n1071), .B2(\mem[4][0] ), 
        .ZN(n1072) );
  INV_X1 U589 ( .A(n1070), .ZN(n777) );
  AOI22_X1 U590 ( .A1(data_in[1]), .A2(n838), .B1(n1071), .B2(\mem[4][1] ), 
        .ZN(n1070) );
  INV_X1 U591 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U592 ( .A1(data_in[2]), .A2(n838), .B1(n1071), .B2(\mem[4][2] ), 
        .ZN(n1069) );
  INV_X1 U593 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U594 ( .A1(data_in[3]), .A2(n838), .B1(n1071), .B2(\mem[4][3] ), 
        .ZN(n1068) );
  INV_X1 U595 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U596 ( .A1(data_in[4]), .A2(n838), .B1(n1071), .B2(\mem[4][4] ), 
        .ZN(n1067) );
  INV_X1 U597 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U598 ( .A1(data_in[5]), .A2(n838), .B1(n1071), .B2(\mem[4][5] ), 
        .ZN(n1066) );
  INV_X1 U599 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U600 ( .A1(data_in[6]), .A2(n838), .B1(n1071), .B2(\mem[4][6] ), 
        .ZN(n1065) );
  INV_X1 U601 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U602 ( .A1(data_in[7]), .A2(n838), .B1(n1071), .B2(\mem[4][7] ), 
        .ZN(n1064) );
  INV_X1 U603 ( .A(N13), .ZN(n843) );
  INV_X1 U604 ( .A(N14), .ZN(n844) );
  MUX2_X1 U605 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n246), .Z(n2) );
  MUX2_X1 U606 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n246), .Z(n3) );
  MUX2_X1 U607 ( .A(n3), .B(n2), .S(n243), .Z(n4) );
  MUX2_X1 U608 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n246), .Z(n5) );
  MUX2_X1 U609 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n246), .Z(n6) );
  MUX2_X1 U610 ( .A(n6), .B(n5), .S(n243), .Z(n7) );
  MUX2_X1 U611 ( .A(n7), .B(n4), .S(n242), .Z(n8) );
  MUX2_X1 U612 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n246), .Z(n9) );
  MUX2_X1 U613 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n246), .Z(n10) );
  MUX2_X1 U614 ( .A(n10), .B(n9), .S(N11), .Z(n11) );
  MUX2_X1 U615 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n246), .Z(n12) );
  MUX2_X1 U616 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n246), .Z(n13) );
  MUX2_X1 U617 ( .A(n13), .B(n12), .S(n245), .Z(n14) );
  MUX2_X1 U618 ( .A(n14), .B(n11), .S(N12), .Z(n15) );
  MUX2_X1 U619 ( .A(n15), .B(n8), .S(N13), .Z(n16) );
  MUX2_X1 U620 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n247), .Z(n17) );
  MUX2_X1 U621 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n247), .Z(n18) );
  MUX2_X1 U622 ( .A(n18), .B(n17), .S(n243), .Z(n19) );
  MUX2_X1 U623 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n247), .Z(n20) );
  MUX2_X1 U624 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n247), .Z(n21) );
  MUX2_X1 U625 ( .A(n21), .B(n20), .S(n243), .Z(n22) );
  MUX2_X1 U626 ( .A(n22), .B(n19), .S(N12), .Z(n23) );
  MUX2_X1 U627 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n247), .Z(n24) );
  MUX2_X1 U628 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n247), .Z(n25) );
  MUX2_X1 U629 ( .A(n25), .B(n24), .S(n243), .Z(n26) );
  MUX2_X1 U630 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n247), .Z(n27) );
  MUX2_X1 U631 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n247), .Z(n28) );
  MUX2_X1 U632 ( .A(n28), .B(n27), .S(n243), .Z(n29) );
  MUX2_X1 U633 ( .A(n29), .B(n26), .S(N12), .Z(n30) );
  MUX2_X1 U634 ( .A(n30), .B(n23), .S(N13), .Z(n31) );
  MUX2_X1 U635 ( .A(n31), .B(n16), .S(N14), .Z(N22) );
  MUX2_X1 U636 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n247), .Z(n32) );
  MUX2_X1 U637 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n247), .Z(n33) );
  MUX2_X1 U638 ( .A(n33), .B(n32), .S(n243), .Z(n34) );
  MUX2_X1 U639 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n247), .Z(n35) );
  MUX2_X1 U640 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n247), .Z(n36) );
  MUX2_X1 U641 ( .A(n36), .B(n35), .S(n243), .Z(n37) );
  MUX2_X1 U642 ( .A(n37), .B(n34), .S(n242), .Z(n38) );
  MUX2_X1 U643 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n248), .Z(n39) );
  MUX2_X1 U644 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n248), .Z(n40) );
  MUX2_X1 U645 ( .A(n40), .B(n39), .S(n243), .Z(n41) );
  MUX2_X1 U646 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n248), .Z(n42) );
  MUX2_X1 U647 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n248), .Z(n43) );
  MUX2_X1 U648 ( .A(n43), .B(n42), .S(n243), .Z(n44) );
  MUX2_X1 U649 ( .A(n44), .B(n41), .S(n242), .Z(n45) );
  MUX2_X1 U650 ( .A(n45), .B(n38), .S(N13), .Z(n46) );
  MUX2_X1 U651 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n248), .Z(n47) );
  MUX2_X1 U652 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n248), .Z(n48) );
  MUX2_X1 U653 ( .A(n48), .B(n47), .S(n243), .Z(n49) );
  MUX2_X1 U654 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n248), .Z(n50) );
  MUX2_X1 U655 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n248), .Z(n51) );
  MUX2_X1 U656 ( .A(n51), .B(n50), .S(n243), .Z(n52) );
  MUX2_X1 U657 ( .A(n52), .B(n49), .S(n242), .Z(n53) );
  MUX2_X1 U658 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n248), .Z(n54) );
  MUX2_X1 U659 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n248), .Z(n55) );
  MUX2_X1 U660 ( .A(n55), .B(n54), .S(n243), .Z(n56) );
  MUX2_X1 U661 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n248), .Z(n57) );
  MUX2_X1 U662 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n248), .Z(n58) );
  MUX2_X1 U663 ( .A(n58), .B(n57), .S(n243), .Z(n59) );
  MUX2_X1 U664 ( .A(n59), .B(n56), .S(n242), .Z(n60) );
  MUX2_X1 U665 ( .A(n60), .B(n53), .S(N13), .Z(n61) );
  MUX2_X1 U666 ( .A(n61), .B(n46), .S(N14), .Z(N21) );
  MUX2_X1 U667 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n249), .Z(n62) );
  MUX2_X1 U668 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n249), .Z(n63) );
  MUX2_X1 U669 ( .A(n63), .B(n62), .S(n244), .Z(n64) );
  MUX2_X1 U670 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n249), .Z(n65) );
  MUX2_X1 U671 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n249), .Z(n66) );
  MUX2_X1 U672 ( .A(n66), .B(n65), .S(n244), .Z(n67) );
  MUX2_X1 U673 ( .A(n67), .B(n64), .S(n242), .Z(n68) );
  MUX2_X1 U674 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n249), .Z(n69) );
  MUX2_X1 U675 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n249), .Z(n70) );
  MUX2_X1 U676 ( .A(n70), .B(n69), .S(n244), .Z(n71) );
  MUX2_X1 U677 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n249), .Z(n72) );
  MUX2_X1 U678 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n249), .Z(n73) );
  MUX2_X1 U679 ( .A(n73), .B(n72), .S(n244), .Z(n74) );
  MUX2_X1 U680 ( .A(n74), .B(n71), .S(n242), .Z(n75) );
  MUX2_X1 U681 ( .A(n75), .B(n68), .S(N13), .Z(n76) );
  MUX2_X1 U682 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n249), .Z(n77) );
  MUX2_X1 U683 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n249), .Z(n78) );
  MUX2_X1 U684 ( .A(n78), .B(n77), .S(n244), .Z(n79) );
  MUX2_X1 U685 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n249), .Z(n80) );
  MUX2_X1 U686 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n249), .Z(n81) );
  MUX2_X1 U687 ( .A(n81), .B(n80), .S(n244), .Z(n82) );
  MUX2_X1 U688 ( .A(n82), .B(n79), .S(n242), .Z(n83) );
  MUX2_X1 U689 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n250), .Z(n84) );
  MUX2_X1 U690 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n250), .Z(n85) );
  MUX2_X1 U691 ( .A(n85), .B(n84), .S(n244), .Z(n86) );
  MUX2_X1 U692 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n250), .Z(n87) );
  MUX2_X1 U693 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n250), .Z(n88) );
  MUX2_X1 U694 ( .A(n88), .B(n87), .S(n244), .Z(n89) );
  MUX2_X1 U695 ( .A(n89), .B(n86), .S(n242), .Z(n90) );
  MUX2_X1 U696 ( .A(n90), .B(n83), .S(N13), .Z(n91) );
  MUX2_X1 U697 ( .A(n91), .B(n76), .S(N14), .Z(N20) );
  MUX2_X1 U698 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n250), .Z(n92) );
  MUX2_X1 U699 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n93) );
  MUX2_X1 U700 ( .A(n93), .B(n92), .S(n244), .Z(n94) );
  MUX2_X1 U701 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n250), .Z(n95) );
  MUX2_X1 U702 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n250), .Z(n96) );
  MUX2_X1 U703 ( .A(n96), .B(n95), .S(n244), .Z(n97) );
  MUX2_X1 U704 ( .A(n97), .B(n94), .S(n242), .Z(n98) );
  MUX2_X1 U705 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n99) );
  MUX2_X1 U706 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n250), .Z(n100) );
  MUX2_X1 U707 ( .A(n100), .B(n99), .S(n244), .Z(n101) );
  MUX2_X1 U708 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n250), .Z(n102) );
  MUX2_X1 U709 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n250), .Z(n103) );
  MUX2_X1 U710 ( .A(n103), .B(n102), .S(n244), .Z(n104) );
  MUX2_X1 U711 ( .A(n104), .B(n101), .S(n242), .Z(n105) );
  MUX2_X1 U712 ( .A(n105), .B(n98), .S(N13), .Z(n106) );
  MUX2_X1 U713 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n248), .Z(n107) );
  MUX2_X1 U714 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(N10), .Z(n108) );
  MUX2_X1 U715 ( .A(n108), .B(n107), .S(n245), .Z(n109) );
  MUX2_X1 U716 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n247), .Z(n110) );
  MUX2_X1 U717 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n251), .Z(n111) );
  MUX2_X1 U718 ( .A(n111), .B(n110), .S(n245), .Z(n112) );
  MUX2_X1 U719 ( .A(n112), .B(n109), .S(n242), .Z(n113) );
  MUX2_X1 U720 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(N10), .Z(n114) );
  MUX2_X1 U721 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n249), .Z(n115) );
  MUX2_X1 U722 ( .A(n115), .B(n114), .S(n245), .Z(n116) );
  MUX2_X1 U723 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n117) );
  MUX2_X1 U724 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n250), .Z(n118) );
  MUX2_X1 U725 ( .A(n118), .B(n117), .S(n245), .Z(n119) );
  MUX2_X1 U726 ( .A(n119), .B(n116), .S(n242), .Z(n120) );
  MUX2_X1 U727 ( .A(n120), .B(n113), .S(N13), .Z(n121) );
  MUX2_X1 U728 ( .A(n121), .B(n106), .S(N14), .Z(N19) );
  MUX2_X1 U729 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n251), .Z(n122) );
  MUX2_X1 U730 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n251), .Z(n123) );
  MUX2_X1 U731 ( .A(n123), .B(n122), .S(n245), .Z(n124) );
  MUX2_X1 U732 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n248), .Z(n125) );
  MUX2_X1 U733 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n251), .Z(n126) );
  MUX2_X1 U734 ( .A(n126), .B(n125), .S(n245), .Z(n127) );
  MUX2_X1 U735 ( .A(n127), .B(n124), .S(n242), .Z(n128) );
  MUX2_X1 U736 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n247), .Z(n129) );
  MUX2_X1 U737 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n251), .Z(n130) );
  MUX2_X1 U738 ( .A(n130), .B(n129), .S(n245), .Z(n131) );
  MUX2_X1 U739 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n250), .Z(n132) );
  MUX2_X1 U740 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(N10), .Z(n133) );
  MUX2_X1 U741 ( .A(n133), .B(n132), .S(n245), .Z(n134) );
  MUX2_X1 U742 ( .A(n134), .B(n131), .S(n242), .Z(n135) );
  MUX2_X1 U743 ( .A(n135), .B(n128), .S(N13), .Z(n136) );
  MUX2_X1 U744 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n246), .Z(n137) );
  MUX2_X1 U745 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n248), .Z(n138) );
  MUX2_X1 U746 ( .A(n138), .B(n137), .S(n245), .Z(n139) );
  MUX2_X1 U747 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n248), .Z(n140) );
  MUX2_X1 U748 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(N10), .Z(n141) );
  MUX2_X1 U749 ( .A(n141), .B(n140), .S(n245), .Z(n142) );
  MUX2_X1 U750 ( .A(n142), .B(n139), .S(n242), .Z(n143) );
  MUX2_X1 U751 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n249), .Z(n144) );
  MUX2_X1 U752 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(N10), .Z(n145) );
  MUX2_X1 U753 ( .A(n145), .B(n144), .S(n245), .Z(n146) );
  MUX2_X1 U754 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(N10), .Z(n147) );
  MUX2_X1 U755 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n148) );
  MUX2_X1 U756 ( .A(n148), .B(n147), .S(n245), .Z(n149) );
  MUX2_X1 U757 ( .A(n149), .B(n146), .S(n242), .Z(n150) );
  MUX2_X1 U758 ( .A(n150), .B(n143), .S(N13), .Z(n151) );
  MUX2_X1 U759 ( .A(n151), .B(n136), .S(N14), .Z(N18) );
  MUX2_X1 U760 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n246), .Z(n152) );
  MUX2_X1 U761 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n246), .Z(n153) );
  MUX2_X1 U762 ( .A(n153), .B(n152), .S(n243), .Z(n154) );
  MUX2_X1 U763 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n246), .Z(n155) );
  MUX2_X1 U764 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(N10), .Z(n156) );
  MUX2_X1 U765 ( .A(n156), .B(n155), .S(N11), .Z(n157) );
  MUX2_X1 U766 ( .A(n157), .B(n154), .S(n242), .Z(n158) );
  MUX2_X1 U767 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(N10), .Z(n159) );
  MUX2_X1 U768 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(N10), .Z(n160) );
  MUX2_X1 U769 ( .A(n160), .B(n159), .S(N11), .Z(n161) );
  MUX2_X1 U770 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n247), .Z(n162) );
  MUX2_X1 U771 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(N10), .Z(n163) );
  MUX2_X1 U772 ( .A(n163), .B(n162), .S(n243), .Z(n164) );
  MUX2_X1 U773 ( .A(n164), .B(n161), .S(N12), .Z(n165) );
  MUX2_X1 U774 ( .A(n165), .B(n158), .S(N13), .Z(n166) );
  MUX2_X1 U775 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n246), .Z(n167) );
  MUX2_X1 U776 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(N10), .Z(n168) );
  MUX2_X1 U777 ( .A(n168), .B(n167), .S(N11), .Z(n169) );
  MUX2_X1 U778 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n251), .Z(n170) );
  MUX2_X1 U779 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(N10), .Z(n171) );
  MUX2_X1 U780 ( .A(n171), .B(n170), .S(n244), .Z(n172) );
  MUX2_X1 U781 ( .A(n172), .B(n169), .S(n242), .Z(n173) );
  MUX2_X1 U782 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n250), .Z(n174) );
  MUX2_X1 U783 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n251), .Z(n175) );
  MUX2_X1 U784 ( .A(n175), .B(n174), .S(N11), .Z(n176) );
  MUX2_X1 U785 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n251), .Z(n177) );
  MUX2_X1 U786 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n251), .Z(n178) );
  MUX2_X1 U787 ( .A(n178), .B(n177), .S(n244), .Z(n179) );
  MUX2_X1 U788 ( .A(n179), .B(n176), .S(N12), .Z(n180) );
  MUX2_X1 U789 ( .A(n180), .B(n173), .S(N13), .Z(n181) );
  MUX2_X1 U790 ( .A(n181), .B(n166), .S(N14), .Z(N17) );
  MUX2_X1 U791 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n251), .Z(n182) );
  MUX2_X1 U792 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n246), .Z(n183) );
  MUX2_X1 U793 ( .A(n183), .B(n182), .S(N11), .Z(n184) );
  MUX2_X1 U794 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n250), .Z(n185) );
  MUX2_X1 U795 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n251), .Z(n186) );
  MUX2_X1 U796 ( .A(n186), .B(n185), .S(N11), .Z(n187) );
  MUX2_X1 U797 ( .A(n187), .B(n184), .S(n242), .Z(n188) );
  MUX2_X1 U798 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n249), .Z(n189) );
  MUX2_X1 U799 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n251), .Z(n190) );
  MUX2_X1 U800 ( .A(n190), .B(n189), .S(N11), .Z(n191) );
  MUX2_X1 U801 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n250), .Z(n192) );
  MUX2_X1 U802 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n251), .Z(n193) );
  MUX2_X1 U803 ( .A(n193), .B(n192), .S(n245), .Z(n194) );
  MUX2_X1 U804 ( .A(n194), .B(n191), .S(N12), .Z(n195) );
  MUX2_X1 U805 ( .A(n195), .B(n188), .S(N13), .Z(n196) );
  MUX2_X1 U806 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n246), .Z(n197) );
  MUX2_X1 U807 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n251), .Z(n198) );
  MUX2_X1 U808 ( .A(n198), .B(n197), .S(n243), .Z(n199) );
  MUX2_X1 U809 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n247), .Z(n200) );
  MUX2_X1 U810 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n249), .Z(n201) );
  MUX2_X1 U811 ( .A(n201), .B(n200), .S(n245), .Z(n202) );
  MUX2_X1 U812 ( .A(n202), .B(n199), .S(n242), .Z(n203) );
  MUX2_X1 U813 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n249), .Z(n204) );
  MUX2_X1 U814 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n251), .Z(n205) );
  MUX2_X1 U815 ( .A(n205), .B(n204), .S(n245), .Z(n206) );
  MUX2_X1 U816 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n251), .Z(n207) );
  MUX2_X1 U817 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n248), .Z(n208) );
  MUX2_X1 U818 ( .A(n208), .B(n207), .S(N11), .Z(n209) );
  MUX2_X1 U819 ( .A(n209), .B(n206), .S(N12), .Z(n210) );
  MUX2_X1 U820 ( .A(n210), .B(n203), .S(N13), .Z(n211) );
  MUX2_X1 U821 ( .A(n211), .B(n196), .S(N14), .Z(N16) );
  MUX2_X1 U822 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(N10), .Z(n212) );
  MUX2_X1 U823 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n249), .Z(n213) );
  MUX2_X1 U824 ( .A(n213), .B(n212), .S(n244), .Z(n214) );
  MUX2_X1 U825 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n248), .Z(n215) );
  MUX2_X1 U826 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n246), .Z(n216) );
  MUX2_X1 U827 ( .A(n216), .B(n215), .S(n245), .Z(n217) );
  MUX2_X1 U828 ( .A(n217), .B(n214), .S(n242), .Z(n218) );
  MUX2_X1 U829 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n247), .Z(n219) );
  MUX2_X1 U830 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n251), .Z(n220) );
  MUX2_X1 U831 ( .A(n220), .B(n219), .S(n244), .Z(n221) );
  MUX2_X1 U832 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n247), .Z(n222) );
  MUX2_X1 U833 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n251), .Z(n223) );
  MUX2_X1 U834 ( .A(n223), .B(n222), .S(N11), .Z(n224) );
  MUX2_X1 U835 ( .A(n224), .B(n221), .S(N12), .Z(n225) );
  MUX2_X1 U836 ( .A(n225), .B(n218), .S(N13), .Z(n226) );
  MUX2_X1 U837 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n251), .Z(n227) );
  MUX2_X1 U838 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n250), .Z(n228) );
  MUX2_X1 U839 ( .A(n228), .B(n227), .S(N11), .Z(n229) );
  MUX2_X1 U840 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n248), .Z(n230) );
  MUX2_X1 U841 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n251), .Z(n231) );
  MUX2_X1 U842 ( .A(n231), .B(n230), .S(N11), .Z(n232) );
  MUX2_X1 U843 ( .A(n232), .B(n229), .S(n242), .Z(n233) );
  MUX2_X1 U844 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n249), .Z(n234) );
  MUX2_X1 U845 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n247), .Z(n235) );
  MUX2_X1 U846 ( .A(n235), .B(n234), .S(n244), .Z(n236) );
  MUX2_X1 U847 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n250), .Z(n237) );
  MUX2_X1 U848 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n246), .Z(n238) );
  MUX2_X1 U849 ( .A(n238), .B(n237), .S(N11), .Z(n239) );
  MUX2_X1 U850 ( .A(n239), .B(n236), .S(N12), .Z(n240) );
  MUX2_X1 U851 ( .A(n240), .B(n233), .S(N13), .Z(n241) );
  MUX2_X1 U852 ( .A(n241), .B(n226), .S(N14), .Z(N15) );
  CLKBUF_X1 U853 ( .A(n251), .Z(n246) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_14 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n255), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n256), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n257), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n258), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n259), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n260), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n261), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n262), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n263), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n264), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n265), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n266), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n267), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n268), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n269), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n270), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n271), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n272), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n273), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n274), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n275), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n276), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n277), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n278), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n279), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n280), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n281), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n282), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n283), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n284), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n285), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n286), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n287), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n288), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n289), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n290), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n291), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n292), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n293), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n594), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n595), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n596), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n597), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n598), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n599), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n600), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n601), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n602), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n603), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n604), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n605), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n606), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n607), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n608), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n609), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n610), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n611), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n612), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n613), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n614), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n615), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n616), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n617), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n618), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n619), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n620), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n621), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n622), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n623), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n624), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n625), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n626), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n627), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n628), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n629), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n630), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n631), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n632), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n633), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n634), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n635), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n636), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n637), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n638), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n639), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n640), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n641), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n642), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n643), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n644), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n645), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n646), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n647), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n648), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n649), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n650), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n651), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n652), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n653), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n654), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n655), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n656), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n657), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n658), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n659), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n660), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n661), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n662), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n663), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n664), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n665), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n666), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n667), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n668), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n669), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n670), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n671), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n672), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n673), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n674), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n675), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n676), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n677), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n678), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n679), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n680), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n681), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n682), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n683), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n684), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n685), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n686), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n687), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n688), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n689), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n690), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n691), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n692), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n693), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n694), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n695), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n696), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n697), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n698), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n699), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n700), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n701), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n702), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n703), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n704), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n705), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n706), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n707), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n708), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n709), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n710), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n711), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n712), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n713), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n714), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n715), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n716), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n717), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n718), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n719), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n720), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n721), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n722), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n723), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n724), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n725), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n726), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n727), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n728), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n729), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n730), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n731), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n732), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n733), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n734), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n735), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n736), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n737), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n738), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n739), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n740), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n741), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n742), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n743), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n744), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n745), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n746), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n747), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n748), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n749), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n750), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n751), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n752), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n753), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n754), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n755), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n756), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n757), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n758), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n759), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n760), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n761), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n762), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n763), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n764), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n765), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n766), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n767), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n768), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n769), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n770), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n771), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n772), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n773), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n774), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n775), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n776), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n777), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n778), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n779), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n780), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n781), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n782), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n783), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n784), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n785), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n786), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n787), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n788), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n789), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n790), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n791), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n792), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n793), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n794), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n795), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n796), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n797), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n798), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n799), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n800), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n801), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n802), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n803), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n804), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n805), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n806), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n807), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n808), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n809), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n810), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  BUF_X1 U3 ( .A(N10), .Z(n248) );
  BUF_X1 U4 ( .A(n251), .Z(n249) );
  BUF_X1 U5 ( .A(n251), .Z(n250) );
  BUF_X1 U6 ( .A(n251), .Z(n247) );
  BUF_X1 U7 ( .A(n251), .Z(n246) );
  BUF_X1 U8 ( .A(N10), .Z(n251) );
  INV_X1 U9 ( .A(n1112), .ZN(n842) );
  INV_X1 U10 ( .A(n1101), .ZN(n841) );
  INV_X1 U11 ( .A(n1091), .ZN(n840) );
  INV_X1 U12 ( .A(n1081), .ZN(n839) );
  INV_X1 U13 ( .A(n1071), .ZN(n838) );
  INV_X1 U14 ( .A(n1061), .ZN(n837) );
  INV_X1 U15 ( .A(n1052), .ZN(n836) );
  INV_X1 U16 ( .A(n1043), .ZN(n835) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1104) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n252), .ZN(n1093) );
  NAND2_X1 U19 ( .A1(n1103), .A2(n1135), .ZN(n1061) );
  NAND2_X1 U20 ( .A1(n1104), .A2(n1103), .ZN(n1112) );
  NAND2_X1 U21 ( .A1(n1093), .A2(n1103), .ZN(n1101) );
  NAND2_X1 U22 ( .A1(n1083), .A2(n1103), .ZN(n1091) );
  NAND2_X1 U23 ( .A1(n1073), .A2(n1103), .ZN(n1081) );
  NAND2_X1 U24 ( .A1(n1063), .A2(n1103), .ZN(n1071) );
  NAND2_X1 U25 ( .A1(n1103), .A2(n1124), .ZN(n1052) );
  NAND2_X1 U26 ( .A1(n1103), .A2(n1114), .ZN(n1043) );
  INV_X1 U27 ( .A(n1132), .ZN(n817) );
  INV_X1 U28 ( .A(n1122), .ZN(n816) );
  INV_X1 U29 ( .A(n888), .ZN(n815) );
  INV_X1 U30 ( .A(n879), .ZN(n814) );
  INV_X1 U31 ( .A(n870), .ZN(n813) );
  INV_X1 U32 ( .A(n861), .ZN(n812) );
  INV_X1 U33 ( .A(n852), .ZN(n811) );
  INV_X1 U34 ( .A(n988), .ZN(n829) );
  INV_X1 U35 ( .A(n979), .ZN(n828) );
  INV_X1 U36 ( .A(n970), .ZN(n827) );
  INV_X1 U37 ( .A(n915), .ZN(n821) );
  INV_X1 U38 ( .A(n906), .ZN(n820) );
  INV_X1 U39 ( .A(n897), .ZN(n819) );
  INV_X1 U40 ( .A(n1034), .ZN(n834) );
  INV_X1 U41 ( .A(n1024), .ZN(n833) );
  INV_X1 U42 ( .A(n1015), .ZN(n832) );
  INV_X1 U43 ( .A(n1006), .ZN(n831) );
  INV_X1 U44 ( .A(n997), .ZN(n830) );
  INV_X1 U45 ( .A(n961), .ZN(n826) );
  INV_X1 U46 ( .A(n951), .ZN(n825) );
  INV_X1 U47 ( .A(n942), .ZN(n824) );
  INV_X1 U48 ( .A(n933), .ZN(n823) );
  INV_X1 U49 ( .A(n924), .ZN(n822) );
  INV_X1 U50 ( .A(n1143), .ZN(n818) );
  BUF_X1 U51 ( .A(N11), .Z(n244) );
  BUF_X1 U52 ( .A(N11), .Z(n245) );
  INV_X1 U53 ( .A(N10), .ZN(n252) );
  BUF_X1 U54 ( .A(N12), .Z(n242) );
  NOR3_X1 U55 ( .A1(n254), .A2(N10), .A3(n253), .ZN(n1124) );
  NOR3_X1 U56 ( .A1(n254), .A2(n252), .A3(n253), .ZN(n1114) );
  NOR3_X1 U57 ( .A1(n252), .A2(N11), .A3(n254), .ZN(n1135) );
  NOR3_X1 U58 ( .A1(N10), .A2(N12), .A3(n253), .ZN(n1083) );
  NOR3_X1 U59 ( .A1(n252), .A2(N12), .A3(n253), .ZN(n1073) );
  NOR3_X1 U60 ( .A1(N10), .A2(N11), .A3(n254), .ZN(n1063) );
  NAND2_X1 U61 ( .A1(n1026), .A2(n1135), .ZN(n988) );
  NAND2_X1 U62 ( .A1(n953), .A2(n1135), .ZN(n915) );
  NAND2_X1 U63 ( .A1(n1026), .A2(n1063), .ZN(n997) );
  NAND2_X1 U64 ( .A1(n953), .A2(n1063), .ZN(n924) );
  NAND2_X1 U65 ( .A1(n1026), .A2(n1104), .ZN(n1034) );
  NAND2_X1 U66 ( .A1(n1026), .A2(n1093), .ZN(n1024) );
  NAND2_X1 U67 ( .A1(n953), .A2(n1104), .ZN(n961) );
  NAND2_X1 U68 ( .A1(n953), .A2(n1093), .ZN(n951) );
  NAND2_X1 U69 ( .A1(n1104), .A2(n1134), .ZN(n888) );
  NAND2_X1 U70 ( .A1(n1093), .A2(n1134), .ZN(n879) );
  NAND2_X1 U71 ( .A1(n1083), .A2(n1134), .ZN(n870) );
  NAND2_X1 U72 ( .A1(n1073), .A2(n1134), .ZN(n861) );
  NAND2_X1 U73 ( .A1(n1063), .A2(n1134), .ZN(n852) );
  NAND2_X1 U74 ( .A1(n1135), .A2(n1134), .ZN(n1143) );
  NAND2_X1 U75 ( .A1(n1124), .A2(n1134), .ZN(n1132) );
  NAND2_X1 U76 ( .A1(n1114), .A2(n1134), .ZN(n1122) );
  NAND2_X1 U77 ( .A1(n1026), .A2(n1083), .ZN(n1015) );
  NAND2_X1 U78 ( .A1(n1026), .A2(n1073), .ZN(n1006) );
  NAND2_X1 U79 ( .A1(n953), .A2(n1083), .ZN(n942) );
  NAND2_X1 U80 ( .A1(n953), .A2(n1073), .ZN(n933) );
  NAND2_X1 U81 ( .A1(n1026), .A2(n1124), .ZN(n979) );
  NAND2_X1 U82 ( .A1(n953), .A2(n1124), .ZN(n906) );
  NAND2_X1 U83 ( .A1(n1026), .A2(n1114), .ZN(n970) );
  NAND2_X1 U84 ( .A1(n953), .A2(n1114), .ZN(n897) );
  AND3_X1 U85 ( .A1(n843), .A2(n844), .A3(wr_en), .ZN(n1103) );
  AND3_X1 U86 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1134) );
  AND3_X1 U87 ( .A1(N13), .A2(n844), .A3(wr_en), .ZN(n1026) );
  AND3_X1 U88 ( .A1(N14), .A2(n843), .A3(wr_en), .ZN(n953) );
  INV_X1 U89 ( .A(n1062), .ZN(n770) );
  AOI22_X1 U90 ( .A1(data_in[0]), .A2(n837), .B1(n1061), .B2(\mem[5][0] ), 
        .ZN(n1062) );
  INV_X1 U91 ( .A(n1060), .ZN(n769) );
  AOI22_X1 U92 ( .A1(data_in[1]), .A2(n837), .B1(n1061), .B2(\mem[5][1] ), 
        .ZN(n1060) );
  INV_X1 U93 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U94 ( .A1(data_in[2]), .A2(n837), .B1(n1061), .B2(\mem[5][2] ), 
        .ZN(n1059) );
  INV_X1 U95 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U96 ( .A1(data_in[3]), .A2(n837), .B1(n1061), .B2(\mem[5][3] ), 
        .ZN(n1058) );
  INV_X1 U97 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U98 ( .A1(data_in[4]), .A2(n837), .B1(n1061), .B2(\mem[5][4] ), 
        .ZN(n1057) );
  INV_X1 U99 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U100 ( .A1(data_in[5]), .A2(n837), .B1(n1061), .B2(\mem[5][5] ), 
        .ZN(n1056) );
  INV_X1 U101 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U102 ( .A1(data_in[6]), .A2(n837), .B1(n1061), .B2(\mem[5][6] ), 
        .ZN(n1055) );
  INV_X1 U103 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U104 ( .A1(data_in[7]), .A2(n837), .B1(n1061), .B2(\mem[5][7] ), 
        .ZN(n1054) );
  INV_X1 U105 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U106 ( .A1(data_in[5]), .A2(n833), .B1(n1024), .B2(\mem[9][5] ), 
        .ZN(n1019) );
  INV_X1 U107 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U108 ( .A1(data_in[6]), .A2(n833), .B1(n1024), .B2(\mem[9][6] ), 
        .ZN(n1018) );
  INV_X1 U109 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U110 ( .A1(data_in[7]), .A2(n833), .B1(n1024), .B2(\mem[9][7] ), 
        .ZN(n1017) );
  INV_X1 U111 ( .A(n989), .ZN(n706) );
  AOI22_X1 U112 ( .A1(data_in[0]), .A2(n829), .B1(n988), .B2(\mem[13][0] ), 
        .ZN(n989) );
  INV_X1 U113 ( .A(n987), .ZN(n705) );
  AOI22_X1 U114 ( .A1(data_in[1]), .A2(n829), .B1(n988), .B2(\mem[13][1] ), 
        .ZN(n987) );
  INV_X1 U115 ( .A(n986), .ZN(n704) );
  AOI22_X1 U116 ( .A1(data_in[2]), .A2(n829), .B1(n988), .B2(\mem[13][2] ), 
        .ZN(n986) );
  INV_X1 U117 ( .A(n985), .ZN(n703) );
  AOI22_X1 U118 ( .A1(data_in[3]), .A2(n829), .B1(n988), .B2(\mem[13][3] ), 
        .ZN(n985) );
  INV_X1 U119 ( .A(n984), .ZN(n702) );
  AOI22_X1 U120 ( .A1(data_in[4]), .A2(n829), .B1(n988), .B2(\mem[13][4] ), 
        .ZN(n984) );
  INV_X1 U121 ( .A(n983), .ZN(n701) );
  AOI22_X1 U122 ( .A1(data_in[5]), .A2(n829), .B1(n988), .B2(\mem[13][5] ), 
        .ZN(n983) );
  INV_X1 U123 ( .A(n982), .ZN(n700) );
  AOI22_X1 U124 ( .A1(data_in[6]), .A2(n829), .B1(n988), .B2(\mem[13][6] ), 
        .ZN(n982) );
  INV_X1 U125 ( .A(n981), .ZN(n699) );
  AOI22_X1 U126 ( .A1(data_in[7]), .A2(n829), .B1(n988), .B2(\mem[13][7] ), 
        .ZN(n981) );
  INV_X1 U127 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U128 ( .A1(data_in[0]), .A2(n832), .B1(n1015), .B2(\mem[10][0] ), 
        .ZN(n1016) );
  INV_X1 U129 ( .A(n1014), .ZN(n729) );
  AOI22_X1 U130 ( .A1(data_in[1]), .A2(n832), .B1(n1015), .B2(\mem[10][1] ), 
        .ZN(n1014) );
  INV_X1 U131 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U132 ( .A1(data_in[2]), .A2(n832), .B1(n1015), .B2(\mem[10][2] ), 
        .ZN(n1013) );
  INV_X1 U133 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U134 ( .A1(data_in[3]), .A2(n832), .B1(n1015), .B2(\mem[10][3] ), 
        .ZN(n1012) );
  INV_X1 U135 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U136 ( .A1(data_in[4]), .A2(n832), .B1(n1015), .B2(\mem[10][4] ), 
        .ZN(n1011) );
  INV_X1 U137 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U138 ( .A1(data_in[5]), .A2(n832), .B1(n1015), .B2(\mem[10][5] ), 
        .ZN(n1010) );
  INV_X1 U139 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U140 ( .A1(data_in[6]), .A2(n832), .B1(n1015), .B2(\mem[10][6] ), 
        .ZN(n1009) );
  INV_X1 U141 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U142 ( .A1(data_in[7]), .A2(n832), .B1(n1015), .B2(\mem[10][7] ), 
        .ZN(n1008) );
  INV_X1 U143 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U144 ( .A1(data_in[0]), .A2(n831), .B1(n1006), .B2(\mem[11][0] ), 
        .ZN(n1007) );
  INV_X1 U145 ( .A(n1005), .ZN(n721) );
  AOI22_X1 U146 ( .A1(data_in[1]), .A2(n831), .B1(n1006), .B2(\mem[11][1] ), 
        .ZN(n1005) );
  INV_X1 U147 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U148 ( .A1(data_in[2]), .A2(n831), .B1(n1006), .B2(\mem[11][2] ), 
        .ZN(n1004) );
  INV_X1 U149 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U150 ( .A1(data_in[3]), .A2(n831), .B1(n1006), .B2(\mem[11][3] ), 
        .ZN(n1003) );
  INV_X1 U151 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U152 ( .A1(data_in[4]), .A2(n831), .B1(n1006), .B2(\mem[11][4] ), 
        .ZN(n1002) );
  INV_X1 U153 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U154 ( .A1(data_in[5]), .A2(n831), .B1(n1006), .B2(\mem[11][5] ), 
        .ZN(n1001) );
  INV_X1 U155 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U156 ( .A1(data_in[6]), .A2(n831), .B1(n1006), .B2(\mem[11][6] ), 
        .ZN(n1000) );
  INV_X1 U157 ( .A(n999), .ZN(n715) );
  AOI22_X1 U158 ( .A1(data_in[7]), .A2(n831), .B1(n1006), .B2(\mem[11][7] ), 
        .ZN(n999) );
  INV_X1 U159 ( .A(n952), .ZN(n674) );
  AOI22_X1 U160 ( .A1(data_in[0]), .A2(n825), .B1(n951), .B2(\mem[17][0] ), 
        .ZN(n952) );
  INV_X1 U161 ( .A(n950), .ZN(n673) );
  AOI22_X1 U162 ( .A1(data_in[1]), .A2(n825), .B1(n951), .B2(\mem[17][1] ), 
        .ZN(n950) );
  INV_X1 U163 ( .A(n949), .ZN(n672) );
  AOI22_X1 U164 ( .A1(data_in[2]), .A2(n825), .B1(n951), .B2(\mem[17][2] ), 
        .ZN(n949) );
  INV_X1 U165 ( .A(n948), .ZN(n671) );
  AOI22_X1 U166 ( .A1(data_in[3]), .A2(n825), .B1(n951), .B2(\mem[17][3] ), 
        .ZN(n948) );
  INV_X1 U167 ( .A(n947), .ZN(n670) );
  AOI22_X1 U168 ( .A1(data_in[4]), .A2(n825), .B1(n951), .B2(\mem[17][4] ), 
        .ZN(n947) );
  INV_X1 U169 ( .A(n946), .ZN(n669) );
  AOI22_X1 U170 ( .A1(data_in[5]), .A2(n825), .B1(n951), .B2(\mem[17][5] ), 
        .ZN(n946) );
  INV_X1 U171 ( .A(n945), .ZN(n668) );
  AOI22_X1 U172 ( .A1(data_in[6]), .A2(n825), .B1(n951), .B2(\mem[17][6] ), 
        .ZN(n945) );
  INV_X1 U173 ( .A(n944), .ZN(n667) );
  AOI22_X1 U174 ( .A1(data_in[7]), .A2(n825), .B1(n951), .B2(\mem[17][7] ), 
        .ZN(n944) );
  INV_X1 U175 ( .A(n916), .ZN(n642) );
  AOI22_X1 U176 ( .A1(data_in[0]), .A2(n821), .B1(n915), .B2(\mem[21][0] ), 
        .ZN(n916) );
  INV_X1 U177 ( .A(n914), .ZN(n641) );
  AOI22_X1 U178 ( .A1(data_in[1]), .A2(n821), .B1(n915), .B2(\mem[21][1] ), 
        .ZN(n914) );
  INV_X1 U179 ( .A(n913), .ZN(n640) );
  AOI22_X1 U180 ( .A1(data_in[2]), .A2(n821), .B1(n915), .B2(\mem[21][2] ), 
        .ZN(n913) );
  INV_X1 U181 ( .A(n912), .ZN(n639) );
  AOI22_X1 U182 ( .A1(data_in[3]), .A2(n821), .B1(n915), .B2(\mem[21][3] ), 
        .ZN(n912) );
  INV_X1 U183 ( .A(n911), .ZN(n638) );
  AOI22_X1 U184 ( .A1(data_in[4]), .A2(n821), .B1(n915), .B2(\mem[21][4] ), 
        .ZN(n911) );
  INV_X1 U185 ( .A(n910), .ZN(n637) );
  AOI22_X1 U186 ( .A1(data_in[5]), .A2(n821), .B1(n915), .B2(\mem[21][5] ), 
        .ZN(n910) );
  INV_X1 U187 ( .A(n909), .ZN(n636) );
  AOI22_X1 U188 ( .A1(data_in[6]), .A2(n821), .B1(n915), .B2(\mem[21][6] ), 
        .ZN(n909) );
  INV_X1 U189 ( .A(n908), .ZN(n635) );
  AOI22_X1 U190 ( .A1(data_in[7]), .A2(n821), .B1(n915), .B2(\mem[21][7] ), 
        .ZN(n908) );
  INV_X1 U191 ( .A(n1025), .ZN(n738) );
  AOI22_X1 U192 ( .A1(data_in[0]), .A2(n833), .B1(n1024), .B2(\mem[9][0] ), 
        .ZN(n1025) );
  INV_X1 U193 ( .A(n1023), .ZN(n737) );
  AOI22_X1 U194 ( .A1(data_in[1]), .A2(n833), .B1(n1024), .B2(\mem[9][1] ), 
        .ZN(n1023) );
  INV_X1 U195 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U196 ( .A1(data_in[2]), .A2(n833), .B1(n1024), .B2(\mem[9][2] ), 
        .ZN(n1022) );
  INV_X1 U197 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U198 ( .A1(data_in[3]), .A2(n833), .B1(n1024), .B2(\mem[9][3] ), 
        .ZN(n1021) );
  INV_X1 U199 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U200 ( .A1(data_in[4]), .A2(n833), .B1(n1024), .B2(\mem[9][4] ), 
        .ZN(n1020) );
  INV_X1 U201 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U202 ( .A1(data_in[0]), .A2(n836), .B1(n1052), .B2(\mem[6][0] ), 
        .ZN(n1053) );
  INV_X1 U203 ( .A(n1051), .ZN(n761) );
  AOI22_X1 U204 ( .A1(data_in[1]), .A2(n836), .B1(n1052), .B2(\mem[6][1] ), 
        .ZN(n1051) );
  INV_X1 U205 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U206 ( .A1(data_in[2]), .A2(n836), .B1(n1052), .B2(\mem[6][2] ), 
        .ZN(n1050) );
  INV_X1 U207 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U208 ( .A1(data_in[3]), .A2(n836), .B1(n1052), .B2(\mem[6][3] ), 
        .ZN(n1049) );
  INV_X1 U209 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U210 ( .A1(data_in[4]), .A2(n836), .B1(n1052), .B2(\mem[6][4] ), 
        .ZN(n1048) );
  INV_X1 U211 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U212 ( .A1(data_in[5]), .A2(n836), .B1(n1052), .B2(\mem[6][5] ), 
        .ZN(n1047) );
  INV_X1 U213 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U214 ( .A1(data_in[6]), .A2(n836), .B1(n1052), .B2(\mem[6][6] ), 
        .ZN(n1046) );
  INV_X1 U215 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U216 ( .A1(data_in[7]), .A2(n836), .B1(n1052), .B2(\mem[6][7] ), 
        .ZN(n1045) );
  INV_X1 U217 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U218 ( .A1(data_in[0]), .A2(n835), .B1(n1043), .B2(\mem[7][0] ), 
        .ZN(n1044) );
  INV_X1 U219 ( .A(n1042), .ZN(n753) );
  AOI22_X1 U220 ( .A1(data_in[1]), .A2(n835), .B1(n1043), .B2(\mem[7][1] ), 
        .ZN(n1042) );
  INV_X1 U221 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U222 ( .A1(data_in[2]), .A2(n835), .B1(n1043), .B2(\mem[7][2] ), 
        .ZN(n1041) );
  INV_X1 U223 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U224 ( .A1(data_in[3]), .A2(n835), .B1(n1043), .B2(\mem[7][3] ), 
        .ZN(n1040) );
  INV_X1 U225 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U226 ( .A1(data_in[4]), .A2(n835), .B1(n1043), .B2(\mem[7][4] ), 
        .ZN(n1039) );
  INV_X1 U227 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U228 ( .A1(data_in[5]), .A2(n835), .B1(n1043), .B2(\mem[7][5] ), 
        .ZN(n1038) );
  INV_X1 U229 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U230 ( .A1(data_in[6]), .A2(n835), .B1(n1043), .B2(\mem[7][6] ), 
        .ZN(n1037) );
  INV_X1 U231 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U232 ( .A1(data_in[7]), .A2(n835), .B1(n1043), .B2(\mem[7][7] ), 
        .ZN(n1036) );
  INV_X1 U233 ( .A(n980), .ZN(n698) );
  AOI22_X1 U234 ( .A1(data_in[0]), .A2(n828), .B1(n979), .B2(\mem[14][0] ), 
        .ZN(n980) );
  INV_X1 U235 ( .A(n978), .ZN(n697) );
  AOI22_X1 U236 ( .A1(data_in[1]), .A2(n828), .B1(n979), .B2(\mem[14][1] ), 
        .ZN(n978) );
  INV_X1 U237 ( .A(n977), .ZN(n696) );
  AOI22_X1 U238 ( .A1(data_in[2]), .A2(n828), .B1(n979), .B2(\mem[14][2] ), 
        .ZN(n977) );
  INV_X1 U239 ( .A(n976), .ZN(n695) );
  AOI22_X1 U240 ( .A1(data_in[3]), .A2(n828), .B1(n979), .B2(\mem[14][3] ), 
        .ZN(n976) );
  INV_X1 U241 ( .A(n975), .ZN(n694) );
  AOI22_X1 U242 ( .A1(data_in[4]), .A2(n828), .B1(n979), .B2(\mem[14][4] ), 
        .ZN(n975) );
  INV_X1 U243 ( .A(n974), .ZN(n693) );
  AOI22_X1 U244 ( .A1(data_in[5]), .A2(n828), .B1(n979), .B2(\mem[14][5] ), 
        .ZN(n974) );
  INV_X1 U245 ( .A(n973), .ZN(n692) );
  AOI22_X1 U246 ( .A1(data_in[6]), .A2(n828), .B1(n979), .B2(\mem[14][6] ), 
        .ZN(n973) );
  INV_X1 U247 ( .A(n972), .ZN(n691) );
  AOI22_X1 U248 ( .A1(data_in[7]), .A2(n828), .B1(n979), .B2(\mem[14][7] ), 
        .ZN(n972) );
  INV_X1 U249 ( .A(n971), .ZN(n690) );
  AOI22_X1 U250 ( .A1(data_in[0]), .A2(n827), .B1(n970), .B2(\mem[15][0] ), 
        .ZN(n971) );
  INV_X1 U251 ( .A(n969), .ZN(n689) );
  AOI22_X1 U252 ( .A1(data_in[1]), .A2(n827), .B1(n970), .B2(\mem[15][1] ), 
        .ZN(n969) );
  INV_X1 U253 ( .A(n968), .ZN(n688) );
  AOI22_X1 U254 ( .A1(data_in[2]), .A2(n827), .B1(n970), .B2(\mem[15][2] ), 
        .ZN(n968) );
  INV_X1 U255 ( .A(n967), .ZN(n687) );
  AOI22_X1 U256 ( .A1(data_in[3]), .A2(n827), .B1(n970), .B2(\mem[15][3] ), 
        .ZN(n967) );
  INV_X1 U257 ( .A(n966), .ZN(n686) );
  AOI22_X1 U258 ( .A1(data_in[4]), .A2(n827), .B1(n970), .B2(\mem[15][4] ), 
        .ZN(n966) );
  INV_X1 U259 ( .A(n965), .ZN(n685) );
  AOI22_X1 U260 ( .A1(data_in[5]), .A2(n827), .B1(n970), .B2(\mem[15][5] ), 
        .ZN(n965) );
  INV_X1 U261 ( .A(n964), .ZN(n684) );
  AOI22_X1 U262 ( .A1(data_in[6]), .A2(n827), .B1(n970), .B2(\mem[15][6] ), 
        .ZN(n964) );
  INV_X1 U263 ( .A(n963), .ZN(n683) );
  AOI22_X1 U264 ( .A1(data_in[7]), .A2(n827), .B1(n970), .B2(\mem[15][7] ), 
        .ZN(n963) );
  INV_X1 U265 ( .A(n943), .ZN(n666) );
  AOI22_X1 U266 ( .A1(data_in[0]), .A2(n824), .B1(n942), .B2(\mem[18][0] ), 
        .ZN(n943) );
  INV_X1 U267 ( .A(n941), .ZN(n665) );
  AOI22_X1 U268 ( .A1(data_in[1]), .A2(n824), .B1(n942), .B2(\mem[18][1] ), 
        .ZN(n941) );
  INV_X1 U269 ( .A(n940), .ZN(n664) );
  AOI22_X1 U270 ( .A1(data_in[2]), .A2(n824), .B1(n942), .B2(\mem[18][2] ), 
        .ZN(n940) );
  INV_X1 U271 ( .A(n939), .ZN(n663) );
  AOI22_X1 U272 ( .A1(data_in[3]), .A2(n824), .B1(n942), .B2(\mem[18][3] ), 
        .ZN(n939) );
  INV_X1 U273 ( .A(n938), .ZN(n662) );
  AOI22_X1 U274 ( .A1(data_in[4]), .A2(n824), .B1(n942), .B2(\mem[18][4] ), 
        .ZN(n938) );
  INV_X1 U275 ( .A(n937), .ZN(n661) );
  AOI22_X1 U276 ( .A1(data_in[5]), .A2(n824), .B1(n942), .B2(\mem[18][5] ), 
        .ZN(n937) );
  INV_X1 U277 ( .A(n936), .ZN(n660) );
  AOI22_X1 U278 ( .A1(data_in[6]), .A2(n824), .B1(n942), .B2(\mem[18][6] ), 
        .ZN(n936) );
  INV_X1 U279 ( .A(n935), .ZN(n659) );
  AOI22_X1 U280 ( .A1(data_in[7]), .A2(n824), .B1(n942), .B2(\mem[18][7] ), 
        .ZN(n935) );
  INV_X1 U281 ( .A(n934), .ZN(n658) );
  AOI22_X1 U282 ( .A1(data_in[0]), .A2(n823), .B1(n933), .B2(\mem[19][0] ), 
        .ZN(n934) );
  INV_X1 U283 ( .A(n932), .ZN(n657) );
  AOI22_X1 U284 ( .A1(data_in[1]), .A2(n823), .B1(n933), .B2(\mem[19][1] ), 
        .ZN(n932) );
  INV_X1 U285 ( .A(n931), .ZN(n656) );
  AOI22_X1 U286 ( .A1(data_in[2]), .A2(n823), .B1(n933), .B2(\mem[19][2] ), 
        .ZN(n931) );
  INV_X1 U287 ( .A(n930), .ZN(n655) );
  AOI22_X1 U288 ( .A1(data_in[3]), .A2(n823), .B1(n933), .B2(\mem[19][3] ), 
        .ZN(n930) );
  INV_X1 U289 ( .A(n929), .ZN(n654) );
  AOI22_X1 U290 ( .A1(data_in[4]), .A2(n823), .B1(n933), .B2(\mem[19][4] ), 
        .ZN(n929) );
  INV_X1 U291 ( .A(n928), .ZN(n653) );
  AOI22_X1 U292 ( .A1(data_in[5]), .A2(n823), .B1(n933), .B2(\mem[19][5] ), 
        .ZN(n928) );
  INV_X1 U293 ( .A(n927), .ZN(n652) );
  AOI22_X1 U294 ( .A1(data_in[6]), .A2(n823), .B1(n933), .B2(\mem[19][6] ), 
        .ZN(n927) );
  INV_X1 U295 ( .A(n926), .ZN(n651) );
  AOI22_X1 U296 ( .A1(data_in[7]), .A2(n823), .B1(n933), .B2(\mem[19][7] ), 
        .ZN(n926) );
  INV_X1 U297 ( .A(n907), .ZN(n634) );
  AOI22_X1 U298 ( .A1(data_in[0]), .A2(n820), .B1(n906), .B2(\mem[22][0] ), 
        .ZN(n907) );
  INV_X1 U299 ( .A(n905), .ZN(n633) );
  AOI22_X1 U300 ( .A1(data_in[1]), .A2(n820), .B1(n906), .B2(\mem[22][1] ), 
        .ZN(n905) );
  INV_X1 U301 ( .A(n904), .ZN(n632) );
  AOI22_X1 U302 ( .A1(data_in[2]), .A2(n820), .B1(n906), .B2(\mem[22][2] ), 
        .ZN(n904) );
  INV_X1 U303 ( .A(n903), .ZN(n631) );
  AOI22_X1 U304 ( .A1(data_in[3]), .A2(n820), .B1(n906), .B2(\mem[22][3] ), 
        .ZN(n903) );
  INV_X1 U305 ( .A(n902), .ZN(n630) );
  AOI22_X1 U306 ( .A1(data_in[4]), .A2(n820), .B1(n906), .B2(\mem[22][4] ), 
        .ZN(n902) );
  INV_X1 U307 ( .A(n901), .ZN(n629) );
  AOI22_X1 U308 ( .A1(data_in[5]), .A2(n820), .B1(n906), .B2(\mem[22][5] ), 
        .ZN(n901) );
  INV_X1 U309 ( .A(n900), .ZN(n628) );
  AOI22_X1 U310 ( .A1(data_in[6]), .A2(n820), .B1(n906), .B2(\mem[22][6] ), 
        .ZN(n900) );
  INV_X1 U311 ( .A(n899), .ZN(n627) );
  AOI22_X1 U312 ( .A1(data_in[7]), .A2(n820), .B1(n906), .B2(\mem[22][7] ), 
        .ZN(n899) );
  INV_X1 U313 ( .A(n896), .ZN(n625) );
  AOI22_X1 U314 ( .A1(data_in[1]), .A2(n819), .B1(n897), .B2(\mem[23][1] ), 
        .ZN(n896) );
  INV_X1 U315 ( .A(n895), .ZN(n624) );
  AOI22_X1 U316 ( .A1(data_in[2]), .A2(n819), .B1(n897), .B2(\mem[23][2] ), 
        .ZN(n895) );
  INV_X1 U317 ( .A(n894), .ZN(n623) );
  AOI22_X1 U318 ( .A1(data_in[3]), .A2(n819), .B1(n897), .B2(\mem[23][3] ), 
        .ZN(n894) );
  INV_X1 U319 ( .A(n893), .ZN(n622) );
  AOI22_X1 U320 ( .A1(data_in[4]), .A2(n819), .B1(n897), .B2(\mem[23][4] ), 
        .ZN(n893) );
  INV_X1 U321 ( .A(n892), .ZN(n621) );
  AOI22_X1 U322 ( .A1(data_in[5]), .A2(n819), .B1(n897), .B2(\mem[23][5] ), 
        .ZN(n892) );
  INV_X1 U323 ( .A(n891), .ZN(n620) );
  AOI22_X1 U324 ( .A1(data_in[6]), .A2(n819), .B1(n897), .B2(\mem[23][6] ), 
        .ZN(n891) );
  INV_X1 U325 ( .A(n890), .ZN(n619) );
  AOI22_X1 U326 ( .A1(data_in[7]), .A2(n819), .B1(n897), .B2(\mem[23][7] ), 
        .ZN(n890) );
  INV_X1 U327 ( .A(n898), .ZN(n626) );
  AOI22_X1 U328 ( .A1(data_in[0]), .A2(n819), .B1(n897), .B2(\mem[23][0] ), 
        .ZN(n898) );
  INV_X1 U329 ( .A(N12), .ZN(n254) );
  INV_X1 U330 ( .A(N11), .ZN(n253) );
  INV_X1 U331 ( .A(n998), .ZN(n714) );
  AOI22_X1 U332 ( .A1(data_in[0]), .A2(n830), .B1(n997), .B2(\mem[12][0] ), 
        .ZN(n998) );
  INV_X1 U333 ( .A(n996), .ZN(n713) );
  AOI22_X1 U334 ( .A1(data_in[1]), .A2(n830), .B1(n997), .B2(\mem[12][1] ), 
        .ZN(n996) );
  INV_X1 U335 ( .A(n995), .ZN(n712) );
  AOI22_X1 U336 ( .A1(data_in[2]), .A2(n830), .B1(n997), .B2(\mem[12][2] ), 
        .ZN(n995) );
  INV_X1 U337 ( .A(n994), .ZN(n711) );
  AOI22_X1 U338 ( .A1(data_in[3]), .A2(n830), .B1(n997), .B2(\mem[12][3] ), 
        .ZN(n994) );
  INV_X1 U339 ( .A(n993), .ZN(n710) );
  AOI22_X1 U340 ( .A1(data_in[4]), .A2(n830), .B1(n997), .B2(\mem[12][4] ), 
        .ZN(n993) );
  INV_X1 U341 ( .A(n992), .ZN(n709) );
  AOI22_X1 U342 ( .A1(data_in[5]), .A2(n830), .B1(n997), .B2(\mem[12][5] ), 
        .ZN(n992) );
  INV_X1 U343 ( .A(n991), .ZN(n708) );
  AOI22_X1 U344 ( .A1(data_in[6]), .A2(n830), .B1(n997), .B2(\mem[12][6] ), 
        .ZN(n991) );
  INV_X1 U345 ( .A(n990), .ZN(n707) );
  AOI22_X1 U346 ( .A1(data_in[7]), .A2(n830), .B1(n997), .B2(\mem[12][7] ), 
        .ZN(n990) );
  INV_X1 U347 ( .A(n925), .ZN(n650) );
  AOI22_X1 U348 ( .A1(data_in[0]), .A2(n822), .B1(n924), .B2(\mem[20][0] ), 
        .ZN(n925) );
  INV_X1 U349 ( .A(n923), .ZN(n649) );
  AOI22_X1 U350 ( .A1(data_in[1]), .A2(n822), .B1(n924), .B2(\mem[20][1] ), 
        .ZN(n923) );
  INV_X1 U351 ( .A(n922), .ZN(n648) );
  AOI22_X1 U352 ( .A1(data_in[2]), .A2(n822), .B1(n924), .B2(\mem[20][2] ), 
        .ZN(n922) );
  INV_X1 U353 ( .A(n921), .ZN(n647) );
  AOI22_X1 U354 ( .A1(data_in[3]), .A2(n822), .B1(n924), .B2(\mem[20][3] ), 
        .ZN(n921) );
  INV_X1 U355 ( .A(n920), .ZN(n646) );
  AOI22_X1 U356 ( .A1(data_in[4]), .A2(n822), .B1(n924), .B2(\mem[20][4] ), 
        .ZN(n920) );
  INV_X1 U357 ( .A(n919), .ZN(n645) );
  AOI22_X1 U358 ( .A1(data_in[5]), .A2(n822), .B1(n924), .B2(\mem[20][5] ), 
        .ZN(n919) );
  INV_X1 U359 ( .A(n918), .ZN(n644) );
  AOI22_X1 U360 ( .A1(data_in[6]), .A2(n822), .B1(n924), .B2(\mem[20][6] ), 
        .ZN(n918) );
  INV_X1 U361 ( .A(n917), .ZN(n643) );
  AOI22_X1 U362 ( .A1(data_in[7]), .A2(n822), .B1(n924), .B2(\mem[20][7] ), 
        .ZN(n917) );
  INV_X1 U363 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U364 ( .A1(data_in[0]), .A2(n834), .B1(n1034), .B2(\mem[8][0] ), 
        .ZN(n1035) );
  INV_X1 U365 ( .A(n1033), .ZN(n745) );
  AOI22_X1 U366 ( .A1(data_in[1]), .A2(n834), .B1(n1034), .B2(\mem[8][1] ), 
        .ZN(n1033) );
  INV_X1 U367 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U368 ( .A1(data_in[2]), .A2(n834), .B1(n1034), .B2(\mem[8][2] ), 
        .ZN(n1032) );
  INV_X1 U369 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U370 ( .A1(data_in[3]), .A2(n834), .B1(n1034), .B2(\mem[8][3] ), 
        .ZN(n1031) );
  INV_X1 U371 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U372 ( .A1(data_in[4]), .A2(n834), .B1(n1034), .B2(\mem[8][4] ), 
        .ZN(n1030) );
  INV_X1 U373 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U374 ( .A1(data_in[5]), .A2(n834), .B1(n1034), .B2(\mem[8][5] ), 
        .ZN(n1029) );
  INV_X1 U375 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U376 ( .A1(data_in[6]), .A2(n834), .B1(n1034), .B2(\mem[8][6] ), 
        .ZN(n1028) );
  INV_X1 U377 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U378 ( .A1(data_in[7]), .A2(n834), .B1(n1034), .B2(\mem[8][7] ), 
        .ZN(n1027) );
  INV_X1 U379 ( .A(n962), .ZN(n682) );
  AOI22_X1 U380 ( .A1(data_in[0]), .A2(n826), .B1(n961), .B2(\mem[16][0] ), 
        .ZN(n962) );
  INV_X1 U381 ( .A(n960), .ZN(n681) );
  AOI22_X1 U382 ( .A1(data_in[1]), .A2(n826), .B1(n961), .B2(\mem[16][1] ), 
        .ZN(n960) );
  INV_X1 U383 ( .A(n959), .ZN(n680) );
  AOI22_X1 U384 ( .A1(data_in[2]), .A2(n826), .B1(n961), .B2(\mem[16][2] ), 
        .ZN(n959) );
  INV_X1 U385 ( .A(n958), .ZN(n679) );
  AOI22_X1 U386 ( .A1(data_in[3]), .A2(n826), .B1(n961), .B2(\mem[16][3] ), 
        .ZN(n958) );
  INV_X1 U387 ( .A(n957), .ZN(n678) );
  AOI22_X1 U388 ( .A1(data_in[4]), .A2(n826), .B1(n961), .B2(\mem[16][4] ), 
        .ZN(n957) );
  INV_X1 U389 ( .A(n956), .ZN(n677) );
  AOI22_X1 U390 ( .A1(data_in[5]), .A2(n826), .B1(n961), .B2(\mem[16][5] ), 
        .ZN(n956) );
  INV_X1 U391 ( .A(n955), .ZN(n676) );
  AOI22_X1 U392 ( .A1(data_in[6]), .A2(n826), .B1(n961), .B2(\mem[16][6] ), 
        .ZN(n955) );
  INV_X1 U393 ( .A(n954), .ZN(n675) );
  AOI22_X1 U394 ( .A1(data_in[7]), .A2(n826), .B1(n961), .B2(\mem[16][7] ), 
        .ZN(n954) );
  INV_X1 U395 ( .A(n889), .ZN(n618) );
  AOI22_X1 U396 ( .A1(data_in[0]), .A2(n815), .B1(n888), .B2(\mem[24][0] ), 
        .ZN(n889) );
  INV_X1 U397 ( .A(n887), .ZN(n617) );
  AOI22_X1 U398 ( .A1(data_in[1]), .A2(n815), .B1(n888), .B2(\mem[24][1] ), 
        .ZN(n887) );
  INV_X1 U399 ( .A(n886), .ZN(n616) );
  AOI22_X1 U400 ( .A1(data_in[2]), .A2(n815), .B1(n888), .B2(\mem[24][2] ), 
        .ZN(n886) );
  INV_X1 U401 ( .A(n885), .ZN(n615) );
  AOI22_X1 U402 ( .A1(data_in[3]), .A2(n815), .B1(n888), .B2(\mem[24][3] ), 
        .ZN(n885) );
  INV_X1 U403 ( .A(n884), .ZN(n614) );
  AOI22_X1 U404 ( .A1(data_in[4]), .A2(n815), .B1(n888), .B2(\mem[24][4] ), 
        .ZN(n884) );
  INV_X1 U405 ( .A(n883), .ZN(n613) );
  AOI22_X1 U406 ( .A1(data_in[5]), .A2(n815), .B1(n888), .B2(\mem[24][5] ), 
        .ZN(n883) );
  INV_X1 U407 ( .A(n882), .ZN(n612) );
  AOI22_X1 U408 ( .A1(data_in[6]), .A2(n815), .B1(n888), .B2(\mem[24][6] ), 
        .ZN(n882) );
  INV_X1 U409 ( .A(n881), .ZN(n611) );
  AOI22_X1 U410 ( .A1(data_in[7]), .A2(n815), .B1(n888), .B2(\mem[24][7] ), 
        .ZN(n881) );
  INV_X1 U411 ( .A(n880), .ZN(n610) );
  AOI22_X1 U412 ( .A1(data_in[0]), .A2(n814), .B1(n879), .B2(\mem[25][0] ), 
        .ZN(n880) );
  INV_X1 U413 ( .A(n878), .ZN(n609) );
  AOI22_X1 U414 ( .A1(data_in[1]), .A2(n814), .B1(n879), .B2(\mem[25][1] ), 
        .ZN(n878) );
  INV_X1 U415 ( .A(n877), .ZN(n608) );
  AOI22_X1 U416 ( .A1(data_in[2]), .A2(n814), .B1(n879), .B2(\mem[25][2] ), 
        .ZN(n877) );
  INV_X1 U417 ( .A(n876), .ZN(n607) );
  AOI22_X1 U418 ( .A1(data_in[3]), .A2(n814), .B1(n879), .B2(\mem[25][3] ), 
        .ZN(n876) );
  INV_X1 U419 ( .A(n875), .ZN(n606) );
  AOI22_X1 U420 ( .A1(data_in[4]), .A2(n814), .B1(n879), .B2(\mem[25][4] ), 
        .ZN(n875) );
  INV_X1 U421 ( .A(n874), .ZN(n605) );
  AOI22_X1 U422 ( .A1(data_in[5]), .A2(n814), .B1(n879), .B2(\mem[25][5] ), 
        .ZN(n874) );
  INV_X1 U423 ( .A(n873), .ZN(n604) );
  AOI22_X1 U424 ( .A1(data_in[6]), .A2(n814), .B1(n879), .B2(\mem[25][6] ), 
        .ZN(n873) );
  INV_X1 U425 ( .A(n872), .ZN(n603) );
  AOI22_X1 U426 ( .A1(data_in[7]), .A2(n814), .B1(n879), .B2(\mem[25][7] ), 
        .ZN(n872) );
  INV_X1 U427 ( .A(n871), .ZN(n602) );
  AOI22_X1 U428 ( .A1(data_in[0]), .A2(n813), .B1(n870), .B2(\mem[26][0] ), 
        .ZN(n871) );
  INV_X1 U429 ( .A(n869), .ZN(n601) );
  AOI22_X1 U430 ( .A1(data_in[1]), .A2(n813), .B1(n870), .B2(\mem[26][1] ), 
        .ZN(n869) );
  INV_X1 U431 ( .A(n868), .ZN(n600) );
  AOI22_X1 U432 ( .A1(data_in[2]), .A2(n813), .B1(n870), .B2(\mem[26][2] ), 
        .ZN(n868) );
  INV_X1 U433 ( .A(n867), .ZN(n599) );
  AOI22_X1 U434 ( .A1(data_in[3]), .A2(n813), .B1(n870), .B2(\mem[26][3] ), 
        .ZN(n867) );
  INV_X1 U435 ( .A(n866), .ZN(n598) );
  AOI22_X1 U436 ( .A1(data_in[4]), .A2(n813), .B1(n870), .B2(\mem[26][4] ), 
        .ZN(n866) );
  INV_X1 U437 ( .A(n865), .ZN(n597) );
  AOI22_X1 U438 ( .A1(data_in[5]), .A2(n813), .B1(n870), .B2(\mem[26][5] ), 
        .ZN(n865) );
  INV_X1 U439 ( .A(n864), .ZN(n596) );
  AOI22_X1 U440 ( .A1(data_in[6]), .A2(n813), .B1(n870), .B2(\mem[26][6] ), 
        .ZN(n864) );
  INV_X1 U441 ( .A(n863), .ZN(n595) );
  AOI22_X1 U442 ( .A1(data_in[7]), .A2(n813), .B1(n870), .B2(\mem[26][7] ), 
        .ZN(n863) );
  INV_X1 U443 ( .A(n862), .ZN(n594) );
  AOI22_X1 U444 ( .A1(data_in[0]), .A2(n812), .B1(n861), .B2(\mem[27][0] ), 
        .ZN(n862) );
  INV_X1 U445 ( .A(n860), .ZN(n293) );
  AOI22_X1 U446 ( .A1(data_in[1]), .A2(n812), .B1(n861), .B2(\mem[27][1] ), 
        .ZN(n860) );
  INV_X1 U447 ( .A(n859), .ZN(n292) );
  AOI22_X1 U448 ( .A1(data_in[2]), .A2(n812), .B1(n861), .B2(\mem[27][2] ), 
        .ZN(n859) );
  INV_X1 U449 ( .A(n858), .ZN(n291) );
  AOI22_X1 U450 ( .A1(data_in[3]), .A2(n812), .B1(n861), .B2(\mem[27][3] ), 
        .ZN(n858) );
  INV_X1 U451 ( .A(n857), .ZN(n290) );
  AOI22_X1 U452 ( .A1(data_in[4]), .A2(n812), .B1(n861), .B2(\mem[27][4] ), 
        .ZN(n857) );
  INV_X1 U453 ( .A(n856), .ZN(n289) );
  AOI22_X1 U454 ( .A1(data_in[5]), .A2(n812), .B1(n861), .B2(\mem[27][5] ), 
        .ZN(n856) );
  INV_X1 U455 ( .A(n855), .ZN(n288) );
  AOI22_X1 U456 ( .A1(data_in[6]), .A2(n812), .B1(n861), .B2(\mem[27][6] ), 
        .ZN(n855) );
  INV_X1 U457 ( .A(n854), .ZN(n287) );
  AOI22_X1 U458 ( .A1(data_in[7]), .A2(n812), .B1(n861), .B2(\mem[27][7] ), 
        .ZN(n854) );
  INV_X1 U459 ( .A(n853), .ZN(n286) );
  AOI22_X1 U460 ( .A1(data_in[0]), .A2(n811), .B1(n852), .B2(\mem[28][0] ), 
        .ZN(n853) );
  INV_X1 U461 ( .A(n851), .ZN(n285) );
  AOI22_X1 U462 ( .A1(data_in[1]), .A2(n811), .B1(n852), .B2(\mem[28][1] ), 
        .ZN(n851) );
  INV_X1 U463 ( .A(n850), .ZN(n284) );
  AOI22_X1 U464 ( .A1(data_in[2]), .A2(n811), .B1(n852), .B2(\mem[28][2] ), 
        .ZN(n850) );
  INV_X1 U465 ( .A(n849), .ZN(n283) );
  AOI22_X1 U466 ( .A1(data_in[3]), .A2(n811), .B1(n852), .B2(\mem[28][3] ), 
        .ZN(n849) );
  INV_X1 U467 ( .A(n848), .ZN(n282) );
  AOI22_X1 U468 ( .A1(data_in[4]), .A2(n811), .B1(n852), .B2(\mem[28][4] ), 
        .ZN(n848) );
  INV_X1 U469 ( .A(n847), .ZN(n281) );
  AOI22_X1 U470 ( .A1(data_in[5]), .A2(n811), .B1(n852), .B2(\mem[28][5] ), 
        .ZN(n847) );
  INV_X1 U471 ( .A(n846), .ZN(n280) );
  AOI22_X1 U472 ( .A1(data_in[6]), .A2(n811), .B1(n852), .B2(\mem[28][6] ), 
        .ZN(n846) );
  INV_X1 U473 ( .A(n845), .ZN(n279) );
  AOI22_X1 U474 ( .A1(data_in[7]), .A2(n811), .B1(n852), .B2(\mem[28][7] ), 
        .ZN(n845) );
  INV_X1 U475 ( .A(n1144), .ZN(n278) );
  AOI22_X1 U476 ( .A1(n818), .A2(data_in[0]), .B1(n1143), .B2(\mem[29][0] ), 
        .ZN(n1144) );
  INV_X1 U477 ( .A(n1142), .ZN(n277) );
  AOI22_X1 U478 ( .A1(n818), .A2(data_in[1]), .B1(n1143), .B2(\mem[29][1] ), 
        .ZN(n1142) );
  INV_X1 U479 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U480 ( .A1(n818), .A2(data_in[2]), .B1(n1143), .B2(\mem[29][2] ), 
        .ZN(n1141) );
  INV_X1 U481 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U482 ( .A1(n818), .A2(data_in[3]), .B1(n1143), .B2(\mem[29][3] ), 
        .ZN(n1140) );
  INV_X1 U483 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U484 ( .A1(n818), .A2(data_in[4]), .B1(n1143), .B2(\mem[29][4] ), 
        .ZN(n1139) );
  INV_X1 U485 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U486 ( .A1(n818), .A2(data_in[5]), .B1(n1143), .B2(\mem[29][5] ), 
        .ZN(n1138) );
  INV_X1 U487 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U488 ( .A1(n818), .A2(data_in[6]), .B1(n1143), .B2(\mem[29][6] ), 
        .ZN(n1137) );
  INV_X1 U489 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U490 ( .A1(n818), .A2(data_in[7]), .B1(n1143), .B2(\mem[29][7] ), 
        .ZN(n1136) );
  INV_X1 U491 ( .A(n1133), .ZN(n270) );
  AOI22_X1 U492 ( .A1(data_in[0]), .A2(n817), .B1(n1132), .B2(\mem[30][0] ), 
        .ZN(n1133) );
  INV_X1 U493 ( .A(n1131), .ZN(n269) );
  AOI22_X1 U494 ( .A1(data_in[1]), .A2(n817), .B1(n1132), .B2(\mem[30][1] ), 
        .ZN(n1131) );
  INV_X1 U495 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U496 ( .A1(data_in[2]), .A2(n817), .B1(n1132), .B2(\mem[30][2] ), 
        .ZN(n1130) );
  INV_X1 U497 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U498 ( .A1(data_in[3]), .A2(n817), .B1(n1132), .B2(\mem[30][3] ), 
        .ZN(n1129) );
  INV_X1 U499 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U500 ( .A1(data_in[4]), .A2(n817), .B1(n1132), .B2(\mem[30][4] ), 
        .ZN(n1128) );
  INV_X1 U501 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U502 ( .A1(data_in[5]), .A2(n817), .B1(n1132), .B2(\mem[30][5] ), 
        .ZN(n1127) );
  INV_X1 U503 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U504 ( .A1(data_in[6]), .A2(n817), .B1(n1132), .B2(\mem[30][6] ), 
        .ZN(n1126) );
  INV_X1 U505 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U506 ( .A1(data_in[7]), .A2(n817), .B1(n1132), .B2(\mem[30][7] ), 
        .ZN(n1125) );
  INV_X1 U507 ( .A(n1123), .ZN(n262) );
  AOI22_X1 U508 ( .A1(data_in[0]), .A2(n816), .B1(n1122), .B2(\mem[31][0] ), 
        .ZN(n1123) );
  INV_X1 U509 ( .A(n1121), .ZN(n261) );
  AOI22_X1 U510 ( .A1(data_in[1]), .A2(n816), .B1(n1122), .B2(\mem[31][1] ), 
        .ZN(n1121) );
  INV_X1 U511 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U512 ( .A1(data_in[2]), .A2(n816), .B1(n1122), .B2(\mem[31][2] ), 
        .ZN(n1120) );
  INV_X1 U513 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U514 ( .A1(data_in[3]), .A2(n816), .B1(n1122), .B2(\mem[31][3] ), 
        .ZN(n1119) );
  INV_X1 U515 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U516 ( .A1(data_in[4]), .A2(n816), .B1(n1122), .B2(\mem[31][4] ), 
        .ZN(n1118) );
  INV_X1 U517 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U518 ( .A1(data_in[5]), .A2(n816), .B1(n1122), .B2(\mem[31][5] ), 
        .ZN(n1117) );
  INV_X1 U519 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U520 ( .A1(data_in[6]), .A2(n816), .B1(n1122), .B2(\mem[31][6] ), 
        .ZN(n1116) );
  INV_X1 U521 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U522 ( .A1(data_in[7]), .A2(n816), .B1(n1122), .B2(\mem[31][7] ), 
        .ZN(n1115) );
  INV_X1 U523 ( .A(n1113), .ZN(n810) );
  AOI22_X1 U524 ( .A1(data_in[0]), .A2(n842), .B1(n1112), .B2(\mem[0][0] ), 
        .ZN(n1113) );
  INV_X1 U525 ( .A(n1111), .ZN(n809) );
  AOI22_X1 U526 ( .A1(data_in[1]), .A2(n842), .B1(n1112), .B2(\mem[0][1] ), 
        .ZN(n1111) );
  INV_X1 U527 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U528 ( .A1(data_in[2]), .A2(n842), .B1(n1112), .B2(\mem[0][2] ), 
        .ZN(n1110) );
  INV_X1 U529 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U530 ( .A1(data_in[3]), .A2(n842), .B1(n1112), .B2(\mem[0][3] ), 
        .ZN(n1109) );
  INV_X1 U531 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U532 ( .A1(data_in[4]), .A2(n842), .B1(n1112), .B2(\mem[0][4] ), 
        .ZN(n1108) );
  INV_X1 U533 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U534 ( .A1(data_in[5]), .A2(n842), .B1(n1112), .B2(\mem[0][5] ), 
        .ZN(n1107) );
  INV_X1 U535 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U536 ( .A1(data_in[6]), .A2(n842), .B1(n1112), .B2(\mem[0][6] ), 
        .ZN(n1106) );
  INV_X1 U537 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U538 ( .A1(data_in[7]), .A2(n842), .B1(n1112), .B2(\mem[0][7] ), 
        .ZN(n1105) );
  INV_X1 U539 ( .A(n1102), .ZN(n802) );
  AOI22_X1 U540 ( .A1(data_in[0]), .A2(n841), .B1(n1101), .B2(\mem[1][0] ), 
        .ZN(n1102) );
  INV_X1 U541 ( .A(n1100), .ZN(n801) );
  AOI22_X1 U542 ( .A1(data_in[1]), .A2(n841), .B1(n1101), .B2(\mem[1][1] ), 
        .ZN(n1100) );
  INV_X1 U543 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U544 ( .A1(data_in[2]), .A2(n841), .B1(n1101), .B2(\mem[1][2] ), 
        .ZN(n1099) );
  INV_X1 U545 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U546 ( .A1(data_in[3]), .A2(n841), .B1(n1101), .B2(\mem[1][3] ), 
        .ZN(n1098) );
  INV_X1 U547 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U548 ( .A1(data_in[4]), .A2(n841), .B1(n1101), .B2(\mem[1][4] ), 
        .ZN(n1097) );
  INV_X1 U549 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U550 ( .A1(data_in[5]), .A2(n841), .B1(n1101), .B2(\mem[1][5] ), 
        .ZN(n1096) );
  INV_X1 U551 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U552 ( .A1(data_in[6]), .A2(n841), .B1(n1101), .B2(\mem[1][6] ), 
        .ZN(n1095) );
  INV_X1 U553 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U554 ( .A1(data_in[7]), .A2(n841), .B1(n1101), .B2(\mem[1][7] ), 
        .ZN(n1094) );
  INV_X1 U555 ( .A(n1092), .ZN(n794) );
  AOI22_X1 U556 ( .A1(data_in[0]), .A2(n840), .B1(n1091), .B2(\mem[2][0] ), 
        .ZN(n1092) );
  INV_X1 U557 ( .A(n1090), .ZN(n793) );
  AOI22_X1 U558 ( .A1(data_in[1]), .A2(n840), .B1(n1091), .B2(\mem[2][1] ), 
        .ZN(n1090) );
  INV_X1 U559 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U560 ( .A1(data_in[2]), .A2(n840), .B1(n1091), .B2(\mem[2][2] ), 
        .ZN(n1089) );
  INV_X1 U561 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U562 ( .A1(data_in[3]), .A2(n840), .B1(n1091), .B2(\mem[2][3] ), 
        .ZN(n1088) );
  INV_X1 U563 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U564 ( .A1(data_in[4]), .A2(n840), .B1(n1091), .B2(\mem[2][4] ), 
        .ZN(n1087) );
  INV_X1 U565 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U566 ( .A1(data_in[5]), .A2(n840), .B1(n1091), .B2(\mem[2][5] ), 
        .ZN(n1086) );
  INV_X1 U567 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U568 ( .A1(data_in[6]), .A2(n840), .B1(n1091), .B2(\mem[2][6] ), 
        .ZN(n1085) );
  INV_X1 U569 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U570 ( .A1(data_in[7]), .A2(n840), .B1(n1091), .B2(\mem[2][7] ), 
        .ZN(n1084) );
  INV_X1 U571 ( .A(n1082), .ZN(n786) );
  AOI22_X1 U572 ( .A1(data_in[0]), .A2(n839), .B1(n1081), .B2(\mem[3][0] ), 
        .ZN(n1082) );
  INV_X1 U573 ( .A(n1080), .ZN(n785) );
  AOI22_X1 U574 ( .A1(data_in[1]), .A2(n839), .B1(n1081), .B2(\mem[3][1] ), 
        .ZN(n1080) );
  INV_X1 U575 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U576 ( .A1(data_in[2]), .A2(n839), .B1(n1081), .B2(\mem[3][2] ), 
        .ZN(n1079) );
  INV_X1 U577 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U578 ( .A1(data_in[3]), .A2(n839), .B1(n1081), .B2(\mem[3][3] ), 
        .ZN(n1078) );
  INV_X1 U579 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U580 ( .A1(data_in[4]), .A2(n839), .B1(n1081), .B2(\mem[3][4] ), 
        .ZN(n1077) );
  INV_X1 U581 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U582 ( .A1(data_in[5]), .A2(n839), .B1(n1081), .B2(\mem[3][5] ), 
        .ZN(n1076) );
  INV_X1 U583 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U584 ( .A1(data_in[6]), .A2(n839), .B1(n1081), .B2(\mem[3][6] ), 
        .ZN(n1075) );
  INV_X1 U585 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U586 ( .A1(data_in[7]), .A2(n839), .B1(n1081), .B2(\mem[3][7] ), 
        .ZN(n1074) );
  INV_X1 U587 ( .A(n1072), .ZN(n778) );
  AOI22_X1 U588 ( .A1(data_in[0]), .A2(n838), .B1(n1071), .B2(\mem[4][0] ), 
        .ZN(n1072) );
  INV_X1 U589 ( .A(n1070), .ZN(n777) );
  AOI22_X1 U590 ( .A1(data_in[1]), .A2(n838), .B1(n1071), .B2(\mem[4][1] ), 
        .ZN(n1070) );
  INV_X1 U591 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U592 ( .A1(data_in[2]), .A2(n838), .B1(n1071), .B2(\mem[4][2] ), 
        .ZN(n1069) );
  INV_X1 U593 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U594 ( .A1(data_in[3]), .A2(n838), .B1(n1071), .B2(\mem[4][3] ), 
        .ZN(n1068) );
  INV_X1 U595 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U596 ( .A1(data_in[4]), .A2(n838), .B1(n1071), .B2(\mem[4][4] ), 
        .ZN(n1067) );
  INV_X1 U597 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U598 ( .A1(data_in[5]), .A2(n838), .B1(n1071), .B2(\mem[4][5] ), 
        .ZN(n1066) );
  INV_X1 U599 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U600 ( .A1(data_in[6]), .A2(n838), .B1(n1071), .B2(\mem[4][6] ), 
        .ZN(n1065) );
  INV_X1 U601 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U602 ( .A1(data_in[7]), .A2(n838), .B1(n1071), .B2(\mem[4][7] ), 
        .ZN(n1064) );
  INV_X1 U603 ( .A(N13), .ZN(n843) );
  INV_X1 U604 ( .A(N14), .ZN(n844) );
  MUX2_X1 U605 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n248), .Z(n2) );
  MUX2_X1 U606 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n248), .Z(n3) );
  MUX2_X1 U607 ( .A(n3), .B(n2), .S(n243), .Z(n4) );
  MUX2_X1 U608 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n248), .Z(n5) );
  MUX2_X1 U609 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n248), .Z(n6) );
  MUX2_X1 U610 ( .A(n6), .B(n5), .S(n243), .Z(n7) );
  MUX2_X1 U611 ( .A(n7), .B(n4), .S(n242), .Z(n8) );
  MUX2_X1 U612 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n248), .Z(n9) );
  MUX2_X1 U613 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n248), .Z(n10) );
  MUX2_X1 U614 ( .A(n10), .B(n9), .S(n243), .Z(n11) );
  MUX2_X1 U615 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n248), .Z(n12) );
  MUX2_X1 U616 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n248), .Z(n13) );
  MUX2_X1 U617 ( .A(n13), .B(n12), .S(n243), .Z(n14) );
  MUX2_X1 U618 ( .A(n14), .B(n11), .S(n242), .Z(n15) );
  MUX2_X1 U619 ( .A(n15), .B(n8), .S(N13), .Z(n16) );
  MUX2_X1 U620 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n246), .Z(n17) );
  MUX2_X1 U621 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n246), .Z(n18) );
  MUX2_X1 U622 ( .A(n18), .B(n17), .S(N11), .Z(n19) );
  MUX2_X1 U623 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n246), .Z(n20) );
  MUX2_X1 U624 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n246), .Z(n21) );
  MUX2_X1 U625 ( .A(n21), .B(n20), .S(N11), .Z(n22) );
  MUX2_X1 U626 ( .A(n22), .B(n19), .S(n242), .Z(n23) );
  MUX2_X1 U627 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n246), .Z(n24) );
  MUX2_X1 U628 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n246), .Z(n25) );
  MUX2_X1 U629 ( .A(n25), .B(n24), .S(N11), .Z(n26) );
  MUX2_X1 U630 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n246), .Z(n27) );
  MUX2_X1 U631 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n246), .Z(n28) );
  MUX2_X1 U632 ( .A(n28), .B(n27), .S(n244), .Z(n29) );
  MUX2_X1 U633 ( .A(n29), .B(n26), .S(n242), .Z(n30) );
  MUX2_X1 U634 ( .A(n30), .B(n23), .S(N13), .Z(n31) );
  MUX2_X1 U635 ( .A(n31), .B(n16), .S(N14), .Z(N22) );
  MUX2_X1 U636 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n246), .Z(n32) );
  MUX2_X1 U637 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n246), .Z(n33) );
  MUX2_X1 U638 ( .A(n33), .B(n32), .S(n244), .Z(n34) );
  MUX2_X1 U639 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n246), .Z(n35) );
  MUX2_X1 U640 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n246), .Z(n36) );
  MUX2_X1 U641 ( .A(n36), .B(n35), .S(N11), .Z(n37) );
  MUX2_X1 U642 ( .A(n37), .B(n34), .S(n242), .Z(n38) );
  MUX2_X1 U643 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n247), .Z(n39) );
  MUX2_X1 U644 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n247), .Z(n40) );
  MUX2_X1 U645 ( .A(n40), .B(n39), .S(N11), .Z(n41) );
  MUX2_X1 U646 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n247), .Z(n42) );
  MUX2_X1 U647 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n247), .Z(n43) );
  MUX2_X1 U648 ( .A(n43), .B(n42), .S(n245), .Z(n44) );
  MUX2_X1 U649 ( .A(n44), .B(n41), .S(N12), .Z(n45) );
  MUX2_X1 U650 ( .A(n45), .B(n38), .S(N13), .Z(n46) );
  MUX2_X1 U651 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n247), .Z(n47) );
  MUX2_X1 U652 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n247), .Z(n48) );
  MUX2_X1 U653 ( .A(n48), .B(n47), .S(N11), .Z(n49) );
  MUX2_X1 U654 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n247), .Z(n50) );
  MUX2_X1 U655 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n247), .Z(n51) );
  MUX2_X1 U656 ( .A(n51), .B(n50), .S(n244), .Z(n52) );
  MUX2_X1 U657 ( .A(n52), .B(n49), .S(N12), .Z(n53) );
  MUX2_X1 U658 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n247), .Z(n54) );
  MUX2_X1 U659 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n247), .Z(n55) );
  MUX2_X1 U660 ( .A(n55), .B(n54), .S(N11), .Z(n56) );
  MUX2_X1 U661 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n247), .Z(n57) );
  MUX2_X1 U662 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n247), .Z(n58) );
  MUX2_X1 U663 ( .A(n58), .B(n57), .S(n245), .Z(n59) );
  MUX2_X1 U664 ( .A(n59), .B(n56), .S(N12), .Z(n60) );
  MUX2_X1 U665 ( .A(n60), .B(n53), .S(N13), .Z(n61) );
  MUX2_X1 U666 ( .A(n61), .B(n46), .S(N14), .Z(N21) );
  MUX2_X1 U667 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n246), .Z(n62) );
  MUX2_X1 U668 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n250), .Z(n63) );
  MUX2_X1 U669 ( .A(n63), .B(n62), .S(n245), .Z(n64) );
  MUX2_X1 U670 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n249), .Z(n65) );
  MUX2_X1 U671 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n250), .Z(n66) );
  MUX2_X1 U672 ( .A(n66), .B(n65), .S(N11), .Z(n67) );
  MUX2_X1 U673 ( .A(n67), .B(n64), .S(n242), .Z(n68) );
  MUX2_X1 U674 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n247), .Z(n69) );
  MUX2_X1 U675 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n246), .Z(n70) );
  MUX2_X1 U676 ( .A(n70), .B(n69), .S(n243), .Z(n71) );
  MUX2_X1 U677 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n249), .Z(n72) );
  MUX2_X1 U678 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n250), .Z(n73) );
  MUX2_X1 U679 ( .A(n73), .B(n72), .S(N11), .Z(n74) );
  MUX2_X1 U680 ( .A(n74), .B(n71), .S(n242), .Z(n75) );
  MUX2_X1 U681 ( .A(n75), .B(n68), .S(N13), .Z(n76) );
  MUX2_X1 U682 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n249), .Z(n77) );
  MUX2_X1 U683 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n247), .Z(n78) );
  MUX2_X1 U684 ( .A(n78), .B(n77), .S(n245), .Z(n79) );
  MUX2_X1 U685 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n246), .Z(n80) );
  MUX2_X1 U686 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n249), .Z(n81) );
  MUX2_X1 U687 ( .A(n81), .B(n80), .S(N11), .Z(n82) );
  MUX2_X1 U688 ( .A(n82), .B(n79), .S(n242), .Z(n83) );
  MUX2_X1 U689 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n251), .Z(n84) );
  MUX2_X1 U690 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n247), .Z(n85) );
  MUX2_X1 U691 ( .A(n85), .B(n84), .S(n243), .Z(n86) );
  MUX2_X1 U692 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n246), .Z(n87) );
  MUX2_X1 U693 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n247), .Z(n88) );
  MUX2_X1 U694 ( .A(n88), .B(n87), .S(N11), .Z(n89) );
  MUX2_X1 U695 ( .A(n89), .B(n86), .S(n242), .Z(n90) );
  MUX2_X1 U696 ( .A(n90), .B(n83), .S(N13), .Z(n91) );
  MUX2_X1 U697 ( .A(n91), .B(n76), .S(N14), .Z(N20) );
  MUX2_X1 U698 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n250), .Z(n92) );
  MUX2_X1 U699 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n251), .Z(n93) );
  MUX2_X1 U700 ( .A(n93), .B(n92), .S(n244), .Z(n94) );
  MUX2_X1 U701 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n249), .Z(n95) );
  MUX2_X1 U702 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n247), .Z(n96) );
  MUX2_X1 U703 ( .A(n96), .B(n95), .S(n244), .Z(n97) );
  MUX2_X1 U704 ( .A(n97), .B(n94), .S(n242), .Z(n98) );
  MUX2_X1 U705 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n251), .Z(n99) );
  MUX2_X1 U706 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n249), .Z(n100) );
  MUX2_X1 U707 ( .A(n100), .B(n99), .S(n245), .Z(n101) );
  MUX2_X1 U708 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n251), .Z(n102) );
  MUX2_X1 U709 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n250), .Z(n103) );
  MUX2_X1 U710 ( .A(n103), .B(n102), .S(N11), .Z(n104) );
  MUX2_X1 U711 ( .A(n104), .B(n101), .S(n242), .Z(n105) );
  MUX2_X1 U712 ( .A(n105), .B(n98), .S(N13), .Z(n106) );
  MUX2_X1 U713 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n248), .Z(n107) );
  MUX2_X1 U714 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n248), .Z(n108) );
  MUX2_X1 U715 ( .A(n108), .B(n107), .S(n243), .Z(n109) );
  MUX2_X1 U716 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n248), .Z(n110) );
  MUX2_X1 U717 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n248), .Z(n111) );
  MUX2_X1 U718 ( .A(n111), .B(n110), .S(n244), .Z(n112) );
  MUX2_X1 U719 ( .A(n112), .B(n109), .S(n242), .Z(n113) );
  MUX2_X1 U720 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n248), .Z(n114) );
  MUX2_X1 U721 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n248), .Z(n115) );
  MUX2_X1 U722 ( .A(n115), .B(n114), .S(n243), .Z(n116) );
  MUX2_X1 U723 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n248), .Z(n117) );
  MUX2_X1 U724 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n248), .Z(n118) );
  MUX2_X1 U725 ( .A(n118), .B(n117), .S(N11), .Z(n119) );
  MUX2_X1 U726 ( .A(n119), .B(n116), .S(n242), .Z(n120) );
  MUX2_X1 U727 ( .A(n120), .B(n113), .S(N13), .Z(n121) );
  MUX2_X1 U728 ( .A(n121), .B(n106), .S(N14), .Z(N19) );
  MUX2_X1 U729 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n248), .Z(n122) );
  MUX2_X1 U730 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n248), .Z(n123) );
  MUX2_X1 U731 ( .A(n123), .B(n122), .S(n243), .Z(n124) );
  MUX2_X1 U732 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n248), .Z(n125) );
  MUX2_X1 U733 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n248), .Z(n126) );
  MUX2_X1 U734 ( .A(n126), .B(n125), .S(n243), .Z(n127) );
  MUX2_X1 U735 ( .A(n127), .B(n124), .S(n242), .Z(n128) );
  MUX2_X1 U736 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n249), .Z(n129) );
  MUX2_X1 U737 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n249), .Z(n130) );
  MUX2_X1 U738 ( .A(n130), .B(n129), .S(n243), .Z(n131) );
  MUX2_X1 U739 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n249), .Z(n132) );
  MUX2_X1 U740 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n249), .Z(n133) );
  MUX2_X1 U741 ( .A(n133), .B(n132), .S(n243), .Z(n134) );
  MUX2_X1 U742 ( .A(n134), .B(n131), .S(n242), .Z(n135) );
  MUX2_X1 U743 ( .A(n135), .B(n128), .S(N13), .Z(n136) );
  MUX2_X1 U744 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n249), .Z(n137) );
  MUX2_X1 U745 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n249), .Z(n138) );
  MUX2_X1 U746 ( .A(n138), .B(n137), .S(n243), .Z(n139) );
  MUX2_X1 U747 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n249), .Z(n140) );
  MUX2_X1 U748 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n249), .Z(n141) );
  MUX2_X1 U749 ( .A(n141), .B(n140), .S(n245), .Z(n142) );
  MUX2_X1 U750 ( .A(n142), .B(n139), .S(n242), .Z(n143) );
  MUX2_X1 U751 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n249), .Z(n144) );
  MUX2_X1 U752 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n249), .Z(n145) );
  MUX2_X1 U753 ( .A(n145), .B(n144), .S(n243), .Z(n146) );
  MUX2_X1 U754 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n249), .Z(n147) );
  MUX2_X1 U755 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n249), .Z(n148) );
  MUX2_X1 U756 ( .A(n148), .B(n147), .S(n243), .Z(n149) );
  MUX2_X1 U757 ( .A(n149), .B(n146), .S(n242), .Z(n150) );
  MUX2_X1 U758 ( .A(n150), .B(n143), .S(N13), .Z(n151) );
  MUX2_X1 U759 ( .A(n151), .B(n136), .S(N14), .Z(N18) );
  MUX2_X1 U760 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n250), .Z(n152) );
  MUX2_X1 U761 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n250), .Z(n153) );
  MUX2_X1 U762 ( .A(n153), .B(n152), .S(n244), .Z(n154) );
  MUX2_X1 U763 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n250), .Z(n155) );
  MUX2_X1 U764 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n250), .Z(n156) );
  MUX2_X1 U765 ( .A(n156), .B(n155), .S(n244), .Z(n157) );
  MUX2_X1 U766 ( .A(n157), .B(n154), .S(n242), .Z(n158) );
  MUX2_X1 U767 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n250), .Z(n159) );
  MUX2_X1 U768 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n250), .Z(n160) );
  MUX2_X1 U769 ( .A(n160), .B(n159), .S(n244), .Z(n161) );
  MUX2_X1 U770 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n250), .Z(n162) );
  MUX2_X1 U771 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n250), .Z(n163) );
  MUX2_X1 U772 ( .A(n163), .B(n162), .S(n244), .Z(n164) );
  MUX2_X1 U773 ( .A(n164), .B(n161), .S(N12), .Z(n165) );
  MUX2_X1 U774 ( .A(n165), .B(n158), .S(N13), .Z(n166) );
  MUX2_X1 U775 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n250), .Z(n167) );
  MUX2_X1 U776 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n250), .Z(n168) );
  MUX2_X1 U777 ( .A(n168), .B(n167), .S(n244), .Z(n169) );
  MUX2_X1 U778 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n250), .Z(n170) );
  MUX2_X1 U779 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n250), .Z(n171) );
  MUX2_X1 U780 ( .A(n171), .B(n170), .S(n244), .Z(n172) );
  MUX2_X1 U781 ( .A(n172), .B(n169), .S(n242), .Z(n173) );
  MUX2_X1 U782 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n251), .Z(n174) );
  MUX2_X1 U783 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n251), .Z(n175) );
  MUX2_X1 U784 ( .A(n175), .B(n174), .S(n244), .Z(n176) );
  MUX2_X1 U785 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n251), .Z(n177) );
  MUX2_X1 U786 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n251), .Z(n178) );
  MUX2_X1 U787 ( .A(n178), .B(n177), .S(n244), .Z(n179) );
  MUX2_X1 U788 ( .A(n179), .B(n176), .S(N12), .Z(n180) );
  MUX2_X1 U789 ( .A(n180), .B(n173), .S(N13), .Z(n181) );
  MUX2_X1 U790 ( .A(n181), .B(n166), .S(N14), .Z(N17) );
  MUX2_X1 U791 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n246), .Z(n182) );
  MUX2_X1 U792 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n251), .Z(n183) );
  MUX2_X1 U793 ( .A(n183), .B(n182), .S(n244), .Z(n184) );
  MUX2_X1 U794 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n251), .Z(n185) );
  MUX2_X1 U795 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n251), .Z(n186) );
  MUX2_X1 U796 ( .A(n186), .B(n185), .S(n244), .Z(n187) );
  MUX2_X1 U797 ( .A(n187), .B(n184), .S(n242), .Z(n188) );
  MUX2_X1 U798 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n251), .Z(n189) );
  MUX2_X1 U799 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n251), .Z(n190) );
  MUX2_X1 U800 ( .A(n190), .B(n189), .S(n244), .Z(n191) );
  MUX2_X1 U801 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n247), .Z(n192) );
  MUX2_X1 U802 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n251), .Z(n193) );
  MUX2_X1 U803 ( .A(n193), .B(n192), .S(n244), .Z(n194) );
  MUX2_X1 U804 ( .A(n194), .B(n191), .S(N12), .Z(n195) );
  MUX2_X1 U805 ( .A(n195), .B(n188), .S(N13), .Z(n196) );
  MUX2_X1 U806 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n251), .Z(n197) );
  MUX2_X1 U807 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(N10), .Z(n198) );
  MUX2_X1 U808 ( .A(n198), .B(n197), .S(n245), .Z(n199) );
  MUX2_X1 U809 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(N10), .Z(n200) );
  MUX2_X1 U810 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n251), .Z(n201) );
  MUX2_X1 U811 ( .A(n201), .B(n200), .S(n245), .Z(n202) );
  MUX2_X1 U812 ( .A(n202), .B(n199), .S(n242), .Z(n203) );
  MUX2_X1 U813 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(N10), .Z(n204) );
  MUX2_X1 U814 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n251), .Z(n205) );
  MUX2_X1 U815 ( .A(n205), .B(n204), .S(n245), .Z(n206) );
  MUX2_X1 U816 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n207) );
  MUX2_X1 U817 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n251), .Z(n208) );
  MUX2_X1 U818 ( .A(n208), .B(n207), .S(n245), .Z(n209) );
  MUX2_X1 U819 ( .A(n209), .B(n206), .S(N12), .Z(n210) );
  MUX2_X1 U820 ( .A(n210), .B(n203), .S(N13), .Z(n211) );
  MUX2_X1 U821 ( .A(n211), .B(n196), .S(N14), .Z(N16) );
  MUX2_X1 U822 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n250), .Z(n212) );
  MUX2_X1 U823 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(N10), .Z(n213) );
  MUX2_X1 U824 ( .A(n213), .B(n212), .S(n245), .Z(n214) );
  MUX2_X1 U825 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(N10), .Z(n215) );
  MUX2_X1 U826 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(N10), .Z(n216) );
  MUX2_X1 U827 ( .A(n216), .B(n215), .S(n245), .Z(n217) );
  MUX2_X1 U828 ( .A(n217), .B(n214), .S(n242), .Z(n218) );
  MUX2_X1 U829 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n248), .Z(n219) );
  MUX2_X1 U830 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(N10), .Z(n220) );
  MUX2_X1 U831 ( .A(n220), .B(n219), .S(n245), .Z(n221) );
  MUX2_X1 U832 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n251), .Z(n222) );
  MUX2_X1 U833 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n223) );
  MUX2_X1 U834 ( .A(n223), .B(n222), .S(n245), .Z(n224) );
  MUX2_X1 U835 ( .A(n224), .B(n221), .S(N12), .Z(n225) );
  MUX2_X1 U836 ( .A(n225), .B(n218), .S(N13), .Z(n226) );
  MUX2_X1 U837 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n248), .Z(n227) );
  MUX2_X1 U838 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n251), .Z(n228) );
  MUX2_X1 U839 ( .A(n228), .B(n227), .S(n245), .Z(n229) );
  MUX2_X1 U840 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n248), .Z(n230) );
  MUX2_X1 U841 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n231) );
  MUX2_X1 U842 ( .A(n231), .B(n230), .S(n245), .Z(n232) );
  MUX2_X1 U843 ( .A(n232), .B(n229), .S(n242), .Z(n233) );
  MUX2_X1 U844 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n234) );
  MUX2_X1 U845 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n235) );
  MUX2_X1 U846 ( .A(n235), .B(n234), .S(n245), .Z(n236) );
  MUX2_X1 U847 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n237) );
  MUX2_X1 U848 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n238) );
  MUX2_X1 U849 ( .A(n238), .B(n237), .S(n245), .Z(n239) );
  MUX2_X1 U850 ( .A(n239), .B(n236), .S(N12), .Z(n240) );
  MUX2_X1 U851 ( .A(n240), .B(n233), .S(N13), .Z(n241) );
  MUX2_X1 U852 ( .A(n241), .B(n226), .S(N14), .Z(N15) );
  CLKBUF_X1 U853 ( .A(N11), .Z(n243) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_13 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  BUF_X1 U3 ( .A(n250), .Z(n246) );
  BUF_X1 U4 ( .A(n250), .Z(n247) );
  BUF_X1 U5 ( .A(n250), .Z(n248) );
  BUF_X1 U6 ( .A(n250), .Z(n249) );
  BUF_X1 U7 ( .A(N10), .Z(n250) );
  INV_X1 U8 ( .A(n1111), .ZN(n841) );
  INV_X1 U9 ( .A(n1100), .ZN(n840) );
  INV_X1 U10 ( .A(n1090), .ZN(n839) );
  INV_X1 U11 ( .A(n1080), .ZN(n838) );
  INV_X1 U12 ( .A(n1070), .ZN(n837) );
  INV_X1 U13 ( .A(n1060), .ZN(n836) );
  INV_X1 U14 ( .A(n1051), .ZN(n835) );
  INV_X1 U15 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U16 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U18 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U19 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U20 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U21 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U22 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U23 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U24 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U26 ( .A(n1131), .ZN(n816) );
  INV_X1 U27 ( .A(n1121), .ZN(n815) );
  INV_X1 U28 ( .A(n887), .ZN(n814) );
  INV_X1 U29 ( .A(n878), .ZN(n813) );
  INV_X1 U30 ( .A(n869), .ZN(n812) );
  INV_X1 U31 ( .A(n860), .ZN(n811) );
  INV_X1 U32 ( .A(n851), .ZN(n810) );
  INV_X1 U33 ( .A(n987), .ZN(n828) );
  INV_X1 U34 ( .A(n978), .ZN(n827) );
  INV_X1 U35 ( .A(n969), .ZN(n826) );
  INV_X1 U36 ( .A(n914), .ZN(n820) );
  INV_X1 U37 ( .A(n905), .ZN(n819) );
  INV_X1 U38 ( .A(n896), .ZN(n818) );
  INV_X1 U39 ( .A(n1033), .ZN(n833) );
  INV_X1 U40 ( .A(n1023), .ZN(n832) );
  INV_X1 U41 ( .A(n1014), .ZN(n831) );
  INV_X1 U42 ( .A(n1005), .ZN(n830) );
  INV_X1 U43 ( .A(n996), .ZN(n829) );
  INV_X1 U44 ( .A(n960), .ZN(n825) );
  INV_X1 U45 ( .A(n950), .ZN(n824) );
  INV_X1 U46 ( .A(n941), .ZN(n823) );
  INV_X1 U47 ( .A(n932), .ZN(n822) );
  INV_X1 U48 ( .A(n923), .ZN(n821) );
  INV_X1 U49 ( .A(n1142), .ZN(n817) );
  BUF_X1 U50 ( .A(N11), .Z(n243) );
  BUF_X1 U51 ( .A(N11), .Z(n244) );
  INV_X1 U52 ( .A(N10), .ZN(n251) );
  BUF_X1 U53 ( .A(N12), .Z(n241) );
  NOR3_X1 U54 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U55 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U56 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U57 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U58 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U59 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U60 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U61 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U62 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U63 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U64 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U65 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U66 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U67 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U68 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U69 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U70 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U71 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U72 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U73 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U74 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U75 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U76 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U77 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U78 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U79 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U80 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U81 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U82 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U83 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U84 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U85 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U86 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U87 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U88 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U89 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U90 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U91 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U92 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U93 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U94 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U95 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U96 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U97 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U98 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U99 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U100 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U101 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U102 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U103 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U104 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U105 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U106 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U107 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U108 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U109 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U110 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U111 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U112 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U113 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U114 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U115 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U116 ( .A(n988), .ZN(n705) );
  AOI22_X1 U117 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U118 ( .A(n986), .ZN(n704) );
  AOI22_X1 U119 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U120 ( .A(n985), .ZN(n703) );
  AOI22_X1 U121 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U122 ( .A(n983), .ZN(n701) );
  AOI22_X1 U123 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U124 ( .A(n982), .ZN(n700) );
  AOI22_X1 U125 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U126 ( .A(n981), .ZN(n699) );
  AOI22_X1 U127 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U128 ( .A(n980), .ZN(n698) );
  AOI22_X1 U129 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U130 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U131 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U132 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U133 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U134 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U135 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U136 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U137 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U138 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U139 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U140 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U141 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U142 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U143 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U144 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U145 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U146 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U147 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U148 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U149 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U150 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U151 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U152 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U153 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U154 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U155 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U156 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U157 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U158 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U159 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U160 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U161 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U162 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U163 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U164 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U165 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U166 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U167 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U168 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U169 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U170 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U171 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U172 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U173 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U174 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U175 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U176 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U177 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U178 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U179 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U180 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U181 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U182 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U183 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U184 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U185 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U186 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U187 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U188 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U189 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U190 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U191 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U192 ( .A(n999), .ZN(n715) );
  AOI22_X1 U193 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U194 ( .A(n998), .ZN(n714) );
  AOI22_X1 U195 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U196 ( .A(n951), .ZN(n673) );
  AOI22_X1 U197 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U198 ( .A(n949), .ZN(n672) );
  AOI22_X1 U199 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U200 ( .A(n948), .ZN(n671) );
  AOI22_X1 U201 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U202 ( .A(n947), .ZN(n670) );
  AOI22_X1 U203 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U204 ( .A(n946), .ZN(n669) );
  AOI22_X1 U205 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U206 ( .A(n913), .ZN(n640) );
  AOI22_X1 U207 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U208 ( .A(n912), .ZN(n639) );
  AOI22_X1 U209 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U210 ( .A(n911), .ZN(n638) );
  AOI22_X1 U211 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U212 ( .A(n910), .ZN(n637) );
  AOI22_X1 U213 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U214 ( .A(n909), .ZN(n636) );
  AOI22_X1 U215 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U216 ( .A(n908), .ZN(n635) );
  AOI22_X1 U217 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U218 ( .A(n907), .ZN(n634) );
  AOI22_X1 U219 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U220 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U221 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U222 ( .A(n984), .ZN(n702) );
  AOI22_X1 U223 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U224 ( .A(n915), .ZN(n641) );
  AOI22_X1 U225 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U226 ( .A(n945), .ZN(n668) );
  AOI22_X1 U227 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U228 ( .A(n944), .ZN(n667) );
  AOI22_X1 U229 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U230 ( .A(n943), .ZN(n666) );
  AOI22_X1 U231 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U232 ( .A(n979), .ZN(n697) );
  AOI22_X1 U233 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U234 ( .A(n977), .ZN(n696) );
  AOI22_X1 U235 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U236 ( .A(n976), .ZN(n695) );
  AOI22_X1 U237 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U238 ( .A(n975), .ZN(n694) );
  AOI22_X1 U239 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U240 ( .A(n974), .ZN(n693) );
  AOI22_X1 U241 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U242 ( .A(n973), .ZN(n692) );
  AOI22_X1 U243 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U244 ( .A(n972), .ZN(n691) );
  AOI22_X1 U245 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U246 ( .A(n971), .ZN(n690) );
  AOI22_X1 U247 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U248 ( .A(n970), .ZN(n689) );
  AOI22_X1 U249 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U250 ( .A(n968), .ZN(n688) );
  AOI22_X1 U251 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U252 ( .A(n967), .ZN(n687) );
  AOI22_X1 U253 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U254 ( .A(n966), .ZN(n686) );
  AOI22_X1 U255 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U256 ( .A(n965), .ZN(n685) );
  AOI22_X1 U257 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U258 ( .A(n964), .ZN(n684) );
  AOI22_X1 U259 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U260 ( .A(n963), .ZN(n683) );
  AOI22_X1 U261 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U262 ( .A(n962), .ZN(n682) );
  AOI22_X1 U263 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U264 ( .A(n942), .ZN(n665) );
  AOI22_X1 U265 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U266 ( .A(n940), .ZN(n664) );
  AOI22_X1 U267 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U268 ( .A(n939), .ZN(n663) );
  AOI22_X1 U269 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U270 ( .A(n938), .ZN(n662) );
  AOI22_X1 U271 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U272 ( .A(n937), .ZN(n661) );
  AOI22_X1 U273 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U274 ( .A(n936), .ZN(n660) );
  AOI22_X1 U275 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U276 ( .A(n935), .ZN(n659) );
  AOI22_X1 U277 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U278 ( .A(n934), .ZN(n658) );
  AOI22_X1 U279 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U280 ( .A(n933), .ZN(n657) );
  AOI22_X1 U281 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U282 ( .A(n931), .ZN(n656) );
  AOI22_X1 U283 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U284 ( .A(n930), .ZN(n655) );
  AOI22_X1 U285 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U286 ( .A(n929), .ZN(n654) );
  AOI22_X1 U287 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U288 ( .A(n928), .ZN(n653) );
  AOI22_X1 U289 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U290 ( .A(n927), .ZN(n652) );
  AOI22_X1 U291 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U292 ( .A(n926), .ZN(n651) );
  AOI22_X1 U293 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U294 ( .A(n925), .ZN(n650) );
  AOI22_X1 U295 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U296 ( .A(n906), .ZN(n633) );
  AOI22_X1 U297 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U298 ( .A(n904), .ZN(n632) );
  AOI22_X1 U299 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U300 ( .A(n903), .ZN(n631) );
  AOI22_X1 U301 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U302 ( .A(n902), .ZN(n630) );
  AOI22_X1 U303 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U304 ( .A(n901), .ZN(n629) );
  AOI22_X1 U305 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U306 ( .A(n900), .ZN(n628) );
  AOI22_X1 U307 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U308 ( .A(n899), .ZN(n627) );
  AOI22_X1 U309 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U310 ( .A(n898), .ZN(n626) );
  AOI22_X1 U311 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U312 ( .A(n897), .ZN(n625) );
  AOI22_X1 U313 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U314 ( .A(n895), .ZN(n624) );
  AOI22_X1 U315 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U316 ( .A(n894), .ZN(n623) );
  AOI22_X1 U317 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U318 ( .A(n893), .ZN(n622) );
  AOI22_X1 U319 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U320 ( .A(n892), .ZN(n621) );
  AOI22_X1 U321 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U322 ( .A(n891), .ZN(n620) );
  AOI22_X1 U323 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U324 ( .A(n890), .ZN(n619) );
  AOI22_X1 U325 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U326 ( .A(n889), .ZN(n618) );
  AOI22_X1 U327 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U328 ( .A(N12), .ZN(n253) );
  INV_X1 U329 ( .A(N11), .ZN(n252) );
  INV_X1 U330 ( .A(n997), .ZN(n713) );
  AOI22_X1 U331 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U332 ( .A(n995), .ZN(n712) );
  AOI22_X1 U333 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U334 ( .A(n994), .ZN(n711) );
  AOI22_X1 U335 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U336 ( .A(n993), .ZN(n710) );
  AOI22_X1 U337 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U338 ( .A(n992), .ZN(n709) );
  AOI22_X1 U339 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U340 ( .A(n991), .ZN(n708) );
  AOI22_X1 U341 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U342 ( .A(n990), .ZN(n707) );
  AOI22_X1 U343 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U344 ( .A(n989), .ZN(n706) );
  AOI22_X1 U345 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U346 ( .A(n924), .ZN(n649) );
  AOI22_X1 U347 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U348 ( .A(n922), .ZN(n648) );
  AOI22_X1 U349 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U350 ( .A(n921), .ZN(n647) );
  AOI22_X1 U351 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U352 ( .A(n920), .ZN(n646) );
  AOI22_X1 U353 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U354 ( .A(n919), .ZN(n645) );
  AOI22_X1 U355 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U356 ( .A(n918), .ZN(n644) );
  AOI22_X1 U357 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U358 ( .A(n917), .ZN(n643) );
  AOI22_X1 U359 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U360 ( .A(n916), .ZN(n642) );
  AOI22_X1 U361 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U362 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U363 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U364 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U365 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U366 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U367 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U368 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U369 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U370 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U371 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U372 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U373 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U374 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U375 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U376 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U377 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U378 ( .A(n961), .ZN(n681) );
  AOI22_X1 U379 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U380 ( .A(n959), .ZN(n680) );
  AOI22_X1 U381 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U382 ( .A(n958), .ZN(n679) );
  AOI22_X1 U383 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U384 ( .A(n957), .ZN(n678) );
  AOI22_X1 U385 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U386 ( .A(n956), .ZN(n677) );
  AOI22_X1 U387 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U388 ( .A(n955), .ZN(n676) );
  AOI22_X1 U389 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U390 ( .A(n954), .ZN(n675) );
  AOI22_X1 U391 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U392 ( .A(n953), .ZN(n674) );
  AOI22_X1 U393 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U394 ( .A(n888), .ZN(n617) );
  AOI22_X1 U395 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U396 ( .A(n886), .ZN(n616) );
  AOI22_X1 U397 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U398 ( .A(n885), .ZN(n615) );
  AOI22_X1 U399 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U400 ( .A(n884), .ZN(n614) );
  AOI22_X1 U401 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U402 ( .A(n883), .ZN(n613) );
  AOI22_X1 U403 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U404 ( .A(n882), .ZN(n612) );
  AOI22_X1 U405 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U406 ( .A(n881), .ZN(n611) );
  AOI22_X1 U407 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U408 ( .A(n880), .ZN(n610) );
  AOI22_X1 U409 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U410 ( .A(n879), .ZN(n609) );
  AOI22_X1 U411 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U412 ( .A(n877), .ZN(n608) );
  AOI22_X1 U413 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U414 ( .A(n876), .ZN(n607) );
  AOI22_X1 U415 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U416 ( .A(n875), .ZN(n606) );
  AOI22_X1 U417 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U418 ( .A(n874), .ZN(n605) );
  AOI22_X1 U419 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U420 ( .A(n873), .ZN(n604) );
  AOI22_X1 U421 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U422 ( .A(n872), .ZN(n603) );
  AOI22_X1 U423 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U424 ( .A(n871), .ZN(n602) );
  AOI22_X1 U425 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U426 ( .A(n870), .ZN(n601) );
  AOI22_X1 U427 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U428 ( .A(n868), .ZN(n600) );
  AOI22_X1 U429 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U430 ( .A(n867), .ZN(n599) );
  AOI22_X1 U431 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U432 ( .A(n866), .ZN(n598) );
  AOI22_X1 U433 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U434 ( .A(n865), .ZN(n597) );
  AOI22_X1 U435 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U436 ( .A(n864), .ZN(n596) );
  AOI22_X1 U437 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U438 ( .A(n863), .ZN(n595) );
  AOI22_X1 U439 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U440 ( .A(n862), .ZN(n594) );
  AOI22_X1 U441 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U442 ( .A(n861), .ZN(n293) );
  AOI22_X1 U443 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U444 ( .A(n859), .ZN(n292) );
  AOI22_X1 U445 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U446 ( .A(n858), .ZN(n291) );
  AOI22_X1 U447 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U448 ( .A(n857), .ZN(n290) );
  AOI22_X1 U449 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U450 ( .A(n856), .ZN(n289) );
  AOI22_X1 U451 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U452 ( .A(n855), .ZN(n288) );
  AOI22_X1 U453 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U454 ( .A(n854), .ZN(n287) );
  AOI22_X1 U455 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U456 ( .A(n853), .ZN(n286) );
  AOI22_X1 U457 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U458 ( .A(n852), .ZN(n285) );
  AOI22_X1 U459 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U460 ( .A(n850), .ZN(n284) );
  AOI22_X1 U461 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U462 ( .A(n849), .ZN(n283) );
  AOI22_X1 U463 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U464 ( .A(n848), .ZN(n282) );
  AOI22_X1 U465 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U466 ( .A(n847), .ZN(n281) );
  AOI22_X1 U467 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U468 ( .A(n846), .ZN(n280) );
  AOI22_X1 U469 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U470 ( .A(n845), .ZN(n279) );
  AOI22_X1 U471 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U472 ( .A(n844), .ZN(n278) );
  AOI22_X1 U473 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U474 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U475 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U476 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U477 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U478 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U479 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U480 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U481 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U482 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U483 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U484 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U485 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U486 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U487 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U488 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U489 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U490 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U491 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U492 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U493 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U494 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U495 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U496 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U497 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U498 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U499 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U500 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U501 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U502 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U503 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U504 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U505 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U506 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U507 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U508 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U509 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U510 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U511 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U512 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U513 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U514 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U515 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U516 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U517 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U518 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U519 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U520 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U521 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U522 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U523 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U524 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U525 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U526 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U527 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U528 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U529 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U530 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U531 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U532 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U533 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U534 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U535 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U536 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U537 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U538 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U539 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U540 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U541 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U542 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U543 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U544 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U545 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U546 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U547 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U548 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U549 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U550 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U551 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U552 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U553 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U554 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U555 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U556 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U557 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U558 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U559 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U560 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U561 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U562 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U563 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U564 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U565 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U566 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U567 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U568 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U569 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U570 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U571 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U572 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U573 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U574 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U575 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U576 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U577 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U578 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U579 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U580 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U581 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U582 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U583 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U584 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U585 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U586 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U587 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U588 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U589 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U590 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U591 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U592 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U593 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U594 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U595 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U596 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U597 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U598 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U599 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U600 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U601 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U602 ( .A(N13), .ZN(n842) );
  INV_X1 U603 ( .A(N14), .ZN(n843) );
  MUX2_X1 U604 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n245), .Z(n1) );
  MUX2_X1 U605 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n245), .Z(n2) );
  MUX2_X1 U606 ( .A(n2), .B(n1), .S(n242), .Z(n3) );
  MUX2_X1 U607 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n245), .Z(n4) );
  MUX2_X1 U608 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n245), .Z(n5) );
  MUX2_X1 U609 ( .A(n5), .B(n4), .S(n242), .Z(n6) );
  MUX2_X1 U610 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U611 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n245), .Z(n8) );
  MUX2_X1 U612 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n245), .Z(n9) );
  MUX2_X1 U613 ( .A(n9), .B(n8), .S(n242), .Z(n10) );
  MUX2_X1 U614 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n245), .Z(n11) );
  MUX2_X1 U615 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n245), .Z(n12) );
  MUX2_X1 U616 ( .A(n12), .B(n11), .S(n242), .Z(n13) );
  MUX2_X1 U617 ( .A(n13), .B(n10), .S(n241), .Z(n14) );
  MUX2_X1 U618 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U619 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n246), .Z(n16) );
  MUX2_X1 U620 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n246), .Z(n17) );
  MUX2_X1 U621 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U622 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n246), .Z(n19) );
  MUX2_X1 U623 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n246), .Z(n20) );
  MUX2_X1 U624 ( .A(n20), .B(n19), .S(n242), .Z(n21) );
  MUX2_X1 U625 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U626 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n246), .Z(n23) );
  MUX2_X1 U627 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n246), .Z(n24) );
  MUX2_X1 U628 ( .A(n24), .B(n23), .S(n244), .Z(n25) );
  MUX2_X1 U629 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n246), .Z(n26) );
  MUX2_X1 U630 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n246), .Z(n27) );
  MUX2_X1 U631 ( .A(n27), .B(n26), .S(n244), .Z(n28) );
  MUX2_X1 U632 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U633 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U634 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U635 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n246), .Z(n31) );
  MUX2_X1 U636 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n246), .Z(n32) );
  MUX2_X1 U637 ( .A(n32), .B(n31), .S(N11), .Z(n33) );
  MUX2_X1 U638 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n246), .Z(n34) );
  MUX2_X1 U639 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n246), .Z(n35) );
  MUX2_X1 U640 ( .A(n35), .B(n34), .S(N11), .Z(n36) );
  MUX2_X1 U641 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U642 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n247), .Z(n38) );
  MUX2_X1 U643 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n247), .Z(n39) );
  MUX2_X1 U644 ( .A(n39), .B(n38), .S(N11), .Z(n40) );
  MUX2_X1 U645 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n247), .Z(n41) );
  MUX2_X1 U646 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n247), .Z(n42) );
  MUX2_X1 U647 ( .A(n42), .B(n41), .S(n242), .Z(n43) );
  MUX2_X1 U648 ( .A(n43), .B(n40), .S(n241), .Z(n44) );
  MUX2_X1 U649 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U650 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n247), .Z(n46) );
  MUX2_X1 U651 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n247), .Z(n47) );
  MUX2_X1 U652 ( .A(n47), .B(n46), .S(N11), .Z(n48) );
  MUX2_X1 U653 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n247), .Z(n49) );
  MUX2_X1 U654 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n247), .Z(n50) );
  MUX2_X1 U655 ( .A(n50), .B(n49), .S(n244), .Z(n51) );
  MUX2_X1 U656 ( .A(n51), .B(n48), .S(n241), .Z(n52) );
  MUX2_X1 U657 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n247), .Z(n53) );
  MUX2_X1 U658 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n247), .Z(n54) );
  MUX2_X1 U659 ( .A(n54), .B(n53), .S(n243), .Z(n55) );
  MUX2_X1 U660 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n247), .Z(n56) );
  MUX2_X1 U661 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n247), .Z(n57) );
  MUX2_X1 U662 ( .A(n57), .B(n56), .S(n243), .Z(n58) );
  MUX2_X1 U663 ( .A(n58), .B(n55), .S(n241), .Z(n59) );
  MUX2_X1 U664 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U665 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U666 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n248), .Z(n61) );
  MUX2_X1 U667 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n248), .Z(n62) );
  MUX2_X1 U668 ( .A(n62), .B(n61), .S(n244), .Z(n63) );
  MUX2_X1 U669 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n248), .Z(n64) );
  MUX2_X1 U670 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n248), .Z(n65) );
  MUX2_X1 U671 ( .A(n65), .B(n64), .S(N11), .Z(n66) );
  MUX2_X1 U672 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U673 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n248), .Z(n68) );
  MUX2_X1 U674 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n248), .Z(n69) );
  MUX2_X1 U675 ( .A(n69), .B(n68), .S(N11), .Z(n70) );
  MUX2_X1 U676 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n248), .Z(n71) );
  MUX2_X1 U677 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n248), .Z(n72) );
  MUX2_X1 U678 ( .A(n72), .B(n71), .S(N11), .Z(n73) );
  MUX2_X1 U679 ( .A(n73), .B(n70), .S(N12), .Z(n74) );
  MUX2_X1 U680 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U681 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n248), .Z(n76) );
  MUX2_X1 U682 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n248), .Z(n77) );
  MUX2_X1 U683 ( .A(n77), .B(n76), .S(n243), .Z(n78) );
  MUX2_X1 U684 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n248), .Z(n79) );
  MUX2_X1 U685 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n248), .Z(n80) );
  MUX2_X1 U686 ( .A(n80), .B(n79), .S(N11), .Z(n81) );
  MUX2_X1 U687 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U688 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n249), .Z(n83) );
  MUX2_X1 U689 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n249), .Z(n84) );
  MUX2_X1 U690 ( .A(n84), .B(n83), .S(N11), .Z(n85) );
  MUX2_X1 U691 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n249), .Z(n86) );
  MUX2_X1 U692 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n249), .Z(n87) );
  MUX2_X1 U693 ( .A(n87), .B(n86), .S(N11), .Z(n88) );
  MUX2_X1 U694 ( .A(n88), .B(n85), .S(N12), .Z(n89) );
  MUX2_X1 U695 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U696 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U697 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n249), .Z(n91) );
  MUX2_X1 U698 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n249), .Z(n92) );
  MUX2_X1 U699 ( .A(n92), .B(n91), .S(N11), .Z(n93) );
  MUX2_X1 U700 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n249), .Z(n94) );
  MUX2_X1 U701 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n249), .Z(n95) );
  MUX2_X1 U702 ( .A(n95), .B(n94), .S(n244), .Z(n96) );
  MUX2_X1 U703 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U704 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n249), .Z(n98) );
  MUX2_X1 U705 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n249), .Z(n99) );
  MUX2_X1 U706 ( .A(n99), .B(n98), .S(n243), .Z(n100) );
  MUX2_X1 U707 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n249), .Z(n101) );
  MUX2_X1 U708 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n249), .Z(n102) );
  MUX2_X1 U709 ( .A(n102), .B(n101), .S(n242), .Z(n103) );
  MUX2_X1 U710 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U711 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U712 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n246), .Z(n106) );
  MUX2_X1 U713 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(N10), .Z(n107) );
  MUX2_X1 U714 ( .A(n107), .B(n106), .S(n242), .Z(n108) );
  MUX2_X1 U715 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n247), .Z(n109) );
  MUX2_X1 U716 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n250), .Z(n110) );
  MUX2_X1 U717 ( .A(n110), .B(n109), .S(n242), .Z(n111) );
  MUX2_X1 U718 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U719 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(N10), .Z(n113) );
  MUX2_X1 U720 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n248), .Z(n114) );
  MUX2_X1 U721 ( .A(n114), .B(n113), .S(n242), .Z(n115) );
  MUX2_X1 U722 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n116) );
  MUX2_X1 U723 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n249), .Z(n117) );
  MUX2_X1 U724 ( .A(n117), .B(n116), .S(n242), .Z(n118) );
  MUX2_X1 U725 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U726 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U727 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U728 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n250), .Z(n121) );
  MUX2_X1 U729 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n250), .Z(n122) );
  MUX2_X1 U730 ( .A(n122), .B(n121), .S(n242), .Z(n123) );
  MUX2_X1 U731 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n246), .Z(n124) );
  MUX2_X1 U732 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n250), .Z(n125) );
  MUX2_X1 U733 ( .A(n125), .B(n124), .S(n243), .Z(n126) );
  MUX2_X1 U734 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U735 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n246), .Z(n128) );
  MUX2_X1 U736 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n250), .Z(n129) );
  MUX2_X1 U737 ( .A(n129), .B(n128), .S(n242), .Z(n130) );
  MUX2_X1 U738 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n249), .Z(n131) );
  MUX2_X1 U739 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(N10), .Z(n132) );
  MUX2_X1 U740 ( .A(n132), .B(n131), .S(N11), .Z(n133) );
  MUX2_X1 U741 ( .A(n133), .B(n130), .S(N12), .Z(n134) );
  MUX2_X1 U742 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U743 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n245), .Z(n136) );
  MUX2_X1 U744 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n246), .Z(n137) );
  MUX2_X1 U745 ( .A(n137), .B(n136), .S(n242), .Z(n138) );
  MUX2_X1 U746 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n247), .Z(n139) );
  MUX2_X1 U747 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(N10), .Z(n140) );
  MUX2_X1 U748 ( .A(n140), .B(n139), .S(n243), .Z(n141) );
  MUX2_X1 U749 ( .A(n141), .B(n138), .S(N12), .Z(n142) );
  MUX2_X1 U750 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n248), .Z(n143) );
  MUX2_X1 U751 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(N10), .Z(n144) );
  MUX2_X1 U752 ( .A(n144), .B(n143), .S(n244), .Z(n145) );
  MUX2_X1 U753 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(N10), .Z(n146) );
  MUX2_X1 U754 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n147) );
  MUX2_X1 U755 ( .A(n147), .B(n146), .S(n242), .Z(n148) );
  MUX2_X1 U756 ( .A(n148), .B(n145), .S(N12), .Z(n149) );
  MUX2_X1 U757 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U758 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U759 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n245), .Z(n151) );
  MUX2_X1 U760 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n245), .Z(n152) );
  MUX2_X1 U761 ( .A(n152), .B(n151), .S(n243), .Z(n153) );
  MUX2_X1 U762 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n245), .Z(n154) );
  MUX2_X1 U763 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(N10), .Z(n155) );
  MUX2_X1 U764 ( .A(n155), .B(n154), .S(n243), .Z(n156) );
  MUX2_X1 U765 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U766 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(N10), .Z(n158) );
  MUX2_X1 U767 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(N10), .Z(n159) );
  MUX2_X1 U768 ( .A(n159), .B(n158), .S(n243), .Z(n160) );
  MUX2_X1 U769 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n247), .Z(n161) );
  MUX2_X1 U770 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(N10), .Z(n162) );
  MUX2_X1 U771 ( .A(n162), .B(n161), .S(n243), .Z(n163) );
  MUX2_X1 U772 ( .A(n163), .B(n160), .S(n241), .Z(n164) );
  MUX2_X1 U773 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U774 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n245), .Z(n166) );
  MUX2_X1 U775 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(N10), .Z(n167) );
  MUX2_X1 U776 ( .A(n167), .B(n166), .S(n243), .Z(n168) );
  MUX2_X1 U777 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n250), .Z(n169) );
  MUX2_X1 U778 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(N10), .Z(n170) );
  MUX2_X1 U779 ( .A(n170), .B(n169), .S(n243), .Z(n171) );
  MUX2_X1 U780 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U781 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n249), .Z(n173) );
  MUX2_X1 U782 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n250), .Z(n174) );
  MUX2_X1 U783 ( .A(n174), .B(n173), .S(n243), .Z(n175) );
  MUX2_X1 U784 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n250), .Z(n176) );
  MUX2_X1 U785 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n250), .Z(n177) );
  MUX2_X1 U786 ( .A(n177), .B(n176), .S(n243), .Z(n178) );
  MUX2_X1 U787 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U788 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U789 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U790 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n250), .Z(n181) );
  MUX2_X1 U791 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n245), .Z(n182) );
  MUX2_X1 U792 ( .A(n182), .B(n181), .S(n243), .Z(n183) );
  MUX2_X1 U793 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n249), .Z(n184) );
  MUX2_X1 U794 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n250), .Z(n185) );
  MUX2_X1 U795 ( .A(n185), .B(n184), .S(n243), .Z(n186) );
  MUX2_X1 U796 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U797 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n248), .Z(n188) );
  MUX2_X1 U798 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n250), .Z(n189) );
  MUX2_X1 U799 ( .A(n189), .B(n188), .S(n243), .Z(n190) );
  MUX2_X1 U800 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n249), .Z(n191) );
  MUX2_X1 U801 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n250), .Z(n192) );
  MUX2_X1 U802 ( .A(n192), .B(n191), .S(n243), .Z(n193) );
  MUX2_X1 U803 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U804 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U805 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n245), .Z(n196) );
  MUX2_X1 U806 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n250), .Z(n197) );
  MUX2_X1 U807 ( .A(n197), .B(n196), .S(n244), .Z(n198) );
  MUX2_X1 U808 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n246), .Z(n199) );
  MUX2_X1 U809 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n248), .Z(n200) );
  MUX2_X1 U810 ( .A(n200), .B(n199), .S(n244), .Z(n201) );
  MUX2_X1 U811 ( .A(n201), .B(n198), .S(n241), .Z(n202) );
  MUX2_X1 U812 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n248), .Z(n203) );
  MUX2_X1 U813 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n250), .Z(n204) );
  MUX2_X1 U814 ( .A(n204), .B(n203), .S(n244), .Z(n205) );
  MUX2_X1 U815 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n250), .Z(n206) );
  MUX2_X1 U816 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n246), .Z(n207) );
  MUX2_X1 U817 ( .A(n207), .B(n206), .S(n244), .Z(n208) );
  MUX2_X1 U818 ( .A(n208), .B(n205), .S(n241), .Z(n209) );
  MUX2_X1 U819 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U820 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U821 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(N10), .Z(n211) );
  MUX2_X1 U822 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n248), .Z(n212) );
  MUX2_X1 U823 ( .A(n212), .B(n211), .S(n244), .Z(n213) );
  MUX2_X1 U824 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n247), .Z(n214) );
  MUX2_X1 U825 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n245), .Z(n215) );
  MUX2_X1 U826 ( .A(n215), .B(n214), .S(n244), .Z(n216) );
  MUX2_X1 U827 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U828 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n247), .Z(n218) );
  MUX2_X1 U829 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n250), .Z(n219) );
  MUX2_X1 U830 ( .A(n219), .B(n218), .S(n244), .Z(n220) );
  MUX2_X1 U831 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n246), .Z(n221) );
  MUX2_X1 U832 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n250), .Z(n222) );
  MUX2_X1 U833 ( .A(n222), .B(n221), .S(n244), .Z(n223) );
  MUX2_X1 U834 ( .A(n223), .B(n220), .S(n241), .Z(n224) );
  MUX2_X1 U835 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U836 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n250), .Z(n226) );
  MUX2_X1 U837 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n249), .Z(n227) );
  MUX2_X1 U838 ( .A(n227), .B(n226), .S(n244), .Z(n228) );
  MUX2_X1 U839 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n247), .Z(n229) );
  MUX2_X1 U840 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n250), .Z(n230) );
  MUX2_X1 U841 ( .A(n230), .B(n229), .S(n244), .Z(n231) );
  MUX2_X1 U842 ( .A(n231), .B(n228), .S(N12), .Z(n232) );
  MUX2_X1 U843 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n248), .Z(n233) );
  MUX2_X1 U844 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n247), .Z(n234) );
  MUX2_X1 U845 ( .A(n234), .B(n233), .S(n244), .Z(n235) );
  MUX2_X1 U846 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n249), .Z(n236) );
  MUX2_X1 U847 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n245), .Z(n237) );
  MUX2_X1 U848 ( .A(n237), .B(n236), .S(n244), .Z(n238) );
  MUX2_X1 U849 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U850 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U851 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U852 ( .A(N11), .Z(n242) );
  CLKBUF_X1 U853 ( .A(n250), .Z(n245) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_12 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X2 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(N10), .Z(n247) );
  BUF_X1 U4 ( .A(N10), .Z(n246) );
  BUF_X1 U5 ( .A(n250), .Z(n248) );
  BUF_X1 U6 ( .A(N10), .Z(n249) );
  BUF_X1 U7 ( .A(N10), .Z(n250) );
  INV_X1 U8 ( .A(n1111), .ZN(n841) );
  INV_X1 U9 ( .A(n1100), .ZN(n840) );
  INV_X1 U10 ( .A(n1090), .ZN(n839) );
  INV_X1 U11 ( .A(n1080), .ZN(n838) );
  INV_X1 U12 ( .A(n1070), .ZN(n837) );
  INV_X1 U13 ( .A(n1060), .ZN(n836) );
  INV_X1 U14 ( .A(n1051), .ZN(n835) );
  INV_X1 U15 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U16 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U18 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U19 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U20 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U21 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U22 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U23 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U24 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U26 ( .A(n1131), .ZN(n816) );
  INV_X1 U27 ( .A(n1121), .ZN(n815) );
  INV_X1 U28 ( .A(n887), .ZN(n814) );
  INV_X1 U29 ( .A(n878), .ZN(n813) );
  INV_X1 U30 ( .A(n869), .ZN(n812) );
  INV_X1 U31 ( .A(n860), .ZN(n811) );
  INV_X1 U32 ( .A(n851), .ZN(n810) );
  INV_X1 U33 ( .A(n987), .ZN(n828) );
  INV_X1 U34 ( .A(n978), .ZN(n827) );
  INV_X1 U35 ( .A(n969), .ZN(n826) );
  INV_X1 U36 ( .A(n914), .ZN(n820) );
  INV_X1 U37 ( .A(n905), .ZN(n819) );
  INV_X1 U38 ( .A(n896), .ZN(n818) );
  INV_X1 U39 ( .A(n1033), .ZN(n833) );
  INV_X1 U40 ( .A(n1023), .ZN(n832) );
  INV_X1 U41 ( .A(n1014), .ZN(n831) );
  INV_X1 U42 ( .A(n1005), .ZN(n830) );
  INV_X1 U43 ( .A(n996), .ZN(n829) );
  INV_X1 U44 ( .A(n960), .ZN(n825) );
  INV_X1 U45 ( .A(n950), .ZN(n824) );
  INV_X1 U46 ( .A(n941), .ZN(n823) );
  INV_X1 U47 ( .A(n932), .ZN(n822) );
  INV_X1 U48 ( .A(n923), .ZN(n821) );
  INV_X1 U49 ( .A(n1142), .ZN(n817) );
  BUF_X1 U50 ( .A(N11), .Z(n242) );
  BUF_X1 U51 ( .A(N11), .Z(n243) );
  BUF_X1 U52 ( .A(N11), .Z(n244) );
  INV_X1 U53 ( .A(N10), .ZN(n251) );
  BUF_X1 U54 ( .A(N12), .Z(n241) );
  NOR3_X1 U55 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U56 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U57 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U58 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U59 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U60 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U61 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U62 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U63 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U64 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U65 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U67 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U69 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U70 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U71 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U72 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U73 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U74 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U75 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U76 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U77 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U79 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U81 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U82 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U83 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U84 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U85 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U86 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U87 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U88 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U89 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U90 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U91 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U92 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U93 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U94 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U95 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U96 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U97 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U98 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U99 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U100 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U101 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U102 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U103 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U104 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U105 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U106 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U107 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U108 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U109 ( .A(n988), .ZN(n705) );
  AOI22_X1 U110 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U111 ( .A(n986), .ZN(n704) );
  AOI22_X1 U112 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U113 ( .A(n985), .ZN(n703) );
  AOI22_X1 U114 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U115 ( .A(n984), .ZN(n702) );
  AOI22_X1 U116 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U117 ( .A(n983), .ZN(n701) );
  AOI22_X1 U118 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U119 ( .A(n982), .ZN(n700) );
  AOI22_X1 U120 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U121 ( .A(n981), .ZN(n699) );
  AOI22_X1 U122 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U123 ( .A(n980), .ZN(n698) );
  AOI22_X1 U124 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U125 ( .A(n949), .ZN(n672) );
  AOI22_X1 U126 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U127 ( .A(n948), .ZN(n671) );
  AOI22_X1 U128 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U129 ( .A(n915), .ZN(n641) );
  AOI22_X1 U130 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U131 ( .A(n913), .ZN(n640) );
  AOI22_X1 U132 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U133 ( .A(n912), .ZN(n639) );
  AOI22_X1 U134 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U135 ( .A(n911), .ZN(n638) );
  AOI22_X1 U136 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U137 ( .A(n910), .ZN(n637) );
  AOI22_X1 U138 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U139 ( .A(n909), .ZN(n636) );
  AOI22_X1 U140 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U141 ( .A(n908), .ZN(n635) );
  AOI22_X1 U142 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U143 ( .A(n907), .ZN(n634) );
  AOI22_X1 U144 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U145 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U146 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U147 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U148 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U149 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U150 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U151 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U152 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U153 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U154 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U155 ( .A(n947), .ZN(n670) );
  AOI22_X1 U156 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U157 ( .A(n946), .ZN(n669) );
  AOI22_X1 U158 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U159 ( .A(n945), .ZN(n668) );
  AOI22_X1 U160 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U161 ( .A(n944), .ZN(n667) );
  AOI22_X1 U162 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U163 ( .A(n943), .ZN(n666) );
  AOI22_X1 U164 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U165 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U166 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U167 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U168 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U169 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U170 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U171 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U172 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U173 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U174 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U175 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U176 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U177 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U178 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U179 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U180 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U181 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U182 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U183 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U184 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U185 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U186 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U187 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U188 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U189 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U190 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U191 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U192 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U193 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U194 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U195 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U196 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U197 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U198 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U199 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U200 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U201 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U202 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U203 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U204 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U205 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U206 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U207 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U208 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U209 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U210 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U211 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U212 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U213 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U214 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U215 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U216 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U217 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U218 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U219 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U220 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U221 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U222 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U223 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U224 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U225 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U226 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U227 ( .A(n999), .ZN(n715) );
  AOI22_X1 U228 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U229 ( .A(n998), .ZN(n714) );
  AOI22_X1 U230 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U231 ( .A(n951), .ZN(n673) );
  AOI22_X1 U232 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U233 ( .A(n979), .ZN(n697) );
  AOI22_X1 U234 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U235 ( .A(n977), .ZN(n696) );
  AOI22_X1 U236 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U237 ( .A(n976), .ZN(n695) );
  AOI22_X1 U238 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U239 ( .A(n975), .ZN(n694) );
  AOI22_X1 U240 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U241 ( .A(n974), .ZN(n693) );
  AOI22_X1 U242 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U243 ( .A(n973), .ZN(n692) );
  AOI22_X1 U244 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U245 ( .A(n972), .ZN(n691) );
  AOI22_X1 U246 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U247 ( .A(n971), .ZN(n690) );
  AOI22_X1 U248 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U249 ( .A(n970), .ZN(n689) );
  AOI22_X1 U250 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U251 ( .A(n968), .ZN(n688) );
  AOI22_X1 U252 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U253 ( .A(n967), .ZN(n687) );
  AOI22_X1 U254 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U255 ( .A(n966), .ZN(n686) );
  AOI22_X1 U256 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U257 ( .A(n965), .ZN(n685) );
  AOI22_X1 U258 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U259 ( .A(n964), .ZN(n684) );
  AOI22_X1 U260 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U261 ( .A(n963), .ZN(n683) );
  AOI22_X1 U262 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U263 ( .A(n962), .ZN(n682) );
  AOI22_X1 U264 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U265 ( .A(n942), .ZN(n665) );
  AOI22_X1 U266 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U267 ( .A(n940), .ZN(n664) );
  AOI22_X1 U268 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U269 ( .A(n939), .ZN(n663) );
  AOI22_X1 U270 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U271 ( .A(n938), .ZN(n662) );
  AOI22_X1 U272 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U273 ( .A(n937), .ZN(n661) );
  AOI22_X1 U274 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U275 ( .A(n936), .ZN(n660) );
  AOI22_X1 U276 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U277 ( .A(n935), .ZN(n659) );
  AOI22_X1 U278 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U279 ( .A(n934), .ZN(n658) );
  AOI22_X1 U280 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U281 ( .A(n933), .ZN(n657) );
  AOI22_X1 U282 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U283 ( .A(n931), .ZN(n656) );
  AOI22_X1 U284 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U285 ( .A(n930), .ZN(n655) );
  AOI22_X1 U286 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U287 ( .A(n929), .ZN(n654) );
  AOI22_X1 U288 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U289 ( .A(n928), .ZN(n653) );
  AOI22_X1 U290 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U291 ( .A(n927), .ZN(n652) );
  AOI22_X1 U292 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U293 ( .A(n926), .ZN(n651) );
  AOI22_X1 U294 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U295 ( .A(n925), .ZN(n650) );
  AOI22_X1 U296 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U297 ( .A(n906), .ZN(n633) );
  AOI22_X1 U298 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U299 ( .A(n904), .ZN(n632) );
  AOI22_X1 U300 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U301 ( .A(n903), .ZN(n631) );
  AOI22_X1 U302 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U303 ( .A(n902), .ZN(n630) );
  AOI22_X1 U304 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U305 ( .A(n901), .ZN(n629) );
  AOI22_X1 U306 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U307 ( .A(n900), .ZN(n628) );
  AOI22_X1 U308 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U309 ( .A(n899), .ZN(n627) );
  AOI22_X1 U310 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U311 ( .A(n898), .ZN(n626) );
  AOI22_X1 U312 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U313 ( .A(n897), .ZN(n625) );
  AOI22_X1 U314 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U315 ( .A(n895), .ZN(n624) );
  AOI22_X1 U316 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U317 ( .A(n894), .ZN(n623) );
  AOI22_X1 U318 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U319 ( .A(n893), .ZN(n622) );
  AOI22_X1 U320 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U321 ( .A(n892), .ZN(n621) );
  AOI22_X1 U322 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U323 ( .A(n891), .ZN(n620) );
  AOI22_X1 U324 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U325 ( .A(n890), .ZN(n619) );
  AOI22_X1 U326 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U327 ( .A(n889), .ZN(n618) );
  AOI22_X1 U328 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U329 ( .A(N12), .ZN(n253) );
  INV_X1 U330 ( .A(N11), .ZN(n252) );
  INV_X1 U331 ( .A(n997), .ZN(n713) );
  AOI22_X1 U332 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U333 ( .A(n995), .ZN(n712) );
  AOI22_X1 U334 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U335 ( .A(n994), .ZN(n711) );
  AOI22_X1 U336 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U337 ( .A(n993), .ZN(n710) );
  AOI22_X1 U338 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U339 ( .A(n992), .ZN(n709) );
  AOI22_X1 U340 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U341 ( .A(n991), .ZN(n708) );
  AOI22_X1 U342 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U343 ( .A(n990), .ZN(n707) );
  AOI22_X1 U344 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U345 ( .A(n989), .ZN(n706) );
  AOI22_X1 U346 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U347 ( .A(n924), .ZN(n649) );
  AOI22_X1 U348 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U349 ( .A(n922), .ZN(n648) );
  AOI22_X1 U350 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U351 ( .A(n921), .ZN(n647) );
  AOI22_X1 U352 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U353 ( .A(n920), .ZN(n646) );
  AOI22_X1 U354 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U355 ( .A(n919), .ZN(n645) );
  AOI22_X1 U356 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U357 ( .A(n918), .ZN(n644) );
  AOI22_X1 U358 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U359 ( .A(n917), .ZN(n643) );
  AOI22_X1 U360 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U361 ( .A(n916), .ZN(n642) );
  AOI22_X1 U362 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U363 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U364 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U365 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U366 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U367 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U368 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U369 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U370 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U371 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U372 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U373 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U374 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U375 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U376 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U377 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U378 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U379 ( .A(n961), .ZN(n681) );
  AOI22_X1 U380 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U381 ( .A(n959), .ZN(n680) );
  AOI22_X1 U382 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U383 ( .A(n958), .ZN(n679) );
  AOI22_X1 U384 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U385 ( .A(n957), .ZN(n678) );
  AOI22_X1 U386 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U387 ( .A(n956), .ZN(n677) );
  AOI22_X1 U388 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U389 ( .A(n955), .ZN(n676) );
  AOI22_X1 U390 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U391 ( .A(n954), .ZN(n675) );
  AOI22_X1 U392 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U393 ( .A(n953), .ZN(n674) );
  AOI22_X1 U394 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U395 ( .A(n888), .ZN(n617) );
  AOI22_X1 U396 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U397 ( .A(n886), .ZN(n616) );
  AOI22_X1 U398 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U399 ( .A(n885), .ZN(n615) );
  AOI22_X1 U400 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U401 ( .A(n884), .ZN(n614) );
  AOI22_X1 U402 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U403 ( .A(n883), .ZN(n613) );
  AOI22_X1 U404 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U405 ( .A(n882), .ZN(n612) );
  AOI22_X1 U406 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U407 ( .A(n881), .ZN(n611) );
  AOI22_X1 U408 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U409 ( .A(n880), .ZN(n610) );
  AOI22_X1 U410 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U411 ( .A(n879), .ZN(n609) );
  AOI22_X1 U412 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U413 ( .A(n877), .ZN(n608) );
  AOI22_X1 U414 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U415 ( .A(n876), .ZN(n607) );
  AOI22_X1 U416 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U417 ( .A(n875), .ZN(n606) );
  AOI22_X1 U418 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U419 ( .A(n874), .ZN(n605) );
  AOI22_X1 U420 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U421 ( .A(n873), .ZN(n604) );
  AOI22_X1 U422 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U423 ( .A(n872), .ZN(n603) );
  AOI22_X1 U424 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U425 ( .A(n871), .ZN(n602) );
  AOI22_X1 U426 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U427 ( .A(n870), .ZN(n601) );
  AOI22_X1 U428 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U429 ( .A(n868), .ZN(n600) );
  AOI22_X1 U430 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U431 ( .A(n867), .ZN(n599) );
  AOI22_X1 U432 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U433 ( .A(n866), .ZN(n598) );
  AOI22_X1 U434 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U435 ( .A(n865), .ZN(n597) );
  AOI22_X1 U436 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U437 ( .A(n864), .ZN(n596) );
  AOI22_X1 U438 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U439 ( .A(n863), .ZN(n595) );
  AOI22_X1 U440 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U441 ( .A(n862), .ZN(n594) );
  AOI22_X1 U442 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U443 ( .A(n861), .ZN(n293) );
  AOI22_X1 U444 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U445 ( .A(n859), .ZN(n292) );
  AOI22_X1 U446 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U447 ( .A(n858), .ZN(n291) );
  AOI22_X1 U448 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U449 ( .A(n857), .ZN(n290) );
  AOI22_X1 U450 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U451 ( .A(n856), .ZN(n289) );
  AOI22_X1 U452 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U453 ( .A(n855), .ZN(n288) );
  AOI22_X1 U454 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U455 ( .A(n854), .ZN(n287) );
  AOI22_X1 U456 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U457 ( .A(n853), .ZN(n286) );
  AOI22_X1 U458 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U459 ( .A(n852), .ZN(n285) );
  AOI22_X1 U460 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U461 ( .A(n850), .ZN(n284) );
  AOI22_X1 U462 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U463 ( .A(n849), .ZN(n283) );
  AOI22_X1 U464 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U465 ( .A(n848), .ZN(n282) );
  AOI22_X1 U466 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U467 ( .A(n847), .ZN(n281) );
  AOI22_X1 U468 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U469 ( .A(n846), .ZN(n280) );
  AOI22_X1 U470 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U471 ( .A(n845), .ZN(n279) );
  AOI22_X1 U472 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U473 ( .A(n844), .ZN(n278) );
  AOI22_X1 U474 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U475 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U476 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U477 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U478 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U479 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U480 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U481 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U482 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U483 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U484 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U485 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U486 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U487 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U488 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U489 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U490 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U491 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U492 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U493 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U494 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U495 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U496 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U497 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U498 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U499 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U500 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U501 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U502 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U503 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U504 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U505 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U506 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U507 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U508 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U509 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U510 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U511 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U512 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U513 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U514 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U515 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U516 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U517 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U518 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U519 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U520 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U521 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U522 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U523 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U524 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U525 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U526 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U527 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U528 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U529 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U530 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U531 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U532 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U533 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U534 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U535 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U536 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U537 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U538 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U539 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U540 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U541 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U542 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U543 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U544 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U545 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U546 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U547 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U548 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U549 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U550 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U551 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U552 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U553 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U554 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U555 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U556 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U557 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U558 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U559 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U560 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U561 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U562 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U563 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U564 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U565 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U566 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U567 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U568 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U569 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U570 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U571 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U572 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U573 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U574 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U575 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U576 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U577 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U578 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U579 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U580 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U581 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U582 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U583 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U584 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U585 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U586 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U587 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U588 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U589 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U590 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U591 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U592 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U593 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U594 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U595 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U596 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U597 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U598 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U599 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U600 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U601 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U602 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U603 ( .A(N13), .ZN(n842) );
  INV_X1 U604 ( .A(N14), .ZN(n843) );
  MUX2_X1 U605 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n245), .Z(n1) );
  MUX2_X1 U606 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n245), .Z(n2) );
  MUX2_X1 U607 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U608 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n245), .Z(n4) );
  MUX2_X1 U609 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n245), .Z(n5) );
  MUX2_X1 U610 ( .A(n5), .B(n4), .S(n243), .Z(n6) );
  MUX2_X1 U611 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U612 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n245), .Z(n8) );
  MUX2_X1 U613 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n245), .Z(n9) );
  MUX2_X1 U614 ( .A(n9), .B(n8), .S(n242), .Z(n10) );
  MUX2_X1 U615 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n245), .Z(n11) );
  MUX2_X1 U616 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n245), .Z(n12) );
  MUX2_X1 U617 ( .A(n12), .B(n11), .S(n244), .Z(n13) );
  MUX2_X1 U618 ( .A(n13), .B(n10), .S(n241), .Z(n14) );
  MUX2_X1 U619 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U620 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n246), .Z(n16) );
  MUX2_X1 U621 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n246), .Z(n17) );
  MUX2_X1 U622 ( .A(n17), .B(n16), .S(n244), .Z(n18) );
  MUX2_X1 U623 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n246), .Z(n19) );
  MUX2_X1 U624 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n246), .Z(n20) );
  MUX2_X1 U625 ( .A(n20), .B(n19), .S(N11), .Z(n21) );
  MUX2_X1 U626 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U627 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n246), .Z(n23) );
  MUX2_X1 U628 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n246), .Z(n24) );
  MUX2_X1 U629 ( .A(n24), .B(n23), .S(n243), .Z(n25) );
  MUX2_X1 U630 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n246), .Z(n26) );
  MUX2_X1 U631 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n246), .Z(n27) );
  MUX2_X1 U632 ( .A(n27), .B(n26), .S(N11), .Z(n28) );
  MUX2_X1 U633 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U634 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U635 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U636 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n246), .Z(n31) );
  MUX2_X1 U637 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n246), .Z(n32) );
  MUX2_X1 U638 ( .A(n32), .B(n31), .S(n243), .Z(n33) );
  MUX2_X1 U639 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n246), .Z(n34) );
  MUX2_X1 U640 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n246), .Z(n35) );
  MUX2_X1 U641 ( .A(n35), .B(n34), .S(n244), .Z(n36) );
  MUX2_X1 U642 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U643 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n247), .Z(n38) );
  MUX2_X1 U644 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n247), .Z(n39) );
  MUX2_X1 U645 ( .A(n39), .B(n38), .S(n243), .Z(n40) );
  MUX2_X1 U646 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n247), .Z(n41) );
  MUX2_X1 U647 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n247), .Z(n42) );
  MUX2_X1 U648 ( .A(n42), .B(n41), .S(N11), .Z(n43) );
  MUX2_X1 U649 ( .A(n43), .B(n40), .S(n241), .Z(n44) );
  MUX2_X1 U650 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U651 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n247), .Z(n46) );
  MUX2_X1 U652 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n247), .Z(n47) );
  MUX2_X1 U653 ( .A(n47), .B(n46), .S(n242), .Z(n48) );
  MUX2_X1 U654 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n247), .Z(n49) );
  MUX2_X1 U655 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n247), .Z(n50) );
  MUX2_X1 U656 ( .A(n50), .B(n49), .S(N11), .Z(n51) );
  MUX2_X1 U657 ( .A(n51), .B(n48), .S(n241), .Z(n52) );
  MUX2_X1 U658 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n247), .Z(n53) );
  MUX2_X1 U659 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n247), .Z(n54) );
  MUX2_X1 U660 ( .A(n54), .B(n53), .S(n242), .Z(n55) );
  MUX2_X1 U661 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n247), .Z(n56) );
  MUX2_X1 U662 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n247), .Z(n57) );
  MUX2_X1 U663 ( .A(n57), .B(n56), .S(N11), .Z(n58) );
  MUX2_X1 U664 ( .A(n58), .B(n55), .S(n241), .Z(n59) );
  MUX2_X1 U665 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U666 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U667 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n248), .Z(n61) );
  MUX2_X1 U668 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n248), .Z(n62) );
  MUX2_X1 U669 ( .A(n62), .B(n61), .S(N11), .Z(n63) );
  MUX2_X1 U670 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n248), .Z(n64) );
  MUX2_X1 U671 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n248), .Z(n65) );
  MUX2_X1 U672 ( .A(n65), .B(n64), .S(n243), .Z(n66) );
  MUX2_X1 U673 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U674 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n248), .Z(n68) );
  MUX2_X1 U675 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n248), .Z(n69) );
  MUX2_X1 U676 ( .A(n69), .B(n68), .S(n244), .Z(n70) );
  MUX2_X1 U677 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n248), .Z(n71) );
  MUX2_X1 U678 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n248), .Z(n72) );
  MUX2_X1 U679 ( .A(n72), .B(n71), .S(n242), .Z(n73) );
  MUX2_X1 U680 ( .A(n73), .B(n70), .S(N12), .Z(n74) );
  MUX2_X1 U681 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U682 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n248), .Z(n76) );
  MUX2_X1 U683 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n248), .Z(n77) );
  MUX2_X1 U684 ( .A(n77), .B(n76), .S(N11), .Z(n78) );
  MUX2_X1 U685 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n248), .Z(n79) );
  MUX2_X1 U686 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n248), .Z(n80) );
  MUX2_X1 U687 ( .A(n80), .B(n79), .S(N11), .Z(n81) );
  MUX2_X1 U688 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U689 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n249), .Z(n83) );
  MUX2_X1 U690 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n249), .Z(n84) );
  MUX2_X1 U691 ( .A(n84), .B(n83), .S(n244), .Z(n85) );
  MUX2_X1 U692 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n249), .Z(n86) );
  MUX2_X1 U693 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n249), .Z(n87) );
  MUX2_X1 U694 ( .A(n87), .B(n86), .S(n242), .Z(n88) );
  MUX2_X1 U695 ( .A(n88), .B(n85), .S(N12), .Z(n89) );
  MUX2_X1 U696 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U697 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U698 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n249), .Z(n91) );
  MUX2_X1 U699 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n249), .Z(n92) );
  MUX2_X1 U700 ( .A(n92), .B(n91), .S(N11), .Z(n93) );
  MUX2_X1 U701 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n249), .Z(n94) );
  MUX2_X1 U702 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n249), .Z(n95) );
  MUX2_X1 U703 ( .A(n95), .B(n94), .S(N11), .Z(n96) );
  MUX2_X1 U704 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U705 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n249), .Z(n98) );
  MUX2_X1 U706 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n249), .Z(n99) );
  MUX2_X1 U707 ( .A(n99), .B(n98), .S(N11), .Z(n100) );
  MUX2_X1 U708 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n249), .Z(n101) );
  MUX2_X1 U709 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n249), .Z(n102) );
  MUX2_X1 U710 ( .A(n102), .B(n101), .S(N11), .Z(n103) );
  MUX2_X1 U711 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U712 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U713 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n246), .Z(n106) );
  MUX2_X1 U714 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n245), .Z(n107) );
  MUX2_X1 U715 ( .A(n107), .B(n106), .S(n242), .Z(n108) );
  MUX2_X1 U716 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n249), .Z(n109) );
  MUX2_X1 U717 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n110) );
  MUX2_X1 U718 ( .A(n110), .B(n109), .S(n242), .Z(n111) );
  MUX2_X1 U719 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U720 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n250), .Z(n113) );
  MUX2_X1 U721 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n114) );
  MUX2_X1 U722 ( .A(n114), .B(n113), .S(n242), .Z(n115) );
  MUX2_X1 U723 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n116) );
  MUX2_X1 U724 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n117) );
  MUX2_X1 U725 ( .A(n117), .B(n116), .S(n242), .Z(n118) );
  MUX2_X1 U726 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U727 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U728 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U729 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(N10), .Z(n121) );
  MUX2_X1 U730 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(N10), .Z(n122) );
  MUX2_X1 U731 ( .A(n122), .B(n121), .S(n242), .Z(n123) );
  MUX2_X1 U732 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(N10), .Z(n124) );
  MUX2_X1 U733 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n125) );
  MUX2_X1 U734 ( .A(n125), .B(n124), .S(n242), .Z(n126) );
  MUX2_X1 U735 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U736 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n249), .Z(n128) );
  MUX2_X1 U737 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n245), .Z(n129) );
  MUX2_X1 U738 ( .A(n129), .B(n128), .S(n242), .Z(n130) );
  MUX2_X1 U739 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n246), .Z(n131) );
  MUX2_X1 U740 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n245), .Z(n132) );
  MUX2_X1 U741 ( .A(n132), .B(n131), .S(n242), .Z(n133) );
  MUX2_X1 U742 ( .A(n133), .B(n130), .S(N12), .Z(n134) );
  MUX2_X1 U743 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U744 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n246), .Z(n136) );
  MUX2_X1 U745 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n249), .Z(n137) );
  MUX2_X1 U746 ( .A(n137), .B(n136), .S(n242), .Z(n138) );
  MUX2_X1 U747 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n245), .Z(n139) );
  MUX2_X1 U748 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n246), .Z(n140) );
  MUX2_X1 U749 ( .A(n140), .B(n139), .S(n242), .Z(n141) );
  MUX2_X1 U750 ( .A(n141), .B(n138), .S(N12), .Z(n142) );
  MUX2_X1 U751 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n247), .Z(n143) );
  MUX2_X1 U752 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n249), .Z(n144) );
  MUX2_X1 U753 ( .A(n144), .B(n143), .S(n242), .Z(n145) );
  MUX2_X1 U754 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n247), .Z(n146) );
  MUX2_X1 U755 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n247), .Z(n147) );
  MUX2_X1 U756 ( .A(n147), .B(n146), .S(n242), .Z(n148) );
  MUX2_X1 U757 ( .A(n148), .B(n145), .S(N12), .Z(n149) );
  MUX2_X1 U758 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U759 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U760 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n245), .Z(n151) );
  MUX2_X1 U761 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n247), .Z(n152) );
  MUX2_X1 U762 ( .A(n152), .B(n151), .S(n243), .Z(n153) );
  MUX2_X1 U763 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n245), .Z(n154) );
  MUX2_X1 U764 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n246), .Z(n155) );
  MUX2_X1 U765 ( .A(n155), .B(n154), .S(n243), .Z(n156) );
  MUX2_X1 U766 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U767 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n246), .Z(n158) );
  MUX2_X1 U768 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n249), .Z(n159) );
  MUX2_X1 U769 ( .A(n159), .B(n158), .S(n243), .Z(n160) );
  MUX2_X1 U770 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n245), .Z(n161) );
  MUX2_X1 U771 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n247), .Z(n162) );
  MUX2_X1 U772 ( .A(n162), .B(n161), .S(n243), .Z(n163) );
  MUX2_X1 U773 ( .A(n163), .B(n160), .S(n241), .Z(n164) );
  MUX2_X1 U774 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U775 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n245), .Z(n166) );
  MUX2_X1 U776 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n247), .Z(n167) );
  MUX2_X1 U777 ( .A(n167), .B(n166), .S(n243), .Z(n168) );
  MUX2_X1 U778 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n249), .Z(n169) );
  MUX2_X1 U779 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n245), .Z(n170) );
  MUX2_X1 U780 ( .A(n170), .B(n169), .S(n243), .Z(n171) );
  MUX2_X1 U781 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U782 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n250), .Z(n173) );
  MUX2_X1 U783 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n250), .Z(n174) );
  MUX2_X1 U784 ( .A(n174), .B(n173), .S(n243), .Z(n175) );
  MUX2_X1 U785 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n245), .Z(n176) );
  MUX2_X1 U786 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n250), .Z(n177) );
  MUX2_X1 U787 ( .A(n177), .B(n176), .S(n243), .Z(n178) );
  MUX2_X1 U788 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U789 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U790 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U791 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n247), .Z(n181) );
  MUX2_X1 U792 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n246), .Z(n182) );
  MUX2_X1 U793 ( .A(n182), .B(n181), .S(n243), .Z(n183) );
  MUX2_X1 U794 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n245), .Z(n184) );
  MUX2_X1 U795 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n250), .Z(n185) );
  MUX2_X1 U796 ( .A(n185), .B(n184), .S(n243), .Z(n186) );
  MUX2_X1 U797 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U798 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n249), .Z(n188) );
  MUX2_X1 U799 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n250), .Z(n189) );
  MUX2_X1 U800 ( .A(n189), .B(n188), .S(n243), .Z(n190) );
  MUX2_X1 U801 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n245), .Z(n191) );
  MUX2_X1 U802 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n245), .Z(n192) );
  MUX2_X1 U803 ( .A(n192), .B(n191), .S(n243), .Z(n193) );
  MUX2_X1 U804 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U805 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U806 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n247), .Z(n196) );
  MUX2_X1 U807 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n247), .Z(n197) );
  MUX2_X1 U808 ( .A(n197), .B(n196), .S(n244), .Z(n198) );
  MUX2_X1 U809 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n249), .Z(n199) );
  MUX2_X1 U810 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n249), .Z(n200) );
  MUX2_X1 U811 ( .A(n200), .B(n199), .S(n244), .Z(n201) );
  MUX2_X1 U812 ( .A(n201), .B(n198), .S(n241), .Z(n202) );
  MUX2_X1 U813 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n246), .Z(n203) );
  MUX2_X1 U814 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n246), .Z(n204) );
  MUX2_X1 U815 ( .A(n204), .B(n203), .S(n244), .Z(n205) );
  MUX2_X1 U816 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n250), .Z(n206) );
  MUX2_X1 U817 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n250), .Z(n207) );
  MUX2_X1 U818 ( .A(n207), .B(n206), .S(n244), .Z(n208) );
  MUX2_X1 U819 ( .A(n208), .B(n205), .S(n241), .Z(n209) );
  MUX2_X1 U820 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U821 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U822 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n250), .Z(n211) );
  MUX2_X1 U823 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n250), .Z(n212) );
  MUX2_X1 U824 ( .A(n212), .B(n211), .S(n244), .Z(n213) );
  MUX2_X1 U825 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n245), .Z(n214) );
  MUX2_X1 U826 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n245), .Z(n215) );
  MUX2_X1 U827 ( .A(n215), .B(n214), .S(n244), .Z(n216) );
  MUX2_X1 U828 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U829 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n247), .Z(n218) );
  MUX2_X1 U830 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n249), .Z(n219) );
  MUX2_X1 U831 ( .A(n219), .B(n218), .S(n244), .Z(n220) );
  MUX2_X1 U832 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n250), .Z(n221) );
  MUX2_X1 U833 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n222) );
  MUX2_X1 U834 ( .A(n222), .B(n221), .S(n244), .Z(n223) );
  MUX2_X1 U835 ( .A(n223), .B(n220), .S(n241), .Z(n224) );
  MUX2_X1 U836 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U837 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n250), .Z(n226) );
  MUX2_X1 U838 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n247), .Z(n227) );
  MUX2_X1 U839 ( .A(n227), .B(n226), .S(n244), .Z(n228) );
  MUX2_X1 U840 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n249), .Z(n229) );
  MUX2_X1 U841 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n230) );
  MUX2_X1 U842 ( .A(n230), .B(n229), .S(n244), .Z(n231) );
  MUX2_X1 U843 ( .A(n231), .B(n228), .S(N12), .Z(n232) );
  MUX2_X1 U844 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n246), .Z(n233) );
  MUX2_X1 U845 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n234) );
  MUX2_X1 U846 ( .A(n234), .B(n233), .S(n244), .Z(n235) );
  MUX2_X1 U847 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n246), .Z(n236) );
  MUX2_X1 U848 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n237) );
  MUX2_X1 U849 ( .A(n237), .B(n236), .S(n244), .Z(n238) );
  MUX2_X1 U850 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U851 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U852 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U853 ( .A(N10), .Z(n245) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_11 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n256), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n257), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n258), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n259), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n260), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n261), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n262), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n263), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n264), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n265), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n266), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n267), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n268), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n269), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n270), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n271), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n272), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n273), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n274), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n275), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n276), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n277), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n278), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n279), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n280), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n281), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n282), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n283), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n284), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n285), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n286), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n287), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n288), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n289), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n290), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n291), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n292), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n293), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n594), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n595), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n596), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n597), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n598), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n599), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n600), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n601), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n602), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n603), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n604), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n605), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n606), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n607), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n608), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n609), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n610), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n611), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n612), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n613), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n614), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n615), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n616), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n617), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n618), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n619), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n620), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n621), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n622), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n623), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n624), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n625), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n626), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n627), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n628), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n629), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n630), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n631), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n632), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n633), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n634), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n635), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n636), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n637), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n638), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n639), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n640), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n641), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n642), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n643), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n644), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n645), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n646), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n647), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n648), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n649), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n650), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n651), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n652), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n653), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n654), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n655), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n656), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n657), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n658), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n659), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n660), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n661), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n662), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n663), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n664), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n665), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n666), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n667), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n668), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n669), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n670), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n671), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n672), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n673), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n674), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n675), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n676), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n677), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n678), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n679), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n680), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n681), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n682), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n683), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n684), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n685), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n686), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n687), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n688), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n689), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n690), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n691), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n692), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n693), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n694), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n695), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n696), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n697), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n698), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n699), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n700), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n701), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n702), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n703), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n704), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n705), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n706), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n707), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n708), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n709), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n710), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n711), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n712), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n713), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n714), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n715), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n716), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n717), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n718), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n719), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n720), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n721), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n722), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n723), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n724), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n725), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n726), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n727), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n728), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n729), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n730), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n731), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n732), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n733), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n734), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n735), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n736), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n737), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n738), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n739), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n740), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n741), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n742), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n743), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n744), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n745), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n746), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n747), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n748), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n749), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n750), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n751), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n752), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n753), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n754), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n755), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n756), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n757), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n758), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n759), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n760), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n761), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n762), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n763), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n764), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n765), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n766), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n767), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n768), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n769), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n770), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n771), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n772), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n773), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n774), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n775), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n776), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n777), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n778), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n779), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n780), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n781), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n782), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n783), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n784), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n785), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n786), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n787), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n788), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n789), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n790), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n791), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n792), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n793), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n794), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n795), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n796), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n797), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n798), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n799), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n800), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n801), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n802), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n803), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n804), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n805), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n806), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n807), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n808), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n809), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n810), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n811), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(n252), .Z(n251) );
  BUF_X1 U5 ( .A(n252), .Z(n248) );
  BUF_X1 U6 ( .A(n252), .Z(n247) );
  BUF_X1 U7 ( .A(n252), .Z(n249) );
  BUF_X1 U8 ( .A(n252), .Z(n250) );
  BUF_X1 U9 ( .A(N10), .Z(n252) );
  INV_X1 U10 ( .A(n1113), .ZN(n843) );
  INV_X1 U11 ( .A(n1102), .ZN(n842) );
  INV_X1 U12 ( .A(n1092), .ZN(n841) );
  INV_X1 U13 ( .A(n1082), .ZN(n840) );
  INV_X1 U14 ( .A(n1072), .ZN(n839) );
  INV_X1 U15 ( .A(n1062), .ZN(n838) );
  INV_X1 U16 ( .A(n1053), .ZN(n837) );
  INV_X1 U17 ( .A(n1044), .ZN(n836) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1105) );
  NOR3_X1 U19 ( .A1(N11), .A2(N12), .A3(n253), .ZN(n1094) );
  NAND2_X1 U20 ( .A1(n1104), .A2(n1136), .ZN(n1062) );
  NAND2_X1 U21 ( .A1(n1105), .A2(n1104), .ZN(n1113) );
  NAND2_X1 U22 ( .A1(n1094), .A2(n1104), .ZN(n1102) );
  NAND2_X1 U23 ( .A1(n1084), .A2(n1104), .ZN(n1092) );
  NAND2_X1 U24 ( .A1(n1074), .A2(n1104), .ZN(n1082) );
  NAND2_X1 U25 ( .A1(n1064), .A2(n1104), .ZN(n1072) );
  NAND2_X1 U26 ( .A1(n1104), .A2(n1125), .ZN(n1053) );
  NAND2_X1 U27 ( .A1(n1104), .A2(n1115), .ZN(n1044) );
  INV_X1 U28 ( .A(n1133), .ZN(n818) );
  INV_X1 U29 ( .A(n1123), .ZN(n817) );
  INV_X1 U30 ( .A(n889), .ZN(n816) );
  INV_X1 U31 ( .A(n880), .ZN(n815) );
  INV_X1 U32 ( .A(n871), .ZN(n814) );
  INV_X1 U33 ( .A(n862), .ZN(n813) );
  INV_X1 U34 ( .A(n853), .ZN(n812) );
  INV_X1 U35 ( .A(n989), .ZN(n830) );
  INV_X1 U36 ( .A(n980), .ZN(n829) );
  INV_X1 U37 ( .A(n971), .ZN(n828) );
  INV_X1 U38 ( .A(n916), .ZN(n822) );
  INV_X1 U39 ( .A(n907), .ZN(n821) );
  INV_X1 U40 ( .A(n898), .ZN(n820) );
  INV_X1 U41 ( .A(n1035), .ZN(n835) );
  INV_X1 U42 ( .A(n1025), .ZN(n834) );
  INV_X1 U43 ( .A(n1016), .ZN(n833) );
  INV_X1 U44 ( .A(n1007), .ZN(n832) );
  INV_X1 U45 ( .A(n998), .ZN(n831) );
  INV_X1 U46 ( .A(n962), .ZN(n827) );
  INV_X1 U47 ( .A(n952), .ZN(n826) );
  INV_X1 U48 ( .A(n943), .ZN(n825) );
  INV_X1 U49 ( .A(n934), .ZN(n824) );
  INV_X1 U50 ( .A(n925), .ZN(n823) );
  INV_X1 U51 ( .A(n1144), .ZN(n819) );
  BUF_X1 U52 ( .A(N11), .Z(n245) );
  BUF_X1 U53 ( .A(N11), .Z(n246) );
  INV_X1 U54 ( .A(N10), .ZN(n253) );
  BUF_X1 U55 ( .A(N12), .Z(n243) );
  NOR3_X1 U56 ( .A1(n255), .A2(N10), .A3(n254), .ZN(n1125) );
  NOR3_X1 U57 ( .A1(n255), .A2(n253), .A3(n254), .ZN(n1115) );
  NOR3_X1 U58 ( .A1(n253), .A2(N11), .A3(n255), .ZN(n1136) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n254), .ZN(n1084) );
  NOR3_X1 U60 ( .A1(n253), .A2(N12), .A3(n254), .ZN(n1074) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n255), .ZN(n1064) );
  NAND2_X1 U62 ( .A1(n1027), .A2(n1136), .ZN(n989) );
  NAND2_X1 U63 ( .A1(n954), .A2(n1136), .ZN(n916) );
  NAND2_X1 U64 ( .A1(n1027), .A2(n1064), .ZN(n998) );
  NAND2_X1 U65 ( .A1(n954), .A2(n1064), .ZN(n925) );
  NAND2_X1 U66 ( .A1(n1027), .A2(n1105), .ZN(n1035) );
  NAND2_X1 U67 ( .A1(n1027), .A2(n1094), .ZN(n1025) );
  NAND2_X1 U68 ( .A1(n954), .A2(n1105), .ZN(n962) );
  NAND2_X1 U69 ( .A1(n954), .A2(n1094), .ZN(n952) );
  NAND2_X1 U70 ( .A1(n1105), .A2(n1135), .ZN(n889) );
  NAND2_X1 U71 ( .A1(n1094), .A2(n1135), .ZN(n880) );
  NAND2_X1 U72 ( .A1(n1084), .A2(n1135), .ZN(n871) );
  NAND2_X1 U73 ( .A1(n1074), .A2(n1135), .ZN(n862) );
  NAND2_X1 U74 ( .A1(n1064), .A2(n1135), .ZN(n853) );
  NAND2_X1 U75 ( .A1(n1136), .A2(n1135), .ZN(n1144) );
  NAND2_X1 U76 ( .A1(n1125), .A2(n1135), .ZN(n1133) );
  NAND2_X1 U77 ( .A1(n1115), .A2(n1135), .ZN(n1123) );
  NAND2_X1 U78 ( .A1(n1027), .A2(n1084), .ZN(n1016) );
  NAND2_X1 U79 ( .A1(n1027), .A2(n1074), .ZN(n1007) );
  NAND2_X1 U80 ( .A1(n954), .A2(n1084), .ZN(n943) );
  NAND2_X1 U81 ( .A1(n954), .A2(n1074), .ZN(n934) );
  NAND2_X1 U82 ( .A1(n1027), .A2(n1125), .ZN(n980) );
  NAND2_X1 U83 ( .A1(n954), .A2(n1125), .ZN(n907) );
  NAND2_X1 U84 ( .A1(n1027), .A2(n1115), .ZN(n971) );
  NAND2_X1 U85 ( .A1(n954), .A2(n1115), .ZN(n898) );
  AND3_X1 U86 ( .A1(n844), .A2(n845), .A3(wr_en), .ZN(n1104) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1135) );
  AND3_X1 U88 ( .A1(N13), .A2(n845), .A3(wr_en), .ZN(n1027) );
  AND3_X1 U89 ( .A1(N14), .A2(n844), .A3(wr_en), .ZN(n954) );
  INV_X1 U90 ( .A(n1063), .ZN(n771) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n838), .B1(n1062), .B2(\mem[5][0] ), 
        .ZN(n1063) );
  INV_X1 U92 ( .A(n1061), .ZN(n770) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n838), .B1(n1062), .B2(\mem[5][1] ), 
        .ZN(n1061) );
  INV_X1 U94 ( .A(n1060), .ZN(n769) );
  AOI22_X1 U95 ( .A1(data_in[2]), .A2(n838), .B1(n1062), .B2(\mem[5][2] ), 
        .ZN(n1060) );
  INV_X1 U96 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U97 ( .A1(data_in[3]), .A2(n838), .B1(n1062), .B2(\mem[5][3] ), 
        .ZN(n1059) );
  INV_X1 U98 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U99 ( .A1(data_in[4]), .A2(n838), .B1(n1062), .B2(\mem[5][4] ), 
        .ZN(n1058) );
  INV_X1 U100 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U101 ( .A1(data_in[5]), .A2(n838), .B1(n1062), .B2(\mem[5][5] ), 
        .ZN(n1057) );
  INV_X1 U102 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U103 ( .A1(data_in[6]), .A2(n838), .B1(n1062), .B2(\mem[5][6] ), 
        .ZN(n1056) );
  INV_X1 U104 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U105 ( .A1(data_in[7]), .A2(n838), .B1(n1062), .B2(\mem[5][7] ), 
        .ZN(n1055) );
  INV_X1 U106 ( .A(n1026), .ZN(n739) );
  AOI22_X1 U107 ( .A1(data_in[0]), .A2(n834), .B1(n1025), .B2(\mem[9][0] ), 
        .ZN(n1026) );
  INV_X1 U108 ( .A(n1024), .ZN(n738) );
  AOI22_X1 U109 ( .A1(data_in[1]), .A2(n834), .B1(n1025), .B2(\mem[9][1] ), 
        .ZN(n1024) );
  INV_X1 U110 ( .A(n1023), .ZN(n737) );
  AOI22_X1 U111 ( .A1(data_in[2]), .A2(n834), .B1(n1025), .B2(\mem[9][2] ), 
        .ZN(n1023) );
  INV_X1 U112 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U113 ( .A1(data_in[3]), .A2(n834), .B1(n1025), .B2(\mem[9][3] ), 
        .ZN(n1022) );
  INV_X1 U114 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U115 ( .A1(data_in[4]), .A2(n834), .B1(n1025), .B2(\mem[9][4] ), 
        .ZN(n1021) );
  INV_X1 U116 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U117 ( .A1(data_in[5]), .A2(n834), .B1(n1025), .B2(\mem[9][5] ), 
        .ZN(n1020) );
  INV_X1 U118 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U119 ( .A1(data_in[6]), .A2(n834), .B1(n1025), .B2(\mem[9][6] ), 
        .ZN(n1019) );
  INV_X1 U120 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U121 ( .A1(data_in[7]), .A2(n834), .B1(n1025), .B2(\mem[9][7] ), 
        .ZN(n1018) );
  INV_X1 U122 ( .A(n990), .ZN(n707) );
  AOI22_X1 U123 ( .A1(data_in[0]), .A2(n830), .B1(n989), .B2(\mem[13][0] ), 
        .ZN(n990) );
  INV_X1 U124 ( .A(n988), .ZN(n706) );
  AOI22_X1 U125 ( .A1(data_in[1]), .A2(n830), .B1(n989), .B2(\mem[13][1] ), 
        .ZN(n988) );
  INV_X1 U126 ( .A(n987), .ZN(n705) );
  AOI22_X1 U127 ( .A1(data_in[2]), .A2(n830), .B1(n989), .B2(\mem[13][2] ), 
        .ZN(n987) );
  INV_X1 U128 ( .A(n986), .ZN(n704) );
  AOI22_X1 U129 ( .A1(data_in[3]), .A2(n830), .B1(n989), .B2(\mem[13][3] ), 
        .ZN(n986) );
  INV_X1 U130 ( .A(n985), .ZN(n703) );
  AOI22_X1 U131 ( .A1(data_in[4]), .A2(n830), .B1(n989), .B2(\mem[13][4] ), 
        .ZN(n985) );
  INV_X1 U132 ( .A(n984), .ZN(n702) );
  AOI22_X1 U133 ( .A1(data_in[5]), .A2(n830), .B1(n989), .B2(\mem[13][5] ), 
        .ZN(n984) );
  INV_X1 U134 ( .A(n983), .ZN(n701) );
  AOI22_X1 U135 ( .A1(data_in[6]), .A2(n830), .B1(n989), .B2(\mem[13][6] ), 
        .ZN(n983) );
  INV_X1 U136 ( .A(n982), .ZN(n700) );
  AOI22_X1 U137 ( .A1(data_in[7]), .A2(n830), .B1(n989), .B2(\mem[13][7] ), 
        .ZN(n982) );
  INV_X1 U138 ( .A(n953), .ZN(n675) );
  AOI22_X1 U139 ( .A1(data_in[0]), .A2(n826), .B1(n952), .B2(\mem[17][0] ), 
        .ZN(n953) );
  INV_X1 U140 ( .A(n915), .ZN(n642) );
  AOI22_X1 U141 ( .A1(data_in[1]), .A2(n822), .B1(n916), .B2(\mem[21][1] ), 
        .ZN(n915) );
  INV_X1 U142 ( .A(n914), .ZN(n641) );
  AOI22_X1 U143 ( .A1(data_in[2]), .A2(n822), .B1(n916), .B2(\mem[21][2] ), 
        .ZN(n914) );
  INV_X1 U144 ( .A(n913), .ZN(n640) );
  AOI22_X1 U145 ( .A1(data_in[3]), .A2(n822), .B1(n916), .B2(\mem[21][3] ), 
        .ZN(n913) );
  INV_X1 U146 ( .A(n912), .ZN(n639) );
  AOI22_X1 U147 ( .A1(data_in[4]), .A2(n822), .B1(n916), .B2(\mem[21][4] ), 
        .ZN(n912) );
  INV_X1 U148 ( .A(n911), .ZN(n638) );
  AOI22_X1 U149 ( .A1(data_in[5]), .A2(n822), .B1(n916), .B2(\mem[21][5] ), 
        .ZN(n911) );
  INV_X1 U150 ( .A(n910), .ZN(n637) );
  AOI22_X1 U151 ( .A1(data_in[6]), .A2(n822), .B1(n916), .B2(\mem[21][6] ), 
        .ZN(n910) );
  INV_X1 U152 ( .A(n909), .ZN(n636) );
  AOI22_X1 U153 ( .A1(data_in[7]), .A2(n822), .B1(n916), .B2(\mem[21][7] ), 
        .ZN(n909) );
  INV_X1 U154 ( .A(n951), .ZN(n674) );
  AOI22_X1 U155 ( .A1(data_in[1]), .A2(n826), .B1(n952), .B2(\mem[17][1] ), 
        .ZN(n951) );
  INV_X1 U156 ( .A(n950), .ZN(n673) );
  AOI22_X1 U157 ( .A1(data_in[2]), .A2(n826), .B1(n952), .B2(\mem[17][2] ), 
        .ZN(n950) );
  INV_X1 U158 ( .A(n949), .ZN(n672) );
  AOI22_X1 U159 ( .A1(data_in[3]), .A2(n826), .B1(n952), .B2(\mem[17][3] ), 
        .ZN(n949) );
  INV_X1 U160 ( .A(n948), .ZN(n671) );
  AOI22_X1 U161 ( .A1(data_in[4]), .A2(n826), .B1(n952), .B2(\mem[17][4] ), 
        .ZN(n948) );
  INV_X1 U162 ( .A(n947), .ZN(n670) );
  AOI22_X1 U163 ( .A1(data_in[5]), .A2(n826), .B1(n952), .B2(\mem[17][5] ), 
        .ZN(n947) );
  INV_X1 U164 ( .A(n946), .ZN(n669) );
  AOI22_X1 U165 ( .A1(data_in[6]), .A2(n826), .B1(n952), .B2(\mem[17][6] ), 
        .ZN(n946) );
  INV_X1 U166 ( .A(n945), .ZN(n668) );
  AOI22_X1 U167 ( .A1(data_in[7]), .A2(n826), .B1(n952), .B2(\mem[17][7] ), 
        .ZN(n945) );
  INV_X1 U168 ( .A(n917), .ZN(n643) );
  AOI22_X1 U169 ( .A1(data_in[0]), .A2(n822), .B1(n916), .B2(\mem[21][0] ), 
        .ZN(n917) );
  INV_X1 U170 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U171 ( .A1(data_in[0]), .A2(n837), .B1(n1053), .B2(\mem[6][0] ), 
        .ZN(n1054) );
  INV_X1 U172 ( .A(n1052), .ZN(n762) );
  AOI22_X1 U173 ( .A1(data_in[1]), .A2(n837), .B1(n1053), .B2(\mem[6][1] ), 
        .ZN(n1052) );
  INV_X1 U174 ( .A(n1051), .ZN(n761) );
  AOI22_X1 U175 ( .A1(data_in[2]), .A2(n837), .B1(n1053), .B2(\mem[6][2] ), 
        .ZN(n1051) );
  INV_X1 U176 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U177 ( .A1(data_in[3]), .A2(n837), .B1(n1053), .B2(\mem[6][3] ), 
        .ZN(n1050) );
  INV_X1 U178 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U179 ( .A1(data_in[4]), .A2(n837), .B1(n1053), .B2(\mem[6][4] ), 
        .ZN(n1049) );
  INV_X1 U180 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U181 ( .A1(data_in[5]), .A2(n837), .B1(n1053), .B2(\mem[6][5] ), 
        .ZN(n1048) );
  INV_X1 U182 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U183 ( .A1(data_in[6]), .A2(n837), .B1(n1053), .B2(\mem[6][6] ), 
        .ZN(n1047) );
  INV_X1 U184 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U185 ( .A1(data_in[7]), .A2(n837), .B1(n1053), .B2(\mem[6][7] ), 
        .ZN(n1046) );
  INV_X1 U186 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U187 ( .A1(data_in[0]), .A2(n836), .B1(n1044), .B2(\mem[7][0] ), 
        .ZN(n1045) );
  INV_X1 U188 ( .A(n1043), .ZN(n754) );
  AOI22_X1 U189 ( .A1(data_in[1]), .A2(n836), .B1(n1044), .B2(\mem[7][1] ), 
        .ZN(n1043) );
  INV_X1 U190 ( .A(n1042), .ZN(n753) );
  AOI22_X1 U191 ( .A1(data_in[2]), .A2(n836), .B1(n1044), .B2(\mem[7][2] ), 
        .ZN(n1042) );
  INV_X1 U192 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U193 ( .A1(data_in[3]), .A2(n836), .B1(n1044), .B2(\mem[7][3] ), 
        .ZN(n1041) );
  INV_X1 U194 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U195 ( .A1(data_in[4]), .A2(n836), .B1(n1044), .B2(\mem[7][4] ), 
        .ZN(n1040) );
  INV_X1 U196 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U197 ( .A1(data_in[5]), .A2(n836), .B1(n1044), .B2(\mem[7][5] ), 
        .ZN(n1039) );
  INV_X1 U198 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U199 ( .A1(data_in[6]), .A2(n836), .B1(n1044), .B2(\mem[7][6] ), 
        .ZN(n1038) );
  INV_X1 U200 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U201 ( .A1(data_in[7]), .A2(n836), .B1(n1044), .B2(\mem[7][7] ), 
        .ZN(n1037) );
  INV_X1 U202 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U203 ( .A1(data_in[0]), .A2(n833), .B1(n1016), .B2(\mem[10][0] ), 
        .ZN(n1017) );
  INV_X1 U204 ( .A(n1015), .ZN(n730) );
  AOI22_X1 U205 ( .A1(data_in[1]), .A2(n833), .B1(n1016), .B2(\mem[10][1] ), 
        .ZN(n1015) );
  INV_X1 U206 ( .A(n1014), .ZN(n729) );
  AOI22_X1 U207 ( .A1(data_in[2]), .A2(n833), .B1(n1016), .B2(\mem[10][2] ), 
        .ZN(n1014) );
  INV_X1 U208 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U209 ( .A1(data_in[3]), .A2(n833), .B1(n1016), .B2(\mem[10][3] ), 
        .ZN(n1013) );
  INV_X1 U210 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U211 ( .A1(data_in[4]), .A2(n833), .B1(n1016), .B2(\mem[10][4] ), 
        .ZN(n1012) );
  INV_X1 U212 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U213 ( .A1(data_in[5]), .A2(n833), .B1(n1016), .B2(\mem[10][5] ), 
        .ZN(n1011) );
  INV_X1 U214 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U215 ( .A1(data_in[6]), .A2(n833), .B1(n1016), .B2(\mem[10][6] ), 
        .ZN(n1010) );
  INV_X1 U216 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U217 ( .A1(data_in[7]), .A2(n833), .B1(n1016), .B2(\mem[10][7] ), 
        .ZN(n1009) );
  INV_X1 U218 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U219 ( .A1(data_in[0]), .A2(n832), .B1(n1007), .B2(\mem[11][0] ), 
        .ZN(n1008) );
  INV_X1 U220 ( .A(n1006), .ZN(n722) );
  AOI22_X1 U221 ( .A1(data_in[1]), .A2(n832), .B1(n1007), .B2(\mem[11][1] ), 
        .ZN(n1006) );
  INV_X1 U222 ( .A(n1005), .ZN(n721) );
  AOI22_X1 U223 ( .A1(data_in[2]), .A2(n832), .B1(n1007), .B2(\mem[11][2] ), 
        .ZN(n1005) );
  INV_X1 U224 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U225 ( .A1(data_in[3]), .A2(n832), .B1(n1007), .B2(\mem[11][3] ), 
        .ZN(n1004) );
  INV_X1 U226 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U227 ( .A1(data_in[4]), .A2(n832), .B1(n1007), .B2(\mem[11][4] ), 
        .ZN(n1003) );
  INV_X1 U228 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U229 ( .A1(data_in[5]), .A2(n832), .B1(n1007), .B2(\mem[11][5] ), 
        .ZN(n1002) );
  INV_X1 U230 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U231 ( .A1(data_in[6]), .A2(n832), .B1(n1007), .B2(\mem[11][6] ), 
        .ZN(n1001) );
  INV_X1 U232 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U233 ( .A1(data_in[7]), .A2(n832), .B1(n1007), .B2(\mem[11][7] ), 
        .ZN(n1000) );
  INV_X1 U234 ( .A(n981), .ZN(n699) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n829), .B1(n980), .B2(\mem[14][0] ), 
        .ZN(n981) );
  INV_X1 U236 ( .A(n979), .ZN(n698) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n829), .B1(n980), .B2(\mem[14][1] ), 
        .ZN(n979) );
  INV_X1 U238 ( .A(n978), .ZN(n697) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n829), .B1(n980), .B2(\mem[14][2] ), 
        .ZN(n978) );
  INV_X1 U240 ( .A(n977), .ZN(n696) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n829), .B1(n980), .B2(\mem[14][3] ), 
        .ZN(n977) );
  INV_X1 U242 ( .A(n976), .ZN(n695) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n829), .B1(n980), .B2(\mem[14][4] ), 
        .ZN(n976) );
  INV_X1 U244 ( .A(n975), .ZN(n694) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n829), .B1(n980), .B2(\mem[14][5] ), 
        .ZN(n975) );
  INV_X1 U246 ( .A(n974), .ZN(n693) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n829), .B1(n980), .B2(\mem[14][6] ), 
        .ZN(n974) );
  INV_X1 U248 ( .A(n973), .ZN(n692) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n829), .B1(n980), .B2(\mem[14][7] ), 
        .ZN(n973) );
  INV_X1 U250 ( .A(n972), .ZN(n691) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n828), .B1(n971), .B2(\mem[15][0] ), 
        .ZN(n972) );
  INV_X1 U252 ( .A(n970), .ZN(n690) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n828), .B1(n971), .B2(\mem[15][1] ), 
        .ZN(n970) );
  INV_X1 U254 ( .A(n969), .ZN(n689) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n828), .B1(n971), .B2(\mem[15][2] ), 
        .ZN(n969) );
  INV_X1 U256 ( .A(n968), .ZN(n688) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n828), .B1(n971), .B2(\mem[15][3] ), 
        .ZN(n968) );
  INV_X1 U258 ( .A(n967), .ZN(n687) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n828), .B1(n971), .B2(\mem[15][4] ), 
        .ZN(n967) );
  INV_X1 U260 ( .A(n966), .ZN(n686) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n828), .B1(n971), .B2(\mem[15][5] ), 
        .ZN(n966) );
  INV_X1 U262 ( .A(n965), .ZN(n685) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n828), .B1(n971), .B2(\mem[15][6] ), 
        .ZN(n965) );
  INV_X1 U264 ( .A(n964), .ZN(n684) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n828), .B1(n971), .B2(\mem[15][7] ), 
        .ZN(n964) );
  INV_X1 U266 ( .A(n944), .ZN(n667) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n825), .B1(n943), .B2(\mem[18][0] ), 
        .ZN(n944) );
  INV_X1 U268 ( .A(n942), .ZN(n666) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n825), .B1(n943), .B2(\mem[18][1] ), 
        .ZN(n942) );
  INV_X1 U270 ( .A(n941), .ZN(n665) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n825), .B1(n943), .B2(\mem[18][2] ), 
        .ZN(n941) );
  INV_X1 U272 ( .A(n940), .ZN(n664) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n825), .B1(n943), .B2(\mem[18][3] ), 
        .ZN(n940) );
  INV_X1 U274 ( .A(n939), .ZN(n663) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n825), .B1(n943), .B2(\mem[18][4] ), 
        .ZN(n939) );
  INV_X1 U276 ( .A(n938), .ZN(n662) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n825), .B1(n943), .B2(\mem[18][5] ), 
        .ZN(n938) );
  INV_X1 U278 ( .A(n937), .ZN(n661) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n825), .B1(n943), .B2(\mem[18][6] ), 
        .ZN(n937) );
  INV_X1 U280 ( .A(n936), .ZN(n660) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n825), .B1(n943), .B2(\mem[18][7] ), 
        .ZN(n936) );
  INV_X1 U282 ( .A(n935), .ZN(n659) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n824), .B1(n934), .B2(\mem[19][0] ), 
        .ZN(n935) );
  INV_X1 U284 ( .A(n933), .ZN(n658) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n824), .B1(n934), .B2(\mem[19][1] ), 
        .ZN(n933) );
  INV_X1 U286 ( .A(n932), .ZN(n657) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n824), .B1(n934), .B2(\mem[19][2] ), 
        .ZN(n932) );
  INV_X1 U288 ( .A(n931), .ZN(n656) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n824), .B1(n934), .B2(\mem[19][3] ), 
        .ZN(n931) );
  INV_X1 U290 ( .A(n930), .ZN(n655) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n824), .B1(n934), .B2(\mem[19][4] ), 
        .ZN(n930) );
  INV_X1 U292 ( .A(n929), .ZN(n654) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n824), .B1(n934), .B2(\mem[19][5] ), 
        .ZN(n929) );
  INV_X1 U294 ( .A(n928), .ZN(n653) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n824), .B1(n934), .B2(\mem[19][6] ), 
        .ZN(n928) );
  INV_X1 U296 ( .A(n927), .ZN(n652) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n824), .B1(n934), .B2(\mem[19][7] ), 
        .ZN(n927) );
  INV_X1 U298 ( .A(n908), .ZN(n635) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n821), .B1(n907), .B2(\mem[22][0] ), 
        .ZN(n908) );
  INV_X1 U300 ( .A(n906), .ZN(n634) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n821), .B1(n907), .B2(\mem[22][1] ), 
        .ZN(n906) );
  INV_X1 U302 ( .A(n905), .ZN(n633) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n821), .B1(n907), .B2(\mem[22][2] ), 
        .ZN(n905) );
  INV_X1 U304 ( .A(n904), .ZN(n632) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n821), .B1(n907), .B2(\mem[22][3] ), 
        .ZN(n904) );
  INV_X1 U306 ( .A(n903), .ZN(n631) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n821), .B1(n907), .B2(\mem[22][4] ), 
        .ZN(n903) );
  INV_X1 U308 ( .A(n902), .ZN(n630) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n821), .B1(n907), .B2(\mem[22][5] ), 
        .ZN(n902) );
  INV_X1 U310 ( .A(n901), .ZN(n629) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n821), .B1(n907), .B2(\mem[22][6] ), 
        .ZN(n901) );
  INV_X1 U312 ( .A(n900), .ZN(n628) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n821), .B1(n907), .B2(\mem[22][7] ), 
        .ZN(n900) );
  INV_X1 U314 ( .A(n899), .ZN(n627) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n820), .B1(n898), .B2(\mem[23][0] ), 
        .ZN(n899) );
  INV_X1 U316 ( .A(n897), .ZN(n626) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n820), .B1(n898), .B2(\mem[23][1] ), 
        .ZN(n897) );
  INV_X1 U318 ( .A(n896), .ZN(n625) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n820), .B1(n898), .B2(\mem[23][2] ), 
        .ZN(n896) );
  INV_X1 U320 ( .A(n895), .ZN(n624) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n820), .B1(n898), .B2(\mem[23][3] ), 
        .ZN(n895) );
  INV_X1 U322 ( .A(n894), .ZN(n623) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n820), .B1(n898), .B2(\mem[23][4] ), 
        .ZN(n894) );
  INV_X1 U324 ( .A(n893), .ZN(n622) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n820), .B1(n898), .B2(\mem[23][5] ), 
        .ZN(n893) );
  INV_X1 U326 ( .A(n892), .ZN(n621) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n820), .B1(n898), .B2(\mem[23][6] ), 
        .ZN(n892) );
  INV_X1 U328 ( .A(n891), .ZN(n620) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n820), .B1(n898), .B2(\mem[23][7] ), 
        .ZN(n891) );
  INV_X1 U330 ( .A(N12), .ZN(n255) );
  INV_X1 U331 ( .A(N11), .ZN(n254) );
  INV_X1 U332 ( .A(n999), .ZN(n715) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n831), .B1(n998), .B2(\mem[12][0] ), 
        .ZN(n999) );
  INV_X1 U334 ( .A(n997), .ZN(n714) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n831), .B1(n998), .B2(\mem[12][1] ), 
        .ZN(n997) );
  INV_X1 U336 ( .A(n996), .ZN(n713) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n831), .B1(n998), .B2(\mem[12][2] ), 
        .ZN(n996) );
  INV_X1 U338 ( .A(n995), .ZN(n712) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n831), .B1(n998), .B2(\mem[12][3] ), 
        .ZN(n995) );
  INV_X1 U340 ( .A(n994), .ZN(n711) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n831), .B1(n998), .B2(\mem[12][4] ), 
        .ZN(n994) );
  INV_X1 U342 ( .A(n993), .ZN(n710) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n831), .B1(n998), .B2(\mem[12][5] ), 
        .ZN(n993) );
  INV_X1 U344 ( .A(n992), .ZN(n709) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n831), .B1(n998), .B2(\mem[12][6] ), 
        .ZN(n992) );
  INV_X1 U346 ( .A(n991), .ZN(n708) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n831), .B1(n998), .B2(\mem[12][7] ), 
        .ZN(n991) );
  INV_X1 U348 ( .A(n926), .ZN(n651) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n823), .B1(n925), .B2(\mem[20][0] ), 
        .ZN(n926) );
  INV_X1 U350 ( .A(n924), .ZN(n650) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n823), .B1(n925), .B2(\mem[20][1] ), 
        .ZN(n924) );
  INV_X1 U352 ( .A(n923), .ZN(n649) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n823), .B1(n925), .B2(\mem[20][2] ), 
        .ZN(n923) );
  INV_X1 U354 ( .A(n922), .ZN(n648) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n823), .B1(n925), .B2(\mem[20][3] ), 
        .ZN(n922) );
  INV_X1 U356 ( .A(n921), .ZN(n647) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n823), .B1(n925), .B2(\mem[20][4] ), 
        .ZN(n921) );
  INV_X1 U358 ( .A(n920), .ZN(n646) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n823), .B1(n925), .B2(\mem[20][5] ), 
        .ZN(n920) );
  INV_X1 U360 ( .A(n919), .ZN(n645) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n823), .B1(n925), .B2(\mem[20][6] ), 
        .ZN(n919) );
  INV_X1 U362 ( .A(n918), .ZN(n644) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n823), .B1(n925), .B2(\mem[20][7] ), 
        .ZN(n918) );
  INV_X1 U364 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n835), .B1(n1035), .B2(\mem[8][0] ), 
        .ZN(n1036) );
  INV_X1 U366 ( .A(n1034), .ZN(n746) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n835), .B1(n1035), .B2(\mem[8][1] ), 
        .ZN(n1034) );
  INV_X1 U368 ( .A(n1033), .ZN(n745) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n835), .B1(n1035), .B2(\mem[8][2] ), 
        .ZN(n1033) );
  INV_X1 U370 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n835), .B1(n1035), .B2(\mem[8][3] ), 
        .ZN(n1032) );
  INV_X1 U372 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n835), .B1(n1035), .B2(\mem[8][4] ), 
        .ZN(n1031) );
  INV_X1 U374 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n835), .B1(n1035), .B2(\mem[8][5] ), 
        .ZN(n1030) );
  INV_X1 U376 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n835), .B1(n1035), .B2(\mem[8][6] ), 
        .ZN(n1029) );
  INV_X1 U378 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n835), .B1(n1035), .B2(\mem[8][7] ), 
        .ZN(n1028) );
  INV_X1 U380 ( .A(n963), .ZN(n683) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n827), .B1(n962), .B2(\mem[16][0] ), 
        .ZN(n963) );
  INV_X1 U382 ( .A(n961), .ZN(n682) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n827), .B1(n962), .B2(\mem[16][1] ), 
        .ZN(n961) );
  INV_X1 U384 ( .A(n960), .ZN(n681) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n827), .B1(n962), .B2(\mem[16][2] ), 
        .ZN(n960) );
  INV_X1 U386 ( .A(n959), .ZN(n680) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n827), .B1(n962), .B2(\mem[16][3] ), 
        .ZN(n959) );
  INV_X1 U388 ( .A(n958), .ZN(n679) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n827), .B1(n962), .B2(\mem[16][4] ), 
        .ZN(n958) );
  INV_X1 U390 ( .A(n957), .ZN(n678) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n827), .B1(n962), .B2(\mem[16][5] ), 
        .ZN(n957) );
  INV_X1 U392 ( .A(n956), .ZN(n677) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n827), .B1(n962), .B2(\mem[16][6] ), 
        .ZN(n956) );
  INV_X1 U394 ( .A(n955), .ZN(n676) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n827), .B1(n962), .B2(\mem[16][7] ), 
        .ZN(n955) );
  INV_X1 U396 ( .A(n890), .ZN(n619) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n816), .B1(n889), .B2(\mem[24][0] ), 
        .ZN(n890) );
  INV_X1 U398 ( .A(n888), .ZN(n618) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n816), .B1(n889), .B2(\mem[24][1] ), 
        .ZN(n888) );
  INV_X1 U400 ( .A(n887), .ZN(n617) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n816), .B1(n889), .B2(\mem[24][2] ), 
        .ZN(n887) );
  INV_X1 U402 ( .A(n886), .ZN(n616) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n816), .B1(n889), .B2(\mem[24][3] ), 
        .ZN(n886) );
  INV_X1 U404 ( .A(n885), .ZN(n615) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n816), .B1(n889), .B2(\mem[24][4] ), 
        .ZN(n885) );
  INV_X1 U406 ( .A(n884), .ZN(n614) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n816), .B1(n889), .B2(\mem[24][5] ), 
        .ZN(n884) );
  INV_X1 U408 ( .A(n883), .ZN(n613) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n816), .B1(n889), .B2(\mem[24][6] ), 
        .ZN(n883) );
  INV_X1 U410 ( .A(n882), .ZN(n612) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n816), .B1(n889), .B2(\mem[24][7] ), 
        .ZN(n882) );
  INV_X1 U412 ( .A(n881), .ZN(n611) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n815), .B1(n880), .B2(\mem[25][0] ), 
        .ZN(n881) );
  INV_X1 U414 ( .A(n879), .ZN(n610) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n815), .B1(n880), .B2(\mem[25][1] ), 
        .ZN(n879) );
  INV_X1 U416 ( .A(n878), .ZN(n609) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n815), .B1(n880), .B2(\mem[25][2] ), 
        .ZN(n878) );
  INV_X1 U418 ( .A(n877), .ZN(n608) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n815), .B1(n880), .B2(\mem[25][3] ), 
        .ZN(n877) );
  INV_X1 U420 ( .A(n876), .ZN(n607) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n815), .B1(n880), .B2(\mem[25][4] ), 
        .ZN(n876) );
  INV_X1 U422 ( .A(n875), .ZN(n606) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n815), .B1(n880), .B2(\mem[25][5] ), 
        .ZN(n875) );
  INV_X1 U424 ( .A(n874), .ZN(n605) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n815), .B1(n880), .B2(\mem[25][6] ), 
        .ZN(n874) );
  INV_X1 U426 ( .A(n873), .ZN(n604) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n815), .B1(n880), .B2(\mem[25][7] ), 
        .ZN(n873) );
  INV_X1 U428 ( .A(n872), .ZN(n603) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n814), .B1(n871), .B2(\mem[26][0] ), 
        .ZN(n872) );
  INV_X1 U430 ( .A(n870), .ZN(n602) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n814), .B1(n871), .B2(\mem[26][1] ), 
        .ZN(n870) );
  INV_X1 U432 ( .A(n869), .ZN(n601) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n814), .B1(n871), .B2(\mem[26][2] ), 
        .ZN(n869) );
  INV_X1 U434 ( .A(n868), .ZN(n600) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n814), .B1(n871), .B2(\mem[26][3] ), 
        .ZN(n868) );
  INV_X1 U436 ( .A(n867), .ZN(n599) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n814), .B1(n871), .B2(\mem[26][4] ), 
        .ZN(n867) );
  INV_X1 U438 ( .A(n866), .ZN(n598) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n814), .B1(n871), .B2(\mem[26][5] ), 
        .ZN(n866) );
  INV_X1 U440 ( .A(n865), .ZN(n597) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n814), .B1(n871), .B2(\mem[26][6] ), 
        .ZN(n865) );
  INV_X1 U442 ( .A(n864), .ZN(n596) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n814), .B1(n871), .B2(\mem[26][7] ), 
        .ZN(n864) );
  INV_X1 U444 ( .A(n863), .ZN(n595) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n813), .B1(n862), .B2(\mem[27][0] ), 
        .ZN(n863) );
  INV_X1 U446 ( .A(n861), .ZN(n594) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n813), .B1(n862), .B2(\mem[27][1] ), 
        .ZN(n861) );
  INV_X1 U448 ( .A(n860), .ZN(n293) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n813), .B1(n862), .B2(\mem[27][2] ), 
        .ZN(n860) );
  INV_X1 U450 ( .A(n859), .ZN(n292) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n813), .B1(n862), .B2(\mem[27][3] ), 
        .ZN(n859) );
  INV_X1 U452 ( .A(n858), .ZN(n291) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n813), .B1(n862), .B2(\mem[27][4] ), 
        .ZN(n858) );
  INV_X1 U454 ( .A(n857), .ZN(n290) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n813), .B1(n862), .B2(\mem[27][5] ), 
        .ZN(n857) );
  INV_X1 U456 ( .A(n856), .ZN(n289) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n813), .B1(n862), .B2(\mem[27][6] ), 
        .ZN(n856) );
  INV_X1 U458 ( .A(n855), .ZN(n288) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n813), .B1(n862), .B2(\mem[27][7] ), 
        .ZN(n855) );
  INV_X1 U460 ( .A(n854), .ZN(n287) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n812), .B1(n853), .B2(\mem[28][0] ), 
        .ZN(n854) );
  INV_X1 U462 ( .A(n852), .ZN(n286) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n812), .B1(n853), .B2(\mem[28][1] ), 
        .ZN(n852) );
  INV_X1 U464 ( .A(n851), .ZN(n285) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n812), .B1(n853), .B2(\mem[28][2] ), 
        .ZN(n851) );
  INV_X1 U466 ( .A(n850), .ZN(n284) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n812), .B1(n853), .B2(\mem[28][3] ), 
        .ZN(n850) );
  INV_X1 U468 ( .A(n849), .ZN(n283) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n812), .B1(n853), .B2(\mem[28][4] ), 
        .ZN(n849) );
  INV_X1 U470 ( .A(n848), .ZN(n282) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n812), .B1(n853), .B2(\mem[28][5] ), 
        .ZN(n848) );
  INV_X1 U472 ( .A(n847), .ZN(n281) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n812), .B1(n853), .B2(\mem[28][6] ), 
        .ZN(n847) );
  INV_X1 U474 ( .A(n846), .ZN(n280) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n812), .B1(n853), .B2(\mem[28][7] ), 
        .ZN(n846) );
  INV_X1 U476 ( .A(n1145), .ZN(n279) );
  AOI22_X1 U477 ( .A1(n819), .A2(data_in[0]), .B1(n1144), .B2(\mem[29][0] ), 
        .ZN(n1145) );
  INV_X1 U478 ( .A(n1143), .ZN(n278) );
  AOI22_X1 U479 ( .A1(n819), .A2(data_in[1]), .B1(n1144), .B2(\mem[29][1] ), 
        .ZN(n1143) );
  INV_X1 U480 ( .A(n1142), .ZN(n277) );
  AOI22_X1 U481 ( .A1(n819), .A2(data_in[2]), .B1(n1144), .B2(\mem[29][2] ), 
        .ZN(n1142) );
  INV_X1 U482 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U483 ( .A1(n819), .A2(data_in[3]), .B1(n1144), .B2(\mem[29][3] ), 
        .ZN(n1141) );
  INV_X1 U484 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U485 ( .A1(n819), .A2(data_in[4]), .B1(n1144), .B2(\mem[29][4] ), 
        .ZN(n1140) );
  INV_X1 U486 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U487 ( .A1(n819), .A2(data_in[5]), .B1(n1144), .B2(\mem[29][5] ), 
        .ZN(n1139) );
  INV_X1 U488 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U489 ( .A1(n819), .A2(data_in[6]), .B1(n1144), .B2(\mem[29][6] ), 
        .ZN(n1138) );
  INV_X1 U490 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U491 ( .A1(n819), .A2(data_in[7]), .B1(n1144), .B2(\mem[29][7] ), 
        .ZN(n1137) );
  INV_X1 U492 ( .A(n1134), .ZN(n271) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n818), .B1(n1133), .B2(\mem[30][0] ), 
        .ZN(n1134) );
  INV_X1 U494 ( .A(n1132), .ZN(n270) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n818), .B1(n1133), .B2(\mem[30][1] ), 
        .ZN(n1132) );
  INV_X1 U496 ( .A(n1131), .ZN(n269) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n818), .B1(n1133), .B2(\mem[30][2] ), 
        .ZN(n1131) );
  INV_X1 U498 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n818), .B1(n1133), .B2(\mem[30][3] ), 
        .ZN(n1130) );
  INV_X1 U500 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n818), .B1(n1133), .B2(\mem[30][4] ), 
        .ZN(n1129) );
  INV_X1 U502 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n818), .B1(n1133), .B2(\mem[30][5] ), 
        .ZN(n1128) );
  INV_X1 U504 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n818), .B1(n1133), .B2(\mem[30][6] ), 
        .ZN(n1127) );
  INV_X1 U506 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n818), .B1(n1133), .B2(\mem[30][7] ), 
        .ZN(n1126) );
  INV_X1 U508 ( .A(n1124), .ZN(n263) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n817), .B1(n1123), .B2(\mem[31][0] ), 
        .ZN(n1124) );
  INV_X1 U510 ( .A(n1122), .ZN(n262) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n817), .B1(n1123), .B2(\mem[31][1] ), 
        .ZN(n1122) );
  INV_X1 U512 ( .A(n1121), .ZN(n261) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n817), .B1(n1123), .B2(\mem[31][2] ), 
        .ZN(n1121) );
  INV_X1 U514 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n817), .B1(n1123), .B2(\mem[31][3] ), 
        .ZN(n1120) );
  INV_X1 U516 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n817), .B1(n1123), .B2(\mem[31][4] ), 
        .ZN(n1119) );
  INV_X1 U518 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n817), .B1(n1123), .B2(\mem[31][5] ), 
        .ZN(n1118) );
  INV_X1 U520 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n817), .B1(n1123), .B2(\mem[31][6] ), 
        .ZN(n1117) );
  INV_X1 U522 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n817), .B1(n1123), .B2(\mem[31][7] ), 
        .ZN(n1116) );
  INV_X1 U524 ( .A(n1114), .ZN(n811) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n843), .B1(n1113), .B2(\mem[0][0] ), 
        .ZN(n1114) );
  INV_X1 U526 ( .A(n1112), .ZN(n810) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n843), .B1(n1113), .B2(\mem[0][1] ), 
        .ZN(n1112) );
  INV_X1 U528 ( .A(n1111), .ZN(n809) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n843), .B1(n1113), .B2(\mem[0][2] ), 
        .ZN(n1111) );
  INV_X1 U530 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n843), .B1(n1113), .B2(\mem[0][3] ), 
        .ZN(n1110) );
  INV_X1 U532 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n843), .B1(n1113), .B2(\mem[0][4] ), 
        .ZN(n1109) );
  INV_X1 U534 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n843), .B1(n1113), .B2(\mem[0][5] ), 
        .ZN(n1108) );
  INV_X1 U536 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n843), .B1(n1113), .B2(\mem[0][6] ), 
        .ZN(n1107) );
  INV_X1 U538 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n843), .B1(n1113), .B2(\mem[0][7] ), 
        .ZN(n1106) );
  INV_X1 U540 ( .A(n1103), .ZN(n803) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[1][0] ), 
        .ZN(n1103) );
  INV_X1 U542 ( .A(n1101), .ZN(n802) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[1][1] ), 
        .ZN(n1101) );
  INV_X1 U544 ( .A(n1100), .ZN(n801) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[1][2] ), 
        .ZN(n1100) );
  INV_X1 U546 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[1][3] ), 
        .ZN(n1099) );
  INV_X1 U548 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[1][4] ), 
        .ZN(n1098) );
  INV_X1 U550 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[1][5] ), 
        .ZN(n1097) );
  INV_X1 U552 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[1][6] ), 
        .ZN(n1096) );
  INV_X1 U554 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[1][7] ), 
        .ZN(n1095) );
  INV_X1 U556 ( .A(n1093), .ZN(n795) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n841), .B1(n1092), .B2(\mem[2][0] ), 
        .ZN(n1093) );
  INV_X1 U558 ( .A(n1091), .ZN(n794) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n841), .B1(n1092), .B2(\mem[2][1] ), 
        .ZN(n1091) );
  INV_X1 U560 ( .A(n1090), .ZN(n793) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n841), .B1(n1092), .B2(\mem[2][2] ), 
        .ZN(n1090) );
  INV_X1 U562 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n841), .B1(n1092), .B2(\mem[2][3] ), 
        .ZN(n1089) );
  INV_X1 U564 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n841), .B1(n1092), .B2(\mem[2][4] ), 
        .ZN(n1088) );
  INV_X1 U566 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n841), .B1(n1092), .B2(\mem[2][5] ), 
        .ZN(n1087) );
  INV_X1 U568 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n841), .B1(n1092), .B2(\mem[2][6] ), 
        .ZN(n1086) );
  INV_X1 U570 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n841), .B1(n1092), .B2(\mem[2][7] ), 
        .ZN(n1085) );
  INV_X1 U572 ( .A(n1083), .ZN(n787) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n840), .B1(n1082), .B2(\mem[3][0] ), 
        .ZN(n1083) );
  INV_X1 U574 ( .A(n1081), .ZN(n786) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n840), .B1(n1082), .B2(\mem[3][1] ), 
        .ZN(n1081) );
  INV_X1 U576 ( .A(n1080), .ZN(n785) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n840), .B1(n1082), .B2(\mem[3][2] ), 
        .ZN(n1080) );
  INV_X1 U578 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n840), .B1(n1082), .B2(\mem[3][3] ), 
        .ZN(n1079) );
  INV_X1 U580 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n840), .B1(n1082), .B2(\mem[3][4] ), 
        .ZN(n1078) );
  INV_X1 U582 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n840), .B1(n1082), .B2(\mem[3][5] ), 
        .ZN(n1077) );
  INV_X1 U584 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n840), .B1(n1082), .B2(\mem[3][6] ), 
        .ZN(n1076) );
  INV_X1 U586 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n840), .B1(n1082), .B2(\mem[3][7] ), 
        .ZN(n1075) );
  INV_X1 U588 ( .A(n1073), .ZN(n779) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n839), .B1(n1072), .B2(\mem[4][0] ), 
        .ZN(n1073) );
  INV_X1 U590 ( .A(n1071), .ZN(n778) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n839), .B1(n1072), .B2(\mem[4][1] ), 
        .ZN(n1071) );
  INV_X1 U592 ( .A(n1070), .ZN(n777) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n839), .B1(n1072), .B2(\mem[4][2] ), 
        .ZN(n1070) );
  INV_X1 U594 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n839), .B1(n1072), .B2(\mem[4][3] ), 
        .ZN(n1069) );
  INV_X1 U596 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n839), .B1(n1072), .B2(\mem[4][4] ), 
        .ZN(n1068) );
  INV_X1 U598 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n839), .B1(n1072), .B2(\mem[4][5] ), 
        .ZN(n1067) );
  INV_X1 U600 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n839), .B1(n1072), .B2(\mem[4][6] ), 
        .ZN(n1066) );
  INV_X1 U602 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n839), .B1(n1072), .B2(\mem[4][7] ), 
        .ZN(n1065) );
  INV_X1 U604 ( .A(N13), .ZN(n844) );
  INV_X1 U605 ( .A(N14), .ZN(n845) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n251), .Z(n3) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n248), .Z(n4) );
  MUX2_X1 U608 ( .A(n4), .B(n3), .S(n244), .Z(n5) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n251), .Z(n6) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n251), .Z(n7) );
  MUX2_X1 U611 ( .A(n7), .B(n6), .S(n244), .Z(n8) );
  MUX2_X1 U612 ( .A(n8), .B(n5), .S(n243), .Z(n9) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n252), .Z(n10) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n250), .Z(n11) );
  MUX2_X1 U615 ( .A(n11), .B(n10), .S(n244), .Z(n12) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n249), .Z(n13) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n249), .Z(n14) );
  MUX2_X1 U618 ( .A(n14), .B(n13), .S(n244), .Z(n15) );
  MUX2_X1 U619 ( .A(n15), .B(n12), .S(n243), .Z(n16) );
  MUX2_X1 U620 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n247), .Z(n18) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n247), .Z(n19) );
  MUX2_X1 U623 ( .A(n19), .B(n18), .S(n245), .Z(n20) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n247), .Z(n21) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n247), .Z(n22) );
  MUX2_X1 U626 ( .A(n22), .B(n21), .S(n245), .Z(n23) );
  MUX2_X1 U627 ( .A(n23), .B(n20), .S(n243), .Z(n24) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n247), .Z(n25) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n247), .Z(n26) );
  MUX2_X1 U630 ( .A(n26), .B(n25), .S(n245), .Z(n27) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n247), .Z(n28) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n247), .Z(n29) );
  MUX2_X1 U633 ( .A(n29), .B(n28), .S(n245), .Z(n30) );
  MUX2_X1 U634 ( .A(n30), .B(n27), .S(n243), .Z(n31) );
  MUX2_X1 U635 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U636 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n247), .Z(n33) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n247), .Z(n34) );
  MUX2_X1 U639 ( .A(n34), .B(n33), .S(n245), .Z(n35) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n247), .Z(n36) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n247), .Z(n37) );
  MUX2_X1 U642 ( .A(n37), .B(n36), .S(n245), .Z(n38) );
  MUX2_X1 U643 ( .A(n38), .B(n35), .S(n243), .Z(n39) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n248), .Z(n40) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n248), .Z(n41) );
  MUX2_X1 U646 ( .A(n41), .B(n40), .S(n245), .Z(n42) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n248), .Z(n43) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n248), .Z(n44) );
  MUX2_X1 U649 ( .A(n44), .B(n43), .S(n245), .Z(n45) );
  MUX2_X1 U650 ( .A(n45), .B(n42), .S(N12), .Z(n46) );
  MUX2_X1 U651 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n248), .Z(n48) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n248), .Z(n49) );
  MUX2_X1 U654 ( .A(n49), .B(n48), .S(n245), .Z(n50) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n248), .Z(n51) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n248), .Z(n52) );
  MUX2_X1 U657 ( .A(n52), .B(n51), .S(n245), .Z(n53) );
  MUX2_X1 U658 ( .A(n53), .B(n50), .S(N12), .Z(n54) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n248), .Z(n55) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n248), .Z(n56) );
  MUX2_X1 U661 ( .A(n56), .B(n55), .S(n245), .Z(n57) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n248), .Z(n58) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n248), .Z(n59) );
  MUX2_X1 U664 ( .A(n59), .B(n58), .S(n245), .Z(n60) );
  MUX2_X1 U665 ( .A(n60), .B(n57), .S(N12), .Z(n61) );
  MUX2_X1 U666 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U667 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n249), .Z(n63) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n249), .Z(n64) );
  MUX2_X1 U670 ( .A(n64), .B(n63), .S(n246), .Z(n65) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n249), .Z(n66) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n249), .Z(n67) );
  MUX2_X1 U673 ( .A(n67), .B(n66), .S(n246), .Z(n68) );
  MUX2_X1 U674 ( .A(n68), .B(n65), .S(n243), .Z(n69) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n249), .Z(n70) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n249), .Z(n71) );
  MUX2_X1 U677 ( .A(n71), .B(n70), .S(n246), .Z(n72) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n249), .Z(n73) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n249), .Z(n74) );
  MUX2_X1 U680 ( .A(n74), .B(n73), .S(n246), .Z(n75) );
  MUX2_X1 U681 ( .A(n75), .B(n72), .S(n243), .Z(n76) );
  MUX2_X1 U682 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n249), .Z(n78) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n249), .Z(n79) );
  MUX2_X1 U685 ( .A(n79), .B(n78), .S(n246), .Z(n80) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n249), .Z(n81) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n249), .Z(n82) );
  MUX2_X1 U688 ( .A(n82), .B(n81), .S(n246), .Z(n83) );
  MUX2_X1 U689 ( .A(n83), .B(n80), .S(n243), .Z(n84) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n250), .Z(n85) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n250), .Z(n86) );
  MUX2_X1 U692 ( .A(n86), .B(n85), .S(n246), .Z(n87) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n250), .Z(n88) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n250), .Z(n89) );
  MUX2_X1 U695 ( .A(n89), .B(n88), .S(n246), .Z(n90) );
  MUX2_X1 U696 ( .A(n90), .B(n87), .S(n243), .Z(n91) );
  MUX2_X1 U697 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U698 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n250), .Z(n93) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U701 ( .A(n94), .B(n93), .S(n246), .Z(n95) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n250), .Z(n96) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n250), .Z(n97) );
  MUX2_X1 U704 ( .A(n97), .B(n96), .S(n246), .Z(n98) );
  MUX2_X1 U705 ( .A(n98), .B(n95), .S(n243), .Z(n99) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n100) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n250), .Z(n101) );
  MUX2_X1 U708 ( .A(n101), .B(n100), .S(n246), .Z(n102) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n250), .Z(n103) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n250), .Z(n104) );
  MUX2_X1 U711 ( .A(n104), .B(n103), .S(n246), .Z(n105) );
  MUX2_X1 U712 ( .A(n105), .B(n102), .S(n243), .Z(n106) );
  MUX2_X1 U713 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n252), .Z(n108) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(N10), .Z(n109) );
  MUX2_X1 U716 ( .A(n109), .B(n108), .S(n246), .Z(n110) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(N10), .Z(n111) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n247), .Z(n112) );
  MUX2_X1 U719 ( .A(n112), .B(n111), .S(N11), .Z(n113) );
  MUX2_X1 U720 ( .A(n113), .B(n110), .S(n243), .Z(n114) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(N10), .Z(n115) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n252), .Z(n116) );
  MUX2_X1 U723 ( .A(n116), .B(n115), .S(N11), .Z(n117) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n118) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n248), .Z(n119) );
  MUX2_X1 U726 ( .A(n119), .B(n118), .S(n245), .Z(n120) );
  MUX2_X1 U727 ( .A(n120), .B(n117), .S(n243), .Z(n121) );
  MUX2_X1 U728 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U729 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n248), .Z(n123) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(N10), .Z(n124) );
  MUX2_X1 U732 ( .A(n124), .B(n123), .S(n245), .Z(n125) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(N10), .Z(n126) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n127) );
  MUX2_X1 U735 ( .A(n127), .B(n126), .S(N11), .Z(n128) );
  MUX2_X1 U736 ( .A(n128), .B(n125), .S(n243), .Z(n129) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n251), .Z(n130) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(N10), .Z(n131) );
  MUX2_X1 U739 ( .A(n131), .B(n130), .S(N11), .Z(n132) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n252), .Z(n133) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(N10), .Z(n134) );
  MUX2_X1 U742 ( .A(n134), .B(n133), .S(n246), .Z(n135) );
  MUX2_X1 U743 ( .A(n135), .B(n132), .S(n243), .Z(n136) );
  MUX2_X1 U744 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n251), .Z(n138) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n252), .Z(n139) );
  MUX2_X1 U747 ( .A(n139), .B(n138), .S(N11), .Z(n140) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n247), .Z(n141) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(N10), .Z(n142) );
  MUX2_X1 U750 ( .A(n142), .B(n141), .S(n245), .Z(n143) );
  MUX2_X1 U751 ( .A(n143), .B(n140), .S(n243), .Z(n144) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(N10), .Z(n145) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(N10), .Z(n146) );
  MUX2_X1 U754 ( .A(n146), .B(n145), .S(N11), .Z(n147) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(N10), .Z(n148) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n149) );
  MUX2_X1 U757 ( .A(n149), .B(n148), .S(n246), .Z(n150) );
  MUX2_X1 U758 ( .A(n150), .B(n147), .S(n243), .Z(n151) );
  MUX2_X1 U759 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U760 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n251), .Z(n153) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n251), .Z(n154) );
  MUX2_X1 U763 ( .A(n154), .B(n153), .S(n245), .Z(n155) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n251), .Z(n156) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n251), .Z(n157) );
  MUX2_X1 U766 ( .A(n157), .B(n156), .S(n246), .Z(n158) );
  MUX2_X1 U767 ( .A(n158), .B(n155), .S(n243), .Z(n159) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n251), .Z(n160) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n251), .Z(n161) );
  MUX2_X1 U770 ( .A(n161), .B(n160), .S(n244), .Z(n162) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n251), .Z(n163) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n251), .Z(n164) );
  MUX2_X1 U773 ( .A(n164), .B(n163), .S(N11), .Z(n165) );
  MUX2_X1 U774 ( .A(n165), .B(n162), .S(N12), .Z(n166) );
  MUX2_X1 U775 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n251), .Z(n168) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n251), .Z(n169) );
  MUX2_X1 U778 ( .A(n169), .B(n168), .S(N11), .Z(n170) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n251), .Z(n171) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n251), .Z(n172) );
  MUX2_X1 U781 ( .A(n172), .B(n171), .S(N11), .Z(n173) );
  MUX2_X1 U782 ( .A(n173), .B(n170), .S(n243), .Z(n174) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n252), .Z(n175) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n247), .Z(n176) );
  MUX2_X1 U785 ( .A(n176), .B(n175), .S(n244), .Z(n177) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n252), .Z(n178) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n247), .Z(n179) );
  MUX2_X1 U788 ( .A(n179), .B(n178), .S(N11), .Z(n180) );
  MUX2_X1 U789 ( .A(n180), .B(n177), .S(N12), .Z(n181) );
  MUX2_X1 U790 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U791 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n247), .Z(n183) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n250), .Z(n184) );
  MUX2_X1 U794 ( .A(n184), .B(n183), .S(n246), .Z(n185) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n251), .Z(n186) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n252), .Z(n187) );
  MUX2_X1 U797 ( .A(n187), .B(n186), .S(N11), .Z(n188) );
  MUX2_X1 U798 ( .A(n188), .B(n185), .S(n243), .Z(n189) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n252), .Z(n190) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n252), .Z(n191) );
  MUX2_X1 U801 ( .A(n191), .B(n190), .S(n245), .Z(n192) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n249), .Z(n193) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n252), .Z(n194) );
  MUX2_X1 U804 ( .A(n194), .B(n193), .S(N11), .Z(n195) );
  MUX2_X1 U805 ( .A(n195), .B(n192), .S(N12), .Z(n196) );
  MUX2_X1 U806 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n250), .Z(n198) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n252), .Z(n199) );
  MUX2_X1 U809 ( .A(n199), .B(n198), .S(n244), .Z(n200) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n248), .Z(n201) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n249), .Z(n202) );
  MUX2_X1 U812 ( .A(n202), .B(n201), .S(n245), .Z(n203) );
  MUX2_X1 U813 ( .A(n203), .B(n200), .S(n243), .Z(n204) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n250), .Z(n205) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n252), .Z(n206) );
  MUX2_X1 U816 ( .A(n206), .B(n205), .S(n244), .Z(n207) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n252), .Z(n208) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n249), .Z(n209) );
  MUX2_X1 U819 ( .A(n209), .B(n208), .S(N11), .Z(n210) );
  MUX2_X1 U820 ( .A(n210), .B(n207), .S(N12), .Z(n211) );
  MUX2_X1 U821 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U822 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n249), .Z(n213) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n249), .Z(n214) );
  MUX2_X1 U825 ( .A(n214), .B(n213), .S(n244), .Z(n215) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n247), .Z(n216) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n250), .Z(n217) );
  MUX2_X1 U828 ( .A(n217), .B(n216), .S(n244), .Z(n218) );
  MUX2_X1 U829 ( .A(n218), .B(n215), .S(n243), .Z(n219) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n252), .Z(n220) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n250), .Z(n221) );
  MUX2_X1 U832 ( .A(n221), .B(n220), .S(n244), .Z(n222) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n252), .Z(n223) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n250), .Z(n224) );
  MUX2_X1 U835 ( .A(n224), .B(n223), .S(n244), .Z(n225) );
  MUX2_X1 U836 ( .A(n225), .B(n222), .S(N12), .Z(n226) );
  MUX2_X1 U837 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(N10), .Z(n228) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n248), .Z(n229) );
  MUX2_X1 U840 ( .A(n229), .B(n228), .S(n244), .Z(n230) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n252), .Z(n231) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n248), .Z(n232) );
  MUX2_X1 U843 ( .A(n232), .B(n231), .S(n246), .Z(n233) );
  MUX2_X1 U844 ( .A(n233), .B(n230), .S(n243), .Z(n234) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n247), .Z(n235) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n252), .Z(n236) );
  MUX2_X1 U847 ( .A(n236), .B(n235), .S(n244), .Z(n237) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n252), .Z(n238) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n252), .Z(n239) );
  MUX2_X1 U850 ( .A(n239), .B(n238), .S(n244), .Z(n240) );
  MUX2_X1 U851 ( .A(n240), .B(n237), .S(N12), .Z(n241) );
  MUX2_X1 U852 ( .A(n241), .B(n234), .S(N13), .Z(n242) );
  MUX2_X1 U853 ( .A(n242), .B(n227), .S(N14), .Z(N15) );
  CLKBUF_X1 U854 ( .A(N11), .Z(n244) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_10 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X2 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  BUF_X1 U3 ( .A(N10), .Z(n247) );
  BUF_X1 U4 ( .A(n250), .Z(n248) );
  BUF_X1 U5 ( .A(n250), .Z(n249) );
  BUF_X1 U6 ( .A(n250), .Z(n246) );
  BUF_X1 U7 ( .A(n250), .Z(n245) );
  BUF_X1 U8 ( .A(N10), .Z(n250) );
  INV_X1 U9 ( .A(n1111), .ZN(n841) );
  INV_X1 U10 ( .A(n1100), .ZN(n840) );
  INV_X1 U11 ( .A(n1090), .ZN(n839) );
  INV_X1 U12 ( .A(n1080), .ZN(n838) );
  INV_X1 U13 ( .A(n1070), .ZN(n837) );
  INV_X1 U14 ( .A(n1060), .ZN(n836) );
  INV_X1 U15 ( .A(n1051), .ZN(n835) );
  INV_X1 U16 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U19 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U20 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U21 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U22 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U23 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U24 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U26 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U27 ( .A(n1131), .ZN(n816) );
  INV_X1 U28 ( .A(n1121), .ZN(n815) );
  INV_X1 U29 ( .A(n887), .ZN(n814) );
  INV_X1 U30 ( .A(n878), .ZN(n813) );
  INV_X1 U31 ( .A(n869), .ZN(n812) );
  INV_X1 U32 ( .A(n860), .ZN(n811) );
  INV_X1 U33 ( .A(n851), .ZN(n810) );
  INV_X1 U34 ( .A(n987), .ZN(n828) );
  INV_X1 U35 ( .A(n978), .ZN(n827) );
  INV_X1 U36 ( .A(n969), .ZN(n826) );
  INV_X1 U37 ( .A(n914), .ZN(n820) );
  INV_X1 U38 ( .A(n905), .ZN(n819) );
  INV_X1 U39 ( .A(n896), .ZN(n818) );
  INV_X1 U40 ( .A(n1033), .ZN(n833) );
  INV_X1 U41 ( .A(n1023), .ZN(n832) );
  INV_X1 U42 ( .A(n1014), .ZN(n831) );
  INV_X1 U43 ( .A(n1005), .ZN(n830) );
  INV_X1 U44 ( .A(n996), .ZN(n829) );
  INV_X1 U45 ( .A(n960), .ZN(n825) );
  INV_X1 U46 ( .A(n950), .ZN(n824) );
  INV_X1 U47 ( .A(n941), .ZN(n823) );
  INV_X1 U48 ( .A(n932), .ZN(n822) );
  INV_X1 U49 ( .A(n923), .ZN(n821) );
  INV_X1 U50 ( .A(n1142), .ZN(n817) );
  BUF_X1 U51 ( .A(N11), .Z(n242) );
  BUF_X1 U52 ( .A(N11), .Z(n243) );
  BUF_X1 U53 ( .A(N11), .Z(n244) );
  INV_X1 U54 ( .A(N10), .ZN(n251) );
  BUF_X1 U55 ( .A(N12), .Z(n241) );
  NOR3_X1 U56 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U57 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U58 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U60 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U62 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U63 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U64 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U65 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U67 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U69 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U70 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U71 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U72 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U73 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U74 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U75 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U76 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U77 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U79 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U81 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U82 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U83 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U84 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U85 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U86 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U88 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U89 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U90 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U91 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U92 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U93 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U94 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U95 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U96 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U97 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U98 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U99 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U100 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U101 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U102 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U103 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U104 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U105 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U106 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U107 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U108 ( .A(n988), .ZN(n705) );
  AOI22_X1 U109 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U110 ( .A(n986), .ZN(n704) );
  AOI22_X1 U111 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U112 ( .A(n985), .ZN(n703) );
  AOI22_X1 U113 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U114 ( .A(n984), .ZN(n702) );
  AOI22_X1 U115 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U116 ( .A(n983), .ZN(n701) );
  AOI22_X1 U117 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U118 ( .A(n982), .ZN(n700) );
  AOI22_X1 U119 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U120 ( .A(n981), .ZN(n699) );
  AOI22_X1 U121 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U122 ( .A(n980), .ZN(n698) );
  AOI22_X1 U123 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U124 ( .A(n949), .ZN(n672) );
  AOI22_X1 U125 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U126 ( .A(n948), .ZN(n671) );
  AOI22_X1 U127 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U128 ( .A(n947), .ZN(n670) );
  AOI22_X1 U129 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U130 ( .A(n946), .ZN(n669) );
  AOI22_X1 U131 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U132 ( .A(n945), .ZN(n668) );
  AOI22_X1 U133 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U134 ( .A(n944), .ZN(n667) );
  AOI22_X1 U135 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U136 ( .A(n943), .ZN(n666) );
  AOI22_X1 U137 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U138 ( .A(n915), .ZN(n641) );
  AOI22_X1 U139 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U140 ( .A(n913), .ZN(n640) );
  AOI22_X1 U141 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U142 ( .A(n912), .ZN(n639) );
  AOI22_X1 U143 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U144 ( .A(n911), .ZN(n638) );
  AOI22_X1 U145 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U146 ( .A(n910), .ZN(n637) );
  AOI22_X1 U147 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U148 ( .A(n909), .ZN(n636) );
  AOI22_X1 U149 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U150 ( .A(n908), .ZN(n635) );
  AOI22_X1 U151 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U152 ( .A(n907), .ZN(n634) );
  AOI22_X1 U153 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U154 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U155 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U156 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U157 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U158 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U159 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U160 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U161 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U162 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U163 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U164 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U165 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U166 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U167 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U168 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U169 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U170 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U171 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U172 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U173 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U174 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U175 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U176 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U177 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U178 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U179 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U180 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U181 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U182 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U183 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U184 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U185 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U186 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U187 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U188 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U189 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U190 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U191 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U192 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U193 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U194 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U195 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U196 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U197 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U198 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U199 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U200 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U201 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U202 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U203 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U204 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U205 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U206 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U207 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U208 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U209 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U210 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U211 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U212 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U213 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U214 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U215 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U216 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U217 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U218 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U219 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U220 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U221 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U222 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U223 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U224 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U225 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U226 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U227 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U228 ( .A(n999), .ZN(n715) );
  AOI22_X1 U229 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U230 ( .A(n998), .ZN(n714) );
  AOI22_X1 U231 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U232 ( .A(n951), .ZN(n673) );
  AOI22_X1 U233 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U234 ( .A(n979), .ZN(n697) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U236 ( .A(n977), .ZN(n696) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U238 ( .A(n976), .ZN(n695) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U240 ( .A(n975), .ZN(n694) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U242 ( .A(n974), .ZN(n693) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U244 ( .A(n973), .ZN(n692) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U246 ( .A(n972), .ZN(n691) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U248 ( .A(n971), .ZN(n690) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U250 ( .A(n970), .ZN(n689) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U252 ( .A(n968), .ZN(n688) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U254 ( .A(n967), .ZN(n687) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U256 ( .A(n966), .ZN(n686) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U258 ( .A(n965), .ZN(n685) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U260 ( .A(n964), .ZN(n684) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U262 ( .A(n963), .ZN(n683) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U264 ( .A(n962), .ZN(n682) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U266 ( .A(n942), .ZN(n665) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U268 ( .A(n940), .ZN(n664) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U270 ( .A(n939), .ZN(n663) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U272 ( .A(n938), .ZN(n662) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U274 ( .A(n937), .ZN(n661) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U276 ( .A(n936), .ZN(n660) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U278 ( .A(n935), .ZN(n659) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U280 ( .A(n934), .ZN(n658) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U282 ( .A(n933), .ZN(n657) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U284 ( .A(n931), .ZN(n656) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U286 ( .A(n930), .ZN(n655) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U288 ( .A(n929), .ZN(n654) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U290 ( .A(n928), .ZN(n653) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U292 ( .A(n927), .ZN(n652) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U294 ( .A(n926), .ZN(n651) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U296 ( .A(n925), .ZN(n650) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U298 ( .A(n906), .ZN(n633) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U300 ( .A(n904), .ZN(n632) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U302 ( .A(n903), .ZN(n631) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U304 ( .A(n902), .ZN(n630) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U306 ( .A(n901), .ZN(n629) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U308 ( .A(n900), .ZN(n628) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U310 ( .A(n899), .ZN(n627) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U312 ( .A(n898), .ZN(n626) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U314 ( .A(n897), .ZN(n625) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U316 ( .A(n895), .ZN(n624) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U318 ( .A(n894), .ZN(n623) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U320 ( .A(n893), .ZN(n622) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U322 ( .A(n892), .ZN(n621) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U324 ( .A(n891), .ZN(n620) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U326 ( .A(n890), .ZN(n619) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U328 ( .A(n889), .ZN(n618) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U330 ( .A(N12), .ZN(n253) );
  INV_X1 U331 ( .A(N11), .ZN(n252) );
  INV_X1 U332 ( .A(n997), .ZN(n713) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U334 ( .A(n995), .ZN(n712) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U336 ( .A(n994), .ZN(n711) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U338 ( .A(n993), .ZN(n710) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U340 ( .A(n992), .ZN(n709) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U342 ( .A(n991), .ZN(n708) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U344 ( .A(n990), .ZN(n707) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U346 ( .A(n989), .ZN(n706) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U348 ( .A(n924), .ZN(n649) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U350 ( .A(n922), .ZN(n648) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U352 ( .A(n921), .ZN(n647) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U354 ( .A(n920), .ZN(n646) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U356 ( .A(n919), .ZN(n645) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U358 ( .A(n918), .ZN(n644) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U360 ( .A(n917), .ZN(n643) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U362 ( .A(n916), .ZN(n642) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U364 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U366 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U368 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U370 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U372 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U374 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U376 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U378 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U380 ( .A(n961), .ZN(n681) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U382 ( .A(n959), .ZN(n680) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U384 ( .A(n958), .ZN(n679) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U386 ( .A(n957), .ZN(n678) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U388 ( .A(n956), .ZN(n677) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U390 ( .A(n955), .ZN(n676) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U392 ( .A(n954), .ZN(n675) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U394 ( .A(n953), .ZN(n674) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U396 ( .A(n888), .ZN(n617) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U398 ( .A(n886), .ZN(n616) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U400 ( .A(n885), .ZN(n615) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U402 ( .A(n884), .ZN(n614) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U404 ( .A(n883), .ZN(n613) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U406 ( .A(n882), .ZN(n612) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U408 ( .A(n881), .ZN(n611) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U410 ( .A(n880), .ZN(n610) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U412 ( .A(n879), .ZN(n609) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U414 ( .A(n877), .ZN(n608) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U416 ( .A(n876), .ZN(n607) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U418 ( .A(n875), .ZN(n606) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U420 ( .A(n874), .ZN(n605) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U422 ( .A(n873), .ZN(n604) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U424 ( .A(n872), .ZN(n603) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U426 ( .A(n871), .ZN(n602) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U428 ( .A(n870), .ZN(n601) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U430 ( .A(n868), .ZN(n600) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U432 ( .A(n867), .ZN(n599) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U434 ( .A(n866), .ZN(n598) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U436 ( .A(n865), .ZN(n597) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U438 ( .A(n864), .ZN(n596) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U440 ( .A(n863), .ZN(n595) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U442 ( .A(n862), .ZN(n594) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U444 ( .A(n861), .ZN(n293) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U446 ( .A(n859), .ZN(n292) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U448 ( .A(n858), .ZN(n291) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U450 ( .A(n857), .ZN(n290) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U452 ( .A(n856), .ZN(n289) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U454 ( .A(n855), .ZN(n288) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U456 ( .A(n854), .ZN(n287) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U458 ( .A(n853), .ZN(n286) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U460 ( .A(n852), .ZN(n285) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U462 ( .A(n850), .ZN(n284) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U464 ( .A(n849), .ZN(n283) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U466 ( .A(n848), .ZN(n282) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U468 ( .A(n847), .ZN(n281) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U470 ( .A(n846), .ZN(n280) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U472 ( .A(n845), .ZN(n279) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U474 ( .A(n844), .ZN(n278) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U476 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U477 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U478 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U479 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U480 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U481 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U482 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U483 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U484 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U485 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U486 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U487 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U488 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U489 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U490 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U491 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U492 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U494 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U496 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U498 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U500 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U502 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U504 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U506 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U508 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U510 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U512 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U514 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U516 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U518 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U520 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U522 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U524 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U526 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U528 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U530 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U532 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U534 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U536 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U538 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U540 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U542 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U544 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U546 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U548 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U550 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U552 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U554 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U556 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U558 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U560 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U562 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U564 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U566 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U568 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U570 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U572 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U574 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U576 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U578 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U580 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U582 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U584 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U586 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U588 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U590 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U592 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U594 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U596 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U598 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U600 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U602 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U604 ( .A(N13), .ZN(n842) );
  INV_X1 U605 ( .A(N14), .ZN(n843) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n247), .Z(n1) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n247), .Z(n2) );
  MUX2_X1 U608 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n247), .Z(n4) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n247), .Z(n5) );
  MUX2_X1 U611 ( .A(n5), .B(n4), .S(n242), .Z(n6) );
  MUX2_X1 U612 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n247), .Z(n8) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n249), .Z(n9) );
  MUX2_X1 U615 ( .A(n9), .B(n8), .S(n243), .Z(n10) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n247), .Z(n11) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n248), .Z(n12) );
  MUX2_X1 U618 ( .A(n12), .B(n11), .S(n244), .Z(n13) );
  MUX2_X1 U619 ( .A(n13), .B(n10), .S(N12), .Z(n14) );
  MUX2_X1 U620 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n245), .Z(n16) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n245), .Z(n17) );
  MUX2_X1 U623 ( .A(n17), .B(n16), .S(N11), .Z(n18) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n245), .Z(n20) );
  MUX2_X1 U626 ( .A(n20), .B(n19), .S(N11), .Z(n21) );
  MUX2_X1 U627 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n245), .Z(n23) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n245), .Z(n24) );
  MUX2_X1 U630 ( .A(n24), .B(n23), .S(N11), .Z(n25) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n245), .Z(n26) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n245), .Z(n27) );
  MUX2_X1 U633 ( .A(n27), .B(n26), .S(N11), .Z(n28) );
  MUX2_X1 U634 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U635 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U636 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n245), .Z(n31) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n245), .Z(n32) );
  MUX2_X1 U639 ( .A(n32), .B(n31), .S(n243), .Z(n33) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U642 ( .A(n35), .B(n34), .S(N11), .Z(n36) );
  MUX2_X1 U643 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n246), .Z(n38) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n246), .Z(n39) );
  MUX2_X1 U646 ( .A(n39), .B(n38), .S(n242), .Z(n40) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n246), .Z(n41) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n246), .Z(n42) );
  MUX2_X1 U649 ( .A(n42), .B(n41), .S(n243), .Z(n43) );
  MUX2_X1 U650 ( .A(n43), .B(n40), .S(n241), .Z(n44) );
  MUX2_X1 U651 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n246), .Z(n46) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n246), .Z(n47) );
  MUX2_X1 U654 ( .A(n47), .B(n46), .S(n244), .Z(n48) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n246), .Z(n49) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n246), .Z(n50) );
  MUX2_X1 U657 ( .A(n50), .B(n49), .S(n242), .Z(n51) );
  MUX2_X1 U658 ( .A(n51), .B(n48), .S(n241), .Z(n52) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n246), .Z(n53) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n246), .Z(n54) );
  MUX2_X1 U661 ( .A(n54), .B(n53), .S(n244), .Z(n55) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n246), .Z(n56) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n246), .Z(n57) );
  MUX2_X1 U664 ( .A(n57), .B(n56), .S(N11), .Z(n58) );
  MUX2_X1 U665 ( .A(n58), .B(n55), .S(n241), .Z(n59) );
  MUX2_X1 U666 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U667 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n249), .Z(n61) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n246), .Z(n62) );
  MUX2_X1 U670 ( .A(n62), .B(n61), .S(N11), .Z(n63) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n248), .Z(n64) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n245), .Z(n65) );
  MUX2_X1 U673 ( .A(n65), .B(n64), .S(n243), .Z(n66) );
  MUX2_X1 U674 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n249), .Z(n68) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n248), .Z(n69) );
  MUX2_X1 U677 ( .A(n69), .B(n68), .S(n244), .Z(n70) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n249), .Z(n71) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n246), .Z(n72) );
  MUX2_X1 U680 ( .A(n72), .B(n71), .S(N11), .Z(n73) );
  MUX2_X1 U681 ( .A(n73), .B(n70), .S(n241), .Z(n74) );
  MUX2_X1 U682 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n245), .Z(n76) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n246), .Z(n77) );
  MUX2_X1 U685 ( .A(n77), .B(n76), .S(n242), .Z(n78) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n245), .Z(n79) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n249), .Z(n80) );
  MUX2_X1 U688 ( .A(n80), .B(n79), .S(n242), .Z(n81) );
  MUX2_X1 U689 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n250), .Z(n83) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n250), .Z(n84) );
  MUX2_X1 U692 ( .A(n84), .B(n83), .S(n244), .Z(n85) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n250), .Z(n86) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n248), .Z(n87) );
  MUX2_X1 U695 ( .A(n87), .B(n86), .S(n243), .Z(n88) );
  MUX2_X1 U696 ( .A(n88), .B(n85), .S(n241), .Z(n89) );
  MUX2_X1 U697 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U698 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n250), .Z(n91) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n92) );
  MUX2_X1 U701 ( .A(n92), .B(n91), .S(N11), .Z(n93) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n250), .Z(n95) );
  MUX2_X1 U704 ( .A(n95), .B(n94), .S(N11), .Z(n96) );
  MUX2_X1 U705 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n98) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n250), .Z(n99) );
  MUX2_X1 U708 ( .A(n99), .B(n98), .S(N11), .Z(n100) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n250), .Z(n101) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n250), .Z(n102) );
  MUX2_X1 U711 ( .A(n102), .B(n101), .S(N11), .Z(n103) );
  MUX2_X1 U712 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U713 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n247), .Z(n106) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n247), .Z(n107) );
  MUX2_X1 U716 ( .A(n107), .B(n106), .S(n242), .Z(n108) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n247), .Z(n109) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n247), .Z(n110) );
  MUX2_X1 U719 ( .A(n110), .B(n109), .S(n242), .Z(n111) );
  MUX2_X1 U720 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n247), .Z(n113) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n247), .Z(n114) );
  MUX2_X1 U723 ( .A(n114), .B(n113), .S(n242), .Z(n115) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n247), .Z(n116) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n247), .Z(n117) );
  MUX2_X1 U726 ( .A(n117), .B(n116), .S(n242), .Z(n118) );
  MUX2_X1 U727 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U728 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U729 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n247), .Z(n121) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n247), .Z(n122) );
  MUX2_X1 U732 ( .A(n122), .B(n121), .S(n242), .Z(n123) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n247), .Z(n124) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n247), .Z(n125) );
  MUX2_X1 U735 ( .A(n125), .B(n124), .S(n242), .Z(n126) );
  MUX2_X1 U736 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n248), .Z(n128) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n248), .Z(n129) );
  MUX2_X1 U739 ( .A(n129), .B(n128), .S(n242), .Z(n130) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n248), .Z(n131) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n248), .Z(n132) );
  MUX2_X1 U742 ( .A(n132), .B(n131), .S(n242), .Z(n133) );
  MUX2_X1 U743 ( .A(n133), .B(n130), .S(n241), .Z(n134) );
  MUX2_X1 U744 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n248), .Z(n136) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n248), .Z(n137) );
  MUX2_X1 U747 ( .A(n137), .B(n136), .S(n242), .Z(n138) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n248), .Z(n139) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n248), .Z(n140) );
  MUX2_X1 U750 ( .A(n140), .B(n139), .S(n242), .Z(n141) );
  MUX2_X1 U751 ( .A(n141), .B(n138), .S(n241), .Z(n142) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n248), .Z(n143) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n248), .Z(n144) );
  MUX2_X1 U754 ( .A(n144), .B(n143), .S(n242), .Z(n145) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n248), .Z(n146) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n248), .Z(n147) );
  MUX2_X1 U757 ( .A(n147), .B(n146), .S(n242), .Z(n148) );
  MUX2_X1 U758 ( .A(n148), .B(n145), .S(n241), .Z(n149) );
  MUX2_X1 U759 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U760 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n249), .Z(n151) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n249), .Z(n152) );
  MUX2_X1 U763 ( .A(n152), .B(n151), .S(n243), .Z(n153) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n249), .Z(n154) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n249), .Z(n155) );
  MUX2_X1 U766 ( .A(n155), .B(n154), .S(n243), .Z(n156) );
  MUX2_X1 U767 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n249), .Z(n158) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n249), .Z(n159) );
  MUX2_X1 U770 ( .A(n159), .B(n158), .S(n243), .Z(n160) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n249), .Z(n161) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n249), .Z(n162) );
  MUX2_X1 U773 ( .A(n162), .B(n161), .S(n243), .Z(n163) );
  MUX2_X1 U774 ( .A(n163), .B(n160), .S(N12), .Z(n164) );
  MUX2_X1 U775 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n249), .Z(n166) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n249), .Z(n167) );
  MUX2_X1 U778 ( .A(n167), .B(n166), .S(n243), .Z(n168) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n249), .Z(n169) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n249), .Z(n170) );
  MUX2_X1 U781 ( .A(n170), .B(n169), .S(n243), .Z(n171) );
  MUX2_X1 U782 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n247), .Z(n173) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n250), .Z(n174) );
  MUX2_X1 U785 ( .A(n174), .B(n173), .S(n243), .Z(n175) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n176) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n250), .Z(n177) );
  MUX2_X1 U788 ( .A(n177), .B(n176), .S(n243), .Z(n178) );
  MUX2_X1 U789 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U790 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U791 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n249), .Z(n181) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n250), .Z(n182) );
  MUX2_X1 U794 ( .A(n182), .B(n181), .S(n243), .Z(n183) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n248), .Z(n184) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(N10), .Z(n185) );
  MUX2_X1 U797 ( .A(n185), .B(n184), .S(n243), .Z(n186) );
  MUX2_X1 U798 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n245), .Z(n188) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(N10), .Z(n189) );
  MUX2_X1 U801 ( .A(n189), .B(n188), .S(n243), .Z(n190) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n248), .Z(n191) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n250), .Z(n192) );
  MUX2_X1 U804 ( .A(n192), .B(n191), .S(n243), .Z(n193) );
  MUX2_X1 U805 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U806 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n246), .Z(n196) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n250), .Z(n197) );
  MUX2_X1 U809 ( .A(n197), .B(n196), .S(n244), .Z(n198) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n250), .Z(n199) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n200) );
  MUX2_X1 U812 ( .A(n200), .B(n199), .S(n244), .Z(n201) );
  MUX2_X1 U813 ( .A(n201), .B(n198), .S(N12), .Z(n202) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n250), .Z(n203) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n204) );
  MUX2_X1 U816 ( .A(n204), .B(n203), .S(n244), .Z(n205) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n206) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n207) );
  MUX2_X1 U819 ( .A(n207), .B(n206), .S(n244), .Z(n208) );
  MUX2_X1 U820 ( .A(n208), .B(n205), .S(N12), .Z(n209) );
  MUX2_X1 U821 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U822 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n246), .Z(n211) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n245), .Z(n212) );
  MUX2_X1 U825 ( .A(n212), .B(n211), .S(n244), .Z(n213) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n246), .Z(n214) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(N10), .Z(n215) );
  MUX2_X1 U828 ( .A(n215), .B(n214), .S(n244), .Z(n216) );
  MUX2_X1 U829 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n247), .Z(n218) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n250), .Z(n219) );
  MUX2_X1 U832 ( .A(n219), .B(n218), .S(n244), .Z(n220) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n247), .Z(n221) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n222) );
  MUX2_X1 U835 ( .A(n222), .B(n221), .S(n244), .Z(n223) );
  MUX2_X1 U836 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U837 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n247), .Z(n226) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n250), .Z(n227) );
  MUX2_X1 U840 ( .A(n227), .B(n226), .S(n244), .Z(n228) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n247), .Z(n229) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n230) );
  MUX2_X1 U843 ( .A(n230), .B(n229), .S(n244), .Z(n231) );
  MUX2_X1 U844 ( .A(n231), .B(n228), .S(N12), .Z(n232) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n233) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n234) );
  MUX2_X1 U847 ( .A(n234), .B(n233), .S(n244), .Z(n235) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n236) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n237) );
  MUX2_X1 U850 ( .A(n237), .B(n236), .S(n244), .Z(n238) );
  MUX2_X1 U851 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U852 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U853 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_9 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(n250), .Z(n248) );
  BUF_X1 U4 ( .A(n250), .Z(n249) );
  BUF_X1 U5 ( .A(N10), .Z(n246) );
  BUF_X1 U6 ( .A(n250), .Z(n247) );
  BUF_X1 U7 ( .A(N10), .Z(n250) );
  INV_X1 U8 ( .A(n1111), .ZN(n841) );
  INV_X1 U9 ( .A(n1100), .ZN(n840) );
  INV_X1 U10 ( .A(n1090), .ZN(n839) );
  INV_X1 U11 ( .A(n1080), .ZN(n838) );
  INV_X1 U12 ( .A(n1070), .ZN(n837) );
  INV_X1 U13 ( .A(n1060), .ZN(n836) );
  INV_X1 U14 ( .A(n1051), .ZN(n835) );
  INV_X1 U15 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U16 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U18 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U19 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U20 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U21 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U22 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U23 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U24 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U26 ( .A(n1131), .ZN(n816) );
  INV_X1 U27 ( .A(n1121), .ZN(n815) );
  INV_X1 U28 ( .A(n887), .ZN(n814) );
  INV_X1 U29 ( .A(n878), .ZN(n813) );
  INV_X1 U30 ( .A(n869), .ZN(n812) );
  INV_X1 U31 ( .A(n860), .ZN(n811) );
  INV_X1 U32 ( .A(n851), .ZN(n810) );
  INV_X1 U33 ( .A(n987), .ZN(n828) );
  INV_X1 U34 ( .A(n978), .ZN(n827) );
  INV_X1 U35 ( .A(n969), .ZN(n826) );
  INV_X1 U36 ( .A(n914), .ZN(n820) );
  INV_X1 U37 ( .A(n905), .ZN(n819) );
  INV_X1 U38 ( .A(n896), .ZN(n818) );
  INV_X1 U39 ( .A(n1033), .ZN(n833) );
  INV_X1 U40 ( .A(n1023), .ZN(n832) );
  INV_X1 U41 ( .A(n1014), .ZN(n831) );
  INV_X1 U42 ( .A(n1005), .ZN(n830) );
  INV_X1 U43 ( .A(n996), .ZN(n829) );
  INV_X1 U44 ( .A(n960), .ZN(n825) );
  INV_X1 U45 ( .A(n950), .ZN(n824) );
  INV_X1 U46 ( .A(n941), .ZN(n823) );
  INV_X1 U47 ( .A(n932), .ZN(n822) );
  INV_X1 U48 ( .A(n923), .ZN(n821) );
  INV_X1 U49 ( .A(n1142), .ZN(n817) );
  BUF_X1 U50 ( .A(N11), .Z(n242) );
  BUF_X1 U51 ( .A(N11), .Z(n243) );
  BUF_X1 U52 ( .A(N11), .Z(n244) );
  INV_X1 U53 ( .A(N10), .ZN(n251) );
  BUF_X1 U54 ( .A(N12), .Z(n241) );
  NOR3_X1 U55 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U56 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U57 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U58 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U59 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U60 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U61 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U62 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U63 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U64 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U65 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U67 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U69 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U70 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U71 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U72 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U73 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U74 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U75 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U76 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U77 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U79 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U81 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U82 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U83 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U84 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U85 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U86 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U87 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U88 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U89 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U90 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U91 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U92 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U93 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U94 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U95 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U96 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U97 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U98 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U99 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U100 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U101 ( .A(n983), .ZN(n701) );
  AOI22_X1 U102 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U103 ( .A(n982), .ZN(n700) );
  AOI22_X1 U104 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U105 ( .A(n981), .ZN(n699) );
  AOI22_X1 U106 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U107 ( .A(n980), .ZN(n698) );
  AOI22_X1 U108 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U109 ( .A(n910), .ZN(n637) );
  AOI22_X1 U110 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U111 ( .A(n909), .ZN(n636) );
  AOI22_X1 U112 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U113 ( .A(n908), .ZN(n635) );
  AOI22_X1 U114 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U115 ( .A(n907), .ZN(n634) );
  AOI22_X1 U116 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U117 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U118 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U119 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U120 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U121 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U122 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U123 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U124 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U125 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U126 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U127 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U128 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U129 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U130 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U131 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U132 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U133 ( .A(n988), .ZN(n705) );
  AOI22_X1 U134 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U135 ( .A(n986), .ZN(n704) );
  AOI22_X1 U136 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U137 ( .A(n985), .ZN(n703) );
  AOI22_X1 U138 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U139 ( .A(n984), .ZN(n702) );
  AOI22_X1 U140 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U141 ( .A(n951), .ZN(n673) );
  AOI22_X1 U142 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U143 ( .A(n949), .ZN(n672) );
  AOI22_X1 U144 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U145 ( .A(n948), .ZN(n671) );
  AOI22_X1 U146 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U147 ( .A(n947), .ZN(n670) );
  AOI22_X1 U148 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U149 ( .A(n946), .ZN(n669) );
  AOI22_X1 U150 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U151 ( .A(n945), .ZN(n668) );
  AOI22_X1 U152 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U153 ( .A(n944), .ZN(n667) );
  AOI22_X1 U154 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U155 ( .A(n943), .ZN(n666) );
  AOI22_X1 U156 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U157 ( .A(n915), .ZN(n641) );
  AOI22_X1 U158 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U159 ( .A(n913), .ZN(n640) );
  AOI22_X1 U160 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U161 ( .A(n912), .ZN(n639) );
  AOI22_X1 U162 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U163 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U164 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U165 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U166 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U167 ( .A(n911), .ZN(n638) );
  AOI22_X1 U168 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U169 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U170 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U171 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U172 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U173 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U174 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U175 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U176 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U177 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U178 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U179 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U180 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U181 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U182 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U183 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U184 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U185 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U186 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U187 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U188 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U189 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U190 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U191 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U192 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U193 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U194 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U195 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U196 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U197 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U198 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U199 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U200 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U201 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U202 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U203 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U204 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U205 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U206 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U207 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U208 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U209 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U210 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U211 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U212 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U213 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U214 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U215 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U216 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U217 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U218 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U219 ( .A(n999), .ZN(n715) );
  AOI22_X1 U220 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U221 ( .A(n998), .ZN(n714) );
  AOI22_X1 U222 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U223 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U224 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U225 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U226 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U227 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U228 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U229 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U230 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U231 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U232 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U233 ( .A(n979), .ZN(n697) );
  AOI22_X1 U234 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U235 ( .A(n977), .ZN(n696) );
  AOI22_X1 U236 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U237 ( .A(n976), .ZN(n695) );
  AOI22_X1 U238 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U239 ( .A(n975), .ZN(n694) );
  AOI22_X1 U240 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U241 ( .A(n974), .ZN(n693) );
  AOI22_X1 U242 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U243 ( .A(n973), .ZN(n692) );
  AOI22_X1 U244 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U245 ( .A(n972), .ZN(n691) );
  AOI22_X1 U246 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U247 ( .A(n971), .ZN(n690) );
  AOI22_X1 U248 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U249 ( .A(n970), .ZN(n689) );
  AOI22_X1 U250 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U251 ( .A(n968), .ZN(n688) );
  AOI22_X1 U252 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U253 ( .A(n967), .ZN(n687) );
  AOI22_X1 U254 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U255 ( .A(n966), .ZN(n686) );
  AOI22_X1 U256 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U257 ( .A(n965), .ZN(n685) );
  AOI22_X1 U258 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U259 ( .A(n964), .ZN(n684) );
  AOI22_X1 U260 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U261 ( .A(n963), .ZN(n683) );
  AOI22_X1 U262 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U263 ( .A(n962), .ZN(n682) );
  AOI22_X1 U264 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U265 ( .A(n942), .ZN(n665) );
  AOI22_X1 U266 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U267 ( .A(n940), .ZN(n664) );
  AOI22_X1 U268 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U269 ( .A(n939), .ZN(n663) );
  AOI22_X1 U270 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U271 ( .A(n935), .ZN(n659) );
  AOI22_X1 U272 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U273 ( .A(n934), .ZN(n658) );
  AOI22_X1 U274 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U275 ( .A(n933), .ZN(n657) );
  AOI22_X1 U276 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U277 ( .A(n931), .ZN(n656) );
  AOI22_X1 U278 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U279 ( .A(n930), .ZN(n655) );
  AOI22_X1 U280 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U281 ( .A(n929), .ZN(n654) );
  AOI22_X1 U282 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U283 ( .A(n928), .ZN(n653) );
  AOI22_X1 U284 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U285 ( .A(n927), .ZN(n652) );
  AOI22_X1 U286 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U287 ( .A(n926), .ZN(n651) );
  AOI22_X1 U288 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U289 ( .A(n925), .ZN(n650) );
  AOI22_X1 U290 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U291 ( .A(n906), .ZN(n633) );
  AOI22_X1 U292 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U293 ( .A(n904), .ZN(n632) );
  AOI22_X1 U294 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U295 ( .A(n903), .ZN(n631) );
  AOI22_X1 U296 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U297 ( .A(n902), .ZN(n630) );
  AOI22_X1 U298 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U299 ( .A(n901), .ZN(n629) );
  AOI22_X1 U300 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U301 ( .A(n900), .ZN(n628) );
  AOI22_X1 U302 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U303 ( .A(n899), .ZN(n627) );
  AOI22_X1 U304 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U305 ( .A(n898), .ZN(n626) );
  AOI22_X1 U306 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U307 ( .A(n897), .ZN(n625) );
  AOI22_X1 U308 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U309 ( .A(n895), .ZN(n624) );
  AOI22_X1 U310 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U311 ( .A(n894), .ZN(n623) );
  AOI22_X1 U312 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U313 ( .A(n893), .ZN(n622) );
  AOI22_X1 U314 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U315 ( .A(n892), .ZN(n621) );
  AOI22_X1 U316 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U317 ( .A(n891), .ZN(n620) );
  AOI22_X1 U318 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U319 ( .A(n890), .ZN(n619) );
  AOI22_X1 U320 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U321 ( .A(n889), .ZN(n618) );
  AOI22_X1 U322 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U323 ( .A(n938), .ZN(n662) );
  AOI22_X1 U324 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U325 ( .A(n937), .ZN(n661) );
  AOI22_X1 U326 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U327 ( .A(n936), .ZN(n660) );
  AOI22_X1 U328 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U329 ( .A(N12), .ZN(n253) );
  INV_X1 U330 ( .A(N11), .ZN(n252) );
  INV_X1 U331 ( .A(n997), .ZN(n713) );
  AOI22_X1 U332 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U333 ( .A(n995), .ZN(n712) );
  AOI22_X1 U334 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U335 ( .A(n994), .ZN(n711) );
  AOI22_X1 U336 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U337 ( .A(n993), .ZN(n710) );
  AOI22_X1 U338 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U339 ( .A(n992), .ZN(n709) );
  AOI22_X1 U340 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U341 ( .A(n991), .ZN(n708) );
  AOI22_X1 U342 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U343 ( .A(n990), .ZN(n707) );
  AOI22_X1 U344 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U345 ( .A(n989), .ZN(n706) );
  AOI22_X1 U346 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U347 ( .A(n924), .ZN(n649) );
  AOI22_X1 U348 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U349 ( .A(n922), .ZN(n648) );
  AOI22_X1 U350 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U351 ( .A(n921), .ZN(n647) );
  AOI22_X1 U352 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U353 ( .A(n920), .ZN(n646) );
  AOI22_X1 U354 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U355 ( .A(n919), .ZN(n645) );
  AOI22_X1 U356 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U357 ( .A(n918), .ZN(n644) );
  AOI22_X1 U358 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U359 ( .A(n917), .ZN(n643) );
  AOI22_X1 U360 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U361 ( .A(n916), .ZN(n642) );
  AOI22_X1 U362 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U363 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U364 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U365 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U366 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U367 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U368 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U369 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U370 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U371 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U372 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U373 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U374 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U375 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U376 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U377 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U378 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U379 ( .A(n961), .ZN(n681) );
  AOI22_X1 U380 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U381 ( .A(n959), .ZN(n680) );
  AOI22_X1 U382 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U383 ( .A(n958), .ZN(n679) );
  AOI22_X1 U384 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U385 ( .A(n957), .ZN(n678) );
  AOI22_X1 U386 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U387 ( .A(n956), .ZN(n677) );
  AOI22_X1 U388 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U389 ( .A(n955), .ZN(n676) );
  AOI22_X1 U390 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U391 ( .A(n954), .ZN(n675) );
  AOI22_X1 U392 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U393 ( .A(n953), .ZN(n674) );
  AOI22_X1 U394 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U395 ( .A(n888), .ZN(n617) );
  AOI22_X1 U396 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U397 ( .A(n886), .ZN(n616) );
  AOI22_X1 U398 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U399 ( .A(n885), .ZN(n615) );
  AOI22_X1 U400 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U401 ( .A(n884), .ZN(n614) );
  AOI22_X1 U402 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U403 ( .A(n883), .ZN(n613) );
  AOI22_X1 U404 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U405 ( .A(n882), .ZN(n612) );
  AOI22_X1 U406 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U407 ( .A(n881), .ZN(n611) );
  AOI22_X1 U408 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U409 ( .A(n880), .ZN(n610) );
  AOI22_X1 U410 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U411 ( .A(n879), .ZN(n609) );
  AOI22_X1 U412 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U413 ( .A(n877), .ZN(n608) );
  AOI22_X1 U414 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U415 ( .A(n876), .ZN(n607) );
  AOI22_X1 U416 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U417 ( .A(n875), .ZN(n606) );
  AOI22_X1 U418 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U419 ( .A(n874), .ZN(n605) );
  AOI22_X1 U420 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U421 ( .A(n873), .ZN(n604) );
  AOI22_X1 U422 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U423 ( .A(n872), .ZN(n603) );
  AOI22_X1 U424 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U425 ( .A(n871), .ZN(n602) );
  AOI22_X1 U426 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U427 ( .A(n870), .ZN(n601) );
  AOI22_X1 U428 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U429 ( .A(n868), .ZN(n600) );
  AOI22_X1 U430 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U431 ( .A(n867), .ZN(n599) );
  AOI22_X1 U432 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U433 ( .A(n866), .ZN(n598) );
  AOI22_X1 U434 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U435 ( .A(n865), .ZN(n597) );
  AOI22_X1 U436 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U437 ( .A(n864), .ZN(n596) );
  AOI22_X1 U438 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U439 ( .A(n863), .ZN(n595) );
  AOI22_X1 U440 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U441 ( .A(n862), .ZN(n594) );
  AOI22_X1 U442 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U443 ( .A(n861), .ZN(n293) );
  AOI22_X1 U444 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U445 ( .A(n859), .ZN(n292) );
  AOI22_X1 U446 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U447 ( .A(n858), .ZN(n291) );
  AOI22_X1 U448 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U449 ( .A(n857), .ZN(n290) );
  AOI22_X1 U450 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U451 ( .A(n856), .ZN(n289) );
  AOI22_X1 U452 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U453 ( .A(n855), .ZN(n288) );
  AOI22_X1 U454 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U455 ( .A(n854), .ZN(n287) );
  AOI22_X1 U456 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U457 ( .A(n853), .ZN(n286) );
  AOI22_X1 U458 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U459 ( .A(n852), .ZN(n285) );
  AOI22_X1 U460 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U461 ( .A(n850), .ZN(n284) );
  AOI22_X1 U462 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U463 ( .A(n849), .ZN(n283) );
  AOI22_X1 U464 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U465 ( .A(n848), .ZN(n282) );
  AOI22_X1 U466 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U467 ( .A(n847), .ZN(n281) );
  AOI22_X1 U468 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U469 ( .A(n846), .ZN(n280) );
  AOI22_X1 U470 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U471 ( .A(n845), .ZN(n279) );
  AOI22_X1 U472 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U473 ( .A(n844), .ZN(n278) );
  AOI22_X1 U474 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U475 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U476 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U477 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U478 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U479 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U480 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U481 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U482 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U483 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U484 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U485 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U486 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U487 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U488 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U489 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U490 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U491 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U492 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U493 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U494 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U495 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U496 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U497 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U498 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U499 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U500 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U501 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U502 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U503 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U504 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U505 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U506 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U507 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U508 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U509 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U510 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U511 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U512 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U513 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U514 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U515 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U516 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U517 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U518 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U519 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U520 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U521 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U522 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U523 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U524 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U525 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U526 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U527 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U528 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U529 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U530 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U531 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U532 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U533 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U534 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U535 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U536 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U537 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U538 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U539 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U540 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U541 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U542 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U543 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U544 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U545 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U546 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U547 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U548 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U549 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U550 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U551 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U552 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U553 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U554 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U555 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U556 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U557 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U558 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U559 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U560 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U561 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U562 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U563 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U564 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U565 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U566 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U567 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U568 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U569 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U570 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U571 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U572 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U573 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U574 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U575 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U576 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U577 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U578 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U579 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U580 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U581 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U582 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U583 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U584 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U585 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U586 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U587 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U588 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U589 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U590 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U591 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U592 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U593 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U594 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U595 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U596 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U597 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U598 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U599 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U600 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U601 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U602 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U603 ( .A(N13), .ZN(n842) );
  INV_X1 U604 ( .A(N14), .ZN(n843) );
  MUX2_X1 U605 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n245), .Z(n1) );
  MUX2_X1 U606 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n245), .Z(n2) );
  MUX2_X1 U607 ( .A(n2), .B(n1), .S(n242), .Z(n3) );
  MUX2_X1 U608 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n245), .Z(n4) );
  MUX2_X1 U609 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n245), .Z(n5) );
  MUX2_X1 U610 ( .A(n5), .B(n4), .S(n244), .Z(n6) );
  MUX2_X1 U611 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U612 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n245), .Z(n8) );
  MUX2_X1 U613 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n245), .Z(n9) );
  MUX2_X1 U614 ( .A(n9), .B(n8), .S(n243), .Z(n10) );
  MUX2_X1 U615 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n245), .Z(n11) );
  MUX2_X1 U616 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n245), .Z(n12) );
  MUX2_X1 U617 ( .A(n12), .B(n11), .S(n243), .Z(n13) );
  MUX2_X1 U618 ( .A(n13), .B(n10), .S(n241), .Z(n14) );
  MUX2_X1 U619 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U620 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n247), .Z(n16) );
  MUX2_X1 U621 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(N10), .Z(n17) );
  MUX2_X1 U622 ( .A(n17), .B(n16), .S(n242), .Z(n18) );
  MUX2_X1 U623 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n248), .Z(n19) );
  MUX2_X1 U624 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n20) );
  MUX2_X1 U625 ( .A(n20), .B(n19), .S(n242), .Z(n21) );
  MUX2_X1 U626 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U627 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(N10), .Z(n23) );
  MUX2_X1 U628 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(N10), .Z(n24) );
  MUX2_X1 U629 ( .A(n24), .B(n23), .S(n242), .Z(n25) );
  MUX2_X1 U630 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(N10), .Z(n26) );
  MUX2_X1 U631 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n27) );
  MUX2_X1 U632 ( .A(n27), .B(n26), .S(n242), .Z(n28) );
  MUX2_X1 U633 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U634 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U635 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U636 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n246), .Z(n31) );
  MUX2_X1 U637 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n249), .Z(n32) );
  MUX2_X1 U638 ( .A(n32), .B(n31), .S(n242), .Z(n33) );
  MUX2_X1 U639 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(N10), .Z(n34) );
  MUX2_X1 U640 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n250), .Z(n35) );
  MUX2_X1 U641 ( .A(n35), .B(n34), .S(n242), .Z(n36) );
  MUX2_X1 U642 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U643 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n245), .Z(n38) );
  MUX2_X1 U644 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(N10), .Z(n39) );
  MUX2_X1 U645 ( .A(n39), .B(n38), .S(n242), .Z(n40) );
  MUX2_X1 U646 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(N10), .Z(n41) );
  MUX2_X1 U647 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n250), .Z(n42) );
  MUX2_X1 U648 ( .A(n42), .B(n41), .S(n242), .Z(n43) );
  MUX2_X1 U649 ( .A(n43), .B(n40), .S(N12), .Z(n44) );
  MUX2_X1 U650 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U651 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n245), .Z(n46) );
  MUX2_X1 U652 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(N10), .Z(n47) );
  MUX2_X1 U653 ( .A(n47), .B(n46), .S(n242), .Z(n48) );
  MUX2_X1 U654 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n245), .Z(n49) );
  MUX2_X1 U655 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n245), .Z(n50) );
  MUX2_X1 U656 ( .A(n50), .B(n49), .S(n242), .Z(n51) );
  MUX2_X1 U657 ( .A(n51), .B(n48), .S(N12), .Z(n52) );
  MUX2_X1 U658 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n245), .Z(n53) );
  MUX2_X1 U659 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n249), .Z(n54) );
  MUX2_X1 U660 ( .A(n54), .B(n53), .S(n242), .Z(n55) );
  MUX2_X1 U661 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n250), .Z(n56) );
  MUX2_X1 U662 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(N10), .Z(n57) );
  MUX2_X1 U663 ( .A(n57), .B(n56), .S(n242), .Z(n58) );
  MUX2_X1 U664 ( .A(n58), .B(n55), .S(N12), .Z(n59) );
  MUX2_X1 U665 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U666 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U667 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n246), .Z(n61) );
  MUX2_X1 U668 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n246), .Z(n62) );
  MUX2_X1 U669 ( .A(n62), .B(n61), .S(n243), .Z(n63) );
  MUX2_X1 U670 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n246), .Z(n64) );
  MUX2_X1 U671 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n246), .Z(n65) );
  MUX2_X1 U672 ( .A(n65), .B(n64), .S(n243), .Z(n66) );
  MUX2_X1 U673 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U674 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n246), .Z(n68) );
  MUX2_X1 U675 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n246), .Z(n69) );
  MUX2_X1 U676 ( .A(n69), .B(n68), .S(n243), .Z(n70) );
  MUX2_X1 U677 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n246), .Z(n71) );
  MUX2_X1 U678 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n246), .Z(n72) );
  MUX2_X1 U679 ( .A(n72), .B(n71), .S(n243), .Z(n73) );
  MUX2_X1 U680 ( .A(n73), .B(n70), .S(n241), .Z(n74) );
  MUX2_X1 U681 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U682 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n246), .Z(n76) );
  MUX2_X1 U683 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n246), .Z(n77) );
  MUX2_X1 U684 ( .A(n77), .B(n76), .S(n243), .Z(n78) );
  MUX2_X1 U685 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n246), .Z(n79) );
  MUX2_X1 U686 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n246), .Z(n80) );
  MUX2_X1 U687 ( .A(n80), .B(n79), .S(n243), .Z(n81) );
  MUX2_X1 U688 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U689 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n247), .Z(n83) );
  MUX2_X1 U690 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n247), .Z(n84) );
  MUX2_X1 U691 ( .A(n84), .B(n83), .S(n243), .Z(n85) );
  MUX2_X1 U692 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n247), .Z(n86) );
  MUX2_X1 U693 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n247), .Z(n87) );
  MUX2_X1 U694 ( .A(n87), .B(n86), .S(n243), .Z(n88) );
  MUX2_X1 U695 ( .A(n88), .B(n85), .S(n241), .Z(n89) );
  MUX2_X1 U696 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U697 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U698 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n247), .Z(n91) );
  MUX2_X1 U699 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n247), .Z(n92) );
  MUX2_X1 U700 ( .A(n92), .B(n91), .S(n243), .Z(n93) );
  MUX2_X1 U701 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n247), .Z(n94) );
  MUX2_X1 U702 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n247), .Z(n95) );
  MUX2_X1 U703 ( .A(n95), .B(n94), .S(n243), .Z(n96) );
  MUX2_X1 U704 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U705 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n247), .Z(n98) );
  MUX2_X1 U706 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n247), .Z(n99) );
  MUX2_X1 U707 ( .A(n99), .B(n98), .S(n243), .Z(n100) );
  MUX2_X1 U708 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n247), .Z(n101) );
  MUX2_X1 U709 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n247), .Z(n102) );
  MUX2_X1 U710 ( .A(n102), .B(n101), .S(n243), .Z(n103) );
  MUX2_X1 U711 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U712 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U713 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n247), .Z(n106) );
  MUX2_X1 U714 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n250), .Z(n107) );
  MUX2_X1 U715 ( .A(n107), .B(n106), .S(n244), .Z(n108) );
  MUX2_X1 U716 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n248), .Z(n109) );
  MUX2_X1 U717 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n250), .Z(n110) );
  MUX2_X1 U718 ( .A(n110), .B(n109), .S(n244), .Z(n111) );
  MUX2_X1 U719 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U720 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n250), .Z(n113) );
  MUX2_X1 U721 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n250), .Z(n114) );
  MUX2_X1 U722 ( .A(n114), .B(n113), .S(n244), .Z(n115) );
  MUX2_X1 U723 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n250), .Z(n116) );
  MUX2_X1 U724 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n250), .Z(n117) );
  MUX2_X1 U725 ( .A(n117), .B(n116), .S(n244), .Z(n118) );
  MUX2_X1 U726 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U727 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U728 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U729 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n250), .Z(n121) );
  MUX2_X1 U730 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n248), .Z(n122) );
  MUX2_X1 U731 ( .A(n122), .B(n121), .S(n244), .Z(n123) );
  MUX2_X1 U732 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n250), .Z(n124) );
  MUX2_X1 U733 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n247), .Z(n125) );
  MUX2_X1 U734 ( .A(n125), .B(n124), .S(n244), .Z(n126) );
  MUX2_X1 U735 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U736 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(N10), .Z(n128) );
  MUX2_X1 U737 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n250), .Z(n129) );
  MUX2_X1 U738 ( .A(n129), .B(n128), .S(n244), .Z(n130) );
  MUX2_X1 U739 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n245), .Z(n131) );
  MUX2_X1 U740 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n250), .Z(n132) );
  MUX2_X1 U741 ( .A(n132), .B(n131), .S(n244), .Z(n133) );
  MUX2_X1 U742 ( .A(n133), .B(n130), .S(n241), .Z(n134) );
  MUX2_X1 U743 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U744 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n250), .Z(n136) );
  MUX2_X1 U745 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n249), .Z(n137) );
  MUX2_X1 U746 ( .A(n137), .B(n136), .S(n244), .Z(n138) );
  MUX2_X1 U747 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(N10), .Z(n139) );
  MUX2_X1 U748 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n250), .Z(n140) );
  MUX2_X1 U749 ( .A(n140), .B(n139), .S(n244), .Z(n141) );
  MUX2_X1 U750 ( .A(n141), .B(n138), .S(n241), .Z(n142) );
  MUX2_X1 U751 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n250), .Z(n143) );
  MUX2_X1 U752 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n250), .Z(n144) );
  MUX2_X1 U753 ( .A(n144), .B(n143), .S(n244), .Z(n145) );
  MUX2_X1 U754 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n250), .Z(n146) );
  MUX2_X1 U755 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n250), .Z(n147) );
  MUX2_X1 U756 ( .A(n147), .B(n146), .S(n244), .Z(n148) );
  MUX2_X1 U757 ( .A(n148), .B(n145), .S(n241), .Z(n149) );
  MUX2_X1 U758 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U759 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U760 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n246), .Z(n151) );
  MUX2_X1 U761 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n246), .Z(n152) );
  MUX2_X1 U762 ( .A(n152), .B(n151), .S(n243), .Z(n153) );
  MUX2_X1 U763 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n246), .Z(n154) );
  MUX2_X1 U764 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n246), .Z(n155) );
  MUX2_X1 U765 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U766 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U767 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n246), .Z(n158) );
  MUX2_X1 U768 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n246), .Z(n159) );
  MUX2_X1 U769 ( .A(n159), .B(n158), .S(N11), .Z(n160) );
  MUX2_X1 U770 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n246), .Z(n161) );
  MUX2_X1 U771 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n250), .Z(n162) );
  MUX2_X1 U772 ( .A(n162), .B(n161), .S(N11), .Z(n163) );
  MUX2_X1 U773 ( .A(n163), .B(n160), .S(n241), .Z(n164) );
  MUX2_X1 U774 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U775 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n246), .Z(n166) );
  MUX2_X1 U776 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(N10), .Z(n167) );
  MUX2_X1 U777 ( .A(n167), .B(n166), .S(n244), .Z(n168) );
  MUX2_X1 U778 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n246), .Z(n169) );
  MUX2_X1 U779 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n246), .Z(n170) );
  MUX2_X1 U780 ( .A(n170), .B(n169), .S(N11), .Z(n171) );
  MUX2_X1 U781 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U782 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n248), .Z(n173) );
  MUX2_X1 U783 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n248), .Z(n174) );
  MUX2_X1 U784 ( .A(n174), .B(n173), .S(N11), .Z(n175) );
  MUX2_X1 U785 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n248), .Z(n176) );
  MUX2_X1 U786 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n248), .Z(n177) );
  MUX2_X1 U787 ( .A(n177), .B(n176), .S(N11), .Z(n178) );
  MUX2_X1 U788 ( .A(n178), .B(n175), .S(n241), .Z(n179) );
  MUX2_X1 U789 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U790 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U791 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n248), .Z(n181) );
  MUX2_X1 U792 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n248), .Z(n182) );
  MUX2_X1 U793 ( .A(n182), .B(n181), .S(N11), .Z(n183) );
  MUX2_X1 U794 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n248), .Z(n184) );
  MUX2_X1 U795 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n248), .Z(n185) );
  MUX2_X1 U796 ( .A(n185), .B(n184), .S(n242), .Z(n186) );
  MUX2_X1 U797 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U798 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n248), .Z(n188) );
  MUX2_X1 U799 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n248), .Z(n189) );
  MUX2_X1 U800 ( .A(n189), .B(n188), .S(N11), .Z(n190) );
  MUX2_X1 U801 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n248), .Z(n191) );
  MUX2_X1 U802 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n248), .Z(n192) );
  MUX2_X1 U803 ( .A(n192), .B(n191), .S(n243), .Z(n193) );
  MUX2_X1 U804 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U805 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U806 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n249), .Z(n196) );
  MUX2_X1 U807 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n249), .Z(n197) );
  MUX2_X1 U808 ( .A(n197), .B(n196), .S(n242), .Z(n198) );
  MUX2_X1 U809 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n249), .Z(n199) );
  MUX2_X1 U810 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n249), .Z(n200) );
  MUX2_X1 U811 ( .A(n200), .B(n199), .S(n243), .Z(n201) );
  MUX2_X1 U812 ( .A(n201), .B(n198), .S(N12), .Z(n202) );
  MUX2_X1 U813 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n249), .Z(n203) );
  MUX2_X1 U814 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n249), .Z(n204) );
  MUX2_X1 U815 ( .A(n204), .B(n203), .S(n244), .Z(n205) );
  MUX2_X1 U816 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n249), .Z(n206) );
  MUX2_X1 U817 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n249), .Z(n207) );
  MUX2_X1 U818 ( .A(n207), .B(n206), .S(N11), .Z(n208) );
  MUX2_X1 U819 ( .A(n208), .B(n205), .S(N12), .Z(n209) );
  MUX2_X1 U820 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U821 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U822 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n249), .Z(n211) );
  MUX2_X1 U823 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n249), .Z(n212) );
  MUX2_X1 U824 ( .A(n212), .B(n211), .S(N11), .Z(n213) );
  MUX2_X1 U825 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n249), .Z(n214) );
  MUX2_X1 U826 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n249), .Z(n215) );
  MUX2_X1 U827 ( .A(n215), .B(n214), .S(n242), .Z(n216) );
  MUX2_X1 U828 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U829 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n247), .Z(n218) );
  MUX2_X1 U830 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n249), .Z(n219) );
  MUX2_X1 U831 ( .A(n219), .B(n218), .S(n244), .Z(n220) );
  MUX2_X1 U832 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n245), .Z(n221) );
  MUX2_X1 U833 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n249), .Z(n222) );
  MUX2_X1 U834 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U835 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U836 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U837 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n248), .Z(n226) );
  MUX2_X1 U838 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n249), .Z(n227) );
  MUX2_X1 U839 ( .A(n227), .B(n226), .S(N11), .Z(n228) );
  MUX2_X1 U840 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n247), .Z(n229) );
  MUX2_X1 U841 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n248), .Z(n230) );
  MUX2_X1 U842 ( .A(n230), .B(n229), .S(n242), .Z(n231) );
  MUX2_X1 U843 ( .A(n231), .B(n228), .S(N12), .Z(n232) );
  MUX2_X1 U844 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n248), .Z(n233) );
  MUX2_X1 U845 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n249), .Z(n234) );
  MUX2_X1 U846 ( .A(n234), .B(n233), .S(n244), .Z(n235) );
  MUX2_X1 U847 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n245), .Z(n236) );
  MUX2_X1 U848 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n247), .Z(n237) );
  MUX2_X1 U849 ( .A(n237), .B(n236), .S(N11), .Z(n238) );
  MUX2_X1 U850 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U851 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U852 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U853 ( .A(n250), .Z(n245) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_8 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  BUF_X1 U3 ( .A(N10), .Z(n247) );
  BUF_X1 U4 ( .A(n250), .Z(n248) );
  BUF_X1 U5 ( .A(n250), .Z(n249) );
  BUF_X1 U6 ( .A(n250), .Z(n246) );
  BUF_X1 U7 ( .A(n250), .Z(n245) );
  BUF_X1 U8 ( .A(N10), .Z(n250) );
  INV_X1 U9 ( .A(n1111), .ZN(n841) );
  INV_X1 U10 ( .A(n1100), .ZN(n840) );
  INV_X1 U11 ( .A(n1090), .ZN(n839) );
  INV_X1 U12 ( .A(n1080), .ZN(n838) );
  INV_X1 U13 ( .A(n1070), .ZN(n837) );
  INV_X1 U14 ( .A(n1060), .ZN(n836) );
  INV_X1 U15 ( .A(n1051), .ZN(n835) );
  INV_X1 U16 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U19 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U20 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U21 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U22 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U23 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U24 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U26 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U27 ( .A(n1131), .ZN(n816) );
  INV_X1 U28 ( .A(n1121), .ZN(n815) );
  INV_X1 U29 ( .A(n887), .ZN(n814) );
  INV_X1 U30 ( .A(n878), .ZN(n813) );
  INV_X1 U31 ( .A(n869), .ZN(n812) );
  INV_X1 U32 ( .A(n860), .ZN(n811) );
  INV_X1 U33 ( .A(n851), .ZN(n810) );
  INV_X1 U34 ( .A(n987), .ZN(n828) );
  INV_X1 U35 ( .A(n978), .ZN(n827) );
  INV_X1 U36 ( .A(n969), .ZN(n826) );
  INV_X1 U37 ( .A(n914), .ZN(n820) );
  INV_X1 U38 ( .A(n905), .ZN(n819) );
  INV_X1 U39 ( .A(n896), .ZN(n818) );
  INV_X1 U40 ( .A(n1033), .ZN(n833) );
  INV_X1 U41 ( .A(n1023), .ZN(n832) );
  INV_X1 U42 ( .A(n1014), .ZN(n831) );
  INV_X1 U43 ( .A(n1005), .ZN(n830) );
  INV_X1 U44 ( .A(n996), .ZN(n829) );
  INV_X1 U45 ( .A(n960), .ZN(n825) );
  INV_X1 U46 ( .A(n950), .ZN(n824) );
  INV_X1 U47 ( .A(n941), .ZN(n823) );
  INV_X1 U48 ( .A(n932), .ZN(n822) );
  INV_X1 U49 ( .A(n923), .ZN(n821) );
  INV_X1 U50 ( .A(n1142), .ZN(n817) );
  BUF_X1 U51 ( .A(N11), .Z(n242) );
  BUF_X1 U52 ( .A(N11), .Z(n243) );
  BUF_X1 U53 ( .A(N11), .Z(n244) );
  INV_X1 U54 ( .A(N10), .ZN(n251) );
  BUF_X1 U55 ( .A(N12), .Z(n241) );
  NOR3_X1 U56 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U57 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U58 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U60 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U62 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U63 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U64 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U65 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U67 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U69 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U70 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U71 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U72 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U73 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U74 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U75 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U76 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U77 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U79 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U81 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U82 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U83 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U84 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U85 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U86 ( .A1(n843), .A2(n842), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U88 ( .A1(N13), .A2(n842), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U89 ( .A1(N14), .A2(n843), .A3(wr_en), .ZN(n952) );
  INV_X1 U90 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U92 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U94 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U95 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U96 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U97 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U98 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U99 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U100 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U101 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U102 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U103 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U104 ( .A(n983), .ZN(n701) );
  AOI22_X1 U105 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U106 ( .A(n982), .ZN(n700) );
  AOI22_X1 U107 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U108 ( .A(n981), .ZN(n699) );
  AOI22_X1 U109 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U110 ( .A(n980), .ZN(n698) );
  AOI22_X1 U111 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U112 ( .A(n910), .ZN(n637) );
  AOI22_X1 U113 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U114 ( .A(n909), .ZN(n636) );
  AOI22_X1 U115 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U116 ( .A(n908), .ZN(n635) );
  AOI22_X1 U117 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U118 ( .A(n907), .ZN(n634) );
  AOI22_X1 U119 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U120 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U121 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U122 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U123 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U124 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U125 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U126 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U127 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U128 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U129 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U130 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U131 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U132 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U133 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U134 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U135 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U136 ( .A(n988), .ZN(n705) );
  AOI22_X1 U137 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U138 ( .A(n986), .ZN(n704) );
  AOI22_X1 U139 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U140 ( .A(n985), .ZN(n703) );
  AOI22_X1 U141 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U142 ( .A(n984), .ZN(n702) );
  AOI22_X1 U143 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U144 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U145 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U146 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U147 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U148 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U149 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U150 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U151 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U152 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U153 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U154 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U155 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U156 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U157 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U158 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U159 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U160 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U161 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U162 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U163 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U164 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U165 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U166 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U167 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U168 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U169 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U170 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U171 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U172 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U173 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U174 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U175 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U176 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U177 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U178 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U179 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U180 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U181 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U182 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U183 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U184 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U185 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U186 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U187 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U188 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U189 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U190 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U191 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U192 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U193 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U194 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U195 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U196 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U197 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U198 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U199 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U200 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U201 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U202 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U203 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U204 ( .A(n999), .ZN(n715) );
  AOI22_X1 U205 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U206 ( .A(n998), .ZN(n714) );
  AOI22_X1 U207 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U208 ( .A(n951), .ZN(n673) );
  AOI22_X1 U209 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U210 ( .A(n949), .ZN(n672) );
  AOI22_X1 U211 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U212 ( .A(n948), .ZN(n671) );
  AOI22_X1 U213 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U214 ( .A(n947), .ZN(n670) );
  AOI22_X1 U215 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U216 ( .A(n946), .ZN(n669) );
  AOI22_X1 U217 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U218 ( .A(n945), .ZN(n668) );
  AOI22_X1 U219 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U220 ( .A(n943), .ZN(n666) );
  AOI22_X1 U221 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U222 ( .A(n915), .ZN(n641) );
  AOI22_X1 U223 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U224 ( .A(n913), .ZN(n640) );
  AOI22_X1 U225 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U226 ( .A(n912), .ZN(n639) );
  AOI22_X1 U227 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U228 ( .A(n944), .ZN(n667) );
  AOI22_X1 U229 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U230 ( .A(n927), .ZN(n652) );
  AOI22_X1 U231 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U232 ( .A(n926), .ZN(n651) );
  AOI22_X1 U233 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U234 ( .A(n925), .ZN(n650) );
  AOI22_X1 U235 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U236 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U237 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U238 ( .A(n911), .ZN(n638) );
  AOI22_X1 U239 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U240 ( .A(n979), .ZN(n697) );
  AOI22_X1 U241 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U242 ( .A(n977), .ZN(n696) );
  AOI22_X1 U243 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U244 ( .A(n976), .ZN(n695) );
  AOI22_X1 U245 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U246 ( .A(n975), .ZN(n694) );
  AOI22_X1 U247 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U248 ( .A(n974), .ZN(n693) );
  AOI22_X1 U249 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U250 ( .A(n973), .ZN(n692) );
  AOI22_X1 U251 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U252 ( .A(n972), .ZN(n691) );
  AOI22_X1 U253 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U254 ( .A(n971), .ZN(n690) );
  AOI22_X1 U255 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U256 ( .A(n970), .ZN(n689) );
  AOI22_X1 U257 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U258 ( .A(n968), .ZN(n688) );
  AOI22_X1 U259 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U260 ( .A(n967), .ZN(n687) );
  AOI22_X1 U261 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U262 ( .A(n966), .ZN(n686) );
  AOI22_X1 U263 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U264 ( .A(n965), .ZN(n685) );
  AOI22_X1 U265 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U266 ( .A(n964), .ZN(n684) );
  AOI22_X1 U267 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U268 ( .A(n963), .ZN(n683) );
  AOI22_X1 U269 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U270 ( .A(n962), .ZN(n682) );
  AOI22_X1 U271 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U272 ( .A(n942), .ZN(n665) );
  AOI22_X1 U273 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U274 ( .A(n940), .ZN(n664) );
  AOI22_X1 U275 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U276 ( .A(n939), .ZN(n663) );
  AOI22_X1 U277 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U278 ( .A(n938), .ZN(n662) );
  AOI22_X1 U279 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U280 ( .A(n937), .ZN(n661) );
  AOI22_X1 U281 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U282 ( .A(n936), .ZN(n660) );
  AOI22_X1 U283 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U284 ( .A(n935), .ZN(n659) );
  AOI22_X1 U285 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U286 ( .A(n934), .ZN(n658) );
  AOI22_X1 U287 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U288 ( .A(n933), .ZN(n657) );
  AOI22_X1 U289 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U290 ( .A(n931), .ZN(n656) );
  AOI22_X1 U291 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U292 ( .A(n930), .ZN(n655) );
  AOI22_X1 U293 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U294 ( .A(n929), .ZN(n654) );
  AOI22_X1 U295 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U296 ( .A(n928), .ZN(n653) );
  AOI22_X1 U297 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U298 ( .A(n906), .ZN(n633) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U300 ( .A(n904), .ZN(n632) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U302 ( .A(n903), .ZN(n631) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U304 ( .A(n902), .ZN(n630) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U306 ( .A(n901), .ZN(n629) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U308 ( .A(n900), .ZN(n628) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U310 ( .A(n899), .ZN(n627) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U312 ( .A(n898), .ZN(n626) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U314 ( .A(n897), .ZN(n625) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U316 ( .A(n895), .ZN(n624) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U318 ( .A(n894), .ZN(n623) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U320 ( .A(n893), .ZN(n622) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U322 ( .A(n892), .ZN(n621) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U324 ( .A(n891), .ZN(n620) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U326 ( .A(n890), .ZN(n619) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U328 ( .A(n889), .ZN(n618) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U330 ( .A(N12), .ZN(n253) );
  INV_X1 U331 ( .A(N11), .ZN(n252) );
  INV_X1 U332 ( .A(n997), .ZN(n713) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U334 ( .A(n995), .ZN(n712) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U336 ( .A(n994), .ZN(n711) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U338 ( .A(n993), .ZN(n710) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U340 ( .A(n992), .ZN(n709) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U342 ( .A(n991), .ZN(n708) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U344 ( .A(n990), .ZN(n707) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U346 ( .A(n989), .ZN(n706) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U348 ( .A(n924), .ZN(n649) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U350 ( .A(n922), .ZN(n648) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U352 ( .A(n921), .ZN(n647) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U354 ( .A(n920), .ZN(n646) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U356 ( .A(n919), .ZN(n645) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U358 ( .A(n918), .ZN(n644) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U360 ( .A(n917), .ZN(n643) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U362 ( .A(n916), .ZN(n642) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U364 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U366 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U368 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U370 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U372 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U374 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U376 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U378 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U380 ( .A(n961), .ZN(n681) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U382 ( .A(n959), .ZN(n680) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U384 ( .A(n958), .ZN(n679) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U386 ( .A(n957), .ZN(n678) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U388 ( .A(n956), .ZN(n677) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U390 ( .A(n955), .ZN(n676) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U392 ( .A(n954), .ZN(n675) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U394 ( .A(n953), .ZN(n674) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U396 ( .A(n888), .ZN(n617) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U398 ( .A(n886), .ZN(n616) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U400 ( .A(n885), .ZN(n615) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U402 ( .A(n884), .ZN(n614) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U404 ( .A(n883), .ZN(n613) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U406 ( .A(n882), .ZN(n612) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U408 ( .A(n881), .ZN(n611) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U410 ( .A(n880), .ZN(n610) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U412 ( .A(n879), .ZN(n609) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U414 ( .A(n877), .ZN(n608) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U416 ( .A(n876), .ZN(n607) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U418 ( .A(n875), .ZN(n606) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U420 ( .A(n874), .ZN(n605) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U422 ( .A(n873), .ZN(n604) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U424 ( .A(n872), .ZN(n603) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U426 ( .A(n871), .ZN(n602) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U428 ( .A(n870), .ZN(n601) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U430 ( .A(n868), .ZN(n600) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U432 ( .A(n867), .ZN(n599) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U434 ( .A(n866), .ZN(n598) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U436 ( .A(n865), .ZN(n597) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U438 ( .A(n864), .ZN(n596) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U440 ( .A(n863), .ZN(n595) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U442 ( .A(n862), .ZN(n594) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U444 ( .A(n861), .ZN(n293) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U446 ( .A(n859), .ZN(n292) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U448 ( .A(n858), .ZN(n291) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U450 ( .A(n857), .ZN(n290) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U452 ( .A(n856), .ZN(n289) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U454 ( .A(n855), .ZN(n288) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U456 ( .A(n854), .ZN(n287) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U458 ( .A(n853), .ZN(n286) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U460 ( .A(n852), .ZN(n285) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U462 ( .A(n850), .ZN(n284) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U464 ( .A(n849), .ZN(n283) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U466 ( .A(n848), .ZN(n282) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U468 ( .A(n847), .ZN(n281) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U470 ( .A(n846), .ZN(n280) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U472 ( .A(n845), .ZN(n279) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U474 ( .A(n844), .ZN(n278) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U476 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U477 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U478 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U479 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U480 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U481 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U482 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U483 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U484 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U485 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U486 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U487 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U488 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U489 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U490 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U491 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U492 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U494 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U496 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U498 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U500 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U502 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U504 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U506 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U508 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U510 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U512 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U514 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U516 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U518 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U520 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U522 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U524 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U526 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U528 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U530 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U532 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U534 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U536 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U538 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U540 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U542 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U544 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U546 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U548 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U550 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U552 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U554 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U556 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U558 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U560 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U562 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U564 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U566 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U568 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U570 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U572 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U574 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U576 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U578 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U580 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U582 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U584 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U586 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U588 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U590 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U592 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U594 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U596 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U598 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U600 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U602 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U604 ( .A(N13), .ZN(n843) );
  INV_X1 U605 ( .A(N14), .ZN(n842) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n247), .Z(n1) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n247), .Z(n2) );
  MUX2_X1 U608 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n247), .Z(n4) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n247), .Z(n5) );
  MUX2_X1 U611 ( .A(n5), .B(n4), .S(n243), .Z(n6) );
  MUX2_X1 U612 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n247), .Z(n8) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n249), .Z(n9) );
  MUX2_X1 U615 ( .A(n9), .B(n8), .S(n242), .Z(n10) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n247), .Z(n11) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n248), .Z(n12) );
  MUX2_X1 U618 ( .A(n12), .B(n11), .S(n244), .Z(n13) );
  MUX2_X1 U619 ( .A(n13), .B(n10), .S(n241), .Z(n14) );
  MUX2_X1 U620 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n245), .Z(n16) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n245), .Z(n17) );
  MUX2_X1 U623 ( .A(n17), .B(n16), .S(n244), .Z(n18) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n245), .Z(n20) );
  MUX2_X1 U626 ( .A(n20), .B(n19), .S(N11), .Z(n21) );
  MUX2_X1 U627 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n245), .Z(n23) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n245), .Z(n24) );
  MUX2_X1 U630 ( .A(n24), .B(n23), .S(n243), .Z(n25) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n245), .Z(n26) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n245), .Z(n27) );
  MUX2_X1 U633 ( .A(n27), .B(n26), .S(N11), .Z(n28) );
  MUX2_X1 U634 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U635 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U636 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n245), .Z(n31) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n245), .Z(n32) );
  MUX2_X1 U639 ( .A(n32), .B(n31), .S(n243), .Z(n33) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U642 ( .A(n35), .B(n34), .S(n244), .Z(n36) );
  MUX2_X1 U643 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n246), .Z(n38) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n246), .Z(n39) );
  MUX2_X1 U646 ( .A(n39), .B(n38), .S(n243), .Z(n40) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n246), .Z(n41) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n246), .Z(n42) );
  MUX2_X1 U649 ( .A(n42), .B(n41), .S(N11), .Z(n43) );
  MUX2_X1 U650 ( .A(n43), .B(n40), .S(n241), .Z(n44) );
  MUX2_X1 U651 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n246), .Z(n46) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n246), .Z(n47) );
  MUX2_X1 U654 ( .A(n47), .B(n46), .S(n242), .Z(n48) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n246), .Z(n49) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n246), .Z(n50) );
  MUX2_X1 U657 ( .A(n50), .B(n49), .S(N11), .Z(n51) );
  MUX2_X1 U658 ( .A(n51), .B(n48), .S(n241), .Z(n52) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n246), .Z(n53) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n246), .Z(n54) );
  MUX2_X1 U661 ( .A(n54), .B(n53), .S(n242), .Z(n55) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n246), .Z(n56) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n246), .Z(n57) );
  MUX2_X1 U664 ( .A(n57), .B(n56), .S(N11), .Z(n58) );
  MUX2_X1 U665 ( .A(n58), .B(n55), .S(n241), .Z(n59) );
  MUX2_X1 U666 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U667 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n245), .Z(n61) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n245), .Z(n62) );
  MUX2_X1 U670 ( .A(n62), .B(n61), .S(N11), .Z(n63) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n246), .Z(n64) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n249), .Z(n65) );
  MUX2_X1 U673 ( .A(n65), .B(n64), .S(n243), .Z(n66) );
  MUX2_X1 U674 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n248), .Z(n68) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n246), .Z(n69) );
  MUX2_X1 U677 ( .A(n69), .B(n68), .S(n244), .Z(n70) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n246), .Z(n71) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n245), .Z(n72) );
  MUX2_X1 U680 ( .A(n72), .B(n71), .S(n242), .Z(n73) );
  MUX2_X1 U681 ( .A(n73), .B(n70), .S(N12), .Z(n74) );
  MUX2_X1 U682 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n248), .Z(n76) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n248), .Z(n77) );
  MUX2_X1 U685 ( .A(n77), .B(n76), .S(N11), .Z(n78) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n249), .Z(n79) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n248), .Z(n80) );
  MUX2_X1 U688 ( .A(n80), .B(n79), .S(N11), .Z(n81) );
  MUX2_X1 U689 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n250), .Z(n83) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n250), .Z(n84) );
  MUX2_X1 U692 ( .A(n84), .B(n83), .S(n244), .Z(n85) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n250), .Z(n86) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n246), .Z(n87) );
  MUX2_X1 U695 ( .A(n87), .B(n86), .S(n242), .Z(n88) );
  MUX2_X1 U696 ( .A(n88), .B(n85), .S(N12), .Z(n89) );
  MUX2_X1 U697 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U698 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n250), .Z(n91) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n92) );
  MUX2_X1 U701 ( .A(n92), .B(n91), .S(N11), .Z(n93) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n250), .Z(n95) );
  MUX2_X1 U704 ( .A(n95), .B(n94), .S(N11), .Z(n96) );
  MUX2_X1 U705 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n98) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n250), .Z(n99) );
  MUX2_X1 U708 ( .A(n99), .B(n98), .S(N11), .Z(n100) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n250), .Z(n101) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n250), .Z(n102) );
  MUX2_X1 U711 ( .A(n102), .B(n101), .S(N11), .Z(n103) );
  MUX2_X1 U712 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U713 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n247), .Z(n106) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n247), .Z(n107) );
  MUX2_X1 U716 ( .A(n107), .B(n106), .S(n242), .Z(n108) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n247), .Z(n109) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n247), .Z(n110) );
  MUX2_X1 U719 ( .A(n110), .B(n109), .S(n242), .Z(n111) );
  MUX2_X1 U720 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n247), .Z(n113) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n247), .Z(n114) );
  MUX2_X1 U723 ( .A(n114), .B(n113), .S(n242), .Z(n115) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n247), .Z(n116) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n247), .Z(n117) );
  MUX2_X1 U726 ( .A(n117), .B(n116), .S(n242), .Z(n118) );
  MUX2_X1 U727 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U728 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U729 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n247), .Z(n121) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n247), .Z(n122) );
  MUX2_X1 U732 ( .A(n122), .B(n121), .S(n242), .Z(n123) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n247), .Z(n124) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n247), .Z(n125) );
  MUX2_X1 U735 ( .A(n125), .B(n124), .S(n242), .Z(n126) );
  MUX2_X1 U736 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n248), .Z(n128) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n248), .Z(n129) );
  MUX2_X1 U739 ( .A(n129), .B(n128), .S(n242), .Z(n130) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n248), .Z(n131) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n248), .Z(n132) );
  MUX2_X1 U742 ( .A(n132), .B(n131), .S(n242), .Z(n133) );
  MUX2_X1 U743 ( .A(n133), .B(n130), .S(N12), .Z(n134) );
  MUX2_X1 U744 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n248), .Z(n136) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n248), .Z(n137) );
  MUX2_X1 U747 ( .A(n137), .B(n136), .S(n242), .Z(n138) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n248), .Z(n139) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n248), .Z(n140) );
  MUX2_X1 U750 ( .A(n140), .B(n139), .S(n242), .Z(n141) );
  MUX2_X1 U751 ( .A(n141), .B(n138), .S(N12), .Z(n142) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n248), .Z(n143) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n248), .Z(n144) );
  MUX2_X1 U754 ( .A(n144), .B(n143), .S(n242), .Z(n145) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n248), .Z(n146) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n248), .Z(n147) );
  MUX2_X1 U757 ( .A(n147), .B(n146), .S(n242), .Z(n148) );
  MUX2_X1 U758 ( .A(n148), .B(n145), .S(N12), .Z(n149) );
  MUX2_X1 U759 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U760 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n249), .Z(n151) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n249), .Z(n152) );
  MUX2_X1 U763 ( .A(n152), .B(n151), .S(n243), .Z(n153) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n249), .Z(n154) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n249), .Z(n155) );
  MUX2_X1 U766 ( .A(n155), .B(n154), .S(n243), .Z(n156) );
  MUX2_X1 U767 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n249), .Z(n158) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n249), .Z(n159) );
  MUX2_X1 U770 ( .A(n159), .B(n158), .S(n243), .Z(n160) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n249), .Z(n161) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n249), .Z(n162) );
  MUX2_X1 U773 ( .A(n162), .B(n161), .S(n243), .Z(n163) );
  MUX2_X1 U774 ( .A(n163), .B(n160), .S(n241), .Z(n164) );
  MUX2_X1 U775 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n249), .Z(n166) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n249), .Z(n167) );
  MUX2_X1 U778 ( .A(n167), .B(n166), .S(n243), .Z(n168) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n249), .Z(n169) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n249), .Z(n170) );
  MUX2_X1 U781 ( .A(n170), .B(n169), .S(n243), .Z(n171) );
  MUX2_X1 U782 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n247), .Z(n173) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(N10), .Z(n174) );
  MUX2_X1 U785 ( .A(n174), .B(n173), .S(n243), .Z(n175) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n176) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n250), .Z(n177) );
  MUX2_X1 U788 ( .A(n177), .B(n176), .S(n243), .Z(n178) );
  MUX2_X1 U789 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U790 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U791 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n249), .Z(n181) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n250), .Z(n182) );
  MUX2_X1 U794 ( .A(n182), .B(n181), .S(n243), .Z(n183) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n248), .Z(n184) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n245), .Z(n185) );
  MUX2_X1 U797 ( .A(n185), .B(n184), .S(n243), .Z(n186) );
  MUX2_X1 U798 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n250), .Z(n188) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n245), .Z(n189) );
  MUX2_X1 U801 ( .A(n189), .B(n188), .S(n243), .Z(n190) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n246), .Z(n191) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(N10), .Z(n192) );
  MUX2_X1 U804 ( .A(n192), .B(n191), .S(n243), .Z(n193) );
  MUX2_X1 U805 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U806 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n245), .Z(n196) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n250), .Z(n197) );
  MUX2_X1 U809 ( .A(n197), .B(n196), .S(n244), .Z(n198) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n250), .Z(n199) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n200) );
  MUX2_X1 U812 ( .A(n200), .B(n199), .S(n244), .Z(n201) );
  MUX2_X1 U813 ( .A(n201), .B(n198), .S(n241), .Z(n202) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n250), .Z(n203) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n204) );
  MUX2_X1 U816 ( .A(n204), .B(n203), .S(n244), .Z(n205) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n206) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n207) );
  MUX2_X1 U819 ( .A(n207), .B(n206), .S(n244), .Z(n208) );
  MUX2_X1 U820 ( .A(n208), .B(n205), .S(n241), .Z(n209) );
  MUX2_X1 U821 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U822 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n250), .Z(n211) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n246), .Z(n212) );
  MUX2_X1 U825 ( .A(n212), .B(n211), .S(n244), .Z(n213) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n249), .Z(n214) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(N10), .Z(n215) );
  MUX2_X1 U828 ( .A(n215), .B(n214), .S(n244), .Z(n216) );
  MUX2_X1 U829 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n247), .Z(n218) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n250), .Z(n219) );
  MUX2_X1 U832 ( .A(n219), .B(n218), .S(n244), .Z(n220) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n247), .Z(n221) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n222) );
  MUX2_X1 U835 ( .A(n222), .B(n221), .S(n244), .Z(n223) );
  MUX2_X1 U836 ( .A(n223), .B(n220), .S(n241), .Z(n224) );
  MUX2_X1 U837 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n247), .Z(n226) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n250), .Z(n227) );
  MUX2_X1 U840 ( .A(n227), .B(n226), .S(n244), .Z(n228) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n247), .Z(n229) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n230) );
  MUX2_X1 U843 ( .A(n230), .B(n229), .S(n244), .Z(n231) );
  MUX2_X1 U844 ( .A(n231), .B(n228), .S(N12), .Z(n232) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n233) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n234) );
  MUX2_X1 U847 ( .A(n234), .B(n233), .S(n244), .Z(n235) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n236) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n237) );
  MUX2_X1 U850 ( .A(n237), .B(n236), .S(n244), .Z(n238) );
  MUX2_X1 U851 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U852 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U853 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_7 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N22, n1, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n257), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n258), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n259), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n260), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n261), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n262), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n263), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n264), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n265), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n266), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n267), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n268), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n269), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n270), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n271), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n272), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n273), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n274), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n275), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n276), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n277), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n278), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n279), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n280), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n281), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n282), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n283), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n284), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n285), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n286), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n287), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n288), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n289), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n290), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n291), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n292), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n293), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n594), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n595), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n596), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n597), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n598), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n599), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n600), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n601), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n602), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n603), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n604), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n605), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n606), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n607), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n608), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n609), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n610), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n611), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n612), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n613), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n614), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n615), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n616), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n617), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n618), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n619), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n620), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n621), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n622), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n623), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n624), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n625), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n626), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n627), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n628), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n629), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n630), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n631), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n632), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n633), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n634), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n635), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n636), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n637), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n638), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n639), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n640), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n641), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n642), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n643), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n644), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n645), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n646), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n647), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n648), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n649), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n650), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n651), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n652), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n653), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n654), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n655), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n656), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n657), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n658), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n659), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n660), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n661), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n662), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n663), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n664), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n665), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n666), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n667), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n668), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n669), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n670), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n671), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n672), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n673), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n674), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n675), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n676), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n677), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n678), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n679), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n680), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n681), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n682), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n683), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n684), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n685), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n686), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n687), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n688), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n689), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n690), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n691), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n692), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n693), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n694), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n695), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n696), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n697), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n698), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n699), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n700), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n701), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n702), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n703), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n704), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n705), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n706), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n707), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n708), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n709), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n710), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n711), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n712), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n713), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n714), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n715), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n716), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n717), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n718), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n719), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n720), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n721), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n722), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n723), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n724), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n725), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n726), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n727), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n728), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n729), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n730), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n731), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n732), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n733), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n734), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n735), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n736), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n737), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n738), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n739), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n740), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n741), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n742), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n743), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n744), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n745), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n746), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n747), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n748), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n749), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n750), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n751), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n752), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n753), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n754), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n755), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n756), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n757), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n758), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n759), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n760), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n761), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n762), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n763), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n764), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n765), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n766), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n767), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n768), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n769), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n770), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n771), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n772), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n773), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n774), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n775), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n776), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n777), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n778), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n779), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n780), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n781), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n782), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n783), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n784), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n785), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n786), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n787), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n788), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n789), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n790), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n791), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n792), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n793), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n794), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n795), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n796), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n797), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n798), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n799), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n800), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n801), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n802), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n803), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n804), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n805), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n806), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n807), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n808), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n809), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n810), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n811), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n812), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  SDFF_X1 \data_out_reg[1]  ( .D(n63), .SI(n48), .SE(N14), .CK(clk), .Q(
        data_out[1]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(n253), .Z(n251) );
  BUF_X1 U5 ( .A(n253), .Z(n252) );
  BUF_X1 U6 ( .A(n253), .Z(n249) );
  BUF_X1 U7 ( .A(n253), .Z(n250) );
  BUF_X1 U8 ( .A(N10), .Z(n253) );
  INV_X1 U9 ( .A(n1114), .ZN(n844) );
  INV_X1 U10 ( .A(n1103), .ZN(n843) );
  INV_X1 U11 ( .A(n1093), .ZN(n842) );
  INV_X1 U12 ( .A(n1083), .ZN(n841) );
  INV_X1 U13 ( .A(n1073), .ZN(n840) );
  INV_X1 U14 ( .A(n1063), .ZN(n839) );
  INV_X1 U15 ( .A(n1054), .ZN(n838) );
  INV_X1 U16 ( .A(n1045), .ZN(n837) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1106) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n254), .ZN(n1095) );
  NAND2_X1 U19 ( .A1(n1105), .A2(n1137), .ZN(n1063) );
  NAND2_X1 U20 ( .A1(n1106), .A2(n1105), .ZN(n1114) );
  NAND2_X1 U21 ( .A1(n1095), .A2(n1105), .ZN(n1103) );
  NAND2_X1 U22 ( .A1(n1085), .A2(n1105), .ZN(n1093) );
  NAND2_X1 U23 ( .A1(n1075), .A2(n1105), .ZN(n1083) );
  NAND2_X1 U24 ( .A1(n1065), .A2(n1105), .ZN(n1073) );
  NAND2_X1 U25 ( .A1(n1105), .A2(n1126), .ZN(n1054) );
  NAND2_X1 U26 ( .A1(n1105), .A2(n1116), .ZN(n1045) );
  INV_X1 U27 ( .A(n1134), .ZN(n819) );
  INV_X1 U28 ( .A(n1124), .ZN(n818) );
  INV_X1 U29 ( .A(n890), .ZN(n817) );
  INV_X1 U30 ( .A(n881), .ZN(n816) );
  INV_X1 U31 ( .A(n872), .ZN(n815) );
  INV_X1 U32 ( .A(n863), .ZN(n814) );
  INV_X1 U33 ( .A(n854), .ZN(n813) );
  INV_X1 U34 ( .A(n990), .ZN(n831) );
  INV_X1 U35 ( .A(n981), .ZN(n830) );
  INV_X1 U36 ( .A(n972), .ZN(n829) );
  INV_X1 U37 ( .A(n917), .ZN(n823) );
  INV_X1 U38 ( .A(n908), .ZN(n822) );
  INV_X1 U39 ( .A(n899), .ZN(n821) );
  INV_X1 U40 ( .A(n1036), .ZN(n836) );
  INV_X1 U41 ( .A(n1026), .ZN(n835) );
  INV_X1 U42 ( .A(n1017), .ZN(n834) );
  INV_X1 U43 ( .A(n1008), .ZN(n833) );
  INV_X1 U44 ( .A(n999), .ZN(n832) );
  INV_X1 U45 ( .A(n963), .ZN(n828) );
  INV_X1 U46 ( .A(n953), .ZN(n827) );
  INV_X1 U47 ( .A(n944), .ZN(n826) );
  INV_X1 U48 ( .A(n935), .ZN(n825) );
  INV_X1 U49 ( .A(n926), .ZN(n824) );
  INV_X1 U50 ( .A(n1145), .ZN(n820) );
  BUF_X1 U51 ( .A(N11), .Z(n245) );
  BUF_X1 U52 ( .A(N11), .Z(n246) );
  BUF_X1 U53 ( .A(N11), .Z(n247) );
  INV_X1 U54 ( .A(N10), .ZN(n254) );
  BUF_X1 U55 ( .A(N12), .Z(n244) );
  NOR3_X1 U56 ( .A1(n256), .A2(N10), .A3(n255), .ZN(n1126) );
  NOR3_X1 U57 ( .A1(n256), .A2(n254), .A3(n255), .ZN(n1116) );
  NOR3_X1 U58 ( .A1(n254), .A2(N11), .A3(n256), .ZN(n1137) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n255), .ZN(n1085) );
  NOR3_X1 U60 ( .A1(n254), .A2(N12), .A3(n255), .ZN(n1075) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n256), .ZN(n1065) );
  NAND2_X1 U62 ( .A1(n1028), .A2(n1137), .ZN(n990) );
  NAND2_X1 U63 ( .A1(n955), .A2(n1137), .ZN(n917) );
  NAND2_X1 U64 ( .A1(n1028), .A2(n1065), .ZN(n999) );
  NAND2_X1 U65 ( .A1(n955), .A2(n1065), .ZN(n926) );
  NAND2_X1 U66 ( .A1(n1028), .A2(n1106), .ZN(n1036) );
  NAND2_X1 U67 ( .A1(n1028), .A2(n1095), .ZN(n1026) );
  NAND2_X1 U68 ( .A1(n955), .A2(n1106), .ZN(n963) );
  NAND2_X1 U69 ( .A1(n955), .A2(n1095), .ZN(n953) );
  NAND2_X1 U70 ( .A1(n1106), .A2(n1136), .ZN(n890) );
  NAND2_X1 U71 ( .A1(n1095), .A2(n1136), .ZN(n881) );
  NAND2_X1 U72 ( .A1(n1085), .A2(n1136), .ZN(n872) );
  NAND2_X1 U73 ( .A1(n1075), .A2(n1136), .ZN(n863) );
  NAND2_X1 U74 ( .A1(n1065), .A2(n1136), .ZN(n854) );
  NAND2_X1 U75 ( .A1(n1137), .A2(n1136), .ZN(n1145) );
  NAND2_X1 U76 ( .A1(n1126), .A2(n1136), .ZN(n1134) );
  NAND2_X1 U77 ( .A1(n1116), .A2(n1136), .ZN(n1124) );
  NAND2_X1 U78 ( .A1(n1028), .A2(n1085), .ZN(n1017) );
  NAND2_X1 U79 ( .A1(n1028), .A2(n1075), .ZN(n1008) );
  NAND2_X1 U80 ( .A1(n955), .A2(n1085), .ZN(n944) );
  NAND2_X1 U81 ( .A1(n955), .A2(n1075), .ZN(n935) );
  NAND2_X1 U82 ( .A1(n1028), .A2(n1126), .ZN(n981) );
  NAND2_X1 U83 ( .A1(n955), .A2(n1126), .ZN(n908) );
  NAND2_X1 U84 ( .A1(n1028), .A2(n1116), .ZN(n972) );
  NAND2_X1 U85 ( .A1(n955), .A2(n1116), .ZN(n899) );
  AND3_X1 U86 ( .A1(n845), .A2(n846), .A3(wr_en), .ZN(n1105) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1136) );
  AND3_X1 U88 ( .A1(N13), .A2(n846), .A3(wr_en), .ZN(n1028) );
  AND3_X1 U89 ( .A1(N14), .A2(n845), .A3(wr_en), .ZN(n955) );
  INV_X1 U90 ( .A(n1064), .ZN(n772) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n839), .B1(n1063), .B2(\mem[5][0] ), 
        .ZN(n1064) );
  INV_X1 U92 ( .A(n1062), .ZN(n771) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n839), .B1(n1063), .B2(\mem[5][1] ), 
        .ZN(n1062) );
  INV_X1 U94 ( .A(n1061), .ZN(n770) );
  AOI22_X1 U95 ( .A1(data_in[2]), .A2(n839), .B1(n1063), .B2(\mem[5][2] ), 
        .ZN(n1061) );
  INV_X1 U96 ( .A(n1060), .ZN(n769) );
  AOI22_X1 U97 ( .A1(data_in[3]), .A2(n839), .B1(n1063), .B2(\mem[5][3] ), 
        .ZN(n1060) );
  INV_X1 U98 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U99 ( .A1(data_in[4]), .A2(n839), .B1(n1063), .B2(\mem[5][4] ), 
        .ZN(n1059) );
  INV_X1 U100 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U101 ( .A1(data_in[5]), .A2(n839), .B1(n1063), .B2(\mem[5][5] ), 
        .ZN(n1058) );
  INV_X1 U102 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U103 ( .A1(data_in[6]), .A2(n839), .B1(n1063), .B2(\mem[5][6] ), 
        .ZN(n1057) );
  INV_X1 U104 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U105 ( .A1(data_in[7]), .A2(n839), .B1(n1063), .B2(\mem[5][7] ), 
        .ZN(n1056) );
  INV_X1 U106 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U107 ( .A1(data_in[5]), .A2(n835), .B1(n1026), .B2(\mem[9][5] ), 
        .ZN(n1021) );
  INV_X1 U108 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U109 ( .A1(data_in[6]), .A2(n835), .B1(n1026), .B2(\mem[9][6] ), 
        .ZN(n1020) );
  INV_X1 U110 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U111 ( .A1(data_in[7]), .A2(n835), .B1(n1026), .B2(\mem[9][7] ), 
        .ZN(n1019) );
  INV_X1 U112 ( .A(n991), .ZN(n708) );
  AOI22_X1 U113 ( .A1(data_in[0]), .A2(n831), .B1(n990), .B2(\mem[13][0] ), 
        .ZN(n991) );
  INV_X1 U114 ( .A(n989), .ZN(n707) );
  AOI22_X1 U115 ( .A1(data_in[1]), .A2(n831), .B1(n990), .B2(\mem[13][1] ), 
        .ZN(n989) );
  INV_X1 U116 ( .A(n988), .ZN(n706) );
  AOI22_X1 U117 ( .A1(data_in[2]), .A2(n831), .B1(n990), .B2(\mem[13][2] ), 
        .ZN(n988) );
  INV_X1 U118 ( .A(n987), .ZN(n705) );
  AOI22_X1 U119 ( .A1(data_in[3]), .A2(n831), .B1(n990), .B2(\mem[13][3] ), 
        .ZN(n987) );
  INV_X1 U120 ( .A(n986), .ZN(n704) );
  AOI22_X1 U121 ( .A1(data_in[4]), .A2(n831), .B1(n990), .B2(\mem[13][4] ), 
        .ZN(n986) );
  INV_X1 U122 ( .A(n985), .ZN(n703) );
  AOI22_X1 U123 ( .A1(data_in[5]), .A2(n831), .B1(n990), .B2(\mem[13][5] ), 
        .ZN(n985) );
  INV_X1 U124 ( .A(n984), .ZN(n702) );
  AOI22_X1 U125 ( .A1(data_in[6]), .A2(n831), .B1(n990), .B2(\mem[13][6] ), 
        .ZN(n984) );
  INV_X1 U126 ( .A(n983), .ZN(n701) );
  AOI22_X1 U127 ( .A1(data_in[7]), .A2(n831), .B1(n990), .B2(\mem[13][7] ), 
        .ZN(n983) );
  INV_X1 U128 ( .A(n954), .ZN(n676) );
  AOI22_X1 U129 ( .A1(data_in[0]), .A2(n827), .B1(n953), .B2(\mem[17][0] ), 
        .ZN(n954) );
  INV_X1 U130 ( .A(n952), .ZN(n675) );
  AOI22_X1 U131 ( .A1(data_in[1]), .A2(n827), .B1(n953), .B2(\mem[17][1] ), 
        .ZN(n952) );
  INV_X1 U132 ( .A(n951), .ZN(n674) );
  AOI22_X1 U133 ( .A1(data_in[2]), .A2(n827), .B1(n953), .B2(\mem[17][2] ), 
        .ZN(n951) );
  INV_X1 U134 ( .A(n950), .ZN(n673) );
  AOI22_X1 U135 ( .A1(data_in[3]), .A2(n827), .B1(n953), .B2(\mem[17][3] ), 
        .ZN(n950) );
  INV_X1 U136 ( .A(n949), .ZN(n672) );
  AOI22_X1 U137 ( .A1(data_in[4]), .A2(n827), .B1(n953), .B2(\mem[17][4] ), 
        .ZN(n949) );
  INV_X1 U138 ( .A(n948), .ZN(n671) );
  AOI22_X1 U139 ( .A1(data_in[5]), .A2(n827), .B1(n953), .B2(\mem[17][5] ), 
        .ZN(n948) );
  INV_X1 U140 ( .A(n947), .ZN(n670) );
  AOI22_X1 U141 ( .A1(data_in[6]), .A2(n827), .B1(n953), .B2(\mem[17][6] ), 
        .ZN(n947) );
  INV_X1 U142 ( .A(n918), .ZN(n644) );
  AOI22_X1 U143 ( .A1(data_in[0]), .A2(n823), .B1(n917), .B2(\mem[21][0] ), 
        .ZN(n918) );
  INV_X1 U144 ( .A(n916), .ZN(n643) );
  AOI22_X1 U145 ( .A1(data_in[1]), .A2(n823), .B1(n917), .B2(\mem[21][1] ), 
        .ZN(n916) );
  INV_X1 U146 ( .A(n915), .ZN(n642) );
  AOI22_X1 U147 ( .A1(data_in[2]), .A2(n823), .B1(n917), .B2(\mem[21][2] ), 
        .ZN(n915) );
  INV_X1 U148 ( .A(n914), .ZN(n641) );
  AOI22_X1 U149 ( .A1(data_in[3]), .A2(n823), .B1(n917), .B2(\mem[21][3] ), 
        .ZN(n914) );
  INV_X1 U150 ( .A(n913), .ZN(n640) );
  AOI22_X1 U151 ( .A1(data_in[4]), .A2(n823), .B1(n917), .B2(\mem[21][4] ), 
        .ZN(n913) );
  INV_X1 U152 ( .A(n912), .ZN(n639) );
  AOI22_X1 U153 ( .A1(data_in[5]), .A2(n823), .B1(n917), .B2(\mem[21][5] ), 
        .ZN(n912) );
  INV_X1 U154 ( .A(n911), .ZN(n638) );
  AOI22_X1 U155 ( .A1(data_in[6]), .A2(n823), .B1(n917), .B2(\mem[21][6] ), 
        .ZN(n911) );
  INV_X1 U156 ( .A(n910), .ZN(n637) );
  AOI22_X1 U157 ( .A1(data_in[7]), .A2(n823), .B1(n917), .B2(\mem[21][7] ), 
        .ZN(n910) );
  INV_X1 U158 ( .A(n1027), .ZN(n740) );
  AOI22_X1 U159 ( .A1(data_in[0]), .A2(n835), .B1(n1026), .B2(\mem[9][0] ), 
        .ZN(n1027) );
  INV_X1 U160 ( .A(n1025), .ZN(n739) );
  AOI22_X1 U161 ( .A1(data_in[1]), .A2(n835), .B1(n1026), .B2(\mem[9][1] ), 
        .ZN(n1025) );
  INV_X1 U162 ( .A(n1024), .ZN(n738) );
  AOI22_X1 U163 ( .A1(data_in[2]), .A2(n835), .B1(n1026), .B2(\mem[9][2] ), 
        .ZN(n1024) );
  INV_X1 U164 ( .A(n1023), .ZN(n737) );
  AOI22_X1 U165 ( .A1(data_in[3]), .A2(n835), .B1(n1026), .B2(\mem[9][3] ), 
        .ZN(n1023) );
  INV_X1 U166 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U167 ( .A1(data_in[4]), .A2(n835), .B1(n1026), .B2(\mem[9][4] ), 
        .ZN(n1022) );
  INV_X1 U168 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U169 ( .A1(data_in[0]), .A2(n838), .B1(n1054), .B2(\mem[6][0] ), 
        .ZN(n1055) );
  INV_X1 U170 ( .A(n1053), .ZN(n763) );
  AOI22_X1 U171 ( .A1(data_in[1]), .A2(n838), .B1(n1054), .B2(\mem[6][1] ), 
        .ZN(n1053) );
  INV_X1 U172 ( .A(n1052), .ZN(n762) );
  AOI22_X1 U173 ( .A1(data_in[2]), .A2(n838), .B1(n1054), .B2(\mem[6][2] ), 
        .ZN(n1052) );
  INV_X1 U174 ( .A(n1051), .ZN(n761) );
  AOI22_X1 U175 ( .A1(data_in[3]), .A2(n838), .B1(n1054), .B2(\mem[6][3] ), 
        .ZN(n1051) );
  INV_X1 U176 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U177 ( .A1(data_in[4]), .A2(n838), .B1(n1054), .B2(\mem[6][4] ), 
        .ZN(n1050) );
  INV_X1 U178 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U179 ( .A1(data_in[5]), .A2(n838), .B1(n1054), .B2(\mem[6][5] ), 
        .ZN(n1049) );
  INV_X1 U180 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U181 ( .A1(data_in[6]), .A2(n838), .B1(n1054), .B2(\mem[6][6] ), 
        .ZN(n1048) );
  INV_X1 U182 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U183 ( .A1(data_in[7]), .A2(n838), .B1(n1054), .B2(\mem[6][7] ), 
        .ZN(n1047) );
  INV_X1 U184 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U185 ( .A1(data_in[0]), .A2(n837), .B1(n1045), .B2(\mem[7][0] ), 
        .ZN(n1046) );
  INV_X1 U186 ( .A(n1044), .ZN(n755) );
  AOI22_X1 U187 ( .A1(data_in[1]), .A2(n837), .B1(n1045), .B2(\mem[7][1] ), 
        .ZN(n1044) );
  INV_X1 U188 ( .A(n1043), .ZN(n754) );
  AOI22_X1 U189 ( .A1(data_in[2]), .A2(n837), .B1(n1045), .B2(\mem[7][2] ), 
        .ZN(n1043) );
  INV_X1 U190 ( .A(n1042), .ZN(n753) );
  AOI22_X1 U191 ( .A1(data_in[3]), .A2(n837), .B1(n1045), .B2(\mem[7][3] ), 
        .ZN(n1042) );
  INV_X1 U192 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U193 ( .A1(data_in[4]), .A2(n837), .B1(n1045), .B2(\mem[7][4] ), 
        .ZN(n1041) );
  INV_X1 U194 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U195 ( .A1(data_in[5]), .A2(n837), .B1(n1045), .B2(\mem[7][5] ), 
        .ZN(n1040) );
  INV_X1 U196 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U197 ( .A1(data_in[6]), .A2(n837), .B1(n1045), .B2(\mem[7][6] ), 
        .ZN(n1039) );
  INV_X1 U198 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U199 ( .A1(data_in[7]), .A2(n837), .B1(n1045), .B2(\mem[7][7] ), 
        .ZN(n1038) );
  INV_X1 U200 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U201 ( .A1(data_in[0]), .A2(n834), .B1(n1017), .B2(\mem[10][0] ), 
        .ZN(n1018) );
  INV_X1 U202 ( .A(n1016), .ZN(n731) );
  AOI22_X1 U203 ( .A1(data_in[1]), .A2(n834), .B1(n1017), .B2(\mem[10][1] ), 
        .ZN(n1016) );
  INV_X1 U204 ( .A(n1015), .ZN(n730) );
  AOI22_X1 U205 ( .A1(data_in[2]), .A2(n834), .B1(n1017), .B2(\mem[10][2] ), 
        .ZN(n1015) );
  INV_X1 U206 ( .A(n1014), .ZN(n729) );
  AOI22_X1 U207 ( .A1(data_in[3]), .A2(n834), .B1(n1017), .B2(\mem[10][3] ), 
        .ZN(n1014) );
  INV_X1 U208 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U209 ( .A1(data_in[4]), .A2(n834), .B1(n1017), .B2(\mem[10][4] ), 
        .ZN(n1013) );
  INV_X1 U210 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U211 ( .A1(data_in[5]), .A2(n834), .B1(n1017), .B2(\mem[10][5] ), 
        .ZN(n1012) );
  INV_X1 U212 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U213 ( .A1(data_in[6]), .A2(n834), .B1(n1017), .B2(\mem[10][6] ), 
        .ZN(n1011) );
  INV_X1 U214 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U215 ( .A1(data_in[7]), .A2(n834), .B1(n1017), .B2(\mem[10][7] ), 
        .ZN(n1010) );
  INV_X1 U216 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U217 ( .A1(data_in[0]), .A2(n833), .B1(n1008), .B2(\mem[11][0] ), 
        .ZN(n1009) );
  INV_X1 U218 ( .A(n1007), .ZN(n723) );
  AOI22_X1 U219 ( .A1(data_in[1]), .A2(n833), .B1(n1008), .B2(\mem[11][1] ), 
        .ZN(n1007) );
  INV_X1 U220 ( .A(n1006), .ZN(n722) );
  AOI22_X1 U221 ( .A1(data_in[2]), .A2(n833), .B1(n1008), .B2(\mem[11][2] ), 
        .ZN(n1006) );
  INV_X1 U222 ( .A(n1005), .ZN(n721) );
  AOI22_X1 U223 ( .A1(data_in[3]), .A2(n833), .B1(n1008), .B2(\mem[11][3] ), 
        .ZN(n1005) );
  INV_X1 U224 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U225 ( .A1(data_in[4]), .A2(n833), .B1(n1008), .B2(\mem[11][4] ), 
        .ZN(n1004) );
  INV_X1 U226 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U227 ( .A1(data_in[5]), .A2(n833), .B1(n1008), .B2(\mem[11][5] ), 
        .ZN(n1003) );
  INV_X1 U228 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U229 ( .A1(data_in[6]), .A2(n833), .B1(n1008), .B2(\mem[11][6] ), 
        .ZN(n1002) );
  INV_X1 U230 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U231 ( .A1(data_in[7]), .A2(n833), .B1(n1008), .B2(\mem[11][7] ), 
        .ZN(n1001) );
  INV_X1 U232 ( .A(n946), .ZN(n669) );
  AOI22_X1 U233 ( .A1(data_in[7]), .A2(n827), .B1(n953), .B2(\mem[17][7] ), 
        .ZN(n946) );
  INV_X1 U234 ( .A(n938), .ZN(n662) );
  AOI22_X1 U235 ( .A1(data_in[6]), .A2(n826), .B1(n944), .B2(\mem[18][6] ), 
        .ZN(n938) );
  INV_X1 U236 ( .A(n937), .ZN(n661) );
  AOI22_X1 U237 ( .A1(data_in[7]), .A2(n826), .B1(n944), .B2(\mem[18][7] ), 
        .ZN(n937) );
  INV_X1 U238 ( .A(n936), .ZN(n660) );
  AOI22_X1 U239 ( .A1(data_in[0]), .A2(n825), .B1(n935), .B2(\mem[19][0] ), 
        .ZN(n936) );
  INV_X1 U240 ( .A(n934), .ZN(n659) );
  AOI22_X1 U241 ( .A1(data_in[1]), .A2(n825), .B1(n935), .B2(\mem[19][1] ), 
        .ZN(n934) );
  INV_X1 U242 ( .A(n933), .ZN(n658) );
  AOI22_X1 U243 ( .A1(data_in[2]), .A2(n825), .B1(n935), .B2(\mem[19][2] ), 
        .ZN(n933) );
  INV_X1 U244 ( .A(n932), .ZN(n657) );
  AOI22_X1 U245 ( .A1(data_in[3]), .A2(n825), .B1(n935), .B2(\mem[19][3] ), 
        .ZN(n932) );
  INV_X1 U246 ( .A(n931), .ZN(n656) );
  AOI22_X1 U247 ( .A1(data_in[4]), .A2(n825), .B1(n935), .B2(\mem[19][4] ), 
        .ZN(n931) );
  INV_X1 U248 ( .A(n930), .ZN(n655) );
  AOI22_X1 U249 ( .A1(data_in[5]), .A2(n825), .B1(n935), .B2(\mem[19][5] ), 
        .ZN(n930) );
  INV_X1 U250 ( .A(n929), .ZN(n654) );
  AOI22_X1 U251 ( .A1(data_in[6]), .A2(n825), .B1(n935), .B2(\mem[19][6] ), 
        .ZN(n929) );
  INV_X1 U252 ( .A(n928), .ZN(n653) );
  AOI22_X1 U253 ( .A1(data_in[7]), .A2(n825), .B1(n935), .B2(\mem[19][7] ), 
        .ZN(n928) );
  INV_X1 U254 ( .A(n982), .ZN(n700) );
  AOI22_X1 U255 ( .A1(data_in[0]), .A2(n830), .B1(n981), .B2(\mem[14][0] ), 
        .ZN(n982) );
  INV_X1 U256 ( .A(n980), .ZN(n699) );
  AOI22_X1 U257 ( .A1(data_in[1]), .A2(n830), .B1(n981), .B2(\mem[14][1] ), 
        .ZN(n980) );
  INV_X1 U258 ( .A(n979), .ZN(n698) );
  AOI22_X1 U259 ( .A1(data_in[2]), .A2(n830), .B1(n981), .B2(\mem[14][2] ), 
        .ZN(n979) );
  INV_X1 U260 ( .A(n978), .ZN(n697) );
  AOI22_X1 U261 ( .A1(data_in[3]), .A2(n830), .B1(n981), .B2(\mem[14][3] ), 
        .ZN(n978) );
  INV_X1 U262 ( .A(n977), .ZN(n696) );
  AOI22_X1 U263 ( .A1(data_in[4]), .A2(n830), .B1(n981), .B2(\mem[14][4] ), 
        .ZN(n977) );
  INV_X1 U264 ( .A(n976), .ZN(n695) );
  AOI22_X1 U265 ( .A1(data_in[5]), .A2(n830), .B1(n981), .B2(\mem[14][5] ), 
        .ZN(n976) );
  INV_X1 U266 ( .A(n975), .ZN(n694) );
  AOI22_X1 U267 ( .A1(data_in[6]), .A2(n830), .B1(n981), .B2(\mem[14][6] ), 
        .ZN(n975) );
  INV_X1 U268 ( .A(n974), .ZN(n693) );
  AOI22_X1 U269 ( .A1(data_in[7]), .A2(n830), .B1(n981), .B2(\mem[14][7] ), 
        .ZN(n974) );
  INV_X1 U270 ( .A(n973), .ZN(n692) );
  AOI22_X1 U271 ( .A1(data_in[0]), .A2(n829), .B1(n972), .B2(\mem[15][0] ), 
        .ZN(n973) );
  INV_X1 U272 ( .A(n971), .ZN(n691) );
  AOI22_X1 U273 ( .A1(data_in[1]), .A2(n829), .B1(n972), .B2(\mem[15][1] ), 
        .ZN(n971) );
  INV_X1 U274 ( .A(n970), .ZN(n690) );
  AOI22_X1 U275 ( .A1(data_in[2]), .A2(n829), .B1(n972), .B2(\mem[15][2] ), 
        .ZN(n970) );
  INV_X1 U276 ( .A(n969), .ZN(n689) );
  AOI22_X1 U277 ( .A1(data_in[3]), .A2(n829), .B1(n972), .B2(\mem[15][3] ), 
        .ZN(n969) );
  INV_X1 U278 ( .A(n968), .ZN(n688) );
  AOI22_X1 U279 ( .A1(data_in[4]), .A2(n829), .B1(n972), .B2(\mem[15][4] ), 
        .ZN(n968) );
  INV_X1 U280 ( .A(n967), .ZN(n687) );
  AOI22_X1 U281 ( .A1(data_in[5]), .A2(n829), .B1(n972), .B2(\mem[15][5] ), 
        .ZN(n967) );
  INV_X1 U282 ( .A(n966), .ZN(n686) );
  AOI22_X1 U283 ( .A1(data_in[6]), .A2(n829), .B1(n972), .B2(\mem[15][6] ), 
        .ZN(n966) );
  INV_X1 U284 ( .A(n965), .ZN(n685) );
  AOI22_X1 U285 ( .A1(data_in[7]), .A2(n829), .B1(n972), .B2(\mem[15][7] ), 
        .ZN(n965) );
  INV_X1 U286 ( .A(n945), .ZN(n668) );
  AOI22_X1 U287 ( .A1(data_in[0]), .A2(n826), .B1(n944), .B2(\mem[18][0] ), 
        .ZN(n945) );
  INV_X1 U288 ( .A(n943), .ZN(n667) );
  AOI22_X1 U289 ( .A1(data_in[1]), .A2(n826), .B1(n944), .B2(\mem[18][1] ), 
        .ZN(n943) );
  INV_X1 U290 ( .A(n942), .ZN(n666) );
  AOI22_X1 U291 ( .A1(data_in[2]), .A2(n826), .B1(n944), .B2(\mem[18][2] ), 
        .ZN(n942) );
  INV_X1 U292 ( .A(n941), .ZN(n665) );
  AOI22_X1 U293 ( .A1(data_in[3]), .A2(n826), .B1(n944), .B2(\mem[18][3] ), 
        .ZN(n941) );
  INV_X1 U294 ( .A(n940), .ZN(n664) );
  AOI22_X1 U295 ( .A1(data_in[4]), .A2(n826), .B1(n944), .B2(\mem[18][4] ), 
        .ZN(n940) );
  INV_X1 U296 ( .A(n939), .ZN(n663) );
  AOI22_X1 U297 ( .A1(data_in[5]), .A2(n826), .B1(n944), .B2(\mem[18][5] ), 
        .ZN(n939) );
  INV_X1 U298 ( .A(n909), .ZN(n636) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n822), .B1(n908), .B2(\mem[22][0] ), 
        .ZN(n909) );
  INV_X1 U300 ( .A(n907), .ZN(n635) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n822), .B1(n908), .B2(\mem[22][1] ), 
        .ZN(n907) );
  INV_X1 U302 ( .A(n906), .ZN(n634) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n822), .B1(n908), .B2(\mem[22][2] ), 
        .ZN(n906) );
  INV_X1 U304 ( .A(n905), .ZN(n633) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n822), .B1(n908), .B2(\mem[22][3] ), 
        .ZN(n905) );
  INV_X1 U306 ( .A(n904), .ZN(n632) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n822), .B1(n908), .B2(\mem[22][4] ), 
        .ZN(n904) );
  INV_X1 U308 ( .A(n903), .ZN(n631) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n822), .B1(n908), .B2(\mem[22][5] ), 
        .ZN(n903) );
  INV_X1 U310 ( .A(n902), .ZN(n630) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n822), .B1(n908), .B2(\mem[22][6] ), 
        .ZN(n902) );
  INV_X1 U312 ( .A(n901), .ZN(n629) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n822), .B1(n908), .B2(\mem[22][7] ), 
        .ZN(n901) );
  INV_X1 U314 ( .A(n900), .ZN(n628) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n821), .B1(n899), .B2(\mem[23][0] ), 
        .ZN(n900) );
  INV_X1 U316 ( .A(n898), .ZN(n627) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n821), .B1(n899), .B2(\mem[23][1] ), 
        .ZN(n898) );
  INV_X1 U318 ( .A(n897), .ZN(n626) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n821), .B1(n899), .B2(\mem[23][2] ), 
        .ZN(n897) );
  INV_X1 U320 ( .A(n896), .ZN(n625) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n821), .B1(n899), .B2(\mem[23][3] ), 
        .ZN(n896) );
  INV_X1 U322 ( .A(n895), .ZN(n624) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n821), .B1(n899), .B2(\mem[23][4] ), 
        .ZN(n895) );
  INV_X1 U324 ( .A(n894), .ZN(n623) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n821), .B1(n899), .B2(\mem[23][5] ), 
        .ZN(n894) );
  INV_X1 U326 ( .A(n893), .ZN(n622) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n821), .B1(n899), .B2(\mem[23][6] ), 
        .ZN(n893) );
  INV_X1 U328 ( .A(n892), .ZN(n621) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n821), .B1(n899), .B2(\mem[23][7] ), 
        .ZN(n892) );
  INV_X1 U330 ( .A(N12), .ZN(n256) );
  INV_X1 U331 ( .A(N11), .ZN(n255) );
  INV_X1 U332 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n832), .B1(n999), .B2(\mem[12][0] ), 
        .ZN(n1000) );
  INV_X1 U334 ( .A(n998), .ZN(n715) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n832), .B1(n999), .B2(\mem[12][1] ), 
        .ZN(n998) );
  INV_X1 U336 ( .A(n997), .ZN(n714) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n832), .B1(n999), .B2(\mem[12][2] ), 
        .ZN(n997) );
  INV_X1 U338 ( .A(n996), .ZN(n713) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n832), .B1(n999), .B2(\mem[12][3] ), 
        .ZN(n996) );
  INV_X1 U340 ( .A(n995), .ZN(n712) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n832), .B1(n999), .B2(\mem[12][4] ), 
        .ZN(n995) );
  INV_X1 U342 ( .A(n994), .ZN(n711) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n832), .B1(n999), .B2(\mem[12][5] ), 
        .ZN(n994) );
  INV_X1 U344 ( .A(n993), .ZN(n710) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n832), .B1(n999), .B2(\mem[12][6] ), 
        .ZN(n993) );
  INV_X1 U346 ( .A(n992), .ZN(n709) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n832), .B1(n999), .B2(\mem[12][7] ), 
        .ZN(n992) );
  INV_X1 U348 ( .A(n927), .ZN(n652) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n824), .B1(n926), .B2(\mem[20][0] ), 
        .ZN(n927) );
  INV_X1 U350 ( .A(n925), .ZN(n651) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n824), .B1(n926), .B2(\mem[20][1] ), 
        .ZN(n925) );
  INV_X1 U352 ( .A(n924), .ZN(n650) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n824), .B1(n926), .B2(\mem[20][2] ), 
        .ZN(n924) );
  INV_X1 U354 ( .A(n923), .ZN(n649) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n824), .B1(n926), .B2(\mem[20][3] ), 
        .ZN(n923) );
  INV_X1 U356 ( .A(n922), .ZN(n648) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n824), .B1(n926), .B2(\mem[20][4] ), 
        .ZN(n922) );
  INV_X1 U358 ( .A(n921), .ZN(n647) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n824), .B1(n926), .B2(\mem[20][5] ), 
        .ZN(n921) );
  INV_X1 U360 ( .A(n920), .ZN(n646) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n824), .B1(n926), .B2(\mem[20][6] ), 
        .ZN(n920) );
  INV_X1 U362 ( .A(n919), .ZN(n645) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n824), .B1(n926), .B2(\mem[20][7] ), 
        .ZN(n919) );
  INV_X1 U364 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n836), .B1(n1036), .B2(\mem[8][0] ), 
        .ZN(n1037) );
  INV_X1 U366 ( .A(n1035), .ZN(n747) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n836), .B1(n1036), .B2(\mem[8][1] ), 
        .ZN(n1035) );
  INV_X1 U368 ( .A(n1034), .ZN(n746) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n836), .B1(n1036), .B2(\mem[8][2] ), 
        .ZN(n1034) );
  INV_X1 U370 ( .A(n1033), .ZN(n745) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n836), .B1(n1036), .B2(\mem[8][3] ), 
        .ZN(n1033) );
  INV_X1 U372 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n836), .B1(n1036), .B2(\mem[8][4] ), 
        .ZN(n1032) );
  INV_X1 U374 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n836), .B1(n1036), .B2(\mem[8][5] ), 
        .ZN(n1031) );
  INV_X1 U376 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n836), .B1(n1036), .B2(\mem[8][6] ), 
        .ZN(n1030) );
  INV_X1 U378 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n836), .B1(n1036), .B2(\mem[8][7] ), 
        .ZN(n1029) );
  INV_X1 U380 ( .A(n964), .ZN(n684) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n828), .B1(n963), .B2(\mem[16][0] ), 
        .ZN(n964) );
  INV_X1 U382 ( .A(n962), .ZN(n683) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n828), .B1(n963), .B2(\mem[16][1] ), 
        .ZN(n962) );
  INV_X1 U384 ( .A(n961), .ZN(n682) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n828), .B1(n963), .B2(\mem[16][2] ), 
        .ZN(n961) );
  INV_X1 U386 ( .A(n960), .ZN(n681) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n828), .B1(n963), .B2(\mem[16][3] ), 
        .ZN(n960) );
  INV_X1 U388 ( .A(n959), .ZN(n680) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n828), .B1(n963), .B2(\mem[16][4] ), 
        .ZN(n959) );
  INV_X1 U390 ( .A(n958), .ZN(n679) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n828), .B1(n963), .B2(\mem[16][5] ), 
        .ZN(n958) );
  INV_X1 U392 ( .A(n957), .ZN(n678) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n828), .B1(n963), .B2(\mem[16][6] ), 
        .ZN(n957) );
  INV_X1 U394 ( .A(n956), .ZN(n677) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n828), .B1(n963), .B2(\mem[16][7] ), 
        .ZN(n956) );
  INV_X1 U396 ( .A(n891), .ZN(n620) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n817), .B1(n890), .B2(\mem[24][0] ), 
        .ZN(n891) );
  INV_X1 U398 ( .A(n889), .ZN(n619) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n817), .B1(n890), .B2(\mem[24][1] ), 
        .ZN(n889) );
  INV_X1 U400 ( .A(n888), .ZN(n618) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n817), .B1(n890), .B2(\mem[24][2] ), 
        .ZN(n888) );
  INV_X1 U402 ( .A(n887), .ZN(n617) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n817), .B1(n890), .B2(\mem[24][3] ), 
        .ZN(n887) );
  INV_X1 U404 ( .A(n886), .ZN(n616) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n817), .B1(n890), .B2(\mem[24][4] ), 
        .ZN(n886) );
  INV_X1 U406 ( .A(n885), .ZN(n615) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n817), .B1(n890), .B2(\mem[24][5] ), 
        .ZN(n885) );
  INV_X1 U408 ( .A(n884), .ZN(n614) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n817), .B1(n890), .B2(\mem[24][6] ), 
        .ZN(n884) );
  INV_X1 U410 ( .A(n883), .ZN(n613) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n817), .B1(n890), .B2(\mem[24][7] ), 
        .ZN(n883) );
  INV_X1 U412 ( .A(n882), .ZN(n612) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n816), .B1(n881), .B2(\mem[25][0] ), 
        .ZN(n882) );
  INV_X1 U414 ( .A(n880), .ZN(n611) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n816), .B1(n881), .B2(\mem[25][1] ), 
        .ZN(n880) );
  INV_X1 U416 ( .A(n879), .ZN(n610) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n816), .B1(n881), .B2(\mem[25][2] ), 
        .ZN(n879) );
  INV_X1 U418 ( .A(n878), .ZN(n609) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n816), .B1(n881), .B2(\mem[25][3] ), 
        .ZN(n878) );
  INV_X1 U420 ( .A(n877), .ZN(n608) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n816), .B1(n881), .B2(\mem[25][4] ), 
        .ZN(n877) );
  INV_X1 U422 ( .A(n876), .ZN(n607) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n816), .B1(n881), .B2(\mem[25][5] ), 
        .ZN(n876) );
  INV_X1 U424 ( .A(n875), .ZN(n606) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n816), .B1(n881), .B2(\mem[25][6] ), 
        .ZN(n875) );
  INV_X1 U426 ( .A(n874), .ZN(n605) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n816), .B1(n881), .B2(\mem[25][7] ), 
        .ZN(n874) );
  INV_X1 U428 ( .A(n873), .ZN(n604) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n815), .B1(n872), .B2(\mem[26][0] ), 
        .ZN(n873) );
  INV_X1 U430 ( .A(n871), .ZN(n603) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n815), .B1(n872), .B2(\mem[26][1] ), 
        .ZN(n871) );
  INV_X1 U432 ( .A(n870), .ZN(n602) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n815), .B1(n872), .B2(\mem[26][2] ), 
        .ZN(n870) );
  INV_X1 U434 ( .A(n869), .ZN(n601) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n815), .B1(n872), .B2(\mem[26][3] ), 
        .ZN(n869) );
  INV_X1 U436 ( .A(n868), .ZN(n600) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n815), .B1(n872), .B2(\mem[26][4] ), 
        .ZN(n868) );
  INV_X1 U438 ( .A(n867), .ZN(n599) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n815), .B1(n872), .B2(\mem[26][5] ), 
        .ZN(n867) );
  INV_X1 U440 ( .A(n866), .ZN(n598) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n815), .B1(n872), .B2(\mem[26][6] ), 
        .ZN(n866) );
  INV_X1 U442 ( .A(n865), .ZN(n597) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n815), .B1(n872), .B2(\mem[26][7] ), 
        .ZN(n865) );
  INV_X1 U444 ( .A(n864), .ZN(n596) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n814), .B1(n863), .B2(\mem[27][0] ), 
        .ZN(n864) );
  INV_X1 U446 ( .A(n862), .ZN(n595) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n814), .B1(n863), .B2(\mem[27][1] ), 
        .ZN(n862) );
  INV_X1 U448 ( .A(n861), .ZN(n594) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n814), .B1(n863), .B2(\mem[27][2] ), 
        .ZN(n861) );
  INV_X1 U450 ( .A(n860), .ZN(n293) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n814), .B1(n863), .B2(\mem[27][3] ), 
        .ZN(n860) );
  INV_X1 U452 ( .A(n859), .ZN(n292) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n814), .B1(n863), .B2(\mem[27][4] ), 
        .ZN(n859) );
  INV_X1 U454 ( .A(n858), .ZN(n291) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n814), .B1(n863), .B2(\mem[27][5] ), 
        .ZN(n858) );
  INV_X1 U456 ( .A(n857), .ZN(n290) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n814), .B1(n863), .B2(\mem[27][6] ), 
        .ZN(n857) );
  INV_X1 U458 ( .A(n856), .ZN(n289) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n814), .B1(n863), .B2(\mem[27][7] ), 
        .ZN(n856) );
  INV_X1 U460 ( .A(n855), .ZN(n288) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n813), .B1(n854), .B2(\mem[28][0] ), 
        .ZN(n855) );
  INV_X1 U462 ( .A(n853), .ZN(n287) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n813), .B1(n854), .B2(\mem[28][1] ), 
        .ZN(n853) );
  INV_X1 U464 ( .A(n852), .ZN(n286) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n813), .B1(n854), .B2(\mem[28][2] ), 
        .ZN(n852) );
  INV_X1 U466 ( .A(n851), .ZN(n285) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n813), .B1(n854), .B2(\mem[28][3] ), 
        .ZN(n851) );
  INV_X1 U468 ( .A(n850), .ZN(n284) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n813), .B1(n854), .B2(\mem[28][4] ), 
        .ZN(n850) );
  INV_X1 U470 ( .A(n849), .ZN(n283) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n813), .B1(n854), .B2(\mem[28][5] ), 
        .ZN(n849) );
  INV_X1 U472 ( .A(n848), .ZN(n282) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n813), .B1(n854), .B2(\mem[28][6] ), 
        .ZN(n848) );
  INV_X1 U474 ( .A(n847), .ZN(n281) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n813), .B1(n854), .B2(\mem[28][7] ), 
        .ZN(n847) );
  INV_X1 U476 ( .A(n1146), .ZN(n280) );
  AOI22_X1 U477 ( .A1(n820), .A2(data_in[0]), .B1(n1145), .B2(\mem[29][0] ), 
        .ZN(n1146) );
  INV_X1 U478 ( .A(n1144), .ZN(n279) );
  AOI22_X1 U479 ( .A1(n820), .A2(data_in[1]), .B1(n1145), .B2(\mem[29][1] ), 
        .ZN(n1144) );
  INV_X1 U480 ( .A(n1143), .ZN(n278) );
  AOI22_X1 U481 ( .A1(n820), .A2(data_in[2]), .B1(n1145), .B2(\mem[29][2] ), 
        .ZN(n1143) );
  INV_X1 U482 ( .A(n1142), .ZN(n277) );
  AOI22_X1 U483 ( .A1(n820), .A2(data_in[3]), .B1(n1145), .B2(\mem[29][3] ), 
        .ZN(n1142) );
  INV_X1 U484 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U485 ( .A1(n820), .A2(data_in[4]), .B1(n1145), .B2(\mem[29][4] ), 
        .ZN(n1141) );
  INV_X1 U486 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U487 ( .A1(n820), .A2(data_in[5]), .B1(n1145), .B2(\mem[29][5] ), 
        .ZN(n1140) );
  INV_X1 U488 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U489 ( .A1(n820), .A2(data_in[6]), .B1(n1145), .B2(\mem[29][6] ), 
        .ZN(n1139) );
  INV_X1 U490 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U491 ( .A1(n820), .A2(data_in[7]), .B1(n1145), .B2(\mem[29][7] ), 
        .ZN(n1138) );
  INV_X1 U492 ( .A(n1135), .ZN(n272) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n819), .B1(n1134), .B2(\mem[30][0] ), 
        .ZN(n1135) );
  INV_X1 U494 ( .A(n1133), .ZN(n271) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n819), .B1(n1134), .B2(\mem[30][1] ), 
        .ZN(n1133) );
  INV_X1 U496 ( .A(n1132), .ZN(n270) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n819), .B1(n1134), .B2(\mem[30][2] ), 
        .ZN(n1132) );
  INV_X1 U498 ( .A(n1131), .ZN(n269) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n819), .B1(n1134), .B2(\mem[30][3] ), 
        .ZN(n1131) );
  INV_X1 U500 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n819), .B1(n1134), .B2(\mem[30][4] ), 
        .ZN(n1130) );
  INV_X1 U502 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n819), .B1(n1134), .B2(\mem[30][5] ), 
        .ZN(n1129) );
  INV_X1 U504 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n819), .B1(n1134), .B2(\mem[30][6] ), 
        .ZN(n1128) );
  INV_X1 U506 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n819), .B1(n1134), .B2(\mem[30][7] ), 
        .ZN(n1127) );
  INV_X1 U508 ( .A(n1125), .ZN(n264) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n818), .B1(n1124), .B2(\mem[31][0] ), 
        .ZN(n1125) );
  INV_X1 U510 ( .A(n1123), .ZN(n263) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n818), .B1(n1124), .B2(\mem[31][1] ), 
        .ZN(n1123) );
  INV_X1 U512 ( .A(n1122), .ZN(n262) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n818), .B1(n1124), .B2(\mem[31][2] ), 
        .ZN(n1122) );
  INV_X1 U514 ( .A(n1121), .ZN(n261) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n818), .B1(n1124), .B2(\mem[31][3] ), 
        .ZN(n1121) );
  INV_X1 U516 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n818), .B1(n1124), .B2(\mem[31][4] ), 
        .ZN(n1120) );
  INV_X1 U518 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n818), .B1(n1124), .B2(\mem[31][5] ), 
        .ZN(n1119) );
  INV_X1 U520 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n818), .B1(n1124), .B2(\mem[31][6] ), 
        .ZN(n1118) );
  INV_X1 U522 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n818), .B1(n1124), .B2(\mem[31][7] ), 
        .ZN(n1117) );
  INV_X1 U524 ( .A(n1115), .ZN(n812) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n844), .B1(n1114), .B2(\mem[0][0] ), 
        .ZN(n1115) );
  INV_X1 U526 ( .A(n1113), .ZN(n811) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n844), .B1(n1114), .B2(\mem[0][1] ), 
        .ZN(n1113) );
  INV_X1 U528 ( .A(n1112), .ZN(n810) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n844), .B1(n1114), .B2(\mem[0][2] ), 
        .ZN(n1112) );
  INV_X1 U530 ( .A(n1111), .ZN(n809) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n844), .B1(n1114), .B2(\mem[0][3] ), 
        .ZN(n1111) );
  INV_X1 U532 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n844), .B1(n1114), .B2(\mem[0][4] ), 
        .ZN(n1110) );
  INV_X1 U534 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n844), .B1(n1114), .B2(\mem[0][5] ), 
        .ZN(n1109) );
  INV_X1 U536 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n844), .B1(n1114), .B2(\mem[0][6] ), 
        .ZN(n1108) );
  INV_X1 U538 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n844), .B1(n1114), .B2(\mem[0][7] ), 
        .ZN(n1107) );
  INV_X1 U540 ( .A(n1104), .ZN(n804) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n843), .B1(n1103), .B2(\mem[1][0] ), 
        .ZN(n1104) );
  INV_X1 U542 ( .A(n1102), .ZN(n803) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n843), .B1(n1103), .B2(\mem[1][1] ), 
        .ZN(n1102) );
  INV_X1 U544 ( .A(n1101), .ZN(n802) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n843), .B1(n1103), .B2(\mem[1][2] ), 
        .ZN(n1101) );
  INV_X1 U546 ( .A(n1100), .ZN(n801) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n843), .B1(n1103), .B2(\mem[1][3] ), 
        .ZN(n1100) );
  INV_X1 U548 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n843), .B1(n1103), .B2(\mem[1][4] ), 
        .ZN(n1099) );
  INV_X1 U550 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n843), .B1(n1103), .B2(\mem[1][5] ), 
        .ZN(n1098) );
  INV_X1 U552 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n843), .B1(n1103), .B2(\mem[1][6] ), 
        .ZN(n1097) );
  INV_X1 U554 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n843), .B1(n1103), .B2(\mem[1][7] ), 
        .ZN(n1096) );
  INV_X1 U556 ( .A(n1094), .ZN(n796) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n842), .B1(n1093), .B2(\mem[2][0] ), 
        .ZN(n1094) );
  INV_X1 U558 ( .A(n1092), .ZN(n795) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n842), .B1(n1093), .B2(\mem[2][1] ), 
        .ZN(n1092) );
  INV_X1 U560 ( .A(n1091), .ZN(n794) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n842), .B1(n1093), .B2(\mem[2][2] ), 
        .ZN(n1091) );
  INV_X1 U562 ( .A(n1090), .ZN(n793) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n842), .B1(n1093), .B2(\mem[2][3] ), 
        .ZN(n1090) );
  INV_X1 U564 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n842), .B1(n1093), .B2(\mem[2][4] ), 
        .ZN(n1089) );
  INV_X1 U566 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n842), .B1(n1093), .B2(\mem[2][5] ), 
        .ZN(n1088) );
  INV_X1 U568 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n842), .B1(n1093), .B2(\mem[2][6] ), 
        .ZN(n1087) );
  INV_X1 U570 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n842), .B1(n1093), .B2(\mem[2][7] ), 
        .ZN(n1086) );
  INV_X1 U572 ( .A(n1084), .ZN(n788) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n841), .B1(n1083), .B2(\mem[3][0] ), 
        .ZN(n1084) );
  INV_X1 U574 ( .A(n1082), .ZN(n787) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n841), .B1(n1083), .B2(\mem[3][1] ), 
        .ZN(n1082) );
  INV_X1 U576 ( .A(n1081), .ZN(n786) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n841), .B1(n1083), .B2(\mem[3][2] ), 
        .ZN(n1081) );
  INV_X1 U578 ( .A(n1080), .ZN(n785) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n841), .B1(n1083), .B2(\mem[3][3] ), 
        .ZN(n1080) );
  INV_X1 U580 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n841), .B1(n1083), .B2(\mem[3][4] ), 
        .ZN(n1079) );
  INV_X1 U582 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n841), .B1(n1083), .B2(\mem[3][5] ), 
        .ZN(n1078) );
  INV_X1 U584 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n841), .B1(n1083), .B2(\mem[3][6] ), 
        .ZN(n1077) );
  INV_X1 U586 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n841), .B1(n1083), .B2(\mem[3][7] ), 
        .ZN(n1076) );
  INV_X1 U588 ( .A(n1074), .ZN(n780) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n840), .B1(n1073), .B2(\mem[4][0] ), 
        .ZN(n1074) );
  INV_X1 U590 ( .A(n1072), .ZN(n779) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n840), .B1(n1073), .B2(\mem[4][1] ), 
        .ZN(n1072) );
  INV_X1 U592 ( .A(n1071), .ZN(n778) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n840), .B1(n1073), .B2(\mem[4][2] ), 
        .ZN(n1071) );
  INV_X1 U594 ( .A(n1070), .ZN(n777) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n840), .B1(n1073), .B2(\mem[4][3] ), 
        .ZN(n1070) );
  INV_X1 U596 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n840), .B1(n1073), .B2(\mem[4][4] ), 
        .ZN(n1069) );
  INV_X1 U598 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n840), .B1(n1073), .B2(\mem[4][5] ), 
        .ZN(n1068) );
  INV_X1 U600 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n840), .B1(n1073), .B2(\mem[4][6] ), 
        .ZN(n1067) );
  INV_X1 U602 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n840), .B1(n1073), .B2(\mem[4][7] ), 
        .ZN(n1066) );
  INV_X1 U604 ( .A(N13), .ZN(n845) );
  INV_X1 U605 ( .A(N14), .ZN(n846) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n248), .Z(n4) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n248), .Z(n5) );
  MUX2_X1 U608 ( .A(n5), .B(n4), .S(n245), .Z(n6) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n248), .Z(n7) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n248), .Z(n8) );
  MUX2_X1 U611 ( .A(n8), .B(n7), .S(n247), .Z(n9) );
  MUX2_X1 U612 ( .A(n9), .B(n6), .S(n244), .Z(n10) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n248), .Z(n11) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n248), .Z(n12) );
  MUX2_X1 U615 ( .A(n12), .B(n11), .S(n246), .Z(n13) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n248), .Z(n14) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n248), .Z(n15) );
  MUX2_X1 U618 ( .A(n15), .B(n14), .S(n246), .Z(n16) );
  MUX2_X1 U619 ( .A(n16), .B(n13), .S(n244), .Z(n17) );
  MUX2_X1 U620 ( .A(n17), .B(n10), .S(N13), .Z(n18) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n248), .Z(n19) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n253), .Z(n20) );
  MUX2_X1 U623 ( .A(n20), .B(n19), .S(n245), .Z(n21) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n248), .Z(n22) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(N10), .Z(n23) );
  MUX2_X1 U626 ( .A(n23), .B(n22), .S(n245), .Z(n24) );
  MUX2_X1 U627 ( .A(n24), .B(n21), .S(n244), .Z(n25) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n248), .Z(n26) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n253), .Z(n27) );
  MUX2_X1 U630 ( .A(n27), .B(n26), .S(n245), .Z(n28) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n253), .Z(n29) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(N10), .Z(n30) );
  MUX2_X1 U633 ( .A(n30), .B(n29), .S(n245), .Z(n31) );
  MUX2_X1 U634 ( .A(n31), .B(n28), .S(N12), .Z(n32) );
  MUX2_X1 U635 ( .A(n32), .B(n25), .S(N13), .Z(n33) );
  MUX2_X1 U636 ( .A(n33), .B(n18), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n253), .Z(n34) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(N10), .Z(n35) );
  MUX2_X1 U639 ( .A(n35), .B(n34), .S(n245), .Z(n36) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n253), .Z(n37) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(N10), .Z(n38) );
  MUX2_X1 U642 ( .A(n38), .B(n37), .S(n245), .Z(n39) );
  MUX2_X1 U643 ( .A(n39), .B(n36), .S(n244), .Z(n40) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n253), .Z(n41) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(N10), .Z(n42) );
  MUX2_X1 U646 ( .A(n42), .B(n41), .S(n245), .Z(n43) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(N10), .Z(n44) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(N10), .Z(n45) );
  MUX2_X1 U649 ( .A(n45), .B(n44), .S(n245), .Z(n46) );
  MUX2_X1 U650 ( .A(n46), .B(n43), .S(N12), .Z(n47) );
  MUX2_X1 U651 ( .A(n47), .B(n40), .S(N13), .Z(n48) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(N10), .Z(n49) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(N10), .Z(n50) );
  MUX2_X1 U654 ( .A(n50), .B(n49), .S(n245), .Z(n51) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(N10), .Z(n52) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(N10), .Z(n53) );
  MUX2_X1 U657 ( .A(n53), .B(n52), .S(n245), .Z(n54) );
  MUX2_X1 U658 ( .A(n54), .B(n51), .S(n244), .Z(n55) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(N10), .Z(n56) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(N10), .Z(n57) );
  MUX2_X1 U661 ( .A(n57), .B(n56), .S(n245), .Z(n58) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(N10), .Z(n59) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n253), .Z(n60) );
  MUX2_X1 U664 ( .A(n60), .B(n59), .S(n245), .Z(n61) );
  MUX2_X1 U665 ( .A(n61), .B(n58), .S(N12), .Z(n62) );
  MUX2_X1 U666 ( .A(n62), .B(n55), .S(N13), .Z(n63) );
  MUX2_X1 U667 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n249), .Z(n64) );
  MUX2_X1 U668 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n249), .Z(n65) );
  MUX2_X1 U669 ( .A(n65), .B(n64), .S(n246), .Z(n66) );
  MUX2_X1 U670 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n249), .Z(n67) );
  MUX2_X1 U671 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n249), .Z(n68) );
  MUX2_X1 U672 ( .A(n68), .B(n67), .S(n246), .Z(n69) );
  MUX2_X1 U673 ( .A(n69), .B(n66), .S(n244), .Z(n70) );
  MUX2_X1 U674 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n249), .Z(n71) );
  MUX2_X1 U675 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n249), .Z(n72) );
  MUX2_X1 U676 ( .A(n72), .B(n71), .S(n246), .Z(n73) );
  MUX2_X1 U677 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n249), .Z(n74) );
  MUX2_X1 U678 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n249), .Z(n75) );
  MUX2_X1 U679 ( .A(n75), .B(n74), .S(n246), .Z(n76) );
  MUX2_X1 U680 ( .A(n76), .B(n73), .S(n244), .Z(n77) );
  MUX2_X1 U681 ( .A(n77), .B(n70), .S(N13), .Z(n78) );
  MUX2_X1 U682 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n249), .Z(n79) );
  MUX2_X1 U683 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n249), .Z(n80) );
  MUX2_X1 U684 ( .A(n80), .B(n79), .S(n246), .Z(n81) );
  MUX2_X1 U685 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n249), .Z(n82) );
  MUX2_X1 U686 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n249), .Z(n83) );
  MUX2_X1 U687 ( .A(n83), .B(n82), .S(n246), .Z(n84) );
  MUX2_X1 U688 ( .A(n84), .B(n81), .S(n244), .Z(n85) );
  MUX2_X1 U689 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n250), .Z(n86) );
  MUX2_X1 U690 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n250), .Z(n87) );
  MUX2_X1 U691 ( .A(n87), .B(n86), .S(n246), .Z(n88) );
  MUX2_X1 U692 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n250), .Z(n89) );
  MUX2_X1 U693 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n250), .Z(n90) );
  MUX2_X1 U694 ( .A(n90), .B(n89), .S(n246), .Z(n91) );
  MUX2_X1 U695 ( .A(n91), .B(n88), .S(n244), .Z(n92) );
  MUX2_X1 U696 ( .A(n92), .B(n85), .S(N13), .Z(n93) );
  MUX2_X1 U697 ( .A(n93), .B(n78), .S(N14), .Z(N20) );
  MUX2_X1 U698 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U699 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n95) );
  MUX2_X1 U700 ( .A(n95), .B(n94), .S(n246), .Z(n96) );
  MUX2_X1 U701 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n250), .Z(n97) );
  MUX2_X1 U702 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n250), .Z(n98) );
  MUX2_X1 U703 ( .A(n98), .B(n97), .S(n246), .Z(n99) );
  MUX2_X1 U704 ( .A(n99), .B(n96), .S(n244), .Z(n100) );
  MUX2_X1 U705 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n101) );
  MUX2_X1 U706 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n250), .Z(n102) );
  MUX2_X1 U707 ( .A(n102), .B(n101), .S(n246), .Z(n103) );
  MUX2_X1 U708 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n250), .Z(n104) );
  MUX2_X1 U709 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n250), .Z(n105) );
  MUX2_X1 U710 ( .A(n105), .B(n104), .S(n246), .Z(n106) );
  MUX2_X1 U711 ( .A(n106), .B(n103), .S(n244), .Z(n107) );
  MUX2_X1 U712 ( .A(n107), .B(n100), .S(N13), .Z(n108) );
  MUX2_X1 U713 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n251), .Z(n109) );
  MUX2_X1 U714 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n250), .Z(n110) );
  MUX2_X1 U715 ( .A(n110), .B(n109), .S(n247), .Z(n111) );
  MUX2_X1 U716 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n251), .Z(n112) );
  MUX2_X1 U717 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n251), .Z(n113) );
  MUX2_X1 U718 ( .A(n113), .B(n112), .S(n247), .Z(n114) );
  MUX2_X1 U719 ( .A(n114), .B(n111), .S(n244), .Z(n115) );
  MUX2_X1 U720 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n252), .Z(n116) );
  MUX2_X1 U721 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n252), .Z(n117) );
  MUX2_X1 U722 ( .A(n117), .B(n116), .S(n247), .Z(n118) );
  MUX2_X1 U723 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n249), .Z(n119) );
  MUX2_X1 U724 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n250), .Z(n120) );
  MUX2_X1 U725 ( .A(n120), .B(n119), .S(n247), .Z(n121) );
  MUX2_X1 U726 ( .A(n121), .B(n118), .S(n244), .Z(n122) );
  MUX2_X1 U727 ( .A(n122), .B(n115), .S(N13), .Z(n123) );
  MUX2_X1 U728 ( .A(n123), .B(n108), .S(N14), .Z(N19) );
  MUX2_X1 U729 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n253), .Z(n124) );
  MUX2_X1 U730 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n250), .Z(n125) );
  MUX2_X1 U731 ( .A(n125), .B(n124), .S(n247), .Z(n126) );
  MUX2_X1 U732 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n249), .Z(n127) );
  MUX2_X1 U733 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n249), .Z(n128) );
  MUX2_X1 U734 ( .A(n128), .B(n127), .S(n247), .Z(n129) );
  MUX2_X1 U735 ( .A(n129), .B(n126), .S(n244), .Z(n130) );
  MUX2_X1 U736 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n253), .Z(n131) );
  MUX2_X1 U737 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n253), .Z(n132) );
  MUX2_X1 U738 ( .A(n132), .B(n131), .S(n247), .Z(n133) );
  MUX2_X1 U739 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n253), .Z(n134) );
  MUX2_X1 U740 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n253), .Z(n135) );
  MUX2_X1 U741 ( .A(n135), .B(n134), .S(n247), .Z(n136) );
  MUX2_X1 U742 ( .A(n136), .B(n133), .S(n244), .Z(n137) );
  MUX2_X1 U743 ( .A(n137), .B(n130), .S(N13), .Z(n138) );
  MUX2_X1 U744 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n253), .Z(n139) );
  MUX2_X1 U745 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n253), .Z(n140) );
  MUX2_X1 U746 ( .A(n140), .B(n139), .S(n247), .Z(n141) );
  MUX2_X1 U747 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n253), .Z(n142) );
  MUX2_X1 U748 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n253), .Z(n143) );
  MUX2_X1 U749 ( .A(n143), .B(n142), .S(n247), .Z(n144) );
  MUX2_X1 U750 ( .A(n144), .B(n141), .S(n244), .Z(n145) );
  MUX2_X1 U751 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n253), .Z(n146) );
  MUX2_X1 U752 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n253), .Z(n147) );
  MUX2_X1 U753 ( .A(n147), .B(n146), .S(n247), .Z(n148) );
  MUX2_X1 U754 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n253), .Z(n149) );
  MUX2_X1 U755 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n253), .Z(n150) );
  MUX2_X1 U756 ( .A(n150), .B(n149), .S(n247), .Z(n151) );
  MUX2_X1 U757 ( .A(n151), .B(n148), .S(n244), .Z(n152) );
  MUX2_X1 U758 ( .A(n152), .B(n145), .S(N13), .Z(n153) );
  MUX2_X1 U759 ( .A(n153), .B(n138), .S(N14), .Z(N18) );
  MUX2_X1 U760 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n248), .Z(n154) );
  MUX2_X1 U761 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n248), .Z(n155) );
  MUX2_X1 U762 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U763 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n248), .Z(n157) );
  MUX2_X1 U764 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n248), .Z(n158) );
  MUX2_X1 U765 ( .A(n158), .B(n157), .S(N11), .Z(n159) );
  MUX2_X1 U766 ( .A(n159), .B(n156), .S(n244), .Z(n160) );
  MUX2_X1 U767 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n248), .Z(n161) );
  MUX2_X1 U768 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n248), .Z(n162) );
  MUX2_X1 U769 ( .A(n162), .B(n161), .S(N11), .Z(n163) );
  MUX2_X1 U770 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n248), .Z(n164) );
  MUX2_X1 U771 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n248), .Z(n165) );
  MUX2_X1 U772 ( .A(n165), .B(n164), .S(n247), .Z(n166) );
  MUX2_X1 U773 ( .A(n166), .B(n163), .S(N12), .Z(n167) );
  MUX2_X1 U774 ( .A(n167), .B(n160), .S(N13), .Z(n168) );
  MUX2_X1 U775 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n248), .Z(n169) );
  MUX2_X1 U776 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n248), .Z(n170) );
  MUX2_X1 U777 ( .A(n170), .B(n169), .S(N11), .Z(n171) );
  MUX2_X1 U778 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n248), .Z(n172) );
  MUX2_X1 U779 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n248), .Z(n173) );
  MUX2_X1 U780 ( .A(n173), .B(n172), .S(n245), .Z(n174) );
  MUX2_X1 U781 ( .A(n174), .B(n171), .S(n244), .Z(n175) );
  MUX2_X1 U782 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n251), .Z(n176) );
  MUX2_X1 U783 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n251), .Z(n177) );
  MUX2_X1 U784 ( .A(n177), .B(n176), .S(N11), .Z(n178) );
  MUX2_X1 U785 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n251), .Z(n179) );
  MUX2_X1 U786 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n251), .Z(n180) );
  MUX2_X1 U787 ( .A(n180), .B(n179), .S(n247), .Z(n181) );
  MUX2_X1 U788 ( .A(n181), .B(n178), .S(N12), .Z(n182) );
  MUX2_X1 U789 ( .A(n182), .B(n175), .S(N13), .Z(n183) );
  MUX2_X1 U790 ( .A(n183), .B(n168), .S(N14), .Z(N17) );
  MUX2_X1 U791 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n251), .Z(n184) );
  MUX2_X1 U792 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n251), .Z(n185) );
  MUX2_X1 U793 ( .A(n185), .B(n184), .S(N11), .Z(n186) );
  MUX2_X1 U794 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n251), .Z(n187) );
  MUX2_X1 U795 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n251), .Z(n188) );
  MUX2_X1 U796 ( .A(n188), .B(n187), .S(N11), .Z(n189) );
  MUX2_X1 U797 ( .A(n189), .B(n186), .S(n244), .Z(n190) );
  MUX2_X1 U798 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n251), .Z(n191) );
  MUX2_X1 U799 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n251), .Z(n192) );
  MUX2_X1 U800 ( .A(n192), .B(n191), .S(N11), .Z(n193) );
  MUX2_X1 U801 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n251), .Z(n194) );
  MUX2_X1 U802 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n251), .Z(n195) );
  MUX2_X1 U803 ( .A(n195), .B(n194), .S(n245), .Z(n196) );
  MUX2_X1 U804 ( .A(n196), .B(n193), .S(N12), .Z(n197) );
  MUX2_X1 U805 ( .A(n197), .B(n190), .S(N13), .Z(n198) );
  MUX2_X1 U806 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n252), .Z(n199) );
  MUX2_X1 U807 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n252), .Z(n200) );
  MUX2_X1 U808 ( .A(n200), .B(n199), .S(n246), .Z(n201) );
  MUX2_X1 U809 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n252), .Z(n202) );
  MUX2_X1 U810 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n252), .Z(n203) );
  MUX2_X1 U811 ( .A(n203), .B(n202), .S(n246), .Z(n204) );
  MUX2_X1 U812 ( .A(n204), .B(n201), .S(n244), .Z(n205) );
  MUX2_X1 U813 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n252), .Z(n206) );
  MUX2_X1 U814 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n252), .Z(n207) );
  MUX2_X1 U815 ( .A(n207), .B(n206), .S(n246), .Z(n208) );
  MUX2_X1 U816 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n252), .Z(n209) );
  MUX2_X1 U817 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n252), .Z(n210) );
  MUX2_X1 U818 ( .A(n210), .B(n209), .S(N11), .Z(n211) );
  MUX2_X1 U819 ( .A(n211), .B(n208), .S(N12), .Z(n212) );
  MUX2_X1 U820 ( .A(n212), .B(n205), .S(N13), .Z(n213) );
  MUX2_X1 U821 ( .A(n213), .B(n198), .S(N14), .Z(N16) );
  MUX2_X1 U822 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n252), .Z(n214) );
  MUX2_X1 U823 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n252), .Z(n215) );
  MUX2_X1 U824 ( .A(n215), .B(n214), .S(n245), .Z(n216) );
  MUX2_X1 U825 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n252), .Z(n217) );
  MUX2_X1 U826 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n252), .Z(n218) );
  MUX2_X1 U827 ( .A(n218), .B(n217), .S(n245), .Z(n219) );
  MUX2_X1 U828 ( .A(n219), .B(n216), .S(n244), .Z(n220) );
  MUX2_X1 U829 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n252), .Z(n221) );
  MUX2_X1 U830 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n250), .Z(n222) );
  MUX2_X1 U831 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U832 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n251), .Z(n224) );
  MUX2_X1 U833 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n249), .Z(n225) );
  MUX2_X1 U834 ( .A(n225), .B(n224), .S(N11), .Z(n226) );
  MUX2_X1 U835 ( .A(n226), .B(n223), .S(N12), .Z(n227) );
  MUX2_X1 U836 ( .A(n227), .B(n220), .S(N13), .Z(n228) );
  MUX2_X1 U837 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n249), .Z(n229) );
  MUX2_X1 U838 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n252), .Z(n230) );
  MUX2_X1 U839 ( .A(n230), .B(n229), .S(n247), .Z(n231) );
  MUX2_X1 U840 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n250), .Z(n232) );
  MUX2_X1 U841 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n252), .Z(n233) );
  MUX2_X1 U842 ( .A(n233), .B(n232), .S(N11), .Z(n234) );
  MUX2_X1 U843 ( .A(n234), .B(n231), .S(n244), .Z(n235) );
  MUX2_X1 U844 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n249), .Z(n236) );
  MUX2_X1 U845 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n250), .Z(n237) );
  MUX2_X1 U846 ( .A(n237), .B(n236), .S(n247), .Z(n238) );
  MUX2_X1 U847 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n251), .Z(n239) );
  MUX2_X1 U848 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n251), .Z(n240) );
  MUX2_X1 U849 ( .A(n240), .B(n239), .S(N11), .Z(n241) );
  MUX2_X1 U850 ( .A(n241), .B(n238), .S(N12), .Z(n242) );
  MUX2_X1 U851 ( .A(n242), .B(n235), .S(N13), .Z(n243) );
  MUX2_X1 U852 ( .A(n243), .B(n228), .S(N14), .Z(N15) );
  CLKBUF_X1 U853 ( .A(N10), .Z(n248) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_6 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X2 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(n250), .Z(n249) );
  BUF_X1 U4 ( .A(n250), .Z(n246) );
  BUF_X1 U5 ( .A(n250), .Z(n247) );
  BUF_X1 U6 ( .A(N10), .Z(n248) );
  BUF_X1 U7 ( .A(n250), .Z(n245) );
  BUF_X1 U8 ( .A(N10), .Z(n250) );
  INV_X1 U9 ( .A(n1111), .ZN(n841) );
  INV_X1 U10 ( .A(n1100), .ZN(n840) );
  INV_X1 U11 ( .A(n1090), .ZN(n839) );
  INV_X1 U12 ( .A(n1080), .ZN(n838) );
  INV_X1 U13 ( .A(n1070), .ZN(n837) );
  INV_X1 U14 ( .A(n1060), .ZN(n836) );
  INV_X1 U15 ( .A(n1051), .ZN(n835) );
  INV_X1 U16 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U19 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U20 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U21 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U22 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U23 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U24 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U26 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U27 ( .A(n1131), .ZN(n816) );
  INV_X1 U28 ( .A(n1121), .ZN(n815) );
  INV_X1 U29 ( .A(n887), .ZN(n814) );
  INV_X1 U30 ( .A(n878), .ZN(n813) );
  INV_X1 U31 ( .A(n869), .ZN(n812) );
  INV_X1 U32 ( .A(n860), .ZN(n811) );
  INV_X1 U33 ( .A(n851), .ZN(n810) );
  INV_X1 U34 ( .A(n987), .ZN(n828) );
  INV_X1 U35 ( .A(n978), .ZN(n827) );
  INV_X1 U36 ( .A(n969), .ZN(n826) );
  INV_X1 U37 ( .A(n914), .ZN(n820) );
  INV_X1 U38 ( .A(n905), .ZN(n819) );
  INV_X1 U39 ( .A(n896), .ZN(n818) );
  INV_X1 U40 ( .A(n1033), .ZN(n833) );
  INV_X1 U41 ( .A(n1023), .ZN(n832) );
  INV_X1 U42 ( .A(n1014), .ZN(n831) );
  INV_X1 U43 ( .A(n1005), .ZN(n830) );
  INV_X1 U44 ( .A(n996), .ZN(n829) );
  INV_X1 U45 ( .A(n960), .ZN(n825) );
  INV_X1 U46 ( .A(n950), .ZN(n824) );
  INV_X1 U47 ( .A(n941), .ZN(n823) );
  INV_X1 U48 ( .A(n932), .ZN(n822) );
  INV_X1 U49 ( .A(n923), .ZN(n821) );
  INV_X1 U50 ( .A(n1142), .ZN(n817) );
  BUF_X1 U51 ( .A(N11), .Z(n242) );
  BUF_X1 U52 ( .A(N11), .Z(n243) );
  BUF_X1 U53 ( .A(N11), .Z(n244) );
  INV_X1 U54 ( .A(N10), .ZN(n251) );
  BUF_X1 U55 ( .A(N12), .Z(n241) );
  NOR3_X1 U56 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U57 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U58 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U60 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U62 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U63 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U64 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U65 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U67 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U69 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U70 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U71 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U72 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U73 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U74 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U75 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U76 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U77 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U79 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U81 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U82 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U83 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U84 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U85 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U86 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U88 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U89 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U90 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U92 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U94 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U95 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U96 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U97 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U98 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U99 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U100 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U101 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U102 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U103 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U104 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U105 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U106 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U107 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U108 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U109 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U110 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U111 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U112 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U113 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U114 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U115 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U116 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U117 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U118 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U119 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U120 ( .A(n988), .ZN(n705) );
  AOI22_X1 U121 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U122 ( .A(n986), .ZN(n704) );
  AOI22_X1 U123 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U124 ( .A(n985), .ZN(n703) );
  AOI22_X1 U125 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U126 ( .A(n984), .ZN(n702) );
  AOI22_X1 U127 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U128 ( .A(n983), .ZN(n701) );
  AOI22_X1 U129 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U130 ( .A(n982), .ZN(n700) );
  AOI22_X1 U131 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U132 ( .A(n981), .ZN(n699) );
  AOI22_X1 U133 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U134 ( .A(n980), .ZN(n698) );
  AOI22_X1 U135 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U136 ( .A(n943), .ZN(n666) );
  AOI22_X1 U137 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U138 ( .A(n915), .ZN(n641) );
  AOI22_X1 U139 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U140 ( .A(n913), .ZN(n640) );
  AOI22_X1 U141 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U142 ( .A(n912), .ZN(n639) );
  AOI22_X1 U143 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U144 ( .A(n911), .ZN(n638) );
  AOI22_X1 U145 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U146 ( .A(n910), .ZN(n637) );
  AOI22_X1 U147 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U148 ( .A(n909), .ZN(n636) );
  AOI22_X1 U149 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U150 ( .A(n908), .ZN(n635) );
  AOI22_X1 U151 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U152 ( .A(n907), .ZN(n634) );
  AOI22_X1 U153 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U154 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U155 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U156 ( .A(n944), .ZN(n667) );
  AOI22_X1 U157 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U158 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U159 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U160 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U161 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U162 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U163 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U164 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U165 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U166 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U167 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U168 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U169 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U170 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U171 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U172 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U173 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U174 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U175 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U176 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U177 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U178 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U179 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U180 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U181 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U182 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U183 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U184 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U185 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U186 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U187 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U188 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U189 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U190 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U191 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U192 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U193 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U194 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U195 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U196 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U197 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U198 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U199 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U200 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U201 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U202 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U203 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U204 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U205 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U206 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U207 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U208 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U209 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U210 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U211 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U212 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U213 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U214 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U215 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U216 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U217 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U218 ( .A(n999), .ZN(n715) );
  AOI22_X1 U219 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U220 ( .A(n998), .ZN(n714) );
  AOI22_X1 U221 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U222 ( .A(n951), .ZN(n673) );
  AOI22_X1 U223 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U224 ( .A(n949), .ZN(n672) );
  AOI22_X1 U225 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U226 ( .A(n948), .ZN(n671) );
  AOI22_X1 U227 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U228 ( .A(n947), .ZN(n670) );
  AOI22_X1 U229 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U230 ( .A(n946), .ZN(n669) );
  AOI22_X1 U231 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U232 ( .A(n945), .ZN(n668) );
  AOI22_X1 U233 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U234 ( .A(n979), .ZN(n697) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U236 ( .A(n977), .ZN(n696) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U238 ( .A(n976), .ZN(n695) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U240 ( .A(n975), .ZN(n694) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U242 ( .A(n974), .ZN(n693) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U244 ( .A(n973), .ZN(n692) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U246 ( .A(n972), .ZN(n691) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U248 ( .A(n971), .ZN(n690) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U250 ( .A(n970), .ZN(n689) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U252 ( .A(n968), .ZN(n688) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U254 ( .A(n967), .ZN(n687) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U256 ( .A(n966), .ZN(n686) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U258 ( .A(n965), .ZN(n685) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U260 ( .A(n964), .ZN(n684) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U262 ( .A(n963), .ZN(n683) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U264 ( .A(n962), .ZN(n682) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U266 ( .A(n942), .ZN(n665) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U268 ( .A(n940), .ZN(n664) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U270 ( .A(n939), .ZN(n663) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U272 ( .A(n938), .ZN(n662) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U274 ( .A(n937), .ZN(n661) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U276 ( .A(n936), .ZN(n660) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U278 ( .A(n935), .ZN(n659) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U280 ( .A(n934), .ZN(n658) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U282 ( .A(n933), .ZN(n657) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U284 ( .A(n931), .ZN(n656) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U286 ( .A(n930), .ZN(n655) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U288 ( .A(n929), .ZN(n654) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U290 ( .A(n928), .ZN(n653) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U292 ( .A(n927), .ZN(n652) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U294 ( .A(n926), .ZN(n651) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U296 ( .A(n925), .ZN(n650) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U298 ( .A(n906), .ZN(n633) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U300 ( .A(n904), .ZN(n632) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U302 ( .A(n903), .ZN(n631) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U304 ( .A(n902), .ZN(n630) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U306 ( .A(n901), .ZN(n629) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U308 ( .A(n900), .ZN(n628) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U310 ( .A(n899), .ZN(n627) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U312 ( .A(n898), .ZN(n626) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U314 ( .A(n897), .ZN(n625) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U316 ( .A(n895), .ZN(n624) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U318 ( .A(n894), .ZN(n623) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U320 ( .A(n893), .ZN(n622) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U322 ( .A(n892), .ZN(n621) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U324 ( .A(n891), .ZN(n620) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U326 ( .A(n890), .ZN(n619) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U328 ( .A(n889), .ZN(n618) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U330 ( .A(N12), .ZN(n253) );
  INV_X1 U331 ( .A(N11), .ZN(n252) );
  INV_X1 U332 ( .A(n997), .ZN(n713) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U334 ( .A(n995), .ZN(n712) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U336 ( .A(n994), .ZN(n711) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U338 ( .A(n993), .ZN(n710) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U340 ( .A(n992), .ZN(n709) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U342 ( .A(n991), .ZN(n708) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U344 ( .A(n990), .ZN(n707) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U346 ( .A(n989), .ZN(n706) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U348 ( .A(n924), .ZN(n649) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U350 ( .A(n922), .ZN(n648) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U352 ( .A(n921), .ZN(n647) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U354 ( .A(n920), .ZN(n646) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U356 ( .A(n919), .ZN(n645) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U358 ( .A(n918), .ZN(n644) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U360 ( .A(n917), .ZN(n643) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U362 ( .A(n916), .ZN(n642) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U364 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U366 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U368 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U370 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U372 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U374 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U376 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U378 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U380 ( .A(n961), .ZN(n681) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U382 ( .A(n959), .ZN(n680) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U384 ( .A(n958), .ZN(n679) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U386 ( .A(n957), .ZN(n678) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U388 ( .A(n956), .ZN(n677) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U390 ( .A(n955), .ZN(n676) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U392 ( .A(n954), .ZN(n675) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U394 ( .A(n953), .ZN(n674) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U396 ( .A(n888), .ZN(n617) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U398 ( .A(n886), .ZN(n616) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U400 ( .A(n885), .ZN(n615) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U402 ( .A(n884), .ZN(n614) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U404 ( .A(n883), .ZN(n613) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U406 ( .A(n882), .ZN(n612) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U408 ( .A(n881), .ZN(n611) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U410 ( .A(n880), .ZN(n610) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U412 ( .A(n879), .ZN(n609) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U414 ( .A(n877), .ZN(n608) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U416 ( .A(n876), .ZN(n607) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U418 ( .A(n875), .ZN(n606) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U420 ( .A(n874), .ZN(n605) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U422 ( .A(n873), .ZN(n604) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U424 ( .A(n872), .ZN(n603) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U426 ( .A(n871), .ZN(n602) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U428 ( .A(n870), .ZN(n601) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U430 ( .A(n868), .ZN(n600) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U432 ( .A(n867), .ZN(n599) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U434 ( .A(n866), .ZN(n598) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U436 ( .A(n865), .ZN(n597) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U438 ( .A(n864), .ZN(n596) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U440 ( .A(n863), .ZN(n595) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U442 ( .A(n862), .ZN(n594) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U444 ( .A(n861), .ZN(n293) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U446 ( .A(n859), .ZN(n292) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U448 ( .A(n858), .ZN(n291) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U450 ( .A(n857), .ZN(n290) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U452 ( .A(n856), .ZN(n289) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U454 ( .A(n855), .ZN(n288) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U456 ( .A(n854), .ZN(n287) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U458 ( .A(n853), .ZN(n286) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U460 ( .A(n852), .ZN(n285) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U462 ( .A(n850), .ZN(n284) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U464 ( .A(n849), .ZN(n283) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U466 ( .A(n848), .ZN(n282) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U468 ( .A(n847), .ZN(n281) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U470 ( .A(n846), .ZN(n280) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U472 ( .A(n845), .ZN(n279) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U474 ( .A(n844), .ZN(n278) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U476 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U477 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U478 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U479 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U480 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U481 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U482 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U483 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U484 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U485 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U486 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U487 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U488 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U489 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U490 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U491 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U492 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U494 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U496 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U498 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U500 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U502 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U504 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U506 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U508 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U510 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U512 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U514 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U516 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U518 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U520 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U522 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U524 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U526 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U528 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U530 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U532 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U534 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U536 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U538 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U540 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U542 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U544 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U546 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U548 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U550 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U552 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U554 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U556 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U558 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U560 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U562 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U564 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U566 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U568 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U570 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U572 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U574 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U576 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U578 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U580 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U582 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U584 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U586 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U588 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U590 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U592 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U594 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U596 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U598 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U600 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U602 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U604 ( .A(N13), .ZN(n842) );
  INV_X1 U605 ( .A(N14), .ZN(n843) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n248), .Z(n1) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n248), .Z(n2) );
  MUX2_X1 U608 ( .A(n2), .B(n1), .S(n242), .Z(n3) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n248), .Z(n4) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n248), .Z(n5) );
  MUX2_X1 U611 ( .A(n5), .B(n4), .S(n244), .Z(n6) );
  MUX2_X1 U612 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n248), .Z(n8) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n248), .Z(n9) );
  MUX2_X1 U615 ( .A(n9), .B(n8), .S(n243), .Z(n10) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n248), .Z(n11) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n248), .Z(n12) );
  MUX2_X1 U618 ( .A(n12), .B(n11), .S(N11), .Z(n13) );
  MUX2_X1 U619 ( .A(n13), .B(n10), .S(n241), .Z(n14) );
  MUX2_X1 U620 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n247), .Z(n16) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n247), .Z(n17) );
  MUX2_X1 U623 ( .A(n17), .B(n16), .S(n242), .Z(n18) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n246), .Z(n20) );
  MUX2_X1 U626 ( .A(n20), .B(n19), .S(n242), .Z(n21) );
  MUX2_X1 U627 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n249), .Z(n23) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n247), .Z(n24) );
  MUX2_X1 U630 ( .A(n24), .B(n23), .S(n242), .Z(n25) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n249), .Z(n26) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n249), .Z(n27) );
  MUX2_X1 U633 ( .A(n27), .B(n26), .S(n242), .Z(n28) );
  MUX2_X1 U634 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U635 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U636 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n246), .Z(n31) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n247), .Z(n32) );
  MUX2_X1 U639 ( .A(n32), .B(n31), .S(n242), .Z(n33) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U642 ( .A(n35), .B(n34), .S(n242), .Z(n36) );
  MUX2_X1 U643 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n245), .Z(n38) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n245), .Z(n39) );
  MUX2_X1 U646 ( .A(n39), .B(n38), .S(n242), .Z(n40) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n245), .Z(n41) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n245), .Z(n42) );
  MUX2_X1 U649 ( .A(n42), .B(n41), .S(n242), .Z(n43) );
  MUX2_X1 U650 ( .A(n43), .B(n40), .S(N12), .Z(n44) );
  MUX2_X1 U651 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n245), .Z(n46) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n245), .Z(n47) );
  MUX2_X1 U654 ( .A(n47), .B(n46), .S(n242), .Z(n48) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n245), .Z(n49) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n245), .Z(n50) );
  MUX2_X1 U657 ( .A(n50), .B(n49), .S(n242), .Z(n51) );
  MUX2_X1 U658 ( .A(n51), .B(n48), .S(N12), .Z(n52) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n245), .Z(n53) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n245), .Z(n54) );
  MUX2_X1 U661 ( .A(n54), .B(n53), .S(n242), .Z(n55) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n245), .Z(n56) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n245), .Z(n57) );
  MUX2_X1 U664 ( .A(n57), .B(n56), .S(n242), .Z(n58) );
  MUX2_X1 U665 ( .A(n58), .B(n55), .S(N12), .Z(n59) );
  MUX2_X1 U666 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U667 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n250), .Z(n61) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n246), .Z(n62) );
  MUX2_X1 U670 ( .A(n62), .B(n61), .S(n243), .Z(n63) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n247), .Z(n64) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n245), .Z(n65) );
  MUX2_X1 U673 ( .A(n65), .B(n64), .S(n243), .Z(n66) );
  MUX2_X1 U674 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n245), .Z(n68) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n246), .Z(n69) );
  MUX2_X1 U677 ( .A(n69), .B(n68), .S(n243), .Z(n70) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n249), .Z(n71) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n249), .Z(n72) );
  MUX2_X1 U680 ( .A(n72), .B(n71), .S(n243), .Z(n73) );
  MUX2_X1 U681 ( .A(n73), .B(n70), .S(n241), .Z(n74) );
  MUX2_X1 U682 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n249), .Z(n76) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n247), .Z(n77) );
  MUX2_X1 U685 ( .A(n77), .B(n76), .S(n243), .Z(n78) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n246), .Z(n79) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n245), .Z(n80) );
  MUX2_X1 U688 ( .A(n80), .B(n79), .S(n243), .Z(n81) );
  MUX2_X1 U689 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n250), .Z(n83) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n250), .Z(n84) );
  MUX2_X1 U692 ( .A(n84), .B(n83), .S(n243), .Z(n85) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n250), .Z(n86) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n250), .Z(n87) );
  MUX2_X1 U695 ( .A(n87), .B(n86), .S(n243), .Z(n88) );
  MUX2_X1 U696 ( .A(n88), .B(n85), .S(n241), .Z(n89) );
  MUX2_X1 U697 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U698 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n250), .Z(n91) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n92) );
  MUX2_X1 U701 ( .A(n92), .B(n91), .S(n243), .Z(n93) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n250), .Z(n95) );
  MUX2_X1 U704 ( .A(n95), .B(n94), .S(n243), .Z(n96) );
  MUX2_X1 U705 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n98) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n250), .Z(n99) );
  MUX2_X1 U708 ( .A(n99), .B(n98), .S(n243), .Z(n100) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n250), .Z(n101) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n250), .Z(n102) );
  MUX2_X1 U711 ( .A(n102), .B(n101), .S(n243), .Z(n103) );
  MUX2_X1 U712 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U713 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n246), .Z(n106) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n246), .Z(n107) );
  MUX2_X1 U716 ( .A(n107), .B(n106), .S(n244), .Z(n108) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n246), .Z(n109) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n246), .Z(n110) );
  MUX2_X1 U719 ( .A(n110), .B(n109), .S(n244), .Z(n111) );
  MUX2_X1 U720 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n246), .Z(n113) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n246), .Z(n114) );
  MUX2_X1 U723 ( .A(n114), .B(n113), .S(n244), .Z(n115) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n246), .Z(n116) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n246), .Z(n117) );
  MUX2_X1 U726 ( .A(n117), .B(n116), .S(n244), .Z(n118) );
  MUX2_X1 U727 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U728 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U729 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n246), .Z(n121) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n246), .Z(n122) );
  MUX2_X1 U732 ( .A(n122), .B(n121), .S(n244), .Z(n123) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n246), .Z(n124) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n246), .Z(n125) );
  MUX2_X1 U735 ( .A(n125), .B(n124), .S(n244), .Z(n126) );
  MUX2_X1 U736 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n247), .Z(n128) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n247), .Z(n129) );
  MUX2_X1 U739 ( .A(n129), .B(n128), .S(n244), .Z(n130) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n247), .Z(n131) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n247), .Z(n132) );
  MUX2_X1 U742 ( .A(n132), .B(n131), .S(n244), .Z(n133) );
  MUX2_X1 U743 ( .A(n133), .B(n130), .S(n241), .Z(n134) );
  MUX2_X1 U744 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n247), .Z(n136) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n247), .Z(n137) );
  MUX2_X1 U747 ( .A(n137), .B(n136), .S(n244), .Z(n138) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n247), .Z(n139) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n247), .Z(n140) );
  MUX2_X1 U750 ( .A(n140), .B(n139), .S(n244), .Z(n141) );
  MUX2_X1 U751 ( .A(n141), .B(n138), .S(n241), .Z(n142) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n247), .Z(n143) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n247), .Z(n144) );
  MUX2_X1 U754 ( .A(n144), .B(n143), .S(n244), .Z(n145) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n247), .Z(n146) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n247), .Z(n147) );
  MUX2_X1 U757 ( .A(n147), .B(n146), .S(n244), .Z(n148) );
  MUX2_X1 U758 ( .A(n148), .B(n145), .S(n241), .Z(n149) );
  MUX2_X1 U759 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U760 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n248), .Z(n151) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n248), .Z(n152) );
  MUX2_X1 U763 ( .A(n152), .B(n151), .S(N11), .Z(n153) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n248), .Z(n154) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n248), .Z(n155) );
  MUX2_X1 U766 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U767 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n248), .Z(n158) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n248), .Z(n159) );
  MUX2_X1 U770 ( .A(n159), .B(n158), .S(N11), .Z(n160) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n248), .Z(n161) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n248), .Z(n162) );
  MUX2_X1 U773 ( .A(n162), .B(n161), .S(N11), .Z(n163) );
  MUX2_X1 U774 ( .A(n163), .B(n160), .S(n241), .Z(n164) );
  MUX2_X1 U775 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n248), .Z(n166) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n248), .Z(n167) );
  MUX2_X1 U778 ( .A(n167), .B(n166), .S(N11), .Z(n168) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n248), .Z(n169) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n248), .Z(n170) );
  MUX2_X1 U781 ( .A(n170), .B(n169), .S(N11), .Z(n171) );
  MUX2_X1 U782 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n250), .Z(n173) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(N10), .Z(n174) );
  MUX2_X1 U785 ( .A(n174), .B(n173), .S(N11), .Z(n175) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n250), .Z(n176) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(N10), .Z(n177) );
  MUX2_X1 U788 ( .A(n177), .B(n176), .S(N11), .Z(n178) );
  MUX2_X1 U789 ( .A(n178), .B(n175), .S(n241), .Z(n179) );
  MUX2_X1 U790 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U791 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(N10), .Z(n181) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(N10), .Z(n182) );
  MUX2_X1 U794 ( .A(n182), .B(n181), .S(N11), .Z(n183) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(N10), .Z(n184) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n250), .Z(n185) );
  MUX2_X1 U797 ( .A(n185), .B(n184), .S(n244), .Z(n186) );
  MUX2_X1 U798 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(N10), .Z(n188) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n250), .Z(n189) );
  MUX2_X1 U801 ( .A(n189), .B(n188), .S(n243), .Z(n190) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(N10), .Z(n191) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n250), .Z(n192) );
  MUX2_X1 U804 ( .A(n192), .B(n191), .S(n244), .Z(n193) );
  MUX2_X1 U805 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U806 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n248), .Z(n196) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(N10), .Z(n197) );
  MUX2_X1 U809 ( .A(n197), .B(n196), .S(n242), .Z(n198) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n250), .Z(n199) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n200) );
  MUX2_X1 U812 ( .A(n200), .B(n199), .S(n244), .Z(n201) );
  MUX2_X1 U813 ( .A(n201), .B(n198), .S(N12), .Z(n202) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n250), .Z(n203) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n204) );
  MUX2_X1 U816 ( .A(n204), .B(n203), .S(n242), .Z(n205) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n206) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n207) );
  MUX2_X1 U819 ( .A(n207), .B(n206), .S(N11), .Z(n208) );
  MUX2_X1 U820 ( .A(n208), .B(n205), .S(N12), .Z(n209) );
  MUX2_X1 U821 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U822 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n248), .Z(n211) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(N10), .Z(n212) );
  MUX2_X1 U825 ( .A(n212), .B(n211), .S(n242), .Z(n213) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n248), .Z(n214) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(N10), .Z(n215) );
  MUX2_X1 U828 ( .A(n215), .B(n214), .S(n242), .Z(n216) );
  MUX2_X1 U829 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n249), .Z(n218) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n249), .Z(n219) );
  MUX2_X1 U832 ( .A(n219), .B(n218), .S(n244), .Z(n220) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n249), .Z(n221) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n249), .Z(n222) );
  MUX2_X1 U835 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U836 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U837 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n249), .Z(n226) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n249), .Z(n227) );
  MUX2_X1 U840 ( .A(n227), .B(n226), .S(n243), .Z(n228) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n249), .Z(n229) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n249), .Z(n230) );
  MUX2_X1 U843 ( .A(n230), .B(n229), .S(n243), .Z(n231) );
  MUX2_X1 U844 ( .A(n231), .B(n228), .S(N12), .Z(n232) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n249), .Z(n233) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n249), .Z(n234) );
  MUX2_X1 U847 ( .A(n234), .B(n233), .S(n243), .Z(n235) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n249), .Z(n236) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n249), .Z(n237) );
  MUX2_X1 U850 ( .A(n237), .B(n236), .S(N11), .Z(n238) );
  MUX2_X1 U851 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U852 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U853 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_5 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  BUF_X1 U3 ( .A(n250), .Z(n248) );
  BUF_X1 U4 ( .A(N10), .Z(n249) );
  BUF_X1 U5 ( .A(n250), .Z(n245) );
  BUF_X1 U6 ( .A(n250), .Z(n246) );
  BUF_X1 U7 ( .A(n250), .Z(n247) );
  BUF_X1 U8 ( .A(N10), .Z(n250) );
  INV_X1 U9 ( .A(n1111), .ZN(n841) );
  INV_X1 U10 ( .A(n1100), .ZN(n840) );
  INV_X1 U11 ( .A(n1090), .ZN(n839) );
  INV_X1 U12 ( .A(n1080), .ZN(n838) );
  INV_X1 U13 ( .A(n1070), .ZN(n837) );
  INV_X1 U14 ( .A(n1060), .ZN(n836) );
  INV_X1 U15 ( .A(n1051), .ZN(n835) );
  INV_X1 U16 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U19 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U20 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U21 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U22 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U23 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U24 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U26 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U27 ( .A(n1131), .ZN(n816) );
  INV_X1 U28 ( .A(n1121), .ZN(n815) );
  INV_X1 U29 ( .A(n887), .ZN(n814) );
  INV_X1 U30 ( .A(n878), .ZN(n813) );
  INV_X1 U31 ( .A(n869), .ZN(n812) );
  INV_X1 U32 ( .A(n860), .ZN(n811) );
  INV_X1 U33 ( .A(n851), .ZN(n810) );
  INV_X1 U34 ( .A(n987), .ZN(n828) );
  INV_X1 U35 ( .A(n978), .ZN(n827) );
  INV_X1 U36 ( .A(n969), .ZN(n826) );
  INV_X1 U37 ( .A(n914), .ZN(n820) );
  INV_X1 U38 ( .A(n905), .ZN(n819) );
  INV_X1 U39 ( .A(n896), .ZN(n818) );
  INV_X1 U40 ( .A(n1033), .ZN(n833) );
  INV_X1 U41 ( .A(n1023), .ZN(n832) );
  INV_X1 U42 ( .A(n1014), .ZN(n831) );
  INV_X1 U43 ( .A(n1005), .ZN(n830) );
  INV_X1 U44 ( .A(n996), .ZN(n829) );
  INV_X1 U45 ( .A(n960), .ZN(n825) );
  INV_X1 U46 ( .A(n950), .ZN(n824) );
  INV_X1 U47 ( .A(n941), .ZN(n823) );
  INV_X1 U48 ( .A(n932), .ZN(n822) );
  INV_X1 U49 ( .A(n923), .ZN(n821) );
  INV_X1 U50 ( .A(n1142), .ZN(n817) );
  BUF_X1 U51 ( .A(N11), .Z(n242) );
  BUF_X1 U52 ( .A(N11), .Z(n243) );
  BUF_X1 U53 ( .A(N11), .Z(n244) );
  INV_X1 U54 ( .A(N10), .ZN(n251) );
  BUF_X1 U55 ( .A(N12), .Z(n241) );
  NOR3_X1 U56 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U57 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U58 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U60 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U62 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U63 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U64 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U65 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U67 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U69 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U70 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U71 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U72 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U73 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U74 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U75 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U76 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U77 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U79 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U81 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U82 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U83 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U84 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U85 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U86 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U88 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U89 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U90 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U92 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U94 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U95 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U96 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U97 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U98 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U99 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U100 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U101 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U102 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U103 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U104 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U105 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U106 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U107 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U108 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U109 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U110 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U111 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U112 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U113 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U114 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U115 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U116 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U117 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U118 ( .A(n988), .ZN(n705) );
  AOI22_X1 U119 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U120 ( .A(n986), .ZN(n704) );
  AOI22_X1 U121 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U122 ( .A(n984), .ZN(n702) );
  AOI22_X1 U123 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U124 ( .A(n983), .ZN(n701) );
  AOI22_X1 U125 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U126 ( .A(n982), .ZN(n700) );
  AOI22_X1 U127 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U128 ( .A(n981), .ZN(n699) );
  AOI22_X1 U129 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U130 ( .A(n980), .ZN(n698) );
  AOI22_X1 U131 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U132 ( .A(n951), .ZN(n673) );
  AOI22_X1 U133 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U134 ( .A(n948), .ZN(n671) );
  AOI22_X1 U135 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U136 ( .A(n947), .ZN(n670) );
  AOI22_X1 U137 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U138 ( .A(n946), .ZN(n669) );
  AOI22_X1 U139 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U140 ( .A(n945), .ZN(n668) );
  AOI22_X1 U141 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U142 ( .A(n944), .ZN(n667) );
  AOI22_X1 U143 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U144 ( .A(n943), .ZN(n666) );
  AOI22_X1 U145 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U146 ( .A(n915), .ZN(n641) );
  AOI22_X1 U147 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U148 ( .A(n913), .ZN(n640) );
  AOI22_X1 U149 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U150 ( .A(n912), .ZN(n639) );
  AOI22_X1 U151 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U152 ( .A(n911), .ZN(n638) );
  AOI22_X1 U153 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U154 ( .A(n910), .ZN(n637) );
  AOI22_X1 U155 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U156 ( .A(n909), .ZN(n636) );
  AOI22_X1 U157 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U158 ( .A(n908), .ZN(n635) );
  AOI22_X1 U159 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U160 ( .A(n907), .ZN(n634) );
  AOI22_X1 U161 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U162 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U163 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U164 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U165 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U166 ( .A(n985), .ZN(n703) );
  AOI22_X1 U167 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U168 ( .A(n949), .ZN(n672) );
  AOI22_X1 U169 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U170 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U171 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U172 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U173 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U174 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U175 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U176 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U177 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U178 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U179 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U180 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U181 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U182 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U183 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U184 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U185 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U186 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U187 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U188 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U189 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U190 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U191 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U192 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U193 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U194 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U195 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U196 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U197 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U198 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U199 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U200 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U201 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U202 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U203 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U204 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U205 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U206 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U207 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U208 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U209 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U210 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U211 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U212 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U213 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U214 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U215 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U216 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U217 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U218 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U219 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U220 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U221 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U222 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U223 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U224 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U225 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U226 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U227 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U228 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U229 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U230 ( .A(n999), .ZN(n715) );
  AOI22_X1 U231 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U232 ( .A(n998), .ZN(n714) );
  AOI22_X1 U233 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U234 ( .A(n979), .ZN(n697) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U236 ( .A(n977), .ZN(n696) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U238 ( .A(n976), .ZN(n695) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U240 ( .A(n975), .ZN(n694) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U242 ( .A(n974), .ZN(n693) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U244 ( .A(n973), .ZN(n692) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U246 ( .A(n972), .ZN(n691) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U248 ( .A(n971), .ZN(n690) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U250 ( .A(n970), .ZN(n689) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U252 ( .A(n968), .ZN(n688) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U254 ( .A(n967), .ZN(n687) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U256 ( .A(n966), .ZN(n686) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U258 ( .A(n965), .ZN(n685) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U260 ( .A(n964), .ZN(n684) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U262 ( .A(n963), .ZN(n683) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U264 ( .A(n962), .ZN(n682) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U266 ( .A(n942), .ZN(n665) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U268 ( .A(n940), .ZN(n664) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U270 ( .A(n939), .ZN(n663) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U272 ( .A(n938), .ZN(n662) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U274 ( .A(n937), .ZN(n661) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U276 ( .A(n936), .ZN(n660) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U278 ( .A(n935), .ZN(n659) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U280 ( .A(n934), .ZN(n658) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U282 ( .A(n933), .ZN(n657) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U284 ( .A(n931), .ZN(n656) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U286 ( .A(n930), .ZN(n655) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U288 ( .A(n929), .ZN(n654) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U290 ( .A(n928), .ZN(n653) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U292 ( .A(n927), .ZN(n652) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U294 ( .A(n926), .ZN(n651) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U296 ( .A(n925), .ZN(n650) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U298 ( .A(n906), .ZN(n633) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U300 ( .A(n904), .ZN(n632) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U302 ( .A(n903), .ZN(n631) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U304 ( .A(n902), .ZN(n630) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U306 ( .A(n901), .ZN(n629) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U308 ( .A(n900), .ZN(n628) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U310 ( .A(n899), .ZN(n627) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U312 ( .A(n898), .ZN(n626) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U314 ( .A(n897), .ZN(n625) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U316 ( .A(n895), .ZN(n624) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U318 ( .A(n894), .ZN(n623) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U320 ( .A(n893), .ZN(n622) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U322 ( .A(n892), .ZN(n621) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U324 ( .A(n891), .ZN(n620) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U326 ( .A(n890), .ZN(n619) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U328 ( .A(n889), .ZN(n618) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U330 ( .A(N12), .ZN(n253) );
  INV_X1 U331 ( .A(N11), .ZN(n252) );
  INV_X1 U332 ( .A(n997), .ZN(n713) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U334 ( .A(n995), .ZN(n712) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U336 ( .A(n994), .ZN(n711) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U338 ( .A(n993), .ZN(n710) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U340 ( .A(n992), .ZN(n709) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U342 ( .A(n991), .ZN(n708) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U344 ( .A(n990), .ZN(n707) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U346 ( .A(n989), .ZN(n706) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U348 ( .A(n924), .ZN(n649) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U350 ( .A(n922), .ZN(n648) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U352 ( .A(n921), .ZN(n647) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U354 ( .A(n920), .ZN(n646) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U356 ( .A(n919), .ZN(n645) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U358 ( .A(n918), .ZN(n644) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U360 ( .A(n917), .ZN(n643) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U362 ( .A(n916), .ZN(n642) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U364 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U366 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U368 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U370 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U372 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U374 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U376 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U378 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U380 ( .A(n961), .ZN(n681) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U382 ( .A(n959), .ZN(n680) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U384 ( .A(n958), .ZN(n679) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U386 ( .A(n957), .ZN(n678) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U388 ( .A(n956), .ZN(n677) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U390 ( .A(n955), .ZN(n676) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U392 ( .A(n954), .ZN(n675) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U394 ( .A(n953), .ZN(n674) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U396 ( .A(n888), .ZN(n617) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U398 ( .A(n886), .ZN(n616) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U400 ( .A(n885), .ZN(n615) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U402 ( .A(n884), .ZN(n614) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U404 ( .A(n883), .ZN(n613) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U406 ( .A(n882), .ZN(n612) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U408 ( .A(n881), .ZN(n611) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U410 ( .A(n880), .ZN(n610) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U412 ( .A(n879), .ZN(n609) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U414 ( .A(n877), .ZN(n608) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U416 ( .A(n876), .ZN(n607) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U418 ( .A(n875), .ZN(n606) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U420 ( .A(n874), .ZN(n605) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U422 ( .A(n873), .ZN(n604) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U424 ( .A(n872), .ZN(n603) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U426 ( .A(n871), .ZN(n602) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U428 ( .A(n870), .ZN(n601) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U430 ( .A(n868), .ZN(n600) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U432 ( .A(n867), .ZN(n599) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U434 ( .A(n866), .ZN(n598) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U436 ( .A(n865), .ZN(n597) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U438 ( .A(n864), .ZN(n596) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U440 ( .A(n863), .ZN(n595) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U442 ( .A(n862), .ZN(n594) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U444 ( .A(n861), .ZN(n293) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U446 ( .A(n859), .ZN(n292) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U448 ( .A(n858), .ZN(n291) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U450 ( .A(n857), .ZN(n290) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U452 ( .A(n856), .ZN(n289) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U454 ( .A(n855), .ZN(n288) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U456 ( .A(n854), .ZN(n287) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U458 ( .A(n853), .ZN(n286) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U460 ( .A(n852), .ZN(n285) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U462 ( .A(n850), .ZN(n284) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U464 ( .A(n849), .ZN(n283) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U466 ( .A(n848), .ZN(n282) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U468 ( .A(n847), .ZN(n281) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U470 ( .A(n846), .ZN(n280) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U472 ( .A(n845), .ZN(n279) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U474 ( .A(n844), .ZN(n278) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U476 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U477 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U478 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U479 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U480 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U481 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U482 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U483 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U484 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U485 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U486 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U487 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U488 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U489 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U490 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U491 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U492 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U494 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U496 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U498 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U500 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U502 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U504 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U506 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U508 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U510 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U512 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U514 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U516 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U518 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U520 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U522 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U524 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U526 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U528 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U530 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U532 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U534 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U536 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U538 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U540 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U542 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U544 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U546 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U548 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U550 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U552 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U554 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U556 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U558 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U560 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U562 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U564 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U566 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U568 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U570 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U572 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U574 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U576 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U578 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U580 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U582 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U584 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U586 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U588 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U590 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U592 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U594 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U596 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U598 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U600 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U602 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U604 ( .A(N13), .ZN(n842) );
  INV_X1 U605 ( .A(N14), .ZN(n843) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n249), .Z(n1) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n249), .Z(n2) );
  MUX2_X1 U608 ( .A(n2), .B(n1), .S(n242), .Z(n3) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n249), .Z(n4) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n249), .Z(n5) );
  MUX2_X1 U611 ( .A(n5), .B(n4), .S(n242), .Z(n6) );
  MUX2_X1 U612 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n249), .Z(n8) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n248), .Z(n9) );
  MUX2_X1 U615 ( .A(n9), .B(n8), .S(N11), .Z(n10) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n249), .Z(n11) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n248), .Z(n12) );
  MUX2_X1 U618 ( .A(n12), .B(n11), .S(n244), .Z(n13) );
  MUX2_X1 U619 ( .A(n13), .B(n10), .S(n241), .Z(n14) );
  MUX2_X1 U620 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n245), .Z(n16) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n245), .Z(n17) );
  MUX2_X1 U623 ( .A(n17), .B(n16), .S(n242), .Z(n18) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n245), .Z(n20) );
  MUX2_X1 U626 ( .A(n20), .B(n19), .S(n242), .Z(n21) );
  MUX2_X1 U627 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n245), .Z(n23) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n245), .Z(n24) );
  MUX2_X1 U630 ( .A(n24), .B(n23), .S(n242), .Z(n25) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n245), .Z(n26) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n245), .Z(n27) );
  MUX2_X1 U633 ( .A(n27), .B(n26), .S(n242), .Z(n28) );
  MUX2_X1 U634 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U635 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U636 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n245), .Z(n31) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n245), .Z(n32) );
  MUX2_X1 U639 ( .A(n32), .B(n31), .S(n242), .Z(n33) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U642 ( .A(n35), .B(n34), .S(n242), .Z(n36) );
  MUX2_X1 U643 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n246), .Z(n38) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n246), .Z(n39) );
  MUX2_X1 U646 ( .A(n39), .B(n38), .S(n242), .Z(n40) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n246), .Z(n41) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n246), .Z(n42) );
  MUX2_X1 U649 ( .A(n42), .B(n41), .S(n242), .Z(n43) );
  MUX2_X1 U650 ( .A(n43), .B(n40), .S(n241), .Z(n44) );
  MUX2_X1 U651 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n246), .Z(n46) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n246), .Z(n47) );
  MUX2_X1 U654 ( .A(n47), .B(n46), .S(n242), .Z(n48) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n246), .Z(n49) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n246), .Z(n50) );
  MUX2_X1 U657 ( .A(n50), .B(n49), .S(n242), .Z(n51) );
  MUX2_X1 U658 ( .A(n51), .B(n48), .S(n241), .Z(n52) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n246), .Z(n53) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n246), .Z(n54) );
  MUX2_X1 U661 ( .A(n54), .B(n53), .S(n242), .Z(n55) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n246), .Z(n56) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n246), .Z(n57) );
  MUX2_X1 U664 ( .A(n57), .B(n56), .S(n242), .Z(n58) );
  MUX2_X1 U665 ( .A(n58), .B(n55), .S(n241), .Z(n59) );
  MUX2_X1 U666 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U667 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n247), .Z(n61) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n247), .Z(n62) );
  MUX2_X1 U670 ( .A(n62), .B(n61), .S(n243), .Z(n63) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n247), .Z(n64) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n247), .Z(n65) );
  MUX2_X1 U673 ( .A(n65), .B(n64), .S(n243), .Z(n66) );
  MUX2_X1 U674 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n247), .Z(n68) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n247), .Z(n69) );
  MUX2_X1 U677 ( .A(n69), .B(n68), .S(n243), .Z(n70) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n247), .Z(n71) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n247), .Z(n72) );
  MUX2_X1 U680 ( .A(n72), .B(n71), .S(n243), .Z(n73) );
  MUX2_X1 U681 ( .A(n73), .B(n70), .S(N12), .Z(n74) );
  MUX2_X1 U682 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n247), .Z(n76) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n247), .Z(n77) );
  MUX2_X1 U685 ( .A(n77), .B(n76), .S(n243), .Z(n78) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n247), .Z(n79) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n247), .Z(n80) );
  MUX2_X1 U688 ( .A(n80), .B(n79), .S(n243), .Z(n81) );
  MUX2_X1 U689 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n245), .Z(n83) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n246), .Z(n84) );
  MUX2_X1 U692 ( .A(n84), .B(n83), .S(n243), .Z(n85) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n247), .Z(n86) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n245), .Z(n87) );
  MUX2_X1 U695 ( .A(n87), .B(n86), .S(n243), .Z(n88) );
  MUX2_X1 U696 ( .A(n88), .B(n85), .S(N12), .Z(n89) );
  MUX2_X1 U697 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U698 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n248), .Z(n91) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n245), .Z(n92) );
  MUX2_X1 U701 ( .A(n92), .B(n91), .S(n243), .Z(n93) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n247), .Z(n95) );
  MUX2_X1 U704 ( .A(n95), .B(n94), .S(n243), .Z(n96) );
  MUX2_X1 U705 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n98) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n248), .Z(n99) );
  MUX2_X1 U708 ( .A(n99), .B(n98), .S(n243), .Z(n100) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n246), .Z(n101) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n247), .Z(n102) );
  MUX2_X1 U711 ( .A(n102), .B(n101), .S(n243), .Z(n103) );
  MUX2_X1 U712 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U713 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n249), .Z(n106) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(N10), .Z(n107) );
  MUX2_X1 U716 ( .A(n107), .B(n106), .S(n244), .Z(n108) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n249), .Z(n109) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n250), .Z(n110) );
  MUX2_X1 U719 ( .A(n110), .B(n109), .S(n244), .Z(n111) );
  MUX2_X1 U720 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n249), .Z(n113) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n114) );
  MUX2_X1 U723 ( .A(n114), .B(n113), .S(n244), .Z(n115) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n249), .Z(n116) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n117) );
  MUX2_X1 U726 ( .A(n117), .B(n116), .S(n244), .Z(n118) );
  MUX2_X1 U727 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U728 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U729 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(N10), .Z(n121) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(N10), .Z(n122) );
  MUX2_X1 U732 ( .A(n122), .B(n121), .S(n244), .Z(n123) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(N10), .Z(n124) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n125) );
  MUX2_X1 U735 ( .A(n125), .B(n124), .S(n244), .Z(n126) );
  MUX2_X1 U736 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n248), .Z(n128) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n248), .Z(n129) );
  MUX2_X1 U739 ( .A(n129), .B(n128), .S(n244), .Z(n130) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n248), .Z(n131) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n248), .Z(n132) );
  MUX2_X1 U742 ( .A(n132), .B(n131), .S(n244), .Z(n133) );
  MUX2_X1 U743 ( .A(n133), .B(n130), .S(N12), .Z(n134) );
  MUX2_X1 U744 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n248), .Z(n136) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n248), .Z(n137) );
  MUX2_X1 U747 ( .A(n137), .B(n136), .S(n244), .Z(n138) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n248), .Z(n139) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n248), .Z(n140) );
  MUX2_X1 U750 ( .A(n140), .B(n139), .S(n244), .Z(n141) );
  MUX2_X1 U751 ( .A(n141), .B(n138), .S(N12), .Z(n142) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n248), .Z(n143) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n248), .Z(n144) );
  MUX2_X1 U754 ( .A(n144), .B(n143), .S(n244), .Z(n145) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n248), .Z(n146) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n248), .Z(n147) );
  MUX2_X1 U757 ( .A(n147), .B(n146), .S(n244), .Z(n148) );
  MUX2_X1 U758 ( .A(n148), .B(n145), .S(N12), .Z(n149) );
  MUX2_X1 U759 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U760 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n249), .Z(n151) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n249), .Z(n152) );
  MUX2_X1 U763 ( .A(n152), .B(n151), .S(n242), .Z(n153) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n249), .Z(n154) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n249), .Z(n155) );
  MUX2_X1 U766 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U767 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n249), .Z(n158) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n249), .Z(n159) );
  MUX2_X1 U770 ( .A(n159), .B(n158), .S(N11), .Z(n160) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n249), .Z(n161) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n249), .Z(n162) );
  MUX2_X1 U773 ( .A(n162), .B(n161), .S(n242), .Z(n163) );
  MUX2_X1 U774 ( .A(n163), .B(n160), .S(n241), .Z(n164) );
  MUX2_X1 U775 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n249), .Z(n166) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n249), .Z(n167) );
  MUX2_X1 U778 ( .A(n167), .B(n166), .S(N11), .Z(n168) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n249), .Z(n169) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n249), .Z(n170) );
  MUX2_X1 U781 ( .A(n170), .B(n169), .S(n243), .Z(n171) );
  MUX2_X1 U782 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n245), .Z(n173) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n250), .Z(n174) );
  MUX2_X1 U785 ( .A(n174), .B(n173), .S(N11), .Z(n175) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n250), .Z(n176) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n250), .Z(n177) );
  MUX2_X1 U788 ( .A(n177), .B(n176), .S(n243), .Z(n178) );
  MUX2_X1 U789 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U790 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U791 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n245), .Z(n181) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n247), .Z(n182) );
  MUX2_X1 U794 ( .A(n182), .B(n181), .S(N11), .Z(n183) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n250), .Z(n184) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n250), .Z(n185) );
  MUX2_X1 U797 ( .A(n185), .B(n184), .S(N11), .Z(n186) );
  MUX2_X1 U798 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n246), .Z(n188) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n250), .Z(n189) );
  MUX2_X1 U801 ( .A(n189), .B(n188), .S(N11), .Z(n190) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n248), .Z(n191) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n250), .Z(n192) );
  MUX2_X1 U804 ( .A(n192), .B(n191), .S(n244), .Z(n193) );
  MUX2_X1 U805 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U806 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n247), .Z(n196) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n250), .Z(n197) );
  MUX2_X1 U809 ( .A(n197), .B(n196), .S(n242), .Z(n198) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n250), .Z(n199) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n250), .Z(n200) );
  MUX2_X1 U812 ( .A(n200), .B(n199), .S(n244), .Z(n201) );
  MUX2_X1 U813 ( .A(n201), .B(n198), .S(n241), .Z(n202) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n250), .Z(n203) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n250), .Z(n204) );
  MUX2_X1 U816 ( .A(n204), .B(n203), .S(n244), .Z(n205) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n250), .Z(n206) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n250), .Z(n207) );
  MUX2_X1 U819 ( .A(n207), .B(n206), .S(N11), .Z(n208) );
  MUX2_X1 U820 ( .A(n208), .B(n205), .S(n241), .Z(n209) );
  MUX2_X1 U821 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U822 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n246), .Z(n211) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n246), .Z(n212) );
  MUX2_X1 U825 ( .A(n212), .B(n211), .S(n243), .Z(n213) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n249), .Z(n214) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n250), .Z(n215) );
  MUX2_X1 U828 ( .A(n215), .B(n214), .S(n244), .Z(n216) );
  MUX2_X1 U829 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n245), .Z(n218) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(N10), .Z(n219) );
  MUX2_X1 U832 ( .A(n219), .B(n218), .S(n243), .Z(n220) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n250), .Z(n221) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n222) );
  MUX2_X1 U835 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U836 ( .A(n223), .B(n220), .S(n241), .Z(n224) );
  MUX2_X1 U837 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n250), .Z(n226) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n227) );
  MUX2_X1 U840 ( .A(n227), .B(n226), .S(N11), .Z(n228) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n246), .Z(n229) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n230) );
  MUX2_X1 U843 ( .A(n230), .B(n229), .S(N11), .Z(n231) );
  MUX2_X1 U844 ( .A(n231), .B(n228), .S(N12), .Z(n232) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n247), .Z(n233) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n234) );
  MUX2_X1 U847 ( .A(n234), .B(n233), .S(n243), .Z(n235) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n236) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n237) );
  MUX2_X1 U850 ( .A(n237), .B(n236), .S(N11), .Z(n238) );
  MUX2_X1 U851 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U852 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U853 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_4 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  BUF_X1 U3 ( .A(N10), .Z(n249) );
  BUF_X1 U4 ( .A(n250), .Z(n246) );
  BUF_X1 U5 ( .A(n250), .Z(n245) );
  BUF_X1 U6 ( .A(n250), .Z(n247) );
  BUF_X1 U7 ( .A(n250), .Z(n248) );
  BUF_X1 U8 ( .A(N10), .Z(n250) );
  INV_X1 U9 ( .A(n1111), .ZN(n841) );
  INV_X1 U10 ( .A(n1100), .ZN(n840) );
  INV_X1 U11 ( .A(n1090), .ZN(n839) );
  INV_X1 U12 ( .A(n1080), .ZN(n838) );
  INV_X1 U13 ( .A(n1070), .ZN(n837) );
  INV_X1 U14 ( .A(n1060), .ZN(n836) );
  INV_X1 U15 ( .A(n1051), .ZN(n835) );
  INV_X1 U16 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U19 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U20 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U21 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U22 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U23 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U24 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U26 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U27 ( .A(n1131), .ZN(n816) );
  INV_X1 U28 ( .A(n1121), .ZN(n815) );
  INV_X1 U29 ( .A(n887), .ZN(n814) );
  INV_X1 U30 ( .A(n878), .ZN(n813) );
  INV_X1 U31 ( .A(n869), .ZN(n812) );
  INV_X1 U32 ( .A(n860), .ZN(n811) );
  INV_X1 U33 ( .A(n851), .ZN(n810) );
  INV_X1 U34 ( .A(n987), .ZN(n828) );
  INV_X1 U35 ( .A(n978), .ZN(n827) );
  INV_X1 U36 ( .A(n969), .ZN(n826) );
  INV_X1 U37 ( .A(n914), .ZN(n820) );
  INV_X1 U38 ( .A(n905), .ZN(n819) );
  INV_X1 U39 ( .A(n896), .ZN(n818) );
  INV_X1 U40 ( .A(n1033), .ZN(n833) );
  INV_X1 U41 ( .A(n1023), .ZN(n832) );
  INV_X1 U42 ( .A(n1014), .ZN(n831) );
  INV_X1 U43 ( .A(n1005), .ZN(n830) );
  INV_X1 U44 ( .A(n996), .ZN(n829) );
  INV_X1 U45 ( .A(n960), .ZN(n825) );
  INV_X1 U46 ( .A(n950), .ZN(n824) );
  INV_X1 U47 ( .A(n941), .ZN(n823) );
  INV_X1 U48 ( .A(n932), .ZN(n822) );
  INV_X1 U49 ( .A(n923), .ZN(n821) );
  INV_X1 U50 ( .A(n1142), .ZN(n817) );
  BUF_X1 U51 ( .A(N11), .Z(n242) );
  BUF_X1 U52 ( .A(N11), .Z(n243) );
  BUF_X1 U53 ( .A(N11), .Z(n244) );
  INV_X1 U54 ( .A(N10), .ZN(n251) );
  BUF_X1 U55 ( .A(N12), .Z(n241) );
  NOR3_X1 U56 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U57 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U58 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U60 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U62 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U63 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U64 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U65 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U67 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U69 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U70 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U71 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U72 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U73 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U74 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U75 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U76 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U77 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U79 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U81 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U82 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U83 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U84 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U85 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U86 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U88 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U89 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U90 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U92 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U94 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U95 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U96 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U97 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U98 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U99 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U100 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U101 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U102 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U103 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U104 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U105 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U106 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U107 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U108 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U109 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U110 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U111 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U112 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U113 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U114 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U115 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U116 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U117 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U118 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U119 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U120 ( .A(n988), .ZN(n705) );
  AOI22_X1 U121 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U122 ( .A(n981), .ZN(n699) );
  AOI22_X1 U123 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U124 ( .A(n980), .ZN(n698) );
  AOI22_X1 U125 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U126 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U127 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U128 ( .A(n986), .ZN(n704) );
  AOI22_X1 U129 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U130 ( .A(n985), .ZN(n703) );
  AOI22_X1 U131 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U132 ( .A(n984), .ZN(n702) );
  AOI22_X1 U133 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U134 ( .A(n983), .ZN(n701) );
  AOI22_X1 U135 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U136 ( .A(n982), .ZN(n700) );
  AOI22_X1 U137 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U138 ( .A(n951), .ZN(n673) );
  AOI22_X1 U139 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U140 ( .A(n948), .ZN(n671) );
  AOI22_X1 U141 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U142 ( .A(n947), .ZN(n670) );
  AOI22_X1 U143 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U144 ( .A(n946), .ZN(n669) );
  AOI22_X1 U145 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U146 ( .A(n945), .ZN(n668) );
  AOI22_X1 U147 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U148 ( .A(n944), .ZN(n667) );
  AOI22_X1 U149 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U150 ( .A(n943), .ZN(n666) );
  AOI22_X1 U151 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U152 ( .A(n915), .ZN(n641) );
  AOI22_X1 U153 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U154 ( .A(n913), .ZN(n640) );
  AOI22_X1 U155 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U156 ( .A(n911), .ZN(n638) );
  AOI22_X1 U157 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U158 ( .A(n910), .ZN(n637) );
  AOI22_X1 U159 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U160 ( .A(n909), .ZN(n636) );
  AOI22_X1 U161 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U162 ( .A(n908), .ZN(n635) );
  AOI22_X1 U163 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U164 ( .A(n907), .ZN(n634) );
  AOI22_X1 U165 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U166 ( .A(n949), .ZN(n672) );
  AOI22_X1 U167 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U168 ( .A(n912), .ZN(n639) );
  AOI22_X1 U169 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U170 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U171 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U172 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U173 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U174 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U175 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U176 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U177 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U178 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U179 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U180 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U181 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U182 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U183 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U184 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U185 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U186 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U187 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U188 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U189 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U190 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U191 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U192 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U193 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U194 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U195 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U196 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U197 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U198 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U199 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U200 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U201 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U202 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U203 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U204 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U205 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U206 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U207 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U208 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U209 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U210 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U211 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U212 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U213 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U214 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U215 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U216 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U217 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U218 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U219 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U220 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U221 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U222 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U223 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U224 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U225 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U226 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U227 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U228 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U229 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U230 ( .A(n999), .ZN(n715) );
  AOI22_X1 U231 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U232 ( .A(n998), .ZN(n714) );
  AOI22_X1 U233 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U234 ( .A(n979), .ZN(n697) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U236 ( .A(n977), .ZN(n696) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U238 ( .A(n976), .ZN(n695) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U240 ( .A(n975), .ZN(n694) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U242 ( .A(n974), .ZN(n693) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U244 ( .A(n973), .ZN(n692) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U246 ( .A(n972), .ZN(n691) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U248 ( .A(n971), .ZN(n690) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U250 ( .A(n970), .ZN(n689) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U252 ( .A(n968), .ZN(n688) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U254 ( .A(n967), .ZN(n687) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U256 ( .A(n966), .ZN(n686) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U258 ( .A(n965), .ZN(n685) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U260 ( .A(n964), .ZN(n684) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U262 ( .A(n963), .ZN(n683) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U264 ( .A(n962), .ZN(n682) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U266 ( .A(n942), .ZN(n665) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U268 ( .A(n940), .ZN(n664) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U270 ( .A(n939), .ZN(n663) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U272 ( .A(n938), .ZN(n662) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U274 ( .A(n937), .ZN(n661) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U276 ( .A(n936), .ZN(n660) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U278 ( .A(n935), .ZN(n659) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U280 ( .A(n934), .ZN(n658) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U282 ( .A(n933), .ZN(n657) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U284 ( .A(n931), .ZN(n656) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U286 ( .A(n930), .ZN(n655) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U288 ( .A(n929), .ZN(n654) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U290 ( .A(n928), .ZN(n653) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U292 ( .A(n927), .ZN(n652) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U294 ( .A(n926), .ZN(n651) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U296 ( .A(n925), .ZN(n650) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U298 ( .A(n906), .ZN(n633) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U300 ( .A(n904), .ZN(n632) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U302 ( .A(n903), .ZN(n631) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U304 ( .A(n902), .ZN(n630) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U306 ( .A(n901), .ZN(n629) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U308 ( .A(n900), .ZN(n628) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U310 ( .A(n899), .ZN(n627) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U312 ( .A(n898), .ZN(n626) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U314 ( .A(n897), .ZN(n625) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U316 ( .A(n895), .ZN(n624) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U318 ( .A(n894), .ZN(n623) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U320 ( .A(n893), .ZN(n622) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U322 ( .A(n892), .ZN(n621) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U324 ( .A(n891), .ZN(n620) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U326 ( .A(n890), .ZN(n619) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U328 ( .A(n889), .ZN(n618) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U330 ( .A(N12), .ZN(n253) );
  INV_X1 U331 ( .A(N11), .ZN(n252) );
  INV_X1 U332 ( .A(n997), .ZN(n713) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U334 ( .A(n995), .ZN(n712) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U336 ( .A(n994), .ZN(n711) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U338 ( .A(n993), .ZN(n710) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U340 ( .A(n992), .ZN(n709) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U342 ( .A(n991), .ZN(n708) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U344 ( .A(n990), .ZN(n707) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U346 ( .A(n989), .ZN(n706) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U348 ( .A(n924), .ZN(n649) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U350 ( .A(n922), .ZN(n648) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U352 ( .A(n921), .ZN(n647) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U354 ( .A(n920), .ZN(n646) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U356 ( .A(n919), .ZN(n645) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U358 ( .A(n918), .ZN(n644) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U360 ( .A(n917), .ZN(n643) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U362 ( .A(n916), .ZN(n642) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U364 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U366 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U368 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U370 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U372 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U374 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U376 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U378 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U380 ( .A(n961), .ZN(n681) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U382 ( .A(n959), .ZN(n680) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U384 ( .A(n958), .ZN(n679) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U386 ( .A(n957), .ZN(n678) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U388 ( .A(n956), .ZN(n677) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U390 ( .A(n955), .ZN(n676) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U392 ( .A(n954), .ZN(n675) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U394 ( .A(n953), .ZN(n674) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U396 ( .A(n888), .ZN(n617) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U398 ( .A(n886), .ZN(n616) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U400 ( .A(n885), .ZN(n615) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U402 ( .A(n884), .ZN(n614) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U404 ( .A(n883), .ZN(n613) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U406 ( .A(n882), .ZN(n612) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U408 ( .A(n881), .ZN(n611) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U410 ( .A(n880), .ZN(n610) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U412 ( .A(n879), .ZN(n609) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U414 ( .A(n877), .ZN(n608) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U416 ( .A(n876), .ZN(n607) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U418 ( .A(n875), .ZN(n606) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U420 ( .A(n874), .ZN(n605) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U422 ( .A(n873), .ZN(n604) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U424 ( .A(n872), .ZN(n603) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U426 ( .A(n871), .ZN(n602) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U428 ( .A(n870), .ZN(n601) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U430 ( .A(n868), .ZN(n600) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U432 ( .A(n867), .ZN(n599) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U434 ( .A(n866), .ZN(n598) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U436 ( .A(n865), .ZN(n597) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U438 ( .A(n864), .ZN(n596) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U440 ( .A(n863), .ZN(n595) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U442 ( .A(n862), .ZN(n594) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U444 ( .A(n861), .ZN(n293) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U446 ( .A(n859), .ZN(n292) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U448 ( .A(n858), .ZN(n291) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U450 ( .A(n857), .ZN(n290) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U452 ( .A(n856), .ZN(n289) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U454 ( .A(n855), .ZN(n288) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U456 ( .A(n854), .ZN(n287) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U458 ( .A(n853), .ZN(n286) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U460 ( .A(n852), .ZN(n285) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U462 ( .A(n850), .ZN(n284) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U464 ( .A(n849), .ZN(n283) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U466 ( .A(n848), .ZN(n282) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U468 ( .A(n847), .ZN(n281) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U470 ( .A(n846), .ZN(n280) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U472 ( .A(n845), .ZN(n279) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U474 ( .A(n844), .ZN(n278) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U476 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U477 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U478 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U479 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U480 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U481 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U482 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U483 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U484 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U485 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U486 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U487 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U488 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U489 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U490 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U491 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U492 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U494 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U496 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U498 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U500 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U502 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U504 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U506 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U508 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U510 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U512 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U514 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U516 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U518 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U520 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U522 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U524 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U526 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U528 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U530 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U532 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U534 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U536 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U538 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U540 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U542 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U544 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U546 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U548 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U550 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U552 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U554 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U556 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U558 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U560 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U562 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U564 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U566 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U568 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U570 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U572 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U574 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U576 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U578 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U580 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U582 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U584 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U586 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U588 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U590 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U592 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U594 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U596 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U598 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U600 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U602 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U604 ( .A(N13), .ZN(n842) );
  INV_X1 U605 ( .A(N14), .ZN(n843) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n249), .Z(n1) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n249), .Z(n2) );
  MUX2_X1 U608 ( .A(n2), .B(n1), .S(n242), .Z(n3) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n249), .Z(n4) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n246), .Z(n5) );
  MUX2_X1 U611 ( .A(n5), .B(n4), .S(n242), .Z(n6) );
  MUX2_X1 U612 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n249), .Z(n8) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n245), .Z(n9) );
  MUX2_X1 U615 ( .A(n9), .B(n8), .S(N11), .Z(n10) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n245), .Z(n11) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n247), .Z(n12) );
  MUX2_X1 U618 ( .A(n12), .B(n11), .S(n244), .Z(n13) );
  MUX2_X1 U619 ( .A(n13), .B(n10), .S(N12), .Z(n14) );
  MUX2_X1 U620 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n245), .Z(n16) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n245), .Z(n17) );
  MUX2_X1 U623 ( .A(n17), .B(n16), .S(n242), .Z(n18) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n245), .Z(n20) );
  MUX2_X1 U626 ( .A(n20), .B(n19), .S(n242), .Z(n21) );
  MUX2_X1 U627 ( .A(n21), .B(n18), .S(N12), .Z(n22) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n245), .Z(n23) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n245), .Z(n24) );
  MUX2_X1 U630 ( .A(n24), .B(n23), .S(n242), .Z(n25) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n245), .Z(n26) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n245), .Z(n27) );
  MUX2_X1 U633 ( .A(n27), .B(n26), .S(n242), .Z(n28) );
  MUX2_X1 U634 ( .A(n28), .B(n25), .S(N12), .Z(n29) );
  MUX2_X1 U635 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U636 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n245), .Z(n31) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n245), .Z(n32) );
  MUX2_X1 U639 ( .A(n32), .B(n31), .S(n242), .Z(n33) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U642 ( .A(n35), .B(n34), .S(n242), .Z(n36) );
  MUX2_X1 U643 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n246), .Z(n38) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n246), .Z(n39) );
  MUX2_X1 U646 ( .A(n39), .B(n38), .S(n242), .Z(n40) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n246), .Z(n41) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n246), .Z(n42) );
  MUX2_X1 U649 ( .A(n42), .B(n41), .S(n242), .Z(n43) );
  MUX2_X1 U650 ( .A(n43), .B(n40), .S(n241), .Z(n44) );
  MUX2_X1 U651 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n246), .Z(n46) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n246), .Z(n47) );
  MUX2_X1 U654 ( .A(n47), .B(n46), .S(n242), .Z(n48) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n246), .Z(n49) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n246), .Z(n50) );
  MUX2_X1 U657 ( .A(n50), .B(n49), .S(n242), .Z(n51) );
  MUX2_X1 U658 ( .A(n51), .B(n48), .S(n241), .Z(n52) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n246), .Z(n53) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n246), .Z(n54) );
  MUX2_X1 U661 ( .A(n54), .B(n53), .S(n242), .Z(n55) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n246), .Z(n56) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n246), .Z(n57) );
  MUX2_X1 U664 ( .A(n57), .B(n56), .S(n242), .Z(n58) );
  MUX2_X1 U665 ( .A(n58), .B(n55), .S(n241), .Z(n59) );
  MUX2_X1 U666 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U667 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n247), .Z(n61) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n247), .Z(n62) );
  MUX2_X1 U670 ( .A(n62), .B(n61), .S(n243), .Z(n63) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n247), .Z(n64) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n247), .Z(n65) );
  MUX2_X1 U673 ( .A(n65), .B(n64), .S(n243), .Z(n66) );
  MUX2_X1 U674 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n247), .Z(n68) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n247), .Z(n69) );
  MUX2_X1 U677 ( .A(n69), .B(n68), .S(n243), .Z(n70) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n247), .Z(n71) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n247), .Z(n72) );
  MUX2_X1 U680 ( .A(n72), .B(n71), .S(n243), .Z(n73) );
  MUX2_X1 U681 ( .A(n73), .B(n70), .S(n241), .Z(n74) );
  MUX2_X1 U682 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n247), .Z(n76) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n247), .Z(n77) );
  MUX2_X1 U685 ( .A(n77), .B(n76), .S(n243), .Z(n78) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n247), .Z(n79) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n247), .Z(n80) );
  MUX2_X1 U688 ( .A(n80), .B(n79), .S(n243), .Z(n81) );
  MUX2_X1 U689 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n248), .Z(n83) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n248), .Z(n84) );
  MUX2_X1 U692 ( .A(n84), .B(n83), .S(n243), .Z(n85) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n248), .Z(n86) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n248), .Z(n87) );
  MUX2_X1 U695 ( .A(n87), .B(n86), .S(n243), .Z(n88) );
  MUX2_X1 U696 ( .A(n88), .B(n85), .S(n241), .Z(n89) );
  MUX2_X1 U697 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U698 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n248), .Z(n91) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n248), .Z(n92) );
  MUX2_X1 U701 ( .A(n92), .B(n91), .S(n243), .Z(n93) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n248), .Z(n94) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n248), .Z(n95) );
  MUX2_X1 U704 ( .A(n95), .B(n94), .S(n243), .Z(n96) );
  MUX2_X1 U705 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n248), .Z(n98) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n248), .Z(n99) );
  MUX2_X1 U708 ( .A(n99), .B(n98), .S(n243), .Z(n100) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n248), .Z(n101) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n248), .Z(n102) );
  MUX2_X1 U711 ( .A(n102), .B(n101), .S(n243), .Z(n103) );
  MUX2_X1 U712 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U713 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n249), .Z(n106) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n247), .Z(n107) );
  MUX2_X1 U716 ( .A(n107), .B(n106), .S(n244), .Z(n108) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n250), .Z(n109) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n248), .Z(n110) );
  MUX2_X1 U719 ( .A(n110), .B(n109), .S(n244), .Z(n111) );
  MUX2_X1 U720 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n245), .Z(n113) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n250), .Z(n114) );
  MUX2_X1 U723 ( .A(n114), .B(n113), .S(n244), .Z(n115) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n246), .Z(n116) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n117) );
  MUX2_X1 U726 ( .A(n117), .B(n116), .S(n244), .Z(n118) );
  MUX2_X1 U727 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U728 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U729 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(N10), .Z(n121) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(N10), .Z(n122) );
  MUX2_X1 U732 ( .A(n122), .B(n121), .S(n244), .Z(n123) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(N10), .Z(n124) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n125) );
  MUX2_X1 U735 ( .A(n125), .B(n124), .S(n244), .Z(n126) );
  MUX2_X1 U736 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n249), .Z(n128) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n250), .Z(n129) );
  MUX2_X1 U739 ( .A(n129), .B(n128), .S(n244), .Z(n130) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n249), .Z(n131) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(N10), .Z(n132) );
  MUX2_X1 U742 ( .A(n132), .B(n131), .S(n244), .Z(n133) );
  MUX2_X1 U743 ( .A(n133), .B(n130), .S(n241), .Z(n134) );
  MUX2_X1 U744 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n249), .Z(n136) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n250), .Z(n137) );
  MUX2_X1 U747 ( .A(n137), .B(n136), .S(n244), .Z(n138) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n249), .Z(n139) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(N10), .Z(n140) );
  MUX2_X1 U750 ( .A(n140), .B(n139), .S(n244), .Z(n141) );
  MUX2_X1 U751 ( .A(n141), .B(n138), .S(n241), .Z(n142) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(N10), .Z(n143) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(N10), .Z(n144) );
  MUX2_X1 U754 ( .A(n144), .B(n143), .S(n244), .Z(n145) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(N10), .Z(n146) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(N10), .Z(n147) );
  MUX2_X1 U757 ( .A(n147), .B(n146), .S(n244), .Z(n148) );
  MUX2_X1 U758 ( .A(n148), .B(n145), .S(n241), .Z(n149) );
  MUX2_X1 U759 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U760 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n249), .Z(n151) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n249), .Z(n152) );
  MUX2_X1 U763 ( .A(n152), .B(n151), .S(n242), .Z(n153) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n249), .Z(n154) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n249), .Z(n155) );
  MUX2_X1 U766 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U767 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n249), .Z(n158) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n249), .Z(n159) );
  MUX2_X1 U770 ( .A(n159), .B(n158), .S(N11), .Z(n160) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n249), .Z(n161) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n249), .Z(n162) );
  MUX2_X1 U773 ( .A(n162), .B(n161), .S(n242), .Z(n163) );
  MUX2_X1 U774 ( .A(n163), .B(n160), .S(N12), .Z(n164) );
  MUX2_X1 U775 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n249), .Z(n166) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n249), .Z(n167) );
  MUX2_X1 U778 ( .A(n167), .B(n166), .S(N11), .Z(n168) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n249), .Z(n169) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n249), .Z(n170) );
  MUX2_X1 U781 ( .A(n170), .B(n169), .S(n243), .Z(n171) );
  MUX2_X1 U782 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n246), .Z(n173) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n250), .Z(n174) );
  MUX2_X1 U785 ( .A(n174), .B(n173), .S(N11), .Z(n175) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n250), .Z(n176) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n250), .Z(n177) );
  MUX2_X1 U788 ( .A(n177), .B(n176), .S(n243), .Z(n178) );
  MUX2_X1 U789 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U790 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U791 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n250), .Z(n181) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n248), .Z(n182) );
  MUX2_X1 U794 ( .A(n182), .B(n181), .S(N11), .Z(n183) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n249), .Z(n184) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n245), .Z(n185) );
  MUX2_X1 U797 ( .A(n185), .B(n184), .S(N11), .Z(n186) );
  MUX2_X1 U798 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n250), .Z(n188) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n250), .Z(n189) );
  MUX2_X1 U801 ( .A(n189), .B(n188), .S(N11), .Z(n190) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n247), .Z(n191) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n246), .Z(n192) );
  MUX2_X1 U804 ( .A(n192), .B(n191), .S(n244), .Z(n193) );
  MUX2_X1 U805 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U806 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n246), .Z(n196) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n250), .Z(n197) );
  MUX2_X1 U809 ( .A(n197), .B(n196), .S(n242), .Z(n198) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n245), .Z(n199) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n248), .Z(n200) );
  MUX2_X1 U812 ( .A(n200), .B(n199), .S(n244), .Z(n201) );
  MUX2_X1 U813 ( .A(n201), .B(n198), .S(n241), .Z(n202) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n250), .Z(n203) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n247), .Z(n204) );
  MUX2_X1 U816 ( .A(n204), .B(n203), .S(n244), .Z(n205) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n246), .Z(n206) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n245), .Z(n207) );
  MUX2_X1 U819 ( .A(n207), .B(n206), .S(N11), .Z(n208) );
  MUX2_X1 U820 ( .A(n208), .B(n205), .S(N12), .Z(n209) );
  MUX2_X1 U821 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U822 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n250), .Z(n211) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n247), .Z(n212) );
  MUX2_X1 U825 ( .A(n212), .B(n211), .S(n243), .Z(n213) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n248), .Z(n214) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n250), .Z(n215) );
  MUX2_X1 U828 ( .A(n215), .B(n214), .S(n244), .Z(n216) );
  MUX2_X1 U829 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n250), .Z(n218) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n250), .Z(n219) );
  MUX2_X1 U832 ( .A(n219), .B(n218), .S(n243), .Z(n220) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(N10), .Z(n221) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n247), .Z(n222) );
  MUX2_X1 U835 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U836 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U837 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n250), .Z(n226) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(N10), .Z(n227) );
  MUX2_X1 U840 ( .A(n227), .B(n226), .S(N11), .Z(n228) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n249), .Z(n229) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n248), .Z(n230) );
  MUX2_X1 U843 ( .A(n230), .B(n229), .S(N11), .Z(n231) );
  MUX2_X1 U844 ( .A(n231), .B(n228), .S(n241), .Z(n232) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n233) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n250), .Z(n234) );
  MUX2_X1 U847 ( .A(n234), .B(n233), .S(n243), .Z(n235) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n250), .Z(n236) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n250), .Z(n237) );
  MUX2_X1 U850 ( .A(n237), .B(n236), .S(N11), .Z(n238) );
  MUX2_X1 U851 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U852 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U853 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_3 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n256), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n257), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n258), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n259), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n260), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n261), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n262), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n263), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n264), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n265), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n266), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n267), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n268), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n269), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n270), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n271), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n272), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n273), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n274), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n275), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n276), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n277), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n278), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n279), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n280), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n281), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n282), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n283), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n284), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n285), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n286), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n287), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n288), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n289), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n290), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n291), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n292), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n293), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n594), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n595), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n596), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n597), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n598), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n599), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n600), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n601), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n602), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n603), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n604), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n605), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n606), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n607), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n608), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n609), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n610), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n611), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n612), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n613), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n614), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n615), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n616), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n617), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n618), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n619), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n620), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n621), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n622), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n623), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n624), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n625), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n626), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n627), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n628), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n629), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n630), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n631), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n632), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n633), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n634), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n635), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n636), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n637), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n638), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n639), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n640), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n641), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n642), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n643), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n644), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n645), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n646), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n647), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n648), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n649), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n650), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n651), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n652), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n653), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n654), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n655), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n656), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n657), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n658), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n659), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n660), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n661), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n662), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n663), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n664), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n665), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n666), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n667), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n668), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n669), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n670), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n671), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n672), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n673), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n674), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n675), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n676), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n677), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n678), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n679), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n680), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n681), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n682), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n683), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n684), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n685), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n686), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n687), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n688), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n689), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n690), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n691), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n692), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n693), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n694), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n695), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n696), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n697), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n698), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n699), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n700), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n701), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n702), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n703), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n704), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n705), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n706), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n707), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n708), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n709), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n710), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n711), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n712), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n713), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n714), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n715), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n716), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n717), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n718), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n719), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n720), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n721), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n722), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n723), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n724), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n725), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n726), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n727), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n728), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n729), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n730), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n731), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n732), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n733), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n734), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n735), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n736), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n737), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n738), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n739), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n740), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n741), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n742), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n743), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n744), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n745), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n746), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n747), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n748), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n749), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n750), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n751), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n752), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n753), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n754), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n755), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n756), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n757), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n758), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n759), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n760), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n761), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n762), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n763), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n764), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n765), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n766), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n767), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n768), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n769), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n770), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n771), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n772), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n773), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n774), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n775), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n776), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n777), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n778), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n779), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n780), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n781), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n782), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n783), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n784), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n785), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n786), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n787), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n788), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n789), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n790), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n791), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n792), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n793), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n794), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n795), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n796), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n797), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n798), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n799), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n800), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n801), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n802), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n803), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n804), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n805), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n806), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n807), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n808), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n809), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n810), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n811), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X2 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .QN(n1) );
  DFF_X2 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  INV_X2 U3 ( .A(n1), .ZN(data_out[3]) );
  BUF_X1 U4 ( .A(n252), .Z(n250) );
  BUF_X1 U5 ( .A(N10), .Z(n251) );
  BUF_X1 U6 ( .A(n252), .Z(n248) );
  BUF_X1 U7 ( .A(n252), .Z(n247) );
  BUF_X1 U8 ( .A(n252), .Z(n249) );
  BUF_X1 U9 ( .A(N10), .Z(n252) );
  INV_X1 U10 ( .A(n1113), .ZN(n843) );
  INV_X1 U11 ( .A(n1102), .ZN(n842) );
  INV_X1 U12 ( .A(n1092), .ZN(n841) );
  INV_X1 U13 ( .A(n1082), .ZN(n840) );
  INV_X1 U14 ( .A(n1072), .ZN(n839) );
  INV_X1 U15 ( .A(n1062), .ZN(n838) );
  INV_X1 U16 ( .A(n1053), .ZN(n837) );
  INV_X1 U17 ( .A(n1044), .ZN(n836) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1105) );
  NOR3_X1 U19 ( .A1(N11), .A2(N12), .A3(n253), .ZN(n1094) );
  NAND2_X1 U20 ( .A1(n1104), .A2(n1136), .ZN(n1062) );
  NAND2_X1 U21 ( .A1(n1105), .A2(n1104), .ZN(n1113) );
  NAND2_X1 U22 ( .A1(n1094), .A2(n1104), .ZN(n1102) );
  NAND2_X1 U23 ( .A1(n1084), .A2(n1104), .ZN(n1092) );
  NAND2_X1 U24 ( .A1(n1074), .A2(n1104), .ZN(n1082) );
  NAND2_X1 U25 ( .A1(n1064), .A2(n1104), .ZN(n1072) );
  NAND2_X1 U26 ( .A1(n1104), .A2(n1125), .ZN(n1053) );
  NAND2_X1 U27 ( .A1(n1104), .A2(n1115), .ZN(n1044) );
  INV_X1 U28 ( .A(n1133), .ZN(n818) );
  INV_X1 U29 ( .A(n1123), .ZN(n817) );
  INV_X1 U30 ( .A(n889), .ZN(n816) );
  INV_X1 U31 ( .A(n880), .ZN(n815) );
  INV_X1 U32 ( .A(n871), .ZN(n814) );
  INV_X1 U33 ( .A(n862), .ZN(n813) );
  INV_X1 U34 ( .A(n853), .ZN(n812) );
  INV_X1 U35 ( .A(n989), .ZN(n830) );
  INV_X1 U36 ( .A(n980), .ZN(n829) );
  INV_X1 U37 ( .A(n971), .ZN(n828) );
  INV_X1 U38 ( .A(n916), .ZN(n822) );
  INV_X1 U39 ( .A(n907), .ZN(n821) );
  INV_X1 U40 ( .A(n898), .ZN(n820) );
  INV_X1 U41 ( .A(n1035), .ZN(n835) );
  INV_X1 U42 ( .A(n1025), .ZN(n834) );
  INV_X1 U43 ( .A(n1016), .ZN(n833) );
  INV_X1 U44 ( .A(n1007), .ZN(n832) );
  INV_X1 U45 ( .A(n998), .ZN(n831) );
  INV_X1 U46 ( .A(n962), .ZN(n827) );
  INV_X1 U47 ( .A(n952), .ZN(n826) );
  INV_X1 U48 ( .A(n943), .ZN(n825) );
  INV_X1 U49 ( .A(n934), .ZN(n824) );
  INV_X1 U50 ( .A(n925), .ZN(n823) );
  INV_X1 U51 ( .A(n1144), .ZN(n819) );
  BUF_X1 U52 ( .A(N11), .Z(n244) );
  BUF_X1 U53 ( .A(N11), .Z(n245) );
  BUF_X1 U54 ( .A(N11), .Z(n246) );
  INV_X1 U55 ( .A(N10), .ZN(n253) );
  BUF_X1 U56 ( .A(N12), .Z(n243) );
  NOR3_X1 U57 ( .A1(n255), .A2(N10), .A3(n254), .ZN(n1125) );
  NOR3_X1 U58 ( .A1(n255), .A2(n253), .A3(n254), .ZN(n1115) );
  NOR3_X1 U59 ( .A1(n253), .A2(N11), .A3(n255), .ZN(n1136) );
  NOR3_X1 U60 ( .A1(N10), .A2(N12), .A3(n254), .ZN(n1084) );
  NOR3_X1 U61 ( .A1(n253), .A2(N12), .A3(n254), .ZN(n1074) );
  NOR3_X1 U62 ( .A1(N10), .A2(N11), .A3(n255), .ZN(n1064) );
  NAND2_X1 U63 ( .A1(n1027), .A2(n1136), .ZN(n989) );
  NAND2_X1 U64 ( .A1(n954), .A2(n1136), .ZN(n916) );
  NAND2_X1 U65 ( .A1(n1027), .A2(n1064), .ZN(n998) );
  NAND2_X1 U66 ( .A1(n954), .A2(n1064), .ZN(n925) );
  NAND2_X1 U67 ( .A1(n1027), .A2(n1105), .ZN(n1035) );
  NAND2_X1 U68 ( .A1(n1027), .A2(n1094), .ZN(n1025) );
  NAND2_X1 U69 ( .A1(n954), .A2(n1105), .ZN(n962) );
  NAND2_X1 U70 ( .A1(n954), .A2(n1094), .ZN(n952) );
  NAND2_X1 U71 ( .A1(n1105), .A2(n1135), .ZN(n889) );
  NAND2_X1 U72 ( .A1(n1094), .A2(n1135), .ZN(n880) );
  NAND2_X1 U73 ( .A1(n1084), .A2(n1135), .ZN(n871) );
  NAND2_X1 U74 ( .A1(n1074), .A2(n1135), .ZN(n862) );
  NAND2_X1 U75 ( .A1(n1064), .A2(n1135), .ZN(n853) );
  NAND2_X1 U76 ( .A1(n1136), .A2(n1135), .ZN(n1144) );
  NAND2_X1 U77 ( .A1(n1125), .A2(n1135), .ZN(n1133) );
  NAND2_X1 U78 ( .A1(n1115), .A2(n1135), .ZN(n1123) );
  NAND2_X1 U79 ( .A1(n1027), .A2(n1084), .ZN(n1016) );
  NAND2_X1 U80 ( .A1(n1027), .A2(n1074), .ZN(n1007) );
  NAND2_X1 U81 ( .A1(n954), .A2(n1084), .ZN(n943) );
  NAND2_X1 U82 ( .A1(n954), .A2(n1074), .ZN(n934) );
  NAND2_X1 U83 ( .A1(n1027), .A2(n1125), .ZN(n980) );
  NAND2_X1 U84 ( .A1(n954), .A2(n1125), .ZN(n907) );
  NAND2_X1 U85 ( .A1(n1027), .A2(n1115), .ZN(n971) );
  NAND2_X1 U86 ( .A1(n954), .A2(n1115), .ZN(n898) );
  AND3_X1 U87 ( .A1(n844), .A2(n845), .A3(wr_en), .ZN(n1104) );
  AND3_X1 U88 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1135) );
  AND3_X1 U89 ( .A1(N13), .A2(n845), .A3(wr_en), .ZN(n1027) );
  AND3_X1 U90 ( .A1(N14), .A2(n844), .A3(wr_en), .ZN(n954) );
  INV_X1 U91 ( .A(n1063), .ZN(n771) );
  AOI22_X1 U92 ( .A1(data_in[0]), .A2(n838), .B1(n1062), .B2(\mem[5][0] ), 
        .ZN(n1063) );
  INV_X1 U93 ( .A(n1061), .ZN(n770) );
  AOI22_X1 U94 ( .A1(data_in[1]), .A2(n838), .B1(n1062), .B2(\mem[5][1] ), 
        .ZN(n1061) );
  INV_X1 U95 ( .A(n1060), .ZN(n769) );
  AOI22_X1 U96 ( .A1(data_in[2]), .A2(n838), .B1(n1062), .B2(\mem[5][2] ), 
        .ZN(n1060) );
  INV_X1 U97 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U98 ( .A1(data_in[3]), .A2(n838), .B1(n1062), .B2(\mem[5][3] ), 
        .ZN(n1059) );
  INV_X1 U99 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U100 ( .A1(data_in[4]), .A2(n838), .B1(n1062), .B2(\mem[5][4] ), 
        .ZN(n1058) );
  INV_X1 U101 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U102 ( .A1(data_in[5]), .A2(n838), .B1(n1062), .B2(\mem[5][5] ), 
        .ZN(n1057) );
  INV_X1 U103 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U104 ( .A1(data_in[6]), .A2(n838), .B1(n1062), .B2(\mem[5][6] ), 
        .ZN(n1056) );
  INV_X1 U105 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U106 ( .A1(data_in[7]), .A2(n838), .B1(n1062), .B2(\mem[5][7] ), 
        .ZN(n1055) );
  INV_X1 U107 ( .A(n1024), .ZN(n738) );
  AOI22_X1 U108 ( .A1(data_in[1]), .A2(n834), .B1(n1025), .B2(\mem[9][1] ), 
        .ZN(n1024) );
  INV_X1 U109 ( .A(n1023), .ZN(n737) );
  AOI22_X1 U110 ( .A1(data_in[2]), .A2(n834), .B1(n1025), .B2(\mem[9][2] ), 
        .ZN(n1023) );
  INV_X1 U111 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U112 ( .A1(data_in[3]), .A2(n834), .B1(n1025), .B2(\mem[9][3] ), 
        .ZN(n1022) );
  INV_X1 U113 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U114 ( .A1(data_in[4]), .A2(n834), .B1(n1025), .B2(\mem[9][4] ), 
        .ZN(n1021) );
  INV_X1 U115 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U116 ( .A1(data_in[5]), .A2(n834), .B1(n1025), .B2(\mem[9][5] ), 
        .ZN(n1020) );
  INV_X1 U117 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U118 ( .A1(data_in[6]), .A2(n834), .B1(n1025), .B2(\mem[9][6] ), 
        .ZN(n1019) );
  INV_X1 U119 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U120 ( .A1(data_in[7]), .A2(n834), .B1(n1025), .B2(\mem[9][7] ), 
        .ZN(n1018) );
  INV_X1 U121 ( .A(n990), .ZN(n707) );
  AOI22_X1 U122 ( .A1(data_in[0]), .A2(n830), .B1(n989), .B2(\mem[13][0] ), 
        .ZN(n990) );
  INV_X1 U123 ( .A(n987), .ZN(n705) );
  AOI22_X1 U124 ( .A1(data_in[2]), .A2(n830), .B1(n989), .B2(\mem[13][2] ), 
        .ZN(n987) );
  INV_X1 U125 ( .A(n986), .ZN(n704) );
  AOI22_X1 U126 ( .A1(data_in[3]), .A2(n830), .B1(n989), .B2(\mem[13][3] ), 
        .ZN(n986) );
  INV_X1 U127 ( .A(n985), .ZN(n703) );
  AOI22_X1 U128 ( .A1(data_in[4]), .A2(n830), .B1(n989), .B2(\mem[13][4] ), 
        .ZN(n985) );
  INV_X1 U129 ( .A(n984), .ZN(n702) );
  AOI22_X1 U130 ( .A1(data_in[5]), .A2(n830), .B1(n989), .B2(\mem[13][5] ), 
        .ZN(n984) );
  INV_X1 U131 ( .A(n983), .ZN(n701) );
  AOI22_X1 U132 ( .A1(data_in[6]), .A2(n830), .B1(n989), .B2(\mem[13][6] ), 
        .ZN(n983) );
  INV_X1 U133 ( .A(n982), .ZN(n700) );
  AOI22_X1 U134 ( .A1(data_in[7]), .A2(n830), .B1(n989), .B2(\mem[13][7] ), 
        .ZN(n982) );
  INV_X1 U135 ( .A(n917), .ZN(n643) );
  AOI22_X1 U136 ( .A1(data_in[0]), .A2(n822), .B1(n916), .B2(\mem[21][0] ), 
        .ZN(n917) );
  INV_X1 U137 ( .A(n915), .ZN(n642) );
  AOI22_X1 U138 ( .A1(data_in[1]), .A2(n822), .B1(n916), .B2(\mem[21][1] ), 
        .ZN(n915) );
  INV_X1 U139 ( .A(n914), .ZN(n641) );
  AOI22_X1 U140 ( .A1(data_in[2]), .A2(n822), .B1(n916), .B2(\mem[21][2] ), 
        .ZN(n914) );
  INV_X1 U141 ( .A(n913), .ZN(n640) );
  AOI22_X1 U142 ( .A1(data_in[3]), .A2(n822), .B1(n916), .B2(\mem[21][3] ), 
        .ZN(n913) );
  INV_X1 U143 ( .A(n912), .ZN(n639) );
  AOI22_X1 U144 ( .A1(data_in[4]), .A2(n822), .B1(n916), .B2(\mem[21][4] ), 
        .ZN(n912) );
  INV_X1 U145 ( .A(n911), .ZN(n638) );
  AOI22_X1 U146 ( .A1(data_in[5]), .A2(n822), .B1(n916), .B2(\mem[21][5] ), 
        .ZN(n911) );
  INV_X1 U147 ( .A(n910), .ZN(n637) );
  AOI22_X1 U148 ( .A1(data_in[6]), .A2(n822), .B1(n916), .B2(\mem[21][6] ), 
        .ZN(n910) );
  INV_X1 U149 ( .A(n909), .ZN(n636) );
  AOI22_X1 U150 ( .A1(data_in[7]), .A2(n822), .B1(n916), .B2(\mem[21][7] ), 
        .ZN(n909) );
  INV_X1 U151 ( .A(n1026), .ZN(n739) );
  AOI22_X1 U152 ( .A1(data_in[0]), .A2(n834), .B1(n1025), .B2(\mem[9][0] ), 
        .ZN(n1026) );
  INV_X1 U153 ( .A(n988), .ZN(n706) );
  AOI22_X1 U154 ( .A1(data_in[1]), .A2(n830), .B1(n989), .B2(\mem[13][1] ), 
        .ZN(n988) );
  INV_X1 U155 ( .A(n953), .ZN(n675) );
  AOI22_X1 U156 ( .A1(data_in[0]), .A2(n826), .B1(n952), .B2(\mem[17][0] ), 
        .ZN(n953) );
  INV_X1 U157 ( .A(n951), .ZN(n674) );
  AOI22_X1 U158 ( .A1(data_in[1]), .A2(n826), .B1(n952), .B2(\mem[17][1] ), 
        .ZN(n951) );
  INV_X1 U159 ( .A(n950), .ZN(n673) );
  AOI22_X1 U160 ( .A1(data_in[2]), .A2(n826), .B1(n952), .B2(\mem[17][2] ), 
        .ZN(n950) );
  INV_X1 U161 ( .A(n949), .ZN(n672) );
  AOI22_X1 U162 ( .A1(data_in[3]), .A2(n826), .B1(n952), .B2(\mem[17][3] ), 
        .ZN(n949) );
  INV_X1 U163 ( .A(n948), .ZN(n671) );
  AOI22_X1 U164 ( .A1(data_in[4]), .A2(n826), .B1(n952), .B2(\mem[17][4] ), 
        .ZN(n948) );
  INV_X1 U165 ( .A(n947), .ZN(n670) );
  AOI22_X1 U166 ( .A1(data_in[5]), .A2(n826), .B1(n952), .B2(\mem[17][5] ), 
        .ZN(n947) );
  INV_X1 U167 ( .A(n946), .ZN(n669) );
  AOI22_X1 U168 ( .A1(data_in[6]), .A2(n826), .B1(n952), .B2(\mem[17][6] ), 
        .ZN(n946) );
  INV_X1 U169 ( .A(n945), .ZN(n668) );
  AOI22_X1 U170 ( .A1(data_in[7]), .A2(n826), .B1(n952), .B2(\mem[17][7] ), 
        .ZN(n945) );
  INV_X1 U171 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U172 ( .A1(data_in[0]), .A2(n837), .B1(n1053), .B2(\mem[6][0] ), 
        .ZN(n1054) );
  INV_X1 U173 ( .A(n1052), .ZN(n762) );
  AOI22_X1 U174 ( .A1(data_in[1]), .A2(n837), .B1(n1053), .B2(\mem[6][1] ), 
        .ZN(n1052) );
  INV_X1 U175 ( .A(n1051), .ZN(n761) );
  AOI22_X1 U176 ( .A1(data_in[2]), .A2(n837), .B1(n1053), .B2(\mem[6][2] ), 
        .ZN(n1051) );
  INV_X1 U177 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U178 ( .A1(data_in[3]), .A2(n837), .B1(n1053), .B2(\mem[6][3] ), 
        .ZN(n1050) );
  INV_X1 U179 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U180 ( .A1(data_in[4]), .A2(n837), .B1(n1053), .B2(\mem[6][4] ), 
        .ZN(n1049) );
  INV_X1 U181 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U182 ( .A1(data_in[5]), .A2(n837), .B1(n1053), .B2(\mem[6][5] ), 
        .ZN(n1048) );
  INV_X1 U183 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U184 ( .A1(data_in[6]), .A2(n837), .B1(n1053), .B2(\mem[6][6] ), 
        .ZN(n1047) );
  INV_X1 U185 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U186 ( .A1(data_in[7]), .A2(n837), .B1(n1053), .B2(\mem[6][7] ), 
        .ZN(n1046) );
  INV_X1 U187 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U188 ( .A1(data_in[0]), .A2(n836), .B1(n1044), .B2(\mem[7][0] ), 
        .ZN(n1045) );
  INV_X1 U189 ( .A(n1043), .ZN(n754) );
  AOI22_X1 U190 ( .A1(data_in[1]), .A2(n836), .B1(n1044), .B2(\mem[7][1] ), 
        .ZN(n1043) );
  INV_X1 U191 ( .A(n1042), .ZN(n753) );
  AOI22_X1 U192 ( .A1(data_in[2]), .A2(n836), .B1(n1044), .B2(\mem[7][2] ), 
        .ZN(n1042) );
  INV_X1 U193 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U194 ( .A1(data_in[3]), .A2(n836), .B1(n1044), .B2(\mem[7][3] ), 
        .ZN(n1041) );
  INV_X1 U195 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U196 ( .A1(data_in[4]), .A2(n836), .B1(n1044), .B2(\mem[7][4] ), 
        .ZN(n1040) );
  INV_X1 U197 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U198 ( .A1(data_in[5]), .A2(n836), .B1(n1044), .B2(\mem[7][5] ), 
        .ZN(n1039) );
  INV_X1 U199 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U200 ( .A1(data_in[6]), .A2(n836), .B1(n1044), .B2(\mem[7][6] ), 
        .ZN(n1038) );
  INV_X1 U201 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U202 ( .A1(data_in[7]), .A2(n836), .B1(n1044), .B2(\mem[7][7] ), 
        .ZN(n1037) );
  INV_X1 U203 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U204 ( .A1(data_in[0]), .A2(n833), .B1(n1016), .B2(\mem[10][0] ), 
        .ZN(n1017) );
  INV_X1 U205 ( .A(n1015), .ZN(n730) );
  AOI22_X1 U206 ( .A1(data_in[1]), .A2(n833), .B1(n1016), .B2(\mem[10][1] ), 
        .ZN(n1015) );
  INV_X1 U207 ( .A(n1014), .ZN(n729) );
  AOI22_X1 U208 ( .A1(data_in[2]), .A2(n833), .B1(n1016), .B2(\mem[10][2] ), 
        .ZN(n1014) );
  INV_X1 U209 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U210 ( .A1(data_in[3]), .A2(n833), .B1(n1016), .B2(\mem[10][3] ), 
        .ZN(n1013) );
  INV_X1 U211 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U212 ( .A1(data_in[4]), .A2(n833), .B1(n1016), .B2(\mem[10][4] ), 
        .ZN(n1012) );
  INV_X1 U213 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U214 ( .A1(data_in[5]), .A2(n833), .B1(n1016), .B2(\mem[10][5] ), 
        .ZN(n1011) );
  INV_X1 U215 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U216 ( .A1(data_in[6]), .A2(n833), .B1(n1016), .B2(\mem[10][6] ), 
        .ZN(n1010) );
  INV_X1 U217 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U218 ( .A1(data_in[7]), .A2(n833), .B1(n1016), .B2(\mem[10][7] ), 
        .ZN(n1009) );
  INV_X1 U219 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U220 ( .A1(data_in[0]), .A2(n832), .B1(n1007), .B2(\mem[11][0] ), 
        .ZN(n1008) );
  INV_X1 U221 ( .A(n1006), .ZN(n722) );
  AOI22_X1 U222 ( .A1(data_in[1]), .A2(n832), .B1(n1007), .B2(\mem[11][1] ), 
        .ZN(n1006) );
  INV_X1 U223 ( .A(n1005), .ZN(n721) );
  AOI22_X1 U224 ( .A1(data_in[2]), .A2(n832), .B1(n1007), .B2(\mem[11][2] ), 
        .ZN(n1005) );
  INV_X1 U225 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U226 ( .A1(data_in[3]), .A2(n832), .B1(n1007), .B2(\mem[11][3] ), 
        .ZN(n1004) );
  INV_X1 U227 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U228 ( .A1(data_in[4]), .A2(n832), .B1(n1007), .B2(\mem[11][4] ), 
        .ZN(n1003) );
  INV_X1 U229 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U230 ( .A1(data_in[5]), .A2(n832), .B1(n1007), .B2(\mem[11][5] ), 
        .ZN(n1002) );
  INV_X1 U231 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U232 ( .A1(data_in[6]), .A2(n832), .B1(n1007), .B2(\mem[11][6] ), 
        .ZN(n1001) );
  INV_X1 U233 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U234 ( .A1(data_in[7]), .A2(n832), .B1(n1007), .B2(\mem[11][7] ), 
        .ZN(n1000) );
  INV_X1 U235 ( .A(n981), .ZN(n699) );
  AOI22_X1 U236 ( .A1(data_in[0]), .A2(n829), .B1(n980), .B2(\mem[14][0] ), 
        .ZN(n981) );
  INV_X1 U237 ( .A(n979), .ZN(n698) );
  AOI22_X1 U238 ( .A1(data_in[1]), .A2(n829), .B1(n980), .B2(\mem[14][1] ), 
        .ZN(n979) );
  INV_X1 U239 ( .A(n978), .ZN(n697) );
  AOI22_X1 U240 ( .A1(data_in[2]), .A2(n829), .B1(n980), .B2(\mem[14][2] ), 
        .ZN(n978) );
  INV_X1 U241 ( .A(n977), .ZN(n696) );
  AOI22_X1 U242 ( .A1(data_in[3]), .A2(n829), .B1(n980), .B2(\mem[14][3] ), 
        .ZN(n977) );
  INV_X1 U243 ( .A(n976), .ZN(n695) );
  AOI22_X1 U244 ( .A1(data_in[4]), .A2(n829), .B1(n980), .B2(\mem[14][4] ), 
        .ZN(n976) );
  INV_X1 U245 ( .A(n975), .ZN(n694) );
  AOI22_X1 U246 ( .A1(data_in[5]), .A2(n829), .B1(n980), .B2(\mem[14][5] ), 
        .ZN(n975) );
  INV_X1 U247 ( .A(n974), .ZN(n693) );
  AOI22_X1 U248 ( .A1(data_in[6]), .A2(n829), .B1(n980), .B2(\mem[14][6] ), 
        .ZN(n974) );
  INV_X1 U249 ( .A(n973), .ZN(n692) );
  AOI22_X1 U250 ( .A1(data_in[7]), .A2(n829), .B1(n980), .B2(\mem[14][7] ), 
        .ZN(n973) );
  INV_X1 U251 ( .A(n972), .ZN(n691) );
  AOI22_X1 U252 ( .A1(data_in[0]), .A2(n828), .B1(n971), .B2(\mem[15][0] ), 
        .ZN(n972) );
  INV_X1 U253 ( .A(n970), .ZN(n690) );
  AOI22_X1 U254 ( .A1(data_in[1]), .A2(n828), .B1(n971), .B2(\mem[15][1] ), 
        .ZN(n970) );
  INV_X1 U255 ( .A(n969), .ZN(n689) );
  AOI22_X1 U256 ( .A1(data_in[2]), .A2(n828), .B1(n971), .B2(\mem[15][2] ), 
        .ZN(n969) );
  INV_X1 U257 ( .A(n968), .ZN(n688) );
  AOI22_X1 U258 ( .A1(data_in[3]), .A2(n828), .B1(n971), .B2(\mem[15][3] ), 
        .ZN(n968) );
  INV_X1 U259 ( .A(n967), .ZN(n687) );
  AOI22_X1 U260 ( .A1(data_in[4]), .A2(n828), .B1(n971), .B2(\mem[15][4] ), 
        .ZN(n967) );
  INV_X1 U261 ( .A(n966), .ZN(n686) );
  AOI22_X1 U262 ( .A1(data_in[5]), .A2(n828), .B1(n971), .B2(\mem[15][5] ), 
        .ZN(n966) );
  INV_X1 U263 ( .A(n965), .ZN(n685) );
  AOI22_X1 U264 ( .A1(data_in[6]), .A2(n828), .B1(n971), .B2(\mem[15][6] ), 
        .ZN(n965) );
  INV_X1 U265 ( .A(n964), .ZN(n684) );
  AOI22_X1 U266 ( .A1(data_in[7]), .A2(n828), .B1(n971), .B2(\mem[15][7] ), 
        .ZN(n964) );
  INV_X1 U267 ( .A(n944), .ZN(n667) );
  AOI22_X1 U268 ( .A1(data_in[0]), .A2(n825), .B1(n943), .B2(\mem[18][0] ), 
        .ZN(n944) );
  INV_X1 U269 ( .A(n942), .ZN(n666) );
  AOI22_X1 U270 ( .A1(data_in[1]), .A2(n825), .B1(n943), .B2(\mem[18][1] ), 
        .ZN(n942) );
  INV_X1 U271 ( .A(n941), .ZN(n665) );
  AOI22_X1 U272 ( .A1(data_in[2]), .A2(n825), .B1(n943), .B2(\mem[18][2] ), 
        .ZN(n941) );
  INV_X1 U273 ( .A(n940), .ZN(n664) );
  AOI22_X1 U274 ( .A1(data_in[3]), .A2(n825), .B1(n943), .B2(\mem[18][3] ), 
        .ZN(n940) );
  INV_X1 U275 ( .A(n939), .ZN(n663) );
  AOI22_X1 U276 ( .A1(data_in[4]), .A2(n825), .B1(n943), .B2(\mem[18][4] ), 
        .ZN(n939) );
  INV_X1 U277 ( .A(n938), .ZN(n662) );
  AOI22_X1 U278 ( .A1(data_in[5]), .A2(n825), .B1(n943), .B2(\mem[18][5] ), 
        .ZN(n938) );
  INV_X1 U279 ( .A(n937), .ZN(n661) );
  AOI22_X1 U280 ( .A1(data_in[6]), .A2(n825), .B1(n943), .B2(\mem[18][6] ), 
        .ZN(n937) );
  INV_X1 U281 ( .A(n936), .ZN(n660) );
  AOI22_X1 U282 ( .A1(data_in[7]), .A2(n825), .B1(n943), .B2(\mem[18][7] ), 
        .ZN(n936) );
  INV_X1 U283 ( .A(n935), .ZN(n659) );
  AOI22_X1 U284 ( .A1(data_in[0]), .A2(n824), .B1(n934), .B2(\mem[19][0] ), 
        .ZN(n935) );
  INV_X1 U285 ( .A(n933), .ZN(n658) );
  AOI22_X1 U286 ( .A1(data_in[1]), .A2(n824), .B1(n934), .B2(\mem[19][1] ), 
        .ZN(n933) );
  INV_X1 U287 ( .A(n932), .ZN(n657) );
  AOI22_X1 U288 ( .A1(data_in[2]), .A2(n824), .B1(n934), .B2(\mem[19][2] ), 
        .ZN(n932) );
  INV_X1 U289 ( .A(n931), .ZN(n656) );
  AOI22_X1 U290 ( .A1(data_in[3]), .A2(n824), .B1(n934), .B2(\mem[19][3] ), 
        .ZN(n931) );
  INV_X1 U291 ( .A(n930), .ZN(n655) );
  AOI22_X1 U292 ( .A1(data_in[4]), .A2(n824), .B1(n934), .B2(\mem[19][4] ), 
        .ZN(n930) );
  INV_X1 U293 ( .A(n929), .ZN(n654) );
  AOI22_X1 U294 ( .A1(data_in[5]), .A2(n824), .B1(n934), .B2(\mem[19][5] ), 
        .ZN(n929) );
  INV_X1 U295 ( .A(n928), .ZN(n653) );
  AOI22_X1 U296 ( .A1(data_in[6]), .A2(n824), .B1(n934), .B2(\mem[19][6] ), 
        .ZN(n928) );
  INV_X1 U297 ( .A(n927), .ZN(n652) );
  AOI22_X1 U298 ( .A1(data_in[7]), .A2(n824), .B1(n934), .B2(\mem[19][7] ), 
        .ZN(n927) );
  INV_X1 U299 ( .A(n908), .ZN(n635) );
  AOI22_X1 U300 ( .A1(data_in[0]), .A2(n821), .B1(n907), .B2(\mem[22][0] ), 
        .ZN(n908) );
  INV_X1 U301 ( .A(n906), .ZN(n634) );
  AOI22_X1 U302 ( .A1(data_in[1]), .A2(n821), .B1(n907), .B2(\mem[22][1] ), 
        .ZN(n906) );
  INV_X1 U303 ( .A(n905), .ZN(n633) );
  AOI22_X1 U304 ( .A1(data_in[2]), .A2(n821), .B1(n907), .B2(\mem[22][2] ), 
        .ZN(n905) );
  INV_X1 U305 ( .A(n904), .ZN(n632) );
  AOI22_X1 U306 ( .A1(data_in[3]), .A2(n821), .B1(n907), .B2(\mem[22][3] ), 
        .ZN(n904) );
  INV_X1 U307 ( .A(n903), .ZN(n631) );
  AOI22_X1 U308 ( .A1(data_in[4]), .A2(n821), .B1(n907), .B2(\mem[22][4] ), 
        .ZN(n903) );
  INV_X1 U309 ( .A(n902), .ZN(n630) );
  AOI22_X1 U310 ( .A1(data_in[5]), .A2(n821), .B1(n907), .B2(\mem[22][5] ), 
        .ZN(n902) );
  INV_X1 U311 ( .A(n901), .ZN(n629) );
  AOI22_X1 U312 ( .A1(data_in[6]), .A2(n821), .B1(n907), .B2(\mem[22][6] ), 
        .ZN(n901) );
  INV_X1 U313 ( .A(n900), .ZN(n628) );
  AOI22_X1 U314 ( .A1(data_in[7]), .A2(n821), .B1(n907), .B2(\mem[22][7] ), 
        .ZN(n900) );
  INV_X1 U315 ( .A(n899), .ZN(n627) );
  AOI22_X1 U316 ( .A1(data_in[0]), .A2(n820), .B1(n898), .B2(\mem[23][0] ), 
        .ZN(n899) );
  INV_X1 U317 ( .A(n897), .ZN(n626) );
  AOI22_X1 U318 ( .A1(data_in[1]), .A2(n820), .B1(n898), .B2(\mem[23][1] ), 
        .ZN(n897) );
  INV_X1 U319 ( .A(n896), .ZN(n625) );
  AOI22_X1 U320 ( .A1(data_in[2]), .A2(n820), .B1(n898), .B2(\mem[23][2] ), 
        .ZN(n896) );
  INV_X1 U321 ( .A(n895), .ZN(n624) );
  AOI22_X1 U322 ( .A1(data_in[3]), .A2(n820), .B1(n898), .B2(\mem[23][3] ), 
        .ZN(n895) );
  INV_X1 U323 ( .A(n894), .ZN(n623) );
  AOI22_X1 U324 ( .A1(data_in[4]), .A2(n820), .B1(n898), .B2(\mem[23][4] ), 
        .ZN(n894) );
  INV_X1 U325 ( .A(n893), .ZN(n622) );
  AOI22_X1 U326 ( .A1(data_in[5]), .A2(n820), .B1(n898), .B2(\mem[23][5] ), 
        .ZN(n893) );
  INV_X1 U327 ( .A(n892), .ZN(n621) );
  AOI22_X1 U328 ( .A1(data_in[6]), .A2(n820), .B1(n898), .B2(\mem[23][6] ), 
        .ZN(n892) );
  INV_X1 U329 ( .A(n891), .ZN(n620) );
  AOI22_X1 U330 ( .A1(data_in[7]), .A2(n820), .B1(n898), .B2(\mem[23][7] ), 
        .ZN(n891) );
  INV_X1 U331 ( .A(N12), .ZN(n255) );
  INV_X1 U332 ( .A(N11), .ZN(n254) );
  INV_X1 U333 ( .A(n999), .ZN(n715) );
  AOI22_X1 U334 ( .A1(data_in[0]), .A2(n831), .B1(n998), .B2(\mem[12][0] ), 
        .ZN(n999) );
  INV_X1 U335 ( .A(n997), .ZN(n714) );
  AOI22_X1 U336 ( .A1(data_in[1]), .A2(n831), .B1(n998), .B2(\mem[12][1] ), 
        .ZN(n997) );
  INV_X1 U337 ( .A(n996), .ZN(n713) );
  AOI22_X1 U338 ( .A1(data_in[2]), .A2(n831), .B1(n998), .B2(\mem[12][2] ), 
        .ZN(n996) );
  INV_X1 U339 ( .A(n995), .ZN(n712) );
  AOI22_X1 U340 ( .A1(data_in[3]), .A2(n831), .B1(n998), .B2(\mem[12][3] ), 
        .ZN(n995) );
  INV_X1 U341 ( .A(n994), .ZN(n711) );
  AOI22_X1 U342 ( .A1(data_in[4]), .A2(n831), .B1(n998), .B2(\mem[12][4] ), 
        .ZN(n994) );
  INV_X1 U343 ( .A(n993), .ZN(n710) );
  AOI22_X1 U344 ( .A1(data_in[5]), .A2(n831), .B1(n998), .B2(\mem[12][5] ), 
        .ZN(n993) );
  INV_X1 U345 ( .A(n992), .ZN(n709) );
  AOI22_X1 U346 ( .A1(data_in[6]), .A2(n831), .B1(n998), .B2(\mem[12][6] ), 
        .ZN(n992) );
  INV_X1 U347 ( .A(n991), .ZN(n708) );
  AOI22_X1 U348 ( .A1(data_in[7]), .A2(n831), .B1(n998), .B2(\mem[12][7] ), 
        .ZN(n991) );
  INV_X1 U349 ( .A(n926), .ZN(n651) );
  AOI22_X1 U350 ( .A1(data_in[0]), .A2(n823), .B1(n925), .B2(\mem[20][0] ), 
        .ZN(n926) );
  INV_X1 U351 ( .A(n924), .ZN(n650) );
  AOI22_X1 U352 ( .A1(data_in[1]), .A2(n823), .B1(n925), .B2(\mem[20][1] ), 
        .ZN(n924) );
  INV_X1 U353 ( .A(n923), .ZN(n649) );
  AOI22_X1 U354 ( .A1(data_in[2]), .A2(n823), .B1(n925), .B2(\mem[20][2] ), 
        .ZN(n923) );
  INV_X1 U355 ( .A(n922), .ZN(n648) );
  AOI22_X1 U356 ( .A1(data_in[3]), .A2(n823), .B1(n925), .B2(\mem[20][3] ), 
        .ZN(n922) );
  INV_X1 U357 ( .A(n921), .ZN(n647) );
  AOI22_X1 U358 ( .A1(data_in[4]), .A2(n823), .B1(n925), .B2(\mem[20][4] ), 
        .ZN(n921) );
  INV_X1 U359 ( .A(n920), .ZN(n646) );
  AOI22_X1 U360 ( .A1(data_in[5]), .A2(n823), .B1(n925), .B2(\mem[20][5] ), 
        .ZN(n920) );
  INV_X1 U361 ( .A(n919), .ZN(n645) );
  AOI22_X1 U362 ( .A1(data_in[6]), .A2(n823), .B1(n925), .B2(\mem[20][6] ), 
        .ZN(n919) );
  INV_X1 U363 ( .A(n918), .ZN(n644) );
  AOI22_X1 U364 ( .A1(data_in[7]), .A2(n823), .B1(n925), .B2(\mem[20][7] ), 
        .ZN(n918) );
  INV_X1 U365 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U366 ( .A1(data_in[0]), .A2(n835), .B1(n1035), .B2(\mem[8][0] ), 
        .ZN(n1036) );
  INV_X1 U367 ( .A(n1034), .ZN(n746) );
  AOI22_X1 U368 ( .A1(data_in[1]), .A2(n835), .B1(n1035), .B2(\mem[8][1] ), 
        .ZN(n1034) );
  INV_X1 U369 ( .A(n1033), .ZN(n745) );
  AOI22_X1 U370 ( .A1(data_in[2]), .A2(n835), .B1(n1035), .B2(\mem[8][2] ), 
        .ZN(n1033) );
  INV_X1 U371 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U372 ( .A1(data_in[3]), .A2(n835), .B1(n1035), .B2(\mem[8][3] ), 
        .ZN(n1032) );
  INV_X1 U373 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U374 ( .A1(data_in[4]), .A2(n835), .B1(n1035), .B2(\mem[8][4] ), 
        .ZN(n1031) );
  INV_X1 U375 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U376 ( .A1(data_in[5]), .A2(n835), .B1(n1035), .B2(\mem[8][5] ), 
        .ZN(n1030) );
  INV_X1 U377 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U378 ( .A1(data_in[6]), .A2(n835), .B1(n1035), .B2(\mem[8][6] ), 
        .ZN(n1029) );
  INV_X1 U379 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U380 ( .A1(data_in[7]), .A2(n835), .B1(n1035), .B2(\mem[8][7] ), 
        .ZN(n1028) );
  INV_X1 U381 ( .A(n963), .ZN(n683) );
  AOI22_X1 U382 ( .A1(data_in[0]), .A2(n827), .B1(n962), .B2(\mem[16][0] ), 
        .ZN(n963) );
  INV_X1 U383 ( .A(n961), .ZN(n682) );
  AOI22_X1 U384 ( .A1(data_in[1]), .A2(n827), .B1(n962), .B2(\mem[16][1] ), 
        .ZN(n961) );
  INV_X1 U385 ( .A(n960), .ZN(n681) );
  AOI22_X1 U386 ( .A1(data_in[2]), .A2(n827), .B1(n962), .B2(\mem[16][2] ), 
        .ZN(n960) );
  INV_X1 U387 ( .A(n959), .ZN(n680) );
  AOI22_X1 U388 ( .A1(data_in[3]), .A2(n827), .B1(n962), .B2(\mem[16][3] ), 
        .ZN(n959) );
  INV_X1 U389 ( .A(n958), .ZN(n679) );
  AOI22_X1 U390 ( .A1(data_in[4]), .A2(n827), .B1(n962), .B2(\mem[16][4] ), 
        .ZN(n958) );
  INV_X1 U391 ( .A(n957), .ZN(n678) );
  AOI22_X1 U392 ( .A1(data_in[5]), .A2(n827), .B1(n962), .B2(\mem[16][5] ), 
        .ZN(n957) );
  INV_X1 U393 ( .A(n956), .ZN(n677) );
  AOI22_X1 U394 ( .A1(data_in[6]), .A2(n827), .B1(n962), .B2(\mem[16][6] ), 
        .ZN(n956) );
  INV_X1 U395 ( .A(n955), .ZN(n676) );
  AOI22_X1 U396 ( .A1(data_in[7]), .A2(n827), .B1(n962), .B2(\mem[16][7] ), 
        .ZN(n955) );
  INV_X1 U397 ( .A(n890), .ZN(n619) );
  AOI22_X1 U398 ( .A1(data_in[0]), .A2(n816), .B1(n889), .B2(\mem[24][0] ), 
        .ZN(n890) );
  INV_X1 U399 ( .A(n888), .ZN(n618) );
  AOI22_X1 U400 ( .A1(data_in[1]), .A2(n816), .B1(n889), .B2(\mem[24][1] ), 
        .ZN(n888) );
  INV_X1 U401 ( .A(n887), .ZN(n617) );
  AOI22_X1 U402 ( .A1(data_in[2]), .A2(n816), .B1(n889), .B2(\mem[24][2] ), 
        .ZN(n887) );
  INV_X1 U403 ( .A(n886), .ZN(n616) );
  AOI22_X1 U404 ( .A1(data_in[3]), .A2(n816), .B1(n889), .B2(\mem[24][3] ), 
        .ZN(n886) );
  INV_X1 U405 ( .A(n885), .ZN(n615) );
  AOI22_X1 U406 ( .A1(data_in[4]), .A2(n816), .B1(n889), .B2(\mem[24][4] ), 
        .ZN(n885) );
  INV_X1 U407 ( .A(n884), .ZN(n614) );
  AOI22_X1 U408 ( .A1(data_in[5]), .A2(n816), .B1(n889), .B2(\mem[24][5] ), 
        .ZN(n884) );
  INV_X1 U409 ( .A(n883), .ZN(n613) );
  AOI22_X1 U410 ( .A1(data_in[6]), .A2(n816), .B1(n889), .B2(\mem[24][6] ), 
        .ZN(n883) );
  INV_X1 U411 ( .A(n882), .ZN(n612) );
  AOI22_X1 U412 ( .A1(data_in[7]), .A2(n816), .B1(n889), .B2(\mem[24][7] ), 
        .ZN(n882) );
  INV_X1 U413 ( .A(n881), .ZN(n611) );
  AOI22_X1 U414 ( .A1(data_in[0]), .A2(n815), .B1(n880), .B2(\mem[25][0] ), 
        .ZN(n881) );
  INV_X1 U415 ( .A(n879), .ZN(n610) );
  AOI22_X1 U416 ( .A1(data_in[1]), .A2(n815), .B1(n880), .B2(\mem[25][1] ), 
        .ZN(n879) );
  INV_X1 U417 ( .A(n878), .ZN(n609) );
  AOI22_X1 U418 ( .A1(data_in[2]), .A2(n815), .B1(n880), .B2(\mem[25][2] ), 
        .ZN(n878) );
  INV_X1 U419 ( .A(n877), .ZN(n608) );
  AOI22_X1 U420 ( .A1(data_in[3]), .A2(n815), .B1(n880), .B2(\mem[25][3] ), 
        .ZN(n877) );
  INV_X1 U421 ( .A(n876), .ZN(n607) );
  AOI22_X1 U422 ( .A1(data_in[4]), .A2(n815), .B1(n880), .B2(\mem[25][4] ), 
        .ZN(n876) );
  INV_X1 U423 ( .A(n875), .ZN(n606) );
  AOI22_X1 U424 ( .A1(data_in[5]), .A2(n815), .B1(n880), .B2(\mem[25][5] ), 
        .ZN(n875) );
  INV_X1 U425 ( .A(n874), .ZN(n605) );
  AOI22_X1 U426 ( .A1(data_in[6]), .A2(n815), .B1(n880), .B2(\mem[25][6] ), 
        .ZN(n874) );
  INV_X1 U427 ( .A(n873), .ZN(n604) );
  AOI22_X1 U428 ( .A1(data_in[7]), .A2(n815), .B1(n880), .B2(\mem[25][7] ), 
        .ZN(n873) );
  INV_X1 U429 ( .A(n872), .ZN(n603) );
  AOI22_X1 U430 ( .A1(data_in[0]), .A2(n814), .B1(n871), .B2(\mem[26][0] ), 
        .ZN(n872) );
  INV_X1 U431 ( .A(n870), .ZN(n602) );
  AOI22_X1 U432 ( .A1(data_in[1]), .A2(n814), .B1(n871), .B2(\mem[26][1] ), 
        .ZN(n870) );
  INV_X1 U433 ( .A(n869), .ZN(n601) );
  AOI22_X1 U434 ( .A1(data_in[2]), .A2(n814), .B1(n871), .B2(\mem[26][2] ), 
        .ZN(n869) );
  INV_X1 U435 ( .A(n868), .ZN(n600) );
  AOI22_X1 U436 ( .A1(data_in[3]), .A2(n814), .B1(n871), .B2(\mem[26][3] ), 
        .ZN(n868) );
  INV_X1 U437 ( .A(n867), .ZN(n599) );
  AOI22_X1 U438 ( .A1(data_in[4]), .A2(n814), .B1(n871), .B2(\mem[26][4] ), 
        .ZN(n867) );
  INV_X1 U439 ( .A(n866), .ZN(n598) );
  AOI22_X1 U440 ( .A1(data_in[5]), .A2(n814), .B1(n871), .B2(\mem[26][5] ), 
        .ZN(n866) );
  INV_X1 U441 ( .A(n865), .ZN(n597) );
  AOI22_X1 U442 ( .A1(data_in[6]), .A2(n814), .B1(n871), .B2(\mem[26][6] ), 
        .ZN(n865) );
  INV_X1 U443 ( .A(n864), .ZN(n596) );
  AOI22_X1 U444 ( .A1(data_in[7]), .A2(n814), .B1(n871), .B2(\mem[26][7] ), 
        .ZN(n864) );
  INV_X1 U445 ( .A(n863), .ZN(n595) );
  AOI22_X1 U446 ( .A1(data_in[0]), .A2(n813), .B1(n862), .B2(\mem[27][0] ), 
        .ZN(n863) );
  INV_X1 U447 ( .A(n861), .ZN(n594) );
  AOI22_X1 U448 ( .A1(data_in[1]), .A2(n813), .B1(n862), .B2(\mem[27][1] ), 
        .ZN(n861) );
  INV_X1 U449 ( .A(n860), .ZN(n293) );
  AOI22_X1 U450 ( .A1(data_in[2]), .A2(n813), .B1(n862), .B2(\mem[27][2] ), 
        .ZN(n860) );
  INV_X1 U451 ( .A(n859), .ZN(n292) );
  AOI22_X1 U452 ( .A1(data_in[3]), .A2(n813), .B1(n862), .B2(\mem[27][3] ), 
        .ZN(n859) );
  INV_X1 U453 ( .A(n858), .ZN(n291) );
  AOI22_X1 U454 ( .A1(data_in[4]), .A2(n813), .B1(n862), .B2(\mem[27][4] ), 
        .ZN(n858) );
  INV_X1 U455 ( .A(n857), .ZN(n290) );
  AOI22_X1 U456 ( .A1(data_in[5]), .A2(n813), .B1(n862), .B2(\mem[27][5] ), 
        .ZN(n857) );
  INV_X1 U457 ( .A(n856), .ZN(n289) );
  AOI22_X1 U458 ( .A1(data_in[6]), .A2(n813), .B1(n862), .B2(\mem[27][6] ), 
        .ZN(n856) );
  INV_X1 U459 ( .A(n855), .ZN(n288) );
  AOI22_X1 U460 ( .A1(data_in[7]), .A2(n813), .B1(n862), .B2(\mem[27][7] ), 
        .ZN(n855) );
  INV_X1 U461 ( .A(n854), .ZN(n287) );
  AOI22_X1 U462 ( .A1(data_in[0]), .A2(n812), .B1(n853), .B2(\mem[28][0] ), 
        .ZN(n854) );
  INV_X1 U463 ( .A(n852), .ZN(n286) );
  AOI22_X1 U464 ( .A1(data_in[1]), .A2(n812), .B1(n853), .B2(\mem[28][1] ), 
        .ZN(n852) );
  INV_X1 U465 ( .A(n851), .ZN(n285) );
  AOI22_X1 U466 ( .A1(data_in[2]), .A2(n812), .B1(n853), .B2(\mem[28][2] ), 
        .ZN(n851) );
  INV_X1 U467 ( .A(n850), .ZN(n284) );
  AOI22_X1 U468 ( .A1(data_in[3]), .A2(n812), .B1(n853), .B2(\mem[28][3] ), 
        .ZN(n850) );
  INV_X1 U469 ( .A(n849), .ZN(n283) );
  AOI22_X1 U470 ( .A1(data_in[4]), .A2(n812), .B1(n853), .B2(\mem[28][4] ), 
        .ZN(n849) );
  INV_X1 U471 ( .A(n848), .ZN(n282) );
  AOI22_X1 U472 ( .A1(data_in[5]), .A2(n812), .B1(n853), .B2(\mem[28][5] ), 
        .ZN(n848) );
  INV_X1 U473 ( .A(n847), .ZN(n281) );
  AOI22_X1 U474 ( .A1(data_in[6]), .A2(n812), .B1(n853), .B2(\mem[28][6] ), 
        .ZN(n847) );
  INV_X1 U475 ( .A(n846), .ZN(n280) );
  AOI22_X1 U476 ( .A1(data_in[7]), .A2(n812), .B1(n853), .B2(\mem[28][7] ), 
        .ZN(n846) );
  INV_X1 U477 ( .A(n1145), .ZN(n279) );
  AOI22_X1 U478 ( .A1(n819), .A2(data_in[0]), .B1(n1144), .B2(\mem[29][0] ), 
        .ZN(n1145) );
  INV_X1 U479 ( .A(n1143), .ZN(n278) );
  AOI22_X1 U480 ( .A1(n819), .A2(data_in[1]), .B1(n1144), .B2(\mem[29][1] ), 
        .ZN(n1143) );
  INV_X1 U481 ( .A(n1142), .ZN(n277) );
  AOI22_X1 U482 ( .A1(n819), .A2(data_in[2]), .B1(n1144), .B2(\mem[29][2] ), 
        .ZN(n1142) );
  INV_X1 U483 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U484 ( .A1(n819), .A2(data_in[3]), .B1(n1144), .B2(\mem[29][3] ), 
        .ZN(n1141) );
  INV_X1 U485 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U486 ( .A1(n819), .A2(data_in[4]), .B1(n1144), .B2(\mem[29][4] ), 
        .ZN(n1140) );
  INV_X1 U487 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U488 ( .A1(n819), .A2(data_in[5]), .B1(n1144), .B2(\mem[29][5] ), 
        .ZN(n1139) );
  INV_X1 U489 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U490 ( .A1(n819), .A2(data_in[6]), .B1(n1144), .B2(\mem[29][6] ), 
        .ZN(n1138) );
  INV_X1 U491 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U492 ( .A1(n819), .A2(data_in[7]), .B1(n1144), .B2(\mem[29][7] ), 
        .ZN(n1137) );
  INV_X1 U493 ( .A(n1134), .ZN(n271) );
  AOI22_X1 U494 ( .A1(data_in[0]), .A2(n818), .B1(n1133), .B2(\mem[30][0] ), 
        .ZN(n1134) );
  INV_X1 U495 ( .A(n1132), .ZN(n270) );
  AOI22_X1 U496 ( .A1(data_in[1]), .A2(n818), .B1(n1133), .B2(\mem[30][1] ), 
        .ZN(n1132) );
  INV_X1 U497 ( .A(n1131), .ZN(n269) );
  AOI22_X1 U498 ( .A1(data_in[2]), .A2(n818), .B1(n1133), .B2(\mem[30][2] ), 
        .ZN(n1131) );
  INV_X1 U499 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U500 ( .A1(data_in[3]), .A2(n818), .B1(n1133), .B2(\mem[30][3] ), 
        .ZN(n1130) );
  INV_X1 U501 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U502 ( .A1(data_in[4]), .A2(n818), .B1(n1133), .B2(\mem[30][4] ), 
        .ZN(n1129) );
  INV_X1 U503 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U504 ( .A1(data_in[5]), .A2(n818), .B1(n1133), .B2(\mem[30][5] ), 
        .ZN(n1128) );
  INV_X1 U505 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U506 ( .A1(data_in[6]), .A2(n818), .B1(n1133), .B2(\mem[30][6] ), 
        .ZN(n1127) );
  INV_X1 U507 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U508 ( .A1(data_in[7]), .A2(n818), .B1(n1133), .B2(\mem[30][7] ), 
        .ZN(n1126) );
  INV_X1 U509 ( .A(n1124), .ZN(n263) );
  AOI22_X1 U510 ( .A1(data_in[0]), .A2(n817), .B1(n1123), .B2(\mem[31][0] ), 
        .ZN(n1124) );
  INV_X1 U511 ( .A(n1122), .ZN(n262) );
  AOI22_X1 U512 ( .A1(data_in[1]), .A2(n817), .B1(n1123), .B2(\mem[31][1] ), 
        .ZN(n1122) );
  INV_X1 U513 ( .A(n1121), .ZN(n261) );
  AOI22_X1 U514 ( .A1(data_in[2]), .A2(n817), .B1(n1123), .B2(\mem[31][2] ), 
        .ZN(n1121) );
  INV_X1 U515 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U516 ( .A1(data_in[3]), .A2(n817), .B1(n1123), .B2(\mem[31][3] ), 
        .ZN(n1120) );
  INV_X1 U517 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U518 ( .A1(data_in[4]), .A2(n817), .B1(n1123), .B2(\mem[31][4] ), 
        .ZN(n1119) );
  INV_X1 U519 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U520 ( .A1(data_in[5]), .A2(n817), .B1(n1123), .B2(\mem[31][5] ), 
        .ZN(n1118) );
  INV_X1 U521 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U522 ( .A1(data_in[6]), .A2(n817), .B1(n1123), .B2(\mem[31][6] ), 
        .ZN(n1117) );
  INV_X1 U523 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U524 ( .A1(data_in[7]), .A2(n817), .B1(n1123), .B2(\mem[31][7] ), 
        .ZN(n1116) );
  INV_X1 U525 ( .A(n1114), .ZN(n811) );
  AOI22_X1 U526 ( .A1(data_in[0]), .A2(n843), .B1(n1113), .B2(\mem[0][0] ), 
        .ZN(n1114) );
  INV_X1 U527 ( .A(n1112), .ZN(n810) );
  AOI22_X1 U528 ( .A1(data_in[1]), .A2(n843), .B1(n1113), .B2(\mem[0][1] ), 
        .ZN(n1112) );
  INV_X1 U529 ( .A(n1111), .ZN(n809) );
  AOI22_X1 U530 ( .A1(data_in[2]), .A2(n843), .B1(n1113), .B2(\mem[0][2] ), 
        .ZN(n1111) );
  INV_X1 U531 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U532 ( .A1(data_in[3]), .A2(n843), .B1(n1113), .B2(\mem[0][3] ), 
        .ZN(n1110) );
  INV_X1 U533 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U534 ( .A1(data_in[4]), .A2(n843), .B1(n1113), .B2(\mem[0][4] ), 
        .ZN(n1109) );
  INV_X1 U535 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U536 ( .A1(data_in[5]), .A2(n843), .B1(n1113), .B2(\mem[0][5] ), 
        .ZN(n1108) );
  INV_X1 U537 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U538 ( .A1(data_in[6]), .A2(n843), .B1(n1113), .B2(\mem[0][6] ), 
        .ZN(n1107) );
  INV_X1 U539 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U540 ( .A1(data_in[7]), .A2(n843), .B1(n1113), .B2(\mem[0][7] ), 
        .ZN(n1106) );
  INV_X1 U541 ( .A(n1103), .ZN(n803) );
  AOI22_X1 U542 ( .A1(data_in[0]), .A2(n842), .B1(n1102), .B2(\mem[1][0] ), 
        .ZN(n1103) );
  INV_X1 U543 ( .A(n1101), .ZN(n802) );
  AOI22_X1 U544 ( .A1(data_in[1]), .A2(n842), .B1(n1102), .B2(\mem[1][1] ), 
        .ZN(n1101) );
  INV_X1 U545 ( .A(n1100), .ZN(n801) );
  AOI22_X1 U546 ( .A1(data_in[2]), .A2(n842), .B1(n1102), .B2(\mem[1][2] ), 
        .ZN(n1100) );
  INV_X1 U547 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U548 ( .A1(data_in[3]), .A2(n842), .B1(n1102), .B2(\mem[1][3] ), 
        .ZN(n1099) );
  INV_X1 U549 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U550 ( .A1(data_in[4]), .A2(n842), .B1(n1102), .B2(\mem[1][4] ), 
        .ZN(n1098) );
  INV_X1 U551 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U552 ( .A1(data_in[5]), .A2(n842), .B1(n1102), .B2(\mem[1][5] ), 
        .ZN(n1097) );
  INV_X1 U553 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U554 ( .A1(data_in[6]), .A2(n842), .B1(n1102), .B2(\mem[1][6] ), 
        .ZN(n1096) );
  INV_X1 U555 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U556 ( .A1(data_in[7]), .A2(n842), .B1(n1102), .B2(\mem[1][7] ), 
        .ZN(n1095) );
  INV_X1 U557 ( .A(n1093), .ZN(n795) );
  AOI22_X1 U558 ( .A1(data_in[0]), .A2(n841), .B1(n1092), .B2(\mem[2][0] ), 
        .ZN(n1093) );
  INV_X1 U559 ( .A(n1091), .ZN(n794) );
  AOI22_X1 U560 ( .A1(data_in[1]), .A2(n841), .B1(n1092), .B2(\mem[2][1] ), 
        .ZN(n1091) );
  INV_X1 U561 ( .A(n1090), .ZN(n793) );
  AOI22_X1 U562 ( .A1(data_in[2]), .A2(n841), .B1(n1092), .B2(\mem[2][2] ), 
        .ZN(n1090) );
  INV_X1 U563 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U564 ( .A1(data_in[3]), .A2(n841), .B1(n1092), .B2(\mem[2][3] ), 
        .ZN(n1089) );
  INV_X1 U565 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U566 ( .A1(data_in[4]), .A2(n841), .B1(n1092), .B2(\mem[2][4] ), 
        .ZN(n1088) );
  INV_X1 U567 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U568 ( .A1(data_in[5]), .A2(n841), .B1(n1092), .B2(\mem[2][5] ), 
        .ZN(n1087) );
  INV_X1 U569 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U570 ( .A1(data_in[6]), .A2(n841), .B1(n1092), .B2(\mem[2][6] ), 
        .ZN(n1086) );
  INV_X1 U571 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U572 ( .A1(data_in[7]), .A2(n841), .B1(n1092), .B2(\mem[2][7] ), 
        .ZN(n1085) );
  INV_X1 U573 ( .A(n1083), .ZN(n787) );
  AOI22_X1 U574 ( .A1(data_in[0]), .A2(n840), .B1(n1082), .B2(\mem[3][0] ), 
        .ZN(n1083) );
  INV_X1 U575 ( .A(n1081), .ZN(n786) );
  AOI22_X1 U576 ( .A1(data_in[1]), .A2(n840), .B1(n1082), .B2(\mem[3][1] ), 
        .ZN(n1081) );
  INV_X1 U577 ( .A(n1080), .ZN(n785) );
  AOI22_X1 U578 ( .A1(data_in[2]), .A2(n840), .B1(n1082), .B2(\mem[3][2] ), 
        .ZN(n1080) );
  INV_X1 U579 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U580 ( .A1(data_in[3]), .A2(n840), .B1(n1082), .B2(\mem[3][3] ), 
        .ZN(n1079) );
  INV_X1 U581 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U582 ( .A1(data_in[4]), .A2(n840), .B1(n1082), .B2(\mem[3][4] ), 
        .ZN(n1078) );
  INV_X1 U583 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U584 ( .A1(data_in[5]), .A2(n840), .B1(n1082), .B2(\mem[3][5] ), 
        .ZN(n1077) );
  INV_X1 U585 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U586 ( .A1(data_in[6]), .A2(n840), .B1(n1082), .B2(\mem[3][6] ), 
        .ZN(n1076) );
  INV_X1 U587 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U588 ( .A1(data_in[7]), .A2(n840), .B1(n1082), .B2(\mem[3][7] ), 
        .ZN(n1075) );
  INV_X1 U589 ( .A(n1073), .ZN(n779) );
  AOI22_X1 U590 ( .A1(data_in[0]), .A2(n839), .B1(n1072), .B2(\mem[4][0] ), 
        .ZN(n1073) );
  INV_X1 U591 ( .A(n1071), .ZN(n778) );
  AOI22_X1 U592 ( .A1(data_in[1]), .A2(n839), .B1(n1072), .B2(\mem[4][1] ), 
        .ZN(n1071) );
  INV_X1 U593 ( .A(n1070), .ZN(n777) );
  AOI22_X1 U594 ( .A1(data_in[2]), .A2(n839), .B1(n1072), .B2(\mem[4][2] ), 
        .ZN(n1070) );
  INV_X1 U595 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U596 ( .A1(data_in[3]), .A2(n839), .B1(n1072), .B2(\mem[4][3] ), 
        .ZN(n1069) );
  INV_X1 U597 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U598 ( .A1(data_in[4]), .A2(n839), .B1(n1072), .B2(\mem[4][4] ), 
        .ZN(n1068) );
  INV_X1 U599 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U600 ( .A1(data_in[5]), .A2(n839), .B1(n1072), .B2(\mem[4][5] ), 
        .ZN(n1067) );
  INV_X1 U601 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U602 ( .A1(data_in[6]), .A2(n839), .B1(n1072), .B2(\mem[4][6] ), 
        .ZN(n1066) );
  INV_X1 U603 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U604 ( .A1(data_in[7]), .A2(n839), .B1(n1072), .B2(\mem[4][7] ), 
        .ZN(n1065) );
  INV_X1 U605 ( .A(N13), .ZN(n844) );
  INV_X1 U606 ( .A(N14), .ZN(n845) );
  MUX2_X1 U607 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n251), .Z(n3) );
  MUX2_X1 U608 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n251), .Z(n4) );
  MUX2_X1 U609 ( .A(n4), .B(n3), .S(n245), .Z(n5) );
  MUX2_X1 U610 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n251), .Z(n6) );
  MUX2_X1 U611 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n250), .Z(n7) );
  MUX2_X1 U612 ( .A(n7), .B(n6), .S(n245), .Z(n8) );
  MUX2_X1 U613 ( .A(n8), .B(n5), .S(n243), .Z(n9) );
  MUX2_X1 U614 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n251), .Z(n10) );
  MUX2_X1 U615 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n250), .Z(n11) );
  MUX2_X1 U616 ( .A(n11), .B(n10), .S(n246), .Z(n12) );
  MUX2_X1 U617 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n251), .Z(n13) );
  MUX2_X1 U618 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n250), .Z(n14) );
  MUX2_X1 U619 ( .A(n14), .B(n13), .S(n244), .Z(n15) );
  MUX2_X1 U620 ( .A(n15), .B(n12), .S(n243), .Z(n16) );
  MUX2_X1 U621 ( .A(n16), .B(n9), .S(N13), .Z(n17) );
  MUX2_X1 U622 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n247), .Z(n18) );
  MUX2_X1 U623 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n247), .Z(n19) );
  MUX2_X1 U624 ( .A(n19), .B(n18), .S(n244), .Z(n20) );
  MUX2_X1 U625 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n247), .Z(n21) );
  MUX2_X1 U626 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n247), .Z(n22) );
  MUX2_X1 U627 ( .A(n22), .B(n21), .S(n244), .Z(n23) );
  MUX2_X1 U628 ( .A(n23), .B(n20), .S(N12), .Z(n24) );
  MUX2_X1 U629 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n247), .Z(n25) );
  MUX2_X1 U630 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n247), .Z(n26) );
  MUX2_X1 U631 ( .A(n26), .B(n25), .S(n244), .Z(n27) );
  MUX2_X1 U632 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n247), .Z(n28) );
  MUX2_X1 U633 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n247), .Z(n29) );
  MUX2_X1 U634 ( .A(n29), .B(n28), .S(n244), .Z(n30) );
  MUX2_X1 U635 ( .A(n30), .B(n27), .S(N12), .Z(n31) );
  MUX2_X1 U636 ( .A(n31), .B(n24), .S(N13), .Z(n32) );
  MUX2_X1 U637 ( .A(n32), .B(n17), .S(N14), .Z(N22) );
  MUX2_X1 U638 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n247), .Z(n33) );
  MUX2_X1 U639 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n247), .Z(n34) );
  MUX2_X1 U640 ( .A(n34), .B(n33), .S(n244), .Z(n35) );
  MUX2_X1 U641 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n247), .Z(n36) );
  MUX2_X1 U642 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n247), .Z(n37) );
  MUX2_X1 U643 ( .A(n37), .B(n36), .S(n244), .Z(n38) );
  MUX2_X1 U644 ( .A(n38), .B(n35), .S(n243), .Z(n39) );
  MUX2_X1 U645 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n248), .Z(n40) );
  MUX2_X1 U646 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n248), .Z(n41) );
  MUX2_X1 U647 ( .A(n41), .B(n40), .S(n244), .Z(n42) );
  MUX2_X1 U648 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n248), .Z(n43) );
  MUX2_X1 U649 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n248), .Z(n44) );
  MUX2_X1 U650 ( .A(n44), .B(n43), .S(n244), .Z(n45) );
  MUX2_X1 U651 ( .A(n45), .B(n42), .S(n243), .Z(n46) );
  MUX2_X1 U652 ( .A(n46), .B(n39), .S(N13), .Z(n47) );
  MUX2_X1 U653 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n248), .Z(n48) );
  MUX2_X1 U654 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n248), .Z(n49) );
  MUX2_X1 U655 ( .A(n49), .B(n48), .S(n244), .Z(n50) );
  MUX2_X1 U656 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n248), .Z(n51) );
  MUX2_X1 U657 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n248), .Z(n52) );
  MUX2_X1 U658 ( .A(n52), .B(n51), .S(n244), .Z(n53) );
  MUX2_X1 U659 ( .A(n53), .B(n50), .S(n243), .Z(n54) );
  MUX2_X1 U660 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n248), .Z(n55) );
  MUX2_X1 U661 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n248), .Z(n56) );
  MUX2_X1 U662 ( .A(n56), .B(n55), .S(n244), .Z(n57) );
  MUX2_X1 U663 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n248), .Z(n58) );
  MUX2_X1 U664 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n248), .Z(n59) );
  MUX2_X1 U665 ( .A(n59), .B(n58), .S(n244), .Z(n60) );
  MUX2_X1 U666 ( .A(n60), .B(n57), .S(n243), .Z(n61) );
  MUX2_X1 U667 ( .A(n61), .B(n54), .S(N13), .Z(n62) );
  MUX2_X1 U668 ( .A(n62), .B(n47), .S(N14), .Z(N21) );
  MUX2_X1 U669 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n249), .Z(n63) );
  MUX2_X1 U670 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n249), .Z(n64) );
  MUX2_X1 U671 ( .A(n64), .B(n63), .S(n245), .Z(n65) );
  MUX2_X1 U672 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n249), .Z(n66) );
  MUX2_X1 U673 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n249), .Z(n67) );
  MUX2_X1 U674 ( .A(n67), .B(n66), .S(n245), .Z(n68) );
  MUX2_X1 U675 ( .A(n68), .B(n65), .S(n243), .Z(n69) );
  MUX2_X1 U676 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n249), .Z(n70) );
  MUX2_X1 U677 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n249), .Z(n71) );
  MUX2_X1 U678 ( .A(n71), .B(n70), .S(n245), .Z(n72) );
  MUX2_X1 U679 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n249), .Z(n73) );
  MUX2_X1 U680 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n249), .Z(n74) );
  MUX2_X1 U681 ( .A(n74), .B(n73), .S(n245), .Z(n75) );
  MUX2_X1 U682 ( .A(n75), .B(n72), .S(n243), .Z(n76) );
  MUX2_X1 U683 ( .A(n76), .B(n69), .S(N13), .Z(n77) );
  MUX2_X1 U684 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n249), .Z(n78) );
  MUX2_X1 U685 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n249), .Z(n79) );
  MUX2_X1 U686 ( .A(n79), .B(n78), .S(n245), .Z(n80) );
  MUX2_X1 U687 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n249), .Z(n81) );
  MUX2_X1 U688 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n249), .Z(n82) );
  MUX2_X1 U689 ( .A(n82), .B(n81), .S(n245), .Z(n83) );
  MUX2_X1 U690 ( .A(n83), .B(n80), .S(n243), .Z(n84) );
  MUX2_X1 U691 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n252), .Z(n85) );
  MUX2_X1 U692 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n249), .Z(n86) );
  MUX2_X1 U693 ( .A(n86), .B(n85), .S(n245), .Z(n87) );
  MUX2_X1 U694 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n247), .Z(n88) );
  MUX2_X1 U695 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n248), .Z(n89) );
  MUX2_X1 U696 ( .A(n89), .B(n88), .S(n245), .Z(n90) );
  MUX2_X1 U697 ( .A(n90), .B(n87), .S(n243), .Z(n91) );
  MUX2_X1 U698 ( .A(n91), .B(n84), .S(N13), .Z(n92) );
  MUX2_X1 U699 ( .A(n92), .B(n77), .S(N14), .Z(N20) );
  MUX2_X1 U700 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n248), .Z(n93) );
  MUX2_X1 U701 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n252), .Z(n94) );
  MUX2_X1 U702 ( .A(n94), .B(n93), .S(n245), .Z(n95) );
  MUX2_X1 U703 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n247), .Z(n96) );
  MUX2_X1 U704 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n250), .Z(n97) );
  MUX2_X1 U705 ( .A(n97), .B(n96), .S(n245), .Z(n98) );
  MUX2_X1 U706 ( .A(n98), .B(n95), .S(n243), .Z(n99) );
  MUX2_X1 U707 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n252), .Z(n100) );
  MUX2_X1 U708 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n248), .Z(n101) );
  MUX2_X1 U709 ( .A(n101), .B(n100), .S(n245), .Z(n102) );
  MUX2_X1 U710 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n249), .Z(n103) );
  MUX2_X1 U711 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n250), .Z(n104) );
  MUX2_X1 U712 ( .A(n104), .B(n103), .S(n245), .Z(n105) );
  MUX2_X1 U713 ( .A(n105), .B(n102), .S(n243), .Z(n106) );
  MUX2_X1 U714 ( .A(n106), .B(n99), .S(N13), .Z(n107) );
  MUX2_X1 U715 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n251), .Z(n108) );
  MUX2_X1 U716 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n252), .Z(n109) );
  MUX2_X1 U717 ( .A(n109), .B(n108), .S(n246), .Z(n110) );
  MUX2_X1 U718 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n251), .Z(n111) );
  MUX2_X1 U719 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(N10), .Z(n112) );
  MUX2_X1 U720 ( .A(n112), .B(n111), .S(n246), .Z(n113) );
  MUX2_X1 U721 ( .A(n113), .B(n110), .S(n243), .Z(n114) );
  MUX2_X1 U722 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n252), .Z(n115) );
  MUX2_X1 U723 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(N10), .Z(n116) );
  MUX2_X1 U724 ( .A(n116), .B(n115), .S(n246), .Z(n117) );
  MUX2_X1 U725 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(N10), .Z(n118) );
  MUX2_X1 U726 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(N10), .Z(n119) );
  MUX2_X1 U727 ( .A(n119), .B(n118), .S(n246), .Z(n120) );
  MUX2_X1 U728 ( .A(n120), .B(n117), .S(n243), .Z(n121) );
  MUX2_X1 U729 ( .A(n121), .B(n114), .S(N13), .Z(n122) );
  MUX2_X1 U730 ( .A(n122), .B(n107), .S(N14), .Z(N19) );
  MUX2_X1 U731 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n251), .Z(n123) );
  MUX2_X1 U732 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(N10), .Z(n124) );
  MUX2_X1 U733 ( .A(n124), .B(n123), .S(n246), .Z(n125) );
  MUX2_X1 U734 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n251), .Z(n126) );
  MUX2_X1 U735 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(N10), .Z(n127) );
  MUX2_X1 U736 ( .A(n127), .B(n126), .S(n246), .Z(n128) );
  MUX2_X1 U737 ( .A(n128), .B(n125), .S(n243), .Z(n129) );
  MUX2_X1 U738 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n250), .Z(n130) );
  MUX2_X1 U739 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n250), .Z(n131) );
  MUX2_X1 U740 ( .A(n131), .B(n130), .S(n246), .Z(n132) );
  MUX2_X1 U741 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n250), .Z(n133) );
  MUX2_X1 U742 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n250), .Z(n134) );
  MUX2_X1 U743 ( .A(n134), .B(n133), .S(n246), .Z(n135) );
  MUX2_X1 U744 ( .A(n135), .B(n132), .S(n243), .Z(n136) );
  MUX2_X1 U745 ( .A(n136), .B(n129), .S(N13), .Z(n137) );
  MUX2_X1 U746 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n250), .Z(n138) );
  MUX2_X1 U747 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n250), .Z(n139) );
  MUX2_X1 U748 ( .A(n139), .B(n138), .S(n246), .Z(n140) );
  MUX2_X1 U749 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n250), .Z(n141) );
  MUX2_X1 U750 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n250), .Z(n142) );
  MUX2_X1 U751 ( .A(n142), .B(n141), .S(n246), .Z(n143) );
  MUX2_X1 U752 ( .A(n143), .B(n140), .S(n243), .Z(n144) );
  MUX2_X1 U753 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n250), .Z(n145) );
  MUX2_X1 U754 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n250), .Z(n146) );
  MUX2_X1 U755 ( .A(n146), .B(n145), .S(n246), .Z(n147) );
  MUX2_X1 U756 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n250), .Z(n148) );
  MUX2_X1 U757 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n250), .Z(n149) );
  MUX2_X1 U758 ( .A(n149), .B(n148), .S(n246), .Z(n150) );
  MUX2_X1 U759 ( .A(n150), .B(n147), .S(n243), .Z(n151) );
  MUX2_X1 U760 ( .A(n151), .B(n144), .S(N13), .Z(n152) );
  MUX2_X1 U761 ( .A(n152), .B(n137), .S(N14), .Z(N18) );
  MUX2_X1 U762 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n251), .Z(n153) );
  MUX2_X1 U763 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n251), .Z(n154) );
  MUX2_X1 U764 ( .A(n154), .B(n153), .S(N11), .Z(n155) );
  MUX2_X1 U765 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n251), .Z(n156) );
  MUX2_X1 U766 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n251), .Z(n157) );
  MUX2_X1 U767 ( .A(n157), .B(n156), .S(N11), .Z(n158) );
  MUX2_X1 U768 ( .A(n158), .B(n155), .S(n243), .Z(n159) );
  MUX2_X1 U769 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n251), .Z(n160) );
  MUX2_X1 U770 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n251), .Z(n161) );
  MUX2_X1 U771 ( .A(n161), .B(n160), .S(N11), .Z(n162) );
  MUX2_X1 U772 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n251), .Z(n163) );
  MUX2_X1 U773 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n251), .Z(n164) );
  MUX2_X1 U774 ( .A(n164), .B(n163), .S(N11), .Z(n165) );
  MUX2_X1 U775 ( .A(n165), .B(n162), .S(n243), .Z(n166) );
  MUX2_X1 U776 ( .A(n166), .B(n159), .S(N13), .Z(n167) );
  MUX2_X1 U777 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n251), .Z(n168) );
  MUX2_X1 U778 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n251), .Z(n169) );
  MUX2_X1 U779 ( .A(n169), .B(n168), .S(N11), .Z(n170) );
  MUX2_X1 U780 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n251), .Z(n171) );
  MUX2_X1 U781 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n251), .Z(n172) );
  MUX2_X1 U782 ( .A(n172), .B(n171), .S(N11), .Z(n173) );
  MUX2_X1 U783 ( .A(n173), .B(n170), .S(n243), .Z(n174) );
  MUX2_X1 U784 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n248), .Z(n175) );
  MUX2_X1 U785 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n252), .Z(n176) );
  MUX2_X1 U786 ( .A(n176), .B(n175), .S(N11), .Z(n177) );
  MUX2_X1 U787 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n247), .Z(n178) );
  MUX2_X1 U788 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n251), .Z(n179) );
  MUX2_X1 U789 ( .A(n179), .B(n178), .S(N11), .Z(n180) );
  MUX2_X1 U790 ( .A(n180), .B(n177), .S(n243), .Z(n181) );
  MUX2_X1 U791 ( .A(n181), .B(n174), .S(N13), .Z(n182) );
  MUX2_X1 U792 ( .A(n182), .B(n167), .S(N14), .Z(N17) );
  MUX2_X1 U793 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n249), .Z(n183) );
  MUX2_X1 U794 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n252), .Z(n184) );
  MUX2_X1 U795 ( .A(n184), .B(n183), .S(N11), .Z(n185) );
  MUX2_X1 U796 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n252), .Z(n186) );
  MUX2_X1 U797 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n252), .Z(n187) );
  MUX2_X1 U798 ( .A(n187), .B(n186), .S(n245), .Z(n188) );
  MUX2_X1 U799 ( .A(n188), .B(n185), .S(n243), .Z(n189) );
  MUX2_X1 U800 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n248), .Z(n190) );
  MUX2_X1 U801 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n252), .Z(n191) );
  MUX2_X1 U802 ( .A(n191), .B(n190), .S(n246), .Z(n192) );
  MUX2_X1 U803 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n252), .Z(n193) );
  MUX2_X1 U804 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n252), .Z(n194) );
  MUX2_X1 U805 ( .A(n194), .B(n193), .S(n244), .Z(n195) );
  MUX2_X1 U806 ( .A(n195), .B(n192), .S(N12), .Z(n196) );
  MUX2_X1 U807 ( .A(n196), .B(n189), .S(N13), .Z(n197) );
  MUX2_X1 U808 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n249), .Z(n198) );
  MUX2_X1 U809 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(N10), .Z(n199) );
  MUX2_X1 U810 ( .A(n199), .B(n198), .S(n245), .Z(n200) );
  MUX2_X1 U811 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n249), .Z(n201) );
  MUX2_X1 U812 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n252), .Z(n202) );
  MUX2_X1 U813 ( .A(n202), .B(n201), .S(n244), .Z(n203) );
  MUX2_X1 U814 ( .A(n203), .B(n200), .S(N12), .Z(n204) );
  MUX2_X1 U815 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n251), .Z(n205) );
  MUX2_X1 U816 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n252), .Z(n206) );
  MUX2_X1 U817 ( .A(n206), .B(n205), .S(n246), .Z(n207) );
  MUX2_X1 U818 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n208) );
  MUX2_X1 U819 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n252), .Z(n209) );
  MUX2_X1 U820 ( .A(n209), .B(n208), .S(N11), .Z(n210) );
  MUX2_X1 U821 ( .A(n210), .B(n207), .S(N12), .Z(n211) );
  MUX2_X1 U822 ( .A(n211), .B(n204), .S(N13), .Z(n212) );
  MUX2_X1 U823 ( .A(n212), .B(n197), .S(N14), .Z(N16) );
  MUX2_X1 U824 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n250), .Z(n213) );
  MUX2_X1 U825 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n252), .Z(n214) );
  MUX2_X1 U826 ( .A(n214), .B(n213), .S(n245), .Z(n215) );
  MUX2_X1 U827 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n252), .Z(n216) );
  MUX2_X1 U828 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(N10), .Z(n217) );
  MUX2_X1 U829 ( .A(n217), .B(n216), .S(n244), .Z(n218) );
  MUX2_X1 U830 ( .A(n218), .B(n215), .S(N12), .Z(n219) );
  MUX2_X1 U831 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n249), .Z(n220) );
  MUX2_X1 U832 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n252), .Z(n221) );
  MUX2_X1 U833 ( .A(n221), .B(n220), .S(n244), .Z(n222) );
  MUX2_X1 U834 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n247), .Z(n223) );
  MUX2_X1 U835 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n224) );
  MUX2_X1 U836 ( .A(n224), .B(n223), .S(N11), .Z(n225) );
  MUX2_X1 U837 ( .A(n225), .B(n222), .S(N12), .Z(n226) );
  MUX2_X1 U838 ( .A(n226), .B(n219), .S(N13), .Z(n227) );
  MUX2_X1 U839 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n247), .Z(n228) );
  MUX2_X1 U840 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n252), .Z(n229) );
  MUX2_X1 U841 ( .A(n229), .B(n228), .S(n246), .Z(n230) );
  MUX2_X1 U842 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n252), .Z(n231) );
  MUX2_X1 U843 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n232) );
  MUX2_X1 U844 ( .A(n232), .B(n231), .S(N11), .Z(n233) );
  MUX2_X1 U845 ( .A(n233), .B(n230), .S(N12), .Z(n234) );
  MUX2_X1 U846 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n248), .Z(n235) );
  MUX2_X1 U847 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n236) );
  MUX2_X1 U848 ( .A(n236), .B(n235), .S(n246), .Z(n237) );
  MUX2_X1 U849 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n238) );
  MUX2_X1 U850 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n239) );
  MUX2_X1 U851 ( .A(n239), .B(n238), .S(N11), .Z(n240) );
  MUX2_X1 U852 ( .A(n240), .B(n237), .S(N12), .Z(n241) );
  MUX2_X1 U853 ( .A(n241), .B(n234), .S(N13), .Z(n242) );
  MUX2_X1 U854 ( .A(n242), .B(n227), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_2 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X2 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  BUF_X1 U3 ( .A(N10), .Z(n247) );
  BUF_X1 U4 ( .A(n250), .Z(n248) );
  BUF_X1 U5 ( .A(n250), .Z(n249) );
  BUF_X1 U6 ( .A(n250), .Z(n245) );
  BUF_X1 U7 ( .A(n250), .Z(n246) );
  BUF_X1 U8 ( .A(N10), .Z(n250) );
  INV_X1 U9 ( .A(n1111), .ZN(n841) );
  INV_X1 U10 ( .A(n1100), .ZN(n840) );
  INV_X1 U11 ( .A(n1090), .ZN(n839) );
  INV_X1 U12 ( .A(n1080), .ZN(n838) );
  INV_X1 U13 ( .A(n1070), .ZN(n837) );
  INV_X1 U14 ( .A(n1060), .ZN(n836) );
  INV_X1 U15 ( .A(n1051), .ZN(n835) );
  INV_X1 U16 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U18 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U19 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U20 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U21 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U22 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U23 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U24 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U26 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U27 ( .A(n1131), .ZN(n816) );
  INV_X1 U28 ( .A(n1121), .ZN(n815) );
  INV_X1 U29 ( .A(n887), .ZN(n814) );
  INV_X1 U30 ( .A(n878), .ZN(n813) );
  INV_X1 U31 ( .A(n869), .ZN(n812) );
  INV_X1 U32 ( .A(n860), .ZN(n811) );
  INV_X1 U33 ( .A(n851), .ZN(n810) );
  INV_X1 U34 ( .A(n987), .ZN(n828) );
  INV_X1 U35 ( .A(n978), .ZN(n827) );
  INV_X1 U36 ( .A(n969), .ZN(n826) );
  INV_X1 U37 ( .A(n914), .ZN(n820) );
  INV_X1 U38 ( .A(n905), .ZN(n819) );
  INV_X1 U39 ( .A(n896), .ZN(n818) );
  INV_X1 U40 ( .A(n1033), .ZN(n833) );
  INV_X1 U41 ( .A(n1023), .ZN(n832) );
  INV_X1 U42 ( .A(n1014), .ZN(n831) );
  INV_X1 U43 ( .A(n1005), .ZN(n830) );
  INV_X1 U44 ( .A(n996), .ZN(n829) );
  INV_X1 U45 ( .A(n960), .ZN(n825) );
  INV_X1 U46 ( .A(n950), .ZN(n824) );
  INV_X1 U47 ( .A(n941), .ZN(n823) );
  INV_X1 U48 ( .A(n932), .ZN(n822) );
  INV_X1 U49 ( .A(n923), .ZN(n821) );
  INV_X1 U50 ( .A(n1142), .ZN(n817) );
  BUF_X1 U51 ( .A(N11), .Z(n242) );
  BUF_X1 U52 ( .A(N11), .Z(n243) );
  BUF_X1 U53 ( .A(N11), .Z(n244) );
  INV_X1 U54 ( .A(N10), .ZN(n251) );
  BUF_X1 U55 ( .A(N12), .Z(n241) );
  NOR3_X1 U56 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U57 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U58 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U59 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U60 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U61 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U62 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U63 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U64 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U65 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U67 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U69 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U70 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U71 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U72 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U73 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U74 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U75 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U76 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U77 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U79 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U81 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U82 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U83 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U84 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U85 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U86 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U87 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U88 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U89 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U90 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U91 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U92 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U93 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U94 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U95 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U96 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U97 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U98 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U99 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U100 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U101 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U102 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U103 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U104 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U105 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U106 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U107 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U108 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U109 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U110 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U111 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U112 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U113 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U114 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U115 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U116 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U117 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U118 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U119 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U120 ( .A(n988), .ZN(n705) );
  AOI22_X1 U121 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U122 ( .A(n986), .ZN(n704) );
  AOI22_X1 U123 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U124 ( .A(n984), .ZN(n702) );
  AOI22_X1 U125 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U126 ( .A(n983), .ZN(n701) );
  AOI22_X1 U127 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U128 ( .A(n951), .ZN(n673) );
  AOI22_X1 U129 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U130 ( .A(n947), .ZN(n670) );
  AOI22_X1 U131 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U132 ( .A(n946), .ZN(n669) );
  AOI22_X1 U133 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U134 ( .A(n913), .ZN(n640) );
  AOI22_X1 U135 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U136 ( .A(n911), .ZN(n638) );
  AOI22_X1 U137 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U138 ( .A(n910), .ZN(n637) );
  AOI22_X1 U139 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U140 ( .A(n909), .ZN(n636) );
  AOI22_X1 U141 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U142 ( .A(n908), .ZN(n635) );
  AOI22_X1 U143 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U144 ( .A(n907), .ZN(n634) );
  AOI22_X1 U145 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U146 ( .A(n985), .ZN(n703) );
  AOI22_X1 U147 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U148 ( .A(n982), .ZN(n700) );
  AOI22_X1 U149 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U150 ( .A(n981), .ZN(n699) );
  AOI22_X1 U151 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U152 ( .A(n980), .ZN(n698) );
  AOI22_X1 U153 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U154 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U155 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U156 ( .A(n948), .ZN(n671) );
  AOI22_X1 U157 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U158 ( .A(n945), .ZN(n668) );
  AOI22_X1 U159 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U160 ( .A(n944), .ZN(n667) );
  AOI22_X1 U161 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U162 ( .A(n943), .ZN(n666) );
  AOI22_X1 U163 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U164 ( .A(n915), .ZN(n641) );
  AOI22_X1 U165 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U166 ( .A(n949), .ZN(n672) );
  AOI22_X1 U167 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U168 ( .A(n912), .ZN(n639) );
  AOI22_X1 U169 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U170 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U171 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U172 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U173 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U174 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U175 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U176 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U177 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U178 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U179 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U180 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U181 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U182 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U183 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U184 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U185 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U186 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U187 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U188 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U189 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U190 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U191 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U192 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U193 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U194 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U195 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U196 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U197 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U198 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U199 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U200 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U201 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U202 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U203 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U204 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U205 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U206 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U207 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U208 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U209 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U210 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U211 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U212 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U213 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U214 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U215 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U216 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U217 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U218 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U219 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U220 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U221 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U222 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U223 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U224 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U225 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U226 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U227 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U228 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U229 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U230 ( .A(n999), .ZN(n715) );
  AOI22_X1 U231 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U232 ( .A(n998), .ZN(n714) );
  AOI22_X1 U233 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U234 ( .A(n979), .ZN(n697) );
  AOI22_X1 U235 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U236 ( .A(n977), .ZN(n696) );
  AOI22_X1 U237 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U238 ( .A(n976), .ZN(n695) );
  AOI22_X1 U239 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U240 ( .A(n975), .ZN(n694) );
  AOI22_X1 U241 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U242 ( .A(n974), .ZN(n693) );
  AOI22_X1 U243 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U244 ( .A(n973), .ZN(n692) );
  AOI22_X1 U245 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U246 ( .A(n972), .ZN(n691) );
  AOI22_X1 U247 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U248 ( .A(n971), .ZN(n690) );
  AOI22_X1 U249 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U250 ( .A(n970), .ZN(n689) );
  AOI22_X1 U251 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U252 ( .A(n968), .ZN(n688) );
  AOI22_X1 U253 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U254 ( .A(n967), .ZN(n687) );
  AOI22_X1 U255 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U256 ( .A(n966), .ZN(n686) );
  AOI22_X1 U257 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U258 ( .A(n965), .ZN(n685) );
  AOI22_X1 U259 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U260 ( .A(n964), .ZN(n684) );
  AOI22_X1 U261 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U262 ( .A(n963), .ZN(n683) );
  AOI22_X1 U263 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U264 ( .A(n962), .ZN(n682) );
  AOI22_X1 U265 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U266 ( .A(n942), .ZN(n665) );
  AOI22_X1 U267 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U268 ( .A(n940), .ZN(n664) );
  AOI22_X1 U269 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U270 ( .A(n939), .ZN(n663) );
  AOI22_X1 U271 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U272 ( .A(n938), .ZN(n662) );
  AOI22_X1 U273 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U274 ( .A(n937), .ZN(n661) );
  AOI22_X1 U275 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U276 ( .A(n936), .ZN(n660) );
  AOI22_X1 U277 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U278 ( .A(n935), .ZN(n659) );
  AOI22_X1 U279 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U280 ( .A(n934), .ZN(n658) );
  AOI22_X1 U281 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U282 ( .A(n933), .ZN(n657) );
  AOI22_X1 U283 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U284 ( .A(n931), .ZN(n656) );
  AOI22_X1 U285 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U286 ( .A(n930), .ZN(n655) );
  AOI22_X1 U287 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U288 ( .A(n929), .ZN(n654) );
  AOI22_X1 U289 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U290 ( .A(n928), .ZN(n653) );
  AOI22_X1 U291 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U292 ( .A(n927), .ZN(n652) );
  AOI22_X1 U293 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U294 ( .A(n926), .ZN(n651) );
  AOI22_X1 U295 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U296 ( .A(n925), .ZN(n650) );
  AOI22_X1 U297 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U298 ( .A(n906), .ZN(n633) );
  AOI22_X1 U299 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U300 ( .A(n904), .ZN(n632) );
  AOI22_X1 U301 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U302 ( .A(n903), .ZN(n631) );
  AOI22_X1 U303 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U304 ( .A(n902), .ZN(n630) );
  AOI22_X1 U305 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U306 ( .A(n901), .ZN(n629) );
  AOI22_X1 U307 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U308 ( .A(n900), .ZN(n628) );
  AOI22_X1 U309 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U310 ( .A(n899), .ZN(n627) );
  AOI22_X1 U311 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U312 ( .A(n898), .ZN(n626) );
  AOI22_X1 U313 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U314 ( .A(n897), .ZN(n625) );
  AOI22_X1 U315 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U316 ( .A(n895), .ZN(n624) );
  AOI22_X1 U317 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U318 ( .A(n894), .ZN(n623) );
  AOI22_X1 U319 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U320 ( .A(n893), .ZN(n622) );
  AOI22_X1 U321 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U322 ( .A(n892), .ZN(n621) );
  AOI22_X1 U323 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U324 ( .A(n891), .ZN(n620) );
  AOI22_X1 U325 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U326 ( .A(n890), .ZN(n619) );
  AOI22_X1 U327 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U328 ( .A(n889), .ZN(n618) );
  AOI22_X1 U329 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U330 ( .A(N12), .ZN(n253) );
  INV_X1 U331 ( .A(N11), .ZN(n252) );
  INV_X1 U332 ( .A(n997), .ZN(n713) );
  AOI22_X1 U333 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U334 ( .A(n995), .ZN(n712) );
  AOI22_X1 U335 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U336 ( .A(n994), .ZN(n711) );
  AOI22_X1 U337 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U338 ( .A(n993), .ZN(n710) );
  AOI22_X1 U339 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U340 ( .A(n992), .ZN(n709) );
  AOI22_X1 U341 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U342 ( .A(n991), .ZN(n708) );
  AOI22_X1 U343 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U344 ( .A(n990), .ZN(n707) );
  AOI22_X1 U345 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U346 ( .A(n989), .ZN(n706) );
  AOI22_X1 U347 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U348 ( .A(n924), .ZN(n649) );
  AOI22_X1 U349 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U350 ( .A(n922), .ZN(n648) );
  AOI22_X1 U351 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U352 ( .A(n921), .ZN(n647) );
  AOI22_X1 U353 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U354 ( .A(n920), .ZN(n646) );
  AOI22_X1 U355 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U356 ( .A(n919), .ZN(n645) );
  AOI22_X1 U357 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U358 ( .A(n918), .ZN(n644) );
  AOI22_X1 U359 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U360 ( .A(n917), .ZN(n643) );
  AOI22_X1 U361 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U362 ( .A(n916), .ZN(n642) );
  AOI22_X1 U363 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U364 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U365 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U366 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U367 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U368 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U369 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U370 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U371 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U372 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U373 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U374 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U375 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U376 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U377 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U378 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U379 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U380 ( .A(n961), .ZN(n681) );
  AOI22_X1 U381 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U382 ( .A(n959), .ZN(n680) );
  AOI22_X1 U383 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U384 ( .A(n958), .ZN(n679) );
  AOI22_X1 U385 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U386 ( .A(n957), .ZN(n678) );
  AOI22_X1 U387 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U388 ( .A(n956), .ZN(n677) );
  AOI22_X1 U389 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U390 ( .A(n955), .ZN(n676) );
  AOI22_X1 U391 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U392 ( .A(n954), .ZN(n675) );
  AOI22_X1 U393 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U394 ( .A(n953), .ZN(n674) );
  AOI22_X1 U395 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U396 ( .A(n888), .ZN(n617) );
  AOI22_X1 U397 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U398 ( .A(n886), .ZN(n616) );
  AOI22_X1 U399 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U400 ( .A(n885), .ZN(n615) );
  AOI22_X1 U401 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U402 ( .A(n884), .ZN(n614) );
  AOI22_X1 U403 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U404 ( .A(n883), .ZN(n613) );
  AOI22_X1 U405 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U406 ( .A(n882), .ZN(n612) );
  AOI22_X1 U407 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U408 ( .A(n881), .ZN(n611) );
  AOI22_X1 U409 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U410 ( .A(n880), .ZN(n610) );
  AOI22_X1 U411 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U412 ( .A(n879), .ZN(n609) );
  AOI22_X1 U413 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U414 ( .A(n877), .ZN(n608) );
  AOI22_X1 U415 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U416 ( .A(n876), .ZN(n607) );
  AOI22_X1 U417 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U418 ( .A(n875), .ZN(n606) );
  AOI22_X1 U419 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U420 ( .A(n874), .ZN(n605) );
  AOI22_X1 U421 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U422 ( .A(n873), .ZN(n604) );
  AOI22_X1 U423 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U424 ( .A(n872), .ZN(n603) );
  AOI22_X1 U425 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U426 ( .A(n871), .ZN(n602) );
  AOI22_X1 U427 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U428 ( .A(n870), .ZN(n601) );
  AOI22_X1 U429 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U430 ( .A(n868), .ZN(n600) );
  AOI22_X1 U431 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U432 ( .A(n867), .ZN(n599) );
  AOI22_X1 U433 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U434 ( .A(n866), .ZN(n598) );
  AOI22_X1 U435 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U436 ( .A(n865), .ZN(n597) );
  AOI22_X1 U437 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U438 ( .A(n864), .ZN(n596) );
  AOI22_X1 U439 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U440 ( .A(n863), .ZN(n595) );
  AOI22_X1 U441 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U442 ( .A(n862), .ZN(n594) );
  AOI22_X1 U443 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U444 ( .A(n861), .ZN(n293) );
  AOI22_X1 U445 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U446 ( .A(n859), .ZN(n292) );
  AOI22_X1 U447 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U448 ( .A(n858), .ZN(n291) );
  AOI22_X1 U449 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U450 ( .A(n857), .ZN(n290) );
  AOI22_X1 U451 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U452 ( .A(n856), .ZN(n289) );
  AOI22_X1 U453 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U454 ( .A(n855), .ZN(n288) );
  AOI22_X1 U455 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U456 ( .A(n854), .ZN(n287) );
  AOI22_X1 U457 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U458 ( .A(n853), .ZN(n286) );
  AOI22_X1 U459 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U460 ( .A(n852), .ZN(n285) );
  AOI22_X1 U461 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U462 ( .A(n850), .ZN(n284) );
  AOI22_X1 U463 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U464 ( .A(n849), .ZN(n283) );
  AOI22_X1 U465 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U466 ( .A(n848), .ZN(n282) );
  AOI22_X1 U467 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U468 ( .A(n847), .ZN(n281) );
  AOI22_X1 U469 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U470 ( .A(n846), .ZN(n280) );
  AOI22_X1 U471 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U472 ( .A(n845), .ZN(n279) );
  AOI22_X1 U473 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U474 ( .A(n844), .ZN(n278) );
  AOI22_X1 U475 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U476 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U477 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U478 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U479 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U480 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U481 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U482 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U483 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U484 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U485 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U486 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U487 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U488 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U489 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U490 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U491 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U492 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U493 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U494 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U495 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U496 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U497 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U498 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U499 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U500 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U501 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U502 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U503 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U504 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U505 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U506 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U507 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U508 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U509 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U510 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U511 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U512 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U513 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U514 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U515 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U516 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U517 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U518 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U519 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U520 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U521 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U522 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U523 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U524 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U525 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U526 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U527 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U528 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U529 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U530 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U531 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U532 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U533 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U534 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U535 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U536 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U537 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U538 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U539 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U540 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U541 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U542 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U543 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U544 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U545 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U546 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U547 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U548 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U549 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U550 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U551 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U552 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U553 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U554 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U555 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U556 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U557 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U558 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U559 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U560 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U561 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U562 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U563 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U564 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U565 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U566 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U567 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U568 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U569 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U570 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U571 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U572 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U573 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U574 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U575 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U576 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U577 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U578 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U579 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U580 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U581 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U582 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U583 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U584 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U585 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U586 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U587 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U588 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U589 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U590 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U591 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U592 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U593 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U594 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U595 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U596 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U597 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U598 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U599 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U600 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U601 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U602 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U603 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U604 ( .A(N13), .ZN(n842) );
  INV_X1 U605 ( .A(N14), .ZN(n843) );
  MUX2_X1 U606 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n247), .Z(n1) );
  MUX2_X1 U607 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n247), .Z(n2) );
  MUX2_X1 U608 ( .A(n2), .B(n1), .S(N11), .Z(n3) );
  MUX2_X1 U609 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n247), .Z(n4) );
  MUX2_X1 U610 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n247), .Z(n5) );
  MUX2_X1 U611 ( .A(n5), .B(n4), .S(n244), .Z(n6) );
  MUX2_X1 U612 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U613 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n247), .Z(n8) );
  MUX2_X1 U614 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n249), .Z(n9) );
  MUX2_X1 U615 ( .A(n9), .B(n8), .S(n242), .Z(n10) );
  MUX2_X1 U616 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n247), .Z(n11) );
  MUX2_X1 U617 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n248), .Z(n12) );
  MUX2_X1 U618 ( .A(n12), .B(n11), .S(n242), .Z(n13) );
  MUX2_X1 U619 ( .A(n13), .B(n10), .S(N12), .Z(n14) );
  MUX2_X1 U620 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U621 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n245), .Z(n16) );
  MUX2_X1 U622 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n245), .Z(n17) );
  MUX2_X1 U623 ( .A(n17), .B(n16), .S(n242), .Z(n18) );
  MUX2_X1 U624 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n245), .Z(n19) );
  MUX2_X1 U625 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n245), .Z(n20) );
  MUX2_X1 U626 ( .A(n20), .B(n19), .S(n242), .Z(n21) );
  MUX2_X1 U627 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U628 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n245), .Z(n23) );
  MUX2_X1 U629 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n245), .Z(n24) );
  MUX2_X1 U630 ( .A(n24), .B(n23), .S(n242), .Z(n25) );
  MUX2_X1 U631 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n245), .Z(n26) );
  MUX2_X1 U632 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n245), .Z(n27) );
  MUX2_X1 U633 ( .A(n27), .B(n26), .S(n242), .Z(n28) );
  MUX2_X1 U634 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U635 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U636 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U637 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n245), .Z(n31) );
  MUX2_X1 U638 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n245), .Z(n32) );
  MUX2_X1 U639 ( .A(n32), .B(n31), .S(n242), .Z(n33) );
  MUX2_X1 U640 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n245), .Z(n34) );
  MUX2_X1 U641 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n245), .Z(n35) );
  MUX2_X1 U642 ( .A(n35), .B(n34), .S(n242), .Z(n36) );
  MUX2_X1 U643 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U644 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n246), .Z(n38) );
  MUX2_X1 U645 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n246), .Z(n39) );
  MUX2_X1 U646 ( .A(n39), .B(n38), .S(n242), .Z(n40) );
  MUX2_X1 U647 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n246), .Z(n41) );
  MUX2_X1 U648 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n246), .Z(n42) );
  MUX2_X1 U649 ( .A(n42), .B(n41), .S(n242), .Z(n43) );
  MUX2_X1 U650 ( .A(n43), .B(n40), .S(n241), .Z(n44) );
  MUX2_X1 U651 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U652 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n246), .Z(n46) );
  MUX2_X1 U653 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n246), .Z(n47) );
  MUX2_X1 U654 ( .A(n47), .B(n46), .S(n242), .Z(n48) );
  MUX2_X1 U655 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n246), .Z(n49) );
  MUX2_X1 U656 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n246), .Z(n50) );
  MUX2_X1 U657 ( .A(n50), .B(n49), .S(n242), .Z(n51) );
  MUX2_X1 U658 ( .A(n51), .B(n48), .S(n241), .Z(n52) );
  MUX2_X1 U659 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n246), .Z(n53) );
  MUX2_X1 U660 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n246), .Z(n54) );
  MUX2_X1 U661 ( .A(n54), .B(n53), .S(n242), .Z(n55) );
  MUX2_X1 U662 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n246), .Z(n56) );
  MUX2_X1 U663 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n246), .Z(n57) );
  MUX2_X1 U664 ( .A(n57), .B(n56), .S(n242), .Z(n58) );
  MUX2_X1 U665 ( .A(n58), .B(n55), .S(n241), .Z(n59) );
  MUX2_X1 U666 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U667 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U668 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n249), .Z(n61) );
  MUX2_X1 U669 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n246), .Z(n62) );
  MUX2_X1 U670 ( .A(n62), .B(n61), .S(n243), .Z(n63) );
  MUX2_X1 U671 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n248), .Z(n64) );
  MUX2_X1 U672 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n245), .Z(n65) );
  MUX2_X1 U673 ( .A(n65), .B(n64), .S(n243), .Z(n66) );
  MUX2_X1 U674 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U675 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n249), .Z(n68) );
  MUX2_X1 U676 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n248), .Z(n69) );
  MUX2_X1 U677 ( .A(n69), .B(n68), .S(n243), .Z(n70) );
  MUX2_X1 U678 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n249), .Z(n71) );
  MUX2_X1 U679 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n246), .Z(n72) );
  MUX2_X1 U680 ( .A(n72), .B(n71), .S(n243), .Z(n73) );
  MUX2_X1 U681 ( .A(n73), .B(n70), .S(n241), .Z(n74) );
  MUX2_X1 U682 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U683 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n245), .Z(n76) );
  MUX2_X1 U684 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n246), .Z(n77) );
  MUX2_X1 U685 ( .A(n77), .B(n76), .S(n243), .Z(n78) );
  MUX2_X1 U686 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n245), .Z(n79) );
  MUX2_X1 U687 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n249), .Z(n80) );
  MUX2_X1 U688 ( .A(n80), .B(n79), .S(n243), .Z(n81) );
  MUX2_X1 U689 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U690 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n250), .Z(n83) );
  MUX2_X1 U691 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n250), .Z(n84) );
  MUX2_X1 U692 ( .A(n84), .B(n83), .S(n243), .Z(n85) );
  MUX2_X1 U693 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n250), .Z(n86) );
  MUX2_X1 U694 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n248), .Z(n87) );
  MUX2_X1 U695 ( .A(n87), .B(n86), .S(n243), .Z(n88) );
  MUX2_X1 U696 ( .A(n88), .B(n85), .S(n241), .Z(n89) );
  MUX2_X1 U697 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U698 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U699 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n250), .Z(n91) );
  MUX2_X1 U700 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n250), .Z(n92) );
  MUX2_X1 U701 ( .A(n92), .B(n91), .S(n243), .Z(n93) );
  MUX2_X1 U702 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n250), .Z(n94) );
  MUX2_X1 U703 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n250), .Z(n95) );
  MUX2_X1 U704 ( .A(n95), .B(n94), .S(n243), .Z(n96) );
  MUX2_X1 U705 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U706 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n250), .Z(n98) );
  MUX2_X1 U707 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n250), .Z(n99) );
  MUX2_X1 U708 ( .A(n99), .B(n98), .S(n243), .Z(n100) );
  MUX2_X1 U709 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n250), .Z(n101) );
  MUX2_X1 U710 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n250), .Z(n102) );
  MUX2_X1 U711 ( .A(n102), .B(n101), .S(n243), .Z(n103) );
  MUX2_X1 U712 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U713 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U714 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n247), .Z(n106) );
  MUX2_X1 U715 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n247), .Z(n107) );
  MUX2_X1 U716 ( .A(n107), .B(n106), .S(n244), .Z(n108) );
  MUX2_X1 U717 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n247), .Z(n109) );
  MUX2_X1 U718 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n247), .Z(n110) );
  MUX2_X1 U719 ( .A(n110), .B(n109), .S(n244), .Z(n111) );
  MUX2_X1 U720 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U721 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n247), .Z(n113) );
  MUX2_X1 U722 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n247), .Z(n114) );
  MUX2_X1 U723 ( .A(n114), .B(n113), .S(n244), .Z(n115) );
  MUX2_X1 U724 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n247), .Z(n116) );
  MUX2_X1 U725 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n247), .Z(n117) );
  MUX2_X1 U726 ( .A(n117), .B(n116), .S(n244), .Z(n118) );
  MUX2_X1 U727 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U728 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U729 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U730 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n247), .Z(n121) );
  MUX2_X1 U731 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n247), .Z(n122) );
  MUX2_X1 U732 ( .A(n122), .B(n121), .S(n244), .Z(n123) );
  MUX2_X1 U733 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n247), .Z(n124) );
  MUX2_X1 U734 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n247), .Z(n125) );
  MUX2_X1 U735 ( .A(n125), .B(n124), .S(n244), .Z(n126) );
  MUX2_X1 U736 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U737 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n248), .Z(n128) );
  MUX2_X1 U738 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n248), .Z(n129) );
  MUX2_X1 U739 ( .A(n129), .B(n128), .S(n244), .Z(n130) );
  MUX2_X1 U740 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n248), .Z(n131) );
  MUX2_X1 U741 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n248), .Z(n132) );
  MUX2_X1 U742 ( .A(n132), .B(n131), .S(n244), .Z(n133) );
  MUX2_X1 U743 ( .A(n133), .B(n130), .S(n241), .Z(n134) );
  MUX2_X1 U744 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U745 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n248), .Z(n136) );
  MUX2_X1 U746 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n248), .Z(n137) );
  MUX2_X1 U747 ( .A(n137), .B(n136), .S(n244), .Z(n138) );
  MUX2_X1 U748 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n248), .Z(n139) );
  MUX2_X1 U749 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n248), .Z(n140) );
  MUX2_X1 U750 ( .A(n140), .B(n139), .S(n244), .Z(n141) );
  MUX2_X1 U751 ( .A(n141), .B(n138), .S(n241), .Z(n142) );
  MUX2_X1 U752 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n248), .Z(n143) );
  MUX2_X1 U753 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n248), .Z(n144) );
  MUX2_X1 U754 ( .A(n144), .B(n143), .S(n244), .Z(n145) );
  MUX2_X1 U755 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n248), .Z(n146) );
  MUX2_X1 U756 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n248), .Z(n147) );
  MUX2_X1 U757 ( .A(n147), .B(n146), .S(n244), .Z(n148) );
  MUX2_X1 U758 ( .A(n148), .B(n145), .S(n241), .Z(n149) );
  MUX2_X1 U759 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U760 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U761 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n249), .Z(n151) );
  MUX2_X1 U762 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n249), .Z(n152) );
  MUX2_X1 U763 ( .A(n152), .B(n151), .S(N11), .Z(n153) );
  MUX2_X1 U764 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n249), .Z(n154) );
  MUX2_X1 U765 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n249), .Z(n155) );
  MUX2_X1 U766 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U767 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U768 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n249), .Z(n158) );
  MUX2_X1 U769 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n249), .Z(n159) );
  MUX2_X1 U770 ( .A(n159), .B(n158), .S(N11), .Z(n160) );
  MUX2_X1 U771 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n249), .Z(n161) );
  MUX2_X1 U772 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n249), .Z(n162) );
  MUX2_X1 U773 ( .A(n162), .B(n161), .S(n244), .Z(n163) );
  MUX2_X1 U774 ( .A(n163), .B(n160), .S(N12), .Z(n164) );
  MUX2_X1 U775 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U776 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n249), .Z(n166) );
  MUX2_X1 U777 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n249), .Z(n167) );
  MUX2_X1 U778 ( .A(n167), .B(n166), .S(N11), .Z(n168) );
  MUX2_X1 U779 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n249), .Z(n169) );
  MUX2_X1 U780 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n249), .Z(n170) );
  MUX2_X1 U781 ( .A(n170), .B(n169), .S(n243), .Z(n171) );
  MUX2_X1 U782 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U783 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n247), .Z(n173) );
  MUX2_X1 U784 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n250), .Z(n174) );
  MUX2_X1 U785 ( .A(n174), .B(n173), .S(n242), .Z(n175) );
  MUX2_X1 U786 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(N10), .Z(n176) );
  MUX2_X1 U787 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n250), .Z(n177) );
  MUX2_X1 U788 ( .A(n177), .B(n176), .S(n243), .Z(n178) );
  MUX2_X1 U789 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U790 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U791 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U792 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n249), .Z(n181) );
  MUX2_X1 U793 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n250), .Z(n182) );
  MUX2_X1 U794 ( .A(n182), .B(n181), .S(N11), .Z(n183) );
  MUX2_X1 U795 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n248), .Z(n184) );
  MUX2_X1 U796 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(N10), .Z(n185) );
  MUX2_X1 U797 ( .A(n185), .B(n184), .S(N11), .Z(n186) );
  MUX2_X1 U798 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U799 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n245), .Z(n188) );
  MUX2_X1 U800 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(N10), .Z(n189) );
  MUX2_X1 U801 ( .A(n189), .B(n188), .S(N11), .Z(n190) );
  MUX2_X1 U802 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n248), .Z(n191) );
  MUX2_X1 U803 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n250), .Z(n192) );
  MUX2_X1 U804 ( .A(n192), .B(n191), .S(n242), .Z(n193) );
  MUX2_X1 U805 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U806 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U807 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n246), .Z(n196) );
  MUX2_X1 U808 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n250), .Z(n197) );
  MUX2_X1 U809 ( .A(n197), .B(n196), .S(N11), .Z(n198) );
  MUX2_X1 U810 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n250), .Z(n199) );
  MUX2_X1 U811 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(N10), .Z(n200) );
  MUX2_X1 U812 ( .A(n200), .B(n199), .S(n242), .Z(n201) );
  MUX2_X1 U813 ( .A(n201), .B(n198), .S(N12), .Z(n202) );
  MUX2_X1 U814 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n250), .Z(n203) );
  MUX2_X1 U815 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(N10), .Z(n204) );
  MUX2_X1 U816 ( .A(n204), .B(n203), .S(n243), .Z(n205) );
  MUX2_X1 U817 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(N10), .Z(n206) );
  MUX2_X1 U818 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(N10), .Z(n207) );
  MUX2_X1 U819 ( .A(n207), .B(n206), .S(N11), .Z(n208) );
  MUX2_X1 U820 ( .A(n208), .B(n205), .S(N12), .Z(n209) );
  MUX2_X1 U821 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U822 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U823 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n246), .Z(n211) );
  MUX2_X1 U824 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n245), .Z(n212) );
  MUX2_X1 U825 ( .A(n212), .B(n211), .S(n243), .Z(n213) );
  MUX2_X1 U826 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n246), .Z(n214) );
  MUX2_X1 U827 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(N10), .Z(n215) );
  MUX2_X1 U828 ( .A(n215), .B(n214), .S(n244), .Z(n216) );
  MUX2_X1 U829 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U830 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n247), .Z(n218) );
  MUX2_X1 U831 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n250), .Z(n219) );
  MUX2_X1 U832 ( .A(n219), .B(n218), .S(n244), .Z(n220) );
  MUX2_X1 U833 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n247), .Z(n221) );
  MUX2_X1 U834 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(N10), .Z(n222) );
  MUX2_X1 U835 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U836 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U837 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U838 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n247), .Z(n226) );
  MUX2_X1 U839 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n250), .Z(n227) );
  MUX2_X1 U840 ( .A(n227), .B(n226), .S(n243), .Z(n228) );
  MUX2_X1 U841 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n247), .Z(n229) );
  MUX2_X1 U842 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(N10), .Z(n230) );
  MUX2_X1 U843 ( .A(n230), .B(n229), .S(N11), .Z(n231) );
  MUX2_X1 U844 ( .A(n231), .B(n228), .S(N12), .Z(n232) );
  MUX2_X1 U845 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(N10), .Z(n233) );
  MUX2_X1 U846 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(N10), .Z(n234) );
  MUX2_X1 U847 ( .A(n234), .B(n233), .S(n244), .Z(n235) );
  MUX2_X1 U848 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(N10), .Z(n236) );
  MUX2_X1 U849 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(N10), .Z(n237) );
  MUX2_X1 U850 ( .A(n237), .B(n236), .S(N11), .Z(n238) );
  MUX2_X1 U851 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U852 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U853 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
endmodule


module memory_WIDTH8_SIZE32_LOGSIZE5_1 ( clk, data_in, data_out, addr, wr_en
 );
  input [7:0] data_in;
  output [7:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][7] , \mem[31][6] , \mem[31][5] ,
         \mem[31][4] , \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] ,
         \mem[30][7] , \mem[30][6] , \mem[30][5] , \mem[30][4] , \mem[30][3] ,
         \mem[30][2] , \mem[30][1] , \mem[30][0] , \mem[29][7] , \mem[29][6] ,
         \mem[29][5] , \mem[29][4] , \mem[29][3] , \mem[29][2] , \mem[29][1] ,
         \mem[29][0] , \mem[28][7] , \mem[28][6] , \mem[28][5] , \mem[28][4] ,
         \mem[28][3] , \mem[28][2] , \mem[28][1] , \mem[28][0] , \mem[27][7] ,
         \mem[27][6] , \mem[27][5] , \mem[27][4] , \mem[27][3] , \mem[27][2] ,
         \mem[27][1] , \mem[27][0] , \mem[26][7] , \mem[26][6] , \mem[26][5] ,
         \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] , \mem[26][0] ,
         \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] , \mem[25][3] ,
         \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][7] ,
         \mem[22][6] , \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] ,
         \mem[22][1] , \mem[22][0] , \mem[21][7] , \mem[21][6] , \mem[21][5] ,
         \mem[21][4] , \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] ,
         \mem[20][7] , \mem[20][6] , \mem[20][5] , \mem[20][4] , \mem[20][3] ,
         \mem[20][2] , \mem[20][1] , \mem[20][0] , \mem[19][7] , \mem[19][6] ,
         \mem[19][5] , \mem[19][4] , \mem[19][3] , \mem[19][2] , \mem[19][1] ,
         \mem[19][0] , \mem[18][7] , \mem[18][6] , \mem[18][5] , \mem[18][4] ,
         \mem[18][3] , \mem[18][2] , \mem[18][1] , \mem[18][0] , \mem[17][7] ,
         \mem[17][6] , \mem[17][5] , \mem[17][4] , \mem[17][3] , \mem[17][2] ,
         \mem[17][1] , \mem[17][0] , \mem[16][7] , \mem[16][6] , \mem[16][5] ,
         \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] , \mem[16][0] ,
         \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] , \mem[15][3] ,
         \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][7] ,
         \mem[12][6] , \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] ,
         \mem[12][1] , \mem[12][0] , \mem[11][7] , \mem[11][6] , \mem[11][5] ,
         \mem[11][4] , \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] ,
         \mem[10][7] , \mem[10][6] , \mem[10][5] , \mem[10][4] , \mem[10][3] ,
         \mem[10][2] , \mem[10][1] , \mem[10][0] , \mem[9][7] , \mem[9][6] ,
         \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] , \mem[9][1] ,
         \mem[9][0] , \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] ,
         \mem[8][3] , \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][7] ,
         \mem[7][6] , \mem[7][5] , \mem[7][4] , \mem[7][3] , \mem[7][2] ,
         \mem[7][1] , \mem[7][0] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][7] , \mem[5][6] , \mem[5][5] , \mem[5][4] , \mem[5][3] ,
         \mem[5][2] , \mem[5][1] , \mem[5][0] , \mem[4][7] , \mem[4][6] ,
         \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] , \mem[4][1] ,
         \mem[4][0] , \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] ,
         \mem[3][3] , \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][7] ,
         \mem[2][6] , \mem[2][5] , \mem[2][4] , \mem[2][3] , \mem[2][2] ,
         \mem[2][1] , \mem[2][0] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][7] , \mem[0][6] , \mem[0][5] , \mem[0][4] , \mem[0][3] ,
         \mem[0][2] , \mem[0][1] , \mem[0][0] , N15, N16, N17, N18, N19, N20,
         N21, N22, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[7]  ( .D(N15), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N16), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N17), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N18), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[2]  ( .D(N20), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[0]  ( .D(N22), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][7]  ( .D(n254), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n255), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n256), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n257), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n258), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n259), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n260), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n261), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n262), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n263), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n264), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n265), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n266), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n267), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n268), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n269), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n270), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n271), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n272), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n273), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n274), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n275), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n276), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n277), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n278), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n279), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n280), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n281), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n282), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n283), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n284), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n285), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n286), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n287), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n288), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n289), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n290), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n291), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n292), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n293), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n594), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n595), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n596), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n597), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n598), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n599), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n600), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n601), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n602), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n603), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n604), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n605), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n606), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n607), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n608), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n609), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n610), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n611), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n612), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n613), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n614), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n615), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n616), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n617), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n618), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n619), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n620), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n621), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n622), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n623), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n624), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n625), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n626), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n627), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n628), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n629), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n630), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n631), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n632), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n633), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n634), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n635), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n636), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n637), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n638), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n639), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n640), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n641), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n642), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n643), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n644), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n645), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n646), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n647), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n648), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n649), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n650), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n651), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n652), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n653), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n654), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n655), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n656), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n657), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n658), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n659), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n660), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n661), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n662), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n663), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n664), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n665), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n666), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n667), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n668), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n669), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n670), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n671), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n672), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n673), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n674), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n675), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n676), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n677), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n678), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n679), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n680), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n681), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n682), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n683), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n684), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n685), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n686), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n687), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n688), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n689), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n690), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n691), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n692), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n693), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n694), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n695), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n696), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n697), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n698), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n699), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n700), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n701), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n702), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n703), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n704), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n705), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n706), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n707), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n708), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n709), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n710), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n711), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n712), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n713), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n714), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n715), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n716), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n717), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n718), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n719), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n720), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n721), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n722), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n723), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n724), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n725), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n726), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n727), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n728), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n729), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n730), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n731), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n732), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n733), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n734), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n735), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n736), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n737), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n738), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n739), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n740), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n741), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n742), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n743), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n744), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n745), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n746), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n747), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n748), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n749), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n750), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n751), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n752), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n753), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n754), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n755), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n756), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n757), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n758), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n759), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n760), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n761), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n762), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n763), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n764), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n765), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n766), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n767), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n768), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n769), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n770), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n771), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n772), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n773), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n774), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n775), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n776), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n777), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n778), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n779), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n780), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n781), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n782), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n783), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n784), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n785), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n786), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n787), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n788), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n789), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n790), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n791), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n792), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n793), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n794), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n795), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n796), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n797), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n798), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n799), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n800), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n801), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n802), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n803), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n804), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n805), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n806), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n807), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n808), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n809), .CK(clk), .Q(\mem[0][0] ) );
  DFF_X1 \data_out_reg[1]  ( .D(N21), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[3]  ( .D(N19), .CK(clk), .Q(data_out[3]) );
  BUF_X1 U3 ( .A(n250), .Z(n247) );
  BUF_X1 U4 ( .A(n250), .Z(n246) );
  BUF_X1 U5 ( .A(n250), .Z(n248) );
  BUF_X1 U6 ( .A(n250), .Z(n249) );
  BUF_X1 U7 ( .A(N10), .Z(n250) );
  INV_X1 U8 ( .A(n1111), .ZN(n841) );
  INV_X1 U9 ( .A(n1100), .ZN(n840) );
  INV_X1 U10 ( .A(n1090), .ZN(n839) );
  INV_X1 U11 ( .A(n1080), .ZN(n838) );
  INV_X1 U12 ( .A(n1070), .ZN(n837) );
  INV_X1 U13 ( .A(n1060), .ZN(n836) );
  INV_X1 U14 ( .A(n1051), .ZN(n835) );
  INV_X1 U15 ( .A(n1042), .ZN(n834) );
  NOR3_X1 U16 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n1103) );
  NOR3_X1 U17 ( .A1(N11), .A2(N12), .A3(n251), .ZN(n1092) );
  NAND2_X1 U18 ( .A1(n1102), .A2(n1134), .ZN(n1060) );
  NAND2_X1 U19 ( .A1(n1103), .A2(n1102), .ZN(n1111) );
  NAND2_X1 U20 ( .A1(n1092), .A2(n1102), .ZN(n1100) );
  NAND2_X1 U21 ( .A1(n1082), .A2(n1102), .ZN(n1090) );
  NAND2_X1 U22 ( .A1(n1072), .A2(n1102), .ZN(n1080) );
  NAND2_X1 U23 ( .A1(n1062), .A2(n1102), .ZN(n1070) );
  NAND2_X1 U24 ( .A1(n1102), .A2(n1123), .ZN(n1051) );
  NAND2_X1 U25 ( .A1(n1102), .A2(n1113), .ZN(n1042) );
  INV_X1 U26 ( .A(n1131), .ZN(n816) );
  INV_X1 U27 ( .A(n1121), .ZN(n815) );
  INV_X1 U28 ( .A(n887), .ZN(n814) );
  INV_X1 U29 ( .A(n878), .ZN(n813) );
  INV_X1 U30 ( .A(n869), .ZN(n812) );
  INV_X1 U31 ( .A(n860), .ZN(n811) );
  INV_X1 U32 ( .A(n851), .ZN(n810) );
  INV_X1 U33 ( .A(n987), .ZN(n828) );
  INV_X1 U34 ( .A(n978), .ZN(n827) );
  INV_X1 U35 ( .A(n969), .ZN(n826) );
  INV_X1 U36 ( .A(n914), .ZN(n820) );
  INV_X1 U37 ( .A(n905), .ZN(n819) );
  INV_X1 U38 ( .A(n896), .ZN(n818) );
  INV_X1 U39 ( .A(n1033), .ZN(n833) );
  INV_X1 U40 ( .A(n1023), .ZN(n832) );
  INV_X1 U41 ( .A(n1014), .ZN(n831) );
  INV_X1 U42 ( .A(n1005), .ZN(n830) );
  INV_X1 U43 ( .A(n996), .ZN(n829) );
  INV_X1 U44 ( .A(n960), .ZN(n825) );
  INV_X1 U45 ( .A(n950), .ZN(n824) );
  INV_X1 U46 ( .A(n941), .ZN(n823) );
  INV_X1 U47 ( .A(n932), .ZN(n822) );
  INV_X1 U48 ( .A(n923), .ZN(n821) );
  INV_X1 U49 ( .A(n1142), .ZN(n817) );
  BUF_X1 U50 ( .A(N11), .Z(n242) );
  BUF_X1 U51 ( .A(N11), .Z(n243) );
  BUF_X1 U52 ( .A(N11), .Z(n244) );
  INV_X1 U53 ( .A(N10), .ZN(n251) );
  BUF_X1 U54 ( .A(N12), .Z(n241) );
  NOR3_X1 U55 ( .A1(n253), .A2(N10), .A3(n252), .ZN(n1123) );
  NOR3_X1 U56 ( .A1(n253), .A2(n251), .A3(n252), .ZN(n1113) );
  NOR3_X1 U57 ( .A1(n251), .A2(N11), .A3(n253), .ZN(n1134) );
  NOR3_X1 U58 ( .A1(N10), .A2(N12), .A3(n252), .ZN(n1082) );
  NOR3_X1 U59 ( .A1(n251), .A2(N12), .A3(n252), .ZN(n1072) );
  NOR3_X1 U60 ( .A1(N10), .A2(N11), .A3(n253), .ZN(n1062) );
  NAND2_X1 U61 ( .A1(n1025), .A2(n1134), .ZN(n987) );
  NAND2_X1 U62 ( .A1(n952), .A2(n1134), .ZN(n914) );
  NAND2_X1 U63 ( .A1(n1025), .A2(n1062), .ZN(n996) );
  NAND2_X1 U64 ( .A1(n952), .A2(n1062), .ZN(n923) );
  NAND2_X1 U65 ( .A1(n1025), .A2(n1103), .ZN(n1033) );
  NAND2_X1 U66 ( .A1(n1025), .A2(n1092), .ZN(n1023) );
  NAND2_X1 U67 ( .A1(n952), .A2(n1103), .ZN(n960) );
  NAND2_X1 U68 ( .A1(n952), .A2(n1092), .ZN(n950) );
  NAND2_X1 U69 ( .A1(n1103), .A2(n1133), .ZN(n887) );
  NAND2_X1 U70 ( .A1(n1092), .A2(n1133), .ZN(n878) );
  NAND2_X1 U71 ( .A1(n1082), .A2(n1133), .ZN(n869) );
  NAND2_X1 U72 ( .A1(n1072), .A2(n1133), .ZN(n860) );
  NAND2_X1 U73 ( .A1(n1062), .A2(n1133), .ZN(n851) );
  NAND2_X1 U74 ( .A1(n1134), .A2(n1133), .ZN(n1142) );
  NAND2_X1 U75 ( .A1(n1123), .A2(n1133), .ZN(n1131) );
  NAND2_X1 U76 ( .A1(n1113), .A2(n1133), .ZN(n1121) );
  NAND2_X1 U77 ( .A1(n1025), .A2(n1082), .ZN(n1014) );
  NAND2_X1 U78 ( .A1(n1025), .A2(n1072), .ZN(n1005) );
  NAND2_X1 U79 ( .A1(n952), .A2(n1082), .ZN(n941) );
  NAND2_X1 U80 ( .A1(n952), .A2(n1072), .ZN(n932) );
  NAND2_X1 U81 ( .A1(n1025), .A2(n1123), .ZN(n978) );
  NAND2_X1 U82 ( .A1(n952), .A2(n1123), .ZN(n905) );
  NAND2_X1 U83 ( .A1(n1025), .A2(n1113), .ZN(n969) );
  NAND2_X1 U84 ( .A1(n952), .A2(n1113), .ZN(n896) );
  AND3_X1 U85 ( .A1(n842), .A2(n843), .A3(wr_en), .ZN(n1102) );
  AND3_X1 U86 ( .A1(N14), .A2(N13), .A3(wr_en), .ZN(n1133) );
  AND3_X1 U87 ( .A1(N13), .A2(n843), .A3(wr_en), .ZN(n1025) );
  AND3_X1 U88 ( .A1(N14), .A2(n842), .A3(wr_en), .ZN(n952) );
  INV_X1 U89 ( .A(n1059), .ZN(n768) );
  AOI22_X1 U90 ( .A1(data_in[1]), .A2(n836), .B1(n1060), .B2(\mem[5][1] ), 
        .ZN(n1059) );
  INV_X1 U91 ( .A(n1058), .ZN(n767) );
  AOI22_X1 U92 ( .A1(data_in[2]), .A2(n836), .B1(n1060), .B2(\mem[5][2] ), 
        .ZN(n1058) );
  INV_X1 U93 ( .A(n1057), .ZN(n766) );
  AOI22_X1 U94 ( .A1(data_in[3]), .A2(n836), .B1(n1060), .B2(\mem[5][3] ), 
        .ZN(n1057) );
  INV_X1 U95 ( .A(n1056), .ZN(n765) );
  AOI22_X1 U96 ( .A1(data_in[4]), .A2(n836), .B1(n1060), .B2(\mem[5][4] ), 
        .ZN(n1056) );
  INV_X1 U97 ( .A(n1055), .ZN(n764) );
  AOI22_X1 U98 ( .A1(data_in[5]), .A2(n836), .B1(n1060), .B2(\mem[5][5] ), 
        .ZN(n1055) );
  INV_X1 U99 ( .A(n1054), .ZN(n763) );
  AOI22_X1 U100 ( .A1(data_in[6]), .A2(n836), .B1(n1060), .B2(\mem[5][6] ), 
        .ZN(n1054) );
  INV_X1 U101 ( .A(n1053), .ZN(n762) );
  AOI22_X1 U102 ( .A1(data_in[7]), .A2(n836), .B1(n1060), .B2(\mem[5][7] ), 
        .ZN(n1053) );
  INV_X1 U103 ( .A(n985), .ZN(n703) );
  AOI22_X1 U104 ( .A1(data_in[2]), .A2(n828), .B1(n987), .B2(\mem[13][2] ), 
        .ZN(n985) );
  INV_X1 U105 ( .A(n984), .ZN(n702) );
  AOI22_X1 U106 ( .A1(data_in[3]), .A2(n828), .B1(n987), .B2(\mem[13][3] ), 
        .ZN(n984) );
  INV_X1 U107 ( .A(n983), .ZN(n701) );
  AOI22_X1 U108 ( .A1(data_in[4]), .A2(n828), .B1(n987), .B2(\mem[13][4] ), 
        .ZN(n983) );
  INV_X1 U109 ( .A(n982), .ZN(n700) );
  AOI22_X1 U110 ( .A1(data_in[5]), .A2(n828), .B1(n987), .B2(\mem[13][5] ), 
        .ZN(n982) );
  INV_X1 U111 ( .A(n981), .ZN(n699) );
  AOI22_X1 U112 ( .A1(data_in[6]), .A2(n828), .B1(n987), .B2(\mem[13][6] ), 
        .ZN(n981) );
  INV_X1 U113 ( .A(n980), .ZN(n698) );
  AOI22_X1 U114 ( .A1(data_in[7]), .A2(n828), .B1(n987), .B2(\mem[13][7] ), 
        .ZN(n980) );
  INV_X1 U115 ( .A(n1061), .ZN(n769) );
  AOI22_X1 U116 ( .A1(data_in[0]), .A2(n836), .B1(n1060), .B2(\mem[5][0] ), 
        .ZN(n1061) );
  INV_X1 U117 ( .A(n945), .ZN(n668) );
  AOI22_X1 U118 ( .A1(data_in[5]), .A2(n824), .B1(n950), .B2(\mem[17][5] ), 
        .ZN(n945) );
  INV_X1 U119 ( .A(n915), .ZN(n641) );
  AOI22_X1 U120 ( .A1(data_in[0]), .A2(n820), .B1(n914), .B2(\mem[21][0] ), 
        .ZN(n915) );
  INV_X1 U121 ( .A(n913), .ZN(n640) );
  AOI22_X1 U122 ( .A1(data_in[1]), .A2(n820), .B1(n914), .B2(\mem[21][1] ), 
        .ZN(n913) );
  INV_X1 U123 ( .A(n912), .ZN(n639) );
  AOI22_X1 U124 ( .A1(data_in[2]), .A2(n820), .B1(n914), .B2(\mem[21][2] ), 
        .ZN(n912) );
  INV_X1 U125 ( .A(n911), .ZN(n638) );
  AOI22_X1 U126 ( .A1(data_in[3]), .A2(n820), .B1(n914), .B2(\mem[21][3] ), 
        .ZN(n911) );
  INV_X1 U127 ( .A(n910), .ZN(n637) );
  AOI22_X1 U128 ( .A1(data_in[4]), .A2(n820), .B1(n914), .B2(\mem[21][4] ), 
        .ZN(n910) );
  INV_X1 U129 ( .A(n909), .ZN(n636) );
  AOI22_X1 U130 ( .A1(data_in[5]), .A2(n820), .B1(n914), .B2(\mem[21][5] ), 
        .ZN(n909) );
  INV_X1 U131 ( .A(n908), .ZN(n635) );
  AOI22_X1 U132 ( .A1(data_in[6]), .A2(n820), .B1(n914), .B2(\mem[21][6] ), 
        .ZN(n908) );
  INV_X1 U133 ( .A(n907), .ZN(n634) );
  AOI22_X1 U134 ( .A1(data_in[7]), .A2(n820), .B1(n914), .B2(\mem[21][7] ), 
        .ZN(n907) );
  INV_X1 U135 ( .A(n951), .ZN(n673) );
  AOI22_X1 U136 ( .A1(data_in[0]), .A2(n824), .B1(n950), .B2(\mem[17][0] ), 
        .ZN(n951) );
  INV_X1 U137 ( .A(n949), .ZN(n672) );
  AOI22_X1 U138 ( .A1(data_in[1]), .A2(n824), .B1(n950), .B2(\mem[17][1] ), 
        .ZN(n949) );
  INV_X1 U139 ( .A(n948), .ZN(n671) );
  AOI22_X1 U140 ( .A1(data_in[2]), .A2(n824), .B1(n950), .B2(\mem[17][2] ), 
        .ZN(n948) );
  INV_X1 U141 ( .A(n947), .ZN(n670) );
  AOI22_X1 U142 ( .A1(data_in[3]), .A2(n824), .B1(n950), .B2(\mem[17][3] ), 
        .ZN(n947) );
  INV_X1 U143 ( .A(n1024), .ZN(n737) );
  AOI22_X1 U144 ( .A1(data_in[0]), .A2(n832), .B1(n1023), .B2(\mem[9][0] ), 
        .ZN(n1024) );
  INV_X1 U145 ( .A(n1022), .ZN(n736) );
  AOI22_X1 U146 ( .A1(data_in[1]), .A2(n832), .B1(n1023), .B2(\mem[9][1] ), 
        .ZN(n1022) );
  INV_X1 U147 ( .A(n1021), .ZN(n735) );
  AOI22_X1 U148 ( .A1(data_in[2]), .A2(n832), .B1(n1023), .B2(\mem[9][2] ), 
        .ZN(n1021) );
  INV_X1 U149 ( .A(n1020), .ZN(n734) );
  AOI22_X1 U150 ( .A1(data_in[3]), .A2(n832), .B1(n1023), .B2(\mem[9][3] ), 
        .ZN(n1020) );
  INV_X1 U151 ( .A(n1018), .ZN(n732) );
  AOI22_X1 U152 ( .A1(data_in[5]), .A2(n832), .B1(n1023), .B2(\mem[9][5] ), 
        .ZN(n1018) );
  INV_X1 U153 ( .A(n1017), .ZN(n731) );
  AOI22_X1 U154 ( .A1(data_in[6]), .A2(n832), .B1(n1023), .B2(\mem[9][6] ), 
        .ZN(n1017) );
  INV_X1 U155 ( .A(n1016), .ZN(n730) );
  AOI22_X1 U156 ( .A1(data_in[7]), .A2(n832), .B1(n1023), .B2(\mem[9][7] ), 
        .ZN(n1016) );
  INV_X1 U157 ( .A(n988), .ZN(n705) );
  AOI22_X1 U158 ( .A1(data_in[0]), .A2(n828), .B1(n987), .B2(\mem[13][0] ), 
        .ZN(n988) );
  INV_X1 U159 ( .A(n986), .ZN(n704) );
  AOI22_X1 U160 ( .A1(data_in[1]), .A2(n828), .B1(n987), .B2(\mem[13][1] ), 
        .ZN(n986) );
  INV_X1 U161 ( .A(n946), .ZN(n669) );
  AOI22_X1 U162 ( .A1(data_in[4]), .A2(n824), .B1(n950), .B2(\mem[17][4] ), 
        .ZN(n946) );
  INV_X1 U163 ( .A(n944), .ZN(n667) );
  AOI22_X1 U164 ( .A1(data_in[6]), .A2(n824), .B1(n950), .B2(\mem[17][6] ), 
        .ZN(n944) );
  INV_X1 U165 ( .A(n943), .ZN(n666) );
  AOI22_X1 U166 ( .A1(data_in[7]), .A2(n824), .B1(n950), .B2(\mem[17][7] ), 
        .ZN(n943) );
  INV_X1 U167 ( .A(n979), .ZN(n697) );
  AOI22_X1 U168 ( .A1(data_in[0]), .A2(n827), .B1(n978), .B2(\mem[14][0] ), 
        .ZN(n979) );
  INV_X1 U169 ( .A(n977), .ZN(n696) );
  AOI22_X1 U170 ( .A1(data_in[1]), .A2(n827), .B1(n978), .B2(\mem[14][1] ), 
        .ZN(n977) );
  INV_X1 U171 ( .A(n976), .ZN(n695) );
  AOI22_X1 U172 ( .A1(data_in[2]), .A2(n827), .B1(n978), .B2(\mem[14][2] ), 
        .ZN(n976) );
  INV_X1 U173 ( .A(n975), .ZN(n694) );
  AOI22_X1 U174 ( .A1(data_in[3]), .A2(n827), .B1(n978), .B2(\mem[14][3] ), 
        .ZN(n975) );
  INV_X1 U175 ( .A(n974), .ZN(n693) );
  AOI22_X1 U176 ( .A1(data_in[4]), .A2(n827), .B1(n978), .B2(\mem[14][4] ), 
        .ZN(n974) );
  INV_X1 U177 ( .A(n973), .ZN(n692) );
  AOI22_X1 U178 ( .A1(data_in[5]), .A2(n827), .B1(n978), .B2(\mem[14][5] ), 
        .ZN(n973) );
  INV_X1 U179 ( .A(n972), .ZN(n691) );
  AOI22_X1 U180 ( .A1(data_in[6]), .A2(n827), .B1(n978), .B2(\mem[14][6] ), 
        .ZN(n972) );
  INV_X1 U181 ( .A(n971), .ZN(n690) );
  AOI22_X1 U182 ( .A1(data_in[7]), .A2(n827), .B1(n978), .B2(\mem[14][7] ), 
        .ZN(n971) );
  INV_X1 U183 ( .A(n970), .ZN(n689) );
  AOI22_X1 U184 ( .A1(data_in[0]), .A2(n826), .B1(n969), .B2(\mem[15][0] ), 
        .ZN(n970) );
  INV_X1 U185 ( .A(n968), .ZN(n688) );
  AOI22_X1 U186 ( .A1(data_in[1]), .A2(n826), .B1(n969), .B2(\mem[15][1] ), 
        .ZN(n968) );
  INV_X1 U187 ( .A(n967), .ZN(n687) );
  AOI22_X1 U188 ( .A1(data_in[2]), .A2(n826), .B1(n969), .B2(\mem[15][2] ), 
        .ZN(n967) );
  INV_X1 U189 ( .A(n966), .ZN(n686) );
  AOI22_X1 U190 ( .A1(data_in[3]), .A2(n826), .B1(n969), .B2(\mem[15][3] ), 
        .ZN(n966) );
  INV_X1 U191 ( .A(n965), .ZN(n685) );
  AOI22_X1 U192 ( .A1(data_in[4]), .A2(n826), .B1(n969), .B2(\mem[15][4] ), 
        .ZN(n965) );
  INV_X1 U193 ( .A(n964), .ZN(n684) );
  AOI22_X1 U194 ( .A1(data_in[5]), .A2(n826), .B1(n969), .B2(\mem[15][5] ), 
        .ZN(n964) );
  INV_X1 U195 ( .A(n963), .ZN(n683) );
  AOI22_X1 U196 ( .A1(data_in[6]), .A2(n826), .B1(n969), .B2(\mem[15][6] ), 
        .ZN(n963) );
  INV_X1 U197 ( .A(n962), .ZN(n682) );
  AOI22_X1 U198 ( .A1(data_in[7]), .A2(n826), .B1(n969), .B2(\mem[15][7] ), 
        .ZN(n962) );
  INV_X1 U199 ( .A(n942), .ZN(n665) );
  AOI22_X1 U200 ( .A1(data_in[0]), .A2(n823), .B1(n941), .B2(\mem[18][0] ), 
        .ZN(n942) );
  INV_X1 U201 ( .A(n940), .ZN(n664) );
  AOI22_X1 U202 ( .A1(data_in[1]), .A2(n823), .B1(n941), .B2(\mem[18][1] ), 
        .ZN(n940) );
  INV_X1 U203 ( .A(n939), .ZN(n663) );
  AOI22_X1 U204 ( .A1(data_in[2]), .A2(n823), .B1(n941), .B2(\mem[18][2] ), 
        .ZN(n939) );
  INV_X1 U205 ( .A(n938), .ZN(n662) );
  AOI22_X1 U206 ( .A1(data_in[3]), .A2(n823), .B1(n941), .B2(\mem[18][3] ), 
        .ZN(n938) );
  INV_X1 U207 ( .A(n937), .ZN(n661) );
  AOI22_X1 U208 ( .A1(data_in[4]), .A2(n823), .B1(n941), .B2(\mem[18][4] ), 
        .ZN(n937) );
  INV_X1 U209 ( .A(n936), .ZN(n660) );
  AOI22_X1 U210 ( .A1(data_in[5]), .A2(n823), .B1(n941), .B2(\mem[18][5] ), 
        .ZN(n936) );
  INV_X1 U211 ( .A(n935), .ZN(n659) );
  AOI22_X1 U212 ( .A1(data_in[6]), .A2(n823), .B1(n941), .B2(\mem[18][6] ), 
        .ZN(n935) );
  INV_X1 U213 ( .A(n934), .ZN(n658) );
  AOI22_X1 U214 ( .A1(data_in[7]), .A2(n823), .B1(n941), .B2(\mem[18][7] ), 
        .ZN(n934) );
  INV_X1 U215 ( .A(n933), .ZN(n657) );
  AOI22_X1 U216 ( .A1(data_in[0]), .A2(n822), .B1(n932), .B2(\mem[19][0] ), 
        .ZN(n933) );
  INV_X1 U217 ( .A(n931), .ZN(n656) );
  AOI22_X1 U218 ( .A1(data_in[1]), .A2(n822), .B1(n932), .B2(\mem[19][1] ), 
        .ZN(n931) );
  INV_X1 U219 ( .A(n930), .ZN(n655) );
  AOI22_X1 U220 ( .A1(data_in[2]), .A2(n822), .B1(n932), .B2(\mem[19][2] ), 
        .ZN(n930) );
  INV_X1 U221 ( .A(n929), .ZN(n654) );
  AOI22_X1 U222 ( .A1(data_in[3]), .A2(n822), .B1(n932), .B2(\mem[19][3] ), 
        .ZN(n929) );
  INV_X1 U223 ( .A(n928), .ZN(n653) );
  AOI22_X1 U224 ( .A1(data_in[4]), .A2(n822), .B1(n932), .B2(\mem[19][4] ), 
        .ZN(n928) );
  INV_X1 U225 ( .A(n927), .ZN(n652) );
  AOI22_X1 U226 ( .A1(data_in[5]), .A2(n822), .B1(n932), .B2(\mem[19][5] ), 
        .ZN(n927) );
  INV_X1 U227 ( .A(n926), .ZN(n651) );
  AOI22_X1 U228 ( .A1(data_in[6]), .A2(n822), .B1(n932), .B2(\mem[19][6] ), 
        .ZN(n926) );
  INV_X1 U229 ( .A(n925), .ZN(n650) );
  AOI22_X1 U230 ( .A1(data_in[7]), .A2(n822), .B1(n932), .B2(\mem[19][7] ), 
        .ZN(n925) );
  INV_X1 U231 ( .A(n906), .ZN(n633) );
  AOI22_X1 U232 ( .A1(data_in[0]), .A2(n819), .B1(n905), .B2(\mem[22][0] ), 
        .ZN(n906) );
  INV_X1 U233 ( .A(n904), .ZN(n632) );
  AOI22_X1 U234 ( .A1(data_in[1]), .A2(n819), .B1(n905), .B2(\mem[22][1] ), 
        .ZN(n904) );
  INV_X1 U235 ( .A(n903), .ZN(n631) );
  AOI22_X1 U236 ( .A1(data_in[2]), .A2(n819), .B1(n905), .B2(\mem[22][2] ), 
        .ZN(n903) );
  INV_X1 U237 ( .A(n902), .ZN(n630) );
  AOI22_X1 U238 ( .A1(data_in[3]), .A2(n819), .B1(n905), .B2(\mem[22][3] ), 
        .ZN(n902) );
  INV_X1 U239 ( .A(n901), .ZN(n629) );
  AOI22_X1 U240 ( .A1(data_in[4]), .A2(n819), .B1(n905), .B2(\mem[22][4] ), 
        .ZN(n901) );
  INV_X1 U241 ( .A(n900), .ZN(n628) );
  AOI22_X1 U242 ( .A1(data_in[5]), .A2(n819), .B1(n905), .B2(\mem[22][5] ), 
        .ZN(n900) );
  INV_X1 U243 ( .A(n899), .ZN(n627) );
  AOI22_X1 U244 ( .A1(data_in[6]), .A2(n819), .B1(n905), .B2(\mem[22][6] ), 
        .ZN(n899) );
  INV_X1 U245 ( .A(n898), .ZN(n626) );
  AOI22_X1 U246 ( .A1(data_in[7]), .A2(n819), .B1(n905), .B2(\mem[22][7] ), 
        .ZN(n898) );
  INV_X1 U247 ( .A(n897), .ZN(n625) );
  AOI22_X1 U248 ( .A1(data_in[0]), .A2(n818), .B1(n896), .B2(\mem[23][0] ), 
        .ZN(n897) );
  INV_X1 U249 ( .A(n895), .ZN(n624) );
  AOI22_X1 U250 ( .A1(data_in[1]), .A2(n818), .B1(n896), .B2(\mem[23][1] ), 
        .ZN(n895) );
  INV_X1 U251 ( .A(n894), .ZN(n623) );
  AOI22_X1 U252 ( .A1(data_in[2]), .A2(n818), .B1(n896), .B2(\mem[23][2] ), 
        .ZN(n894) );
  INV_X1 U253 ( .A(n893), .ZN(n622) );
  AOI22_X1 U254 ( .A1(data_in[3]), .A2(n818), .B1(n896), .B2(\mem[23][3] ), 
        .ZN(n893) );
  INV_X1 U255 ( .A(n892), .ZN(n621) );
  AOI22_X1 U256 ( .A1(data_in[4]), .A2(n818), .B1(n896), .B2(\mem[23][4] ), 
        .ZN(n892) );
  INV_X1 U257 ( .A(n891), .ZN(n620) );
  AOI22_X1 U258 ( .A1(data_in[5]), .A2(n818), .B1(n896), .B2(\mem[23][5] ), 
        .ZN(n891) );
  INV_X1 U259 ( .A(n890), .ZN(n619) );
  AOI22_X1 U260 ( .A1(data_in[6]), .A2(n818), .B1(n896), .B2(\mem[23][6] ), 
        .ZN(n890) );
  INV_X1 U261 ( .A(n889), .ZN(n618) );
  AOI22_X1 U262 ( .A1(data_in[7]), .A2(n818), .B1(n896), .B2(\mem[23][7] ), 
        .ZN(n889) );
  INV_X1 U263 ( .A(n1019), .ZN(n733) );
  AOI22_X1 U264 ( .A1(data_in[4]), .A2(n832), .B1(n1023), .B2(\mem[9][4] ), 
        .ZN(n1019) );
  INV_X1 U265 ( .A(n1052), .ZN(n761) );
  AOI22_X1 U266 ( .A1(data_in[0]), .A2(n835), .B1(n1051), .B2(\mem[6][0] ), 
        .ZN(n1052) );
  INV_X1 U267 ( .A(n1050), .ZN(n760) );
  AOI22_X1 U268 ( .A1(data_in[1]), .A2(n835), .B1(n1051), .B2(\mem[6][1] ), 
        .ZN(n1050) );
  INV_X1 U269 ( .A(n1049), .ZN(n759) );
  AOI22_X1 U270 ( .A1(data_in[2]), .A2(n835), .B1(n1051), .B2(\mem[6][2] ), 
        .ZN(n1049) );
  INV_X1 U271 ( .A(n1048), .ZN(n758) );
  AOI22_X1 U272 ( .A1(data_in[3]), .A2(n835), .B1(n1051), .B2(\mem[6][3] ), 
        .ZN(n1048) );
  INV_X1 U273 ( .A(n1047), .ZN(n757) );
  AOI22_X1 U274 ( .A1(data_in[4]), .A2(n835), .B1(n1051), .B2(\mem[6][4] ), 
        .ZN(n1047) );
  INV_X1 U275 ( .A(n1046), .ZN(n756) );
  AOI22_X1 U276 ( .A1(data_in[5]), .A2(n835), .B1(n1051), .B2(\mem[6][5] ), 
        .ZN(n1046) );
  INV_X1 U277 ( .A(n1045), .ZN(n755) );
  AOI22_X1 U278 ( .A1(data_in[6]), .A2(n835), .B1(n1051), .B2(\mem[6][6] ), 
        .ZN(n1045) );
  INV_X1 U279 ( .A(n1044), .ZN(n754) );
  AOI22_X1 U280 ( .A1(data_in[7]), .A2(n835), .B1(n1051), .B2(\mem[6][7] ), 
        .ZN(n1044) );
  INV_X1 U281 ( .A(n1043), .ZN(n753) );
  AOI22_X1 U282 ( .A1(data_in[0]), .A2(n834), .B1(n1042), .B2(\mem[7][0] ), 
        .ZN(n1043) );
  INV_X1 U283 ( .A(n1041), .ZN(n752) );
  AOI22_X1 U284 ( .A1(data_in[1]), .A2(n834), .B1(n1042), .B2(\mem[7][1] ), 
        .ZN(n1041) );
  INV_X1 U285 ( .A(n1040), .ZN(n751) );
  AOI22_X1 U286 ( .A1(data_in[2]), .A2(n834), .B1(n1042), .B2(\mem[7][2] ), 
        .ZN(n1040) );
  INV_X1 U287 ( .A(n1039), .ZN(n750) );
  AOI22_X1 U288 ( .A1(data_in[3]), .A2(n834), .B1(n1042), .B2(\mem[7][3] ), 
        .ZN(n1039) );
  INV_X1 U289 ( .A(n1038), .ZN(n749) );
  AOI22_X1 U290 ( .A1(data_in[4]), .A2(n834), .B1(n1042), .B2(\mem[7][4] ), 
        .ZN(n1038) );
  INV_X1 U291 ( .A(n1037), .ZN(n748) );
  AOI22_X1 U292 ( .A1(data_in[5]), .A2(n834), .B1(n1042), .B2(\mem[7][5] ), 
        .ZN(n1037) );
  INV_X1 U293 ( .A(n1036), .ZN(n747) );
  AOI22_X1 U294 ( .A1(data_in[6]), .A2(n834), .B1(n1042), .B2(\mem[7][6] ), 
        .ZN(n1036) );
  INV_X1 U295 ( .A(n1035), .ZN(n746) );
  AOI22_X1 U296 ( .A1(data_in[7]), .A2(n834), .B1(n1042), .B2(\mem[7][7] ), 
        .ZN(n1035) );
  INV_X1 U297 ( .A(n1015), .ZN(n729) );
  AOI22_X1 U298 ( .A1(data_in[0]), .A2(n831), .B1(n1014), .B2(\mem[10][0] ), 
        .ZN(n1015) );
  INV_X1 U299 ( .A(n1013), .ZN(n728) );
  AOI22_X1 U300 ( .A1(data_in[1]), .A2(n831), .B1(n1014), .B2(\mem[10][1] ), 
        .ZN(n1013) );
  INV_X1 U301 ( .A(n1012), .ZN(n727) );
  AOI22_X1 U302 ( .A1(data_in[2]), .A2(n831), .B1(n1014), .B2(\mem[10][2] ), 
        .ZN(n1012) );
  INV_X1 U303 ( .A(n1011), .ZN(n726) );
  AOI22_X1 U304 ( .A1(data_in[3]), .A2(n831), .B1(n1014), .B2(\mem[10][3] ), 
        .ZN(n1011) );
  INV_X1 U305 ( .A(n1010), .ZN(n725) );
  AOI22_X1 U306 ( .A1(data_in[4]), .A2(n831), .B1(n1014), .B2(\mem[10][4] ), 
        .ZN(n1010) );
  INV_X1 U307 ( .A(n1009), .ZN(n724) );
  AOI22_X1 U308 ( .A1(data_in[5]), .A2(n831), .B1(n1014), .B2(\mem[10][5] ), 
        .ZN(n1009) );
  INV_X1 U309 ( .A(n1008), .ZN(n723) );
  AOI22_X1 U310 ( .A1(data_in[6]), .A2(n831), .B1(n1014), .B2(\mem[10][6] ), 
        .ZN(n1008) );
  INV_X1 U311 ( .A(n1007), .ZN(n722) );
  AOI22_X1 U312 ( .A1(data_in[7]), .A2(n831), .B1(n1014), .B2(\mem[10][7] ), 
        .ZN(n1007) );
  INV_X1 U313 ( .A(n1006), .ZN(n721) );
  AOI22_X1 U314 ( .A1(data_in[0]), .A2(n830), .B1(n1005), .B2(\mem[11][0] ), 
        .ZN(n1006) );
  INV_X1 U315 ( .A(n1004), .ZN(n720) );
  AOI22_X1 U316 ( .A1(data_in[1]), .A2(n830), .B1(n1005), .B2(\mem[11][1] ), 
        .ZN(n1004) );
  INV_X1 U317 ( .A(n1003), .ZN(n719) );
  AOI22_X1 U318 ( .A1(data_in[2]), .A2(n830), .B1(n1005), .B2(\mem[11][2] ), 
        .ZN(n1003) );
  INV_X1 U319 ( .A(n1002), .ZN(n718) );
  AOI22_X1 U320 ( .A1(data_in[3]), .A2(n830), .B1(n1005), .B2(\mem[11][3] ), 
        .ZN(n1002) );
  INV_X1 U321 ( .A(n1001), .ZN(n717) );
  AOI22_X1 U322 ( .A1(data_in[4]), .A2(n830), .B1(n1005), .B2(\mem[11][4] ), 
        .ZN(n1001) );
  INV_X1 U323 ( .A(n1000), .ZN(n716) );
  AOI22_X1 U324 ( .A1(data_in[5]), .A2(n830), .B1(n1005), .B2(\mem[11][5] ), 
        .ZN(n1000) );
  INV_X1 U325 ( .A(n999), .ZN(n715) );
  AOI22_X1 U326 ( .A1(data_in[6]), .A2(n830), .B1(n1005), .B2(\mem[11][6] ), 
        .ZN(n999) );
  INV_X1 U327 ( .A(n998), .ZN(n714) );
  AOI22_X1 U328 ( .A1(data_in[7]), .A2(n830), .B1(n1005), .B2(\mem[11][7] ), 
        .ZN(n998) );
  INV_X1 U329 ( .A(N12), .ZN(n253) );
  INV_X1 U330 ( .A(N11), .ZN(n252) );
  INV_X1 U331 ( .A(n997), .ZN(n713) );
  AOI22_X1 U332 ( .A1(data_in[0]), .A2(n829), .B1(n996), .B2(\mem[12][0] ), 
        .ZN(n997) );
  INV_X1 U333 ( .A(n995), .ZN(n712) );
  AOI22_X1 U334 ( .A1(data_in[1]), .A2(n829), .B1(n996), .B2(\mem[12][1] ), 
        .ZN(n995) );
  INV_X1 U335 ( .A(n994), .ZN(n711) );
  AOI22_X1 U336 ( .A1(data_in[2]), .A2(n829), .B1(n996), .B2(\mem[12][2] ), 
        .ZN(n994) );
  INV_X1 U337 ( .A(n993), .ZN(n710) );
  AOI22_X1 U338 ( .A1(data_in[3]), .A2(n829), .B1(n996), .B2(\mem[12][3] ), 
        .ZN(n993) );
  INV_X1 U339 ( .A(n992), .ZN(n709) );
  AOI22_X1 U340 ( .A1(data_in[4]), .A2(n829), .B1(n996), .B2(\mem[12][4] ), 
        .ZN(n992) );
  INV_X1 U341 ( .A(n991), .ZN(n708) );
  AOI22_X1 U342 ( .A1(data_in[5]), .A2(n829), .B1(n996), .B2(\mem[12][5] ), 
        .ZN(n991) );
  INV_X1 U343 ( .A(n990), .ZN(n707) );
  AOI22_X1 U344 ( .A1(data_in[6]), .A2(n829), .B1(n996), .B2(\mem[12][6] ), 
        .ZN(n990) );
  INV_X1 U345 ( .A(n989), .ZN(n706) );
  AOI22_X1 U346 ( .A1(data_in[7]), .A2(n829), .B1(n996), .B2(\mem[12][7] ), 
        .ZN(n989) );
  INV_X1 U347 ( .A(n924), .ZN(n649) );
  AOI22_X1 U348 ( .A1(data_in[0]), .A2(n821), .B1(n923), .B2(\mem[20][0] ), 
        .ZN(n924) );
  INV_X1 U349 ( .A(n922), .ZN(n648) );
  AOI22_X1 U350 ( .A1(data_in[1]), .A2(n821), .B1(n923), .B2(\mem[20][1] ), 
        .ZN(n922) );
  INV_X1 U351 ( .A(n921), .ZN(n647) );
  AOI22_X1 U352 ( .A1(data_in[2]), .A2(n821), .B1(n923), .B2(\mem[20][2] ), 
        .ZN(n921) );
  INV_X1 U353 ( .A(n920), .ZN(n646) );
  AOI22_X1 U354 ( .A1(data_in[3]), .A2(n821), .B1(n923), .B2(\mem[20][3] ), 
        .ZN(n920) );
  INV_X1 U355 ( .A(n919), .ZN(n645) );
  AOI22_X1 U356 ( .A1(data_in[4]), .A2(n821), .B1(n923), .B2(\mem[20][4] ), 
        .ZN(n919) );
  INV_X1 U357 ( .A(n918), .ZN(n644) );
  AOI22_X1 U358 ( .A1(data_in[5]), .A2(n821), .B1(n923), .B2(\mem[20][5] ), 
        .ZN(n918) );
  INV_X1 U359 ( .A(n917), .ZN(n643) );
  AOI22_X1 U360 ( .A1(data_in[6]), .A2(n821), .B1(n923), .B2(\mem[20][6] ), 
        .ZN(n917) );
  INV_X1 U361 ( .A(n916), .ZN(n642) );
  AOI22_X1 U362 ( .A1(data_in[7]), .A2(n821), .B1(n923), .B2(\mem[20][7] ), 
        .ZN(n916) );
  INV_X1 U363 ( .A(n1034), .ZN(n745) );
  AOI22_X1 U364 ( .A1(data_in[0]), .A2(n833), .B1(n1033), .B2(\mem[8][0] ), 
        .ZN(n1034) );
  INV_X1 U365 ( .A(n1032), .ZN(n744) );
  AOI22_X1 U366 ( .A1(data_in[1]), .A2(n833), .B1(n1033), .B2(\mem[8][1] ), 
        .ZN(n1032) );
  INV_X1 U367 ( .A(n1031), .ZN(n743) );
  AOI22_X1 U368 ( .A1(data_in[2]), .A2(n833), .B1(n1033), .B2(\mem[8][2] ), 
        .ZN(n1031) );
  INV_X1 U369 ( .A(n1030), .ZN(n742) );
  AOI22_X1 U370 ( .A1(data_in[3]), .A2(n833), .B1(n1033), .B2(\mem[8][3] ), 
        .ZN(n1030) );
  INV_X1 U371 ( .A(n1029), .ZN(n741) );
  AOI22_X1 U372 ( .A1(data_in[4]), .A2(n833), .B1(n1033), .B2(\mem[8][4] ), 
        .ZN(n1029) );
  INV_X1 U373 ( .A(n1028), .ZN(n740) );
  AOI22_X1 U374 ( .A1(data_in[5]), .A2(n833), .B1(n1033), .B2(\mem[8][5] ), 
        .ZN(n1028) );
  INV_X1 U375 ( .A(n1027), .ZN(n739) );
  AOI22_X1 U376 ( .A1(data_in[6]), .A2(n833), .B1(n1033), .B2(\mem[8][6] ), 
        .ZN(n1027) );
  INV_X1 U377 ( .A(n1026), .ZN(n738) );
  AOI22_X1 U378 ( .A1(data_in[7]), .A2(n833), .B1(n1033), .B2(\mem[8][7] ), 
        .ZN(n1026) );
  INV_X1 U379 ( .A(n961), .ZN(n681) );
  AOI22_X1 U380 ( .A1(data_in[0]), .A2(n825), .B1(n960), .B2(\mem[16][0] ), 
        .ZN(n961) );
  INV_X1 U381 ( .A(n959), .ZN(n680) );
  AOI22_X1 U382 ( .A1(data_in[1]), .A2(n825), .B1(n960), .B2(\mem[16][1] ), 
        .ZN(n959) );
  INV_X1 U383 ( .A(n958), .ZN(n679) );
  AOI22_X1 U384 ( .A1(data_in[2]), .A2(n825), .B1(n960), .B2(\mem[16][2] ), 
        .ZN(n958) );
  INV_X1 U385 ( .A(n957), .ZN(n678) );
  AOI22_X1 U386 ( .A1(data_in[3]), .A2(n825), .B1(n960), .B2(\mem[16][3] ), 
        .ZN(n957) );
  INV_X1 U387 ( .A(n956), .ZN(n677) );
  AOI22_X1 U388 ( .A1(data_in[4]), .A2(n825), .B1(n960), .B2(\mem[16][4] ), 
        .ZN(n956) );
  INV_X1 U389 ( .A(n955), .ZN(n676) );
  AOI22_X1 U390 ( .A1(data_in[5]), .A2(n825), .B1(n960), .B2(\mem[16][5] ), 
        .ZN(n955) );
  INV_X1 U391 ( .A(n954), .ZN(n675) );
  AOI22_X1 U392 ( .A1(data_in[6]), .A2(n825), .B1(n960), .B2(\mem[16][6] ), 
        .ZN(n954) );
  INV_X1 U393 ( .A(n953), .ZN(n674) );
  AOI22_X1 U394 ( .A1(data_in[7]), .A2(n825), .B1(n960), .B2(\mem[16][7] ), 
        .ZN(n953) );
  INV_X1 U395 ( .A(n888), .ZN(n617) );
  AOI22_X1 U396 ( .A1(data_in[0]), .A2(n814), .B1(n887), .B2(\mem[24][0] ), 
        .ZN(n888) );
  INV_X1 U397 ( .A(n886), .ZN(n616) );
  AOI22_X1 U398 ( .A1(data_in[1]), .A2(n814), .B1(n887), .B2(\mem[24][1] ), 
        .ZN(n886) );
  INV_X1 U399 ( .A(n885), .ZN(n615) );
  AOI22_X1 U400 ( .A1(data_in[2]), .A2(n814), .B1(n887), .B2(\mem[24][2] ), 
        .ZN(n885) );
  INV_X1 U401 ( .A(n884), .ZN(n614) );
  AOI22_X1 U402 ( .A1(data_in[3]), .A2(n814), .B1(n887), .B2(\mem[24][3] ), 
        .ZN(n884) );
  INV_X1 U403 ( .A(n883), .ZN(n613) );
  AOI22_X1 U404 ( .A1(data_in[4]), .A2(n814), .B1(n887), .B2(\mem[24][4] ), 
        .ZN(n883) );
  INV_X1 U405 ( .A(n882), .ZN(n612) );
  AOI22_X1 U406 ( .A1(data_in[5]), .A2(n814), .B1(n887), .B2(\mem[24][5] ), 
        .ZN(n882) );
  INV_X1 U407 ( .A(n881), .ZN(n611) );
  AOI22_X1 U408 ( .A1(data_in[6]), .A2(n814), .B1(n887), .B2(\mem[24][6] ), 
        .ZN(n881) );
  INV_X1 U409 ( .A(n880), .ZN(n610) );
  AOI22_X1 U410 ( .A1(data_in[7]), .A2(n814), .B1(n887), .B2(\mem[24][7] ), 
        .ZN(n880) );
  INV_X1 U411 ( .A(n879), .ZN(n609) );
  AOI22_X1 U412 ( .A1(data_in[0]), .A2(n813), .B1(n878), .B2(\mem[25][0] ), 
        .ZN(n879) );
  INV_X1 U413 ( .A(n877), .ZN(n608) );
  AOI22_X1 U414 ( .A1(data_in[1]), .A2(n813), .B1(n878), .B2(\mem[25][1] ), 
        .ZN(n877) );
  INV_X1 U415 ( .A(n876), .ZN(n607) );
  AOI22_X1 U416 ( .A1(data_in[2]), .A2(n813), .B1(n878), .B2(\mem[25][2] ), 
        .ZN(n876) );
  INV_X1 U417 ( .A(n875), .ZN(n606) );
  AOI22_X1 U418 ( .A1(data_in[3]), .A2(n813), .B1(n878), .B2(\mem[25][3] ), 
        .ZN(n875) );
  INV_X1 U419 ( .A(n874), .ZN(n605) );
  AOI22_X1 U420 ( .A1(data_in[4]), .A2(n813), .B1(n878), .B2(\mem[25][4] ), 
        .ZN(n874) );
  INV_X1 U421 ( .A(n873), .ZN(n604) );
  AOI22_X1 U422 ( .A1(data_in[5]), .A2(n813), .B1(n878), .B2(\mem[25][5] ), 
        .ZN(n873) );
  INV_X1 U423 ( .A(n872), .ZN(n603) );
  AOI22_X1 U424 ( .A1(data_in[6]), .A2(n813), .B1(n878), .B2(\mem[25][6] ), 
        .ZN(n872) );
  INV_X1 U425 ( .A(n871), .ZN(n602) );
  AOI22_X1 U426 ( .A1(data_in[7]), .A2(n813), .B1(n878), .B2(\mem[25][7] ), 
        .ZN(n871) );
  INV_X1 U427 ( .A(n870), .ZN(n601) );
  AOI22_X1 U428 ( .A1(data_in[0]), .A2(n812), .B1(n869), .B2(\mem[26][0] ), 
        .ZN(n870) );
  INV_X1 U429 ( .A(n868), .ZN(n600) );
  AOI22_X1 U430 ( .A1(data_in[1]), .A2(n812), .B1(n869), .B2(\mem[26][1] ), 
        .ZN(n868) );
  INV_X1 U431 ( .A(n867), .ZN(n599) );
  AOI22_X1 U432 ( .A1(data_in[2]), .A2(n812), .B1(n869), .B2(\mem[26][2] ), 
        .ZN(n867) );
  INV_X1 U433 ( .A(n866), .ZN(n598) );
  AOI22_X1 U434 ( .A1(data_in[3]), .A2(n812), .B1(n869), .B2(\mem[26][3] ), 
        .ZN(n866) );
  INV_X1 U435 ( .A(n865), .ZN(n597) );
  AOI22_X1 U436 ( .A1(data_in[4]), .A2(n812), .B1(n869), .B2(\mem[26][4] ), 
        .ZN(n865) );
  INV_X1 U437 ( .A(n864), .ZN(n596) );
  AOI22_X1 U438 ( .A1(data_in[5]), .A2(n812), .B1(n869), .B2(\mem[26][5] ), 
        .ZN(n864) );
  INV_X1 U439 ( .A(n863), .ZN(n595) );
  AOI22_X1 U440 ( .A1(data_in[6]), .A2(n812), .B1(n869), .B2(\mem[26][6] ), 
        .ZN(n863) );
  INV_X1 U441 ( .A(n862), .ZN(n594) );
  AOI22_X1 U442 ( .A1(data_in[7]), .A2(n812), .B1(n869), .B2(\mem[26][7] ), 
        .ZN(n862) );
  INV_X1 U443 ( .A(n861), .ZN(n293) );
  AOI22_X1 U444 ( .A1(data_in[0]), .A2(n811), .B1(n860), .B2(\mem[27][0] ), 
        .ZN(n861) );
  INV_X1 U445 ( .A(n859), .ZN(n292) );
  AOI22_X1 U446 ( .A1(data_in[1]), .A2(n811), .B1(n860), .B2(\mem[27][1] ), 
        .ZN(n859) );
  INV_X1 U447 ( .A(n858), .ZN(n291) );
  AOI22_X1 U448 ( .A1(data_in[2]), .A2(n811), .B1(n860), .B2(\mem[27][2] ), 
        .ZN(n858) );
  INV_X1 U449 ( .A(n857), .ZN(n290) );
  AOI22_X1 U450 ( .A1(data_in[3]), .A2(n811), .B1(n860), .B2(\mem[27][3] ), 
        .ZN(n857) );
  INV_X1 U451 ( .A(n856), .ZN(n289) );
  AOI22_X1 U452 ( .A1(data_in[4]), .A2(n811), .B1(n860), .B2(\mem[27][4] ), 
        .ZN(n856) );
  INV_X1 U453 ( .A(n855), .ZN(n288) );
  AOI22_X1 U454 ( .A1(data_in[5]), .A2(n811), .B1(n860), .B2(\mem[27][5] ), 
        .ZN(n855) );
  INV_X1 U455 ( .A(n854), .ZN(n287) );
  AOI22_X1 U456 ( .A1(data_in[6]), .A2(n811), .B1(n860), .B2(\mem[27][6] ), 
        .ZN(n854) );
  INV_X1 U457 ( .A(n853), .ZN(n286) );
  AOI22_X1 U458 ( .A1(data_in[7]), .A2(n811), .B1(n860), .B2(\mem[27][7] ), 
        .ZN(n853) );
  INV_X1 U459 ( .A(n852), .ZN(n285) );
  AOI22_X1 U460 ( .A1(data_in[0]), .A2(n810), .B1(n851), .B2(\mem[28][0] ), 
        .ZN(n852) );
  INV_X1 U461 ( .A(n850), .ZN(n284) );
  AOI22_X1 U462 ( .A1(data_in[1]), .A2(n810), .B1(n851), .B2(\mem[28][1] ), 
        .ZN(n850) );
  INV_X1 U463 ( .A(n849), .ZN(n283) );
  AOI22_X1 U464 ( .A1(data_in[2]), .A2(n810), .B1(n851), .B2(\mem[28][2] ), 
        .ZN(n849) );
  INV_X1 U465 ( .A(n848), .ZN(n282) );
  AOI22_X1 U466 ( .A1(data_in[3]), .A2(n810), .B1(n851), .B2(\mem[28][3] ), 
        .ZN(n848) );
  INV_X1 U467 ( .A(n847), .ZN(n281) );
  AOI22_X1 U468 ( .A1(data_in[4]), .A2(n810), .B1(n851), .B2(\mem[28][4] ), 
        .ZN(n847) );
  INV_X1 U469 ( .A(n846), .ZN(n280) );
  AOI22_X1 U470 ( .A1(data_in[5]), .A2(n810), .B1(n851), .B2(\mem[28][5] ), 
        .ZN(n846) );
  INV_X1 U471 ( .A(n845), .ZN(n279) );
  AOI22_X1 U472 ( .A1(data_in[6]), .A2(n810), .B1(n851), .B2(\mem[28][6] ), 
        .ZN(n845) );
  INV_X1 U473 ( .A(n844), .ZN(n278) );
  AOI22_X1 U474 ( .A1(data_in[7]), .A2(n810), .B1(n851), .B2(\mem[28][7] ), 
        .ZN(n844) );
  INV_X1 U475 ( .A(n1143), .ZN(n277) );
  AOI22_X1 U476 ( .A1(n817), .A2(data_in[0]), .B1(n1142), .B2(\mem[29][0] ), 
        .ZN(n1143) );
  INV_X1 U477 ( .A(n1141), .ZN(n276) );
  AOI22_X1 U478 ( .A1(n817), .A2(data_in[1]), .B1(n1142), .B2(\mem[29][1] ), 
        .ZN(n1141) );
  INV_X1 U479 ( .A(n1140), .ZN(n275) );
  AOI22_X1 U480 ( .A1(n817), .A2(data_in[2]), .B1(n1142), .B2(\mem[29][2] ), 
        .ZN(n1140) );
  INV_X1 U481 ( .A(n1139), .ZN(n274) );
  AOI22_X1 U482 ( .A1(n817), .A2(data_in[3]), .B1(n1142), .B2(\mem[29][3] ), 
        .ZN(n1139) );
  INV_X1 U483 ( .A(n1138), .ZN(n273) );
  AOI22_X1 U484 ( .A1(n817), .A2(data_in[4]), .B1(n1142), .B2(\mem[29][4] ), 
        .ZN(n1138) );
  INV_X1 U485 ( .A(n1137), .ZN(n272) );
  AOI22_X1 U486 ( .A1(n817), .A2(data_in[5]), .B1(n1142), .B2(\mem[29][5] ), 
        .ZN(n1137) );
  INV_X1 U487 ( .A(n1136), .ZN(n271) );
  AOI22_X1 U488 ( .A1(n817), .A2(data_in[6]), .B1(n1142), .B2(\mem[29][6] ), 
        .ZN(n1136) );
  INV_X1 U489 ( .A(n1135), .ZN(n270) );
  AOI22_X1 U490 ( .A1(n817), .A2(data_in[7]), .B1(n1142), .B2(\mem[29][7] ), 
        .ZN(n1135) );
  INV_X1 U491 ( .A(n1132), .ZN(n269) );
  AOI22_X1 U492 ( .A1(data_in[0]), .A2(n816), .B1(n1131), .B2(\mem[30][0] ), 
        .ZN(n1132) );
  INV_X1 U493 ( .A(n1130), .ZN(n268) );
  AOI22_X1 U494 ( .A1(data_in[1]), .A2(n816), .B1(n1131), .B2(\mem[30][1] ), 
        .ZN(n1130) );
  INV_X1 U495 ( .A(n1129), .ZN(n267) );
  AOI22_X1 U496 ( .A1(data_in[2]), .A2(n816), .B1(n1131), .B2(\mem[30][2] ), 
        .ZN(n1129) );
  INV_X1 U497 ( .A(n1128), .ZN(n266) );
  AOI22_X1 U498 ( .A1(data_in[3]), .A2(n816), .B1(n1131), .B2(\mem[30][3] ), 
        .ZN(n1128) );
  INV_X1 U499 ( .A(n1127), .ZN(n265) );
  AOI22_X1 U500 ( .A1(data_in[4]), .A2(n816), .B1(n1131), .B2(\mem[30][4] ), 
        .ZN(n1127) );
  INV_X1 U501 ( .A(n1126), .ZN(n264) );
  AOI22_X1 U502 ( .A1(data_in[5]), .A2(n816), .B1(n1131), .B2(\mem[30][5] ), 
        .ZN(n1126) );
  INV_X1 U503 ( .A(n1125), .ZN(n263) );
  AOI22_X1 U504 ( .A1(data_in[6]), .A2(n816), .B1(n1131), .B2(\mem[30][6] ), 
        .ZN(n1125) );
  INV_X1 U505 ( .A(n1124), .ZN(n262) );
  AOI22_X1 U506 ( .A1(data_in[7]), .A2(n816), .B1(n1131), .B2(\mem[30][7] ), 
        .ZN(n1124) );
  INV_X1 U507 ( .A(n1122), .ZN(n261) );
  AOI22_X1 U508 ( .A1(data_in[0]), .A2(n815), .B1(n1121), .B2(\mem[31][0] ), 
        .ZN(n1122) );
  INV_X1 U509 ( .A(n1120), .ZN(n260) );
  AOI22_X1 U510 ( .A1(data_in[1]), .A2(n815), .B1(n1121), .B2(\mem[31][1] ), 
        .ZN(n1120) );
  INV_X1 U511 ( .A(n1119), .ZN(n259) );
  AOI22_X1 U512 ( .A1(data_in[2]), .A2(n815), .B1(n1121), .B2(\mem[31][2] ), 
        .ZN(n1119) );
  INV_X1 U513 ( .A(n1118), .ZN(n258) );
  AOI22_X1 U514 ( .A1(data_in[3]), .A2(n815), .B1(n1121), .B2(\mem[31][3] ), 
        .ZN(n1118) );
  INV_X1 U515 ( .A(n1117), .ZN(n257) );
  AOI22_X1 U516 ( .A1(data_in[4]), .A2(n815), .B1(n1121), .B2(\mem[31][4] ), 
        .ZN(n1117) );
  INV_X1 U517 ( .A(n1116), .ZN(n256) );
  AOI22_X1 U518 ( .A1(data_in[5]), .A2(n815), .B1(n1121), .B2(\mem[31][5] ), 
        .ZN(n1116) );
  INV_X1 U519 ( .A(n1115), .ZN(n255) );
  AOI22_X1 U520 ( .A1(data_in[6]), .A2(n815), .B1(n1121), .B2(\mem[31][6] ), 
        .ZN(n1115) );
  INV_X1 U521 ( .A(n1114), .ZN(n254) );
  AOI22_X1 U522 ( .A1(data_in[7]), .A2(n815), .B1(n1121), .B2(\mem[31][7] ), 
        .ZN(n1114) );
  INV_X1 U523 ( .A(n1112), .ZN(n809) );
  AOI22_X1 U524 ( .A1(data_in[0]), .A2(n841), .B1(n1111), .B2(\mem[0][0] ), 
        .ZN(n1112) );
  INV_X1 U525 ( .A(n1110), .ZN(n808) );
  AOI22_X1 U526 ( .A1(data_in[1]), .A2(n841), .B1(n1111), .B2(\mem[0][1] ), 
        .ZN(n1110) );
  INV_X1 U527 ( .A(n1109), .ZN(n807) );
  AOI22_X1 U528 ( .A1(data_in[2]), .A2(n841), .B1(n1111), .B2(\mem[0][2] ), 
        .ZN(n1109) );
  INV_X1 U529 ( .A(n1108), .ZN(n806) );
  AOI22_X1 U530 ( .A1(data_in[3]), .A2(n841), .B1(n1111), .B2(\mem[0][3] ), 
        .ZN(n1108) );
  INV_X1 U531 ( .A(n1107), .ZN(n805) );
  AOI22_X1 U532 ( .A1(data_in[4]), .A2(n841), .B1(n1111), .B2(\mem[0][4] ), 
        .ZN(n1107) );
  INV_X1 U533 ( .A(n1106), .ZN(n804) );
  AOI22_X1 U534 ( .A1(data_in[5]), .A2(n841), .B1(n1111), .B2(\mem[0][5] ), 
        .ZN(n1106) );
  INV_X1 U535 ( .A(n1105), .ZN(n803) );
  AOI22_X1 U536 ( .A1(data_in[6]), .A2(n841), .B1(n1111), .B2(\mem[0][6] ), 
        .ZN(n1105) );
  INV_X1 U537 ( .A(n1104), .ZN(n802) );
  AOI22_X1 U538 ( .A1(data_in[7]), .A2(n841), .B1(n1111), .B2(\mem[0][7] ), 
        .ZN(n1104) );
  INV_X1 U539 ( .A(n1101), .ZN(n801) );
  AOI22_X1 U540 ( .A1(data_in[0]), .A2(n840), .B1(n1100), .B2(\mem[1][0] ), 
        .ZN(n1101) );
  INV_X1 U541 ( .A(n1099), .ZN(n800) );
  AOI22_X1 U542 ( .A1(data_in[1]), .A2(n840), .B1(n1100), .B2(\mem[1][1] ), 
        .ZN(n1099) );
  INV_X1 U543 ( .A(n1098), .ZN(n799) );
  AOI22_X1 U544 ( .A1(data_in[2]), .A2(n840), .B1(n1100), .B2(\mem[1][2] ), 
        .ZN(n1098) );
  INV_X1 U545 ( .A(n1097), .ZN(n798) );
  AOI22_X1 U546 ( .A1(data_in[3]), .A2(n840), .B1(n1100), .B2(\mem[1][3] ), 
        .ZN(n1097) );
  INV_X1 U547 ( .A(n1096), .ZN(n797) );
  AOI22_X1 U548 ( .A1(data_in[4]), .A2(n840), .B1(n1100), .B2(\mem[1][4] ), 
        .ZN(n1096) );
  INV_X1 U549 ( .A(n1095), .ZN(n796) );
  AOI22_X1 U550 ( .A1(data_in[5]), .A2(n840), .B1(n1100), .B2(\mem[1][5] ), 
        .ZN(n1095) );
  INV_X1 U551 ( .A(n1094), .ZN(n795) );
  AOI22_X1 U552 ( .A1(data_in[6]), .A2(n840), .B1(n1100), .B2(\mem[1][6] ), 
        .ZN(n1094) );
  INV_X1 U553 ( .A(n1093), .ZN(n794) );
  AOI22_X1 U554 ( .A1(data_in[7]), .A2(n840), .B1(n1100), .B2(\mem[1][7] ), 
        .ZN(n1093) );
  INV_X1 U555 ( .A(n1091), .ZN(n793) );
  AOI22_X1 U556 ( .A1(data_in[0]), .A2(n839), .B1(n1090), .B2(\mem[2][0] ), 
        .ZN(n1091) );
  INV_X1 U557 ( .A(n1089), .ZN(n792) );
  AOI22_X1 U558 ( .A1(data_in[1]), .A2(n839), .B1(n1090), .B2(\mem[2][1] ), 
        .ZN(n1089) );
  INV_X1 U559 ( .A(n1088), .ZN(n791) );
  AOI22_X1 U560 ( .A1(data_in[2]), .A2(n839), .B1(n1090), .B2(\mem[2][2] ), 
        .ZN(n1088) );
  INV_X1 U561 ( .A(n1087), .ZN(n790) );
  AOI22_X1 U562 ( .A1(data_in[3]), .A2(n839), .B1(n1090), .B2(\mem[2][3] ), 
        .ZN(n1087) );
  INV_X1 U563 ( .A(n1086), .ZN(n789) );
  AOI22_X1 U564 ( .A1(data_in[4]), .A2(n839), .B1(n1090), .B2(\mem[2][4] ), 
        .ZN(n1086) );
  INV_X1 U565 ( .A(n1085), .ZN(n788) );
  AOI22_X1 U566 ( .A1(data_in[5]), .A2(n839), .B1(n1090), .B2(\mem[2][5] ), 
        .ZN(n1085) );
  INV_X1 U567 ( .A(n1084), .ZN(n787) );
  AOI22_X1 U568 ( .A1(data_in[6]), .A2(n839), .B1(n1090), .B2(\mem[2][6] ), 
        .ZN(n1084) );
  INV_X1 U569 ( .A(n1083), .ZN(n786) );
  AOI22_X1 U570 ( .A1(data_in[7]), .A2(n839), .B1(n1090), .B2(\mem[2][7] ), 
        .ZN(n1083) );
  INV_X1 U571 ( .A(n1081), .ZN(n785) );
  AOI22_X1 U572 ( .A1(data_in[0]), .A2(n838), .B1(n1080), .B2(\mem[3][0] ), 
        .ZN(n1081) );
  INV_X1 U573 ( .A(n1079), .ZN(n784) );
  AOI22_X1 U574 ( .A1(data_in[1]), .A2(n838), .B1(n1080), .B2(\mem[3][1] ), 
        .ZN(n1079) );
  INV_X1 U575 ( .A(n1078), .ZN(n783) );
  AOI22_X1 U576 ( .A1(data_in[2]), .A2(n838), .B1(n1080), .B2(\mem[3][2] ), 
        .ZN(n1078) );
  INV_X1 U577 ( .A(n1077), .ZN(n782) );
  AOI22_X1 U578 ( .A1(data_in[3]), .A2(n838), .B1(n1080), .B2(\mem[3][3] ), 
        .ZN(n1077) );
  INV_X1 U579 ( .A(n1076), .ZN(n781) );
  AOI22_X1 U580 ( .A1(data_in[4]), .A2(n838), .B1(n1080), .B2(\mem[3][4] ), 
        .ZN(n1076) );
  INV_X1 U581 ( .A(n1075), .ZN(n780) );
  AOI22_X1 U582 ( .A1(data_in[5]), .A2(n838), .B1(n1080), .B2(\mem[3][5] ), 
        .ZN(n1075) );
  INV_X1 U583 ( .A(n1074), .ZN(n779) );
  AOI22_X1 U584 ( .A1(data_in[6]), .A2(n838), .B1(n1080), .B2(\mem[3][6] ), 
        .ZN(n1074) );
  INV_X1 U585 ( .A(n1073), .ZN(n778) );
  AOI22_X1 U586 ( .A1(data_in[7]), .A2(n838), .B1(n1080), .B2(\mem[3][7] ), 
        .ZN(n1073) );
  INV_X1 U587 ( .A(n1071), .ZN(n777) );
  AOI22_X1 U588 ( .A1(data_in[0]), .A2(n837), .B1(n1070), .B2(\mem[4][0] ), 
        .ZN(n1071) );
  INV_X1 U589 ( .A(n1069), .ZN(n776) );
  AOI22_X1 U590 ( .A1(data_in[1]), .A2(n837), .B1(n1070), .B2(\mem[4][1] ), 
        .ZN(n1069) );
  INV_X1 U591 ( .A(n1068), .ZN(n775) );
  AOI22_X1 U592 ( .A1(data_in[2]), .A2(n837), .B1(n1070), .B2(\mem[4][2] ), 
        .ZN(n1068) );
  INV_X1 U593 ( .A(n1067), .ZN(n774) );
  AOI22_X1 U594 ( .A1(data_in[3]), .A2(n837), .B1(n1070), .B2(\mem[4][3] ), 
        .ZN(n1067) );
  INV_X1 U595 ( .A(n1066), .ZN(n773) );
  AOI22_X1 U596 ( .A1(data_in[4]), .A2(n837), .B1(n1070), .B2(\mem[4][4] ), 
        .ZN(n1066) );
  INV_X1 U597 ( .A(n1065), .ZN(n772) );
  AOI22_X1 U598 ( .A1(data_in[5]), .A2(n837), .B1(n1070), .B2(\mem[4][5] ), 
        .ZN(n1065) );
  INV_X1 U599 ( .A(n1064), .ZN(n771) );
  AOI22_X1 U600 ( .A1(data_in[6]), .A2(n837), .B1(n1070), .B2(\mem[4][6] ), 
        .ZN(n1064) );
  INV_X1 U601 ( .A(n1063), .ZN(n770) );
  AOI22_X1 U602 ( .A1(data_in[7]), .A2(n837), .B1(n1070), .B2(\mem[4][7] ), 
        .ZN(n1063) );
  INV_X1 U603 ( .A(N13), .ZN(n842) );
  INV_X1 U604 ( .A(N14), .ZN(n843) );
  MUX2_X1 U605 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n245), .Z(n1) );
  MUX2_X1 U606 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n245), .Z(n2) );
  MUX2_X1 U607 ( .A(n2), .B(n1), .S(n242), .Z(n3) );
  MUX2_X1 U608 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n245), .Z(n4) );
  MUX2_X1 U609 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n245), .Z(n5) );
  MUX2_X1 U610 ( .A(n5), .B(n4), .S(n244), .Z(n6) );
  MUX2_X1 U611 ( .A(n6), .B(n3), .S(n241), .Z(n7) );
  MUX2_X1 U612 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n245), .Z(n8) );
  MUX2_X1 U613 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n245), .Z(n9) );
  MUX2_X1 U614 ( .A(n9), .B(n8), .S(n243), .Z(n10) );
  MUX2_X1 U615 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n245), .Z(n11) );
  MUX2_X1 U616 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n245), .Z(n12) );
  MUX2_X1 U617 ( .A(n12), .B(n11), .S(n243), .Z(n13) );
  MUX2_X1 U618 ( .A(n13), .B(n10), .S(n241), .Z(n14) );
  MUX2_X1 U619 ( .A(n14), .B(n7), .S(N13), .Z(n15) );
  MUX2_X1 U620 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n246), .Z(n16) );
  MUX2_X1 U621 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n246), .Z(n17) );
  MUX2_X1 U622 ( .A(n17), .B(n16), .S(n242), .Z(n18) );
  MUX2_X1 U623 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n246), .Z(n19) );
  MUX2_X1 U624 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n246), .Z(n20) );
  MUX2_X1 U625 ( .A(n20), .B(n19), .S(n242), .Z(n21) );
  MUX2_X1 U626 ( .A(n21), .B(n18), .S(n241), .Z(n22) );
  MUX2_X1 U627 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n246), .Z(n23) );
  MUX2_X1 U628 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n246), .Z(n24) );
  MUX2_X1 U629 ( .A(n24), .B(n23), .S(n242), .Z(n25) );
  MUX2_X1 U630 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n246), .Z(n26) );
  MUX2_X1 U631 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n246), .Z(n27) );
  MUX2_X1 U632 ( .A(n27), .B(n26), .S(n242), .Z(n28) );
  MUX2_X1 U633 ( .A(n28), .B(n25), .S(n241), .Z(n29) );
  MUX2_X1 U634 ( .A(n29), .B(n22), .S(N13), .Z(n30) );
  MUX2_X1 U635 ( .A(n30), .B(n15), .S(N14), .Z(N22) );
  MUX2_X1 U636 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n246), .Z(n31) );
  MUX2_X1 U637 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n246), .Z(n32) );
  MUX2_X1 U638 ( .A(n32), .B(n31), .S(n242), .Z(n33) );
  MUX2_X1 U639 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n246), .Z(n34) );
  MUX2_X1 U640 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n246), .Z(n35) );
  MUX2_X1 U641 ( .A(n35), .B(n34), .S(n242), .Z(n36) );
  MUX2_X1 U642 ( .A(n36), .B(n33), .S(n241), .Z(n37) );
  MUX2_X1 U643 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n247), .Z(n38) );
  MUX2_X1 U644 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n247), .Z(n39) );
  MUX2_X1 U645 ( .A(n39), .B(n38), .S(n242), .Z(n40) );
  MUX2_X1 U646 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n247), .Z(n41) );
  MUX2_X1 U647 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n247), .Z(n42) );
  MUX2_X1 U648 ( .A(n42), .B(n41), .S(n242), .Z(n43) );
  MUX2_X1 U649 ( .A(n43), .B(n40), .S(N12), .Z(n44) );
  MUX2_X1 U650 ( .A(n44), .B(n37), .S(N13), .Z(n45) );
  MUX2_X1 U651 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n247), .Z(n46) );
  MUX2_X1 U652 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n247), .Z(n47) );
  MUX2_X1 U653 ( .A(n47), .B(n46), .S(n242), .Z(n48) );
  MUX2_X1 U654 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n247), .Z(n49) );
  MUX2_X1 U655 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n247), .Z(n50) );
  MUX2_X1 U656 ( .A(n50), .B(n49), .S(n242), .Z(n51) );
  MUX2_X1 U657 ( .A(n51), .B(n48), .S(N12), .Z(n52) );
  MUX2_X1 U658 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n247), .Z(n53) );
  MUX2_X1 U659 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n247), .Z(n54) );
  MUX2_X1 U660 ( .A(n54), .B(n53), .S(n242), .Z(n55) );
  MUX2_X1 U661 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n247), .Z(n56) );
  MUX2_X1 U662 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n247), .Z(n57) );
  MUX2_X1 U663 ( .A(n57), .B(n56), .S(n242), .Z(n58) );
  MUX2_X1 U664 ( .A(n58), .B(n55), .S(N12), .Z(n59) );
  MUX2_X1 U665 ( .A(n59), .B(n52), .S(N13), .Z(n60) );
  MUX2_X1 U666 ( .A(n60), .B(n45), .S(N14), .Z(N21) );
  MUX2_X1 U667 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n248), .Z(n61) );
  MUX2_X1 U668 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n248), .Z(n62) );
  MUX2_X1 U669 ( .A(n62), .B(n61), .S(n243), .Z(n63) );
  MUX2_X1 U670 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n248), .Z(n64) );
  MUX2_X1 U671 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n248), .Z(n65) );
  MUX2_X1 U672 ( .A(n65), .B(n64), .S(n243), .Z(n66) );
  MUX2_X1 U673 ( .A(n66), .B(n63), .S(n241), .Z(n67) );
  MUX2_X1 U674 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n248), .Z(n68) );
  MUX2_X1 U675 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n248), .Z(n69) );
  MUX2_X1 U676 ( .A(n69), .B(n68), .S(n243), .Z(n70) );
  MUX2_X1 U677 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n248), .Z(n71) );
  MUX2_X1 U678 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n248), .Z(n72) );
  MUX2_X1 U679 ( .A(n72), .B(n71), .S(n243), .Z(n73) );
  MUX2_X1 U680 ( .A(n73), .B(n70), .S(n241), .Z(n74) );
  MUX2_X1 U681 ( .A(n74), .B(n67), .S(N13), .Z(n75) );
  MUX2_X1 U682 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n248), .Z(n76) );
  MUX2_X1 U683 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(n248), .Z(n77) );
  MUX2_X1 U684 ( .A(n77), .B(n76), .S(n243), .Z(n78) );
  MUX2_X1 U685 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(n248), .Z(n79) );
  MUX2_X1 U686 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(n248), .Z(n80) );
  MUX2_X1 U687 ( .A(n80), .B(n79), .S(n243), .Z(n81) );
  MUX2_X1 U688 ( .A(n81), .B(n78), .S(n241), .Z(n82) );
  MUX2_X1 U689 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(n249), .Z(n83) );
  MUX2_X1 U690 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(n249), .Z(n84) );
  MUX2_X1 U691 ( .A(n84), .B(n83), .S(n243), .Z(n85) );
  MUX2_X1 U692 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(n249), .Z(n86) );
  MUX2_X1 U693 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(n249), .Z(n87) );
  MUX2_X1 U694 ( .A(n87), .B(n86), .S(n243), .Z(n88) );
  MUX2_X1 U695 ( .A(n88), .B(n85), .S(n241), .Z(n89) );
  MUX2_X1 U696 ( .A(n89), .B(n82), .S(N13), .Z(n90) );
  MUX2_X1 U697 ( .A(n90), .B(n75), .S(N14), .Z(N20) );
  MUX2_X1 U698 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n249), .Z(n91) );
  MUX2_X1 U699 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(n249), .Z(n92) );
  MUX2_X1 U700 ( .A(n92), .B(n91), .S(n243), .Z(n93) );
  MUX2_X1 U701 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n249), .Z(n94) );
  MUX2_X1 U702 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(n249), .Z(n95) );
  MUX2_X1 U703 ( .A(n95), .B(n94), .S(n243), .Z(n96) );
  MUX2_X1 U704 ( .A(n96), .B(n93), .S(n241), .Z(n97) );
  MUX2_X1 U705 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n249), .Z(n98) );
  MUX2_X1 U706 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n249), .Z(n99) );
  MUX2_X1 U707 ( .A(n99), .B(n98), .S(n243), .Z(n100) );
  MUX2_X1 U708 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n249), .Z(n101) );
  MUX2_X1 U709 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n249), .Z(n102) );
  MUX2_X1 U710 ( .A(n102), .B(n101), .S(n243), .Z(n103) );
  MUX2_X1 U711 ( .A(n103), .B(n100), .S(n241), .Z(n104) );
  MUX2_X1 U712 ( .A(n104), .B(n97), .S(N13), .Z(n105) );
  MUX2_X1 U713 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n250), .Z(n106) );
  MUX2_X1 U714 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n245), .Z(n107) );
  MUX2_X1 U715 ( .A(n107), .B(n106), .S(n244), .Z(n108) );
  MUX2_X1 U716 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n250), .Z(n109) );
  MUX2_X1 U717 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n250), .Z(n110) );
  MUX2_X1 U718 ( .A(n110), .B(n109), .S(n244), .Z(n111) );
  MUX2_X1 U719 ( .A(n111), .B(n108), .S(n241), .Z(n112) );
  MUX2_X1 U720 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n246), .Z(n113) );
  MUX2_X1 U721 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n249), .Z(n114) );
  MUX2_X1 U722 ( .A(n114), .B(n113), .S(n244), .Z(n115) );
  MUX2_X1 U723 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n246), .Z(n116) );
  MUX2_X1 U724 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n250), .Z(n117) );
  MUX2_X1 U725 ( .A(n117), .B(n116), .S(n244), .Z(n118) );
  MUX2_X1 U726 ( .A(n118), .B(n115), .S(n241), .Z(n119) );
  MUX2_X1 U727 ( .A(n119), .B(n112), .S(N13), .Z(n120) );
  MUX2_X1 U728 ( .A(n120), .B(n105), .S(N14), .Z(N19) );
  MUX2_X1 U729 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(N10), .Z(n121) );
  MUX2_X1 U730 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n249), .Z(n122) );
  MUX2_X1 U731 ( .A(n122), .B(n121), .S(n244), .Z(n123) );
  MUX2_X1 U732 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n250), .Z(n124) );
  MUX2_X1 U733 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n250), .Z(n125) );
  MUX2_X1 U734 ( .A(n125), .B(n124), .S(n244), .Z(n126) );
  MUX2_X1 U735 ( .A(n126), .B(n123), .S(n241), .Z(n127) );
  MUX2_X1 U736 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n250), .Z(n128) );
  MUX2_X1 U737 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(N10), .Z(n129) );
  MUX2_X1 U738 ( .A(n129), .B(n128), .S(n244), .Z(n130) );
  MUX2_X1 U739 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(N10), .Z(n131) );
  MUX2_X1 U740 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n250), .Z(n132) );
  MUX2_X1 U741 ( .A(n132), .B(n131), .S(n244), .Z(n133) );
  MUX2_X1 U742 ( .A(n133), .B(n130), .S(n241), .Z(n134) );
  MUX2_X1 U743 ( .A(n134), .B(n127), .S(N13), .Z(n135) );
  MUX2_X1 U744 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n247), .Z(n136) );
  MUX2_X1 U745 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(N10), .Z(n137) );
  MUX2_X1 U746 ( .A(n137), .B(n136), .S(n244), .Z(n138) );
  MUX2_X1 U747 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(N10), .Z(n139) );
  MUX2_X1 U748 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(N10), .Z(n140) );
  MUX2_X1 U749 ( .A(n140), .B(n139), .S(n244), .Z(n141) );
  MUX2_X1 U750 ( .A(n141), .B(n138), .S(n241), .Z(n142) );
  MUX2_X1 U751 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(N10), .Z(n143) );
  MUX2_X1 U752 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n247), .Z(n144) );
  MUX2_X1 U753 ( .A(n144), .B(n143), .S(n244), .Z(n145) );
  MUX2_X1 U754 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(N10), .Z(n146) );
  MUX2_X1 U755 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n245), .Z(n147) );
  MUX2_X1 U756 ( .A(n147), .B(n146), .S(n244), .Z(n148) );
  MUX2_X1 U757 ( .A(n148), .B(n145), .S(n241), .Z(n149) );
  MUX2_X1 U758 ( .A(n149), .B(n142), .S(N13), .Z(n150) );
  MUX2_X1 U759 ( .A(n150), .B(n135), .S(N14), .Z(N18) );
  MUX2_X1 U760 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n245), .Z(n151) );
  MUX2_X1 U761 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n250), .Z(n152) );
  MUX2_X1 U762 ( .A(n152), .B(n151), .S(N11), .Z(n153) );
  MUX2_X1 U763 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n245), .Z(n154) );
  MUX2_X1 U764 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(N10), .Z(n155) );
  MUX2_X1 U765 ( .A(n155), .B(n154), .S(N11), .Z(n156) );
  MUX2_X1 U766 ( .A(n156), .B(n153), .S(n241), .Z(n157) );
  MUX2_X1 U767 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(N10), .Z(n158) );
  MUX2_X1 U768 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(N10), .Z(n159) );
  MUX2_X1 U769 ( .A(n159), .B(n158), .S(N11), .Z(n160) );
  MUX2_X1 U770 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(N10), .Z(n161) );
  MUX2_X1 U771 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(N10), .Z(n162) );
  MUX2_X1 U772 ( .A(n162), .B(n161), .S(n244), .Z(n163) );
  MUX2_X1 U773 ( .A(n163), .B(n160), .S(N12), .Z(n164) );
  MUX2_X1 U774 ( .A(n164), .B(n157), .S(N13), .Z(n165) );
  MUX2_X1 U775 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n245), .Z(n166) );
  MUX2_X1 U776 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(N10), .Z(n167) );
  MUX2_X1 U777 ( .A(n167), .B(n166), .S(N11), .Z(n168) );
  MUX2_X1 U778 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n248), .Z(n169) );
  MUX2_X1 U779 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(N10), .Z(n170) );
  MUX2_X1 U780 ( .A(n170), .B(n169), .S(n242), .Z(n171) );
  MUX2_X1 U781 ( .A(n171), .B(n168), .S(n241), .Z(n172) );
  MUX2_X1 U782 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n246), .Z(n173) );
  MUX2_X1 U783 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n248), .Z(n174) );
  MUX2_X1 U784 ( .A(n174), .B(n173), .S(N11), .Z(n175) );
  MUX2_X1 U785 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n246), .Z(n176) );
  MUX2_X1 U786 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n250), .Z(n177) );
  MUX2_X1 U787 ( .A(n177), .B(n176), .S(n244), .Z(n178) );
  MUX2_X1 U788 ( .A(n178), .B(n175), .S(N12), .Z(n179) );
  MUX2_X1 U789 ( .A(n179), .B(n172), .S(N13), .Z(n180) );
  MUX2_X1 U790 ( .A(n180), .B(n165), .S(N14), .Z(N17) );
  MUX2_X1 U791 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n245), .Z(n181) );
  MUX2_X1 U792 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n247), .Z(n182) );
  MUX2_X1 U793 ( .A(n182), .B(n181), .S(N11), .Z(n183) );
  MUX2_X1 U794 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n246), .Z(n184) );
  MUX2_X1 U795 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n249), .Z(n185) );
  MUX2_X1 U796 ( .A(n185), .B(n184), .S(N11), .Z(n186) );
  MUX2_X1 U797 ( .A(n186), .B(n183), .S(n241), .Z(n187) );
  MUX2_X1 U798 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n249), .Z(n188) );
  MUX2_X1 U799 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(n247), .Z(n189) );
  MUX2_X1 U800 ( .A(n189), .B(n188), .S(N11), .Z(n190) );
  MUX2_X1 U801 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(n248), .Z(n191) );
  MUX2_X1 U802 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n250), .Z(n192) );
  MUX2_X1 U803 ( .A(n192), .B(n191), .S(n242), .Z(n193) );
  MUX2_X1 U804 ( .A(n193), .B(n190), .S(N12), .Z(n194) );
  MUX2_X1 U805 ( .A(n194), .B(n187), .S(N13), .Z(n195) );
  MUX2_X1 U806 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n245), .Z(n196) );
  MUX2_X1 U807 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(n250), .Z(n197) );
  MUX2_X1 U808 ( .A(n197), .B(n196), .S(n243), .Z(n198) );
  MUX2_X1 U809 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(n250), .Z(n199) );
  MUX2_X1 U810 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n248), .Z(n200) );
  MUX2_X1 U811 ( .A(n200), .B(n199), .S(n243), .Z(n201) );
  MUX2_X1 U812 ( .A(n201), .B(n198), .S(n241), .Z(n202) );
  MUX2_X1 U813 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n247), .Z(n203) );
  MUX2_X1 U814 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n250), .Z(n204) );
  MUX2_X1 U815 ( .A(n204), .B(n203), .S(n243), .Z(n205) );
  MUX2_X1 U816 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n250), .Z(n206) );
  MUX2_X1 U817 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n246), .Z(n207) );
  MUX2_X1 U818 ( .A(n207), .B(n206), .S(N11), .Z(n208) );
  MUX2_X1 U819 ( .A(n208), .B(n205), .S(N12), .Z(n209) );
  MUX2_X1 U820 ( .A(n209), .B(n202), .S(N13), .Z(n210) );
  MUX2_X1 U821 ( .A(n210), .B(n195), .S(N14), .Z(N16) );
  MUX2_X1 U822 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n250), .Z(n211) );
  MUX2_X1 U823 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n245), .Z(n212) );
  MUX2_X1 U824 ( .A(n212), .B(n211), .S(n242), .Z(n213) );
  MUX2_X1 U825 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n250), .Z(n214) );
  MUX2_X1 U826 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n249), .Z(n215) );
  MUX2_X1 U827 ( .A(n215), .B(n214), .S(n242), .Z(n216) );
  MUX2_X1 U828 ( .A(n216), .B(n213), .S(n241), .Z(n217) );
  MUX2_X1 U829 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n248), .Z(n218) );
  MUX2_X1 U830 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n250), .Z(n219) );
  MUX2_X1 U831 ( .A(n219), .B(n218), .S(N11), .Z(n220) );
  MUX2_X1 U832 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n248), .Z(n221) );
  MUX2_X1 U833 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n250), .Z(n222) );
  MUX2_X1 U834 ( .A(n222), .B(n221), .S(N11), .Z(n223) );
  MUX2_X1 U835 ( .A(n223), .B(n220), .S(N12), .Z(n224) );
  MUX2_X1 U836 ( .A(n224), .B(n217), .S(N13), .Z(n225) );
  MUX2_X1 U837 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n249), .Z(n226) );
  MUX2_X1 U838 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n249), .Z(n227) );
  MUX2_X1 U839 ( .A(n227), .B(n226), .S(n244), .Z(n228) );
  MUX2_X1 U840 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n247), .Z(n229) );
  MUX2_X1 U841 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n250), .Z(n230) );
  MUX2_X1 U842 ( .A(n230), .B(n229), .S(N11), .Z(n231) );
  MUX2_X1 U843 ( .A(n231), .B(n228), .S(n241), .Z(n232) );
  MUX2_X1 U844 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n246), .Z(n233) );
  MUX2_X1 U845 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n245), .Z(n234) );
  MUX2_X1 U846 ( .A(n234), .B(n233), .S(n244), .Z(n235) );
  MUX2_X1 U847 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n247), .Z(n236) );
  MUX2_X1 U848 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n248), .Z(n237) );
  MUX2_X1 U849 ( .A(n237), .B(n236), .S(N11), .Z(n238) );
  MUX2_X1 U850 ( .A(n238), .B(n235), .S(N12), .Z(n239) );
  MUX2_X1 U851 ( .A(n239), .B(n232), .S(N13), .Z(n240) );
  MUX2_X1 U852 ( .A(n240), .B(n225), .S(N14), .Z(N15) );
  CLKBUF_X1 U853 ( .A(n250), .Z(n245) );
endmodule


module memory_WIDTH16_SIZE32_LOGSIZE5 ( clk, data_in, data_out, addr, wr_en );
  input [15:0] data_in;
  output [15:0] data_out;
  input [4:0] addr;
  input clk, wr_en;
  wire   N10, N11, N12, N13, N14, \mem[31][15] , \mem[31][14] , \mem[31][13] ,
         \mem[31][12] , \mem[31][11] , \mem[31][10] , \mem[31][9] ,
         \mem[31][8] , \mem[31][7] , \mem[31][6] , \mem[31][5] , \mem[31][4] ,
         \mem[31][3] , \mem[31][2] , \mem[31][1] , \mem[31][0] , \mem[30][15] ,
         \mem[30][14] , \mem[30][13] , \mem[30][12] , \mem[30][11] ,
         \mem[30][10] , \mem[30][9] , \mem[30][8] , \mem[30][7] , \mem[30][6] ,
         \mem[30][5] , \mem[30][4] , \mem[30][3] , \mem[30][2] , \mem[30][1] ,
         \mem[30][0] , \mem[29][15] , \mem[29][14] , \mem[29][13] ,
         \mem[29][12] , \mem[29][11] , \mem[29][10] , \mem[29][9] ,
         \mem[29][8] , \mem[29][7] , \mem[29][6] , \mem[29][5] , \mem[29][4] ,
         \mem[29][3] , \mem[29][2] , \mem[29][1] , \mem[29][0] , \mem[28][15] ,
         \mem[28][14] , \mem[28][13] , \mem[28][12] , \mem[28][11] ,
         \mem[28][10] , \mem[28][9] , \mem[28][8] , \mem[28][7] , \mem[28][6] ,
         \mem[28][5] , \mem[28][4] , \mem[28][3] , \mem[28][2] , \mem[28][1] ,
         \mem[28][0] , \mem[27][15] , \mem[27][14] , \mem[27][13] ,
         \mem[27][12] , \mem[27][11] , \mem[27][10] , \mem[27][9] ,
         \mem[27][8] , \mem[27][7] , \mem[27][6] , \mem[27][5] , \mem[27][4] ,
         \mem[27][3] , \mem[27][2] , \mem[27][1] , \mem[27][0] , \mem[26][15] ,
         \mem[26][14] , \mem[26][13] , \mem[26][12] , \mem[26][11] ,
         \mem[26][10] , \mem[26][9] , \mem[26][8] , \mem[26][7] , \mem[26][6] ,
         \mem[26][5] , \mem[26][4] , \mem[26][3] , \mem[26][2] , \mem[26][1] ,
         \mem[26][0] , \mem[25][15] , \mem[25][14] , \mem[25][13] ,
         \mem[25][12] , \mem[25][11] , \mem[25][10] , \mem[25][9] ,
         \mem[25][8] , \mem[25][7] , \mem[25][6] , \mem[25][5] , \mem[25][4] ,
         \mem[25][3] , \mem[25][2] , \mem[25][1] , \mem[25][0] , \mem[24][15] ,
         \mem[24][14] , \mem[24][13] , \mem[24][12] , \mem[24][11] ,
         \mem[24][10] , \mem[24][9] , \mem[24][8] , \mem[24][7] , \mem[24][6] ,
         \mem[24][5] , \mem[24][4] , \mem[24][3] , \mem[24][2] , \mem[24][1] ,
         \mem[24][0] , \mem[23][15] , \mem[23][14] , \mem[23][13] ,
         \mem[23][12] , \mem[23][11] , \mem[23][10] , \mem[23][9] ,
         \mem[23][8] , \mem[23][7] , \mem[23][6] , \mem[23][5] , \mem[23][4] ,
         \mem[23][3] , \mem[23][2] , \mem[23][1] , \mem[23][0] , \mem[22][15] ,
         \mem[22][14] , \mem[22][13] , \mem[22][12] , \mem[22][11] ,
         \mem[22][10] , \mem[22][9] , \mem[22][8] , \mem[22][7] , \mem[22][6] ,
         \mem[22][5] , \mem[22][4] , \mem[22][3] , \mem[22][2] , \mem[22][1] ,
         \mem[22][0] , \mem[21][15] , \mem[21][14] , \mem[21][13] ,
         \mem[21][12] , \mem[21][11] , \mem[21][10] , \mem[21][9] ,
         \mem[21][8] , \mem[21][7] , \mem[21][6] , \mem[21][5] , \mem[21][4] ,
         \mem[21][3] , \mem[21][2] , \mem[21][1] , \mem[21][0] , \mem[20][15] ,
         \mem[20][14] , \mem[20][13] , \mem[20][12] , \mem[20][11] ,
         \mem[20][10] , \mem[20][9] , \mem[20][8] , \mem[20][7] , \mem[20][6] ,
         \mem[20][5] , \mem[20][4] , \mem[20][3] , \mem[20][2] , \mem[20][1] ,
         \mem[20][0] , \mem[19][15] , \mem[19][14] , \mem[19][13] ,
         \mem[19][12] , \mem[19][11] , \mem[19][10] , \mem[19][9] ,
         \mem[19][8] , \mem[19][7] , \mem[19][6] , \mem[19][5] , \mem[19][4] ,
         \mem[19][3] , \mem[19][2] , \mem[19][1] , \mem[19][0] , \mem[18][15] ,
         \mem[18][14] , \mem[18][13] , \mem[18][12] , \mem[18][11] ,
         \mem[18][10] , \mem[18][9] , \mem[18][8] , \mem[18][7] , \mem[18][6] ,
         \mem[18][5] , \mem[18][4] , \mem[18][3] , \mem[18][2] , \mem[18][1] ,
         \mem[18][0] , \mem[17][15] , \mem[17][14] , \mem[17][13] ,
         \mem[17][12] , \mem[17][11] , \mem[17][10] , \mem[17][9] ,
         \mem[17][8] , \mem[17][7] , \mem[17][6] , \mem[17][5] , \mem[17][4] ,
         \mem[17][3] , \mem[17][2] , \mem[17][1] , \mem[17][0] , \mem[16][15] ,
         \mem[16][14] , \mem[16][13] , \mem[16][12] , \mem[16][11] ,
         \mem[16][10] , \mem[16][9] , \mem[16][8] , \mem[16][7] , \mem[16][6] ,
         \mem[16][5] , \mem[16][4] , \mem[16][3] , \mem[16][2] , \mem[16][1] ,
         \mem[16][0] , \mem[15][15] , \mem[15][14] , \mem[15][13] ,
         \mem[15][12] , \mem[15][11] , \mem[15][10] , \mem[15][9] ,
         \mem[15][8] , \mem[15][7] , \mem[15][6] , \mem[15][5] , \mem[15][4] ,
         \mem[15][3] , \mem[15][2] , \mem[15][1] , \mem[15][0] , \mem[14][15] ,
         \mem[14][14] , \mem[14][13] , \mem[14][12] , \mem[14][11] ,
         \mem[14][10] , \mem[14][9] , \mem[14][8] , \mem[14][7] , \mem[14][6] ,
         \mem[14][5] , \mem[14][4] , \mem[14][3] , \mem[14][2] , \mem[14][1] ,
         \mem[14][0] , \mem[13][15] , \mem[13][14] , \mem[13][13] ,
         \mem[13][12] , \mem[13][11] , \mem[13][10] , \mem[13][9] ,
         \mem[13][8] , \mem[13][7] , \mem[13][6] , \mem[13][5] , \mem[13][4] ,
         \mem[13][3] , \mem[13][2] , \mem[13][1] , \mem[13][0] , \mem[12][15] ,
         \mem[12][14] , \mem[12][13] , \mem[12][12] , \mem[12][11] ,
         \mem[12][10] , \mem[12][9] , \mem[12][8] , \mem[12][7] , \mem[12][6] ,
         \mem[12][5] , \mem[12][4] , \mem[12][3] , \mem[12][2] , \mem[12][1] ,
         \mem[12][0] , \mem[11][15] , \mem[11][14] , \mem[11][13] ,
         \mem[11][12] , \mem[11][11] , \mem[11][10] , \mem[11][9] ,
         \mem[11][8] , \mem[11][7] , \mem[11][6] , \mem[11][5] , \mem[11][4] ,
         \mem[11][3] , \mem[11][2] , \mem[11][1] , \mem[11][0] , \mem[10][15] ,
         \mem[10][14] , \mem[10][13] , \mem[10][12] , \mem[10][11] ,
         \mem[10][10] , \mem[10][9] , \mem[10][8] , \mem[10][7] , \mem[10][6] ,
         \mem[10][5] , \mem[10][4] , \mem[10][3] , \mem[10][2] , \mem[10][1] ,
         \mem[10][0] , \mem[9][15] , \mem[9][14] , \mem[9][13] , \mem[9][12] ,
         \mem[9][11] , \mem[9][10] , \mem[9][9] , \mem[9][8] , \mem[9][7] ,
         \mem[9][6] , \mem[9][5] , \mem[9][4] , \mem[9][3] , \mem[9][2] ,
         \mem[9][1] , \mem[9][0] , \mem[8][15] , \mem[8][14] , \mem[8][13] ,
         \mem[8][12] , \mem[8][11] , \mem[8][10] , \mem[8][9] , \mem[8][8] ,
         \mem[8][7] , \mem[8][6] , \mem[8][5] , \mem[8][4] , \mem[8][3] ,
         \mem[8][2] , \mem[8][1] , \mem[8][0] , \mem[7][15] , \mem[7][14] ,
         \mem[7][13] , \mem[7][12] , \mem[7][11] , \mem[7][10] , \mem[7][9] ,
         \mem[7][8] , \mem[7][7] , \mem[7][6] , \mem[7][5] , \mem[7][4] ,
         \mem[7][3] , \mem[7][2] , \mem[7][1] , \mem[7][0] , \mem[6][15] ,
         \mem[6][14] , \mem[6][13] , \mem[6][12] , \mem[6][11] , \mem[6][10] ,
         \mem[6][9] , \mem[6][8] , \mem[6][7] , \mem[6][6] , \mem[6][5] ,
         \mem[6][4] , \mem[6][3] , \mem[6][2] , \mem[6][1] , \mem[6][0] ,
         \mem[5][15] , \mem[5][14] , \mem[5][13] , \mem[5][12] , \mem[5][11] ,
         \mem[5][10] , \mem[5][9] , \mem[5][8] , \mem[5][7] , \mem[5][6] ,
         \mem[5][5] , \mem[5][4] , \mem[5][3] , \mem[5][2] , \mem[5][1] ,
         \mem[5][0] , \mem[4][15] , \mem[4][14] , \mem[4][13] , \mem[4][12] ,
         \mem[4][11] , \mem[4][10] , \mem[4][9] , \mem[4][8] , \mem[4][7] ,
         \mem[4][6] , \mem[4][5] , \mem[4][4] , \mem[4][3] , \mem[4][2] ,
         \mem[4][1] , \mem[4][0] , \mem[3][15] , \mem[3][14] , \mem[3][13] ,
         \mem[3][12] , \mem[3][11] , \mem[3][10] , \mem[3][9] , \mem[3][8] ,
         \mem[3][7] , \mem[3][6] , \mem[3][5] , \mem[3][4] , \mem[3][3] ,
         \mem[3][2] , \mem[3][1] , \mem[3][0] , \mem[2][15] , \mem[2][14] ,
         \mem[2][13] , \mem[2][12] , \mem[2][11] , \mem[2][10] , \mem[2][9] ,
         \mem[2][8] , \mem[2][7] , \mem[2][6] , \mem[2][5] , \mem[2][4] ,
         \mem[2][3] , \mem[2][2] , \mem[2][1] , \mem[2][0] , \mem[1][15] ,
         \mem[1][14] , \mem[1][13] , \mem[1][12] , \mem[1][11] , \mem[1][10] ,
         \mem[1][9] , \mem[1][8] , \mem[1][7] , \mem[1][6] , \mem[1][5] ,
         \mem[1][4] , \mem[1][3] , \mem[1][2] , \mem[1][1] , \mem[1][0] ,
         \mem[0][15] , \mem[0][14] , \mem[0][13] , \mem[0][12] , \mem[0][11] ,
         \mem[0][10] , \mem[0][9] , \mem[0][8] , \mem[0][7] , \mem[0][6] ,
         \mem[0][5] , \mem[0][4] , \mem[0][3] , \mem[0][2] , \mem[0][1] ,
         \mem[0][0] , N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25,
         N26, N27, N28, N29, N30, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637;
  assign N10 = addr[0];
  assign N11 = addr[1];
  assign N12 = addr[2];
  assign N13 = addr[3];
  assign N14 = addr[4];

  DFF_X1 \data_out_reg[15]  ( .D(N15), .CK(clk), .Q(data_out[15]) );
  DFF_X1 \data_out_reg[14]  ( .D(N16), .CK(clk), .Q(data_out[14]) );
  DFF_X1 \data_out_reg[13]  ( .D(N17), .CK(clk), .Q(data_out[13]) );
  DFF_X1 \data_out_reg[12]  ( .D(N18), .CK(clk), .Q(data_out[12]) );
  DFF_X1 \data_out_reg[11]  ( .D(N19), .CK(clk), .Q(data_out[11]) );
  DFF_X1 \data_out_reg[10]  ( .D(N20), .CK(clk), .Q(data_out[10]) );
  DFF_X1 \data_out_reg[9]  ( .D(N21), .CK(clk), .Q(data_out[9]) );
  DFF_X1 \data_out_reg[8]  ( .D(N22), .CK(clk), .Q(data_out[8]) );
  DFF_X1 \data_out_reg[7]  ( .D(N23), .CK(clk), .Q(data_out[7]) );
  DFF_X1 \data_out_reg[6]  ( .D(N24), .CK(clk), .Q(data_out[6]) );
  DFF_X1 \data_out_reg[5]  ( .D(N25), .CK(clk), .Q(data_out[5]) );
  DFF_X1 \data_out_reg[4]  ( .D(N26), .CK(clk), .Q(data_out[4]) );
  DFF_X1 \data_out_reg[3]  ( .D(N27), .CK(clk), .Q(data_out[3]) );
  DFF_X1 \data_out_reg[2]  ( .D(N28), .CK(clk), .Q(data_out[2]) );
  DFF_X1 \data_out_reg[1]  ( .D(N29), .CK(clk), .Q(data_out[1]) );
  DFF_X1 \data_out_reg[0]  ( .D(N30), .CK(clk), .Q(data_out[0]) );
  DFF_X1 \mem_reg[31][15]  ( .D(n1605), .CK(clk), .Q(\mem[31][15] ) );
  DFF_X1 \mem_reg[31][14]  ( .D(n1606), .CK(clk), .Q(\mem[31][14] ) );
  DFF_X1 \mem_reg[31][13]  ( .D(n1607), .CK(clk), .Q(\mem[31][13] ) );
  DFF_X1 \mem_reg[31][12]  ( .D(n1608), .CK(clk), .Q(\mem[31][12] ) );
  DFF_X1 \mem_reg[31][11]  ( .D(n1609), .CK(clk), .Q(\mem[31][11] ) );
  DFF_X1 \mem_reg[31][10]  ( .D(n1610), .CK(clk), .Q(\mem[31][10] ) );
  DFF_X1 \mem_reg[31][9]  ( .D(n1611), .CK(clk), .Q(\mem[31][9] ) );
  DFF_X1 \mem_reg[31][8]  ( .D(n1612), .CK(clk), .Q(\mem[31][8] ) );
  DFF_X1 \mem_reg[31][7]  ( .D(n1613), .CK(clk), .Q(\mem[31][7] ) );
  DFF_X1 \mem_reg[31][6]  ( .D(n1614), .CK(clk), .Q(\mem[31][6] ) );
  DFF_X1 \mem_reg[31][5]  ( .D(n1615), .CK(clk), .Q(\mem[31][5] ) );
  DFF_X1 \mem_reg[31][4]  ( .D(n1616), .CK(clk), .Q(\mem[31][4] ) );
  DFF_X1 \mem_reg[31][3]  ( .D(n1617), .CK(clk), .Q(\mem[31][3] ) );
  DFF_X1 \mem_reg[31][2]  ( .D(n1618), .CK(clk), .Q(\mem[31][2] ) );
  DFF_X1 \mem_reg[31][1]  ( .D(n1619), .CK(clk), .Q(\mem[31][1] ) );
  DFF_X1 \mem_reg[31][0]  ( .D(n1620), .CK(clk), .Q(\mem[31][0] ) );
  DFF_X1 \mem_reg[30][15]  ( .D(n1089), .CK(clk), .Q(\mem[30][15] ) );
  DFF_X1 \mem_reg[30][14]  ( .D(n1088), .CK(clk), .Q(\mem[30][14] ) );
  DFF_X1 \mem_reg[30][13]  ( .D(n1087), .CK(clk), .Q(\mem[30][13] ) );
  DFF_X1 \mem_reg[30][12]  ( .D(n1086), .CK(clk), .Q(\mem[30][12] ) );
  DFF_X1 \mem_reg[30][11]  ( .D(n1085), .CK(clk), .Q(\mem[30][11] ) );
  DFF_X1 \mem_reg[30][10]  ( .D(n1084), .CK(clk), .Q(\mem[30][10] ) );
  DFF_X1 \mem_reg[30][9]  ( .D(n1083), .CK(clk), .Q(\mem[30][9] ) );
  DFF_X1 \mem_reg[30][8]  ( .D(n1082), .CK(clk), .Q(\mem[30][8] ) );
  DFF_X1 \mem_reg[30][7]  ( .D(n1081), .CK(clk), .Q(\mem[30][7] ) );
  DFF_X1 \mem_reg[30][6]  ( .D(n1080), .CK(clk), .Q(\mem[30][6] ) );
  DFF_X1 \mem_reg[30][5]  ( .D(n1079), .CK(clk), .Q(\mem[30][5] ) );
  DFF_X1 \mem_reg[30][4]  ( .D(n1078), .CK(clk), .Q(\mem[30][4] ) );
  DFF_X1 \mem_reg[30][3]  ( .D(n1077), .CK(clk), .Q(\mem[30][3] ) );
  DFF_X1 \mem_reg[30][2]  ( .D(n1076), .CK(clk), .Q(\mem[30][2] ) );
  DFF_X1 \mem_reg[30][1]  ( .D(n1075), .CK(clk), .Q(\mem[30][1] ) );
  DFF_X1 \mem_reg[30][0]  ( .D(n1074), .CK(clk), .Q(\mem[30][0] ) );
  DFF_X1 \mem_reg[29][15]  ( .D(n1073), .CK(clk), .Q(\mem[29][15] ) );
  DFF_X1 \mem_reg[29][14]  ( .D(n1072), .CK(clk), .Q(\mem[29][14] ) );
  DFF_X1 \mem_reg[29][13]  ( .D(n1071), .CK(clk), .Q(\mem[29][13] ) );
  DFF_X1 \mem_reg[29][12]  ( .D(n1070), .CK(clk), .Q(\mem[29][12] ) );
  DFF_X1 \mem_reg[29][11]  ( .D(n1069), .CK(clk), .Q(\mem[29][11] ) );
  DFF_X1 \mem_reg[29][10]  ( .D(n1068), .CK(clk), .Q(\mem[29][10] ) );
  DFF_X1 \mem_reg[29][9]  ( .D(n1067), .CK(clk), .Q(\mem[29][9] ) );
  DFF_X1 \mem_reg[29][8]  ( .D(n1066), .CK(clk), .Q(\mem[29][8] ) );
  DFF_X1 \mem_reg[29][7]  ( .D(n1065), .CK(clk), .Q(\mem[29][7] ) );
  DFF_X1 \mem_reg[29][6]  ( .D(n1064), .CK(clk), .Q(\mem[29][6] ) );
  DFF_X1 \mem_reg[29][5]  ( .D(n1063), .CK(clk), .Q(\mem[29][5] ) );
  DFF_X1 \mem_reg[29][4]  ( .D(n1062), .CK(clk), .Q(\mem[29][4] ) );
  DFF_X1 \mem_reg[29][3]  ( .D(n1061), .CK(clk), .Q(\mem[29][3] ) );
  DFF_X1 \mem_reg[29][2]  ( .D(n1060), .CK(clk), .Q(\mem[29][2] ) );
  DFF_X1 \mem_reg[29][1]  ( .D(n1059), .CK(clk), .Q(\mem[29][1] ) );
  DFF_X1 \mem_reg[29][0]  ( .D(n1058), .CK(clk), .Q(\mem[29][0] ) );
  DFF_X1 \mem_reg[28][15]  ( .D(n1057), .CK(clk), .Q(\mem[28][15] ) );
  DFF_X1 \mem_reg[28][14]  ( .D(n1056), .CK(clk), .Q(\mem[28][14] ) );
  DFF_X1 \mem_reg[28][13]  ( .D(n1055), .CK(clk), .Q(\mem[28][13] ) );
  DFF_X1 \mem_reg[28][12]  ( .D(n1054), .CK(clk), .Q(\mem[28][12] ) );
  DFF_X1 \mem_reg[28][11]  ( .D(n1053), .CK(clk), .Q(\mem[28][11] ) );
  DFF_X1 \mem_reg[28][10]  ( .D(n1052), .CK(clk), .Q(\mem[28][10] ) );
  DFF_X1 \mem_reg[28][9]  ( .D(n1051), .CK(clk), .Q(\mem[28][9] ) );
  DFF_X1 \mem_reg[28][8]  ( .D(n1050), .CK(clk), .Q(\mem[28][8] ) );
  DFF_X1 \mem_reg[28][7]  ( .D(n1049), .CK(clk), .Q(\mem[28][7] ) );
  DFF_X1 \mem_reg[28][6]  ( .D(n1048), .CK(clk), .Q(\mem[28][6] ) );
  DFF_X1 \mem_reg[28][5]  ( .D(n1047), .CK(clk), .Q(\mem[28][5] ) );
  DFF_X1 \mem_reg[28][4]  ( .D(n1046), .CK(clk), .Q(\mem[28][4] ) );
  DFF_X1 \mem_reg[28][3]  ( .D(n1045), .CK(clk), .Q(\mem[28][3] ) );
  DFF_X1 \mem_reg[28][2]  ( .D(n1044), .CK(clk), .Q(\mem[28][2] ) );
  DFF_X1 \mem_reg[28][1]  ( .D(n1043), .CK(clk), .Q(\mem[28][1] ) );
  DFF_X1 \mem_reg[28][0]  ( .D(n1042), .CK(clk), .Q(\mem[28][0] ) );
  DFF_X1 \mem_reg[27][15]  ( .D(n1041), .CK(clk), .Q(\mem[27][15] ) );
  DFF_X1 \mem_reg[27][14]  ( .D(n1040), .CK(clk), .Q(\mem[27][14] ) );
  DFF_X1 \mem_reg[27][13]  ( .D(n1039), .CK(clk), .Q(\mem[27][13] ) );
  DFF_X1 \mem_reg[27][12]  ( .D(n1038), .CK(clk), .Q(\mem[27][12] ) );
  DFF_X1 \mem_reg[27][11]  ( .D(n1037), .CK(clk), .Q(\mem[27][11] ) );
  DFF_X1 \mem_reg[27][10]  ( .D(n1036), .CK(clk), .Q(\mem[27][10] ) );
  DFF_X1 \mem_reg[27][9]  ( .D(n1035), .CK(clk), .Q(\mem[27][9] ) );
  DFF_X1 \mem_reg[27][8]  ( .D(n1034), .CK(clk), .Q(\mem[27][8] ) );
  DFF_X1 \mem_reg[27][7]  ( .D(n1033), .CK(clk), .Q(\mem[27][7] ) );
  DFF_X1 \mem_reg[27][6]  ( .D(n1032), .CK(clk), .Q(\mem[27][6] ) );
  DFF_X1 \mem_reg[27][5]  ( .D(n1031), .CK(clk), .Q(\mem[27][5] ) );
  DFF_X1 \mem_reg[27][4]  ( .D(n1030), .CK(clk), .Q(\mem[27][4] ) );
  DFF_X1 \mem_reg[27][3]  ( .D(n1029), .CK(clk), .Q(\mem[27][3] ) );
  DFF_X1 \mem_reg[27][2]  ( .D(n1028), .CK(clk), .Q(\mem[27][2] ) );
  DFF_X1 \mem_reg[27][1]  ( .D(n1027), .CK(clk), .Q(\mem[27][1] ) );
  DFF_X1 \mem_reg[27][0]  ( .D(n1026), .CK(clk), .Q(\mem[27][0] ) );
  DFF_X1 \mem_reg[26][15]  ( .D(n1025), .CK(clk), .Q(\mem[26][15] ) );
  DFF_X1 \mem_reg[26][14]  ( .D(n1024), .CK(clk), .Q(\mem[26][14] ) );
  DFF_X1 \mem_reg[26][13]  ( .D(n1023), .CK(clk), .Q(\mem[26][13] ) );
  DFF_X1 \mem_reg[26][12]  ( .D(n1022), .CK(clk), .Q(\mem[26][12] ) );
  DFF_X1 \mem_reg[26][11]  ( .D(n1021), .CK(clk), .Q(\mem[26][11] ) );
  DFF_X1 \mem_reg[26][10]  ( .D(n1020), .CK(clk), .Q(\mem[26][10] ) );
  DFF_X1 \mem_reg[26][9]  ( .D(n1019), .CK(clk), .Q(\mem[26][9] ) );
  DFF_X1 \mem_reg[26][8]  ( .D(n1018), .CK(clk), .Q(\mem[26][8] ) );
  DFF_X1 \mem_reg[26][7]  ( .D(n1017), .CK(clk), .Q(\mem[26][7] ) );
  DFF_X1 \mem_reg[26][6]  ( .D(n1016), .CK(clk), .Q(\mem[26][6] ) );
  DFF_X1 \mem_reg[26][5]  ( .D(n1015), .CK(clk), .Q(\mem[26][5] ) );
  DFF_X1 \mem_reg[26][4]  ( .D(n1014), .CK(clk), .Q(\mem[26][4] ) );
  DFF_X1 \mem_reg[26][3]  ( .D(n1013), .CK(clk), .Q(\mem[26][3] ) );
  DFF_X1 \mem_reg[26][2]  ( .D(n1012), .CK(clk), .Q(\mem[26][2] ) );
  DFF_X1 \mem_reg[26][1]  ( .D(n1011), .CK(clk), .Q(\mem[26][1] ) );
  DFF_X1 \mem_reg[26][0]  ( .D(n1010), .CK(clk), .Q(\mem[26][0] ) );
  DFF_X1 \mem_reg[25][15]  ( .D(n1009), .CK(clk), .Q(\mem[25][15] ) );
  DFF_X1 \mem_reg[25][14]  ( .D(n1008), .CK(clk), .Q(\mem[25][14] ) );
  DFF_X1 \mem_reg[25][13]  ( .D(n1007), .CK(clk), .Q(\mem[25][13] ) );
  DFF_X1 \mem_reg[25][12]  ( .D(n1006), .CK(clk), .Q(\mem[25][12] ) );
  DFF_X1 \mem_reg[25][11]  ( .D(n1005), .CK(clk), .Q(\mem[25][11] ) );
  DFF_X1 \mem_reg[25][10]  ( .D(n1004), .CK(clk), .Q(\mem[25][10] ) );
  DFF_X1 \mem_reg[25][9]  ( .D(n1003), .CK(clk), .Q(\mem[25][9] ) );
  DFF_X1 \mem_reg[25][8]  ( .D(n1002), .CK(clk), .Q(\mem[25][8] ) );
  DFF_X1 \mem_reg[25][7]  ( .D(n1001), .CK(clk), .Q(\mem[25][7] ) );
  DFF_X1 \mem_reg[25][6]  ( .D(n1000), .CK(clk), .Q(\mem[25][6] ) );
  DFF_X1 \mem_reg[25][5]  ( .D(n999), .CK(clk), .Q(\mem[25][5] ) );
  DFF_X1 \mem_reg[25][4]  ( .D(n998), .CK(clk), .Q(\mem[25][4] ) );
  DFF_X1 \mem_reg[25][3]  ( .D(n997), .CK(clk), .Q(\mem[25][3] ) );
  DFF_X1 \mem_reg[25][2]  ( .D(n996), .CK(clk), .Q(\mem[25][2] ) );
  DFF_X1 \mem_reg[25][1]  ( .D(n995), .CK(clk), .Q(\mem[25][1] ) );
  DFF_X1 \mem_reg[25][0]  ( .D(n994), .CK(clk), .Q(\mem[25][0] ) );
  DFF_X1 \mem_reg[24][15]  ( .D(n993), .CK(clk), .Q(\mem[24][15] ) );
  DFF_X1 \mem_reg[24][14]  ( .D(n992), .CK(clk), .Q(\mem[24][14] ) );
  DFF_X1 \mem_reg[24][13]  ( .D(n991), .CK(clk), .Q(\mem[24][13] ) );
  DFF_X1 \mem_reg[24][12]  ( .D(n990), .CK(clk), .Q(\mem[24][12] ) );
  DFF_X1 \mem_reg[24][11]  ( .D(n989), .CK(clk), .Q(\mem[24][11] ) );
  DFF_X1 \mem_reg[24][10]  ( .D(n988), .CK(clk), .Q(\mem[24][10] ) );
  DFF_X1 \mem_reg[24][9]  ( .D(n987), .CK(clk), .Q(\mem[24][9] ) );
  DFF_X1 \mem_reg[24][8]  ( .D(n986), .CK(clk), .Q(\mem[24][8] ) );
  DFF_X1 \mem_reg[24][7]  ( .D(n985), .CK(clk), .Q(\mem[24][7] ) );
  DFF_X1 \mem_reg[24][6]  ( .D(n984), .CK(clk), .Q(\mem[24][6] ) );
  DFF_X1 \mem_reg[24][5]  ( .D(n983), .CK(clk), .Q(\mem[24][5] ) );
  DFF_X1 \mem_reg[24][4]  ( .D(n982), .CK(clk), .Q(\mem[24][4] ) );
  DFF_X1 \mem_reg[24][3]  ( .D(n981), .CK(clk), .Q(\mem[24][3] ) );
  DFF_X1 \mem_reg[24][2]  ( .D(n980), .CK(clk), .Q(\mem[24][2] ) );
  DFF_X1 \mem_reg[24][1]  ( .D(n979), .CK(clk), .Q(\mem[24][1] ) );
  DFF_X1 \mem_reg[24][0]  ( .D(n978), .CK(clk), .Q(\mem[24][0] ) );
  DFF_X1 \mem_reg[23][15]  ( .D(n977), .CK(clk), .Q(\mem[23][15] ) );
  DFF_X1 \mem_reg[23][14]  ( .D(n976), .CK(clk), .Q(\mem[23][14] ) );
  DFF_X1 \mem_reg[23][13]  ( .D(n975), .CK(clk), .Q(\mem[23][13] ) );
  DFF_X1 \mem_reg[23][12]  ( .D(n974), .CK(clk), .Q(\mem[23][12] ) );
  DFF_X1 \mem_reg[23][11]  ( .D(n973), .CK(clk), .Q(\mem[23][11] ) );
  DFF_X1 \mem_reg[23][10]  ( .D(n972), .CK(clk), .Q(\mem[23][10] ) );
  DFF_X1 \mem_reg[23][9]  ( .D(n971), .CK(clk), .Q(\mem[23][9] ) );
  DFF_X1 \mem_reg[23][8]  ( .D(n970), .CK(clk), .Q(\mem[23][8] ) );
  DFF_X1 \mem_reg[23][7]  ( .D(n969), .CK(clk), .Q(\mem[23][7] ) );
  DFF_X1 \mem_reg[23][6]  ( .D(n968), .CK(clk), .Q(\mem[23][6] ) );
  DFF_X1 \mem_reg[23][5]  ( .D(n967), .CK(clk), .Q(\mem[23][5] ) );
  DFF_X1 \mem_reg[23][4]  ( .D(n966), .CK(clk), .Q(\mem[23][4] ) );
  DFF_X1 \mem_reg[23][3]  ( .D(n965), .CK(clk), .Q(\mem[23][3] ) );
  DFF_X1 \mem_reg[23][2]  ( .D(n964), .CK(clk), .Q(\mem[23][2] ) );
  DFF_X1 \mem_reg[23][1]  ( .D(n963), .CK(clk), .Q(\mem[23][1] ) );
  DFF_X1 \mem_reg[23][0]  ( .D(n962), .CK(clk), .Q(\mem[23][0] ) );
  DFF_X1 \mem_reg[22][15]  ( .D(n961), .CK(clk), .Q(\mem[22][15] ) );
  DFF_X1 \mem_reg[22][14]  ( .D(n960), .CK(clk), .Q(\mem[22][14] ) );
  DFF_X1 \mem_reg[22][13]  ( .D(n959), .CK(clk), .Q(\mem[22][13] ) );
  DFF_X1 \mem_reg[22][12]  ( .D(n958), .CK(clk), .Q(\mem[22][12] ) );
  DFF_X1 \mem_reg[22][11]  ( .D(n957), .CK(clk), .Q(\mem[22][11] ) );
  DFF_X1 \mem_reg[22][10]  ( .D(n956), .CK(clk), .Q(\mem[22][10] ) );
  DFF_X1 \mem_reg[22][9]  ( .D(n955), .CK(clk), .Q(\mem[22][9] ) );
  DFF_X1 \mem_reg[22][8]  ( .D(n954), .CK(clk), .Q(\mem[22][8] ) );
  DFF_X1 \mem_reg[22][7]  ( .D(n953), .CK(clk), .Q(\mem[22][7] ) );
  DFF_X1 \mem_reg[22][6]  ( .D(n952), .CK(clk), .Q(\mem[22][6] ) );
  DFF_X1 \mem_reg[22][5]  ( .D(n951), .CK(clk), .Q(\mem[22][5] ) );
  DFF_X1 \mem_reg[22][4]  ( .D(n950), .CK(clk), .Q(\mem[22][4] ) );
  DFF_X1 \mem_reg[22][3]  ( .D(n949), .CK(clk), .Q(\mem[22][3] ) );
  DFF_X1 \mem_reg[22][2]  ( .D(n948), .CK(clk), .Q(\mem[22][2] ) );
  DFF_X1 \mem_reg[22][1]  ( .D(n947), .CK(clk), .Q(\mem[22][1] ) );
  DFF_X1 \mem_reg[22][0]  ( .D(n946), .CK(clk), .Q(\mem[22][0] ) );
  DFF_X1 \mem_reg[21][15]  ( .D(n945), .CK(clk), .Q(\mem[21][15] ) );
  DFF_X1 \mem_reg[21][14]  ( .D(n944), .CK(clk), .Q(\mem[21][14] ) );
  DFF_X1 \mem_reg[21][13]  ( .D(n943), .CK(clk), .Q(\mem[21][13] ) );
  DFF_X1 \mem_reg[21][12]  ( .D(n942), .CK(clk), .Q(\mem[21][12] ) );
  DFF_X1 \mem_reg[21][11]  ( .D(n941), .CK(clk), .Q(\mem[21][11] ) );
  DFF_X1 \mem_reg[21][10]  ( .D(n940), .CK(clk), .Q(\mem[21][10] ) );
  DFF_X1 \mem_reg[21][9]  ( .D(n939), .CK(clk), .Q(\mem[21][9] ) );
  DFF_X1 \mem_reg[21][8]  ( .D(n938), .CK(clk), .Q(\mem[21][8] ) );
  DFF_X1 \mem_reg[21][7]  ( .D(n937), .CK(clk), .Q(\mem[21][7] ) );
  DFF_X1 \mem_reg[21][6]  ( .D(n936), .CK(clk), .Q(\mem[21][6] ) );
  DFF_X1 \mem_reg[21][5]  ( .D(n935), .CK(clk), .Q(\mem[21][5] ) );
  DFF_X1 \mem_reg[21][4]  ( .D(n934), .CK(clk), .Q(\mem[21][4] ) );
  DFF_X1 \mem_reg[21][3]  ( .D(n933), .CK(clk), .Q(\mem[21][3] ) );
  DFF_X1 \mem_reg[21][2]  ( .D(n932), .CK(clk), .Q(\mem[21][2] ) );
  DFF_X1 \mem_reg[21][1]  ( .D(n931), .CK(clk), .Q(\mem[21][1] ) );
  DFF_X1 \mem_reg[21][0]  ( .D(n930), .CK(clk), .Q(\mem[21][0] ) );
  DFF_X1 \mem_reg[20][15]  ( .D(n929), .CK(clk), .Q(\mem[20][15] ) );
  DFF_X1 \mem_reg[20][14]  ( .D(n928), .CK(clk), .Q(\mem[20][14] ) );
  DFF_X1 \mem_reg[20][13]  ( .D(n927), .CK(clk), .Q(\mem[20][13] ) );
  DFF_X1 \mem_reg[20][12]  ( .D(n926), .CK(clk), .Q(\mem[20][12] ) );
  DFF_X1 \mem_reg[20][11]  ( .D(n925), .CK(clk), .Q(\mem[20][11] ) );
  DFF_X1 \mem_reg[20][10]  ( .D(n924), .CK(clk), .Q(\mem[20][10] ) );
  DFF_X1 \mem_reg[20][9]  ( .D(n923), .CK(clk), .Q(\mem[20][9] ) );
  DFF_X1 \mem_reg[20][8]  ( .D(n922), .CK(clk), .Q(\mem[20][8] ) );
  DFF_X1 \mem_reg[20][7]  ( .D(n921), .CK(clk), .Q(\mem[20][7] ) );
  DFF_X1 \mem_reg[20][6]  ( .D(n920), .CK(clk), .Q(\mem[20][6] ) );
  DFF_X1 \mem_reg[20][5]  ( .D(n919), .CK(clk), .Q(\mem[20][5] ) );
  DFF_X1 \mem_reg[20][4]  ( .D(n918), .CK(clk), .Q(\mem[20][4] ) );
  DFF_X1 \mem_reg[20][3]  ( .D(n917), .CK(clk), .Q(\mem[20][3] ) );
  DFF_X1 \mem_reg[20][2]  ( .D(n916), .CK(clk), .Q(\mem[20][2] ) );
  DFF_X1 \mem_reg[20][1]  ( .D(n915), .CK(clk), .Q(\mem[20][1] ) );
  DFF_X1 \mem_reg[20][0]  ( .D(n914), .CK(clk), .Q(\mem[20][0] ) );
  DFF_X1 \mem_reg[19][15]  ( .D(n913), .CK(clk), .Q(\mem[19][15] ) );
  DFF_X1 \mem_reg[19][14]  ( .D(n912), .CK(clk), .Q(\mem[19][14] ) );
  DFF_X1 \mem_reg[19][13]  ( .D(n911), .CK(clk), .Q(\mem[19][13] ) );
  DFF_X1 \mem_reg[19][12]  ( .D(n910), .CK(clk), .Q(\mem[19][12] ) );
  DFF_X1 \mem_reg[19][11]  ( .D(n909), .CK(clk), .Q(\mem[19][11] ) );
  DFF_X1 \mem_reg[19][10]  ( .D(n908), .CK(clk), .Q(\mem[19][10] ) );
  DFF_X1 \mem_reg[19][9]  ( .D(n907), .CK(clk), .Q(\mem[19][9] ) );
  DFF_X1 \mem_reg[19][8]  ( .D(n906), .CK(clk), .Q(\mem[19][8] ) );
  DFF_X1 \mem_reg[19][7]  ( .D(n905), .CK(clk), .Q(\mem[19][7] ) );
  DFF_X1 \mem_reg[19][6]  ( .D(n904), .CK(clk), .Q(\mem[19][6] ) );
  DFF_X1 \mem_reg[19][5]  ( .D(n903), .CK(clk), .Q(\mem[19][5] ) );
  DFF_X1 \mem_reg[19][4]  ( .D(n902), .CK(clk), .Q(\mem[19][4] ) );
  DFF_X1 \mem_reg[19][3]  ( .D(n901), .CK(clk), .Q(\mem[19][3] ) );
  DFF_X1 \mem_reg[19][2]  ( .D(n900), .CK(clk), .Q(\mem[19][2] ) );
  DFF_X1 \mem_reg[19][1]  ( .D(n899), .CK(clk), .Q(\mem[19][1] ) );
  DFF_X1 \mem_reg[19][0]  ( .D(n898), .CK(clk), .Q(\mem[19][0] ) );
  DFF_X1 \mem_reg[18][15]  ( .D(n897), .CK(clk), .Q(\mem[18][15] ) );
  DFF_X1 \mem_reg[18][14]  ( .D(n896), .CK(clk), .Q(\mem[18][14] ) );
  DFF_X1 \mem_reg[18][13]  ( .D(n895), .CK(clk), .Q(\mem[18][13] ) );
  DFF_X1 \mem_reg[18][12]  ( .D(n894), .CK(clk), .Q(\mem[18][12] ) );
  DFF_X1 \mem_reg[18][11]  ( .D(n893), .CK(clk), .Q(\mem[18][11] ) );
  DFF_X1 \mem_reg[18][10]  ( .D(n892), .CK(clk), .Q(\mem[18][10] ) );
  DFF_X1 \mem_reg[18][9]  ( .D(n891), .CK(clk), .Q(\mem[18][9] ) );
  DFF_X1 \mem_reg[18][8]  ( .D(n890), .CK(clk), .Q(\mem[18][8] ) );
  DFF_X1 \mem_reg[18][7]  ( .D(n889), .CK(clk), .Q(\mem[18][7] ) );
  DFF_X1 \mem_reg[18][6]  ( .D(n888), .CK(clk), .Q(\mem[18][6] ) );
  DFF_X1 \mem_reg[18][5]  ( .D(n887), .CK(clk), .Q(\mem[18][5] ) );
  DFF_X1 \mem_reg[18][4]  ( .D(n886), .CK(clk), .Q(\mem[18][4] ) );
  DFF_X1 \mem_reg[18][3]  ( .D(n885), .CK(clk), .Q(\mem[18][3] ) );
  DFF_X1 \mem_reg[18][2]  ( .D(n884), .CK(clk), .Q(\mem[18][2] ) );
  DFF_X1 \mem_reg[18][1]  ( .D(n883), .CK(clk), .Q(\mem[18][1] ) );
  DFF_X1 \mem_reg[18][0]  ( .D(n882), .CK(clk), .Q(\mem[18][0] ) );
  DFF_X1 \mem_reg[17][15]  ( .D(n881), .CK(clk), .Q(\mem[17][15] ) );
  DFF_X1 \mem_reg[17][14]  ( .D(n880), .CK(clk), .Q(\mem[17][14] ) );
  DFF_X1 \mem_reg[17][13]  ( .D(n879), .CK(clk), .Q(\mem[17][13] ) );
  DFF_X1 \mem_reg[17][12]  ( .D(n878), .CK(clk), .Q(\mem[17][12] ) );
  DFF_X1 \mem_reg[17][11]  ( .D(n877), .CK(clk), .Q(\mem[17][11] ) );
  DFF_X1 \mem_reg[17][10]  ( .D(n876), .CK(clk), .Q(\mem[17][10] ) );
  DFF_X1 \mem_reg[17][9]  ( .D(n875), .CK(clk), .Q(\mem[17][9] ) );
  DFF_X1 \mem_reg[17][8]  ( .D(n874), .CK(clk), .Q(\mem[17][8] ) );
  DFF_X1 \mem_reg[17][7]  ( .D(n873), .CK(clk), .Q(\mem[17][7] ) );
  DFF_X1 \mem_reg[17][6]  ( .D(n872), .CK(clk), .Q(\mem[17][6] ) );
  DFF_X1 \mem_reg[17][5]  ( .D(n871), .CK(clk), .Q(\mem[17][5] ) );
  DFF_X1 \mem_reg[17][4]  ( .D(n870), .CK(clk), .Q(\mem[17][4] ) );
  DFF_X1 \mem_reg[17][3]  ( .D(n869), .CK(clk), .Q(\mem[17][3] ) );
  DFF_X1 \mem_reg[17][2]  ( .D(n868), .CK(clk), .Q(\mem[17][2] ) );
  DFF_X1 \mem_reg[17][1]  ( .D(n867), .CK(clk), .Q(\mem[17][1] ) );
  DFF_X1 \mem_reg[17][0]  ( .D(n866), .CK(clk), .Q(\mem[17][0] ) );
  DFF_X1 \mem_reg[16][15]  ( .D(n865), .CK(clk), .Q(\mem[16][15] ) );
  DFF_X1 \mem_reg[16][14]  ( .D(n864), .CK(clk), .Q(\mem[16][14] ) );
  DFF_X1 \mem_reg[16][13]  ( .D(n863), .CK(clk), .Q(\mem[16][13] ) );
  DFF_X1 \mem_reg[16][12]  ( .D(n862), .CK(clk), .Q(\mem[16][12] ) );
  DFF_X1 \mem_reg[16][11]  ( .D(n861), .CK(clk), .Q(\mem[16][11] ) );
  DFF_X1 \mem_reg[16][10]  ( .D(n860), .CK(clk), .Q(\mem[16][10] ) );
  DFF_X1 \mem_reg[16][9]  ( .D(n859), .CK(clk), .Q(\mem[16][9] ) );
  DFF_X1 \mem_reg[16][8]  ( .D(n858), .CK(clk), .Q(\mem[16][8] ) );
  DFF_X1 \mem_reg[16][7]  ( .D(n857), .CK(clk), .Q(\mem[16][7] ) );
  DFF_X1 \mem_reg[16][6]  ( .D(n856), .CK(clk), .Q(\mem[16][6] ) );
  DFF_X1 \mem_reg[16][5]  ( .D(n855), .CK(clk), .Q(\mem[16][5] ) );
  DFF_X1 \mem_reg[16][4]  ( .D(n854), .CK(clk), .Q(\mem[16][4] ) );
  DFF_X1 \mem_reg[16][3]  ( .D(n853), .CK(clk), .Q(\mem[16][3] ) );
  DFF_X1 \mem_reg[16][2]  ( .D(n852), .CK(clk), .Q(\mem[16][2] ) );
  DFF_X1 \mem_reg[16][1]  ( .D(n851), .CK(clk), .Q(\mem[16][1] ) );
  DFF_X1 \mem_reg[16][0]  ( .D(n850), .CK(clk), .Q(\mem[16][0] ) );
  DFF_X1 \mem_reg[15][15]  ( .D(n849), .CK(clk), .Q(\mem[15][15] ) );
  DFF_X1 \mem_reg[15][14]  ( .D(n848), .CK(clk), .Q(\mem[15][14] ) );
  DFF_X1 \mem_reg[15][13]  ( .D(n847), .CK(clk), .Q(\mem[15][13] ) );
  DFF_X1 \mem_reg[15][12]  ( .D(n846), .CK(clk), .Q(\mem[15][12] ) );
  DFF_X1 \mem_reg[15][11]  ( .D(n845), .CK(clk), .Q(\mem[15][11] ) );
  DFF_X1 \mem_reg[15][10]  ( .D(n844), .CK(clk), .Q(\mem[15][10] ) );
  DFF_X1 \mem_reg[15][9]  ( .D(n843), .CK(clk), .Q(\mem[15][9] ) );
  DFF_X1 \mem_reg[15][8]  ( .D(n842), .CK(clk), .Q(\mem[15][8] ) );
  DFF_X1 \mem_reg[15][7]  ( .D(n841), .CK(clk), .Q(\mem[15][7] ) );
  DFF_X1 \mem_reg[15][6]  ( .D(n840), .CK(clk), .Q(\mem[15][6] ) );
  DFF_X1 \mem_reg[15][5]  ( .D(n839), .CK(clk), .Q(\mem[15][5] ) );
  DFF_X1 \mem_reg[15][4]  ( .D(n838), .CK(clk), .Q(\mem[15][4] ) );
  DFF_X1 \mem_reg[15][3]  ( .D(n837), .CK(clk), .Q(\mem[15][3] ) );
  DFF_X1 \mem_reg[15][2]  ( .D(n836), .CK(clk), .Q(\mem[15][2] ) );
  DFF_X1 \mem_reg[15][1]  ( .D(n835), .CK(clk), .Q(\mem[15][1] ) );
  DFF_X1 \mem_reg[15][0]  ( .D(n834), .CK(clk), .Q(\mem[15][0] ) );
  DFF_X1 \mem_reg[14][15]  ( .D(n833), .CK(clk), .Q(\mem[14][15] ) );
  DFF_X1 \mem_reg[14][14]  ( .D(n832), .CK(clk), .Q(\mem[14][14] ) );
  DFF_X1 \mem_reg[14][13]  ( .D(n831), .CK(clk), .Q(\mem[14][13] ) );
  DFF_X1 \mem_reg[14][12]  ( .D(n830), .CK(clk), .Q(\mem[14][12] ) );
  DFF_X1 \mem_reg[14][11]  ( .D(n829), .CK(clk), .Q(\mem[14][11] ) );
  DFF_X1 \mem_reg[14][10]  ( .D(n828), .CK(clk), .Q(\mem[14][10] ) );
  DFF_X1 \mem_reg[14][9]  ( .D(n827), .CK(clk), .Q(\mem[14][9] ) );
  DFF_X1 \mem_reg[14][8]  ( .D(n826), .CK(clk), .Q(\mem[14][8] ) );
  DFF_X1 \mem_reg[14][7]  ( .D(n825), .CK(clk), .Q(\mem[14][7] ) );
  DFF_X1 \mem_reg[14][6]  ( .D(n824), .CK(clk), .Q(\mem[14][6] ) );
  DFF_X1 \mem_reg[14][5]  ( .D(n823), .CK(clk), .Q(\mem[14][5] ) );
  DFF_X1 \mem_reg[14][4]  ( .D(n822), .CK(clk), .Q(\mem[14][4] ) );
  DFF_X1 \mem_reg[14][3]  ( .D(n821), .CK(clk), .Q(\mem[14][3] ) );
  DFF_X1 \mem_reg[14][2]  ( .D(n820), .CK(clk), .Q(\mem[14][2] ) );
  DFF_X1 \mem_reg[14][1]  ( .D(n819), .CK(clk), .Q(\mem[14][1] ) );
  DFF_X1 \mem_reg[14][0]  ( .D(n818), .CK(clk), .Q(\mem[14][0] ) );
  DFF_X1 \mem_reg[13][15]  ( .D(n817), .CK(clk), .Q(\mem[13][15] ) );
  DFF_X1 \mem_reg[13][14]  ( .D(n816), .CK(clk), .Q(\mem[13][14] ) );
  DFF_X1 \mem_reg[13][13]  ( .D(n815), .CK(clk), .Q(\mem[13][13] ) );
  DFF_X1 \mem_reg[13][12]  ( .D(n814), .CK(clk), .Q(\mem[13][12] ) );
  DFF_X1 \mem_reg[13][11]  ( .D(n813), .CK(clk), .Q(\mem[13][11] ) );
  DFF_X1 \mem_reg[13][10]  ( .D(n812), .CK(clk), .Q(\mem[13][10] ) );
  DFF_X1 \mem_reg[13][9]  ( .D(n811), .CK(clk), .Q(\mem[13][9] ) );
  DFF_X1 \mem_reg[13][8]  ( .D(n810), .CK(clk), .Q(\mem[13][8] ) );
  DFF_X1 \mem_reg[13][7]  ( .D(n809), .CK(clk), .Q(\mem[13][7] ) );
  DFF_X1 \mem_reg[13][6]  ( .D(n808), .CK(clk), .Q(\mem[13][6] ) );
  DFF_X1 \mem_reg[13][5]  ( .D(n807), .CK(clk), .Q(\mem[13][5] ) );
  DFF_X1 \mem_reg[13][4]  ( .D(n806), .CK(clk), .Q(\mem[13][4] ) );
  DFF_X1 \mem_reg[13][3]  ( .D(n805), .CK(clk), .Q(\mem[13][3] ) );
  DFF_X1 \mem_reg[13][2]  ( .D(n804), .CK(clk), .Q(\mem[13][2] ) );
  DFF_X1 \mem_reg[13][1]  ( .D(n803), .CK(clk), .Q(\mem[13][1] ) );
  DFF_X1 \mem_reg[13][0]  ( .D(n802), .CK(clk), .Q(\mem[13][0] ) );
  DFF_X1 \mem_reg[12][15]  ( .D(n801), .CK(clk), .Q(\mem[12][15] ) );
  DFF_X1 \mem_reg[12][14]  ( .D(n800), .CK(clk), .Q(\mem[12][14] ) );
  DFF_X1 \mem_reg[12][13]  ( .D(n799), .CK(clk), .Q(\mem[12][13] ) );
  DFF_X1 \mem_reg[12][12]  ( .D(n798), .CK(clk), .Q(\mem[12][12] ) );
  DFF_X1 \mem_reg[12][11]  ( .D(n797), .CK(clk), .Q(\mem[12][11] ) );
  DFF_X1 \mem_reg[12][10]  ( .D(n796), .CK(clk), .Q(\mem[12][10] ) );
  DFF_X1 \mem_reg[12][9]  ( .D(n795), .CK(clk), .Q(\mem[12][9] ) );
  DFF_X1 \mem_reg[12][8]  ( .D(n794), .CK(clk), .Q(\mem[12][8] ) );
  DFF_X1 \mem_reg[12][7]  ( .D(n793), .CK(clk), .Q(\mem[12][7] ) );
  DFF_X1 \mem_reg[12][6]  ( .D(n792), .CK(clk), .Q(\mem[12][6] ) );
  DFF_X1 \mem_reg[12][5]  ( .D(n791), .CK(clk), .Q(\mem[12][5] ) );
  DFF_X1 \mem_reg[12][4]  ( .D(n790), .CK(clk), .Q(\mem[12][4] ) );
  DFF_X1 \mem_reg[12][3]  ( .D(n789), .CK(clk), .Q(\mem[12][3] ) );
  DFF_X1 \mem_reg[12][2]  ( .D(n788), .CK(clk), .Q(\mem[12][2] ) );
  DFF_X1 \mem_reg[12][1]  ( .D(n787), .CK(clk), .Q(\mem[12][1] ) );
  DFF_X1 \mem_reg[12][0]  ( .D(n786), .CK(clk), .Q(\mem[12][0] ) );
  DFF_X1 \mem_reg[11][15]  ( .D(n785), .CK(clk), .Q(\mem[11][15] ) );
  DFF_X1 \mem_reg[11][14]  ( .D(n784), .CK(clk), .Q(\mem[11][14] ) );
  DFF_X1 \mem_reg[11][13]  ( .D(n783), .CK(clk), .Q(\mem[11][13] ) );
  DFF_X1 \mem_reg[11][12]  ( .D(n782), .CK(clk), .Q(\mem[11][12] ) );
  DFF_X1 \mem_reg[11][11]  ( .D(n781), .CK(clk), .Q(\mem[11][11] ) );
  DFF_X1 \mem_reg[11][10]  ( .D(n780), .CK(clk), .Q(\mem[11][10] ) );
  DFF_X1 \mem_reg[11][9]  ( .D(n779), .CK(clk), .Q(\mem[11][9] ) );
  DFF_X1 \mem_reg[11][8]  ( .D(n778), .CK(clk), .Q(\mem[11][8] ) );
  DFF_X1 \mem_reg[11][7]  ( .D(n777), .CK(clk), .Q(\mem[11][7] ) );
  DFF_X1 \mem_reg[11][6]  ( .D(n776), .CK(clk), .Q(\mem[11][6] ) );
  DFF_X1 \mem_reg[11][5]  ( .D(n775), .CK(clk), .Q(\mem[11][5] ) );
  DFF_X1 \mem_reg[11][4]  ( .D(n774), .CK(clk), .Q(\mem[11][4] ) );
  DFF_X1 \mem_reg[11][3]  ( .D(n773), .CK(clk), .Q(\mem[11][3] ) );
  DFF_X1 \mem_reg[11][2]  ( .D(n772), .CK(clk), .Q(\mem[11][2] ) );
  DFF_X1 \mem_reg[11][1]  ( .D(n771), .CK(clk), .Q(\mem[11][1] ) );
  DFF_X1 \mem_reg[11][0]  ( .D(n770), .CK(clk), .Q(\mem[11][0] ) );
  DFF_X1 \mem_reg[10][15]  ( .D(n769), .CK(clk), .Q(\mem[10][15] ) );
  DFF_X1 \mem_reg[10][14]  ( .D(n768), .CK(clk), .Q(\mem[10][14] ) );
  DFF_X1 \mem_reg[10][13]  ( .D(n767), .CK(clk), .Q(\mem[10][13] ) );
  DFF_X1 \mem_reg[10][12]  ( .D(n766), .CK(clk), .Q(\mem[10][12] ) );
  DFF_X1 \mem_reg[10][11]  ( .D(n765), .CK(clk), .Q(\mem[10][11] ) );
  DFF_X1 \mem_reg[10][10]  ( .D(n764), .CK(clk), .Q(\mem[10][10] ) );
  DFF_X1 \mem_reg[10][9]  ( .D(n763), .CK(clk), .Q(\mem[10][9] ) );
  DFF_X1 \mem_reg[10][8]  ( .D(n762), .CK(clk), .Q(\mem[10][8] ) );
  DFF_X1 \mem_reg[10][7]  ( .D(n761), .CK(clk), .Q(\mem[10][7] ) );
  DFF_X1 \mem_reg[10][6]  ( .D(n760), .CK(clk), .Q(\mem[10][6] ) );
  DFF_X1 \mem_reg[10][5]  ( .D(n759), .CK(clk), .Q(\mem[10][5] ) );
  DFF_X1 \mem_reg[10][4]  ( .D(n758), .CK(clk), .Q(\mem[10][4] ) );
  DFF_X1 \mem_reg[10][3]  ( .D(n757), .CK(clk), .Q(\mem[10][3] ) );
  DFF_X1 \mem_reg[10][2]  ( .D(n756), .CK(clk), .Q(\mem[10][2] ) );
  DFF_X1 \mem_reg[10][1]  ( .D(n755), .CK(clk), .Q(\mem[10][1] ) );
  DFF_X1 \mem_reg[10][0]  ( .D(n754), .CK(clk), .Q(\mem[10][0] ) );
  DFF_X1 \mem_reg[9][15]  ( .D(n753), .CK(clk), .Q(\mem[9][15] ) );
  DFF_X1 \mem_reg[9][14]  ( .D(n752), .CK(clk), .Q(\mem[9][14] ) );
  DFF_X1 \mem_reg[9][13]  ( .D(n751), .CK(clk), .Q(\mem[9][13] ) );
  DFF_X1 \mem_reg[9][12]  ( .D(n750), .CK(clk), .Q(\mem[9][12] ) );
  DFF_X1 \mem_reg[9][11]  ( .D(n749), .CK(clk), .Q(\mem[9][11] ) );
  DFF_X1 \mem_reg[9][10]  ( .D(n748), .CK(clk), .Q(\mem[9][10] ) );
  DFF_X1 \mem_reg[9][9]  ( .D(n747), .CK(clk), .Q(\mem[9][9] ) );
  DFF_X1 \mem_reg[9][8]  ( .D(n746), .CK(clk), .Q(\mem[9][8] ) );
  DFF_X1 \mem_reg[9][7]  ( .D(n745), .CK(clk), .Q(\mem[9][7] ) );
  DFF_X1 \mem_reg[9][6]  ( .D(n744), .CK(clk), .Q(\mem[9][6] ) );
  DFF_X1 \mem_reg[9][5]  ( .D(n743), .CK(clk), .Q(\mem[9][5] ) );
  DFF_X1 \mem_reg[9][4]  ( .D(n742), .CK(clk), .Q(\mem[9][4] ) );
  DFF_X1 \mem_reg[9][3]  ( .D(n741), .CK(clk), .Q(\mem[9][3] ) );
  DFF_X1 \mem_reg[9][2]  ( .D(n740), .CK(clk), .Q(\mem[9][2] ) );
  DFF_X1 \mem_reg[9][1]  ( .D(n739), .CK(clk), .Q(\mem[9][1] ) );
  DFF_X1 \mem_reg[9][0]  ( .D(n738), .CK(clk), .Q(\mem[9][0] ) );
  DFF_X1 \mem_reg[8][15]  ( .D(n737), .CK(clk), .Q(\mem[8][15] ) );
  DFF_X1 \mem_reg[8][14]  ( .D(n736), .CK(clk), .Q(\mem[8][14] ) );
  DFF_X1 \mem_reg[8][13]  ( .D(n735), .CK(clk), .Q(\mem[8][13] ) );
  DFF_X1 \mem_reg[8][12]  ( .D(n734), .CK(clk), .Q(\mem[8][12] ) );
  DFF_X1 \mem_reg[8][11]  ( .D(n733), .CK(clk), .Q(\mem[8][11] ) );
  DFF_X1 \mem_reg[8][10]  ( .D(n732), .CK(clk), .Q(\mem[8][10] ) );
  DFF_X1 \mem_reg[8][9]  ( .D(n731), .CK(clk), .Q(\mem[8][9] ) );
  DFF_X1 \mem_reg[8][8]  ( .D(n730), .CK(clk), .Q(\mem[8][8] ) );
  DFF_X1 \mem_reg[8][7]  ( .D(n729), .CK(clk), .Q(\mem[8][7] ) );
  DFF_X1 \mem_reg[8][6]  ( .D(n728), .CK(clk), .Q(\mem[8][6] ) );
  DFF_X1 \mem_reg[8][5]  ( .D(n727), .CK(clk), .Q(\mem[8][5] ) );
  DFF_X1 \mem_reg[8][4]  ( .D(n726), .CK(clk), .Q(\mem[8][4] ) );
  DFF_X1 \mem_reg[8][3]  ( .D(n725), .CK(clk), .Q(\mem[8][3] ) );
  DFF_X1 \mem_reg[8][2]  ( .D(n724), .CK(clk), .Q(\mem[8][2] ) );
  DFF_X1 \mem_reg[8][1]  ( .D(n723), .CK(clk), .Q(\mem[8][1] ) );
  DFF_X1 \mem_reg[8][0]  ( .D(n722), .CK(clk), .Q(\mem[8][0] ) );
  DFF_X1 \mem_reg[7][15]  ( .D(n721), .CK(clk), .Q(\mem[7][15] ) );
  DFF_X1 \mem_reg[7][14]  ( .D(n720), .CK(clk), .Q(\mem[7][14] ) );
  DFF_X1 \mem_reg[7][13]  ( .D(n719), .CK(clk), .Q(\mem[7][13] ) );
  DFF_X1 \mem_reg[7][12]  ( .D(n718), .CK(clk), .Q(\mem[7][12] ) );
  DFF_X1 \mem_reg[7][11]  ( .D(n717), .CK(clk), .Q(\mem[7][11] ) );
  DFF_X1 \mem_reg[7][10]  ( .D(n716), .CK(clk), .Q(\mem[7][10] ) );
  DFF_X1 \mem_reg[7][9]  ( .D(n715), .CK(clk), .Q(\mem[7][9] ) );
  DFF_X1 \mem_reg[7][8]  ( .D(n714), .CK(clk), .Q(\mem[7][8] ) );
  DFF_X1 \mem_reg[7][7]  ( .D(n713), .CK(clk), .Q(\mem[7][7] ) );
  DFF_X1 \mem_reg[7][6]  ( .D(n712), .CK(clk), .Q(\mem[7][6] ) );
  DFF_X1 \mem_reg[7][5]  ( .D(n711), .CK(clk), .Q(\mem[7][5] ) );
  DFF_X1 \mem_reg[7][4]  ( .D(n710), .CK(clk), .Q(\mem[7][4] ) );
  DFF_X1 \mem_reg[7][3]  ( .D(n709), .CK(clk), .Q(\mem[7][3] ) );
  DFF_X1 \mem_reg[7][2]  ( .D(n708), .CK(clk), .Q(\mem[7][2] ) );
  DFF_X1 \mem_reg[7][1]  ( .D(n707), .CK(clk), .Q(\mem[7][1] ) );
  DFF_X1 \mem_reg[7][0]  ( .D(n706), .CK(clk), .Q(\mem[7][0] ) );
  DFF_X1 \mem_reg[6][15]  ( .D(n705), .CK(clk), .Q(\mem[6][15] ) );
  DFF_X1 \mem_reg[6][14]  ( .D(n704), .CK(clk), .Q(\mem[6][14] ) );
  DFF_X1 \mem_reg[6][13]  ( .D(n703), .CK(clk), .Q(\mem[6][13] ) );
  DFF_X1 \mem_reg[6][12]  ( .D(n702), .CK(clk), .Q(\mem[6][12] ) );
  DFF_X1 \mem_reg[6][11]  ( .D(n701), .CK(clk), .Q(\mem[6][11] ) );
  DFF_X1 \mem_reg[6][10]  ( .D(n700), .CK(clk), .Q(\mem[6][10] ) );
  DFF_X1 \mem_reg[6][9]  ( .D(n699), .CK(clk), .Q(\mem[6][9] ) );
  DFF_X1 \mem_reg[6][8]  ( .D(n698), .CK(clk), .Q(\mem[6][8] ) );
  DFF_X1 \mem_reg[6][7]  ( .D(n697), .CK(clk), .Q(\mem[6][7] ) );
  DFF_X1 \mem_reg[6][6]  ( .D(n696), .CK(clk), .Q(\mem[6][6] ) );
  DFF_X1 \mem_reg[6][5]  ( .D(n695), .CK(clk), .Q(\mem[6][5] ) );
  DFF_X1 \mem_reg[6][4]  ( .D(n694), .CK(clk), .Q(\mem[6][4] ) );
  DFF_X1 \mem_reg[6][3]  ( .D(n693), .CK(clk), .Q(\mem[6][3] ) );
  DFF_X1 \mem_reg[6][2]  ( .D(n692), .CK(clk), .Q(\mem[6][2] ) );
  DFF_X1 \mem_reg[6][1]  ( .D(n691), .CK(clk), .Q(\mem[6][1] ) );
  DFF_X1 \mem_reg[6][0]  ( .D(n690), .CK(clk), .Q(\mem[6][0] ) );
  DFF_X1 \mem_reg[5][15]  ( .D(n689), .CK(clk), .Q(\mem[5][15] ) );
  DFF_X1 \mem_reg[5][14]  ( .D(n688), .CK(clk), .Q(\mem[5][14] ) );
  DFF_X1 \mem_reg[5][13]  ( .D(n687), .CK(clk), .Q(\mem[5][13] ) );
  DFF_X1 \mem_reg[5][12]  ( .D(n686), .CK(clk), .Q(\mem[5][12] ) );
  DFF_X1 \mem_reg[5][11]  ( .D(n685), .CK(clk), .Q(\mem[5][11] ) );
  DFF_X1 \mem_reg[5][10]  ( .D(n684), .CK(clk), .Q(\mem[5][10] ) );
  DFF_X1 \mem_reg[5][9]  ( .D(n683), .CK(clk), .Q(\mem[5][9] ) );
  DFF_X1 \mem_reg[5][8]  ( .D(n682), .CK(clk), .Q(\mem[5][8] ) );
  DFF_X1 \mem_reg[5][7]  ( .D(n681), .CK(clk), .Q(\mem[5][7] ) );
  DFF_X1 \mem_reg[5][6]  ( .D(n680), .CK(clk), .Q(\mem[5][6] ) );
  DFF_X1 \mem_reg[5][5]  ( .D(n679), .CK(clk), .Q(\mem[5][5] ) );
  DFF_X1 \mem_reg[5][4]  ( .D(n678), .CK(clk), .Q(\mem[5][4] ) );
  DFF_X1 \mem_reg[5][3]  ( .D(n677), .CK(clk), .Q(\mem[5][3] ) );
  DFF_X1 \mem_reg[5][2]  ( .D(n676), .CK(clk), .Q(\mem[5][2] ) );
  DFF_X1 \mem_reg[5][1]  ( .D(n675), .CK(clk), .Q(\mem[5][1] ) );
  DFF_X1 \mem_reg[5][0]  ( .D(n674), .CK(clk), .Q(\mem[5][0] ) );
  DFF_X1 \mem_reg[4][15]  ( .D(n673), .CK(clk), .Q(\mem[4][15] ) );
  DFF_X1 \mem_reg[4][14]  ( .D(n672), .CK(clk), .Q(\mem[4][14] ) );
  DFF_X1 \mem_reg[4][13]  ( .D(n671), .CK(clk), .Q(\mem[4][13] ) );
  DFF_X1 \mem_reg[4][12]  ( .D(n670), .CK(clk), .Q(\mem[4][12] ) );
  DFF_X1 \mem_reg[4][11]  ( .D(n669), .CK(clk), .Q(\mem[4][11] ) );
  DFF_X1 \mem_reg[4][10]  ( .D(n668), .CK(clk), .Q(\mem[4][10] ) );
  DFF_X1 \mem_reg[4][9]  ( .D(n667), .CK(clk), .Q(\mem[4][9] ) );
  DFF_X1 \mem_reg[4][8]  ( .D(n666), .CK(clk), .Q(\mem[4][8] ) );
  DFF_X1 \mem_reg[4][7]  ( .D(n665), .CK(clk), .Q(\mem[4][7] ) );
  DFF_X1 \mem_reg[4][6]  ( .D(n664), .CK(clk), .Q(\mem[4][6] ) );
  DFF_X1 \mem_reg[4][5]  ( .D(n663), .CK(clk), .Q(\mem[4][5] ) );
  DFF_X1 \mem_reg[4][4]  ( .D(n662), .CK(clk), .Q(\mem[4][4] ) );
  DFF_X1 \mem_reg[4][3]  ( .D(n661), .CK(clk), .Q(\mem[4][3] ) );
  DFF_X1 \mem_reg[4][2]  ( .D(n660), .CK(clk), .Q(\mem[4][2] ) );
  DFF_X1 \mem_reg[4][1]  ( .D(n659), .CK(clk), .Q(\mem[4][1] ) );
  DFF_X1 \mem_reg[4][0]  ( .D(n658), .CK(clk), .Q(\mem[4][0] ) );
  DFF_X1 \mem_reg[3][15]  ( .D(n657), .CK(clk), .Q(\mem[3][15] ) );
  DFF_X1 \mem_reg[3][14]  ( .D(n656), .CK(clk), .Q(\mem[3][14] ) );
  DFF_X1 \mem_reg[3][13]  ( .D(n655), .CK(clk), .Q(\mem[3][13] ) );
  DFF_X1 \mem_reg[3][12]  ( .D(n654), .CK(clk), .Q(\mem[3][12] ) );
  DFF_X1 \mem_reg[3][11]  ( .D(n653), .CK(clk), .Q(\mem[3][11] ) );
  DFF_X1 \mem_reg[3][10]  ( .D(n652), .CK(clk), .Q(\mem[3][10] ) );
  DFF_X1 \mem_reg[3][9]  ( .D(n651), .CK(clk), .Q(\mem[3][9] ) );
  DFF_X1 \mem_reg[3][8]  ( .D(n650), .CK(clk), .Q(\mem[3][8] ) );
  DFF_X1 \mem_reg[3][7]  ( .D(n649), .CK(clk), .Q(\mem[3][7] ) );
  DFF_X1 \mem_reg[3][6]  ( .D(n648), .CK(clk), .Q(\mem[3][6] ) );
  DFF_X1 \mem_reg[3][5]  ( .D(n647), .CK(clk), .Q(\mem[3][5] ) );
  DFF_X1 \mem_reg[3][4]  ( .D(n646), .CK(clk), .Q(\mem[3][4] ) );
  DFF_X1 \mem_reg[3][3]  ( .D(n645), .CK(clk), .Q(\mem[3][3] ) );
  DFF_X1 \mem_reg[3][2]  ( .D(n644), .CK(clk), .Q(\mem[3][2] ) );
  DFF_X1 \mem_reg[3][1]  ( .D(n643), .CK(clk), .Q(\mem[3][1] ) );
  DFF_X1 \mem_reg[3][0]  ( .D(n642), .CK(clk), .Q(\mem[3][0] ) );
  DFF_X1 \mem_reg[2][15]  ( .D(n641), .CK(clk), .Q(\mem[2][15] ) );
  DFF_X1 \mem_reg[2][14]  ( .D(n640), .CK(clk), .Q(\mem[2][14] ) );
  DFF_X1 \mem_reg[2][13]  ( .D(n639), .CK(clk), .Q(\mem[2][13] ) );
  DFF_X1 \mem_reg[2][12]  ( .D(n638), .CK(clk), .Q(\mem[2][12] ) );
  DFF_X1 \mem_reg[2][11]  ( .D(n637), .CK(clk), .Q(\mem[2][11] ) );
  DFF_X1 \mem_reg[2][10]  ( .D(n636), .CK(clk), .Q(\mem[2][10] ) );
  DFF_X1 \mem_reg[2][9]  ( .D(n635), .CK(clk), .Q(\mem[2][9] ) );
  DFF_X1 \mem_reg[2][8]  ( .D(n634), .CK(clk), .Q(\mem[2][8] ) );
  DFF_X1 \mem_reg[2][7]  ( .D(n633), .CK(clk), .Q(\mem[2][7] ) );
  DFF_X1 \mem_reg[2][6]  ( .D(n632), .CK(clk), .Q(\mem[2][6] ) );
  DFF_X1 \mem_reg[2][5]  ( .D(n631), .CK(clk), .Q(\mem[2][5] ) );
  DFF_X1 \mem_reg[2][4]  ( .D(n630), .CK(clk), .Q(\mem[2][4] ) );
  DFF_X1 \mem_reg[2][3]  ( .D(n629), .CK(clk), .Q(\mem[2][3] ) );
  DFF_X1 \mem_reg[2][2]  ( .D(n628), .CK(clk), .Q(\mem[2][2] ) );
  DFF_X1 \mem_reg[2][1]  ( .D(n627), .CK(clk), .Q(\mem[2][1] ) );
  DFF_X1 \mem_reg[2][0]  ( .D(n626), .CK(clk), .Q(\mem[2][0] ) );
  DFF_X1 \mem_reg[1][15]  ( .D(n625), .CK(clk), .Q(\mem[1][15] ) );
  DFF_X1 \mem_reg[1][14]  ( .D(n624), .CK(clk), .Q(\mem[1][14] ) );
  DFF_X1 \mem_reg[1][13]  ( .D(n623), .CK(clk), .Q(\mem[1][13] ) );
  DFF_X1 \mem_reg[1][12]  ( .D(n622), .CK(clk), .Q(\mem[1][12] ) );
  DFF_X1 \mem_reg[1][11]  ( .D(n621), .CK(clk), .Q(\mem[1][11] ) );
  DFF_X1 \mem_reg[1][10]  ( .D(n620), .CK(clk), .Q(\mem[1][10] ) );
  DFF_X1 \mem_reg[1][9]  ( .D(n619), .CK(clk), .Q(\mem[1][9] ) );
  DFF_X1 \mem_reg[1][8]  ( .D(n618), .CK(clk), .Q(\mem[1][8] ) );
  DFF_X1 \mem_reg[1][7]  ( .D(n617), .CK(clk), .Q(\mem[1][7] ) );
  DFF_X1 \mem_reg[1][6]  ( .D(n616), .CK(clk), .Q(\mem[1][6] ) );
  DFF_X1 \mem_reg[1][5]  ( .D(n615), .CK(clk), .Q(\mem[1][5] ) );
  DFF_X1 \mem_reg[1][4]  ( .D(n614), .CK(clk), .Q(\mem[1][4] ) );
  DFF_X1 \mem_reg[1][3]  ( .D(n613), .CK(clk), .Q(\mem[1][3] ) );
  DFF_X1 \mem_reg[1][2]  ( .D(n612), .CK(clk), .Q(\mem[1][2] ) );
  DFF_X1 \mem_reg[1][1]  ( .D(n611), .CK(clk), .Q(\mem[1][1] ) );
  DFF_X1 \mem_reg[1][0]  ( .D(n610), .CK(clk), .Q(\mem[1][0] ) );
  DFF_X1 \mem_reg[0][15]  ( .D(n609), .CK(clk), .Q(\mem[0][15] ) );
  DFF_X1 \mem_reg[0][14]  ( .D(n608), .CK(clk), .Q(\mem[0][14] ) );
  DFF_X1 \mem_reg[0][13]  ( .D(n607), .CK(clk), .Q(\mem[0][13] ) );
  DFF_X1 \mem_reg[0][12]  ( .D(n606), .CK(clk), .Q(\mem[0][12] ) );
  DFF_X1 \mem_reg[0][11]  ( .D(n605), .CK(clk), .Q(\mem[0][11] ) );
  DFF_X1 \mem_reg[0][10]  ( .D(n604), .CK(clk), .Q(\mem[0][10] ) );
  DFF_X1 \mem_reg[0][9]  ( .D(n603), .CK(clk), .Q(\mem[0][9] ) );
  DFF_X1 \mem_reg[0][8]  ( .D(n602), .CK(clk), .Q(\mem[0][8] ) );
  DFF_X1 \mem_reg[0][7]  ( .D(n601), .CK(clk), .Q(\mem[0][7] ) );
  DFF_X1 \mem_reg[0][6]  ( .D(n600), .CK(clk), .Q(\mem[0][6] ) );
  DFF_X1 \mem_reg[0][5]  ( .D(n599), .CK(clk), .Q(\mem[0][5] ) );
  DFF_X1 \mem_reg[0][4]  ( .D(n598), .CK(clk), .Q(\mem[0][4] ) );
  DFF_X1 \mem_reg[0][3]  ( .D(n597), .CK(clk), .Q(\mem[0][3] ) );
  DFF_X1 \mem_reg[0][2]  ( .D(n596), .CK(clk), .Q(\mem[0][2] ) );
  DFF_X1 \mem_reg[0][1]  ( .D(n595), .CK(clk), .Q(\mem[0][1] ) );
  DFF_X1 \mem_reg[0][0]  ( .D(n594), .CK(clk), .Q(\mem[0][0] ) );
  CLKBUF_X1 U3 ( .A(n1553), .Z(n1548) );
  BUF_X1 U4 ( .A(n1553), .Z(n1550) );
  CLKBUF_X1 U5 ( .A(n1553), .Z(n1549) );
  BUF_X1 U6 ( .A(n1543), .Z(n1545) );
  BUF_X1 U7 ( .A(n1553), .Z(n1551) );
  BUF_X1 U8 ( .A(n1552), .Z(n1543) );
  BUF_X1 U9 ( .A(n1550), .Z(n1544) );
  BUF_X1 U10 ( .A(n1553), .Z(n1546) );
  BUF_X1 U11 ( .A(n1553), .Z(n1547) );
  BUF_X1 U12 ( .A(n1542), .Z(n1540) );
  BUF_X1 U13 ( .A(n1542), .Z(n1541) );
  BUF_X1 U14 ( .A(N11), .Z(n1538) );
  BUF_X1 U15 ( .A(N11), .Z(n1539) );
  BUF_X1 U16 ( .A(n1552), .Z(n1553) );
  INV_X1 U17 ( .A(n578), .ZN(n1621) );
  BUF_X1 U18 ( .A(n338), .Z(n1583) );
  BUF_X1 U19 ( .A(n355), .Z(n1582) );
  BUF_X1 U20 ( .A(n372), .Z(n1581) );
  BUF_X1 U21 ( .A(n457), .Z(n1576) );
  BUF_X1 U22 ( .A(n475), .Z(n1575) );
  BUF_X1 U23 ( .A(n492), .Z(n1574) );
  BUF_X1 U24 ( .A(n509), .Z(n1573) );
  BUF_X1 U25 ( .A(n389), .Z(n1580) );
  BUF_X1 U26 ( .A(n406), .Z(n1579) );
  BUF_X1 U27 ( .A(n440), .Z(n1577) );
  BUF_X1 U28 ( .A(n543), .Z(n1571) );
  BUF_X1 U29 ( .A(n560), .Z(n1570) );
  BUF_X1 U30 ( .A(n320), .Z(n1584) );
  BUF_X1 U31 ( .A(n423), .Z(n1578) );
  BUF_X1 U32 ( .A(n526), .Z(n1572) );
  BUF_X1 U33 ( .A(N11), .Z(n1542) );
  BUF_X1 U34 ( .A(N10), .Z(n1552) );
  BUF_X1 U35 ( .A(N13), .Z(n1533) );
  NAND2_X1 U36 ( .A1(n474), .A2(n182), .ZN(n578) );
  BUF_X1 U37 ( .A(n38), .Z(n1600) );
  BUF_X1 U38 ( .A(n218), .Z(n1590) );
  BUF_X1 U39 ( .A(n235), .Z(n1589) );
  BUF_X1 U40 ( .A(n57), .Z(n1599) );
  BUF_X1 U41 ( .A(n75), .Z(n1598) );
  BUF_X1 U42 ( .A(n93), .Z(n1597) );
  BUF_X1 U43 ( .A(n111), .Z(n1596) );
  BUF_X1 U44 ( .A(n165), .Z(n1593) );
  BUF_X1 U45 ( .A(n252), .Z(n1588) );
  BUF_X1 U46 ( .A(n269), .Z(n1587) );
  BUF_X1 U47 ( .A(n286), .Z(n1586) );
  BUF_X1 U48 ( .A(n303), .Z(n1585) );
  BUF_X1 U49 ( .A(n201), .Z(n1591) );
  BUF_X1 U50 ( .A(n129), .Z(n1595) );
  BUF_X1 U51 ( .A(n183), .Z(n1592) );
  BUF_X1 U52 ( .A(n147), .Z(n1594) );
  NAND2_X1 U53 ( .A1(n337), .A2(n55), .ZN(n320) );
  NAND2_X1 U54 ( .A1(n337), .A2(n74), .ZN(n338) );
  NAND2_X1 U55 ( .A1(n337), .A2(n92), .ZN(n355) );
  NAND2_X1 U56 ( .A1(n337), .A2(n110), .ZN(n372) );
  NAND2_X1 U57 ( .A1(n474), .A2(n55), .ZN(n457) );
  NAND2_X1 U58 ( .A1(n474), .A2(n74), .ZN(n475) );
  NAND2_X1 U59 ( .A1(n474), .A2(n92), .ZN(n492) );
  NAND2_X1 U60 ( .A1(n474), .A2(n110), .ZN(n509) );
  NAND2_X1 U61 ( .A1(n337), .A2(n128), .ZN(n389) );
  NAND2_X1 U62 ( .A1(n337), .A2(n146), .ZN(n406) );
  NAND2_X1 U63 ( .A1(n337), .A2(n164), .ZN(n423) );
  NAND2_X1 U64 ( .A1(n337), .A2(n182), .ZN(n440) );
  NAND2_X1 U65 ( .A1(n474), .A2(n128), .ZN(n526) );
  NAND2_X1 U66 ( .A1(n474), .A2(n146), .ZN(n543) );
  NAND2_X1 U67 ( .A1(n474), .A2(n164), .ZN(n560) );
  AND3_X1 U68 ( .A1(wr_en), .A2(n1603), .A3(N14), .ZN(n337) );
  AND3_X1 U69 ( .A1(N13), .A2(wr_en), .A3(N14), .ZN(n474) );
  AND3_X1 U70 ( .A1(N11), .A2(N10), .A3(N12), .ZN(n182) );
  NAND2_X1 U71 ( .A1(n55), .A2(n56), .ZN(n38) );
  NAND2_X1 U72 ( .A1(n74), .A2(n56), .ZN(n57) );
  NAND2_X1 U73 ( .A1(n92), .A2(n56), .ZN(n75) );
  NAND2_X1 U74 ( .A1(n110), .A2(n56), .ZN(n93) );
  NAND2_X1 U75 ( .A1(n200), .A2(n55), .ZN(n183) );
  NAND2_X1 U76 ( .A1(n200), .A2(n74), .ZN(n201) );
  NAND2_X1 U77 ( .A1(n200), .A2(n92), .ZN(n218) );
  NAND2_X1 U78 ( .A1(n200), .A2(n110), .ZN(n235) );
  NAND2_X1 U79 ( .A1(n128), .A2(n56), .ZN(n111) );
  NAND2_X1 U80 ( .A1(n146), .A2(n56), .ZN(n129) );
  NAND2_X1 U81 ( .A1(n164), .A2(n56), .ZN(n147) );
  NAND2_X1 U82 ( .A1(n182), .A2(n56), .ZN(n165) );
  NAND2_X1 U83 ( .A1(n200), .A2(n128), .ZN(n252) );
  NAND2_X1 U84 ( .A1(n200), .A2(n146), .ZN(n269) );
  NAND2_X1 U85 ( .A1(n200), .A2(n164), .ZN(n286) );
  NAND2_X1 U86 ( .A1(n200), .A2(n182), .ZN(n303) );
  NOR3_X1 U87 ( .A1(N11), .A2(N12), .A3(N10), .ZN(n55) );
  NOR3_X1 U88 ( .A1(N11), .A2(N12), .A3(n1601), .ZN(n74) );
  NOR3_X1 U89 ( .A1(N10), .A2(N12), .A3(n1602), .ZN(n92) );
  NOR3_X1 U90 ( .A1(n1601), .A2(N12), .A3(n1602), .ZN(n110) );
  AND3_X1 U91 ( .A1(n1601), .A2(n1602), .A3(N12), .ZN(n128) );
  AND3_X1 U92 ( .A1(N10), .A2(n1602), .A3(N12), .ZN(n146) );
  AND3_X1 U93 ( .A1(N11), .A2(n1601), .A3(N12), .ZN(n164) );
  AND3_X1 U94 ( .A1(n1603), .A2(n1604), .A3(wr_en), .ZN(n56) );
  AND3_X1 U95 ( .A1(wr_en), .A2(n1604), .A3(N13), .ZN(n200) );
  BUF_X1 U96 ( .A(n1637), .Z(n1569) );
  BUF_X1 U97 ( .A(n1636), .Z(n1568) );
  BUF_X1 U98 ( .A(n1635), .Z(n1567) );
  BUF_X1 U99 ( .A(n1634), .Z(n1566) );
  BUF_X1 U100 ( .A(n1633), .Z(n1565) );
  BUF_X1 U101 ( .A(n1632), .Z(n1564) );
  BUF_X1 U102 ( .A(n1631), .Z(n1563) );
  BUF_X1 U103 ( .A(n1630), .Z(n1562) );
  BUF_X1 U104 ( .A(n1628), .Z(n1560) );
  BUF_X1 U105 ( .A(n1627), .Z(n1559) );
  BUF_X1 U106 ( .A(n1626), .Z(n1558) );
  BUF_X1 U107 ( .A(n1625), .Z(n1557) );
  BUF_X1 U108 ( .A(n1624), .Z(n1556) );
  BUF_X1 U109 ( .A(n1623), .Z(n1555) );
  BUF_X1 U110 ( .A(n1622), .Z(n1554) );
  BUF_X1 U111 ( .A(n1629), .Z(n1561) );
  OAI21_X1 U112 ( .B1(n1562), .B2(n57), .A(n65), .ZN(n617) );
  NAND2_X1 U113 ( .A1(\mem[1][7] ), .A2(n1599), .ZN(n65) );
  OAI21_X1 U114 ( .B1(n1629), .B2(n1599), .A(n66), .ZN(n618) );
  NAND2_X1 U115 ( .A1(\mem[1][8] ), .A2(n1599), .ZN(n66) );
  OAI21_X1 U116 ( .B1(n1560), .B2(n57), .A(n67), .ZN(n619) );
  NAND2_X1 U117 ( .A1(\mem[1][9] ), .A2(n1599), .ZN(n67) );
  OAI21_X1 U118 ( .B1(n1559), .B2(n57), .A(n68), .ZN(n620) );
  NAND2_X1 U119 ( .A1(\mem[1][10] ), .A2(n1599), .ZN(n68) );
  OAI21_X1 U120 ( .B1(n1558), .B2(n57), .A(n69), .ZN(n621) );
  NAND2_X1 U121 ( .A1(\mem[1][11] ), .A2(n1599), .ZN(n69) );
  OAI21_X1 U122 ( .B1(n1557), .B2(n57), .A(n70), .ZN(n622) );
  NAND2_X1 U123 ( .A1(\mem[1][12] ), .A2(n1599), .ZN(n70) );
  OAI21_X1 U124 ( .B1(n1556), .B2(n57), .A(n71), .ZN(n623) );
  NAND2_X1 U125 ( .A1(\mem[1][13] ), .A2(n1599), .ZN(n71) );
  OAI21_X1 U126 ( .B1(n1555), .B2(n57), .A(n72), .ZN(n624) );
  NAND2_X1 U127 ( .A1(\mem[1][14] ), .A2(n1599), .ZN(n72) );
  OAI21_X1 U128 ( .B1(n1562), .B2(n75), .A(n83), .ZN(n633) );
  NAND2_X1 U129 ( .A1(\mem[2][7] ), .A2(n1598), .ZN(n83) );
  OAI21_X1 U130 ( .B1(n1629), .B2(n1598), .A(n84), .ZN(n634) );
  NAND2_X1 U131 ( .A1(\mem[2][8] ), .A2(n1598), .ZN(n84) );
  OAI21_X1 U132 ( .B1(n1560), .B2(n75), .A(n85), .ZN(n635) );
  NAND2_X1 U133 ( .A1(\mem[2][9] ), .A2(n1598), .ZN(n85) );
  OAI21_X1 U134 ( .B1(n1559), .B2(n75), .A(n86), .ZN(n636) );
  NAND2_X1 U135 ( .A1(\mem[2][10] ), .A2(n1598), .ZN(n86) );
  OAI21_X1 U136 ( .B1(n1558), .B2(n75), .A(n87), .ZN(n637) );
  NAND2_X1 U137 ( .A1(\mem[2][11] ), .A2(n1598), .ZN(n87) );
  OAI21_X1 U138 ( .B1(n1557), .B2(n75), .A(n88), .ZN(n638) );
  NAND2_X1 U139 ( .A1(\mem[2][12] ), .A2(n1598), .ZN(n88) );
  OAI21_X1 U140 ( .B1(n1556), .B2(n75), .A(n89), .ZN(n639) );
  NAND2_X1 U141 ( .A1(\mem[2][13] ), .A2(n1598), .ZN(n89) );
  OAI21_X1 U142 ( .B1(n1555), .B2(n75), .A(n90), .ZN(n640) );
  NAND2_X1 U143 ( .A1(\mem[2][14] ), .A2(n1598), .ZN(n90) );
  OAI21_X1 U144 ( .B1(n1562), .B2(n93), .A(n101), .ZN(n649) );
  NAND2_X1 U145 ( .A1(\mem[3][7] ), .A2(n1597), .ZN(n101) );
  OAI21_X1 U146 ( .B1(n1629), .B2(n1597), .A(n102), .ZN(n650) );
  NAND2_X1 U147 ( .A1(\mem[3][8] ), .A2(n1597), .ZN(n102) );
  OAI21_X1 U148 ( .B1(n1560), .B2(n93), .A(n103), .ZN(n651) );
  NAND2_X1 U149 ( .A1(\mem[3][9] ), .A2(n1597), .ZN(n103) );
  OAI21_X1 U150 ( .B1(n1559), .B2(n93), .A(n104), .ZN(n652) );
  NAND2_X1 U151 ( .A1(\mem[3][10] ), .A2(n1597), .ZN(n104) );
  OAI21_X1 U152 ( .B1(n1558), .B2(n93), .A(n105), .ZN(n653) );
  NAND2_X1 U153 ( .A1(\mem[3][11] ), .A2(n1597), .ZN(n105) );
  OAI21_X1 U154 ( .B1(n1557), .B2(n93), .A(n106), .ZN(n654) );
  NAND2_X1 U155 ( .A1(\mem[3][12] ), .A2(n1597), .ZN(n106) );
  OAI21_X1 U156 ( .B1(n1556), .B2(n93), .A(n107), .ZN(n655) );
  NAND2_X1 U157 ( .A1(\mem[3][13] ), .A2(n1597), .ZN(n107) );
  OAI21_X1 U158 ( .B1(n1555), .B2(n93), .A(n108), .ZN(n656) );
  NAND2_X1 U159 ( .A1(\mem[3][14] ), .A2(n1597), .ZN(n108) );
  OAI21_X1 U160 ( .B1(n1562), .B2(n1592), .A(n191), .ZN(n729) );
  NAND2_X1 U161 ( .A1(\mem[8][7] ), .A2(n1592), .ZN(n191) );
  OAI21_X1 U162 ( .B1(n1629), .B2(n1592), .A(n192), .ZN(n730) );
  NAND2_X1 U163 ( .A1(\mem[8][8] ), .A2(n183), .ZN(n192) );
  OAI21_X1 U164 ( .B1(n1560), .B2(n1592), .A(n193), .ZN(n731) );
  NAND2_X1 U165 ( .A1(\mem[8][9] ), .A2(n183), .ZN(n193) );
  OAI21_X1 U166 ( .B1(n1559), .B2(n1592), .A(n194), .ZN(n732) );
  NAND2_X1 U167 ( .A1(\mem[8][10] ), .A2(n183), .ZN(n194) );
  OAI21_X1 U168 ( .B1(n1558), .B2(n1592), .A(n195), .ZN(n733) );
  NAND2_X1 U169 ( .A1(\mem[8][11] ), .A2(n183), .ZN(n195) );
  OAI21_X1 U170 ( .B1(n1557), .B2(n1592), .A(n196), .ZN(n734) );
  NAND2_X1 U171 ( .A1(\mem[8][12] ), .A2(n183), .ZN(n196) );
  OAI21_X1 U172 ( .B1(n1556), .B2(n1592), .A(n197), .ZN(n735) );
  NAND2_X1 U173 ( .A1(\mem[8][13] ), .A2(n183), .ZN(n197) );
  OAI21_X1 U174 ( .B1(n1555), .B2(n1592), .A(n198), .ZN(n736) );
  NAND2_X1 U175 ( .A1(\mem[8][14] ), .A2(n183), .ZN(n198) );
  OAI21_X1 U176 ( .B1(n1562), .B2(n201), .A(n209), .ZN(n745) );
  NAND2_X1 U177 ( .A1(\mem[9][7] ), .A2(n1591), .ZN(n209) );
  OAI21_X1 U178 ( .B1(n1629), .B2(n201), .A(n210), .ZN(n746) );
  NAND2_X1 U179 ( .A1(\mem[9][8] ), .A2(n1591), .ZN(n210) );
  OAI21_X1 U180 ( .B1(n1560), .B2(n201), .A(n211), .ZN(n747) );
  NAND2_X1 U181 ( .A1(\mem[9][9] ), .A2(n201), .ZN(n211) );
  OAI21_X1 U182 ( .B1(n1559), .B2(n201), .A(n212), .ZN(n748) );
  NAND2_X1 U183 ( .A1(\mem[9][10] ), .A2(n201), .ZN(n212) );
  OAI21_X1 U184 ( .B1(n1558), .B2(n201), .A(n213), .ZN(n749) );
  NAND2_X1 U185 ( .A1(\mem[9][11] ), .A2(n201), .ZN(n213) );
  OAI21_X1 U186 ( .B1(n1557), .B2(n201), .A(n214), .ZN(n750) );
  NAND2_X1 U187 ( .A1(\mem[9][12] ), .A2(n1591), .ZN(n214) );
  OAI21_X1 U188 ( .B1(n1556), .B2(n201), .A(n215), .ZN(n751) );
  NAND2_X1 U189 ( .A1(\mem[9][13] ), .A2(n201), .ZN(n215) );
  OAI21_X1 U190 ( .B1(n1555), .B2(n201), .A(n216), .ZN(n752) );
  NAND2_X1 U191 ( .A1(\mem[9][14] ), .A2(n201), .ZN(n216) );
  OAI21_X1 U192 ( .B1(n1562), .B2(n218), .A(n226), .ZN(n761) );
  NAND2_X1 U193 ( .A1(\mem[10][7] ), .A2(n1590), .ZN(n226) );
  OAI21_X1 U194 ( .B1(n1629), .B2(n1590), .A(n227), .ZN(n762) );
  NAND2_X1 U195 ( .A1(\mem[10][8] ), .A2(n1590), .ZN(n227) );
  OAI21_X1 U196 ( .B1(n1560), .B2(n218), .A(n228), .ZN(n763) );
  NAND2_X1 U197 ( .A1(\mem[10][9] ), .A2(n1590), .ZN(n228) );
  OAI21_X1 U198 ( .B1(n1559), .B2(n218), .A(n229), .ZN(n764) );
  NAND2_X1 U199 ( .A1(\mem[10][10] ), .A2(n1590), .ZN(n229) );
  OAI21_X1 U200 ( .B1(n1558), .B2(n218), .A(n230), .ZN(n765) );
  NAND2_X1 U201 ( .A1(\mem[10][11] ), .A2(n1590), .ZN(n230) );
  OAI21_X1 U202 ( .B1(n1557), .B2(n218), .A(n231), .ZN(n766) );
  NAND2_X1 U203 ( .A1(\mem[10][12] ), .A2(n1590), .ZN(n231) );
  OAI21_X1 U204 ( .B1(n1556), .B2(n218), .A(n232), .ZN(n767) );
  NAND2_X1 U205 ( .A1(\mem[10][13] ), .A2(n1590), .ZN(n232) );
  OAI21_X1 U206 ( .B1(n1555), .B2(n218), .A(n233), .ZN(n768) );
  NAND2_X1 U207 ( .A1(\mem[10][14] ), .A2(n1590), .ZN(n233) );
  OAI21_X1 U208 ( .B1(n1562), .B2(n235), .A(n243), .ZN(n777) );
  NAND2_X1 U209 ( .A1(\mem[11][7] ), .A2(n1589), .ZN(n243) );
  OAI21_X1 U210 ( .B1(n1629), .B2(n1589), .A(n244), .ZN(n778) );
  NAND2_X1 U211 ( .A1(\mem[11][8] ), .A2(n1589), .ZN(n244) );
  OAI21_X1 U212 ( .B1(n1560), .B2(n235), .A(n245), .ZN(n779) );
  NAND2_X1 U213 ( .A1(\mem[11][9] ), .A2(n1589), .ZN(n245) );
  OAI21_X1 U214 ( .B1(n1559), .B2(n235), .A(n246), .ZN(n780) );
  NAND2_X1 U215 ( .A1(\mem[11][10] ), .A2(n1589), .ZN(n246) );
  OAI21_X1 U216 ( .B1(n1558), .B2(n235), .A(n247), .ZN(n781) );
  NAND2_X1 U217 ( .A1(\mem[11][11] ), .A2(n1589), .ZN(n247) );
  OAI21_X1 U218 ( .B1(n1557), .B2(n235), .A(n248), .ZN(n782) );
  NAND2_X1 U219 ( .A1(\mem[11][12] ), .A2(n1589), .ZN(n248) );
  OAI21_X1 U220 ( .B1(n1556), .B2(n235), .A(n249), .ZN(n783) );
  NAND2_X1 U221 ( .A1(\mem[11][13] ), .A2(n1589), .ZN(n249) );
  OAI21_X1 U222 ( .B1(n1555), .B2(n235), .A(n250), .ZN(n784) );
  NAND2_X1 U223 ( .A1(\mem[11][14] ), .A2(n1589), .ZN(n250) );
  OAI21_X1 U224 ( .B1(n1630), .B2(n320), .A(n328), .ZN(n857) );
  NAND2_X1 U225 ( .A1(\mem[16][7] ), .A2(n1584), .ZN(n328) );
  OAI21_X1 U226 ( .B1(n1561), .B2(n320), .A(n329), .ZN(n858) );
  NAND2_X1 U227 ( .A1(\mem[16][8] ), .A2(n1584), .ZN(n329) );
  OAI21_X1 U228 ( .B1(n1628), .B2(n320), .A(n330), .ZN(n859) );
  NAND2_X1 U229 ( .A1(\mem[16][9] ), .A2(n320), .ZN(n330) );
  OAI21_X1 U230 ( .B1(n1627), .B2(n320), .A(n331), .ZN(n860) );
  NAND2_X1 U231 ( .A1(\mem[16][10] ), .A2(n320), .ZN(n331) );
  OAI21_X1 U232 ( .B1(n1626), .B2(n320), .A(n332), .ZN(n861) );
  NAND2_X1 U233 ( .A1(\mem[16][11] ), .A2(n320), .ZN(n332) );
  OAI21_X1 U234 ( .B1(n1625), .B2(n320), .A(n333), .ZN(n862) );
  NAND2_X1 U235 ( .A1(\mem[16][12] ), .A2(n1584), .ZN(n333) );
  OAI21_X1 U236 ( .B1(n1624), .B2(n320), .A(n334), .ZN(n863) );
  NAND2_X1 U237 ( .A1(\mem[16][13] ), .A2(n320), .ZN(n334) );
  OAI21_X1 U238 ( .B1(n1623), .B2(n320), .A(n335), .ZN(n864) );
  NAND2_X1 U239 ( .A1(\mem[16][14] ), .A2(n320), .ZN(n335) );
  OAI21_X1 U240 ( .B1(n1630), .B2(n338), .A(n346), .ZN(n873) );
  NAND2_X1 U241 ( .A1(\mem[17][7] ), .A2(n1583), .ZN(n346) );
  OAI21_X1 U242 ( .B1(n1561), .B2(n1583), .A(n347), .ZN(n874) );
  NAND2_X1 U243 ( .A1(\mem[17][8] ), .A2(n1583), .ZN(n347) );
  OAI21_X1 U244 ( .B1(n1628), .B2(n338), .A(n348), .ZN(n875) );
  NAND2_X1 U245 ( .A1(\mem[17][9] ), .A2(n1583), .ZN(n348) );
  OAI21_X1 U246 ( .B1(n1627), .B2(n338), .A(n349), .ZN(n876) );
  NAND2_X1 U247 ( .A1(\mem[17][10] ), .A2(n1583), .ZN(n349) );
  OAI21_X1 U248 ( .B1(n1626), .B2(n338), .A(n350), .ZN(n877) );
  NAND2_X1 U249 ( .A1(\mem[17][11] ), .A2(n1583), .ZN(n350) );
  OAI21_X1 U250 ( .B1(n1625), .B2(n338), .A(n351), .ZN(n878) );
  NAND2_X1 U251 ( .A1(\mem[17][12] ), .A2(n1583), .ZN(n351) );
  OAI21_X1 U252 ( .B1(n1624), .B2(n338), .A(n352), .ZN(n879) );
  NAND2_X1 U253 ( .A1(\mem[17][13] ), .A2(n1583), .ZN(n352) );
  OAI21_X1 U254 ( .B1(n1623), .B2(n338), .A(n353), .ZN(n880) );
  NAND2_X1 U255 ( .A1(\mem[17][14] ), .A2(n1583), .ZN(n353) );
  OAI21_X1 U256 ( .B1(n1630), .B2(n355), .A(n363), .ZN(n889) );
  NAND2_X1 U257 ( .A1(\mem[18][7] ), .A2(n1582), .ZN(n363) );
  OAI21_X1 U258 ( .B1(n1561), .B2(n1582), .A(n364), .ZN(n890) );
  NAND2_X1 U259 ( .A1(\mem[18][8] ), .A2(n1582), .ZN(n364) );
  OAI21_X1 U260 ( .B1(n1628), .B2(n355), .A(n365), .ZN(n891) );
  NAND2_X1 U261 ( .A1(\mem[18][9] ), .A2(n1582), .ZN(n365) );
  OAI21_X1 U262 ( .B1(n1627), .B2(n355), .A(n366), .ZN(n892) );
  NAND2_X1 U263 ( .A1(\mem[18][10] ), .A2(n1582), .ZN(n366) );
  OAI21_X1 U264 ( .B1(n1626), .B2(n355), .A(n367), .ZN(n893) );
  NAND2_X1 U265 ( .A1(\mem[18][11] ), .A2(n1582), .ZN(n367) );
  OAI21_X1 U266 ( .B1(n1625), .B2(n355), .A(n368), .ZN(n894) );
  NAND2_X1 U267 ( .A1(\mem[18][12] ), .A2(n1582), .ZN(n368) );
  OAI21_X1 U268 ( .B1(n1624), .B2(n355), .A(n369), .ZN(n895) );
  NAND2_X1 U269 ( .A1(\mem[18][13] ), .A2(n1582), .ZN(n369) );
  OAI21_X1 U270 ( .B1(n1623), .B2(n355), .A(n370), .ZN(n896) );
  NAND2_X1 U271 ( .A1(\mem[18][14] ), .A2(n1582), .ZN(n370) );
  OAI21_X1 U272 ( .B1(n1630), .B2(n372), .A(n380), .ZN(n905) );
  NAND2_X1 U273 ( .A1(\mem[19][7] ), .A2(n1581), .ZN(n380) );
  OAI21_X1 U274 ( .B1(n1561), .B2(n1581), .A(n381), .ZN(n906) );
  NAND2_X1 U275 ( .A1(\mem[19][8] ), .A2(n1581), .ZN(n381) );
  OAI21_X1 U276 ( .B1(n1628), .B2(n372), .A(n382), .ZN(n907) );
  NAND2_X1 U277 ( .A1(\mem[19][9] ), .A2(n1581), .ZN(n382) );
  OAI21_X1 U278 ( .B1(n1627), .B2(n372), .A(n383), .ZN(n908) );
  NAND2_X1 U279 ( .A1(\mem[19][10] ), .A2(n1581), .ZN(n383) );
  OAI21_X1 U280 ( .B1(n1626), .B2(n372), .A(n384), .ZN(n909) );
  NAND2_X1 U281 ( .A1(\mem[19][11] ), .A2(n1581), .ZN(n384) );
  OAI21_X1 U282 ( .B1(n1625), .B2(n372), .A(n385), .ZN(n910) );
  NAND2_X1 U283 ( .A1(\mem[19][12] ), .A2(n1581), .ZN(n385) );
  OAI21_X1 U284 ( .B1(n1624), .B2(n372), .A(n386), .ZN(n911) );
  NAND2_X1 U285 ( .A1(\mem[19][13] ), .A2(n1581), .ZN(n386) );
  OAI21_X1 U286 ( .B1(n1623), .B2(n372), .A(n387), .ZN(n912) );
  NAND2_X1 U287 ( .A1(\mem[19][14] ), .A2(n1581), .ZN(n387) );
  OAI21_X1 U288 ( .B1(n1630), .B2(n457), .A(n465), .ZN(n985) );
  NAND2_X1 U289 ( .A1(\mem[24][7] ), .A2(n1576), .ZN(n465) );
  OAI21_X1 U290 ( .B1(n1561), .B2(n1576), .A(n466), .ZN(n986) );
  NAND2_X1 U291 ( .A1(\mem[24][8] ), .A2(n1576), .ZN(n466) );
  OAI21_X1 U292 ( .B1(n1628), .B2(n457), .A(n467), .ZN(n987) );
  NAND2_X1 U293 ( .A1(\mem[24][9] ), .A2(n1576), .ZN(n467) );
  OAI21_X1 U294 ( .B1(n1627), .B2(n457), .A(n468), .ZN(n988) );
  NAND2_X1 U295 ( .A1(\mem[24][10] ), .A2(n1576), .ZN(n468) );
  OAI21_X1 U296 ( .B1(n1626), .B2(n457), .A(n469), .ZN(n989) );
  NAND2_X1 U297 ( .A1(\mem[24][11] ), .A2(n1576), .ZN(n469) );
  OAI21_X1 U298 ( .B1(n1625), .B2(n457), .A(n470), .ZN(n990) );
  NAND2_X1 U299 ( .A1(\mem[24][12] ), .A2(n1576), .ZN(n470) );
  OAI21_X1 U300 ( .B1(n1624), .B2(n457), .A(n471), .ZN(n991) );
  NAND2_X1 U301 ( .A1(\mem[24][13] ), .A2(n1576), .ZN(n471) );
  OAI21_X1 U302 ( .B1(n1623), .B2(n457), .A(n472), .ZN(n992) );
  NAND2_X1 U303 ( .A1(\mem[24][14] ), .A2(n1576), .ZN(n472) );
  OAI21_X1 U304 ( .B1(n1630), .B2(n475), .A(n483), .ZN(n1001) );
  NAND2_X1 U305 ( .A1(\mem[25][7] ), .A2(n1575), .ZN(n483) );
  OAI21_X1 U306 ( .B1(n1561), .B2(n1575), .A(n484), .ZN(n1002) );
  NAND2_X1 U307 ( .A1(\mem[25][8] ), .A2(n1575), .ZN(n484) );
  OAI21_X1 U308 ( .B1(n1628), .B2(n475), .A(n485), .ZN(n1003) );
  NAND2_X1 U309 ( .A1(\mem[25][9] ), .A2(n1575), .ZN(n485) );
  OAI21_X1 U310 ( .B1(n1627), .B2(n475), .A(n486), .ZN(n1004) );
  NAND2_X1 U311 ( .A1(\mem[25][10] ), .A2(n1575), .ZN(n486) );
  OAI21_X1 U312 ( .B1(n1626), .B2(n475), .A(n487), .ZN(n1005) );
  NAND2_X1 U313 ( .A1(\mem[25][11] ), .A2(n1575), .ZN(n487) );
  OAI21_X1 U314 ( .B1(n1625), .B2(n475), .A(n488), .ZN(n1006) );
  NAND2_X1 U315 ( .A1(\mem[25][12] ), .A2(n1575), .ZN(n488) );
  OAI21_X1 U316 ( .B1(n1624), .B2(n475), .A(n489), .ZN(n1007) );
  NAND2_X1 U317 ( .A1(\mem[25][13] ), .A2(n1575), .ZN(n489) );
  OAI21_X1 U318 ( .B1(n1623), .B2(n475), .A(n490), .ZN(n1008) );
  NAND2_X1 U319 ( .A1(\mem[25][14] ), .A2(n1575), .ZN(n490) );
  OAI21_X1 U320 ( .B1(n1630), .B2(n492), .A(n500), .ZN(n1017) );
  NAND2_X1 U321 ( .A1(\mem[26][7] ), .A2(n1574), .ZN(n500) );
  OAI21_X1 U322 ( .B1(n1629), .B2(n1574), .A(n501), .ZN(n1018) );
  NAND2_X1 U323 ( .A1(\mem[26][8] ), .A2(n1574), .ZN(n501) );
  OAI21_X1 U324 ( .B1(n1628), .B2(n492), .A(n502), .ZN(n1019) );
  NAND2_X1 U325 ( .A1(\mem[26][9] ), .A2(n1574), .ZN(n502) );
  OAI21_X1 U326 ( .B1(n1627), .B2(n492), .A(n503), .ZN(n1020) );
  NAND2_X1 U327 ( .A1(\mem[26][10] ), .A2(n1574), .ZN(n503) );
  OAI21_X1 U328 ( .B1(n1626), .B2(n492), .A(n504), .ZN(n1021) );
  NAND2_X1 U329 ( .A1(\mem[26][11] ), .A2(n1574), .ZN(n504) );
  OAI21_X1 U330 ( .B1(n1625), .B2(n492), .A(n505), .ZN(n1022) );
  NAND2_X1 U331 ( .A1(\mem[26][12] ), .A2(n1574), .ZN(n505) );
  OAI21_X1 U332 ( .B1(n1624), .B2(n492), .A(n506), .ZN(n1023) );
  NAND2_X1 U333 ( .A1(\mem[26][13] ), .A2(n1574), .ZN(n506) );
  OAI21_X1 U334 ( .B1(n1623), .B2(n492), .A(n507), .ZN(n1024) );
  NAND2_X1 U335 ( .A1(\mem[26][14] ), .A2(n1574), .ZN(n507) );
  OAI21_X1 U336 ( .B1(n1630), .B2(n509), .A(n517), .ZN(n1033) );
  NAND2_X1 U337 ( .A1(\mem[27][7] ), .A2(n509), .ZN(n517) );
  OAI21_X1 U338 ( .B1(n1629), .B2(n1573), .A(n518), .ZN(n1034) );
  NAND2_X1 U339 ( .A1(\mem[27][8] ), .A2(n1573), .ZN(n518) );
  OAI21_X1 U340 ( .B1(n1628), .B2(n509), .A(n519), .ZN(n1035) );
  NAND2_X1 U341 ( .A1(\mem[27][9] ), .A2(n1573), .ZN(n519) );
  OAI21_X1 U342 ( .B1(n1627), .B2(n509), .A(n520), .ZN(n1036) );
  NAND2_X1 U343 ( .A1(\mem[27][10] ), .A2(n1573), .ZN(n520) );
  OAI21_X1 U344 ( .B1(n1626), .B2(n509), .A(n521), .ZN(n1037) );
  NAND2_X1 U345 ( .A1(\mem[27][11] ), .A2(n1573), .ZN(n521) );
  OAI21_X1 U346 ( .B1(n1625), .B2(n509), .A(n522), .ZN(n1038) );
  NAND2_X1 U347 ( .A1(\mem[27][12] ), .A2(n1573), .ZN(n522) );
  OAI21_X1 U348 ( .B1(n1624), .B2(n509), .A(n523), .ZN(n1039) );
  NAND2_X1 U349 ( .A1(\mem[27][13] ), .A2(n1573), .ZN(n523) );
  OAI21_X1 U350 ( .B1(n1623), .B2(n509), .A(n524), .ZN(n1040) );
  NAND2_X1 U351 ( .A1(\mem[27][14] ), .A2(n1573), .ZN(n524) );
  OAI21_X1 U352 ( .B1(n1562), .B2(n111), .A(n119), .ZN(n665) );
  NAND2_X1 U353 ( .A1(\mem[4][7] ), .A2(n1596), .ZN(n119) );
  OAI21_X1 U354 ( .B1(n1629), .B2(n1596), .A(n120), .ZN(n666) );
  NAND2_X1 U355 ( .A1(\mem[4][8] ), .A2(n1596), .ZN(n120) );
  OAI21_X1 U356 ( .B1(n1560), .B2(n111), .A(n121), .ZN(n667) );
  NAND2_X1 U357 ( .A1(\mem[4][9] ), .A2(n1596), .ZN(n121) );
  OAI21_X1 U358 ( .B1(n1559), .B2(n111), .A(n122), .ZN(n668) );
  NAND2_X1 U359 ( .A1(\mem[4][10] ), .A2(n1596), .ZN(n122) );
  OAI21_X1 U360 ( .B1(n1558), .B2(n111), .A(n123), .ZN(n669) );
  NAND2_X1 U361 ( .A1(\mem[4][11] ), .A2(n1596), .ZN(n123) );
  OAI21_X1 U362 ( .B1(n1557), .B2(n111), .A(n124), .ZN(n670) );
  NAND2_X1 U363 ( .A1(\mem[4][12] ), .A2(n1596), .ZN(n124) );
  OAI21_X1 U364 ( .B1(n1556), .B2(n111), .A(n125), .ZN(n671) );
  NAND2_X1 U365 ( .A1(\mem[4][13] ), .A2(n1596), .ZN(n125) );
  OAI21_X1 U366 ( .B1(n1555), .B2(n111), .A(n126), .ZN(n672) );
  NAND2_X1 U367 ( .A1(\mem[4][14] ), .A2(n1596), .ZN(n126) );
  OAI21_X1 U368 ( .B1(n1562), .B2(n129), .A(n137), .ZN(n681) );
  NAND2_X1 U369 ( .A1(\mem[5][7] ), .A2(n1595), .ZN(n137) );
  OAI21_X1 U370 ( .B1(n1629), .B2(n129), .A(n138), .ZN(n682) );
  NAND2_X1 U371 ( .A1(\mem[5][8] ), .A2(n1595), .ZN(n138) );
  OAI21_X1 U372 ( .B1(n1560), .B2(n129), .A(n139), .ZN(n683) );
  NAND2_X1 U373 ( .A1(\mem[5][9] ), .A2(n129), .ZN(n139) );
  OAI21_X1 U374 ( .B1(n1559), .B2(n129), .A(n140), .ZN(n684) );
  NAND2_X1 U375 ( .A1(\mem[5][10] ), .A2(n129), .ZN(n140) );
  OAI21_X1 U376 ( .B1(n1558), .B2(n129), .A(n141), .ZN(n685) );
  NAND2_X1 U377 ( .A1(\mem[5][11] ), .A2(n129), .ZN(n141) );
  OAI21_X1 U378 ( .B1(n1557), .B2(n129), .A(n142), .ZN(n686) );
  NAND2_X1 U379 ( .A1(\mem[5][12] ), .A2(n1595), .ZN(n142) );
  OAI21_X1 U380 ( .B1(n1556), .B2(n129), .A(n143), .ZN(n687) );
  NAND2_X1 U381 ( .A1(\mem[5][13] ), .A2(n129), .ZN(n143) );
  OAI21_X1 U382 ( .B1(n1555), .B2(n129), .A(n144), .ZN(n688) );
  NAND2_X1 U383 ( .A1(\mem[5][14] ), .A2(n129), .ZN(n144) );
  OAI21_X1 U384 ( .B1(n1562), .B2(n1594), .A(n155), .ZN(n697) );
  NAND2_X1 U385 ( .A1(\mem[6][7] ), .A2(n1594), .ZN(n155) );
  OAI21_X1 U386 ( .B1(n1629), .B2(n1594), .A(n156), .ZN(n698) );
  NAND2_X1 U387 ( .A1(\mem[6][8] ), .A2(n147), .ZN(n156) );
  OAI21_X1 U388 ( .B1(n1560), .B2(n1594), .A(n157), .ZN(n699) );
  NAND2_X1 U389 ( .A1(\mem[6][9] ), .A2(n147), .ZN(n157) );
  OAI21_X1 U390 ( .B1(n1559), .B2(n1594), .A(n158), .ZN(n700) );
  NAND2_X1 U391 ( .A1(\mem[6][10] ), .A2(n147), .ZN(n158) );
  OAI21_X1 U392 ( .B1(n1558), .B2(n1594), .A(n159), .ZN(n701) );
  NAND2_X1 U393 ( .A1(\mem[6][11] ), .A2(n147), .ZN(n159) );
  OAI21_X1 U394 ( .B1(n1557), .B2(n1594), .A(n160), .ZN(n702) );
  NAND2_X1 U395 ( .A1(\mem[6][12] ), .A2(n147), .ZN(n160) );
  OAI21_X1 U396 ( .B1(n1556), .B2(n1594), .A(n161), .ZN(n703) );
  NAND2_X1 U397 ( .A1(\mem[6][13] ), .A2(n147), .ZN(n161) );
  OAI21_X1 U398 ( .B1(n1555), .B2(n1594), .A(n162), .ZN(n704) );
  NAND2_X1 U399 ( .A1(\mem[6][14] ), .A2(n147), .ZN(n162) );
  OAI21_X1 U400 ( .B1(n1562), .B2(n165), .A(n173), .ZN(n713) );
  NAND2_X1 U401 ( .A1(\mem[7][7] ), .A2(n1593), .ZN(n173) );
  OAI21_X1 U402 ( .B1(n1629), .B2(n1593), .A(n174), .ZN(n714) );
  NAND2_X1 U403 ( .A1(\mem[7][8] ), .A2(n1593), .ZN(n174) );
  OAI21_X1 U404 ( .B1(n1560), .B2(n165), .A(n175), .ZN(n715) );
  NAND2_X1 U405 ( .A1(\mem[7][9] ), .A2(n1593), .ZN(n175) );
  OAI21_X1 U406 ( .B1(n1559), .B2(n165), .A(n176), .ZN(n716) );
  NAND2_X1 U407 ( .A1(\mem[7][10] ), .A2(n1593), .ZN(n176) );
  OAI21_X1 U408 ( .B1(n1558), .B2(n165), .A(n177), .ZN(n717) );
  NAND2_X1 U409 ( .A1(\mem[7][11] ), .A2(n1593), .ZN(n177) );
  OAI21_X1 U410 ( .B1(n1557), .B2(n165), .A(n178), .ZN(n718) );
  NAND2_X1 U411 ( .A1(\mem[7][12] ), .A2(n1593), .ZN(n178) );
  OAI21_X1 U412 ( .B1(n1556), .B2(n165), .A(n179), .ZN(n719) );
  NAND2_X1 U413 ( .A1(\mem[7][13] ), .A2(n1593), .ZN(n179) );
  OAI21_X1 U414 ( .B1(n1555), .B2(n165), .A(n180), .ZN(n720) );
  NAND2_X1 U415 ( .A1(\mem[7][14] ), .A2(n1593), .ZN(n180) );
  OAI21_X1 U416 ( .B1(n1562), .B2(n252), .A(n260), .ZN(n793) );
  NAND2_X1 U417 ( .A1(\mem[12][7] ), .A2(n1588), .ZN(n260) );
  OAI21_X1 U418 ( .B1(n1629), .B2(n1588), .A(n261), .ZN(n794) );
  NAND2_X1 U419 ( .A1(\mem[12][8] ), .A2(n1588), .ZN(n261) );
  OAI21_X1 U420 ( .B1(n1560), .B2(n252), .A(n262), .ZN(n795) );
  NAND2_X1 U421 ( .A1(\mem[12][9] ), .A2(n1588), .ZN(n262) );
  OAI21_X1 U422 ( .B1(n1559), .B2(n252), .A(n263), .ZN(n796) );
  NAND2_X1 U423 ( .A1(\mem[12][10] ), .A2(n1588), .ZN(n263) );
  OAI21_X1 U424 ( .B1(n1558), .B2(n252), .A(n264), .ZN(n797) );
  NAND2_X1 U425 ( .A1(\mem[12][11] ), .A2(n1588), .ZN(n264) );
  OAI21_X1 U426 ( .B1(n1557), .B2(n252), .A(n265), .ZN(n798) );
  NAND2_X1 U427 ( .A1(\mem[12][12] ), .A2(n1588), .ZN(n265) );
  OAI21_X1 U428 ( .B1(n1556), .B2(n252), .A(n266), .ZN(n799) );
  NAND2_X1 U429 ( .A1(\mem[12][13] ), .A2(n1588), .ZN(n266) );
  OAI21_X1 U430 ( .B1(n1555), .B2(n252), .A(n267), .ZN(n800) );
  NAND2_X1 U431 ( .A1(\mem[12][14] ), .A2(n1588), .ZN(n267) );
  OAI21_X1 U432 ( .B1(n1630), .B2(n269), .A(n277), .ZN(n809) );
  NAND2_X1 U433 ( .A1(\mem[13][7] ), .A2(n1587), .ZN(n277) );
  OAI21_X1 U434 ( .B1(n1561), .B2(n1587), .A(n278), .ZN(n810) );
  NAND2_X1 U435 ( .A1(\mem[13][8] ), .A2(n1587), .ZN(n278) );
  OAI21_X1 U436 ( .B1(n1628), .B2(n269), .A(n279), .ZN(n811) );
  NAND2_X1 U437 ( .A1(\mem[13][9] ), .A2(n1587), .ZN(n279) );
  OAI21_X1 U438 ( .B1(n1627), .B2(n269), .A(n280), .ZN(n812) );
  NAND2_X1 U439 ( .A1(\mem[13][10] ), .A2(n1587), .ZN(n280) );
  OAI21_X1 U440 ( .B1(n1626), .B2(n269), .A(n281), .ZN(n813) );
  NAND2_X1 U441 ( .A1(\mem[13][11] ), .A2(n1587), .ZN(n281) );
  OAI21_X1 U442 ( .B1(n1625), .B2(n269), .A(n282), .ZN(n814) );
  NAND2_X1 U443 ( .A1(\mem[13][12] ), .A2(n1587), .ZN(n282) );
  OAI21_X1 U444 ( .B1(n1624), .B2(n269), .A(n283), .ZN(n815) );
  NAND2_X1 U445 ( .A1(\mem[13][13] ), .A2(n1587), .ZN(n283) );
  OAI21_X1 U446 ( .B1(n1623), .B2(n269), .A(n284), .ZN(n816) );
  NAND2_X1 U447 ( .A1(\mem[13][14] ), .A2(n1587), .ZN(n284) );
  OAI21_X1 U448 ( .B1(n1630), .B2(n1586), .A(n294), .ZN(n825) );
  NAND2_X1 U449 ( .A1(\mem[14][7] ), .A2(n1586), .ZN(n294) );
  OAI21_X1 U450 ( .B1(n1561), .B2(n286), .A(n295), .ZN(n826) );
  NAND2_X1 U451 ( .A1(\mem[14][8] ), .A2(n1586), .ZN(n295) );
  OAI21_X1 U452 ( .B1(n1628), .B2(n286), .A(n296), .ZN(n827) );
  NAND2_X1 U453 ( .A1(\mem[14][9] ), .A2(n1586), .ZN(n296) );
  OAI21_X1 U454 ( .B1(n1627), .B2(n286), .A(n297), .ZN(n828) );
  NAND2_X1 U455 ( .A1(\mem[14][10] ), .A2(n1586), .ZN(n297) );
  OAI21_X1 U456 ( .B1(n1626), .B2(n286), .A(n298), .ZN(n829) );
  NAND2_X1 U457 ( .A1(\mem[14][11] ), .A2(n1586), .ZN(n298) );
  OAI21_X1 U458 ( .B1(n1625), .B2(n286), .A(n299), .ZN(n830) );
  NAND2_X1 U459 ( .A1(\mem[14][12] ), .A2(n1586), .ZN(n299) );
  OAI21_X1 U460 ( .B1(n1624), .B2(n286), .A(n300), .ZN(n831) );
  NAND2_X1 U461 ( .A1(\mem[14][13] ), .A2(n1586), .ZN(n300) );
  OAI21_X1 U462 ( .B1(n1623), .B2(n286), .A(n301), .ZN(n832) );
  NAND2_X1 U463 ( .A1(\mem[14][14] ), .A2(n1586), .ZN(n301) );
  OAI21_X1 U464 ( .B1(n1630), .B2(n303), .A(n311), .ZN(n841) );
  NAND2_X1 U465 ( .A1(\mem[15][7] ), .A2(n1585), .ZN(n311) );
  OAI21_X1 U466 ( .B1(n1561), .B2(n1585), .A(n312), .ZN(n842) );
  NAND2_X1 U467 ( .A1(\mem[15][8] ), .A2(n1585), .ZN(n312) );
  OAI21_X1 U468 ( .B1(n1628), .B2(n303), .A(n313), .ZN(n843) );
  NAND2_X1 U469 ( .A1(\mem[15][9] ), .A2(n1585), .ZN(n313) );
  OAI21_X1 U470 ( .B1(n1627), .B2(n303), .A(n314), .ZN(n844) );
  NAND2_X1 U471 ( .A1(\mem[15][10] ), .A2(n1585), .ZN(n314) );
  OAI21_X1 U472 ( .B1(n1626), .B2(n303), .A(n315), .ZN(n845) );
  NAND2_X1 U473 ( .A1(\mem[15][11] ), .A2(n1585), .ZN(n315) );
  OAI21_X1 U474 ( .B1(n1625), .B2(n303), .A(n316), .ZN(n846) );
  NAND2_X1 U475 ( .A1(\mem[15][12] ), .A2(n1585), .ZN(n316) );
  OAI21_X1 U476 ( .B1(n1624), .B2(n303), .A(n317), .ZN(n847) );
  NAND2_X1 U477 ( .A1(\mem[15][13] ), .A2(n1585), .ZN(n317) );
  OAI21_X1 U478 ( .B1(n1623), .B2(n303), .A(n318), .ZN(n848) );
  NAND2_X1 U479 ( .A1(\mem[15][14] ), .A2(n1585), .ZN(n318) );
  OAI21_X1 U480 ( .B1(n1630), .B2(n389), .A(n397), .ZN(n921) );
  NAND2_X1 U481 ( .A1(\mem[20][7] ), .A2(n1580), .ZN(n397) );
  OAI21_X1 U482 ( .B1(n1561), .B2(n1580), .A(n398), .ZN(n922) );
  NAND2_X1 U483 ( .A1(\mem[20][8] ), .A2(n1580), .ZN(n398) );
  OAI21_X1 U484 ( .B1(n1628), .B2(n389), .A(n399), .ZN(n923) );
  NAND2_X1 U485 ( .A1(\mem[20][9] ), .A2(n1580), .ZN(n399) );
  OAI21_X1 U486 ( .B1(n1627), .B2(n389), .A(n400), .ZN(n924) );
  NAND2_X1 U487 ( .A1(\mem[20][10] ), .A2(n1580), .ZN(n400) );
  OAI21_X1 U488 ( .B1(n1626), .B2(n389), .A(n401), .ZN(n925) );
  NAND2_X1 U489 ( .A1(\mem[20][11] ), .A2(n1580), .ZN(n401) );
  OAI21_X1 U490 ( .B1(n1625), .B2(n389), .A(n402), .ZN(n926) );
  NAND2_X1 U491 ( .A1(\mem[20][12] ), .A2(n1580), .ZN(n402) );
  OAI21_X1 U492 ( .B1(n1624), .B2(n389), .A(n403), .ZN(n927) );
  NAND2_X1 U493 ( .A1(\mem[20][13] ), .A2(n1580), .ZN(n403) );
  OAI21_X1 U494 ( .B1(n1623), .B2(n389), .A(n404), .ZN(n928) );
  NAND2_X1 U495 ( .A1(\mem[20][14] ), .A2(n1580), .ZN(n404) );
  OAI21_X1 U496 ( .B1(n1630), .B2(n406), .A(n414), .ZN(n937) );
  NAND2_X1 U497 ( .A1(\mem[21][7] ), .A2(n1579), .ZN(n414) );
  OAI21_X1 U498 ( .B1(n1561), .B2(n1579), .A(n415), .ZN(n938) );
  NAND2_X1 U499 ( .A1(\mem[21][8] ), .A2(n1579), .ZN(n415) );
  OAI21_X1 U500 ( .B1(n1628), .B2(n406), .A(n416), .ZN(n939) );
  NAND2_X1 U501 ( .A1(\mem[21][9] ), .A2(n1579), .ZN(n416) );
  OAI21_X1 U502 ( .B1(n1627), .B2(n406), .A(n417), .ZN(n940) );
  NAND2_X1 U503 ( .A1(\mem[21][10] ), .A2(n1579), .ZN(n417) );
  OAI21_X1 U504 ( .B1(n1626), .B2(n406), .A(n418), .ZN(n941) );
  NAND2_X1 U505 ( .A1(\mem[21][11] ), .A2(n1579), .ZN(n418) );
  OAI21_X1 U506 ( .B1(n1625), .B2(n406), .A(n419), .ZN(n942) );
  NAND2_X1 U507 ( .A1(\mem[21][12] ), .A2(n1579), .ZN(n419) );
  OAI21_X1 U508 ( .B1(n1624), .B2(n406), .A(n420), .ZN(n943) );
  NAND2_X1 U509 ( .A1(\mem[21][13] ), .A2(n1579), .ZN(n420) );
  OAI21_X1 U510 ( .B1(n1623), .B2(n406), .A(n421), .ZN(n944) );
  NAND2_X1 U511 ( .A1(\mem[21][14] ), .A2(n1579), .ZN(n421) );
  OAI21_X1 U512 ( .B1(n1630), .B2(n423), .A(n431), .ZN(n953) );
  NAND2_X1 U513 ( .A1(\mem[22][7] ), .A2(n1578), .ZN(n431) );
  OAI21_X1 U514 ( .B1(n1561), .B2(n423), .A(n432), .ZN(n954) );
  NAND2_X1 U515 ( .A1(\mem[22][8] ), .A2(n1578), .ZN(n432) );
  OAI21_X1 U516 ( .B1(n1628), .B2(n423), .A(n433), .ZN(n955) );
  NAND2_X1 U517 ( .A1(\mem[22][9] ), .A2(n423), .ZN(n433) );
  OAI21_X1 U518 ( .B1(n1627), .B2(n423), .A(n434), .ZN(n956) );
  NAND2_X1 U519 ( .A1(\mem[22][10] ), .A2(n423), .ZN(n434) );
  OAI21_X1 U520 ( .B1(n1626), .B2(n423), .A(n435), .ZN(n957) );
  NAND2_X1 U521 ( .A1(\mem[22][11] ), .A2(n423), .ZN(n435) );
  OAI21_X1 U522 ( .B1(n1625), .B2(n423), .A(n436), .ZN(n958) );
  NAND2_X1 U523 ( .A1(\mem[22][12] ), .A2(n1578), .ZN(n436) );
  OAI21_X1 U524 ( .B1(n1624), .B2(n423), .A(n437), .ZN(n959) );
  NAND2_X1 U525 ( .A1(\mem[22][13] ), .A2(n423), .ZN(n437) );
  OAI21_X1 U526 ( .B1(n1623), .B2(n423), .A(n438), .ZN(n960) );
  NAND2_X1 U527 ( .A1(\mem[22][14] ), .A2(n423), .ZN(n438) );
  OAI21_X1 U528 ( .B1(n1630), .B2(n440), .A(n448), .ZN(n969) );
  NAND2_X1 U529 ( .A1(\mem[23][7] ), .A2(n1577), .ZN(n448) );
  OAI21_X1 U530 ( .B1(n1561), .B2(n1577), .A(n449), .ZN(n970) );
  NAND2_X1 U531 ( .A1(\mem[23][8] ), .A2(n1577), .ZN(n449) );
  OAI21_X1 U532 ( .B1(n1628), .B2(n440), .A(n450), .ZN(n971) );
  NAND2_X1 U533 ( .A1(\mem[23][9] ), .A2(n1577), .ZN(n450) );
  OAI21_X1 U534 ( .B1(n1627), .B2(n440), .A(n451), .ZN(n972) );
  NAND2_X1 U535 ( .A1(\mem[23][10] ), .A2(n1577), .ZN(n451) );
  OAI21_X1 U536 ( .B1(n1626), .B2(n440), .A(n452), .ZN(n973) );
  NAND2_X1 U537 ( .A1(\mem[23][11] ), .A2(n1577), .ZN(n452) );
  OAI21_X1 U538 ( .B1(n1625), .B2(n440), .A(n453), .ZN(n974) );
  NAND2_X1 U539 ( .A1(\mem[23][12] ), .A2(n1577), .ZN(n453) );
  OAI21_X1 U540 ( .B1(n1624), .B2(n440), .A(n454), .ZN(n975) );
  NAND2_X1 U541 ( .A1(\mem[23][13] ), .A2(n1577), .ZN(n454) );
  OAI21_X1 U542 ( .B1(n1623), .B2(n440), .A(n455), .ZN(n976) );
  NAND2_X1 U543 ( .A1(\mem[23][14] ), .A2(n1577), .ZN(n455) );
  OAI21_X1 U544 ( .B1(n1630), .B2(n1572), .A(n534), .ZN(n1049) );
  NAND2_X1 U545 ( .A1(\mem[28][7] ), .A2(n1572), .ZN(n534) );
  OAI21_X1 U546 ( .B1(n1629), .B2(n1572), .A(n535), .ZN(n1050) );
  NAND2_X1 U547 ( .A1(\mem[28][8] ), .A2(n526), .ZN(n535) );
  OAI21_X1 U548 ( .B1(n1628), .B2(n1572), .A(n536), .ZN(n1051) );
  NAND2_X1 U549 ( .A1(\mem[28][9] ), .A2(n526), .ZN(n536) );
  OAI21_X1 U550 ( .B1(n1627), .B2(n1572), .A(n537), .ZN(n1052) );
  NAND2_X1 U551 ( .A1(\mem[28][10] ), .A2(n526), .ZN(n537) );
  OAI21_X1 U552 ( .B1(n1626), .B2(n1572), .A(n538), .ZN(n1053) );
  NAND2_X1 U553 ( .A1(\mem[28][11] ), .A2(n526), .ZN(n538) );
  OAI21_X1 U554 ( .B1(n1625), .B2(n1572), .A(n539), .ZN(n1054) );
  NAND2_X1 U555 ( .A1(\mem[28][12] ), .A2(n526), .ZN(n539) );
  OAI21_X1 U556 ( .B1(n1624), .B2(n1572), .A(n540), .ZN(n1055) );
  NAND2_X1 U557 ( .A1(\mem[28][13] ), .A2(n526), .ZN(n540) );
  OAI21_X1 U558 ( .B1(n1623), .B2(n1572), .A(n541), .ZN(n1056) );
  NAND2_X1 U559 ( .A1(\mem[28][14] ), .A2(n526), .ZN(n541) );
  OAI21_X1 U560 ( .B1(n1630), .B2(n543), .A(n551), .ZN(n1065) );
  NAND2_X1 U561 ( .A1(\mem[29][7] ), .A2(n1571), .ZN(n551) );
  OAI21_X1 U562 ( .B1(n1629), .B2(n1571), .A(n552), .ZN(n1066) );
  NAND2_X1 U563 ( .A1(\mem[29][8] ), .A2(n1571), .ZN(n552) );
  OAI21_X1 U564 ( .B1(n1628), .B2(n543), .A(n553), .ZN(n1067) );
  NAND2_X1 U565 ( .A1(\mem[29][9] ), .A2(n1571), .ZN(n553) );
  OAI21_X1 U566 ( .B1(n1627), .B2(n543), .A(n554), .ZN(n1068) );
  NAND2_X1 U567 ( .A1(\mem[29][10] ), .A2(n1571), .ZN(n554) );
  OAI21_X1 U568 ( .B1(n1626), .B2(n543), .A(n555), .ZN(n1069) );
  NAND2_X1 U569 ( .A1(\mem[29][11] ), .A2(n1571), .ZN(n555) );
  OAI21_X1 U570 ( .B1(n1625), .B2(n543), .A(n556), .ZN(n1070) );
  NAND2_X1 U571 ( .A1(\mem[29][12] ), .A2(n1571), .ZN(n556) );
  OAI21_X1 U572 ( .B1(n1624), .B2(n543), .A(n557), .ZN(n1071) );
  NAND2_X1 U573 ( .A1(\mem[29][13] ), .A2(n1571), .ZN(n557) );
  OAI21_X1 U574 ( .B1(n1623), .B2(n543), .A(n558), .ZN(n1072) );
  NAND2_X1 U575 ( .A1(\mem[29][14] ), .A2(n1571), .ZN(n558) );
  OAI21_X1 U576 ( .B1(n1630), .B2(n560), .A(n568), .ZN(n1081) );
  NAND2_X1 U577 ( .A1(\mem[30][7] ), .A2(n560), .ZN(n568) );
  OAI21_X1 U578 ( .B1(n1629), .B2(n1570), .A(n569), .ZN(n1082) );
  NAND2_X1 U579 ( .A1(\mem[30][8] ), .A2(n1570), .ZN(n569) );
  OAI21_X1 U580 ( .B1(n1628), .B2(n560), .A(n570), .ZN(n1083) );
  NAND2_X1 U581 ( .A1(\mem[30][9] ), .A2(n1570), .ZN(n570) );
  OAI21_X1 U582 ( .B1(n1627), .B2(n560), .A(n571), .ZN(n1084) );
  NAND2_X1 U583 ( .A1(\mem[30][10] ), .A2(n1570), .ZN(n571) );
  OAI21_X1 U584 ( .B1(n1626), .B2(n560), .A(n572), .ZN(n1085) );
  NAND2_X1 U585 ( .A1(\mem[30][11] ), .A2(n1570), .ZN(n572) );
  OAI21_X1 U586 ( .B1(n1625), .B2(n560), .A(n573), .ZN(n1086) );
  NAND2_X1 U587 ( .A1(\mem[30][12] ), .A2(n1570), .ZN(n573) );
  OAI21_X1 U588 ( .B1(n1624), .B2(n560), .A(n574), .ZN(n1087) );
  NAND2_X1 U589 ( .A1(\mem[30][13] ), .A2(n1570), .ZN(n574) );
  OAI21_X1 U590 ( .B1(n1623), .B2(n560), .A(n575), .ZN(n1088) );
  NAND2_X1 U591 ( .A1(\mem[30][14] ), .A2(n1570), .ZN(n575) );
  OAI21_X1 U592 ( .B1(n38), .B2(n1629), .A(n47), .ZN(n602) );
  NAND2_X1 U593 ( .A1(\mem[0][8] ), .A2(n1600), .ZN(n47) );
  OAI21_X1 U594 ( .B1(n38), .B2(n1560), .A(n48), .ZN(n603) );
  NAND2_X1 U595 ( .A1(\mem[0][9] ), .A2(n38), .ZN(n48) );
  OAI21_X1 U596 ( .B1(n1600), .B2(n1559), .A(n49), .ZN(n604) );
  NAND2_X1 U597 ( .A1(\mem[0][10] ), .A2(n38), .ZN(n49) );
  OAI21_X1 U598 ( .B1(n38), .B2(n1558), .A(n50), .ZN(n605) );
  NAND2_X1 U599 ( .A1(\mem[0][11] ), .A2(n38), .ZN(n50) );
  OAI21_X1 U600 ( .B1(n38), .B2(n1557), .A(n51), .ZN(n606) );
  NAND2_X1 U601 ( .A1(\mem[0][12] ), .A2(n38), .ZN(n51) );
  OAI21_X1 U602 ( .B1(n38), .B2(n1556), .A(n52), .ZN(n607) );
  NAND2_X1 U603 ( .A1(\mem[0][13] ), .A2(n38), .ZN(n52) );
  OAI21_X1 U604 ( .B1(n38), .B2(n1555), .A(n53), .ZN(n608) );
  NAND2_X1 U605 ( .A1(\mem[0][14] ), .A2(n38), .ZN(n53) );
  OAI21_X1 U606 ( .B1(n1637), .B2(n492), .A(n493), .ZN(n1010) );
  NAND2_X1 U607 ( .A1(\mem[26][0] ), .A2(n1574), .ZN(n493) );
  OAI21_X1 U608 ( .B1(n1636), .B2(n492), .A(n494), .ZN(n1011) );
  NAND2_X1 U609 ( .A1(\mem[26][1] ), .A2(n1574), .ZN(n494) );
  OAI21_X1 U610 ( .B1(n1635), .B2(n492), .A(n495), .ZN(n1012) );
  NAND2_X1 U611 ( .A1(\mem[26][2] ), .A2(n1574), .ZN(n495) );
  OAI21_X1 U612 ( .B1(n1634), .B2(n492), .A(n496), .ZN(n1013) );
  NAND2_X1 U613 ( .A1(\mem[26][3] ), .A2(n1574), .ZN(n496) );
  OAI21_X1 U614 ( .B1(n1633), .B2(n492), .A(n497), .ZN(n1014) );
  NAND2_X1 U615 ( .A1(\mem[26][4] ), .A2(n492), .ZN(n497) );
  OAI21_X1 U616 ( .B1(n1632), .B2(n492), .A(n498), .ZN(n1015) );
  NAND2_X1 U617 ( .A1(\mem[26][5] ), .A2(n492), .ZN(n498) );
  OAI21_X1 U618 ( .B1(n1631), .B2(n492), .A(n499), .ZN(n1016) );
  NAND2_X1 U619 ( .A1(\mem[26][6] ), .A2(n492), .ZN(n499) );
  OAI21_X1 U620 ( .B1(n1622), .B2(n492), .A(n508), .ZN(n1025) );
  NAND2_X1 U621 ( .A1(\mem[26][15] ), .A2(n1574), .ZN(n508) );
  OAI21_X1 U622 ( .B1(n1637), .B2(n509), .A(n510), .ZN(n1026) );
  NAND2_X1 U623 ( .A1(\mem[27][0] ), .A2(n1573), .ZN(n510) );
  OAI21_X1 U624 ( .B1(n1636), .B2(n509), .A(n511), .ZN(n1027) );
  NAND2_X1 U625 ( .A1(\mem[27][1] ), .A2(n1573), .ZN(n511) );
  OAI21_X1 U626 ( .B1(n1635), .B2(n509), .A(n512), .ZN(n1028) );
  NAND2_X1 U627 ( .A1(\mem[27][2] ), .A2(n1573), .ZN(n512) );
  OAI21_X1 U628 ( .B1(n1634), .B2(n509), .A(n513), .ZN(n1029) );
  NAND2_X1 U629 ( .A1(\mem[27][3] ), .A2(n1573), .ZN(n513) );
  OAI21_X1 U630 ( .B1(n1633), .B2(n509), .A(n514), .ZN(n1030) );
  NAND2_X1 U631 ( .A1(\mem[27][4] ), .A2(n1573), .ZN(n514) );
  OAI21_X1 U632 ( .B1(n1632), .B2(n509), .A(n515), .ZN(n1031) );
  NAND2_X1 U633 ( .A1(\mem[27][5] ), .A2(n509), .ZN(n515) );
  OAI21_X1 U634 ( .B1(n1631), .B2(n509), .A(n516), .ZN(n1032) );
  NAND2_X1 U635 ( .A1(\mem[27][6] ), .A2(n509), .ZN(n516) );
  OAI21_X1 U636 ( .B1(n1622), .B2(n509), .A(n525), .ZN(n1041) );
  NAND2_X1 U637 ( .A1(\mem[27][15] ), .A2(n1573), .ZN(n525) );
  OAI21_X1 U638 ( .B1(n1637), .B2(n1572), .A(n527), .ZN(n1042) );
  NAND2_X1 U639 ( .A1(\mem[28][0] ), .A2(n1572), .ZN(n527) );
  OAI21_X1 U640 ( .B1(n1636), .B2(n526), .A(n528), .ZN(n1043) );
  NAND2_X1 U641 ( .A1(\mem[28][1] ), .A2(n526), .ZN(n528) );
  OAI21_X1 U642 ( .B1(n1635), .B2(n526), .A(n529), .ZN(n1044) );
  NAND2_X1 U643 ( .A1(\mem[28][2] ), .A2(n526), .ZN(n529) );
  OAI21_X1 U644 ( .B1(n1634), .B2(n526), .A(n530), .ZN(n1045) );
  NAND2_X1 U645 ( .A1(\mem[28][3] ), .A2(n526), .ZN(n530) );
  OAI21_X1 U646 ( .B1(n1633), .B2(n526), .A(n531), .ZN(n1046) );
  NAND2_X1 U647 ( .A1(\mem[28][4] ), .A2(n1572), .ZN(n531) );
  OAI21_X1 U648 ( .B1(n1632), .B2(n526), .A(n532), .ZN(n1047) );
  NAND2_X1 U649 ( .A1(\mem[28][5] ), .A2(n1572), .ZN(n532) );
  OAI21_X1 U650 ( .B1(n1631), .B2(n526), .A(n533), .ZN(n1048) );
  NAND2_X1 U651 ( .A1(\mem[28][6] ), .A2(n1572), .ZN(n533) );
  OAI21_X1 U652 ( .B1(n1622), .B2(n526), .A(n542), .ZN(n1057) );
  NAND2_X1 U653 ( .A1(\mem[28][15] ), .A2(n526), .ZN(n542) );
  OAI21_X1 U654 ( .B1(n1637), .B2(n543), .A(n544), .ZN(n1058) );
  NAND2_X1 U655 ( .A1(\mem[29][0] ), .A2(n1571), .ZN(n544) );
  OAI21_X1 U656 ( .B1(n1636), .B2(n543), .A(n545), .ZN(n1059) );
  NAND2_X1 U657 ( .A1(\mem[29][1] ), .A2(n1571), .ZN(n545) );
  OAI21_X1 U658 ( .B1(n1635), .B2(n543), .A(n546), .ZN(n1060) );
  NAND2_X1 U659 ( .A1(\mem[29][2] ), .A2(n1571), .ZN(n546) );
  OAI21_X1 U660 ( .B1(n1634), .B2(n543), .A(n547), .ZN(n1061) );
  NAND2_X1 U661 ( .A1(\mem[29][3] ), .A2(n1571), .ZN(n547) );
  OAI21_X1 U662 ( .B1(n1633), .B2(n543), .A(n548), .ZN(n1062) );
  NAND2_X1 U663 ( .A1(\mem[29][4] ), .A2(n543), .ZN(n548) );
  OAI21_X1 U664 ( .B1(n1632), .B2(n543), .A(n549), .ZN(n1063) );
  NAND2_X1 U665 ( .A1(\mem[29][5] ), .A2(n543), .ZN(n549) );
  OAI21_X1 U666 ( .B1(n1631), .B2(n543), .A(n550), .ZN(n1064) );
  NAND2_X1 U667 ( .A1(\mem[29][6] ), .A2(n543), .ZN(n550) );
  OAI21_X1 U668 ( .B1(n1622), .B2(n543), .A(n559), .ZN(n1073) );
  NAND2_X1 U669 ( .A1(\mem[29][15] ), .A2(n1571), .ZN(n559) );
  OAI21_X1 U670 ( .B1(n1637), .B2(n560), .A(n561), .ZN(n1074) );
  NAND2_X1 U671 ( .A1(\mem[30][0] ), .A2(n1570), .ZN(n561) );
  OAI21_X1 U672 ( .B1(n1636), .B2(n560), .A(n562), .ZN(n1075) );
  NAND2_X1 U673 ( .A1(\mem[30][1] ), .A2(n1570), .ZN(n562) );
  OAI21_X1 U674 ( .B1(n1635), .B2(n560), .A(n563), .ZN(n1076) );
  NAND2_X1 U675 ( .A1(\mem[30][2] ), .A2(n1570), .ZN(n563) );
  OAI21_X1 U676 ( .B1(n1634), .B2(n560), .A(n564), .ZN(n1077) );
  NAND2_X1 U677 ( .A1(\mem[30][3] ), .A2(n1570), .ZN(n564) );
  OAI21_X1 U678 ( .B1(n1633), .B2(n560), .A(n565), .ZN(n1078) );
  NAND2_X1 U679 ( .A1(\mem[30][4] ), .A2(n1570), .ZN(n565) );
  OAI21_X1 U680 ( .B1(n1632), .B2(n560), .A(n566), .ZN(n1079) );
  NAND2_X1 U681 ( .A1(\mem[30][5] ), .A2(n560), .ZN(n566) );
  OAI21_X1 U682 ( .B1(n1631), .B2(n560), .A(n567), .ZN(n1080) );
  NAND2_X1 U683 ( .A1(\mem[30][6] ), .A2(n560), .ZN(n567) );
  OAI21_X1 U684 ( .B1(n1622), .B2(n560), .A(n576), .ZN(n1089) );
  NAND2_X1 U685 ( .A1(\mem[30][15] ), .A2(n1570), .ZN(n576) );
  OAI21_X1 U686 ( .B1(n1600), .B2(n1569), .A(n39), .ZN(n594) );
  NAND2_X1 U687 ( .A1(\mem[0][0] ), .A2(n38), .ZN(n39) );
  OAI21_X1 U688 ( .B1(n1600), .B2(n1568), .A(n40), .ZN(n595) );
  NAND2_X1 U689 ( .A1(\mem[0][1] ), .A2(n38), .ZN(n40) );
  OAI21_X1 U690 ( .B1(n1600), .B2(n1567), .A(n41), .ZN(n596) );
  NAND2_X1 U691 ( .A1(\mem[0][2] ), .A2(n38), .ZN(n41) );
  OAI21_X1 U692 ( .B1(n1600), .B2(n1566), .A(n42), .ZN(n597) );
  NAND2_X1 U693 ( .A1(\mem[0][3] ), .A2(n38), .ZN(n42) );
  OAI21_X1 U694 ( .B1(n1600), .B2(n1565), .A(n43), .ZN(n598) );
  NAND2_X1 U695 ( .A1(\mem[0][4] ), .A2(n1600), .ZN(n43) );
  OAI21_X1 U696 ( .B1(n1600), .B2(n1564), .A(n44), .ZN(n599) );
  NAND2_X1 U697 ( .A1(\mem[0][5] ), .A2(n1600), .ZN(n44) );
  OAI21_X1 U698 ( .B1(n1600), .B2(n1563), .A(n45), .ZN(n600) );
  NAND2_X1 U699 ( .A1(\mem[0][6] ), .A2(n1600), .ZN(n45) );
  OAI21_X1 U700 ( .B1(n1600), .B2(n1562), .A(n46), .ZN(n601) );
  NAND2_X1 U701 ( .A1(\mem[0][7] ), .A2(n1600), .ZN(n46) );
  OAI21_X1 U702 ( .B1(n1600), .B2(n1554), .A(n54), .ZN(n609) );
  NAND2_X1 U703 ( .A1(\mem[0][15] ), .A2(n38), .ZN(n54) );
  OAI21_X1 U704 ( .B1(n1569), .B2(n57), .A(n58), .ZN(n610) );
  NAND2_X1 U705 ( .A1(\mem[1][0] ), .A2(n1599), .ZN(n58) );
  OAI21_X1 U706 ( .B1(n1568), .B2(n57), .A(n59), .ZN(n611) );
  NAND2_X1 U707 ( .A1(\mem[1][1] ), .A2(n1599), .ZN(n59) );
  OAI21_X1 U708 ( .B1(n1567), .B2(n57), .A(n60), .ZN(n612) );
  NAND2_X1 U709 ( .A1(\mem[1][2] ), .A2(n1599), .ZN(n60) );
  OAI21_X1 U710 ( .B1(n1566), .B2(n57), .A(n61), .ZN(n613) );
  NAND2_X1 U711 ( .A1(\mem[1][3] ), .A2(n1599), .ZN(n61) );
  OAI21_X1 U712 ( .B1(n1565), .B2(n57), .A(n62), .ZN(n614) );
  NAND2_X1 U713 ( .A1(\mem[1][4] ), .A2(n57), .ZN(n62) );
  OAI21_X1 U714 ( .B1(n1564), .B2(n57), .A(n63), .ZN(n615) );
  NAND2_X1 U715 ( .A1(\mem[1][5] ), .A2(n57), .ZN(n63) );
  OAI21_X1 U716 ( .B1(n1563), .B2(n57), .A(n64), .ZN(n616) );
  NAND2_X1 U717 ( .A1(\mem[1][6] ), .A2(n57), .ZN(n64) );
  OAI21_X1 U718 ( .B1(n1554), .B2(n57), .A(n73), .ZN(n625) );
  NAND2_X1 U719 ( .A1(\mem[1][15] ), .A2(n1599), .ZN(n73) );
  OAI21_X1 U720 ( .B1(n1569), .B2(n75), .A(n76), .ZN(n626) );
  NAND2_X1 U721 ( .A1(\mem[2][0] ), .A2(n1598), .ZN(n76) );
  OAI21_X1 U722 ( .B1(n1568), .B2(n75), .A(n77), .ZN(n627) );
  NAND2_X1 U723 ( .A1(\mem[2][1] ), .A2(n1598), .ZN(n77) );
  OAI21_X1 U724 ( .B1(n1567), .B2(n75), .A(n78), .ZN(n628) );
  NAND2_X1 U725 ( .A1(\mem[2][2] ), .A2(n1598), .ZN(n78) );
  OAI21_X1 U726 ( .B1(n1566), .B2(n75), .A(n79), .ZN(n629) );
  NAND2_X1 U727 ( .A1(\mem[2][3] ), .A2(n1598), .ZN(n79) );
  OAI21_X1 U728 ( .B1(n1565), .B2(n75), .A(n80), .ZN(n630) );
  NAND2_X1 U729 ( .A1(\mem[2][4] ), .A2(n75), .ZN(n80) );
  OAI21_X1 U730 ( .B1(n1564), .B2(n75), .A(n81), .ZN(n631) );
  NAND2_X1 U731 ( .A1(\mem[2][5] ), .A2(n75), .ZN(n81) );
  OAI21_X1 U732 ( .B1(n1563), .B2(n75), .A(n82), .ZN(n632) );
  NAND2_X1 U733 ( .A1(\mem[2][6] ), .A2(n75), .ZN(n82) );
  OAI21_X1 U734 ( .B1(n1554), .B2(n75), .A(n91), .ZN(n641) );
  NAND2_X1 U735 ( .A1(\mem[2][15] ), .A2(n1598), .ZN(n91) );
  OAI21_X1 U736 ( .B1(n1569), .B2(n93), .A(n94), .ZN(n642) );
  NAND2_X1 U737 ( .A1(\mem[3][0] ), .A2(n1597), .ZN(n94) );
  OAI21_X1 U738 ( .B1(n1568), .B2(n93), .A(n95), .ZN(n643) );
  NAND2_X1 U739 ( .A1(\mem[3][1] ), .A2(n1597), .ZN(n95) );
  OAI21_X1 U740 ( .B1(n1567), .B2(n93), .A(n96), .ZN(n644) );
  NAND2_X1 U741 ( .A1(\mem[3][2] ), .A2(n1597), .ZN(n96) );
  OAI21_X1 U742 ( .B1(n1566), .B2(n93), .A(n97), .ZN(n645) );
  NAND2_X1 U743 ( .A1(\mem[3][3] ), .A2(n1597), .ZN(n97) );
  OAI21_X1 U744 ( .B1(n1565), .B2(n93), .A(n98), .ZN(n646) );
  NAND2_X1 U745 ( .A1(\mem[3][4] ), .A2(n93), .ZN(n98) );
  OAI21_X1 U746 ( .B1(n1564), .B2(n93), .A(n99), .ZN(n647) );
  NAND2_X1 U747 ( .A1(\mem[3][5] ), .A2(n93), .ZN(n99) );
  OAI21_X1 U748 ( .B1(n1563), .B2(n93), .A(n100), .ZN(n648) );
  NAND2_X1 U749 ( .A1(\mem[3][6] ), .A2(n93), .ZN(n100) );
  OAI21_X1 U750 ( .B1(n1554), .B2(n93), .A(n109), .ZN(n657) );
  NAND2_X1 U751 ( .A1(\mem[3][15] ), .A2(n1597), .ZN(n109) );
  OAI21_X1 U752 ( .B1(n1569), .B2(n111), .A(n112), .ZN(n658) );
  NAND2_X1 U753 ( .A1(\mem[4][0] ), .A2(n1596), .ZN(n112) );
  OAI21_X1 U754 ( .B1(n1568), .B2(n111), .A(n113), .ZN(n659) );
  NAND2_X1 U755 ( .A1(\mem[4][1] ), .A2(n1596), .ZN(n113) );
  OAI21_X1 U756 ( .B1(n1567), .B2(n111), .A(n114), .ZN(n660) );
  NAND2_X1 U757 ( .A1(\mem[4][2] ), .A2(n1596), .ZN(n114) );
  OAI21_X1 U758 ( .B1(n1566), .B2(n111), .A(n115), .ZN(n661) );
  NAND2_X1 U759 ( .A1(\mem[4][3] ), .A2(n1596), .ZN(n115) );
  OAI21_X1 U760 ( .B1(n1565), .B2(n111), .A(n116), .ZN(n662) );
  NAND2_X1 U761 ( .A1(\mem[4][4] ), .A2(n111), .ZN(n116) );
  OAI21_X1 U762 ( .B1(n1564), .B2(n111), .A(n117), .ZN(n663) );
  NAND2_X1 U763 ( .A1(\mem[4][5] ), .A2(n111), .ZN(n117) );
  OAI21_X1 U764 ( .B1(n1563), .B2(n111), .A(n118), .ZN(n664) );
  NAND2_X1 U765 ( .A1(\mem[4][6] ), .A2(n111), .ZN(n118) );
  OAI21_X1 U766 ( .B1(n1554), .B2(n111), .A(n127), .ZN(n673) );
  NAND2_X1 U767 ( .A1(\mem[4][15] ), .A2(n1596), .ZN(n127) );
  OAI21_X1 U768 ( .B1(n1569), .B2(n1595), .A(n130), .ZN(n674) );
  NAND2_X1 U769 ( .A1(\mem[5][0] ), .A2(n129), .ZN(n130) );
  OAI21_X1 U770 ( .B1(n1568), .B2(n1595), .A(n131), .ZN(n675) );
  NAND2_X1 U771 ( .A1(\mem[5][1] ), .A2(n129), .ZN(n131) );
  OAI21_X1 U772 ( .B1(n1567), .B2(n1595), .A(n132), .ZN(n676) );
  NAND2_X1 U773 ( .A1(\mem[5][2] ), .A2(n129), .ZN(n132) );
  OAI21_X1 U774 ( .B1(n1566), .B2(n1595), .A(n133), .ZN(n677) );
  NAND2_X1 U775 ( .A1(\mem[5][3] ), .A2(n129), .ZN(n133) );
  OAI21_X1 U776 ( .B1(n1565), .B2(n1595), .A(n134), .ZN(n678) );
  NAND2_X1 U777 ( .A1(\mem[5][4] ), .A2(n1595), .ZN(n134) );
  OAI21_X1 U778 ( .B1(n1564), .B2(n1595), .A(n135), .ZN(n679) );
  NAND2_X1 U779 ( .A1(\mem[5][5] ), .A2(n1595), .ZN(n135) );
  OAI21_X1 U780 ( .B1(n1563), .B2(n1595), .A(n136), .ZN(n680) );
  NAND2_X1 U781 ( .A1(\mem[5][6] ), .A2(n1595), .ZN(n136) );
  OAI21_X1 U782 ( .B1(n1554), .B2(n1595), .A(n145), .ZN(n689) );
  NAND2_X1 U783 ( .A1(\mem[5][15] ), .A2(n129), .ZN(n145) );
  OAI21_X1 U784 ( .B1(n1569), .B2(n147), .A(n148), .ZN(n690) );
  NAND2_X1 U785 ( .A1(\mem[6][0] ), .A2(n1594), .ZN(n148) );
  OAI21_X1 U786 ( .B1(n1568), .B2(n147), .A(n149), .ZN(n691) );
  NAND2_X1 U787 ( .A1(\mem[6][1] ), .A2(n147), .ZN(n149) );
  OAI21_X1 U788 ( .B1(n1567), .B2(n147), .A(n150), .ZN(n692) );
  NAND2_X1 U789 ( .A1(\mem[6][2] ), .A2(n147), .ZN(n150) );
  OAI21_X1 U790 ( .B1(n1566), .B2(n147), .A(n151), .ZN(n693) );
  NAND2_X1 U791 ( .A1(\mem[6][3] ), .A2(n147), .ZN(n151) );
  OAI21_X1 U792 ( .B1(n1565), .B2(n147), .A(n152), .ZN(n694) );
  NAND2_X1 U793 ( .A1(\mem[6][4] ), .A2(n1594), .ZN(n152) );
  OAI21_X1 U794 ( .B1(n1564), .B2(n1594), .A(n153), .ZN(n695) );
  NAND2_X1 U795 ( .A1(\mem[6][5] ), .A2(n1594), .ZN(n153) );
  OAI21_X1 U796 ( .B1(n1563), .B2(n147), .A(n154), .ZN(n696) );
  NAND2_X1 U797 ( .A1(\mem[6][6] ), .A2(n1594), .ZN(n154) );
  OAI21_X1 U798 ( .B1(n1554), .B2(n147), .A(n163), .ZN(n705) );
  NAND2_X1 U799 ( .A1(\mem[6][15] ), .A2(n147), .ZN(n163) );
  OAI21_X1 U800 ( .B1(n1569), .B2(n165), .A(n166), .ZN(n706) );
  NAND2_X1 U801 ( .A1(\mem[7][0] ), .A2(n1593), .ZN(n166) );
  OAI21_X1 U802 ( .B1(n1568), .B2(n165), .A(n167), .ZN(n707) );
  NAND2_X1 U803 ( .A1(\mem[7][1] ), .A2(n1593), .ZN(n167) );
  OAI21_X1 U804 ( .B1(n1567), .B2(n165), .A(n168), .ZN(n708) );
  NAND2_X1 U805 ( .A1(\mem[7][2] ), .A2(n1593), .ZN(n168) );
  OAI21_X1 U806 ( .B1(n1566), .B2(n165), .A(n169), .ZN(n709) );
  NAND2_X1 U807 ( .A1(\mem[7][3] ), .A2(n1593), .ZN(n169) );
  OAI21_X1 U808 ( .B1(n1565), .B2(n165), .A(n170), .ZN(n710) );
  NAND2_X1 U809 ( .A1(\mem[7][4] ), .A2(n165), .ZN(n170) );
  OAI21_X1 U810 ( .B1(n1564), .B2(n165), .A(n171), .ZN(n711) );
  NAND2_X1 U811 ( .A1(\mem[7][5] ), .A2(n165), .ZN(n171) );
  OAI21_X1 U812 ( .B1(n1563), .B2(n165), .A(n172), .ZN(n712) );
  NAND2_X1 U813 ( .A1(\mem[7][6] ), .A2(n165), .ZN(n172) );
  OAI21_X1 U814 ( .B1(n1554), .B2(n165), .A(n181), .ZN(n721) );
  NAND2_X1 U815 ( .A1(\mem[7][15] ), .A2(n1593), .ZN(n181) );
  OAI21_X1 U816 ( .B1(n1569), .B2(n1592), .A(n184), .ZN(n722) );
  NAND2_X1 U817 ( .A1(\mem[8][0] ), .A2(n183), .ZN(n184) );
  OAI21_X1 U818 ( .B1(n1568), .B2(n183), .A(n185), .ZN(n723) );
  NAND2_X1 U819 ( .A1(\mem[8][1] ), .A2(n1592), .ZN(n185) );
  OAI21_X1 U820 ( .B1(n1567), .B2(n183), .A(n186), .ZN(n724) );
  NAND2_X1 U821 ( .A1(\mem[8][2] ), .A2(n183), .ZN(n186) );
  OAI21_X1 U822 ( .B1(n1566), .B2(n183), .A(n187), .ZN(n725) );
  NAND2_X1 U823 ( .A1(\mem[8][3] ), .A2(n183), .ZN(n187) );
  OAI21_X1 U824 ( .B1(n1565), .B2(n183), .A(n188), .ZN(n726) );
  NAND2_X1 U825 ( .A1(\mem[8][4] ), .A2(n1592), .ZN(n188) );
  OAI21_X1 U826 ( .B1(n1564), .B2(n183), .A(n189), .ZN(n727) );
  NAND2_X1 U827 ( .A1(\mem[8][5] ), .A2(n1592), .ZN(n189) );
  OAI21_X1 U828 ( .B1(n1563), .B2(n183), .A(n190), .ZN(n728) );
  NAND2_X1 U829 ( .A1(\mem[8][6] ), .A2(n1592), .ZN(n190) );
  OAI21_X1 U830 ( .B1(n1554), .B2(n183), .A(n199), .ZN(n737) );
  NAND2_X1 U831 ( .A1(\mem[8][15] ), .A2(n183), .ZN(n199) );
  OAI21_X1 U832 ( .B1(n1569), .B2(n1591), .A(n202), .ZN(n738) );
  NAND2_X1 U833 ( .A1(\mem[9][0] ), .A2(n201), .ZN(n202) );
  OAI21_X1 U834 ( .B1(n1568), .B2(n1591), .A(n203), .ZN(n739) );
  NAND2_X1 U835 ( .A1(\mem[9][1] ), .A2(n201), .ZN(n203) );
  OAI21_X1 U836 ( .B1(n1567), .B2(n1591), .A(n204), .ZN(n740) );
  NAND2_X1 U837 ( .A1(\mem[9][2] ), .A2(n201), .ZN(n204) );
  OAI21_X1 U838 ( .B1(n1566), .B2(n1591), .A(n205), .ZN(n741) );
  NAND2_X1 U839 ( .A1(\mem[9][3] ), .A2(n201), .ZN(n205) );
  OAI21_X1 U840 ( .B1(n1565), .B2(n1591), .A(n206), .ZN(n742) );
  NAND2_X1 U841 ( .A1(\mem[9][4] ), .A2(n1591), .ZN(n206) );
  OAI21_X1 U842 ( .B1(n1564), .B2(n1591), .A(n207), .ZN(n743) );
  NAND2_X1 U843 ( .A1(\mem[9][5] ), .A2(n1591), .ZN(n207) );
  OAI21_X1 U844 ( .B1(n1563), .B2(n1591), .A(n208), .ZN(n744) );
  NAND2_X1 U845 ( .A1(\mem[9][6] ), .A2(n1591), .ZN(n208) );
  OAI21_X1 U846 ( .B1(n1554), .B2(n1591), .A(n217), .ZN(n753) );
  NAND2_X1 U847 ( .A1(\mem[9][15] ), .A2(n201), .ZN(n217) );
  OAI21_X1 U848 ( .B1(n1569), .B2(n218), .A(n219), .ZN(n754) );
  NAND2_X1 U849 ( .A1(\mem[10][0] ), .A2(n1590), .ZN(n219) );
  OAI21_X1 U850 ( .B1(n1568), .B2(n218), .A(n220), .ZN(n755) );
  NAND2_X1 U851 ( .A1(\mem[10][1] ), .A2(n1590), .ZN(n220) );
  OAI21_X1 U852 ( .B1(n1567), .B2(n218), .A(n221), .ZN(n756) );
  NAND2_X1 U853 ( .A1(\mem[10][2] ), .A2(n1590), .ZN(n221) );
  OAI21_X1 U854 ( .B1(n1566), .B2(n218), .A(n222), .ZN(n757) );
  NAND2_X1 U855 ( .A1(\mem[10][3] ), .A2(n1590), .ZN(n222) );
  OAI21_X1 U856 ( .B1(n1565), .B2(n218), .A(n223), .ZN(n758) );
  NAND2_X1 U857 ( .A1(\mem[10][4] ), .A2(n218), .ZN(n223) );
  OAI21_X1 U858 ( .B1(n1564), .B2(n218), .A(n224), .ZN(n759) );
  NAND2_X1 U859 ( .A1(\mem[10][5] ), .A2(n218), .ZN(n224) );
  OAI21_X1 U860 ( .B1(n1563), .B2(n218), .A(n225), .ZN(n760) );
  NAND2_X1 U861 ( .A1(\mem[10][6] ), .A2(n218), .ZN(n225) );
  OAI21_X1 U862 ( .B1(n1554), .B2(n218), .A(n234), .ZN(n769) );
  NAND2_X1 U863 ( .A1(\mem[10][15] ), .A2(n1590), .ZN(n234) );
  OAI21_X1 U864 ( .B1(n1569), .B2(n235), .A(n236), .ZN(n770) );
  NAND2_X1 U865 ( .A1(\mem[11][0] ), .A2(n1589), .ZN(n236) );
  OAI21_X1 U866 ( .B1(n1568), .B2(n235), .A(n237), .ZN(n771) );
  NAND2_X1 U867 ( .A1(\mem[11][1] ), .A2(n1589), .ZN(n237) );
  OAI21_X1 U868 ( .B1(n1567), .B2(n235), .A(n238), .ZN(n772) );
  NAND2_X1 U869 ( .A1(\mem[11][2] ), .A2(n1589), .ZN(n238) );
  OAI21_X1 U870 ( .B1(n1566), .B2(n235), .A(n239), .ZN(n773) );
  NAND2_X1 U871 ( .A1(\mem[11][3] ), .A2(n1589), .ZN(n239) );
  OAI21_X1 U872 ( .B1(n1565), .B2(n235), .A(n240), .ZN(n774) );
  NAND2_X1 U873 ( .A1(\mem[11][4] ), .A2(n235), .ZN(n240) );
  OAI21_X1 U874 ( .B1(n1564), .B2(n235), .A(n241), .ZN(n775) );
  NAND2_X1 U875 ( .A1(\mem[11][5] ), .A2(n235), .ZN(n241) );
  OAI21_X1 U876 ( .B1(n1563), .B2(n235), .A(n242), .ZN(n776) );
  NAND2_X1 U877 ( .A1(\mem[11][6] ), .A2(n235), .ZN(n242) );
  OAI21_X1 U878 ( .B1(n1554), .B2(n235), .A(n251), .ZN(n785) );
  NAND2_X1 U879 ( .A1(\mem[11][15] ), .A2(n1589), .ZN(n251) );
  OAI21_X1 U880 ( .B1(n1569), .B2(n252), .A(n253), .ZN(n786) );
  NAND2_X1 U881 ( .A1(\mem[12][0] ), .A2(n1588), .ZN(n253) );
  OAI21_X1 U882 ( .B1(n1568), .B2(n252), .A(n254), .ZN(n787) );
  NAND2_X1 U883 ( .A1(\mem[12][1] ), .A2(n1588), .ZN(n254) );
  OAI21_X1 U884 ( .B1(n1567), .B2(n252), .A(n255), .ZN(n788) );
  NAND2_X1 U885 ( .A1(\mem[12][2] ), .A2(n1588), .ZN(n255) );
  OAI21_X1 U886 ( .B1(n1566), .B2(n252), .A(n256), .ZN(n789) );
  NAND2_X1 U887 ( .A1(\mem[12][3] ), .A2(n1588), .ZN(n256) );
  OAI21_X1 U888 ( .B1(n1565), .B2(n252), .A(n257), .ZN(n790) );
  NAND2_X1 U889 ( .A1(\mem[12][4] ), .A2(n252), .ZN(n257) );
  OAI21_X1 U890 ( .B1(n1564), .B2(n252), .A(n258), .ZN(n791) );
  NAND2_X1 U891 ( .A1(\mem[12][5] ), .A2(n252), .ZN(n258) );
  OAI21_X1 U892 ( .B1(n1563), .B2(n252), .A(n259), .ZN(n792) );
  NAND2_X1 U893 ( .A1(\mem[12][6] ), .A2(n252), .ZN(n259) );
  OAI21_X1 U894 ( .B1(n1554), .B2(n252), .A(n268), .ZN(n801) );
  NAND2_X1 U895 ( .A1(\mem[12][15] ), .A2(n1588), .ZN(n268) );
  OAI21_X1 U896 ( .B1(n1637), .B2(n269), .A(n270), .ZN(n802) );
  NAND2_X1 U897 ( .A1(\mem[13][0] ), .A2(n1587), .ZN(n270) );
  OAI21_X1 U898 ( .B1(n1636), .B2(n269), .A(n271), .ZN(n803) );
  NAND2_X1 U899 ( .A1(\mem[13][1] ), .A2(n1587), .ZN(n271) );
  OAI21_X1 U900 ( .B1(n1635), .B2(n269), .A(n272), .ZN(n804) );
  NAND2_X1 U901 ( .A1(\mem[13][2] ), .A2(n1587), .ZN(n272) );
  OAI21_X1 U902 ( .B1(n1634), .B2(n269), .A(n273), .ZN(n805) );
  NAND2_X1 U903 ( .A1(\mem[13][3] ), .A2(n1587), .ZN(n273) );
  OAI21_X1 U904 ( .B1(n1633), .B2(n269), .A(n274), .ZN(n806) );
  NAND2_X1 U905 ( .A1(\mem[13][4] ), .A2(n269), .ZN(n274) );
  OAI21_X1 U906 ( .B1(n1632), .B2(n269), .A(n275), .ZN(n807) );
  NAND2_X1 U907 ( .A1(\mem[13][5] ), .A2(n269), .ZN(n275) );
  OAI21_X1 U908 ( .B1(n1631), .B2(n269), .A(n276), .ZN(n808) );
  NAND2_X1 U909 ( .A1(\mem[13][6] ), .A2(n269), .ZN(n276) );
  OAI21_X1 U910 ( .B1(n1622), .B2(n269), .A(n285), .ZN(n817) );
  NAND2_X1 U911 ( .A1(\mem[13][15] ), .A2(n1587), .ZN(n285) );
  OAI21_X1 U912 ( .B1(n1637), .B2(n286), .A(n287), .ZN(n818) );
  NAND2_X1 U913 ( .A1(\mem[14][0] ), .A2(n1586), .ZN(n287) );
  OAI21_X1 U914 ( .B1(n1636), .B2(n286), .A(n288), .ZN(n819) );
  NAND2_X1 U915 ( .A1(\mem[14][1] ), .A2(n1586), .ZN(n288) );
  OAI21_X1 U916 ( .B1(n1635), .B2(n286), .A(n289), .ZN(n820) );
  NAND2_X1 U917 ( .A1(\mem[14][2] ), .A2(n1586), .ZN(n289) );
  OAI21_X1 U918 ( .B1(n1634), .B2(n286), .A(n290), .ZN(n821) );
  NAND2_X1 U919 ( .A1(\mem[14][3] ), .A2(n1586), .ZN(n290) );
  OAI21_X1 U920 ( .B1(n1633), .B2(n286), .A(n291), .ZN(n822) );
  NAND2_X1 U921 ( .A1(\mem[14][4] ), .A2(n286), .ZN(n291) );
  OAI21_X1 U922 ( .B1(n1632), .B2(n286), .A(n292), .ZN(n823) );
  NAND2_X1 U923 ( .A1(\mem[14][5] ), .A2(n286), .ZN(n292) );
  OAI21_X1 U924 ( .B1(n1631), .B2(n286), .A(n293), .ZN(n824) );
  NAND2_X1 U925 ( .A1(\mem[14][6] ), .A2(n286), .ZN(n293) );
  OAI21_X1 U926 ( .B1(n1622), .B2(n286), .A(n302), .ZN(n833) );
  NAND2_X1 U927 ( .A1(\mem[14][15] ), .A2(n1586), .ZN(n302) );
  OAI21_X1 U928 ( .B1(n1637), .B2(n303), .A(n304), .ZN(n834) );
  NAND2_X1 U929 ( .A1(\mem[15][0] ), .A2(n1585), .ZN(n304) );
  OAI21_X1 U930 ( .B1(n1636), .B2(n303), .A(n305), .ZN(n835) );
  NAND2_X1 U931 ( .A1(\mem[15][1] ), .A2(n1585), .ZN(n305) );
  OAI21_X1 U932 ( .B1(n1635), .B2(n303), .A(n306), .ZN(n836) );
  NAND2_X1 U933 ( .A1(\mem[15][2] ), .A2(n1585), .ZN(n306) );
  OAI21_X1 U934 ( .B1(n1634), .B2(n303), .A(n307), .ZN(n837) );
  NAND2_X1 U935 ( .A1(\mem[15][3] ), .A2(n1585), .ZN(n307) );
  OAI21_X1 U936 ( .B1(n1633), .B2(n303), .A(n308), .ZN(n838) );
  NAND2_X1 U937 ( .A1(\mem[15][4] ), .A2(n303), .ZN(n308) );
  OAI21_X1 U938 ( .B1(n1632), .B2(n303), .A(n309), .ZN(n839) );
  NAND2_X1 U939 ( .A1(\mem[15][5] ), .A2(n303), .ZN(n309) );
  OAI21_X1 U940 ( .B1(n1631), .B2(n303), .A(n310), .ZN(n840) );
  NAND2_X1 U941 ( .A1(\mem[15][6] ), .A2(n303), .ZN(n310) );
  OAI21_X1 U942 ( .B1(n1622), .B2(n303), .A(n319), .ZN(n849) );
  NAND2_X1 U943 ( .A1(\mem[15][15] ), .A2(n1585), .ZN(n319) );
  OAI21_X1 U944 ( .B1(n1637), .B2(n1584), .A(n321), .ZN(n850) );
  NAND2_X1 U945 ( .A1(\mem[16][0] ), .A2(n320), .ZN(n321) );
  OAI21_X1 U946 ( .B1(n1636), .B2(n1584), .A(n322), .ZN(n851) );
  NAND2_X1 U947 ( .A1(\mem[16][1] ), .A2(n320), .ZN(n322) );
  OAI21_X1 U948 ( .B1(n1635), .B2(n1584), .A(n323), .ZN(n852) );
  NAND2_X1 U949 ( .A1(\mem[16][2] ), .A2(n320), .ZN(n323) );
  OAI21_X1 U950 ( .B1(n1634), .B2(n1584), .A(n324), .ZN(n853) );
  NAND2_X1 U951 ( .A1(\mem[16][3] ), .A2(n320), .ZN(n324) );
  OAI21_X1 U952 ( .B1(n1633), .B2(n1584), .A(n325), .ZN(n854) );
  NAND2_X1 U953 ( .A1(\mem[16][4] ), .A2(n1584), .ZN(n325) );
  OAI21_X1 U954 ( .B1(n1632), .B2(n1584), .A(n326), .ZN(n855) );
  NAND2_X1 U955 ( .A1(\mem[16][5] ), .A2(n1584), .ZN(n326) );
  OAI21_X1 U956 ( .B1(n1631), .B2(n1584), .A(n327), .ZN(n856) );
  NAND2_X1 U957 ( .A1(\mem[16][6] ), .A2(n1584), .ZN(n327) );
  OAI21_X1 U958 ( .B1(n1622), .B2(n1584), .A(n336), .ZN(n865) );
  NAND2_X1 U959 ( .A1(\mem[16][15] ), .A2(n320), .ZN(n336) );
  OAI21_X1 U960 ( .B1(n1637), .B2(n338), .A(n339), .ZN(n866) );
  NAND2_X1 U961 ( .A1(\mem[17][0] ), .A2(n1583), .ZN(n339) );
  OAI21_X1 U962 ( .B1(n1636), .B2(n338), .A(n340), .ZN(n867) );
  NAND2_X1 U963 ( .A1(\mem[17][1] ), .A2(n1583), .ZN(n340) );
  OAI21_X1 U964 ( .B1(n1635), .B2(n338), .A(n341), .ZN(n868) );
  NAND2_X1 U965 ( .A1(\mem[17][2] ), .A2(n1583), .ZN(n341) );
  OAI21_X1 U966 ( .B1(n1634), .B2(n338), .A(n342), .ZN(n869) );
  NAND2_X1 U967 ( .A1(\mem[17][3] ), .A2(n1583), .ZN(n342) );
  OAI21_X1 U968 ( .B1(n1633), .B2(n338), .A(n343), .ZN(n870) );
  NAND2_X1 U969 ( .A1(\mem[17][4] ), .A2(n338), .ZN(n343) );
  OAI21_X1 U970 ( .B1(n1632), .B2(n338), .A(n344), .ZN(n871) );
  NAND2_X1 U971 ( .A1(\mem[17][5] ), .A2(n338), .ZN(n344) );
  OAI21_X1 U972 ( .B1(n1631), .B2(n338), .A(n345), .ZN(n872) );
  NAND2_X1 U973 ( .A1(\mem[17][6] ), .A2(n338), .ZN(n345) );
  OAI21_X1 U974 ( .B1(n1622), .B2(n338), .A(n354), .ZN(n881) );
  NAND2_X1 U975 ( .A1(\mem[17][15] ), .A2(n1583), .ZN(n354) );
  OAI21_X1 U976 ( .B1(n1637), .B2(n355), .A(n356), .ZN(n882) );
  NAND2_X1 U977 ( .A1(\mem[18][0] ), .A2(n1582), .ZN(n356) );
  OAI21_X1 U978 ( .B1(n1636), .B2(n355), .A(n357), .ZN(n883) );
  NAND2_X1 U979 ( .A1(\mem[18][1] ), .A2(n1582), .ZN(n357) );
  OAI21_X1 U980 ( .B1(n1635), .B2(n355), .A(n358), .ZN(n884) );
  NAND2_X1 U981 ( .A1(\mem[18][2] ), .A2(n1582), .ZN(n358) );
  OAI21_X1 U982 ( .B1(n1634), .B2(n355), .A(n359), .ZN(n885) );
  NAND2_X1 U983 ( .A1(\mem[18][3] ), .A2(n1582), .ZN(n359) );
  OAI21_X1 U984 ( .B1(n1633), .B2(n355), .A(n360), .ZN(n886) );
  NAND2_X1 U985 ( .A1(\mem[18][4] ), .A2(n355), .ZN(n360) );
  OAI21_X1 U986 ( .B1(n1632), .B2(n355), .A(n361), .ZN(n887) );
  NAND2_X1 U987 ( .A1(\mem[18][5] ), .A2(n355), .ZN(n361) );
  OAI21_X1 U988 ( .B1(n1631), .B2(n355), .A(n362), .ZN(n888) );
  NAND2_X1 U989 ( .A1(\mem[18][6] ), .A2(n355), .ZN(n362) );
  OAI21_X1 U990 ( .B1(n1622), .B2(n355), .A(n371), .ZN(n897) );
  NAND2_X1 U991 ( .A1(\mem[18][15] ), .A2(n1582), .ZN(n371) );
  OAI21_X1 U992 ( .B1(n1637), .B2(n372), .A(n373), .ZN(n898) );
  NAND2_X1 U993 ( .A1(\mem[19][0] ), .A2(n1581), .ZN(n373) );
  OAI21_X1 U994 ( .B1(n1636), .B2(n372), .A(n374), .ZN(n899) );
  NAND2_X1 U995 ( .A1(\mem[19][1] ), .A2(n1581), .ZN(n374) );
  OAI21_X1 U996 ( .B1(n1635), .B2(n372), .A(n375), .ZN(n900) );
  NAND2_X1 U997 ( .A1(\mem[19][2] ), .A2(n1581), .ZN(n375) );
  OAI21_X1 U998 ( .B1(n1634), .B2(n372), .A(n376), .ZN(n901) );
  NAND2_X1 U999 ( .A1(\mem[19][3] ), .A2(n1581), .ZN(n376) );
  OAI21_X1 U1000 ( .B1(n1633), .B2(n372), .A(n377), .ZN(n902) );
  NAND2_X1 U1001 ( .A1(\mem[19][4] ), .A2(n372), .ZN(n377) );
  OAI21_X1 U1002 ( .B1(n1632), .B2(n372), .A(n378), .ZN(n903) );
  NAND2_X1 U1003 ( .A1(\mem[19][5] ), .A2(n372), .ZN(n378) );
  OAI21_X1 U1004 ( .B1(n1631), .B2(n372), .A(n379), .ZN(n904) );
  NAND2_X1 U1005 ( .A1(\mem[19][6] ), .A2(n372), .ZN(n379) );
  OAI21_X1 U1006 ( .B1(n1622), .B2(n372), .A(n388), .ZN(n913) );
  NAND2_X1 U1007 ( .A1(\mem[19][15] ), .A2(n1581), .ZN(n388) );
  OAI21_X1 U1008 ( .B1(n1637), .B2(n389), .A(n390), .ZN(n914) );
  NAND2_X1 U1009 ( .A1(\mem[20][0] ), .A2(n1580), .ZN(n390) );
  OAI21_X1 U1010 ( .B1(n1636), .B2(n389), .A(n391), .ZN(n915) );
  NAND2_X1 U1011 ( .A1(\mem[20][1] ), .A2(n1580), .ZN(n391) );
  OAI21_X1 U1012 ( .B1(n1635), .B2(n389), .A(n392), .ZN(n916) );
  NAND2_X1 U1013 ( .A1(\mem[20][2] ), .A2(n1580), .ZN(n392) );
  OAI21_X1 U1014 ( .B1(n1634), .B2(n389), .A(n393), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(\mem[20][3] ), .A2(n1580), .ZN(n393) );
  OAI21_X1 U1016 ( .B1(n1633), .B2(n389), .A(n394), .ZN(n918) );
  NAND2_X1 U1017 ( .A1(\mem[20][4] ), .A2(n389), .ZN(n394) );
  OAI21_X1 U1018 ( .B1(n1632), .B2(n389), .A(n395), .ZN(n919) );
  NAND2_X1 U1019 ( .A1(\mem[20][5] ), .A2(n389), .ZN(n395) );
  OAI21_X1 U1020 ( .B1(n1631), .B2(n389), .A(n396), .ZN(n920) );
  NAND2_X1 U1021 ( .A1(\mem[20][6] ), .A2(n389), .ZN(n396) );
  OAI21_X1 U1022 ( .B1(n1622), .B2(n389), .A(n405), .ZN(n929) );
  NAND2_X1 U1023 ( .A1(\mem[20][15] ), .A2(n1580), .ZN(n405) );
  OAI21_X1 U1024 ( .B1(n1637), .B2(n406), .A(n407), .ZN(n930) );
  NAND2_X1 U1025 ( .A1(\mem[21][0] ), .A2(n1579), .ZN(n407) );
  OAI21_X1 U1026 ( .B1(n1636), .B2(n406), .A(n408), .ZN(n931) );
  NAND2_X1 U1027 ( .A1(\mem[21][1] ), .A2(n1579), .ZN(n408) );
  OAI21_X1 U1028 ( .B1(n1635), .B2(n406), .A(n409), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(\mem[21][2] ), .A2(n1579), .ZN(n409) );
  OAI21_X1 U1030 ( .B1(n1634), .B2(n406), .A(n410), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(\mem[21][3] ), .A2(n1579), .ZN(n410) );
  OAI21_X1 U1032 ( .B1(n1633), .B2(n406), .A(n411), .ZN(n934) );
  NAND2_X1 U1033 ( .A1(\mem[21][4] ), .A2(n406), .ZN(n411) );
  OAI21_X1 U1034 ( .B1(n1632), .B2(n406), .A(n412), .ZN(n935) );
  NAND2_X1 U1035 ( .A1(\mem[21][5] ), .A2(n406), .ZN(n412) );
  OAI21_X1 U1036 ( .B1(n1631), .B2(n406), .A(n413), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(\mem[21][6] ), .A2(n406), .ZN(n413) );
  OAI21_X1 U1038 ( .B1(n1622), .B2(n406), .A(n422), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(\mem[21][15] ), .A2(n1579), .ZN(n422) );
  OAI21_X1 U1040 ( .B1(n1637), .B2(n1578), .A(n424), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(\mem[22][0] ), .A2(n423), .ZN(n424) );
  OAI21_X1 U1042 ( .B1(n1636), .B2(n1578), .A(n425), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(\mem[22][1] ), .A2(n423), .ZN(n425) );
  OAI21_X1 U1044 ( .B1(n1635), .B2(n1578), .A(n426), .ZN(n948) );
  NAND2_X1 U1045 ( .A1(\mem[22][2] ), .A2(n423), .ZN(n426) );
  OAI21_X1 U1046 ( .B1(n1634), .B2(n1578), .A(n427), .ZN(n949) );
  NAND2_X1 U1047 ( .A1(\mem[22][3] ), .A2(n423), .ZN(n427) );
  OAI21_X1 U1048 ( .B1(n1633), .B2(n1578), .A(n428), .ZN(n950) );
  NAND2_X1 U1049 ( .A1(\mem[22][4] ), .A2(n1578), .ZN(n428) );
  OAI21_X1 U1050 ( .B1(n1632), .B2(n1578), .A(n429), .ZN(n951) );
  NAND2_X1 U1051 ( .A1(\mem[22][5] ), .A2(n1578), .ZN(n429) );
  OAI21_X1 U1052 ( .B1(n1631), .B2(n1578), .A(n430), .ZN(n952) );
  NAND2_X1 U1053 ( .A1(\mem[22][6] ), .A2(n1578), .ZN(n430) );
  OAI21_X1 U1054 ( .B1(n1622), .B2(n1578), .A(n439), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(\mem[22][15] ), .A2(n423), .ZN(n439) );
  OAI21_X1 U1056 ( .B1(n1637), .B2(n440), .A(n441), .ZN(n962) );
  NAND2_X1 U1057 ( .A1(\mem[23][0] ), .A2(n1577), .ZN(n441) );
  OAI21_X1 U1058 ( .B1(n1636), .B2(n440), .A(n442), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(\mem[23][1] ), .A2(n1577), .ZN(n442) );
  OAI21_X1 U1060 ( .B1(n1635), .B2(n440), .A(n443), .ZN(n964) );
  NAND2_X1 U1061 ( .A1(\mem[23][2] ), .A2(n1577), .ZN(n443) );
  OAI21_X1 U1062 ( .B1(n1634), .B2(n440), .A(n444), .ZN(n965) );
  NAND2_X1 U1063 ( .A1(\mem[23][3] ), .A2(n1577), .ZN(n444) );
  OAI21_X1 U1064 ( .B1(n1633), .B2(n440), .A(n445), .ZN(n966) );
  NAND2_X1 U1065 ( .A1(\mem[23][4] ), .A2(n440), .ZN(n445) );
  OAI21_X1 U1066 ( .B1(n1632), .B2(n440), .A(n446), .ZN(n967) );
  NAND2_X1 U1067 ( .A1(\mem[23][5] ), .A2(n440), .ZN(n446) );
  OAI21_X1 U1068 ( .B1(n1631), .B2(n440), .A(n447), .ZN(n968) );
  NAND2_X1 U1069 ( .A1(\mem[23][6] ), .A2(n440), .ZN(n447) );
  OAI21_X1 U1070 ( .B1(n1622), .B2(n440), .A(n456), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(\mem[23][15] ), .A2(n1577), .ZN(n456) );
  OAI21_X1 U1072 ( .B1(n1637), .B2(n457), .A(n458), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(\mem[24][0] ), .A2(n1576), .ZN(n458) );
  OAI21_X1 U1074 ( .B1(n1636), .B2(n457), .A(n459), .ZN(n979) );
  NAND2_X1 U1075 ( .A1(\mem[24][1] ), .A2(n1576), .ZN(n459) );
  OAI21_X1 U1076 ( .B1(n1635), .B2(n457), .A(n460), .ZN(n980) );
  NAND2_X1 U1077 ( .A1(\mem[24][2] ), .A2(n1576), .ZN(n460) );
  OAI21_X1 U1078 ( .B1(n1634), .B2(n457), .A(n461), .ZN(n981) );
  NAND2_X1 U1079 ( .A1(\mem[24][3] ), .A2(n1576), .ZN(n461) );
  OAI21_X1 U1080 ( .B1(n1633), .B2(n457), .A(n462), .ZN(n982) );
  NAND2_X1 U1081 ( .A1(\mem[24][4] ), .A2(n457), .ZN(n462) );
  OAI21_X1 U1082 ( .B1(n1632), .B2(n457), .A(n463), .ZN(n983) );
  NAND2_X1 U1083 ( .A1(\mem[24][5] ), .A2(n457), .ZN(n463) );
  OAI21_X1 U1084 ( .B1(n1631), .B2(n457), .A(n464), .ZN(n984) );
  NAND2_X1 U1085 ( .A1(\mem[24][6] ), .A2(n457), .ZN(n464) );
  OAI21_X1 U1086 ( .B1(n1622), .B2(n457), .A(n473), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(\mem[24][15] ), .A2(n1576), .ZN(n473) );
  OAI21_X1 U1088 ( .B1(n1637), .B2(n475), .A(n476), .ZN(n994) );
  NAND2_X1 U1089 ( .A1(\mem[25][0] ), .A2(n1575), .ZN(n476) );
  OAI21_X1 U1090 ( .B1(n1636), .B2(n475), .A(n477), .ZN(n995) );
  NAND2_X1 U1091 ( .A1(\mem[25][1] ), .A2(n1575), .ZN(n477) );
  OAI21_X1 U1092 ( .B1(n1635), .B2(n475), .A(n478), .ZN(n996) );
  NAND2_X1 U1093 ( .A1(\mem[25][2] ), .A2(n1575), .ZN(n478) );
  OAI21_X1 U1094 ( .B1(n1634), .B2(n475), .A(n479), .ZN(n997) );
  NAND2_X1 U1095 ( .A1(\mem[25][3] ), .A2(n1575), .ZN(n479) );
  OAI21_X1 U1096 ( .B1(n1633), .B2(n475), .A(n480), .ZN(n998) );
  NAND2_X1 U1097 ( .A1(\mem[25][4] ), .A2(n475), .ZN(n480) );
  OAI21_X1 U1098 ( .B1(n1632), .B2(n475), .A(n481), .ZN(n999) );
  NAND2_X1 U1099 ( .A1(\mem[25][5] ), .A2(n475), .ZN(n481) );
  OAI21_X1 U1100 ( .B1(n1631), .B2(n475), .A(n482), .ZN(n1000) );
  NAND2_X1 U1101 ( .A1(\mem[25][6] ), .A2(n475), .ZN(n482) );
  OAI21_X1 U1102 ( .B1(n1622), .B2(n475), .A(n491), .ZN(n1009) );
  NAND2_X1 U1103 ( .A1(\mem[25][15] ), .A2(n1575), .ZN(n491) );
  INV_X1 U1104 ( .A(n577), .ZN(n1620) );
  AOI22_X1 U1105 ( .A1(data_in[0]), .A2(n1621), .B1(n578), .B2(\mem[31][0] ), 
        .ZN(n577) );
  INV_X1 U1106 ( .A(n579), .ZN(n1619) );
  AOI22_X1 U1107 ( .A1(data_in[1]), .A2(n1621), .B1(n578), .B2(\mem[31][1] ), 
        .ZN(n579) );
  INV_X1 U1108 ( .A(n580), .ZN(n1618) );
  AOI22_X1 U1109 ( .A1(data_in[2]), .A2(n1621), .B1(n578), .B2(\mem[31][2] ), 
        .ZN(n580) );
  INV_X1 U1110 ( .A(n581), .ZN(n1617) );
  AOI22_X1 U1111 ( .A1(data_in[3]), .A2(n1621), .B1(n578), .B2(\mem[31][3] ), 
        .ZN(n581) );
  INV_X1 U1112 ( .A(n582), .ZN(n1616) );
  AOI22_X1 U1113 ( .A1(data_in[4]), .A2(n1621), .B1(n578), .B2(\mem[31][4] ), 
        .ZN(n582) );
  INV_X1 U1114 ( .A(n583), .ZN(n1615) );
  AOI22_X1 U1115 ( .A1(data_in[5]), .A2(n1621), .B1(n578), .B2(\mem[31][5] ), 
        .ZN(n583) );
  INV_X1 U1116 ( .A(n584), .ZN(n1614) );
  AOI22_X1 U1117 ( .A1(data_in[6]), .A2(n1621), .B1(n578), .B2(\mem[31][6] ), 
        .ZN(n584) );
  INV_X1 U1118 ( .A(n585), .ZN(n1613) );
  AOI22_X1 U1119 ( .A1(data_in[7]), .A2(n1621), .B1(n578), .B2(\mem[31][7] ), 
        .ZN(n585) );
  INV_X1 U1120 ( .A(n586), .ZN(n1612) );
  AOI22_X1 U1121 ( .A1(data_in[8]), .A2(n1621), .B1(n578), .B2(\mem[31][8] ), 
        .ZN(n586) );
  INV_X1 U1122 ( .A(n587), .ZN(n1611) );
  AOI22_X1 U1123 ( .A1(data_in[9]), .A2(n1621), .B1(n578), .B2(\mem[31][9] ), 
        .ZN(n587) );
  INV_X1 U1124 ( .A(n588), .ZN(n1610) );
  AOI22_X1 U1125 ( .A1(data_in[10]), .A2(n1621), .B1(n578), .B2(\mem[31][10] ), 
        .ZN(n588) );
  INV_X1 U1126 ( .A(n589), .ZN(n1609) );
  AOI22_X1 U1127 ( .A1(data_in[11]), .A2(n1621), .B1(n578), .B2(\mem[31][11] ), 
        .ZN(n589) );
  INV_X1 U1128 ( .A(n590), .ZN(n1608) );
  AOI22_X1 U1129 ( .A1(data_in[12]), .A2(n1621), .B1(n578), .B2(\mem[31][12] ), 
        .ZN(n590) );
  INV_X1 U1130 ( .A(n591), .ZN(n1607) );
  AOI22_X1 U1131 ( .A1(data_in[13]), .A2(n1621), .B1(n578), .B2(\mem[31][13] ), 
        .ZN(n591) );
  INV_X1 U1132 ( .A(n592), .ZN(n1606) );
  AOI22_X1 U1133 ( .A1(data_in[14]), .A2(n1621), .B1(n578), .B2(\mem[31][14] ), 
        .ZN(n592) );
  INV_X1 U1134 ( .A(n593), .ZN(n1605) );
  AOI22_X1 U1135 ( .A1(data_in[15]), .A2(n1621), .B1(n578), .B2(\mem[31][15] ), 
        .ZN(n593) );
  INV_X1 U1136 ( .A(data_in[0]), .ZN(n1637) );
  INV_X1 U1137 ( .A(data_in[1]), .ZN(n1636) );
  INV_X1 U1138 ( .A(data_in[2]), .ZN(n1635) );
  INV_X1 U1139 ( .A(data_in[3]), .ZN(n1634) );
  INV_X1 U1140 ( .A(data_in[4]), .ZN(n1633) );
  INV_X1 U1141 ( .A(data_in[5]), .ZN(n1632) );
  INV_X1 U1142 ( .A(data_in[6]), .ZN(n1631) );
  INV_X1 U1143 ( .A(data_in[7]), .ZN(n1630) );
  INV_X1 U1144 ( .A(data_in[8]), .ZN(n1629) );
  INV_X1 U1145 ( .A(data_in[9]), .ZN(n1628) );
  INV_X1 U1146 ( .A(data_in[10]), .ZN(n1627) );
  INV_X1 U1147 ( .A(data_in[11]), .ZN(n1626) );
  INV_X1 U1148 ( .A(data_in[12]), .ZN(n1625) );
  INV_X1 U1149 ( .A(data_in[13]), .ZN(n1624) );
  INV_X1 U1150 ( .A(data_in[14]), .ZN(n1623) );
  INV_X1 U1151 ( .A(data_in[15]), .ZN(n1622) );
  MUX2_X1 U1152 ( .A(\mem[30][0] ), .B(\mem[31][0] ), .S(n1543), .Z(n1) );
  MUX2_X1 U1153 ( .A(\mem[28][0] ), .B(\mem[29][0] ), .S(n1546), .Z(n2) );
  MUX2_X1 U1154 ( .A(n2), .B(n1), .S(n1537), .Z(n3) );
  MUX2_X1 U1155 ( .A(\mem[26][0] ), .B(\mem[27][0] ), .S(n1547), .Z(n4) );
  MUX2_X1 U1156 ( .A(\mem[24][0] ), .B(\mem[25][0] ), .S(n1547), .Z(n5) );
  MUX2_X1 U1157 ( .A(n5), .B(n4), .S(n1537), .Z(n6) );
  MUX2_X1 U1158 ( .A(n6), .B(n3), .S(n1534), .Z(n7) );
  MUX2_X1 U1159 ( .A(\mem[22][0] ), .B(\mem[23][0] ), .S(n1553), .Z(n8) );
  MUX2_X1 U1160 ( .A(\mem[20][0] ), .B(\mem[21][0] ), .S(n1551), .Z(n9) );
  MUX2_X1 U1161 ( .A(n9), .B(n8), .S(n1537), .Z(n10) );
  MUX2_X1 U1162 ( .A(\mem[18][0] ), .B(\mem[19][0] ), .S(n1553), .Z(n11) );
  MUX2_X1 U1163 ( .A(\mem[16][0] ), .B(\mem[17][0] ), .S(n1549), .Z(n12) );
  MUX2_X1 U1164 ( .A(n12), .B(n11), .S(n1537), .Z(n13) );
  MUX2_X1 U1165 ( .A(n13), .B(n10), .S(n1534), .Z(n14) );
  MUX2_X1 U1166 ( .A(n14), .B(n7), .S(n1533), .Z(n15) );
  MUX2_X1 U1167 ( .A(\mem[14][0] ), .B(\mem[15][0] ), .S(n1551), .Z(n16) );
  MUX2_X1 U1168 ( .A(\mem[12][0] ), .B(\mem[13][0] ), .S(n1553), .Z(n17) );
  MUX2_X1 U1169 ( .A(n17), .B(n16), .S(n1537), .Z(n18) );
  MUX2_X1 U1170 ( .A(\mem[10][0] ), .B(\mem[11][0] ), .S(n1549), .Z(n19) );
  MUX2_X1 U1171 ( .A(\mem[8][0] ), .B(\mem[9][0] ), .S(n1553), .Z(n20) );
  MUX2_X1 U1172 ( .A(n20), .B(n19), .S(n1537), .Z(n21) );
  MUX2_X1 U1173 ( .A(n21), .B(n18), .S(n1534), .Z(n22) );
  MUX2_X1 U1174 ( .A(\mem[6][0] ), .B(\mem[7][0] ), .S(n1547), .Z(n23) );
  MUX2_X1 U1175 ( .A(\mem[4][0] ), .B(\mem[5][0] ), .S(n1553), .Z(n24) );
  MUX2_X1 U1176 ( .A(n24), .B(n23), .S(n1537), .Z(n25) );
  MUX2_X1 U1177 ( .A(\mem[2][0] ), .B(\mem[3][0] ), .S(n1546), .Z(n26) );
  MUX2_X1 U1178 ( .A(\mem[0][0] ), .B(\mem[1][0] ), .S(n1547), .Z(n27) );
  MUX2_X1 U1179 ( .A(n27), .B(n26), .S(n1537), .Z(n28) );
  MUX2_X1 U1180 ( .A(n28), .B(n25), .S(n1534), .Z(n29) );
  MUX2_X1 U1181 ( .A(n29), .B(n22), .S(n1533), .Z(n30) );
  MUX2_X1 U1182 ( .A(n30), .B(n15), .S(N14), .Z(N30) );
  MUX2_X1 U1183 ( .A(\mem[30][1] ), .B(\mem[31][1] ), .S(n1545), .Z(n31) );
  MUX2_X1 U1184 ( .A(\mem[28][1] ), .B(\mem[29][1] ), .S(n1545), .Z(n32) );
  MUX2_X1 U1185 ( .A(n32), .B(n31), .S(N11), .Z(n33) );
  MUX2_X1 U1186 ( .A(\mem[26][1] ), .B(\mem[27][1] ), .S(n1545), .Z(n34) );
  MUX2_X1 U1187 ( .A(\mem[24][1] ), .B(\mem[25][1] ), .S(n1550), .Z(n35) );
  MUX2_X1 U1188 ( .A(n35), .B(n34), .S(N11), .Z(n36) );
  MUX2_X1 U1189 ( .A(n36), .B(n33), .S(n1535), .Z(n37) );
  MUX2_X1 U1190 ( .A(\mem[22][1] ), .B(\mem[23][1] ), .S(n1551), .Z(n1090) );
  MUX2_X1 U1191 ( .A(\mem[20][1] ), .B(\mem[21][1] ), .S(n1551), .Z(n1091) );
  MUX2_X1 U1192 ( .A(n1091), .B(n1090), .S(N11), .Z(n1092) );
  MUX2_X1 U1193 ( .A(\mem[18][1] ), .B(\mem[19][1] ), .S(n1551), .Z(n1093) );
  MUX2_X1 U1194 ( .A(\mem[16][1] ), .B(\mem[17][1] ), .S(n1548), .Z(n1094) );
  MUX2_X1 U1195 ( .A(n1094), .B(n1093), .S(n1542), .Z(n1095) );
  MUX2_X1 U1196 ( .A(n1095), .B(n1092), .S(n1535), .Z(n1096) );
  MUX2_X1 U1197 ( .A(n1096), .B(n37), .S(n1533), .Z(n1097) );
  MUX2_X1 U1198 ( .A(\mem[14][1] ), .B(\mem[15][1] ), .S(n1545), .Z(n1098) );
  MUX2_X1 U1199 ( .A(\mem[12][1] ), .B(\mem[13][1] ), .S(n1549), .Z(n1099) );
  MUX2_X1 U1200 ( .A(n1099), .B(n1098), .S(n1542), .Z(n1100) );
  MUX2_X1 U1201 ( .A(\mem[10][1] ), .B(\mem[11][1] ), .S(n1553), .Z(n1101) );
  MUX2_X1 U1202 ( .A(\mem[8][1] ), .B(\mem[9][1] ), .S(n1548), .Z(n1102) );
  MUX2_X1 U1203 ( .A(n1102), .B(n1101), .S(N11), .Z(n1103) );
  MUX2_X1 U1204 ( .A(n1103), .B(n1100), .S(n1535), .Z(n1104) );
  MUX2_X1 U1205 ( .A(\mem[6][1] ), .B(\mem[7][1] ), .S(n1543), .Z(n1105) );
  MUX2_X1 U1206 ( .A(\mem[4][1] ), .B(\mem[5][1] ), .S(n1548), .Z(n1106) );
  MUX2_X1 U1207 ( .A(n1106), .B(n1105), .S(N11), .Z(n1107) );
  MUX2_X1 U1208 ( .A(\mem[2][1] ), .B(\mem[3][1] ), .S(n1546), .Z(n1108) );
  MUX2_X1 U1209 ( .A(\mem[0][1] ), .B(\mem[1][1] ), .S(n1553), .Z(n1109) );
  MUX2_X1 U1210 ( .A(n1109), .B(n1108), .S(N11), .Z(n1110) );
  MUX2_X1 U1211 ( .A(n1110), .B(n1107), .S(n1535), .Z(n1111) );
  MUX2_X1 U1212 ( .A(n1111), .B(n1104), .S(N13), .Z(n1112) );
  MUX2_X1 U1213 ( .A(n1112), .B(n1097), .S(N14), .Z(N29) );
  MUX2_X1 U1214 ( .A(\mem[30][2] ), .B(\mem[31][2] ), .S(n1543), .Z(n1113) );
  MUX2_X1 U1215 ( .A(\mem[28][2] ), .B(\mem[29][2] ), .S(n1551), .Z(n1114) );
  MUX2_X1 U1216 ( .A(n1114), .B(n1113), .S(n1542), .Z(n1115) );
  MUX2_X1 U1217 ( .A(\mem[26][2] ), .B(\mem[27][2] ), .S(n1549), .Z(n1116) );
  MUX2_X1 U1218 ( .A(\mem[24][2] ), .B(\mem[25][2] ), .S(n1553), .Z(n1117) );
  MUX2_X1 U1219 ( .A(n1117), .B(n1116), .S(n1542), .Z(n1118) );
  MUX2_X1 U1220 ( .A(n1118), .B(n1115), .S(n1535), .Z(n1119) );
  MUX2_X1 U1221 ( .A(\mem[22][2] ), .B(\mem[23][2] ), .S(n1546), .Z(n1120) );
  MUX2_X1 U1222 ( .A(\mem[20][2] ), .B(\mem[21][2] ), .S(n1548), .Z(n1121) );
  MUX2_X1 U1223 ( .A(n1121), .B(n1120), .S(N11), .Z(n1122) );
  MUX2_X1 U1224 ( .A(\mem[18][2] ), .B(\mem[19][2] ), .S(n1553), .Z(n1123) );
  MUX2_X1 U1225 ( .A(\mem[16][2] ), .B(\mem[17][2] ), .S(n1553), .Z(n1124) );
  MUX2_X1 U1226 ( .A(n1124), .B(n1123), .S(N11), .Z(n1125) );
  MUX2_X1 U1227 ( .A(n1125), .B(n1122), .S(n1535), .Z(n1126) );
  MUX2_X1 U1228 ( .A(n1126), .B(n1119), .S(n1533), .Z(n1127) );
  MUX2_X1 U1229 ( .A(\mem[14][2] ), .B(\mem[15][2] ), .S(n1552), .Z(n1128) );
  MUX2_X1 U1230 ( .A(\mem[12][2] ), .B(\mem[13][2] ), .S(N10), .Z(n1129) );
  MUX2_X1 U1231 ( .A(n1129), .B(n1128), .S(n1537), .Z(n1130) );
  MUX2_X1 U1232 ( .A(\mem[10][2] ), .B(\mem[11][2] ), .S(N10), .Z(n1131) );
  MUX2_X1 U1233 ( .A(\mem[8][2] ), .B(\mem[9][2] ), .S(N10), .Z(n1132) );
  MUX2_X1 U1234 ( .A(n1132), .B(n1131), .S(n1542), .Z(n1133) );
  MUX2_X1 U1235 ( .A(n1133), .B(n1130), .S(n1535), .Z(n1134) );
  MUX2_X1 U1236 ( .A(\mem[6][2] ), .B(\mem[7][2] ), .S(N10), .Z(n1135) );
  MUX2_X1 U1237 ( .A(\mem[4][2] ), .B(\mem[5][2] ), .S(N10), .Z(n1136) );
  MUX2_X1 U1238 ( .A(n1136), .B(n1135), .S(n1542), .Z(n1137) );
  MUX2_X1 U1239 ( .A(\mem[2][2] ), .B(\mem[3][2] ), .S(N10), .Z(n1138) );
  MUX2_X1 U1240 ( .A(\mem[0][2] ), .B(\mem[1][2] ), .S(N10), .Z(n1139) );
  MUX2_X1 U1241 ( .A(n1139), .B(n1138), .S(n1542), .Z(n1140) );
  MUX2_X1 U1242 ( .A(n1140), .B(n1137), .S(n1535), .Z(n1141) );
  MUX2_X1 U1243 ( .A(n1141), .B(n1134), .S(n1533), .Z(n1142) );
  MUX2_X1 U1244 ( .A(n1142), .B(n1127), .S(N14), .Z(N28) );
  MUX2_X1 U1245 ( .A(\mem[30][3] ), .B(\mem[31][3] ), .S(n1552), .Z(n1143) );
  MUX2_X1 U1246 ( .A(\mem[28][3] ), .B(\mem[29][3] ), .S(N10), .Z(n1144) );
  MUX2_X1 U1247 ( .A(n1144), .B(n1143), .S(n1537), .Z(n1145) );
  MUX2_X1 U1248 ( .A(\mem[26][3] ), .B(\mem[27][3] ), .S(n1552), .Z(n1146) );
  MUX2_X1 U1249 ( .A(\mem[24][3] ), .B(\mem[25][3] ), .S(N10), .Z(n1147) );
  MUX2_X1 U1250 ( .A(n1147), .B(n1146), .S(N11), .Z(n1148) );
  MUX2_X1 U1251 ( .A(n1148), .B(n1145), .S(n1535), .Z(n1149) );
  MUX2_X1 U1252 ( .A(\mem[22][3] ), .B(\mem[23][3] ), .S(n1543), .Z(n1150) );
  MUX2_X1 U1253 ( .A(\mem[20][3] ), .B(\mem[21][3] ), .S(n1547), .Z(n1151) );
  MUX2_X1 U1254 ( .A(n1151), .B(n1150), .S(n1537), .Z(n1152) );
  MUX2_X1 U1255 ( .A(\mem[18][3] ), .B(\mem[19][3] ), .S(n1546), .Z(n1153) );
  MUX2_X1 U1256 ( .A(\mem[16][3] ), .B(\mem[17][3] ), .S(n1549), .Z(n1154) );
  MUX2_X1 U1257 ( .A(n1154), .B(n1153), .S(n1542), .Z(n1155) );
  MUX2_X1 U1258 ( .A(n1155), .B(n1152), .S(n1535), .Z(n1156) );
  MUX2_X1 U1259 ( .A(n1156), .B(n1149), .S(N13), .Z(n1157) );
  MUX2_X1 U1260 ( .A(\mem[14][3] ), .B(\mem[15][3] ), .S(n1543), .Z(n1158) );
  MUX2_X1 U1261 ( .A(\mem[12][3] ), .B(\mem[13][3] ), .S(n1549), .Z(n1159) );
  MUX2_X1 U1262 ( .A(n1159), .B(n1158), .S(N11), .Z(n1160) );
  MUX2_X1 U1263 ( .A(\mem[10][3] ), .B(\mem[11][3] ), .S(n1543), .Z(n1161) );
  MUX2_X1 U1264 ( .A(\mem[8][3] ), .B(\mem[9][3] ), .S(n1546), .Z(n1162) );
  MUX2_X1 U1265 ( .A(n1162), .B(n1161), .S(n1542), .Z(n1163) );
  MUX2_X1 U1266 ( .A(n1163), .B(n1160), .S(n1535), .Z(n1164) );
  MUX2_X1 U1267 ( .A(\mem[6][3] ), .B(\mem[7][3] ), .S(n1551), .Z(n1165) );
  MUX2_X1 U1268 ( .A(\mem[4][3] ), .B(\mem[5][3] ), .S(n1547), .Z(n1166) );
  MUX2_X1 U1269 ( .A(n1166), .B(n1165), .S(n1542), .Z(n1167) );
  MUX2_X1 U1270 ( .A(\mem[2][3] ), .B(\mem[3][3] ), .S(n1551), .Z(n1168) );
  MUX2_X1 U1271 ( .A(\mem[0][3] ), .B(\mem[1][3] ), .S(n1552), .Z(n1169) );
  MUX2_X1 U1272 ( .A(n1169), .B(n1168), .S(n1542), .Z(n1170) );
  MUX2_X1 U1273 ( .A(n1170), .B(n1167), .S(n1535), .Z(n1171) );
  MUX2_X1 U1274 ( .A(n1171), .B(n1164), .S(N13), .Z(n1172) );
  MUX2_X1 U1275 ( .A(n1172), .B(n1157), .S(N14), .Z(N27) );
  MUX2_X1 U1276 ( .A(\mem[30][4] ), .B(\mem[31][4] ), .S(n1545), .Z(n1173) );
  MUX2_X1 U1277 ( .A(\mem[28][4] ), .B(\mem[29][4] ), .S(n1545), .Z(n1174) );
  MUX2_X1 U1278 ( .A(n1174), .B(n1173), .S(n1538), .Z(n1175) );
  MUX2_X1 U1279 ( .A(\mem[26][4] ), .B(\mem[27][4] ), .S(n1545), .Z(n1176) );
  MUX2_X1 U1280 ( .A(\mem[24][4] ), .B(\mem[25][4] ), .S(n1548), .Z(n1177) );
  MUX2_X1 U1281 ( .A(n1177), .B(n1176), .S(n1538), .Z(n1178) );
  MUX2_X1 U1282 ( .A(n1178), .B(n1175), .S(n1534), .Z(n1179) );
  MUX2_X1 U1283 ( .A(\mem[22][4] ), .B(\mem[23][4] ), .S(n1545), .Z(n1180) );
  MUX2_X1 U1284 ( .A(\mem[20][4] ), .B(\mem[21][4] ), .S(n1547), .Z(n1181) );
  MUX2_X1 U1285 ( .A(n1181), .B(n1180), .S(n1538), .Z(n1182) );
  MUX2_X1 U1286 ( .A(\mem[18][4] ), .B(\mem[19][4] ), .S(n1547), .Z(n1183) );
  MUX2_X1 U1287 ( .A(\mem[16][4] ), .B(\mem[17][4] ), .S(n1550), .Z(n1184) );
  MUX2_X1 U1288 ( .A(n1184), .B(n1183), .S(n1538), .Z(n1185) );
  MUX2_X1 U1289 ( .A(n1185), .B(n1182), .S(n1534), .Z(n1186) );
  MUX2_X1 U1290 ( .A(n1186), .B(n1179), .S(n1533), .Z(n1187) );
  MUX2_X1 U1291 ( .A(\mem[14][4] ), .B(\mem[15][4] ), .S(n1545), .Z(n1188) );
  MUX2_X1 U1292 ( .A(\mem[12][4] ), .B(\mem[13][4] ), .S(n1550), .Z(n1189) );
  MUX2_X1 U1293 ( .A(n1189), .B(n1188), .S(n1538), .Z(n1190) );
  MUX2_X1 U1294 ( .A(\mem[10][4] ), .B(\mem[11][4] ), .S(n1549), .Z(n1191) );
  MUX2_X1 U1295 ( .A(\mem[8][4] ), .B(\mem[9][4] ), .S(n1550), .Z(n1192) );
  MUX2_X1 U1296 ( .A(n1192), .B(n1191), .S(n1538), .Z(n1193) );
  MUX2_X1 U1297 ( .A(n1193), .B(n1190), .S(n1534), .Z(n1194) );
  MUX2_X1 U1298 ( .A(\mem[6][4] ), .B(\mem[7][4] ), .S(n1552), .Z(n1195) );
  MUX2_X1 U1299 ( .A(\mem[4][4] ), .B(\mem[5][4] ), .S(n1552), .Z(n1196) );
  MUX2_X1 U1300 ( .A(n1196), .B(n1195), .S(n1538), .Z(n1197) );
  MUX2_X1 U1301 ( .A(\mem[2][4] ), .B(\mem[3][4] ), .S(n1553), .Z(n1198) );
  MUX2_X1 U1302 ( .A(\mem[0][4] ), .B(\mem[1][4] ), .S(n1552), .Z(n1199) );
  MUX2_X1 U1303 ( .A(n1199), .B(n1198), .S(n1538), .Z(n1200) );
  MUX2_X1 U1304 ( .A(n1200), .B(n1197), .S(n1536), .Z(n1201) );
  MUX2_X1 U1305 ( .A(n1201), .B(n1194), .S(n1533), .Z(n1202) );
  MUX2_X1 U1306 ( .A(n1202), .B(n1187), .S(N14), .Z(N26) );
  MUX2_X1 U1307 ( .A(\mem[30][5] ), .B(\mem[31][5] ), .S(n1543), .Z(n1203) );
  MUX2_X1 U1308 ( .A(\mem[28][5] ), .B(\mem[29][5] ), .S(n1552), .Z(n1204) );
  MUX2_X1 U1309 ( .A(n1204), .B(n1203), .S(n1538), .Z(n1205) );
  MUX2_X1 U1310 ( .A(\mem[26][5] ), .B(\mem[27][5] ), .S(n1553), .Z(n1206) );
  MUX2_X1 U1311 ( .A(\mem[24][5] ), .B(\mem[25][5] ), .S(n1552), .Z(n1207) );
  MUX2_X1 U1312 ( .A(n1207), .B(n1206), .S(n1538), .Z(n1208) );
  MUX2_X1 U1313 ( .A(n1208), .B(n1205), .S(n1534), .Z(n1209) );
  MUX2_X1 U1314 ( .A(\mem[22][5] ), .B(\mem[23][5] ), .S(n1546), .Z(n1210) );
  MUX2_X1 U1315 ( .A(\mem[20][5] ), .B(\mem[21][5] ), .S(n1553), .Z(n1211) );
  MUX2_X1 U1316 ( .A(n1211), .B(n1210), .S(n1538), .Z(n1212) );
  MUX2_X1 U1317 ( .A(\mem[18][5] ), .B(\mem[19][5] ), .S(n1549), .Z(n1213) );
  MUX2_X1 U1318 ( .A(\mem[16][5] ), .B(\mem[17][5] ), .S(n1553), .Z(n1214) );
  MUX2_X1 U1319 ( .A(n1214), .B(n1213), .S(n1538), .Z(n1215) );
  MUX2_X1 U1320 ( .A(n1215), .B(n1212), .S(n1534), .Z(n1216) );
  MUX2_X1 U1321 ( .A(n1216), .B(n1209), .S(n1533), .Z(n1217) );
  MUX2_X1 U1322 ( .A(\mem[14][5] ), .B(\mem[15][5] ), .S(n1543), .Z(n1218) );
  MUX2_X1 U1323 ( .A(\mem[12][5] ), .B(\mem[13][5] ), .S(n1552), .Z(n1219) );
  MUX2_X1 U1324 ( .A(n1219), .B(n1218), .S(n1539), .Z(n1220) );
  MUX2_X1 U1325 ( .A(\mem[10][5] ), .B(\mem[11][5] ), .S(n1549), .Z(n1221) );
  MUX2_X1 U1326 ( .A(\mem[8][5] ), .B(\mem[9][5] ), .S(n1551), .Z(n1222) );
  MUX2_X1 U1327 ( .A(n1222), .B(n1221), .S(n1539), .Z(n1223) );
  MUX2_X1 U1328 ( .A(n1223), .B(n1220), .S(n1534), .Z(n1224) );
  MUX2_X1 U1329 ( .A(\mem[6][5] ), .B(\mem[7][5] ), .S(n1552), .Z(n1225) );
  MUX2_X1 U1330 ( .A(\mem[4][5] ), .B(\mem[5][5] ), .S(n1552), .Z(n1226) );
  MUX2_X1 U1331 ( .A(n1226), .B(n1225), .S(n1539), .Z(n1227) );
  MUX2_X1 U1332 ( .A(\mem[2][5] ), .B(\mem[3][5] ), .S(n1549), .Z(n1228) );
  MUX2_X1 U1333 ( .A(\mem[0][5] ), .B(\mem[1][5] ), .S(n1552), .Z(n1229) );
  MUX2_X1 U1334 ( .A(n1229), .B(n1228), .S(n1539), .Z(n1230) );
  MUX2_X1 U1335 ( .A(n1230), .B(n1227), .S(n1536), .Z(n1231) );
  MUX2_X1 U1336 ( .A(n1231), .B(n1224), .S(n1533), .Z(n1232) );
  MUX2_X1 U1337 ( .A(n1232), .B(n1217), .S(N14), .Z(N25) );
  MUX2_X1 U1338 ( .A(\mem[30][6] ), .B(\mem[31][6] ), .S(n1552), .Z(n1233) );
  MUX2_X1 U1339 ( .A(\mem[28][6] ), .B(\mem[29][6] ), .S(n1552), .Z(n1234) );
  MUX2_X1 U1340 ( .A(n1234), .B(n1233), .S(n1539), .Z(n1235) );
  MUX2_X1 U1341 ( .A(\mem[26][6] ), .B(\mem[27][6] ), .S(n1552), .Z(n1236) );
  MUX2_X1 U1342 ( .A(\mem[24][6] ), .B(\mem[25][6] ), .S(n1547), .Z(n1237) );
  MUX2_X1 U1343 ( .A(n1237), .B(n1236), .S(n1539), .Z(n1238) );
  MUX2_X1 U1344 ( .A(n1238), .B(n1235), .S(n1534), .Z(n1239) );
  MUX2_X1 U1345 ( .A(\mem[22][6] ), .B(\mem[23][6] ), .S(n1552), .Z(n1240) );
  MUX2_X1 U1346 ( .A(\mem[20][6] ), .B(\mem[21][6] ), .S(N10), .Z(n1241) );
  MUX2_X1 U1347 ( .A(n1241), .B(n1240), .S(n1539), .Z(n1242) );
  MUX2_X1 U1348 ( .A(\mem[18][6] ), .B(\mem[19][6] ), .S(N10), .Z(n1243) );
  MUX2_X1 U1349 ( .A(\mem[16][6] ), .B(\mem[17][6] ), .S(n1552), .Z(n1244) );
  MUX2_X1 U1350 ( .A(n1244), .B(n1243), .S(n1539), .Z(n1245) );
  MUX2_X1 U1351 ( .A(n1245), .B(n1242), .S(n1535), .Z(n1246) );
  MUX2_X1 U1352 ( .A(n1246), .B(n1239), .S(n1533), .Z(n1247) );
  MUX2_X1 U1353 ( .A(\mem[14][6] ), .B(\mem[15][6] ), .S(n1552), .Z(n1248) );
  MUX2_X1 U1354 ( .A(\mem[12][6] ), .B(\mem[13][6] ), .S(N10), .Z(n1249) );
  MUX2_X1 U1355 ( .A(n1249), .B(n1248), .S(n1539), .Z(n1250) );
  MUX2_X1 U1356 ( .A(\mem[10][6] ), .B(\mem[11][6] ), .S(N10), .Z(n1251) );
  MUX2_X1 U1357 ( .A(\mem[8][6] ), .B(\mem[9][6] ), .S(n1553), .Z(n1252) );
  MUX2_X1 U1358 ( .A(n1252), .B(n1251), .S(n1539), .Z(n1253) );
  MUX2_X1 U1359 ( .A(n1253), .B(n1250), .S(n1534), .Z(n1254) );
  MUX2_X1 U1360 ( .A(\mem[6][6] ), .B(\mem[7][6] ), .S(n1552), .Z(n1255) );
  MUX2_X1 U1361 ( .A(\mem[4][6] ), .B(\mem[5][6] ), .S(n1553), .Z(n1256) );
  MUX2_X1 U1362 ( .A(n1256), .B(n1255), .S(n1539), .Z(n1257) );
  MUX2_X1 U1363 ( .A(\mem[2][6] ), .B(\mem[3][6] ), .S(n1552), .Z(n1258) );
  MUX2_X1 U1364 ( .A(\mem[0][6] ), .B(\mem[1][6] ), .S(n1552), .Z(n1259) );
  MUX2_X1 U1365 ( .A(n1259), .B(n1258), .S(n1539), .Z(n1260) );
  MUX2_X1 U1366 ( .A(n1260), .B(n1257), .S(n1534), .Z(n1261) );
  MUX2_X1 U1367 ( .A(n1261), .B(n1254), .S(n1533), .Z(n1262) );
  MUX2_X1 U1368 ( .A(n1262), .B(n1247), .S(N14), .Z(N24) );
  MUX2_X1 U1369 ( .A(\mem[30][7] ), .B(\mem[31][7] ), .S(n1543), .Z(n1263) );
  MUX2_X1 U1370 ( .A(\mem[28][7] ), .B(\mem[29][7] ), .S(n1543), .Z(n1264) );
  MUX2_X1 U1371 ( .A(n1264), .B(n1263), .S(n1538), .Z(n1265) );
  MUX2_X1 U1372 ( .A(\mem[26][7] ), .B(\mem[27][7] ), .S(n1543), .Z(n1266) );
  MUX2_X1 U1373 ( .A(\mem[24][7] ), .B(\mem[25][7] ), .S(n1543), .Z(n1267) );
  MUX2_X1 U1374 ( .A(n1267), .B(n1266), .S(n1538), .Z(n1268) );
  MUX2_X1 U1375 ( .A(n1268), .B(n1265), .S(n1534), .Z(n1269) );
  MUX2_X1 U1376 ( .A(\mem[22][7] ), .B(\mem[23][7] ), .S(n1543), .Z(n1270) );
  MUX2_X1 U1377 ( .A(\mem[20][7] ), .B(\mem[21][7] ), .S(n1543), .Z(n1271) );
  MUX2_X1 U1378 ( .A(n1271), .B(n1270), .S(n1538), .Z(n1272) );
  MUX2_X1 U1379 ( .A(\mem[18][7] ), .B(\mem[19][7] ), .S(n1543), .Z(n1273) );
  MUX2_X1 U1380 ( .A(\mem[16][7] ), .B(\mem[17][7] ), .S(n1543), .Z(n1274) );
  MUX2_X1 U1381 ( .A(n1274), .B(n1273), .S(n1537), .Z(n1275) );
  MUX2_X1 U1382 ( .A(n1275), .B(n1272), .S(n1536), .Z(n1276) );
  MUX2_X1 U1383 ( .A(n1276), .B(n1269), .S(n1533), .Z(n1277) );
  MUX2_X1 U1384 ( .A(\mem[14][7] ), .B(\mem[15][7] ), .S(n1543), .Z(n1278) );
  MUX2_X1 U1385 ( .A(\mem[12][7] ), .B(\mem[13][7] ), .S(n1543), .Z(n1279) );
  MUX2_X1 U1386 ( .A(n1279), .B(n1278), .S(n1537), .Z(n1280) );
  MUX2_X1 U1387 ( .A(\mem[10][7] ), .B(\mem[11][7] ), .S(n1543), .Z(n1281) );
  MUX2_X1 U1388 ( .A(\mem[8][7] ), .B(\mem[9][7] ), .S(n1543), .Z(n1282) );
  MUX2_X1 U1389 ( .A(n1282), .B(n1281), .S(n1542), .Z(n1283) );
  MUX2_X1 U1390 ( .A(n1283), .B(n1280), .S(n1535), .Z(n1284) );
  MUX2_X1 U1391 ( .A(\mem[6][7] ), .B(\mem[7][7] ), .S(n1550), .Z(n1285) );
  MUX2_X1 U1392 ( .A(\mem[4][7] ), .B(\mem[5][7] ), .S(n1544), .Z(n1286) );
  MUX2_X1 U1393 ( .A(n1286), .B(n1285), .S(n1537), .Z(n1287) );
  MUX2_X1 U1394 ( .A(\mem[2][7] ), .B(\mem[3][7] ), .S(n1544), .Z(n1288) );
  MUX2_X1 U1395 ( .A(\mem[0][7] ), .B(\mem[1][7] ), .S(n1544), .Z(n1289) );
  MUX2_X1 U1396 ( .A(n1289), .B(n1288), .S(n1542), .Z(n1290) );
  MUX2_X1 U1397 ( .A(n1290), .B(n1287), .S(n1535), .Z(n1291) );
  MUX2_X1 U1398 ( .A(n1291), .B(n1284), .S(n1533), .Z(n1292) );
  MUX2_X1 U1399 ( .A(n1292), .B(n1277), .S(N14), .Z(N23) );
  MUX2_X1 U1400 ( .A(\mem[30][8] ), .B(\mem[31][8] ), .S(n1548), .Z(n1293) );
  MUX2_X1 U1401 ( .A(\mem[28][8] ), .B(\mem[29][8] ), .S(n1548), .Z(n1294) );
  MUX2_X1 U1402 ( .A(n1294), .B(n1293), .S(n1537), .Z(n1295) );
  MUX2_X1 U1403 ( .A(\mem[26][8] ), .B(\mem[27][8] ), .S(n1548), .Z(n1296) );
  MUX2_X1 U1404 ( .A(\mem[24][8] ), .B(\mem[25][8] ), .S(n1544), .Z(n1297) );
  MUX2_X1 U1405 ( .A(n1297), .B(n1296), .S(n1539), .Z(n1298) );
  MUX2_X1 U1406 ( .A(n1298), .B(n1295), .S(n1536), .Z(n1299) );
  MUX2_X1 U1407 ( .A(\mem[22][8] ), .B(\mem[23][8] ), .S(n1548), .Z(n1300) );
  MUX2_X1 U1408 ( .A(\mem[20][8] ), .B(\mem[21][8] ), .S(n1544), .Z(n1301) );
  MUX2_X1 U1409 ( .A(n1301), .B(n1300), .S(n1539), .Z(n1302) );
  MUX2_X1 U1410 ( .A(\mem[18][8] ), .B(\mem[19][8] ), .S(n1550), .Z(n1303) );
  MUX2_X1 U1411 ( .A(\mem[16][8] ), .B(\mem[17][8] ), .S(n1544), .Z(n1304) );
  MUX2_X1 U1412 ( .A(n1304), .B(n1303), .S(n1537), .Z(n1305) );
  MUX2_X1 U1413 ( .A(n1305), .B(n1302), .S(n1534), .Z(n1306) );
  MUX2_X1 U1414 ( .A(n1306), .B(n1299), .S(n1533), .Z(n1307) );
  MUX2_X1 U1415 ( .A(\mem[14][8] ), .B(\mem[15][8] ), .S(n1544), .Z(n1308) );
  MUX2_X1 U1416 ( .A(\mem[12][8] ), .B(\mem[13][8] ), .S(n1544), .Z(n1309) );
  MUX2_X1 U1417 ( .A(n1309), .B(n1308), .S(n1539), .Z(n1310) );
  MUX2_X1 U1418 ( .A(\mem[10][8] ), .B(\mem[11][8] ), .S(n1544), .Z(n1311) );
  MUX2_X1 U1419 ( .A(\mem[8][8] ), .B(\mem[9][8] ), .S(n1544), .Z(n1312) );
  MUX2_X1 U1420 ( .A(n1312), .B(n1311), .S(n1539), .Z(n1313) );
  MUX2_X1 U1421 ( .A(n1313), .B(n1310), .S(n1534), .Z(n1314) );
  MUX2_X1 U1422 ( .A(\mem[6][8] ), .B(\mem[7][8] ), .S(n1544), .Z(n1315) );
  MUX2_X1 U1423 ( .A(\mem[4][8] ), .B(\mem[5][8] ), .S(n1544), .Z(n1316) );
  MUX2_X1 U1424 ( .A(n1316), .B(n1315), .S(n1539), .Z(n1317) );
  MUX2_X1 U1425 ( .A(\mem[2][8] ), .B(\mem[3][8] ), .S(n1544), .Z(n1318) );
  MUX2_X1 U1426 ( .A(\mem[0][8] ), .B(\mem[1][8] ), .S(n1544), .Z(n1319) );
  MUX2_X1 U1427 ( .A(n1319), .B(n1318), .S(n1537), .Z(n1320) );
  MUX2_X1 U1428 ( .A(n1320), .B(n1317), .S(n1536), .Z(n1321) );
  MUX2_X1 U1429 ( .A(n1321), .B(n1314), .S(n1533), .Z(n1322) );
  MUX2_X1 U1430 ( .A(n1322), .B(n1307), .S(N14), .Z(N22) );
  MUX2_X1 U1431 ( .A(\mem[30][9] ), .B(\mem[31][9] ), .S(n1544), .Z(n1323) );
  MUX2_X1 U1432 ( .A(\mem[28][9] ), .B(\mem[29][9] ), .S(n1544), .Z(n1324) );
  MUX2_X1 U1433 ( .A(n1324), .B(n1323), .S(n1539), .Z(n1325) );
  MUX2_X1 U1434 ( .A(\mem[26][9] ), .B(\mem[27][9] ), .S(n1544), .Z(n1326) );
  MUX2_X1 U1435 ( .A(\mem[24][9] ), .B(\mem[25][9] ), .S(n1544), .Z(n1327) );
  MUX2_X1 U1436 ( .A(n1327), .B(n1326), .S(n1537), .Z(n1328) );
  MUX2_X1 U1437 ( .A(n1328), .B(n1325), .S(n1536), .Z(n1329) );
  MUX2_X1 U1438 ( .A(\mem[22][9] ), .B(\mem[23][9] ), .S(n1545), .Z(n1330) );
  MUX2_X1 U1439 ( .A(\mem[20][9] ), .B(\mem[21][9] ), .S(n1550), .Z(n1331) );
  MUX2_X1 U1440 ( .A(n1331), .B(n1330), .S(n1537), .Z(n1332) );
  MUX2_X1 U1441 ( .A(\mem[18][9] ), .B(\mem[19][9] ), .S(n1544), .Z(n1333) );
  MUX2_X1 U1442 ( .A(\mem[16][9] ), .B(\mem[17][9] ), .S(n1550), .Z(n1334) );
  MUX2_X1 U1443 ( .A(n1334), .B(n1333), .S(n1537), .Z(n1335) );
  MUX2_X1 U1444 ( .A(n1335), .B(n1332), .S(n1534), .Z(n1336) );
  MUX2_X1 U1445 ( .A(n1336), .B(n1329), .S(n1533), .Z(n1337) );
  MUX2_X1 U1446 ( .A(\mem[14][9] ), .B(\mem[15][9] ), .S(n1543), .Z(n1338) );
  MUX2_X1 U1447 ( .A(\mem[12][9] ), .B(\mem[13][9] ), .S(n1544), .Z(n1339) );
  MUX2_X1 U1448 ( .A(n1339), .B(n1338), .S(n1538), .Z(n1340) );
  MUX2_X1 U1449 ( .A(\mem[10][9] ), .B(\mem[11][9] ), .S(n1548), .Z(n1341) );
  MUX2_X1 U1450 ( .A(\mem[8][9] ), .B(\mem[9][9] ), .S(n1546), .Z(n1342) );
  MUX2_X1 U1451 ( .A(n1342), .B(n1341), .S(n1538), .Z(n1343) );
  MUX2_X1 U1452 ( .A(n1343), .B(n1340), .S(n1535), .Z(n1344) );
  MUX2_X1 U1453 ( .A(\mem[6][9] ), .B(\mem[7][9] ), .S(n1550), .Z(n1345) );
  MUX2_X1 U1454 ( .A(\mem[4][9] ), .B(\mem[5][9] ), .S(n1545), .Z(n1346) );
  MUX2_X1 U1455 ( .A(n1346), .B(n1345), .S(n1538), .Z(n1347) );
  MUX2_X1 U1456 ( .A(\mem[2][9] ), .B(\mem[3][9] ), .S(n1543), .Z(n1348) );
  MUX2_X1 U1457 ( .A(\mem[0][9] ), .B(\mem[1][9] ), .S(n1548), .Z(n1349) );
  MUX2_X1 U1458 ( .A(n1349), .B(n1348), .S(n1539), .Z(n1350) );
  MUX2_X1 U1459 ( .A(n1350), .B(n1347), .S(n1535), .Z(n1351) );
  MUX2_X1 U1460 ( .A(n1351), .B(n1344), .S(n1533), .Z(n1352) );
  MUX2_X1 U1461 ( .A(n1352), .B(n1337), .S(N14), .Z(N21) );
  MUX2_X1 U1462 ( .A(\mem[30][10] ), .B(\mem[31][10] ), .S(n1546), .Z(n1353)
         );
  MUX2_X1 U1463 ( .A(\mem[28][10] ), .B(\mem[29][10] ), .S(n1547), .Z(n1354)
         );
  MUX2_X1 U1464 ( .A(n1354), .B(n1353), .S(n1538), .Z(n1355) );
  MUX2_X1 U1465 ( .A(\mem[26][10] ), .B(\mem[27][10] ), .S(n1553), .Z(n1356)
         );
  MUX2_X1 U1466 ( .A(\mem[24][10] ), .B(\mem[25][10] ), .S(n1549), .Z(n1357)
         );
  MUX2_X1 U1467 ( .A(n1357), .B(n1356), .S(n1538), .Z(n1358) );
  MUX2_X1 U1468 ( .A(n1358), .B(n1355), .S(n1536), .Z(n1359) );
  MUX2_X1 U1469 ( .A(\mem[22][10] ), .B(\mem[23][10] ), .S(n1553), .Z(n1360)
         );
  MUX2_X1 U1470 ( .A(\mem[20][10] ), .B(\mem[21][10] ), .S(n1551), .Z(n1361)
         );
  MUX2_X1 U1471 ( .A(n1361), .B(n1360), .S(n1538), .Z(n1362) );
  MUX2_X1 U1472 ( .A(\mem[18][10] ), .B(\mem[19][10] ), .S(n1553), .Z(n1363)
         );
  MUX2_X1 U1473 ( .A(\mem[16][10] ), .B(\mem[17][10] ), .S(n1550), .Z(n1364)
         );
  MUX2_X1 U1474 ( .A(n1364), .B(n1363), .S(n1538), .Z(n1365) );
  MUX2_X1 U1475 ( .A(n1365), .B(n1362), .S(n1534), .Z(n1366) );
  MUX2_X1 U1476 ( .A(n1366), .B(n1359), .S(n1533), .Z(n1367) );
  MUX2_X1 U1477 ( .A(\mem[14][10] ), .B(\mem[15][10] ), .S(n1551), .Z(n1368)
         );
  MUX2_X1 U1478 ( .A(\mem[12][10] ), .B(\mem[13][10] ), .S(n1547), .Z(n1369)
         );
  MUX2_X1 U1479 ( .A(n1369), .B(n1368), .S(n1537), .Z(n1370) );
  MUX2_X1 U1480 ( .A(\mem[10][10] ), .B(\mem[11][10] ), .S(n1546), .Z(n1371)
         );
  MUX2_X1 U1481 ( .A(\mem[8][10] ), .B(\mem[9][10] ), .S(n1546), .Z(n1372) );
  MUX2_X1 U1482 ( .A(n1372), .B(n1371), .S(n1537), .Z(n1373) );
  MUX2_X1 U1483 ( .A(n1373), .B(n1370), .S(n1534), .Z(n1374) );
  MUX2_X1 U1484 ( .A(\mem[6][10] ), .B(\mem[7][10] ), .S(n1545), .Z(n1375) );
  MUX2_X1 U1485 ( .A(\mem[4][10] ), .B(\mem[5][10] ), .S(n1545), .Z(n1376) );
  MUX2_X1 U1486 ( .A(n1376), .B(n1375), .S(n1537), .Z(n1377) );
  MUX2_X1 U1487 ( .A(\mem[2][10] ), .B(\mem[3][10] ), .S(n1545), .Z(n1378) );
  MUX2_X1 U1488 ( .A(\mem[0][10] ), .B(\mem[1][10] ), .S(n1545), .Z(n1379) );
  MUX2_X1 U1489 ( .A(n1379), .B(n1378), .S(n1538), .Z(n1380) );
  MUX2_X1 U1490 ( .A(n1380), .B(n1377), .S(n1534), .Z(n1381) );
  MUX2_X1 U1491 ( .A(n1381), .B(n1374), .S(N13), .Z(n1382) );
  MUX2_X1 U1492 ( .A(n1382), .B(n1367), .S(N14), .Z(N20) );
  MUX2_X1 U1493 ( .A(\mem[30][11] ), .B(\mem[31][11] ), .S(n1545), .Z(n1383)
         );
  MUX2_X1 U1494 ( .A(\mem[28][11] ), .B(\mem[29][11] ), .S(n1545), .Z(n1384)
         );
  MUX2_X1 U1495 ( .A(n1384), .B(n1383), .S(n1539), .Z(n1385) );
  MUX2_X1 U1496 ( .A(\mem[26][11] ), .B(\mem[27][11] ), .S(n1545), .Z(n1386)
         );
  MUX2_X1 U1497 ( .A(\mem[24][11] ), .B(\mem[25][11] ), .S(n1545), .Z(n1387)
         );
  MUX2_X1 U1498 ( .A(n1387), .B(n1386), .S(n1539), .Z(n1388) );
  MUX2_X1 U1499 ( .A(n1388), .B(n1385), .S(n1534), .Z(n1389) );
  MUX2_X1 U1500 ( .A(\mem[22][11] ), .B(\mem[23][11] ), .S(n1545), .Z(n1390)
         );
  MUX2_X1 U1501 ( .A(\mem[20][11] ), .B(\mem[21][11] ), .S(n1545), .Z(n1391)
         );
  MUX2_X1 U1502 ( .A(n1391), .B(n1390), .S(n1539), .Z(n1392) );
  MUX2_X1 U1503 ( .A(\mem[18][11] ), .B(\mem[19][11] ), .S(n1545), .Z(n1393)
         );
  MUX2_X1 U1504 ( .A(\mem[16][11] ), .B(\mem[17][11] ), .S(n1545), .Z(n1394)
         );
  MUX2_X1 U1505 ( .A(n1394), .B(n1393), .S(n1539), .Z(n1395) );
  MUX2_X1 U1506 ( .A(n1395), .B(n1392), .S(n1535), .Z(n1396) );
  MUX2_X1 U1507 ( .A(n1396), .B(n1389), .S(n1533), .Z(n1397) );
  MUX2_X1 U1508 ( .A(\mem[14][11] ), .B(\mem[15][11] ), .S(n1546), .Z(n1398)
         );
  MUX2_X1 U1509 ( .A(\mem[12][11] ), .B(\mem[13][11] ), .S(n1546), .Z(n1399)
         );
  MUX2_X1 U1510 ( .A(n1399), .B(n1398), .S(n1540), .Z(n1400) );
  MUX2_X1 U1511 ( .A(\mem[10][11] ), .B(\mem[11][11] ), .S(n1546), .Z(n1401)
         );
  MUX2_X1 U1512 ( .A(\mem[8][11] ), .B(\mem[9][11] ), .S(n1546), .Z(n1402) );
  MUX2_X1 U1513 ( .A(n1402), .B(n1401), .S(n1540), .Z(n1403) );
  MUX2_X1 U1514 ( .A(n1403), .B(n1400), .S(n1535), .Z(n1404) );
  MUX2_X1 U1515 ( .A(\mem[6][11] ), .B(\mem[7][11] ), .S(n1546), .Z(n1405) );
  MUX2_X1 U1516 ( .A(\mem[4][11] ), .B(\mem[5][11] ), .S(n1546), .Z(n1406) );
  MUX2_X1 U1517 ( .A(n1406), .B(n1405), .S(n1540), .Z(n1407) );
  MUX2_X1 U1518 ( .A(\mem[2][11] ), .B(\mem[3][11] ), .S(n1546), .Z(n1408) );
  MUX2_X1 U1519 ( .A(\mem[0][11] ), .B(\mem[1][11] ), .S(n1546), .Z(n1409) );
  MUX2_X1 U1520 ( .A(n1409), .B(n1408), .S(n1540), .Z(n1410) );
  MUX2_X1 U1521 ( .A(n1410), .B(n1407), .S(n1535), .Z(n1411) );
  MUX2_X1 U1522 ( .A(n1411), .B(n1404), .S(N13), .Z(n1412) );
  MUX2_X1 U1523 ( .A(n1412), .B(n1397), .S(N14), .Z(N19) );
  MUX2_X1 U1524 ( .A(\mem[30][12] ), .B(\mem[31][12] ), .S(n1546), .Z(n1413)
         );
  MUX2_X1 U1525 ( .A(\mem[28][12] ), .B(\mem[29][12] ), .S(n1546), .Z(n1414)
         );
  MUX2_X1 U1526 ( .A(n1414), .B(n1413), .S(n1540), .Z(n1415) );
  MUX2_X1 U1527 ( .A(\mem[26][12] ), .B(\mem[27][12] ), .S(n1546), .Z(n1416)
         );
  MUX2_X1 U1528 ( .A(\mem[24][12] ), .B(\mem[25][12] ), .S(n1546), .Z(n1417)
         );
  MUX2_X1 U1529 ( .A(n1417), .B(n1416), .S(n1540), .Z(n1418) );
  MUX2_X1 U1530 ( .A(n1418), .B(n1415), .S(n1535), .Z(n1419) );
  MUX2_X1 U1531 ( .A(\mem[22][12] ), .B(\mem[23][12] ), .S(n1547), .Z(n1420)
         );
  MUX2_X1 U1532 ( .A(\mem[20][12] ), .B(\mem[21][12] ), .S(n1547), .Z(n1421)
         );
  MUX2_X1 U1533 ( .A(n1421), .B(n1420), .S(n1540), .Z(n1422) );
  MUX2_X1 U1534 ( .A(\mem[18][12] ), .B(\mem[19][12] ), .S(n1547), .Z(n1423)
         );
  MUX2_X1 U1535 ( .A(\mem[16][12] ), .B(\mem[17][12] ), .S(n1547), .Z(n1424)
         );
  MUX2_X1 U1536 ( .A(n1424), .B(n1423), .S(n1540), .Z(n1425) );
  MUX2_X1 U1537 ( .A(n1425), .B(n1422), .S(n1536), .Z(n1426) );
  MUX2_X1 U1538 ( .A(n1426), .B(n1419), .S(n1533), .Z(n1427) );
  MUX2_X1 U1539 ( .A(\mem[14][12] ), .B(\mem[15][12] ), .S(n1547), .Z(n1428)
         );
  MUX2_X1 U1540 ( .A(\mem[12][12] ), .B(\mem[13][12] ), .S(n1547), .Z(n1429)
         );
  MUX2_X1 U1541 ( .A(n1429), .B(n1428), .S(n1540), .Z(n1430) );
  MUX2_X1 U1542 ( .A(\mem[10][12] ), .B(\mem[11][12] ), .S(n1547), .Z(n1431)
         );
  MUX2_X1 U1543 ( .A(\mem[8][12] ), .B(\mem[9][12] ), .S(n1547), .Z(n1432) );
  MUX2_X1 U1544 ( .A(n1432), .B(n1431), .S(n1540), .Z(n1433) );
  MUX2_X1 U1545 ( .A(n1433), .B(n1430), .S(n1536), .Z(n1434) );
  MUX2_X1 U1546 ( .A(\mem[6][12] ), .B(\mem[7][12] ), .S(n1547), .Z(n1435) );
  MUX2_X1 U1547 ( .A(\mem[4][12] ), .B(\mem[5][12] ), .S(n1547), .Z(n1436) );
  MUX2_X1 U1548 ( .A(n1436), .B(n1435), .S(n1540), .Z(n1437) );
  MUX2_X1 U1549 ( .A(\mem[2][12] ), .B(\mem[3][12] ), .S(n1547), .Z(n1438) );
  MUX2_X1 U1550 ( .A(\mem[0][12] ), .B(\mem[1][12] ), .S(n1547), .Z(n1439) );
  MUX2_X1 U1551 ( .A(n1439), .B(n1438), .S(n1540), .Z(n1440) );
  MUX2_X1 U1552 ( .A(n1440), .B(n1437), .S(n1536), .Z(n1441) );
  MUX2_X1 U1553 ( .A(n1441), .B(n1434), .S(N13), .Z(n1442) );
  MUX2_X1 U1554 ( .A(n1442), .B(n1427), .S(N14), .Z(N18) );
  MUX2_X1 U1555 ( .A(\mem[30][13] ), .B(\mem[31][13] ), .S(n1548), .Z(n1443)
         );
  MUX2_X1 U1556 ( .A(\mem[28][13] ), .B(\mem[29][13] ), .S(n1548), .Z(n1444)
         );
  MUX2_X1 U1557 ( .A(n1444), .B(n1443), .S(n1541), .Z(n1445) );
  MUX2_X1 U1558 ( .A(\mem[26][13] ), .B(\mem[27][13] ), .S(n1548), .Z(n1446)
         );
  MUX2_X1 U1559 ( .A(\mem[24][13] ), .B(\mem[25][13] ), .S(n1548), .Z(n1447)
         );
  MUX2_X1 U1560 ( .A(n1447), .B(n1446), .S(n1541), .Z(n1448) );
  MUX2_X1 U1561 ( .A(n1448), .B(n1445), .S(n1536), .Z(n1449) );
  MUX2_X1 U1562 ( .A(\mem[22][13] ), .B(\mem[23][13] ), .S(n1548), .Z(n1450)
         );
  MUX2_X1 U1563 ( .A(\mem[20][13] ), .B(\mem[21][13] ), .S(n1548), .Z(n1451)
         );
  MUX2_X1 U1564 ( .A(n1451), .B(n1450), .S(n1541), .Z(n1452) );
  MUX2_X1 U1565 ( .A(\mem[18][13] ), .B(\mem[19][13] ), .S(n1548), .Z(n1453)
         );
  MUX2_X1 U1566 ( .A(\mem[16][13] ), .B(\mem[17][13] ), .S(n1548), .Z(n1454)
         );
  MUX2_X1 U1567 ( .A(n1454), .B(n1453), .S(n1541), .Z(n1455) );
  MUX2_X1 U1568 ( .A(n1455), .B(n1452), .S(n1536), .Z(n1456) );
  MUX2_X1 U1569 ( .A(n1456), .B(n1449), .S(n1533), .Z(n1457) );
  MUX2_X1 U1570 ( .A(\mem[14][13] ), .B(\mem[15][13] ), .S(n1548), .Z(n1458)
         );
  MUX2_X1 U1571 ( .A(\mem[12][13] ), .B(\mem[13][13] ), .S(n1548), .Z(n1459)
         );
  MUX2_X1 U1572 ( .A(n1459), .B(n1458), .S(n1541), .Z(n1460) );
  MUX2_X1 U1573 ( .A(\mem[10][13] ), .B(\mem[11][13] ), .S(n1548), .Z(n1461)
         );
  MUX2_X1 U1574 ( .A(\mem[8][13] ), .B(\mem[9][13] ), .S(n1548), .Z(n1462) );
  MUX2_X1 U1575 ( .A(n1462), .B(n1461), .S(n1541), .Z(n1463) );
  MUX2_X1 U1576 ( .A(n1463), .B(n1460), .S(n1536), .Z(n1464) );
  MUX2_X1 U1577 ( .A(\mem[6][13] ), .B(\mem[7][13] ), .S(n1549), .Z(n1465) );
  MUX2_X1 U1578 ( .A(\mem[4][13] ), .B(\mem[5][13] ), .S(n1549), .Z(n1466) );
  MUX2_X1 U1579 ( .A(n1466), .B(n1465), .S(n1541), .Z(n1467) );
  MUX2_X1 U1580 ( .A(\mem[2][13] ), .B(\mem[3][13] ), .S(n1549), .Z(n1468) );
  MUX2_X1 U1581 ( .A(\mem[0][13] ), .B(\mem[1][13] ), .S(n1549), .Z(n1469) );
  MUX2_X1 U1582 ( .A(n1469), .B(n1468), .S(n1541), .Z(n1470) );
  MUX2_X1 U1583 ( .A(n1470), .B(n1467), .S(n1536), .Z(n1471) );
  MUX2_X1 U1584 ( .A(n1471), .B(n1464), .S(N13), .Z(n1472) );
  MUX2_X1 U1585 ( .A(n1472), .B(n1457), .S(N14), .Z(N17) );
  MUX2_X1 U1586 ( .A(\mem[30][14] ), .B(\mem[31][14] ), .S(n1549), .Z(n1473)
         );
  MUX2_X1 U1587 ( .A(\mem[28][14] ), .B(\mem[29][14] ), .S(n1549), .Z(n1474)
         );
  MUX2_X1 U1588 ( .A(n1474), .B(n1473), .S(n1541), .Z(n1475) );
  MUX2_X1 U1589 ( .A(\mem[26][14] ), .B(\mem[27][14] ), .S(n1549), .Z(n1476)
         );
  MUX2_X1 U1590 ( .A(\mem[24][14] ), .B(\mem[25][14] ), .S(n1549), .Z(n1477)
         );
  MUX2_X1 U1591 ( .A(n1477), .B(n1476), .S(n1541), .Z(n1478) );
  MUX2_X1 U1592 ( .A(n1478), .B(n1475), .S(n1536), .Z(n1479) );
  MUX2_X1 U1593 ( .A(\mem[22][14] ), .B(\mem[23][14] ), .S(n1549), .Z(n1480)
         );
  MUX2_X1 U1594 ( .A(\mem[20][14] ), .B(\mem[21][14] ), .S(n1549), .Z(n1481)
         );
  MUX2_X1 U1595 ( .A(n1481), .B(n1480), .S(n1541), .Z(n1482) );
  MUX2_X1 U1596 ( .A(\mem[18][14] ), .B(\mem[19][14] ), .S(n1549), .Z(n1483)
         );
  MUX2_X1 U1597 ( .A(\mem[16][14] ), .B(\mem[17][14] ), .S(n1549), .Z(n1484)
         );
  MUX2_X1 U1598 ( .A(n1484), .B(n1483), .S(n1541), .Z(n1485) );
  MUX2_X1 U1599 ( .A(n1485), .B(n1482), .S(n1536), .Z(n1486) );
  MUX2_X1 U1600 ( .A(n1486), .B(n1479), .S(n1533), .Z(n1487) );
  MUX2_X1 U1601 ( .A(\mem[14][14] ), .B(\mem[15][14] ), .S(n1550), .Z(n1488)
         );
  MUX2_X1 U1602 ( .A(\mem[12][14] ), .B(\mem[13][14] ), .S(n1550), .Z(n1489)
         );
  MUX2_X1 U1603 ( .A(n1489), .B(n1488), .S(n1542), .Z(n1490) );
  MUX2_X1 U1604 ( .A(\mem[10][14] ), .B(\mem[11][14] ), .S(n1550), .Z(n1491)
         );
  MUX2_X1 U1605 ( .A(\mem[8][14] ), .B(\mem[9][14] ), .S(n1550), .Z(n1492) );
  MUX2_X1 U1606 ( .A(n1492), .B(n1491), .S(n1542), .Z(n1493) );
  MUX2_X1 U1607 ( .A(n1493), .B(n1490), .S(n1536), .Z(n1494) );
  MUX2_X1 U1608 ( .A(\mem[6][14] ), .B(\mem[7][14] ), .S(n1550), .Z(n1495) );
  MUX2_X1 U1609 ( .A(\mem[4][14] ), .B(\mem[5][14] ), .S(n1550), .Z(n1496) );
  MUX2_X1 U1610 ( .A(n1496), .B(n1495), .S(n1542), .Z(n1497) );
  MUX2_X1 U1611 ( .A(\mem[2][14] ), .B(\mem[3][14] ), .S(n1550), .Z(n1498) );
  MUX2_X1 U1612 ( .A(\mem[0][14] ), .B(\mem[1][14] ), .S(n1550), .Z(n1499) );
  MUX2_X1 U1613 ( .A(n1499), .B(n1498), .S(n1541), .Z(n1500) );
  MUX2_X1 U1614 ( .A(n1500), .B(n1497), .S(n1536), .Z(n1501) );
  MUX2_X1 U1615 ( .A(n1501), .B(n1494), .S(N13), .Z(n1502) );
  MUX2_X1 U1616 ( .A(n1502), .B(n1487), .S(N14), .Z(N16) );
  MUX2_X1 U1617 ( .A(\mem[30][15] ), .B(\mem[31][15] ), .S(n1550), .Z(n1503)
         );
  MUX2_X1 U1618 ( .A(\mem[28][15] ), .B(\mem[29][15] ), .S(n1550), .Z(n1504)
         );
  MUX2_X1 U1619 ( .A(n1504), .B(n1503), .S(n1542), .Z(n1505) );
  MUX2_X1 U1620 ( .A(\mem[26][15] ), .B(\mem[27][15] ), .S(n1550), .Z(n1506)
         );
  MUX2_X1 U1621 ( .A(\mem[24][15] ), .B(\mem[25][15] ), .S(n1550), .Z(n1507)
         );
  MUX2_X1 U1622 ( .A(n1507), .B(n1506), .S(n1542), .Z(n1508) );
  MUX2_X1 U1623 ( .A(n1508), .B(n1505), .S(n1536), .Z(n1509) );
  MUX2_X1 U1624 ( .A(\mem[22][15] ), .B(\mem[23][15] ), .S(n1551), .Z(n1510)
         );
  MUX2_X1 U1625 ( .A(\mem[20][15] ), .B(\mem[21][15] ), .S(n1551), .Z(n1511)
         );
  MUX2_X1 U1626 ( .A(n1511), .B(n1510), .S(n1542), .Z(n1512) );
  MUX2_X1 U1627 ( .A(\mem[18][15] ), .B(\mem[19][15] ), .S(n1551), .Z(n1513)
         );
  MUX2_X1 U1628 ( .A(\mem[16][15] ), .B(\mem[17][15] ), .S(n1551), .Z(n1514)
         );
  MUX2_X1 U1629 ( .A(n1514), .B(n1513), .S(n1542), .Z(n1515) );
  MUX2_X1 U1630 ( .A(n1515), .B(n1512), .S(n1536), .Z(n1516) );
  MUX2_X1 U1631 ( .A(n1516), .B(n1509), .S(n1533), .Z(n1517) );
  MUX2_X1 U1632 ( .A(\mem[14][15] ), .B(\mem[15][15] ), .S(n1551), .Z(n1518)
         );
  MUX2_X1 U1633 ( .A(\mem[12][15] ), .B(\mem[13][15] ), .S(n1551), .Z(n1519)
         );
  MUX2_X1 U1634 ( .A(n1519), .B(n1518), .S(n1542), .Z(n1520) );
  MUX2_X1 U1635 ( .A(\mem[10][15] ), .B(\mem[11][15] ), .S(n1551), .Z(n1521)
         );
  MUX2_X1 U1636 ( .A(\mem[8][15] ), .B(\mem[9][15] ), .S(n1551), .Z(n1522) );
  MUX2_X1 U1637 ( .A(n1522), .B(n1521), .S(n1540), .Z(n1523) );
  MUX2_X1 U1638 ( .A(n1523), .B(n1520), .S(n1536), .Z(n1524) );
  MUX2_X1 U1639 ( .A(\mem[6][15] ), .B(\mem[7][15] ), .S(n1551), .Z(n1525) );
  MUX2_X1 U1640 ( .A(\mem[4][15] ), .B(\mem[5][15] ), .S(n1551), .Z(n1526) );
  MUX2_X1 U1641 ( .A(n1526), .B(n1525), .S(n1542), .Z(n1527) );
  MUX2_X1 U1642 ( .A(\mem[2][15] ), .B(\mem[3][15] ), .S(n1551), .Z(n1528) );
  MUX2_X1 U1643 ( .A(\mem[0][15] ), .B(\mem[1][15] ), .S(n1551), .Z(n1529) );
  MUX2_X1 U1644 ( .A(n1529), .B(n1528), .S(n1540), .Z(n1530) );
  MUX2_X1 U1645 ( .A(n1530), .B(n1527), .S(n1536), .Z(n1531) );
  MUX2_X1 U1646 ( .A(n1531), .B(n1524), .S(N13), .Z(n1532) );
  MUX2_X1 U1647 ( .A(n1532), .B(n1517), .S(N14), .Z(N15) );
  CLKBUF_X1 U1648 ( .A(N12), .Z(n1534) );
  CLKBUF_X1 U1649 ( .A(N12), .Z(n1535) );
  CLKBUF_X1 U1650 ( .A(N12), .Z(n1536) );
  CLKBUF_X1 U1651 ( .A(N11), .Z(n1537) );
  INV_X1 U1652 ( .A(N10), .ZN(n1601) );
  INV_X1 U1653 ( .A(N11), .ZN(n1602) );
  INV_X1 U1654 ( .A(N13), .ZN(n1603) );
  INV_X1 U1655 ( .A(N14), .ZN(n1604) );
endmodule


module datapath_DW_mult_tc_31 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333;

  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n278), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n277), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n281), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n280), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n282), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  CLKBUF_X1 U157 ( .A(a[3]), .Z(n206) );
  AND2_X1 U158 ( .A1(n95), .A2(n102), .ZN(n207) );
  XNOR2_X1 U159 ( .A(n275), .B(n15), .ZN(n208) );
  AND3_X1 U160 ( .A1(n229), .A2(n230), .A3(n231), .ZN(product[15]) );
  XNOR2_X1 U161 ( .A(n210), .B(n233), .ZN(product[5]) );
  XNOR2_X1 U162 ( .A(n50), .B(n53), .ZN(n210) );
  XNOR2_X1 U163 ( .A(n211), .B(n220), .ZN(product[4]) );
  XNOR2_X1 U164 ( .A(n54), .B(n207), .ZN(n211) );
  XOR2_X1 U165 ( .A(n17), .B(n274), .Z(n212) );
  XOR2_X1 U166 ( .A(n3), .B(n212), .Z(product[13]) );
  NAND2_X1 U167 ( .A1(n3), .A2(n17), .ZN(n213) );
  NAND2_X1 U168 ( .A1(n3), .A2(n274), .ZN(n214) );
  NAND2_X1 U169 ( .A1(n17), .A2(n274), .ZN(n215) );
  NAND3_X1 U170 ( .A1(n213), .A2(n214), .A3(n215), .ZN(n2) );
  XNOR2_X1 U171 ( .A(n2), .B(n208), .ZN(product[14]) );
  XOR2_X1 U172 ( .A(n33), .B(n28), .Z(n216) );
  XOR2_X1 U173 ( .A(n7), .B(n216), .Z(product[9]) );
  NAND2_X1 U174 ( .A1(n7), .A2(n33), .ZN(n217) );
  NAND2_X1 U175 ( .A1(n7), .A2(n28), .ZN(n218) );
  NAND2_X1 U176 ( .A1(n33), .A2(n28), .ZN(n219) );
  NAND3_X1 U177 ( .A1(n217), .A2(n218), .A3(n219), .ZN(n6) );
  CLKBUF_X1 U178 ( .A(n12), .Z(n220) );
  NAND3_X1 U179 ( .A1(n258), .A2(n257), .A3(n259), .ZN(n221) );
  NAND3_X1 U180 ( .A1(n225), .A2(n224), .A3(n226), .ZN(n222) );
  NAND2_X2 U181 ( .A1(n311), .A2(n330), .ZN(n313) );
  XOR2_X2 U182 ( .A(a[6]), .B(n279), .Z(n311) );
  XOR2_X1 U183 ( .A(n27), .B(n24), .Z(n223) );
  XOR2_X1 U184 ( .A(n6), .B(n223), .Z(product[10]) );
  NAND2_X1 U185 ( .A1(n6), .A2(n27), .ZN(n224) );
  NAND2_X1 U186 ( .A1(n6), .A2(n24), .ZN(n225) );
  NAND2_X1 U187 ( .A1(n27), .A2(n24), .ZN(n226) );
  NAND3_X1 U188 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n5) );
  NAND3_X1 U189 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n227) );
  NAND3_X1 U190 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n228) );
  CLKBUF_X1 U191 ( .A(b[1]), .Z(n264) );
  NAND2_X1 U192 ( .A1(n2), .A2(n275), .ZN(n229) );
  NAND2_X1 U193 ( .A1(n2), .A2(n15), .ZN(n230) );
  NAND2_X1 U194 ( .A1(n275), .A2(n15), .ZN(n231) );
  NAND3_X1 U195 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n232) );
  NAND3_X1 U196 ( .A1(n235), .A2(n237), .A3(n236), .ZN(n233) );
  NAND3_X1 U197 ( .A1(n240), .A2(n239), .A3(n238), .ZN(n234) );
  NAND2_X1 U198 ( .A1(n54), .A2(n207), .ZN(n235) );
  NAND2_X1 U199 ( .A1(n12), .A2(n54), .ZN(n236) );
  NAND2_X1 U200 ( .A1(n207), .A2(n12), .ZN(n237) );
  NAND3_X1 U201 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n11) );
  NAND2_X1 U202 ( .A1(n50), .A2(n53), .ZN(n238) );
  NAND2_X1 U203 ( .A1(n232), .A2(n50), .ZN(n239) );
  NAND2_X1 U204 ( .A1(n53), .A2(n11), .ZN(n240) );
  NAND3_X1 U205 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n10) );
  NAND3_X1 U206 ( .A1(n258), .A2(n257), .A3(n259), .ZN(n241) );
  NAND3_X1 U207 ( .A1(n250), .A2(n249), .A3(n251), .ZN(n242) );
  XOR2_X1 U208 ( .A(n34), .B(n39), .Z(n243) );
  XOR2_X1 U209 ( .A(n228), .B(n243), .Z(product[8]) );
  NAND2_X1 U210 ( .A1(n227), .A2(n34), .ZN(n244) );
  NAND2_X1 U211 ( .A1(n8), .A2(n39), .ZN(n245) );
  NAND2_X1 U212 ( .A1(n34), .A2(n39), .ZN(n246) );
  NAND3_X1 U213 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n7) );
  XNOR2_X1 U214 ( .A(b[2]), .B(n272), .ZN(n247) );
  NAND2_X2 U215 ( .A1(n290), .A2(n328), .ZN(n292) );
  XOR2_X1 U216 ( .A(n46), .B(n49), .Z(n248) );
  XOR2_X1 U217 ( .A(n248), .B(n10), .Z(product[6]) );
  NAND2_X1 U218 ( .A1(n46), .A2(n49), .ZN(n249) );
  NAND2_X1 U219 ( .A1(n46), .A2(n234), .ZN(n250) );
  NAND2_X1 U220 ( .A1(n49), .A2(n234), .ZN(n251) );
  NAND3_X1 U221 ( .A1(n251), .A2(n250), .A3(n249), .ZN(n9) );
  XOR2_X1 U222 ( .A(n40), .B(n45), .Z(n252) );
  XOR2_X1 U223 ( .A(n252), .B(n9), .Z(product[7]) );
  NAND2_X1 U224 ( .A1(n40), .A2(n45), .ZN(n253) );
  NAND2_X1 U225 ( .A1(n40), .A2(n242), .ZN(n254) );
  NAND2_X1 U226 ( .A1(n45), .A2(n9), .ZN(n255) );
  NAND3_X1 U227 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n8) );
  XOR2_X1 U228 ( .A(n23), .B(n20), .Z(n256) );
  XOR2_X1 U229 ( .A(n222), .B(n256), .Z(product[11]) );
  NAND2_X1 U230 ( .A1(n5), .A2(n23), .ZN(n257) );
  NAND2_X1 U231 ( .A1(n222), .A2(n20), .ZN(n258) );
  NAND2_X1 U232 ( .A1(n23), .A2(n20), .ZN(n259) );
  NAND3_X1 U233 ( .A1(n258), .A2(n257), .A3(n259), .ZN(n4) );
  XOR2_X1 U234 ( .A(n18), .B(n19), .Z(n260) );
  XOR2_X1 U235 ( .A(n221), .B(n260), .Z(product[12]) );
  NAND2_X1 U236 ( .A1(n241), .A2(n18), .ZN(n261) );
  NAND2_X1 U237 ( .A1(n4), .A2(n19), .ZN(n262) );
  NAND2_X1 U238 ( .A1(n18), .A2(n19), .ZN(n263) );
  NAND3_X1 U239 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n3) );
  INV_X2 U240 ( .A(n271), .ZN(n272) );
  XOR2_X1 U241 ( .A(n95), .B(n102), .Z(n56) );
  CLKBUF_X1 U242 ( .A(b[0]), .Z(n265) );
  NAND2_X1 U243 ( .A1(a[4]), .A2(a[3]), .ZN(n268) );
  NAND2_X1 U244 ( .A1(n266), .A2(n267), .ZN(n269) );
  NAND2_X2 U245 ( .A1(n268), .A2(n269), .ZN(n300) );
  INV_X1 U246 ( .A(a[4]), .ZN(n266) );
  INV_X1 U247 ( .A(a[3]), .ZN(n267) );
  NAND2_X2 U248 ( .A1(n300), .A2(n329), .ZN(n302) );
  BUF_X1 U249 ( .A(n290), .Z(n270) );
  XOR2_X1 U250 ( .A(a[2]), .B(n283), .Z(n290) );
  INV_X1 U251 ( .A(n15), .ZN(n274) );
  INV_X1 U252 ( .A(n21), .ZN(n277) );
  INV_X1 U253 ( .A(n309), .ZN(n278) );
  INV_X1 U254 ( .A(n320), .ZN(n275) );
  INV_X1 U255 ( .A(b[0]), .ZN(n273) );
  INV_X1 U256 ( .A(n289), .ZN(n282) );
  INV_X1 U257 ( .A(n298), .ZN(n281) );
  INV_X1 U258 ( .A(n31), .ZN(n280) );
  INV_X1 U259 ( .A(a[0]), .ZN(n284) );
  INV_X1 U260 ( .A(a[5]), .ZN(n279) );
  INV_X1 U261 ( .A(a[7]), .ZN(n276) );
  INV_X1 U262 ( .A(a[1]), .ZN(n271) );
  INV_X1 U263 ( .A(a[1]), .ZN(n283) );
  NOR2_X1 U264 ( .A1(n284), .A2(n273), .ZN(product[0]) );
  OAI22_X1 U265 ( .A1(n285), .A2(n286), .B1(n287), .B2(n284), .ZN(n99) );
  OAI22_X1 U266 ( .A1(n287), .A2(n286), .B1(n288), .B2(n284), .ZN(n98) );
  XNOR2_X1 U267 ( .A(b[6]), .B(n272), .ZN(n287) );
  OAI22_X1 U268 ( .A1(n284), .A2(n288), .B1(n286), .B2(n288), .ZN(n289) );
  XNOR2_X1 U269 ( .A(b[7]), .B(n272), .ZN(n288) );
  NOR2_X1 U270 ( .A1(n290), .A2(n273), .ZN(n96) );
  OAI22_X1 U271 ( .A1(n291), .A2(n292), .B1(n293), .B2(n290), .ZN(n95) );
  XNOR2_X1 U272 ( .A(a[3]), .B(n265), .ZN(n291) );
  OAI22_X1 U273 ( .A1(n293), .A2(n292), .B1(n270), .B2(n294), .ZN(n94) );
  XNOR2_X1 U274 ( .A(n264), .B(a[3]), .ZN(n293) );
  OAI22_X1 U275 ( .A1(n294), .A2(n292), .B1(n270), .B2(n295), .ZN(n93) );
  XNOR2_X1 U276 ( .A(b[2]), .B(a[3]), .ZN(n294) );
  OAI22_X1 U277 ( .A1(n295), .A2(n292), .B1(n270), .B2(n296), .ZN(n92) );
  XNOR2_X1 U278 ( .A(b[3]), .B(n206), .ZN(n295) );
  OAI22_X1 U279 ( .A1(n296), .A2(n292), .B1(n270), .B2(n297), .ZN(n91) );
  XNOR2_X1 U280 ( .A(b[4]), .B(a[3]), .ZN(n296) );
  OAI22_X1 U281 ( .A1(n299), .A2(n270), .B1(n292), .B2(n299), .ZN(n298) );
  NOR2_X1 U282 ( .A1(n300), .A2(n273), .ZN(n88) );
  OAI22_X1 U283 ( .A1(n301), .A2(n302), .B1(n300), .B2(n303), .ZN(n87) );
  XNOR2_X1 U284 ( .A(a[5]), .B(n265), .ZN(n301) );
  OAI22_X1 U285 ( .A1(n303), .A2(n302), .B1(n300), .B2(n304), .ZN(n86) );
  XNOR2_X1 U286 ( .A(n264), .B(a[5]), .ZN(n303) );
  OAI22_X1 U287 ( .A1(n304), .A2(n302), .B1(n300), .B2(n305), .ZN(n85) );
  XNOR2_X1 U288 ( .A(b[2]), .B(a[5]), .ZN(n304) );
  OAI22_X1 U289 ( .A1(n305), .A2(n302), .B1(n300), .B2(n306), .ZN(n84) );
  XNOR2_X1 U290 ( .A(b[3]), .B(a[5]), .ZN(n305) );
  OAI22_X1 U291 ( .A1(n306), .A2(n302), .B1(n300), .B2(n307), .ZN(n83) );
  XNOR2_X1 U292 ( .A(b[4]), .B(a[5]), .ZN(n306) );
  OAI22_X1 U293 ( .A1(n307), .A2(n302), .B1(n300), .B2(n308), .ZN(n82) );
  XNOR2_X1 U294 ( .A(b[5]), .B(a[5]), .ZN(n307) );
  OAI22_X1 U295 ( .A1(n310), .A2(n300), .B1(n302), .B2(n310), .ZN(n309) );
  NOR2_X1 U296 ( .A1(n311), .A2(n273), .ZN(n80) );
  OAI22_X1 U297 ( .A1(n312), .A2(n313), .B1(n311), .B2(n314), .ZN(n79) );
  XNOR2_X1 U298 ( .A(a[7]), .B(n265), .ZN(n312) );
  OAI22_X1 U299 ( .A1(n315), .A2(n313), .B1(n311), .B2(n316), .ZN(n77) );
  OAI22_X1 U300 ( .A1(n316), .A2(n313), .B1(n311), .B2(n317), .ZN(n76) );
  XNOR2_X1 U301 ( .A(b[3]), .B(a[7]), .ZN(n316) );
  OAI22_X1 U302 ( .A1(n317), .A2(n313), .B1(n311), .B2(n318), .ZN(n75) );
  XNOR2_X1 U303 ( .A(b[4]), .B(a[7]), .ZN(n317) );
  OAI22_X1 U304 ( .A1(n318), .A2(n313), .B1(n311), .B2(n319), .ZN(n74) );
  XNOR2_X1 U305 ( .A(b[5]), .B(a[7]), .ZN(n318) );
  OAI22_X1 U306 ( .A1(n321), .A2(n311), .B1(n313), .B2(n321), .ZN(n320) );
  OAI21_X1 U307 ( .B1(n265), .B2(n283), .A(n286), .ZN(n72) );
  OAI21_X1 U308 ( .B1(n267), .B2(n292), .A(n322), .ZN(n71) );
  OR3_X1 U309 ( .A1(n270), .A2(n265), .A3(n267), .ZN(n322) );
  OAI21_X1 U310 ( .B1(n279), .B2(n302), .A(n323), .ZN(n70) );
  OR3_X1 U311 ( .A1(n300), .A2(n265), .A3(n279), .ZN(n323) );
  OAI21_X1 U312 ( .B1(n276), .B2(n313), .A(n324), .ZN(n69) );
  OR3_X1 U313 ( .A1(n311), .A2(n265), .A3(n276), .ZN(n324) );
  XNOR2_X1 U314 ( .A(n325), .B(n326), .ZN(n38) );
  OR2_X1 U315 ( .A1(n325), .A2(n326), .ZN(n37) );
  OAI22_X1 U316 ( .A1(n297), .A2(n292), .B1(n270), .B2(n327), .ZN(n326) );
  XNOR2_X1 U317 ( .A(b[5]), .B(n206), .ZN(n297) );
  OAI22_X1 U318 ( .A1(n314), .A2(n313), .B1(n311), .B2(n315), .ZN(n325) );
  XNOR2_X1 U319 ( .A(b[2]), .B(a[7]), .ZN(n315) );
  XNOR2_X1 U320 ( .A(n264), .B(a[7]), .ZN(n314) );
  OAI22_X1 U321 ( .A1(n327), .A2(n292), .B1(n270), .B2(n299), .ZN(n31) );
  XNOR2_X1 U322 ( .A(b[7]), .B(n206), .ZN(n299) );
  XNOR2_X1 U323 ( .A(n267), .B(a[2]), .ZN(n328) );
  XNOR2_X1 U324 ( .A(b[6]), .B(n206), .ZN(n327) );
  OAI22_X1 U325 ( .A1(n308), .A2(n302), .B1(n300), .B2(n310), .ZN(n21) );
  XNOR2_X1 U326 ( .A(b[7]), .B(a[5]), .ZN(n310) );
  XNOR2_X1 U327 ( .A(n279), .B(a[4]), .ZN(n329) );
  XNOR2_X1 U328 ( .A(b[6]), .B(a[5]), .ZN(n308) );
  OAI22_X1 U329 ( .A1(n319), .A2(n313), .B1(n311), .B2(n321), .ZN(n15) );
  XNOR2_X1 U330 ( .A(b[7]), .B(a[7]), .ZN(n321) );
  XNOR2_X1 U331 ( .A(n276), .B(a[6]), .ZN(n330) );
  XNOR2_X1 U332 ( .A(b[6]), .B(a[7]), .ZN(n319) );
  OAI22_X1 U333 ( .A1(n265), .A2(n286), .B1(n331), .B2(n284), .ZN(n104) );
  OAI22_X1 U334 ( .A1(n331), .A2(n286), .B1(n247), .B2(n284), .ZN(n103) );
  XNOR2_X1 U335 ( .A(b[1]), .B(n272), .ZN(n331) );
  OAI22_X1 U336 ( .A1(n247), .A2(n286), .B1(n332), .B2(n284), .ZN(n102) );
  OAI22_X1 U337 ( .A1(n332), .A2(n286), .B1(n333), .B2(n284), .ZN(n101) );
  XNOR2_X1 U338 ( .A(b[3]), .B(n272), .ZN(n332) );
  OAI22_X1 U339 ( .A1(n333), .A2(n286), .B1(n285), .B2(n284), .ZN(n100) );
  XNOR2_X1 U340 ( .A(b[5]), .B(n272), .ZN(n285) );
  NAND2_X1 U341 ( .A1(a[1]), .A2(n284), .ZN(n286) );
  XNOR2_X1 U342 ( .A(b[4]), .B(n272), .ZN(n333) );
endmodule


module datapath_DW01_add_31 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n70;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n70), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(n59), .Z(n1) );
  NAND3_X1 U2 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n2) );
  NAND3_X1 U3 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n3) );
  CLKBUF_X1 U4 ( .A(B[3]), .Z(n4) );
  NAND3_X1 U5 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n5) );
  NAND3_X1 U6 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n6) );
  NAND3_X1 U7 ( .A1(n13), .A2(n14), .A3(n15), .ZN(n7) );
  NAND3_X1 U8 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n8) );
  NAND3_X1 U9 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n9) );
  NAND3_X1 U10 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n10) );
  NAND3_X1 U11 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n11) );
  XOR2_X1 U12 ( .A(B[8]), .B(A[8]), .Z(n12) );
  XOR2_X1 U13 ( .A(n5), .B(n12), .Z(SUM[8]) );
  NAND2_X1 U14 ( .A1(n5), .A2(B[8]), .ZN(n13) );
  NAND2_X1 U15 ( .A1(carry[8]), .A2(A[8]), .ZN(n14) );
  NAND2_X1 U16 ( .A1(B[8]), .A2(A[8]), .ZN(n15) );
  NAND3_X1 U17 ( .A1(n13), .A2(n14), .A3(n15), .ZN(carry[9]) );
  XOR2_X1 U18 ( .A(carry[2]), .B(A[2]), .Z(n16) );
  XOR2_X1 U19 ( .A(B[2]), .B(n16), .Z(SUM[2]) );
  NAND2_X1 U20 ( .A1(B[2]), .A2(carry[2]), .ZN(n17) );
  NAND2_X1 U21 ( .A1(B[2]), .A2(A[2]), .ZN(n18) );
  NAND2_X1 U22 ( .A1(carry[2]), .A2(A[2]), .ZN(n19) );
  NAND3_X1 U23 ( .A1(n17), .A2(n18), .A3(n19), .ZN(carry[3]) );
  XOR2_X1 U24 ( .A(B[6]), .B(A[6]), .Z(n20) );
  XOR2_X1 U25 ( .A(n9), .B(n20), .Z(SUM[6]) );
  NAND2_X1 U26 ( .A1(n8), .A2(B[6]), .ZN(n21) );
  NAND2_X1 U27 ( .A1(carry[6]), .A2(A[6]), .ZN(n22) );
  NAND2_X1 U28 ( .A1(B[6]), .A2(A[6]), .ZN(n23) );
  NAND3_X1 U29 ( .A1(n21), .A2(n22), .A3(n23), .ZN(carry[7]) );
  NAND3_X1 U30 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n24) );
  XOR2_X1 U31 ( .A(B[12]), .B(A[12]), .Z(n25) );
  XOR2_X1 U32 ( .A(carry[12]), .B(n25), .Z(SUM[12]) );
  NAND2_X1 U33 ( .A1(n24), .A2(B[12]), .ZN(n26) );
  NAND2_X1 U34 ( .A1(carry[12]), .A2(A[12]), .ZN(n27) );
  NAND2_X1 U35 ( .A1(B[12]), .A2(A[12]), .ZN(n28) );
  NAND3_X1 U36 ( .A1(n26), .A2(n27), .A3(n28), .ZN(carry[13]) );
  XOR2_X1 U37 ( .A(B[13]), .B(A[13]), .Z(n29) );
  XOR2_X1 U38 ( .A(n11), .B(n29), .Z(SUM[13]) );
  NAND2_X1 U39 ( .A1(B[13]), .A2(carry[13]), .ZN(n30) );
  NAND2_X1 U40 ( .A1(n10), .A2(A[13]), .ZN(n31) );
  NAND2_X1 U41 ( .A1(B[13]), .A2(A[13]), .ZN(n32) );
  NAND3_X1 U42 ( .A1(n30), .A2(n31), .A3(n32), .ZN(carry[14]) );
  CLKBUF_X1 U43 ( .A(n7), .Z(n33) );
  NAND3_X1 U44 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n34) );
  NAND3_X1 U45 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n35) );
  NAND3_X1 U46 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n36) );
  XOR2_X1 U47 ( .A(n4), .B(A[3]), .Z(n37) );
  XOR2_X1 U48 ( .A(carry[3]), .B(n37), .Z(SUM[3]) );
  NAND2_X1 U49 ( .A1(n3), .A2(B[3]), .ZN(n38) );
  NAND2_X1 U50 ( .A1(n2), .A2(A[3]), .ZN(n39) );
  NAND2_X1 U51 ( .A1(B[3]), .A2(A[3]), .ZN(n40) );
  NAND3_X1 U52 ( .A1(n38), .A2(n39), .A3(n40), .ZN(carry[4]) );
  NAND3_X1 U53 ( .A1(n63), .A2(n62), .A3(n61), .ZN(n41) );
  NAND3_X1 U54 ( .A1(n59), .A2(n58), .A3(n57), .ZN(n42) );
  NAND3_X1 U55 ( .A1(n57), .A2(n58), .A3(n1), .ZN(n43) );
  XOR2_X1 U56 ( .A(B[11]), .B(A[11]), .Z(n44) );
  XOR2_X1 U57 ( .A(n41), .B(n44), .Z(SUM[11]) );
  NAND2_X1 U58 ( .A1(n41), .A2(B[11]), .ZN(n45) );
  NAND2_X1 U59 ( .A1(carry[11]), .A2(A[11]), .ZN(n46) );
  NAND2_X1 U60 ( .A1(B[11]), .A2(A[11]), .ZN(n47) );
  NAND3_X1 U61 ( .A1(n45), .A2(n46), .A3(n47), .ZN(carry[12]) );
  XOR2_X1 U62 ( .A(B[4]), .B(A[4]), .Z(n48) );
  XOR2_X1 U63 ( .A(n36), .B(n48), .Z(SUM[4]) );
  NAND2_X1 U64 ( .A1(n35), .A2(B[4]), .ZN(n49) );
  NAND2_X1 U65 ( .A1(carry[4]), .A2(A[4]), .ZN(n50) );
  NAND2_X1 U66 ( .A1(B[4]), .A2(A[4]), .ZN(n51) );
  NAND3_X1 U67 ( .A1(n49), .A2(n50), .A3(n51), .ZN(carry[5]) );
  XOR2_X1 U68 ( .A(B[5]), .B(A[5]), .Z(n52) );
  XOR2_X1 U69 ( .A(n34), .B(n52), .Z(SUM[5]) );
  NAND2_X1 U70 ( .A1(n34), .A2(B[5]), .ZN(n53) );
  NAND2_X1 U71 ( .A1(carry[5]), .A2(A[5]), .ZN(n54) );
  NAND2_X1 U72 ( .A1(B[5]), .A2(A[5]), .ZN(n55) );
  NAND3_X1 U73 ( .A1(n53), .A2(n54), .A3(n55), .ZN(carry[6]) );
  XOR2_X1 U74 ( .A(A[9]), .B(B[9]), .Z(n56) );
  XOR2_X1 U75 ( .A(n56), .B(n33), .Z(SUM[9]) );
  NAND2_X1 U76 ( .A1(A[9]), .A2(B[9]), .ZN(n57) );
  NAND2_X1 U77 ( .A1(A[9]), .A2(carry[9]), .ZN(n58) );
  NAND2_X1 U78 ( .A1(B[9]), .A2(n7), .ZN(n59) );
  NAND3_X1 U79 ( .A1(n59), .A2(n58), .A3(n57), .ZN(carry[10]) );
  XOR2_X1 U80 ( .A(A[10]), .B(B[10]), .Z(n60) );
  XOR2_X1 U81 ( .A(n60), .B(n43), .Z(SUM[10]) );
  NAND2_X1 U82 ( .A1(A[10]), .A2(B[10]), .ZN(n61) );
  NAND2_X1 U83 ( .A1(A[10]), .A2(carry[10]), .ZN(n62) );
  NAND2_X1 U84 ( .A1(B[10]), .A2(n42), .ZN(n63) );
  NAND3_X1 U85 ( .A1(n63), .A2(n62), .A3(n61), .ZN(carry[11]) );
  XOR2_X1 U86 ( .A(B[7]), .B(A[7]), .Z(n64) );
  XOR2_X1 U87 ( .A(carry[7]), .B(n64), .Z(SUM[7]) );
  NAND2_X1 U88 ( .A1(n6), .A2(B[7]), .ZN(n65) );
  NAND2_X1 U89 ( .A1(carry[7]), .A2(A[7]), .ZN(n66) );
  NAND2_X1 U90 ( .A1(B[7]), .A2(A[7]), .ZN(n67) );
  NAND3_X1 U91 ( .A1(n65), .A2(n66), .A3(n67), .ZN(carry[8]) );
  XNOR2_X1 U92 ( .A(carry[15]), .B(n68), .ZN(SUM[15]) );
  XNOR2_X1 U93 ( .A(B[15]), .B(A[15]), .ZN(n68) );
  XOR2_X1 U94 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U95 ( .A1(B[0]), .A2(A[0]), .ZN(n70) );
endmodule


module datapath_DW_mult_tc_30 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331;

  FA_X1 U10 ( .A(n46), .B(n49), .CI(n10), .CO(n9), .S(product[6]) );
  FA_X1 U11 ( .A(n50), .B(n53), .CI(n11), .CO(n10), .S(product[5]) );
  FA_X1 U12 ( .A(n54), .B(n207), .CI(n12), .CO(n11), .S(product[4]) );
  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n274), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n273), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n277), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n276), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n279), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  CLKBUF_X3 U157 ( .A(a[1]), .Z(n206) );
  NAND2_X1 U158 ( .A1(n297), .A2(n326), .ZN(n299) );
  BUF_X1 U159 ( .A(n269), .Z(n224) );
  XNOR2_X1 U160 ( .A(n254), .B(n210), .ZN(product[10]) );
  AND2_X1 U161 ( .A1(n214), .A2(n225), .ZN(n207) );
  AND3_X1 U162 ( .A1(n259), .A2(n260), .A3(n261), .ZN(product[15]) );
  CLKBUF_X1 U163 ( .A(b[1]), .Z(n209) );
  AND3_X1 U164 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n213) );
  AND3_X1 U165 ( .A1(n253), .A2(n252), .A3(n251), .ZN(n210) );
  CLKBUF_X1 U166 ( .A(b[4]), .Z(n211) );
  NAND2_X2 U167 ( .A1(n308), .A2(n327), .ZN(n310) );
  XOR2_X2 U168 ( .A(a[6]), .B(n275), .Z(n308) );
  NAND3_X1 U169 ( .A1(n219), .A2(n218), .A3(n220), .ZN(n212) );
  XNOR2_X1 U170 ( .A(n213), .B(n258), .ZN(product[14]) );
  OAI22_X1 U171 ( .A1(n288), .A2(n289), .B1(n266), .B2(n290), .ZN(n214) );
  NAND3_X1 U172 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n215) );
  NAND3_X1 U173 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n216) );
  XOR2_X1 U174 ( .A(n23), .B(n20), .Z(n217) );
  XOR2_X1 U175 ( .A(n216), .B(n217), .Z(product[11]) );
  NAND2_X1 U176 ( .A1(n5), .A2(n23), .ZN(n218) );
  NAND2_X1 U177 ( .A1(n215), .A2(n20), .ZN(n219) );
  NAND2_X1 U178 ( .A1(n23), .A2(n20), .ZN(n220) );
  NAND3_X1 U179 ( .A1(n219), .A2(n218), .A3(n220), .ZN(n4) );
  NAND3_X1 U180 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n221) );
  NAND3_X1 U181 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n222) );
  NAND3_X1 U182 ( .A1(n231), .A2(n232), .A3(n233), .ZN(n223) );
  CLKBUF_X1 U183 ( .A(n102), .Z(n225) );
  XOR2_X1 U184 ( .A(n103), .B(n96), .Z(n226) );
  XOR2_X1 U185 ( .A(n226), .B(n14), .Z(product[2]) );
  NAND2_X1 U186 ( .A1(n14), .A2(n103), .ZN(n227) );
  NAND2_X1 U187 ( .A1(n14), .A2(n96), .ZN(n228) );
  NAND2_X1 U188 ( .A1(n103), .A2(n96), .ZN(n229) );
  NAND3_X1 U189 ( .A1(n227), .A2(n228), .A3(n229), .ZN(n13) );
  NAND2_X2 U190 ( .A1(n287), .A2(n325), .ZN(n289) );
  INV_X2 U191 ( .A(n269), .ZN(n268) );
  XOR2_X1 U192 ( .A(a[3]), .B(n269), .Z(n288) );
  XOR2_X1 U193 ( .A(n19), .B(n18), .Z(n230) );
  XOR2_X1 U194 ( .A(n230), .B(n4), .Z(product[12]) );
  NAND2_X1 U195 ( .A1(n19), .A2(n18), .ZN(n231) );
  NAND2_X1 U196 ( .A1(n19), .A2(n212), .ZN(n232) );
  NAND2_X1 U197 ( .A1(n18), .A2(n4), .ZN(n233) );
  NAND3_X1 U198 ( .A1(n231), .A2(n232), .A3(n233), .ZN(n3) );
  XOR2_X1 U199 ( .A(n17), .B(n270), .Z(n234) );
  XOR2_X1 U200 ( .A(n234), .B(n223), .Z(product[13]) );
  NAND2_X1 U201 ( .A1(n17), .A2(n270), .ZN(n235) );
  NAND2_X1 U202 ( .A1(n17), .A2(n3), .ZN(n236) );
  NAND2_X1 U203 ( .A1(n270), .A2(n3), .ZN(n237) );
  NAND3_X1 U204 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n238) );
  NAND3_X1 U205 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n239) );
  XOR2_X1 U206 ( .A(n95), .B(n102), .Z(n56) );
  XOR2_X1 U207 ( .A(n40), .B(n45), .Z(n240) );
  XOR2_X1 U208 ( .A(n9), .B(n240), .Z(product[7]) );
  NAND2_X1 U209 ( .A1(n9), .A2(n40), .ZN(n241) );
  NAND2_X1 U210 ( .A1(n9), .A2(n45), .ZN(n242) );
  NAND2_X1 U211 ( .A1(n40), .A2(n45), .ZN(n243) );
  NAND3_X1 U212 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n8) );
  NAND3_X1 U213 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n244) );
  XOR2_X1 U214 ( .A(n34), .B(n39), .Z(n245) );
  XOR2_X1 U215 ( .A(n239), .B(n245), .Z(product[8]) );
  NAND2_X1 U216 ( .A1(n238), .A2(n34), .ZN(n246) );
  NAND2_X1 U217 ( .A1(n8), .A2(n39), .ZN(n247) );
  NAND2_X1 U218 ( .A1(n34), .A2(n39), .ZN(n248) );
  NAND3_X1 U219 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n7) );
  NAND3_X1 U220 ( .A1(n253), .A2(n252), .A3(n251), .ZN(n249) );
  XOR2_X1 U221 ( .A(n28), .B(n33), .Z(n250) );
  XOR2_X1 U222 ( .A(n250), .B(n244), .Z(product[9]) );
  NAND2_X1 U223 ( .A1(n28), .A2(n33), .ZN(n251) );
  NAND2_X1 U224 ( .A1(n28), .A2(n7), .ZN(n252) );
  NAND2_X1 U225 ( .A1(n33), .A2(n7), .ZN(n253) );
  NAND3_X1 U226 ( .A1(n252), .A2(n251), .A3(n253), .ZN(n6) );
  XOR2_X1 U227 ( .A(n24), .B(n27), .Z(n254) );
  NAND2_X1 U228 ( .A1(n24), .A2(n27), .ZN(n255) );
  NAND2_X1 U229 ( .A1(n24), .A2(n249), .ZN(n256) );
  NAND2_X1 U230 ( .A1(n27), .A2(n6), .ZN(n257) );
  NAND3_X1 U231 ( .A1(n257), .A2(n256), .A3(n255), .ZN(n5) );
  XOR2_X1 U232 ( .A(n271), .B(n15), .Z(n258) );
  NAND2_X1 U233 ( .A1(n222), .A2(n271), .ZN(n259) );
  NAND2_X1 U234 ( .A1(n221), .A2(n15), .ZN(n260) );
  NAND2_X1 U235 ( .A1(n271), .A2(n15), .ZN(n261) );
  NAND2_X1 U236 ( .A1(a[4]), .A2(a[3]), .ZN(n264) );
  NAND2_X1 U237 ( .A1(n262), .A2(n263), .ZN(n265) );
  NAND2_X2 U238 ( .A1(n264), .A2(n265), .ZN(n297) );
  INV_X1 U239 ( .A(a[4]), .ZN(n262) );
  INV_X1 U240 ( .A(a[3]), .ZN(n263) );
  INV_X1 U241 ( .A(a[0]), .ZN(n281) );
  INV_X1 U242 ( .A(n15), .ZN(n270) );
  INV_X1 U243 ( .A(n21), .ZN(n273) );
  INV_X1 U244 ( .A(n306), .ZN(n274) );
  INV_X1 U245 ( .A(n317), .ZN(n271) );
  INV_X1 U246 ( .A(b[0]), .ZN(n269) );
  INV_X1 U247 ( .A(n286), .ZN(n279) );
  INV_X1 U248 ( .A(n295), .ZN(n277) );
  INV_X1 U249 ( .A(n31), .ZN(n276) );
  INV_X1 U250 ( .A(a[5]), .ZN(n275) );
  INV_X1 U251 ( .A(a[7]), .ZN(n272) );
  BUF_X1 U252 ( .A(n287), .Z(n266) );
  BUF_X1 U253 ( .A(n287), .Z(n267) );
  XNOR2_X1 U254 ( .A(a[2]), .B(n206), .ZN(n287) );
  INV_X1 U255 ( .A(a[3]), .ZN(n278) );
  INV_X1 U256 ( .A(n206), .ZN(n280) );
  NOR2_X1 U257 ( .A1(n281), .A2(n224), .ZN(product[0]) );
  OAI22_X1 U258 ( .A1(n282), .A2(n283), .B1(n284), .B2(n281), .ZN(n99) );
  OAI22_X1 U259 ( .A1(n284), .A2(n283), .B1(n285), .B2(n281), .ZN(n98) );
  XNOR2_X1 U260 ( .A(b[6]), .B(n206), .ZN(n284) );
  OAI22_X1 U261 ( .A1(n281), .A2(n285), .B1(n283), .B2(n285), .ZN(n286) );
  XNOR2_X1 U262 ( .A(b[7]), .B(n206), .ZN(n285) );
  NOR2_X1 U263 ( .A1(n267), .A2(n224), .ZN(n96) );
  OAI22_X1 U264 ( .A1(n288), .A2(n289), .B1(n266), .B2(n290), .ZN(n95) );
  OAI22_X1 U265 ( .A1(n290), .A2(n289), .B1(n266), .B2(n291), .ZN(n94) );
  XNOR2_X1 U266 ( .A(b[1]), .B(a[3]), .ZN(n290) );
  OAI22_X1 U267 ( .A1(n291), .A2(n289), .B1(n266), .B2(n292), .ZN(n93) );
  XNOR2_X1 U268 ( .A(b[2]), .B(a[3]), .ZN(n291) );
  OAI22_X1 U269 ( .A1(n292), .A2(n289), .B1(n267), .B2(n293), .ZN(n92) );
  XNOR2_X1 U270 ( .A(b[3]), .B(a[3]), .ZN(n292) );
  OAI22_X1 U271 ( .A1(n293), .A2(n289), .B1(n267), .B2(n294), .ZN(n91) );
  XNOR2_X1 U272 ( .A(n211), .B(a[3]), .ZN(n293) );
  OAI22_X1 U273 ( .A1(n296), .A2(n266), .B1(n289), .B2(n296), .ZN(n295) );
  NOR2_X1 U274 ( .A1(n297), .A2(n224), .ZN(n88) );
  OAI22_X1 U275 ( .A1(n298), .A2(n299), .B1(n297), .B2(n300), .ZN(n87) );
  XNOR2_X1 U276 ( .A(a[5]), .B(n268), .ZN(n298) );
  OAI22_X1 U277 ( .A1(n300), .A2(n299), .B1(n297), .B2(n301), .ZN(n86) );
  XNOR2_X1 U278 ( .A(n209), .B(a[5]), .ZN(n300) );
  OAI22_X1 U279 ( .A1(n301), .A2(n299), .B1(n297), .B2(n302), .ZN(n85) );
  XNOR2_X1 U280 ( .A(b[2]), .B(a[5]), .ZN(n301) );
  OAI22_X1 U281 ( .A1(n302), .A2(n299), .B1(n297), .B2(n303), .ZN(n84) );
  XNOR2_X1 U282 ( .A(b[3]), .B(a[5]), .ZN(n302) );
  OAI22_X1 U283 ( .A1(n303), .A2(n299), .B1(n297), .B2(n304), .ZN(n83) );
  XNOR2_X1 U284 ( .A(n211), .B(a[5]), .ZN(n303) );
  OAI22_X1 U285 ( .A1(n304), .A2(n299), .B1(n297), .B2(n305), .ZN(n82) );
  XNOR2_X1 U286 ( .A(b[5]), .B(a[5]), .ZN(n304) );
  OAI22_X1 U287 ( .A1(n307), .A2(n297), .B1(n299), .B2(n307), .ZN(n306) );
  NOR2_X1 U288 ( .A1(n308), .A2(n224), .ZN(n80) );
  OAI22_X1 U289 ( .A1(n309), .A2(n310), .B1(n308), .B2(n311), .ZN(n79) );
  XNOR2_X1 U290 ( .A(a[7]), .B(n268), .ZN(n309) );
  OAI22_X1 U291 ( .A1(n312), .A2(n310), .B1(n308), .B2(n313), .ZN(n77) );
  OAI22_X1 U292 ( .A1(n313), .A2(n310), .B1(n308), .B2(n314), .ZN(n76) );
  XNOR2_X1 U293 ( .A(b[3]), .B(a[7]), .ZN(n313) );
  OAI22_X1 U294 ( .A1(n314), .A2(n310), .B1(n308), .B2(n315), .ZN(n75) );
  XNOR2_X1 U295 ( .A(n211), .B(a[7]), .ZN(n314) );
  OAI22_X1 U296 ( .A1(n315), .A2(n310), .B1(n308), .B2(n316), .ZN(n74) );
  XNOR2_X1 U297 ( .A(b[5]), .B(a[7]), .ZN(n315) );
  OAI22_X1 U298 ( .A1(n318), .A2(n308), .B1(n310), .B2(n318), .ZN(n317) );
  OAI21_X1 U299 ( .B1(n268), .B2(n280), .A(n283), .ZN(n72) );
  OAI21_X1 U300 ( .B1(n278), .B2(n289), .A(n319), .ZN(n71) );
  OR3_X1 U301 ( .A1(n267), .A2(n268), .A3(n278), .ZN(n319) );
  OAI21_X1 U302 ( .B1(n275), .B2(n299), .A(n320), .ZN(n70) );
  OR3_X1 U303 ( .A1(n297), .A2(n268), .A3(n275), .ZN(n320) );
  OAI21_X1 U304 ( .B1(n272), .B2(n310), .A(n321), .ZN(n69) );
  OR3_X1 U305 ( .A1(n308), .A2(n268), .A3(n272), .ZN(n321) );
  XNOR2_X1 U306 ( .A(n322), .B(n323), .ZN(n38) );
  OR2_X1 U307 ( .A1(n322), .A2(n323), .ZN(n37) );
  OAI22_X1 U308 ( .A1(n294), .A2(n289), .B1(n267), .B2(n324), .ZN(n323) );
  XNOR2_X1 U309 ( .A(b[5]), .B(a[3]), .ZN(n294) );
  OAI22_X1 U310 ( .A1(n311), .A2(n310), .B1(n308), .B2(n312), .ZN(n322) );
  XNOR2_X1 U311 ( .A(b[2]), .B(a[7]), .ZN(n312) );
  XNOR2_X1 U312 ( .A(n209), .B(a[7]), .ZN(n311) );
  OAI22_X1 U313 ( .A1(n324), .A2(n289), .B1(n266), .B2(n296), .ZN(n31) );
  XNOR2_X1 U314 ( .A(b[7]), .B(a[3]), .ZN(n296) );
  XNOR2_X1 U315 ( .A(n278), .B(a[2]), .ZN(n325) );
  XNOR2_X1 U316 ( .A(b[6]), .B(a[3]), .ZN(n324) );
  OAI22_X1 U317 ( .A1(n305), .A2(n299), .B1(n297), .B2(n307), .ZN(n21) );
  XNOR2_X1 U318 ( .A(b[7]), .B(a[5]), .ZN(n307) );
  XNOR2_X1 U319 ( .A(n275), .B(a[4]), .ZN(n326) );
  XNOR2_X1 U320 ( .A(b[6]), .B(a[5]), .ZN(n305) );
  OAI22_X1 U321 ( .A1(n316), .A2(n310), .B1(n308), .B2(n318), .ZN(n15) );
  XNOR2_X1 U322 ( .A(b[7]), .B(a[7]), .ZN(n318) );
  XNOR2_X1 U323 ( .A(n272), .B(a[6]), .ZN(n327) );
  XNOR2_X1 U324 ( .A(b[6]), .B(a[7]), .ZN(n316) );
  OAI22_X1 U325 ( .A1(n268), .A2(n283), .B1(n328), .B2(n281), .ZN(n104) );
  OAI22_X1 U326 ( .A1(n328), .A2(n283), .B1(n329), .B2(n281), .ZN(n103) );
  XNOR2_X1 U327 ( .A(b[1]), .B(n206), .ZN(n328) );
  OAI22_X1 U328 ( .A1(n329), .A2(n283), .B1(n330), .B2(n281), .ZN(n102) );
  XNOR2_X1 U329 ( .A(b[2]), .B(n206), .ZN(n329) );
  OAI22_X1 U330 ( .A1(n330), .A2(n283), .B1(n331), .B2(n281), .ZN(n101) );
  XNOR2_X1 U331 ( .A(b[3]), .B(n206), .ZN(n330) );
  OAI22_X1 U332 ( .A1(n331), .A2(n283), .B1(n282), .B2(n281), .ZN(n100) );
  XNOR2_X1 U333 ( .A(b[5]), .B(n206), .ZN(n282) );
  NAND2_X1 U334 ( .A1(n206), .A2(n281), .ZN(n283) );
  XNOR2_X1 U335 ( .A(b[4]), .B(n206), .ZN(n331) );
endmodule


module datapath_DW01_add_30 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n70;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n70), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(B[13]), .Z(n1) );
  NAND3_X1 U2 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n2) );
  NAND3_X1 U3 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n3) );
  XOR2_X1 U4 ( .A(n3), .B(A[4]), .Z(n4) );
  XOR2_X1 U5 ( .A(B[4]), .B(n4), .Z(SUM[4]) );
  NAND2_X1 U6 ( .A1(B[4]), .A2(n2), .ZN(n5) );
  NAND2_X1 U7 ( .A1(B[4]), .A2(A[4]), .ZN(n6) );
  NAND2_X1 U8 ( .A1(carry[4]), .A2(A[4]), .ZN(n7) );
  NAND3_X1 U9 ( .A1(n5), .A2(n6), .A3(n7), .ZN(carry[5]) );
  CLKBUF_X1 U10 ( .A(n43), .Z(n8) );
  CLKBUF_X1 U11 ( .A(B[12]), .Z(n9) );
  CLKBUF_X1 U12 ( .A(n21), .Z(n10) );
  NAND3_X1 U13 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n11) );
  NAND3_X1 U14 ( .A1(n67), .A2(n68), .A3(n66), .ZN(n12) );
  XOR2_X1 U15 ( .A(B[5]), .B(A[5]), .Z(n13) );
  XOR2_X1 U16 ( .A(carry[5]), .B(n13), .Z(SUM[5]) );
  NAND2_X1 U17 ( .A1(carry[5]), .A2(B[5]), .ZN(n14) );
  NAND2_X1 U18 ( .A1(carry[5]), .A2(A[5]), .ZN(n15) );
  NAND2_X1 U19 ( .A1(B[5]), .A2(A[5]), .ZN(n16) );
  NAND3_X1 U20 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[6]) );
  CLKBUF_X1 U21 ( .A(carry[10]), .Z(n17) );
  NAND3_X1 U22 ( .A1(n26), .A2(n28), .A3(n27), .ZN(n18) );
  NAND3_X1 U23 ( .A1(n10), .A2(n22), .A3(n23), .ZN(n19) );
  XOR2_X1 U24 ( .A(B[10]), .B(A[10]), .Z(n20) );
  XOR2_X1 U25 ( .A(n17), .B(n20), .Z(SUM[10]) );
  NAND2_X1 U26 ( .A1(carry[10]), .A2(B[10]), .ZN(n21) );
  NAND2_X1 U27 ( .A1(n12), .A2(A[10]), .ZN(n22) );
  NAND2_X1 U28 ( .A1(B[10]), .A2(A[10]), .ZN(n23) );
  NAND3_X1 U29 ( .A1(n21), .A2(n22), .A3(n23), .ZN(carry[11]) );
  NAND3_X1 U30 ( .A1(n31), .A2(n32), .A3(n33), .ZN(n24) );
  XOR2_X1 U31 ( .A(n19), .B(A[11]), .Z(n25) );
  XOR2_X1 U32 ( .A(B[11]), .B(n25), .Z(SUM[11]) );
  NAND2_X1 U33 ( .A1(B[11]), .A2(n11), .ZN(n26) );
  NAND2_X1 U34 ( .A1(B[11]), .A2(A[11]), .ZN(n27) );
  NAND2_X1 U35 ( .A1(carry[11]), .A2(A[11]), .ZN(n28) );
  NAND3_X1 U36 ( .A1(n26), .A2(n28), .A3(n27), .ZN(carry[12]) );
  CLKBUF_X1 U37 ( .A(n64), .Z(n29) );
  XOR2_X1 U38 ( .A(B[6]), .B(A[6]), .Z(n30) );
  XOR2_X1 U39 ( .A(carry[6]), .B(n30), .Z(SUM[6]) );
  NAND2_X1 U40 ( .A1(carry[6]), .A2(B[6]), .ZN(n31) );
  NAND2_X1 U41 ( .A1(carry[6]), .A2(A[6]), .ZN(n32) );
  NAND2_X1 U42 ( .A1(B[6]), .A2(A[6]), .ZN(n33) );
  NAND3_X1 U43 ( .A1(n31), .A2(n32), .A3(n33), .ZN(carry[7]) );
  XOR2_X1 U44 ( .A(carry[2]), .B(A[2]), .Z(n34) );
  XOR2_X1 U45 ( .A(B[2]), .B(n34), .Z(SUM[2]) );
  NAND2_X1 U46 ( .A1(B[2]), .A2(carry[2]), .ZN(n35) );
  NAND2_X1 U47 ( .A1(B[2]), .A2(A[2]), .ZN(n36) );
  NAND2_X1 U48 ( .A1(carry[2]), .A2(A[2]), .ZN(n37) );
  NAND3_X1 U49 ( .A1(n35), .A2(n36), .A3(n37), .ZN(carry[3]) );
  NAND3_X1 U50 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n38) );
  CLKBUF_X1 U51 ( .A(n63), .Z(n39) );
  XOR2_X1 U52 ( .A(n9), .B(A[12]), .Z(n40) );
  XOR2_X1 U53 ( .A(n18), .B(n40), .Z(SUM[12]) );
  NAND2_X1 U54 ( .A1(n18), .A2(B[12]), .ZN(n41) );
  NAND2_X1 U55 ( .A1(carry[12]), .A2(A[12]), .ZN(n42) );
  NAND2_X1 U56 ( .A1(B[12]), .A2(A[12]), .ZN(n43) );
  NAND3_X1 U57 ( .A1(n41), .A2(n42), .A3(n8), .ZN(carry[13]) );
  NAND3_X1 U58 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n44) );
  NAND3_X1 U59 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n45) );
  XOR2_X1 U60 ( .A(carry[3]), .B(A[3]), .Z(n46) );
  XOR2_X1 U61 ( .A(B[3]), .B(n46), .Z(SUM[3]) );
  NAND2_X1 U62 ( .A1(carry[3]), .A2(B[3]), .ZN(n47) );
  NAND2_X1 U63 ( .A1(B[3]), .A2(A[3]), .ZN(n48) );
  NAND2_X1 U64 ( .A1(carry[3]), .A2(A[3]), .ZN(n49) );
  NAND3_X1 U65 ( .A1(n47), .A2(n48), .A3(n49), .ZN(carry[4]) );
  XNOR2_X1 U66 ( .A(carry[15]), .B(n50), .ZN(SUM[15]) );
  XNOR2_X1 U67 ( .A(B[15]), .B(A[15]), .ZN(n50) );
  XOR2_X1 U68 ( .A(n1), .B(A[13]), .Z(n51) );
  XOR2_X1 U69 ( .A(carry[13]), .B(n51), .Z(SUM[13]) );
  NAND2_X1 U70 ( .A1(n38), .A2(B[13]), .ZN(n52) );
  NAND2_X1 U71 ( .A1(n38), .A2(A[13]), .ZN(n53) );
  NAND2_X1 U72 ( .A1(B[13]), .A2(A[13]), .ZN(n54) );
  NAND3_X1 U73 ( .A1(n52), .A2(n53), .A3(n54), .ZN(carry[14]) );
  XOR2_X1 U74 ( .A(B[7]), .B(A[7]), .Z(n55) );
  XOR2_X1 U75 ( .A(carry[7]), .B(n55), .Z(SUM[7]) );
  NAND2_X1 U76 ( .A1(n24), .A2(B[7]), .ZN(n56) );
  NAND2_X1 U77 ( .A1(n24), .A2(A[7]), .ZN(n57) );
  NAND2_X1 U78 ( .A1(B[7]), .A2(A[7]), .ZN(n58) );
  NAND3_X1 U79 ( .A1(n56), .A2(n57), .A3(n58), .ZN(carry[8]) );
  NAND3_X1 U80 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n59) );
  NAND3_X1 U81 ( .A1(n62), .A2(n39), .A3(n29), .ZN(n60) );
  XOR2_X1 U82 ( .A(A[8]), .B(B[8]), .Z(n61) );
  XOR2_X1 U83 ( .A(n61), .B(n45), .Z(SUM[8]) );
  NAND2_X1 U84 ( .A1(A[8]), .A2(B[8]), .ZN(n62) );
  NAND2_X1 U85 ( .A1(A[8]), .A2(n44), .ZN(n63) );
  NAND2_X1 U86 ( .A1(B[8]), .A2(carry[8]), .ZN(n64) );
  NAND3_X1 U87 ( .A1(n62), .A2(n63), .A3(n64), .ZN(carry[9]) );
  XOR2_X1 U88 ( .A(A[9]), .B(B[9]), .Z(n65) );
  XOR2_X1 U89 ( .A(n65), .B(n60), .Z(SUM[9]) );
  NAND2_X1 U90 ( .A1(A[9]), .A2(B[9]), .ZN(n66) );
  NAND2_X1 U91 ( .A1(carry[9]), .A2(A[9]), .ZN(n67) );
  NAND2_X1 U92 ( .A1(B[9]), .A2(n59), .ZN(n68) );
  NAND3_X1 U93 ( .A1(n68), .A2(n67), .A3(n66), .ZN(carry[10]) );
  XOR2_X1 U94 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U95 ( .A1(B[0]), .A2(A[0]), .ZN(n70) );
endmodule


module datapath_DW_mult_tc_29 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329;

  FA_X1 U5 ( .A(n20), .B(n23), .CI(n5), .CO(n4), .S(product[11]) );
  FA_X1 U11 ( .A(n50), .B(n53), .CI(n11), .CO(n10), .S(product[5]) );
  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n272), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n271), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n275), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n274), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n277), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  NAND2_X1 U157 ( .A1(n295), .A2(n324), .ZN(n297) );
  NAND2_X2 U158 ( .A1(n306), .A2(n325), .ZN(n308) );
  INV_X1 U159 ( .A(n15), .ZN(n268) );
  AND2_X1 U160 ( .A1(n233), .A2(n102), .ZN(n206) );
  XNOR2_X1 U161 ( .A(n269), .B(n15), .ZN(n207) );
  AND3_X1 U162 ( .A1(n254), .A2(n255), .A3(n256), .ZN(product[15]) );
  INV_X1 U163 ( .A(n253), .ZN(n209) );
  XOR2_X1 U164 ( .A(n27), .B(n24), .Z(n210) );
  XOR2_X1 U165 ( .A(n6), .B(n210), .Z(product[10]) );
  NAND2_X1 U166 ( .A1(n6), .A2(n27), .ZN(n211) );
  NAND2_X1 U167 ( .A1(n6), .A2(n24), .ZN(n212) );
  NAND2_X1 U168 ( .A1(n27), .A2(n24), .ZN(n213) );
  NAND3_X1 U169 ( .A1(n211), .A2(n212), .A3(n213), .ZN(n5) );
  XOR2_X1 U170 ( .A(n54), .B(n206), .Z(n214) );
  XOR2_X1 U171 ( .A(n12), .B(n214), .Z(product[4]) );
  NAND2_X1 U172 ( .A1(n12), .A2(n54), .ZN(n215) );
  NAND2_X1 U173 ( .A1(n12), .A2(n206), .ZN(n216) );
  NAND2_X1 U174 ( .A1(n54), .A2(n206), .ZN(n217) );
  NAND3_X1 U175 ( .A1(n215), .A2(n216), .A3(n217), .ZN(n11) );
  NAND2_X1 U176 ( .A1(n9), .A2(n45), .ZN(n218) );
  CLKBUF_X1 U177 ( .A(n231), .Z(n219) );
  NAND3_X1 U178 ( .A1(n230), .A2(n231), .A3(n232), .ZN(n220) );
  NAND3_X1 U179 ( .A1(n230), .A2(n219), .A3(n232), .ZN(n221) );
  INV_X1 U180 ( .A(n278), .ZN(n222) );
  INV_X2 U181 ( .A(a[0]), .ZN(n279) );
  XOR2_X1 U182 ( .A(n18), .B(n19), .Z(n223) );
  XOR2_X1 U183 ( .A(n4), .B(n223), .Z(product[12]) );
  NAND2_X1 U184 ( .A1(n4), .A2(n18), .ZN(n224) );
  NAND2_X1 U185 ( .A1(n4), .A2(n19), .ZN(n225) );
  NAND2_X1 U186 ( .A1(n18), .A2(n19), .ZN(n226) );
  NAND3_X1 U187 ( .A1(n225), .A2(n224), .A3(n226), .ZN(n3) );
  NAND3_X1 U188 ( .A1(n235), .A2(n218), .A3(n237), .ZN(n227) );
  NAND3_X1 U189 ( .A1(n235), .A2(n218), .A3(n237), .ZN(n228) );
  XOR2_X1 U190 ( .A(n46), .B(n49), .Z(n229) );
  XOR2_X1 U191 ( .A(n10), .B(n229), .Z(product[6]) );
  NAND2_X1 U192 ( .A1(n10), .A2(n46), .ZN(n230) );
  NAND2_X1 U193 ( .A1(n10), .A2(n49), .ZN(n231) );
  NAND2_X1 U194 ( .A1(n46), .A2(n49), .ZN(n232) );
  NAND3_X1 U195 ( .A1(n230), .A2(n231), .A3(n232), .ZN(n9) );
  OAI22_X1 U196 ( .A1(n286), .A2(n287), .B1(n285), .B2(n288), .ZN(n233) );
  XOR2_X1 U197 ( .A(n40), .B(n45), .Z(n234) );
  XOR2_X1 U198 ( .A(n221), .B(n234), .Z(product[7]) );
  NAND2_X1 U199 ( .A1(n220), .A2(n40), .ZN(n235) );
  NAND2_X1 U200 ( .A1(n9), .A2(n45), .ZN(n236) );
  NAND2_X1 U201 ( .A1(n40), .A2(n45), .ZN(n237) );
  NAND3_X1 U202 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n8) );
  CLKBUF_X1 U203 ( .A(b[2]), .Z(n238) );
  NAND2_X1 U204 ( .A1(n264), .A2(n265), .ZN(n239) );
  XNOR2_X1 U205 ( .A(n2), .B(n207), .ZN(product[14]) );
  NAND2_X2 U206 ( .A1(n285), .A2(n323), .ZN(n287) );
  NAND3_X1 U207 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n240) );
  XOR2_X1 U208 ( .A(n95), .B(n102), .Z(n56) );
  XOR2_X1 U209 ( .A(n34), .B(n39), .Z(n241) );
  XOR2_X1 U210 ( .A(n241), .B(n228), .Z(product[8]) );
  NAND2_X1 U211 ( .A1(n34), .A2(n39), .ZN(n242) );
  NAND2_X1 U212 ( .A1(n34), .A2(n8), .ZN(n243) );
  NAND2_X1 U213 ( .A1(n39), .A2(n227), .ZN(n244) );
  NAND3_X1 U214 ( .A1(n244), .A2(n243), .A3(n242), .ZN(n7) );
  XOR2_X1 U215 ( .A(n28), .B(n33), .Z(n245) );
  XOR2_X1 U216 ( .A(n245), .B(n240), .Z(product[9]) );
  NAND2_X1 U217 ( .A1(n28), .A2(n33), .ZN(n246) );
  NAND2_X1 U218 ( .A1(n28), .A2(n7), .ZN(n247) );
  NAND2_X1 U219 ( .A1(n33), .A2(n7), .ZN(n248) );
  NAND3_X1 U220 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n6) );
  XOR2_X1 U221 ( .A(n17), .B(n268), .Z(n249) );
  XOR2_X1 U222 ( .A(n3), .B(n249), .Z(product[13]) );
  NAND2_X1 U223 ( .A1(n3), .A2(n17), .ZN(n250) );
  NAND2_X1 U224 ( .A1(n3), .A2(n268), .ZN(n251) );
  NAND2_X1 U225 ( .A1(n17), .A2(n268), .ZN(n252) );
  NAND3_X1 U226 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n2) );
  INV_X1 U227 ( .A(n267), .ZN(n253) );
  NAND2_X1 U228 ( .A1(n2), .A2(n269), .ZN(n254) );
  NAND2_X1 U229 ( .A1(n2), .A2(n15), .ZN(n255) );
  NAND2_X1 U230 ( .A1(n269), .A2(n15), .ZN(n256) );
  NAND2_X1 U231 ( .A1(a[4]), .A2(a[3]), .ZN(n259) );
  NAND2_X1 U232 ( .A1(n257), .A2(n258), .ZN(n260) );
  NAND2_X2 U233 ( .A1(n259), .A2(n260), .ZN(n295) );
  INV_X1 U234 ( .A(a[4]), .ZN(n257) );
  INV_X1 U235 ( .A(a[3]), .ZN(n258) );
  OR2_X1 U236 ( .A1(n326), .A2(n281), .ZN(n261) );
  OR2_X1 U237 ( .A1(n327), .A2(n279), .ZN(n262) );
  NAND2_X1 U238 ( .A1(n261), .A2(n262), .ZN(n103) );
  NAND2_X1 U239 ( .A1(n264), .A2(n265), .ZN(n285) );
  NAND2_X1 U240 ( .A1(a[2]), .A2(a[1]), .ZN(n264) );
  NAND2_X1 U241 ( .A1(n263), .A2(n278), .ZN(n265) );
  INV_X1 U242 ( .A(a[2]), .ZN(n263) );
  INV_X1 U243 ( .A(n21), .ZN(n271) );
  INV_X1 U244 ( .A(n304), .ZN(n272) );
  INV_X1 U245 ( .A(n315), .ZN(n269) );
  INV_X1 U246 ( .A(b[0]), .ZN(n267) );
  INV_X1 U247 ( .A(n284), .ZN(n277) );
  INV_X1 U248 ( .A(n293), .ZN(n275) );
  INV_X1 U249 ( .A(n31), .ZN(n274) );
  XOR2_X1 U250 ( .A(a[6]), .B(n273), .Z(n306) );
  INV_X1 U251 ( .A(a[5]), .ZN(n273) );
  INV_X1 U252 ( .A(a[7]), .ZN(n270) );
  INV_X1 U253 ( .A(a[3]), .ZN(n276) );
  INV_X1 U254 ( .A(a[1]), .ZN(n278) );
  INV_X1 U255 ( .A(n267), .ZN(n266) );
  NOR2_X1 U256 ( .A1(n279), .A2(n209), .ZN(product[0]) );
  OAI22_X1 U257 ( .A1(n280), .A2(n281), .B1(n282), .B2(n279), .ZN(n99) );
  OAI22_X1 U258 ( .A1(n282), .A2(n281), .B1(n283), .B2(n279), .ZN(n98) );
  XNOR2_X1 U259 ( .A(b[6]), .B(n222), .ZN(n282) );
  OAI22_X1 U260 ( .A1(n279), .A2(n283), .B1(n281), .B2(n283), .ZN(n284) );
  XNOR2_X1 U261 ( .A(b[7]), .B(n222), .ZN(n283) );
  NOR2_X1 U262 ( .A1(n239), .A2(n267), .ZN(n96) );
  OAI22_X1 U263 ( .A1(n286), .A2(n287), .B1(n285), .B2(n288), .ZN(n95) );
  XNOR2_X1 U264 ( .A(a[3]), .B(n266), .ZN(n286) );
  OAI22_X1 U265 ( .A1(n288), .A2(n287), .B1(n239), .B2(n289), .ZN(n94) );
  XNOR2_X1 U266 ( .A(b[1]), .B(a[3]), .ZN(n288) );
  OAI22_X1 U267 ( .A1(n289), .A2(n287), .B1(n239), .B2(n290), .ZN(n93) );
  XNOR2_X1 U268 ( .A(n238), .B(a[3]), .ZN(n289) );
  OAI22_X1 U269 ( .A1(n290), .A2(n287), .B1(n239), .B2(n291), .ZN(n92) );
  XNOR2_X1 U270 ( .A(b[3]), .B(a[3]), .ZN(n290) );
  OAI22_X1 U271 ( .A1(n291), .A2(n287), .B1(n239), .B2(n292), .ZN(n91) );
  XNOR2_X1 U272 ( .A(b[4]), .B(a[3]), .ZN(n291) );
  OAI22_X1 U273 ( .A1(n294), .A2(n239), .B1(n287), .B2(n294), .ZN(n293) );
  NOR2_X1 U274 ( .A1(n295), .A2(n267), .ZN(n88) );
  OAI22_X1 U275 ( .A1(n296), .A2(n297), .B1(n295), .B2(n298), .ZN(n87) );
  XNOR2_X1 U276 ( .A(a[5]), .B(n253), .ZN(n296) );
  OAI22_X1 U277 ( .A1(n298), .A2(n297), .B1(n295), .B2(n299), .ZN(n86) );
  XNOR2_X1 U278 ( .A(b[1]), .B(a[5]), .ZN(n298) );
  OAI22_X1 U279 ( .A1(n299), .A2(n297), .B1(n295), .B2(n300), .ZN(n85) );
  XNOR2_X1 U280 ( .A(n238), .B(a[5]), .ZN(n299) );
  OAI22_X1 U281 ( .A1(n300), .A2(n297), .B1(n295), .B2(n301), .ZN(n84) );
  XNOR2_X1 U282 ( .A(b[3]), .B(a[5]), .ZN(n300) );
  OAI22_X1 U283 ( .A1(n301), .A2(n297), .B1(n295), .B2(n302), .ZN(n83) );
  XNOR2_X1 U284 ( .A(b[4]), .B(a[5]), .ZN(n301) );
  OAI22_X1 U285 ( .A1(n302), .A2(n297), .B1(n295), .B2(n303), .ZN(n82) );
  XNOR2_X1 U286 ( .A(b[5]), .B(a[5]), .ZN(n302) );
  OAI22_X1 U287 ( .A1(n305), .A2(n295), .B1(n297), .B2(n305), .ZN(n304) );
  NOR2_X1 U288 ( .A1(n306), .A2(n209), .ZN(n80) );
  OAI22_X1 U289 ( .A1(n307), .A2(n308), .B1(n306), .B2(n309), .ZN(n79) );
  XNOR2_X1 U290 ( .A(a[7]), .B(n253), .ZN(n307) );
  OAI22_X1 U291 ( .A1(n310), .A2(n308), .B1(n306), .B2(n311), .ZN(n77) );
  OAI22_X1 U292 ( .A1(n311), .A2(n308), .B1(n306), .B2(n312), .ZN(n76) );
  XNOR2_X1 U293 ( .A(b[3]), .B(a[7]), .ZN(n311) );
  OAI22_X1 U294 ( .A1(n312), .A2(n308), .B1(n306), .B2(n313), .ZN(n75) );
  XNOR2_X1 U295 ( .A(b[4]), .B(a[7]), .ZN(n312) );
  OAI22_X1 U296 ( .A1(n313), .A2(n308), .B1(n306), .B2(n314), .ZN(n74) );
  XNOR2_X1 U297 ( .A(b[5]), .B(a[7]), .ZN(n313) );
  OAI22_X1 U298 ( .A1(n316), .A2(n306), .B1(n308), .B2(n316), .ZN(n315) );
  OAI21_X1 U299 ( .B1(n266), .B2(n278), .A(n281), .ZN(n72) );
  OAI21_X1 U300 ( .B1(n276), .B2(n287), .A(n317), .ZN(n71) );
  OR3_X1 U301 ( .A1(n285), .A2(n253), .A3(n276), .ZN(n317) );
  OAI21_X1 U302 ( .B1(n273), .B2(n297), .A(n318), .ZN(n70) );
  OR3_X1 U303 ( .A1(n295), .A2(n253), .A3(n273), .ZN(n318) );
  OAI21_X1 U304 ( .B1(n270), .B2(n308), .A(n319), .ZN(n69) );
  OR3_X1 U305 ( .A1(n306), .A2(n253), .A3(n270), .ZN(n319) );
  XNOR2_X1 U306 ( .A(n320), .B(n321), .ZN(n38) );
  OR2_X1 U307 ( .A1(n320), .A2(n321), .ZN(n37) );
  OAI22_X1 U308 ( .A1(n292), .A2(n287), .B1(n239), .B2(n322), .ZN(n321) );
  XNOR2_X1 U309 ( .A(b[5]), .B(a[3]), .ZN(n292) );
  OAI22_X1 U310 ( .A1(n309), .A2(n308), .B1(n306), .B2(n310), .ZN(n320) );
  XNOR2_X1 U311 ( .A(n238), .B(a[7]), .ZN(n310) );
  XNOR2_X1 U312 ( .A(b[1]), .B(a[7]), .ZN(n309) );
  OAI22_X1 U313 ( .A1(n322), .A2(n287), .B1(n239), .B2(n294), .ZN(n31) );
  XNOR2_X1 U314 ( .A(b[7]), .B(a[3]), .ZN(n294) );
  XNOR2_X1 U315 ( .A(n276), .B(a[2]), .ZN(n323) );
  XNOR2_X1 U316 ( .A(b[6]), .B(a[3]), .ZN(n322) );
  OAI22_X1 U317 ( .A1(n303), .A2(n297), .B1(n295), .B2(n305), .ZN(n21) );
  XNOR2_X1 U318 ( .A(b[7]), .B(a[5]), .ZN(n305) );
  XNOR2_X1 U319 ( .A(n273), .B(a[4]), .ZN(n324) );
  XNOR2_X1 U320 ( .A(b[6]), .B(a[5]), .ZN(n303) );
  OAI22_X1 U321 ( .A1(n314), .A2(n308), .B1(n306), .B2(n316), .ZN(n15) );
  XNOR2_X1 U322 ( .A(b[7]), .B(a[7]), .ZN(n316) );
  XNOR2_X1 U323 ( .A(n270), .B(a[6]), .ZN(n325) );
  XNOR2_X1 U324 ( .A(b[6]), .B(a[7]), .ZN(n314) );
  OAI22_X1 U325 ( .A1(n266), .A2(n281), .B1(n326), .B2(n279), .ZN(n104) );
  XNOR2_X1 U326 ( .A(b[1]), .B(a[1]), .ZN(n326) );
  OAI22_X1 U327 ( .A1(n281), .A2(n327), .B1(n328), .B2(n279), .ZN(n102) );
  XNOR2_X1 U328 ( .A(b[2]), .B(a[1]), .ZN(n327) );
  OAI22_X1 U329 ( .A1(n328), .A2(n281), .B1(n329), .B2(n279), .ZN(n101) );
  XNOR2_X1 U330 ( .A(b[3]), .B(n222), .ZN(n328) );
  OAI22_X1 U331 ( .A1(n329), .A2(n281), .B1(n280), .B2(n279), .ZN(n100) );
  XNOR2_X1 U332 ( .A(b[5]), .B(n222), .ZN(n280) );
  NAND2_X1 U333 ( .A1(a[1]), .A2(n279), .ZN(n281) );
  XNOR2_X1 U334 ( .A(b[4]), .B(n222), .ZN(n329) );
endmodule


module datapath_DW01_add_29 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n77;
  wire   [15:1] carry;

  FA_X1 U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n77), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(n51), .Z(n1) );
  CLKBUF_X1 U2 ( .A(n63), .Z(n2) );
  XOR2_X1 U3 ( .A(B[3]), .B(A[3]), .Z(n3) );
  XOR2_X1 U4 ( .A(carry[3]), .B(n3), .Z(SUM[3]) );
  NAND2_X1 U5 ( .A1(carry[3]), .A2(B[3]), .ZN(n4) );
  NAND2_X1 U6 ( .A1(carry[3]), .A2(A[3]), .ZN(n5) );
  NAND2_X1 U7 ( .A1(B[3]), .A2(A[3]), .ZN(n6) );
  NAND3_X1 U8 ( .A1(n4), .A2(n5), .A3(n6), .ZN(carry[4]) );
  CLKBUF_X1 U9 ( .A(n36), .Z(n7) );
  NAND3_X1 U10 ( .A1(n12), .A2(n13), .A3(n14), .ZN(n8) );
  CLKBUF_X1 U11 ( .A(n74), .Z(n9) );
  CLKBUF_X1 U12 ( .A(n71), .Z(n10) );
  XOR2_X1 U13 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR2_X1 U14 ( .A(carry[4]), .B(n11), .Z(SUM[4]) );
  NAND2_X1 U15 ( .A1(carry[4]), .A2(B[4]), .ZN(n12) );
  NAND2_X1 U16 ( .A1(carry[4]), .A2(A[4]), .ZN(n13) );
  NAND2_X1 U17 ( .A1(B[4]), .A2(A[4]), .ZN(n14) );
  NAND3_X1 U18 ( .A1(n12), .A2(n13), .A3(n14), .ZN(carry[5]) );
  NAND3_X1 U19 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n15) );
  NAND3_X1 U20 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n16) );
  CLKBUF_X1 U21 ( .A(B[11]), .Z(n17) );
  CLKBUF_X1 U22 ( .A(n62), .Z(n18) );
  CLKBUF_X1 U23 ( .A(n47), .Z(n19) );
  XOR2_X1 U24 ( .A(B[5]), .B(A[5]), .Z(n20) );
  XOR2_X1 U25 ( .A(n8), .B(n20), .Z(SUM[5]) );
  NAND2_X1 U26 ( .A1(n8), .A2(B[5]), .ZN(n21) );
  NAND2_X1 U27 ( .A1(carry[5]), .A2(A[5]), .ZN(n22) );
  NAND2_X1 U28 ( .A1(B[5]), .A2(A[5]), .ZN(n23) );
  NAND3_X1 U29 ( .A1(n21), .A2(n22), .A3(n23), .ZN(carry[6]) );
  CLKBUF_X1 U30 ( .A(n50), .Z(n24) );
  CLKBUF_X1 U31 ( .A(n46), .Z(n25) );
  XOR2_X1 U32 ( .A(B[6]), .B(A[6]), .Z(n26) );
  XOR2_X1 U33 ( .A(n16), .B(n26), .Z(SUM[6]) );
  NAND2_X1 U34 ( .A1(n16), .A2(B[6]), .ZN(n27) );
  NAND2_X1 U35 ( .A1(carry[6]), .A2(A[6]), .ZN(n28) );
  NAND2_X1 U36 ( .A1(B[6]), .A2(A[6]), .ZN(n29) );
  NAND3_X1 U37 ( .A1(n27), .A2(n28), .A3(n29), .ZN(carry[7]) );
  NAND3_X1 U38 ( .A1(n75), .A2(n74), .A3(n73), .ZN(n30) );
  NAND3_X1 U39 ( .A1(n75), .A2(n9), .A3(n73), .ZN(n31) );
  NAND3_X1 U40 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n32) );
  NAND3_X1 U41 ( .A1(n36), .A2(n37), .A3(n38), .ZN(n33) );
  NAND3_X1 U42 ( .A1(n7), .A2(n37), .A3(n38), .ZN(n34) );
  XOR2_X1 U43 ( .A(n31), .B(A[10]), .Z(n35) );
  XOR2_X1 U44 ( .A(B[10]), .B(n35), .Z(SUM[10]) );
  NAND2_X1 U45 ( .A1(B[10]), .A2(n30), .ZN(n36) );
  NAND2_X1 U46 ( .A1(B[10]), .A2(A[10]), .ZN(n37) );
  NAND2_X1 U47 ( .A1(carry[10]), .A2(A[10]), .ZN(n38) );
  NAND3_X1 U48 ( .A1(n38), .A2(n37), .A3(n36), .ZN(carry[11]) );
  NAND3_X1 U49 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n39) );
  NAND3_X1 U50 ( .A1(n49), .A2(n24), .A3(n1), .ZN(n40) );
  NAND3_X1 U51 ( .A1(n47), .A2(n46), .A3(n45), .ZN(n41) );
  NAND3_X1 U52 ( .A1(n45), .A2(n25), .A3(n19), .ZN(n42) );
  XNOR2_X1 U53 ( .A(n43), .B(n59), .ZN(SUM[14]) );
  XNOR2_X1 U54 ( .A(B[14]), .B(A[14]), .ZN(n43) );
  XOR2_X1 U55 ( .A(A[11]), .B(n17), .Z(n44) );
  XOR2_X1 U56 ( .A(n44), .B(n34), .Z(SUM[11]) );
  NAND2_X1 U57 ( .A1(A[11]), .A2(B[11]), .ZN(n45) );
  NAND2_X1 U58 ( .A1(A[11]), .A2(carry[11]), .ZN(n46) );
  NAND2_X1 U59 ( .A1(B[11]), .A2(n33), .ZN(n47) );
  NAND3_X1 U60 ( .A1(n46), .A2(n45), .A3(n47), .ZN(carry[12]) );
  XOR2_X1 U61 ( .A(A[12]), .B(B[12]), .Z(n48) );
  XOR2_X1 U62 ( .A(n48), .B(n42), .Z(SUM[12]) );
  NAND2_X1 U63 ( .A1(A[12]), .A2(B[12]), .ZN(n49) );
  NAND2_X1 U64 ( .A1(A[12]), .A2(n41), .ZN(n50) );
  NAND2_X1 U65 ( .A1(B[12]), .A2(carry[12]), .ZN(n51) );
  NAND3_X1 U66 ( .A1(n51), .A2(n50), .A3(n49), .ZN(carry[13]) );
  XOR2_X1 U67 ( .A(B[7]), .B(A[7]), .Z(n52) );
  XOR2_X1 U68 ( .A(carry[7]), .B(n52), .Z(SUM[7]) );
  NAND2_X1 U69 ( .A1(n15), .A2(B[7]), .ZN(n53) );
  NAND2_X1 U70 ( .A1(carry[7]), .A2(A[7]), .ZN(n54) );
  NAND2_X1 U71 ( .A1(B[7]), .A2(A[7]), .ZN(n55) );
  NAND3_X1 U72 ( .A1(n53), .A2(n54), .A3(n55), .ZN(carry[8]) );
  NAND3_X1 U73 ( .A1(n71), .A2(n70), .A3(n69), .ZN(n56) );
  NAND3_X1 U74 ( .A1(n69), .A2(n70), .A3(n10), .ZN(n57) );
  NAND3_X1 U75 ( .A1(n63), .A2(n62), .A3(n61), .ZN(n58) );
  NAND3_X1 U76 ( .A1(n61), .A2(n18), .A3(n2), .ZN(n59) );
  XOR2_X1 U77 ( .A(A[13]), .B(B[13]), .Z(n60) );
  XOR2_X1 U78 ( .A(n60), .B(n40), .Z(SUM[13]) );
  NAND2_X1 U79 ( .A1(A[13]), .A2(B[13]), .ZN(n61) );
  NAND2_X1 U80 ( .A1(A[13]), .A2(carry[13]), .ZN(n62) );
  NAND2_X1 U81 ( .A1(B[13]), .A2(n39), .ZN(n63) );
  NAND3_X1 U82 ( .A1(n63), .A2(n62), .A3(n61), .ZN(carry[14]) );
  NAND2_X1 U83 ( .A1(A[14]), .A2(B[14]), .ZN(n64) );
  NAND2_X1 U84 ( .A1(A[14]), .A2(carry[14]), .ZN(n65) );
  NAND2_X1 U85 ( .A1(B[14]), .A2(n58), .ZN(n66) );
  NAND3_X1 U86 ( .A1(n66), .A2(n65), .A3(n64), .ZN(carry[15]) );
  XNOR2_X1 U87 ( .A(carry[15]), .B(n67), .ZN(SUM[15]) );
  XNOR2_X1 U88 ( .A(B[15]), .B(A[15]), .ZN(n67) );
  XOR2_X1 U89 ( .A(A[8]), .B(B[8]), .Z(n68) );
  XOR2_X1 U90 ( .A(n68), .B(n32), .Z(SUM[8]) );
  NAND2_X1 U91 ( .A1(B[8]), .A2(A[8]), .ZN(n69) );
  NAND2_X1 U92 ( .A1(A[8]), .A2(carry[8]), .ZN(n70) );
  NAND2_X1 U93 ( .A1(n32), .A2(B[8]), .ZN(n71) );
  NAND3_X1 U94 ( .A1(n71), .A2(n70), .A3(n69), .ZN(carry[9]) );
  XOR2_X1 U95 ( .A(A[9]), .B(B[9]), .Z(n72) );
  XOR2_X1 U96 ( .A(n72), .B(n57), .Z(SUM[9]) );
  NAND2_X1 U97 ( .A1(A[9]), .A2(B[9]), .ZN(n73) );
  NAND2_X1 U98 ( .A1(A[9]), .A2(carry[9]), .ZN(n74) );
  NAND2_X1 U99 ( .A1(B[9]), .A2(n56), .ZN(n75) );
  NAND3_X1 U100 ( .A1(n75), .A2(n74), .A3(n73), .ZN(carry[10]) );
  XOR2_X1 U101 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U102 ( .A1(B[0]), .A2(A[0]), .ZN(n77) );
endmodule


module datapath_DW_mult_tc_28 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n286), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n285), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n289), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n288), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n291), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  INV_X1 U157 ( .A(n15), .ZN(n282) );
  AND2_X1 U158 ( .A1(n95), .A2(n102), .ZN(n206) );
  XNOR2_X1 U159 ( .A(n283), .B(n15), .ZN(n207) );
  AND3_X1 U160 ( .A1(n226), .A2(n227), .A3(n228), .ZN(product[15]) );
  XOR2_X1 U161 ( .A(n95), .B(n102), .Z(n209) );
  XOR2_X1 U162 ( .A(n103), .B(n96), .Z(n210) );
  XOR2_X1 U163 ( .A(n14), .B(n210), .Z(product[2]) );
  NAND2_X1 U164 ( .A1(n14), .A2(n103), .ZN(n211) );
  NAND2_X1 U165 ( .A1(n14), .A2(n96), .ZN(n212) );
  NAND2_X1 U166 ( .A1(n103), .A2(n96), .ZN(n213) );
  NAND3_X1 U167 ( .A1(n211), .A2(n212), .A3(n213), .ZN(n13) );
  NAND3_X1 U168 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n214) );
  NAND3_X1 U169 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n215) );
  NAND3_X1 U170 ( .A1(n223), .A2(n224), .A3(n225), .ZN(n216) );
  NAND3_X1 U171 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n217) );
  XNOR2_X1 U172 ( .A(n2), .B(n207), .ZN(product[14]) );
  XOR2_X1 U173 ( .A(n56), .B(n71), .Z(n218) );
  XOR2_X1 U174 ( .A(n218), .B(n13), .Z(product[3]) );
  NAND2_X1 U175 ( .A1(n13), .A2(n209), .ZN(n219) );
  NAND2_X1 U176 ( .A1(n13), .A2(n71), .ZN(n220) );
  NAND2_X1 U177 ( .A1(n209), .A2(n71), .ZN(n221) );
  NAND3_X1 U178 ( .A1(n219), .A2(n220), .A3(n221), .ZN(n12) );
  XOR2_X1 U179 ( .A(n27), .B(n24), .Z(n222) );
  XOR2_X1 U180 ( .A(n215), .B(n222), .Z(product[10]) );
  NAND2_X1 U181 ( .A1(n214), .A2(n27), .ZN(n223) );
  NAND2_X1 U182 ( .A1(n6), .A2(n24), .ZN(n224) );
  NAND2_X1 U183 ( .A1(n27), .A2(n24), .ZN(n225) );
  NAND3_X1 U184 ( .A1(n223), .A2(n224), .A3(n225), .ZN(n5) );
  NAND2_X1 U185 ( .A1(n217), .A2(n283), .ZN(n226) );
  NAND2_X1 U186 ( .A1(n217), .A2(n15), .ZN(n227) );
  NAND2_X1 U187 ( .A1(n283), .A2(n15), .ZN(n228) );
  NAND3_X1 U188 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n229) );
  NAND3_X1 U189 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n230) );
  NAND3_X1 U190 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n231) );
  XOR2_X1 U191 ( .A(n23), .B(n20), .Z(n232) );
  XOR2_X1 U192 ( .A(n216), .B(n232), .Z(product[11]) );
  NAND2_X1 U193 ( .A1(n216), .A2(n23), .ZN(n233) );
  NAND2_X1 U194 ( .A1(n5), .A2(n20), .ZN(n234) );
  NAND2_X1 U195 ( .A1(n23), .A2(n20), .ZN(n235) );
  NAND3_X1 U196 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n4) );
  XOR2_X1 U197 ( .A(n34), .B(n39), .Z(n236) );
  XOR2_X1 U198 ( .A(n230), .B(n236), .Z(product[8]) );
  NAND2_X1 U199 ( .A1(n229), .A2(n34), .ZN(n237) );
  NAND2_X1 U200 ( .A1(n8), .A2(n39), .ZN(n238) );
  NAND2_X1 U201 ( .A1(n34), .A2(n39), .ZN(n239) );
  NAND3_X1 U202 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n7) );
  NAND3_X1 U203 ( .A1(n249), .A2(n250), .A3(n251), .ZN(n240) );
  NAND3_X1 U204 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n241) );
  XNOR2_X1 U205 ( .A(b[1]), .B(n279), .ZN(n242) );
  NAND3_X1 U206 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n243) );
  XOR2_X1 U207 ( .A(n33), .B(n28), .Z(n244) );
  XOR2_X1 U208 ( .A(n231), .B(n244), .Z(product[9]) );
  NAND2_X1 U209 ( .A1(n231), .A2(n33), .ZN(n245) );
  NAND2_X1 U210 ( .A1(n7), .A2(n28), .ZN(n246) );
  NAND2_X1 U211 ( .A1(n33), .A2(n28), .ZN(n247) );
  NAND3_X1 U212 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n6) );
  XOR2_X1 U213 ( .A(n18), .B(n19), .Z(n248) );
  XOR2_X1 U214 ( .A(n4), .B(n248), .Z(product[12]) );
  NAND2_X1 U215 ( .A1(n4), .A2(n18), .ZN(n249) );
  NAND2_X1 U216 ( .A1(n4), .A2(n19), .ZN(n250) );
  NAND2_X1 U217 ( .A1(n18), .A2(n19), .ZN(n251) );
  NAND3_X1 U218 ( .A1(n249), .A2(n250), .A3(n251), .ZN(n3) );
  XOR2_X1 U219 ( .A(n54), .B(n206), .Z(n252) );
  XOR2_X1 U220 ( .A(n12), .B(n252), .Z(product[4]) );
  NAND2_X1 U221 ( .A1(n12), .A2(n54), .ZN(n253) );
  NAND2_X1 U222 ( .A1(n12), .A2(n206), .ZN(n254) );
  NAND2_X1 U223 ( .A1(n54), .A2(n206), .ZN(n255) );
  NAND3_X1 U224 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n11) );
  XOR2_X1 U225 ( .A(n17), .B(n282), .Z(n256) );
  XOR2_X1 U226 ( .A(n3), .B(n256), .Z(product[13]) );
  NAND2_X1 U227 ( .A1(n240), .A2(n17), .ZN(n257) );
  NAND2_X1 U228 ( .A1(n240), .A2(n282), .ZN(n258) );
  NAND2_X1 U229 ( .A1(n17), .A2(n282), .ZN(n259) );
  NAND3_X1 U230 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n2) );
  CLKBUF_X1 U231 ( .A(b[1]), .Z(n260) );
  XOR2_X1 U232 ( .A(n50), .B(n53), .Z(n261) );
  XOR2_X1 U233 ( .A(n243), .B(n261), .Z(product[5]) );
  NAND2_X1 U234 ( .A1(n11), .A2(n50), .ZN(n262) );
  NAND2_X1 U235 ( .A1(n11), .A2(n53), .ZN(n263) );
  NAND2_X1 U236 ( .A1(n50), .A2(n53), .ZN(n264) );
  NAND3_X1 U237 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n10) );
  NAND3_X1 U238 ( .A1(n267), .A2(n268), .A3(n269), .ZN(n265) );
  XOR2_X1 U239 ( .A(n95), .B(n102), .Z(n56) );
  XOR2_X1 U240 ( .A(n46), .B(n49), .Z(n266) );
  XOR2_X1 U241 ( .A(n241), .B(n266), .Z(product[6]) );
  NAND2_X1 U242 ( .A1(n241), .A2(n46), .ZN(n267) );
  NAND2_X1 U243 ( .A1(n10), .A2(n49), .ZN(n268) );
  NAND2_X1 U244 ( .A1(n46), .A2(n49), .ZN(n269) );
  NAND3_X1 U245 ( .A1(n267), .A2(n268), .A3(n269), .ZN(n9) );
  XOR2_X1 U246 ( .A(n40), .B(n45), .Z(n270) );
  XOR2_X1 U247 ( .A(n9), .B(n270), .Z(product[7]) );
  NAND2_X1 U248 ( .A1(n265), .A2(n40), .ZN(n271) );
  NAND2_X1 U249 ( .A1(n265), .A2(n45), .ZN(n272) );
  NAND2_X1 U250 ( .A1(n40), .A2(n45), .ZN(n273) );
  NAND3_X1 U251 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n8) );
  INV_X2 U252 ( .A(n281), .ZN(n280) );
  NAND2_X1 U253 ( .A1(a[4]), .A2(a[3]), .ZN(n275) );
  NAND2_X1 U254 ( .A1(n274), .A2(n290), .ZN(n276) );
  NAND2_X2 U255 ( .A1(n275), .A2(n276), .ZN(n308) );
  INV_X1 U256 ( .A(a[4]), .ZN(n274) );
  NAND2_X2 U257 ( .A1(n308), .A2(n337), .ZN(n310) );
  BUF_X1 U258 ( .A(n298), .Z(n277) );
  XOR2_X1 U259 ( .A(a[2]), .B(n278), .Z(n298) );
  INV_X1 U260 ( .A(n21), .ZN(n285) );
  INV_X1 U261 ( .A(n317), .ZN(n286) );
  INV_X1 U262 ( .A(n328), .ZN(n283) );
  INV_X1 U263 ( .A(b[0]), .ZN(n281) );
  INV_X1 U264 ( .A(n297), .ZN(n291) );
  INV_X1 U265 ( .A(n306), .ZN(n289) );
  INV_X1 U266 ( .A(n31), .ZN(n288) );
  XOR2_X1 U267 ( .A(a[6]), .B(n287), .Z(n319) );
  NAND2_X1 U268 ( .A1(n298), .A2(n336), .ZN(n300) );
  INV_X1 U269 ( .A(n278), .ZN(n279) );
  INV_X1 U270 ( .A(a[0]), .ZN(n292) );
  INV_X1 U271 ( .A(a[5]), .ZN(n287) );
  INV_X1 U272 ( .A(a[7]), .ZN(n284) );
  INV_X1 U273 ( .A(a[3]), .ZN(n290) );
  INV_X1 U274 ( .A(a[1]), .ZN(n278) );
  NOR2_X1 U275 ( .A1(n292), .A2(n281), .ZN(product[0]) );
  OAI22_X1 U276 ( .A1(n293), .A2(n294), .B1(n295), .B2(n292), .ZN(n99) );
  OAI22_X1 U277 ( .A1(n295), .A2(n294), .B1(n296), .B2(n292), .ZN(n98) );
  XNOR2_X1 U278 ( .A(b[6]), .B(n279), .ZN(n295) );
  OAI22_X1 U279 ( .A1(n292), .A2(n296), .B1(n294), .B2(n296), .ZN(n297) );
  XNOR2_X1 U280 ( .A(b[7]), .B(n279), .ZN(n296) );
  NOR2_X1 U281 ( .A1(n298), .A2(n281), .ZN(n96) );
  OAI22_X1 U282 ( .A1(n299), .A2(n300), .B1(n298), .B2(n301), .ZN(n95) );
  XNOR2_X1 U283 ( .A(a[3]), .B(n280), .ZN(n299) );
  OAI22_X1 U284 ( .A1(n301), .A2(n300), .B1(n277), .B2(n302), .ZN(n94) );
  XNOR2_X1 U285 ( .A(b[1]), .B(a[3]), .ZN(n301) );
  OAI22_X1 U286 ( .A1(n302), .A2(n300), .B1(n277), .B2(n303), .ZN(n93) );
  XNOR2_X1 U287 ( .A(b[2]), .B(a[3]), .ZN(n302) );
  OAI22_X1 U288 ( .A1(n303), .A2(n300), .B1(n277), .B2(n304), .ZN(n92) );
  XNOR2_X1 U289 ( .A(b[3]), .B(a[3]), .ZN(n303) );
  OAI22_X1 U290 ( .A1(n304), .A2(n300), .B1(n277), .B2(n305), .ZN(n91) );
  XNOR2_X1 U291 ( .A(b[4]), .B(a[3]), .ZN(n304) );
  OAI22_X1 U292 ( .A1(n307), .A2(n277), .B1(n300), .B2(n307), .ZN(n306) );
  NOR2_X1 U293 ( .A1(n308), .A2(n281), .ZN(n88) );
  OAI22_X1 U294 ( .A1(n309), .A2(n310), .B1(n308), .B2(n311), .ZN(n87) );
  XNOR2_X1 U295 ( .A(a[5]), .B(n280), .ZN(n309) );
  OAI22_X1 U296 ( .A1(n311), .A2(n310), .B1(n308), .B2(n312), .ZN(n86) );
  XNOR2_X1 U297 ( .A(n260), .B(a[5]), .ZN(n311) );
  OAI22_X1 U298 ( .A1(n312), .A2(n310), .B1(n308), .B2(n313), .ZN(n85) );
  XNOR2_X1 U299 ( .A(b[2]), .B(a[5]), .ZN(n312) );
  OAI22_X1 U300 ( .A1(n313), .A2(n310), .B1(n308), .B2(n314), .ZN(n84) );
  XNOR2_X1 U301 ( .A(b[3]), .B(a[5]), .ZN(n313) );
  OAI22_X1 U302 ( .A1(n314), .A2(n310), .B1(n308), .B2(n315), .ZN(n83) );
  XNOR2_X1 U303 ( .A(b[4]), .B(a[5]), .ZN(n314) );
  OAI22_X1 U304 ( .A1(n315), .A2(n310), .B1(n308), .B2(n316), .ZN(n82) );
  XNOR2_X1 U305 ( .A(b[5]), .B(a[5]), .ZN(n315) );
  OAI22_X1 U306 ( .A1(n318), .A2(n308), .B1(n310), .B2(n318), .ZN(n317) );
  NOR2_X1 U307 ( .A1(n319), .A2(n281), .ZN(n80) );
  OAI22_X1 U308 ( .A1(n320), .A2(n321), .B1(n319), .B2(n322), .ZN(n79) );
  XNOR2_X1 U309 ( .A(a[7]), .B(n280), .ZN(n320) );
  OAI22_X1 U310 ( .A1(n323), .A2(n321), .B1(n319), .B2(n324), .ZN(n77) );
  OAI22_X1 U311 ( .A1(n324), .A2(n321), .B1(n319), .B2(n325), .ZN(n76) );
  XNOR2_X1 U312 ( .A(b[3]), .B(a[7]), .ZN(n324) );
  OAI22_X1 U313 ( .A1(n325), .A2(n321), .B1(n319), .B2(n326), .ZN(n75) );
  XNOR2_X1 U314 ( .A(b[4]), .B(a[7]), .ZN(n325) );
  OAI22_X1 U315 ( .A1(n326), .A2(n321), .B1(n319), .B2(n327), .ZN(n74) );
  XNOR2_X1 U316 ( .A(b[5]), .B(a[7]), .ZN(n326) );
  OAI22_X1 U317 ( .A1(n329), .A2(n319), .B1(n321), .B2(n329), .ZN(n328) );
  OAI21_X1 U318 ( .B1(n280), .B2(n278), .A(n294), .ZN(n72) );
  OAI21_X1 U319 ( .B1(n290), .B2(n300), .A(n330), .ZN(n71) );
  OR3_X1 U320 ( .A1(n277), .A2(n280), .A3(n290), .ZN(n330) );
  OAI21_X1 U321 ( .B1(n287), .B2(n310), .A(n331), .ZN(n70) );
  OR3_X1 U322 ( .A1(n308), .A2(n280), .A3(n287), .ZN(n331) );
  OAI21_X1 U323 ( .B1(n284), .B2(n321), .A(n332), .ZN(n69) );
  OR3_X1 U324 ( .A1(n319), .A2(n280), .A3(n284), .ZN(n332) );
  XNOR2_X1 U325 ( .A(n333), .B(n334), .ZN(n38) );
  OR2_X1 U326 ( .A1(n333), .A2(n334), .ZN(n37) );
  OAI22_X1 U327 ( .A1(n305), .A2(n300), .B1(n277), .B2(n335), .ZN(n334) );
  XNOR2_X1 U328 ( .A(b[5]), .B(a[3]), .ZN(n305) );
  OAI22_X1 U329 ( .A1(n322), .A2(n321), .B1(n319), .B2(n323), .ZN(n333) );
  XNOR2_X1 U330 ( .A(b[2]), .B(a[7]), .ZN(n323) );
  XNOR2_X1 U331 ( .A(n260), .B(a[7]), .ZN(n322) );
  OAI22_X1 U332 ( .A1(n335), .A2(n300), .B1(n277), .B2(n307), .ZN(n31) );
  XNOR2_X1 U333 ( .A(b[7]), .B(a[3]), .ZN(n307) );
  XNOR2_X1 U334 ( .A(n290), .B(a[2]), .ZN(n336) );
  XNOR2_X1 U335 ( .A(b[6]), .B(a[3]), .ZN(n335) );
  OAI22_X1 U336 ( .A1(n316), .A2(n310), .B1(n308), .B2(n318), .ZN(n21) );
  XNOR2_X1 U337 ( .A(b[7]), .B(a[5]), .ZN(n318) );
  XNOR2_X1 U338 ( .A(n287), .B(a[4]), .ZN(n337) );
  XNOR2_X1 U339 ( .A(b[6]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U340 ( .A1(n327), .A2(n321), .B1(n319), .B2(n329), .ZN(n15) );
  XNOR2_X1 U341 ( .A(b[7]), .B(a[7]), .ZN(n329) );
  NAND2_X1 U342 ( .A1(n338), .A2(n319), .ZN(n321) );
  XNOR2_X1 U343 ( .A(n284), .B(a[6]), .ZN(n338) );
  XNOR2_X1 U344 ( .A(b[6]), .B(a[7]), .ZN(n327) );
  OAI22_X1 U345 ( .A1(n280), .A2(n294), .B1(n339), .B2(n292), .ZN(n104) );
  OAI22_X1 U346 ( .A1(n242), .A2(n294), .B1(n340), .B2(n292), .ZN(n103) );
  XNOR2_X1 U347 ( .A(b[1]), .B(n279), .ZN(n339) );
  OAI22_X1 U348 ( .A1(n340), .A2(n294), .B1(n341), .B2(n292), .ZN(n102) );
  XNOR2_X1 U349 ( .A(b[2]), .B(n279), .ZN(n340) );
  OAI22_X1 U350 ( .A1(n341), .A2(n294), .B1(n342), .B2(n292), .ZN(n101) );
  XNOR2_X1 U351 ( .A(b[3]), .B(n279), .ZN(n341) );
  OAI22_X1 U352 ( .A1(n342), .A2(n294), .B1(n293), .B2(n292), .ZN(n100) );
  XNOR2_X1 U353 ( .A(b[5]), .B(n279), .ZN(n293) );
  NAND2_X1 U354 ( .A1(a[1]), .A2(n292), .ZN(n294) );
  XNOR2_X1 U355 ( .A(b[4]), .B(n279), .ZN(n342) );
endmodule


module datapath_DW01_add_28 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n77;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n77), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(n64), .Z(n1) );
  CLKBUF_X1 U2 ( .A(n10), .Z(n2) );
  CLKBUF_X1 U3 ( .A(n51), .Z(n3) );
  CLKBUF_X1 U4 ( .A(n71), .Z(n4) );
  CLKBUF_X1 U5 ( .A(n24), .Z(n5) );
  NAND3_X1 U6 ( .A1(n32), .A2(n33), .A3(n34), .ZN(n6) );
  CLKBUF_X1 U7 ( .A(n35), .Z(n7) );
  NAND3_X1 U8 ( .A1(n73), .A2(n74), .A3(n75), .ZN(n8) );
  NAND3_X1 U9 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n9) );
  NAND3_X1 U10 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n10) );
  NAND3_X1 U11 ( .A1(n24), .A2(n25), .A3(n26), .ZN(n11) );
  NAND3_X1 U12 ( .A1(n5), .A2(n25), .A3(n26), .ZN(n12) );
  XOR2_X1 U13 ( .A(B[11]), .B(A[11]), .Z(n13) );
  XOR2_X1 U14 ( .A(n12), .B(n13), .Z(SUM[11]) );
  NAND2_X1 U15 ( .A1(n11), .A2(B[11]), .ZN(n14) );
  NAND2_X1 U16 ( .A1(carry[11]), .A2(A[11]), .ZN(n15) );
  NAND2_X1 U17 ( .A1(B[11]), .A2(A[11]), .ZN(n16) );
  NAND3_X1 U18 ( .A1(n15), .A2(n14), .A3(n16), .ZN(carry[12]) );
  CLKBUF_X1 U19 ( .A(n9), .Z(n17) );
  NAND3_X1 U20 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n18) );
  NAND3_X1 U21 ( .A1(n3), .A2(n52), .A3(n53), .ZN(n19) );
  CLKBUF_X1 U22 ( .A(n6), .Z(n20) );
  NAND3_X1 U23 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n21) );
  NAND3_X1 U24 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n22) );
  XOR2_X1 U25 ( .A(B[10]), .B(A[10]), .Z(n23) );
  XOR2_X1 U26 ( .A(n17), .B(n23), .Z(SUM[10]) );
  NAND2_X1 U27 ( .A1(n9), .A2(B[10]), .ZN(n24) );
  NAND2_X1 U28 ( .A1(carry[10]), .A2(A[10]), .ZN(n25) );
  NAND2_X1 U29 ( .A1(B[10]), .A2(A[10]), .ZN(n26) );
  NAND3_X1 U30 ( .A1(n24), .A2(n25), .A3(n26), .ZN(carry[11]) );
  XOR2_X1 U31 ( .A(carry[2]), .B(A[2]), .Z(n27) );
  XOR2_X1 U32 ( .A(B[2]), .B(n27), .Z(SUM[2]) );
  NAND2_X1 U33 ( .A1(B[2]), .A2(carry[2]), .ZN(n28) );
  NAND2_X1 U34 ( .A1(B[2]), .A2(A[2]), .ZN(n29) );
  NAND2_X1 U35 ( .A1(carry[2]), .A2(A[2]), .ZN(n30) );
  NAND3_X1 U36 ( .A1(n28), .A2(n29), .A3(n30), .ZN(carry[3]) );
  XOR2_X1 U37 ( .A(B[8]), .B(A[8]), .Z(n31) );
  XOR2_X1 U38 ( .A(n19), .B(n31), .Z(SUM[8]) );
  NAND2_X1 U39 ( .A1(n18), .A2(B[8]), .ZN(n32) );
  NAND2_X1 U40 ( .A1(carry[8]), .A2(A[8]), .ZN(n33) );
  NAND2_X1 U41 ( .A1(B[8]), .A2(A[8]), .ZN(n34) );
  NAND3_X1 U42 ( .A1(n32), .A2(n33), .A3(n34), .ZN(carry[9]) );
  NAND3_X1 U43 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n35) );
  XOR2_X1 U44 ( .A(B[9]), .B(A[9]), .Z(n36) );
  XOR2_X1 U45 ( .A(n20), .B(n36), .Z(SUM[9]) );
  NAND2_X1 U46 ( .A1(n6), .A2(B[9]), .ZN(n37) );
  NAND2_X1 U47 ( .A1(carry[9]), .A2(A[9]), .ZN(n38) );
  NAND2_X1 U48 ( .A1(B[9]), .A2(A[9]), .ZN(n39) );
  NAND3_X1 U49 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[10]) );
  XOR2_X1 U50 ( .A(B[12]), .B(A[12]), .Z(n40) );
  XOR2_X1 U51 ( .A(n2), .B(n40), .Z(SUM[12]) );
  NAND2_X1 U52 ( .A1(n10), .A2(B[12]), .ZN(n41) );
  NAND2_X1 U53 ( .A1(carry[12]), .A2(A[12]), .ZN(n42) );
  NAND2_X1 U54 ( .A1(B[12]), .A2(A[12]), .ZN(n43) );
  NAND3_X1 U55 ( .A1(n41), .A2(n42), .A3(n43), .ZN(carry[13]) );
  CLKBUF_X1 U56 ( .A(n8), .Z(n44) );
  NAND3_X1 U57 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n45) );
  XOR2_X1 U58 ( .A(B[13]), .B(A[13]), .Z(n46) );
  XOR2_X1 U59 ( .A(n7), .B(n46), .Z(SUM[13]) );
  NAND2_X1 U60 ( .A1(n35), .A2(B[13]), .ZN(n47) );
  NAND2_X1 U61 ( .A1(carry[13]), .A2(A[13]), .ZN(n48) );
  NAND2_X1 U62 ( .A1(B[13]), .A2(A[13]), .ZN(n49) );
  NAND3_X1 U63 ( .A1(n47), .A2(n48), .A3(n49), .ZN(carry[14]) );
  XOR2_X1 U64 ( .A(B[7]), .B(A[7]), .Z(n50) );
  XOR2_X1 U65 ( .A(n44), .B(n50), .Z(SUM[7]) );
  NAND2_X1 U66 ( .A1(n8), .A2(B[7]), .ZN(n51) );
  NAND2_X1 U67 ( .A1(carry[7]), .A2(A[7]), .ZN(n52) );
  NAND2_X1 U68 ( .A1(B[7]), .A2(A[7]), .ZN(n53) );
  NAND3_X1 U69 ( .A1(n51), .A2(n52), .A3(n53), .ZN(carry[8]) );
  XOR2_X1 U70 ( .A(B[3]), .B(A[3]), .Z(n54) );
  XOR2_X1 U71 ( .A(n22), .B(n54), .Z(SUM[3]) );
  NAND2_X1 U72 ( .A1(n21), .A2(B[3]), .ZN(n55) );
  NAND2_X1 U73 ( .A1(carry[3]), .A2(A[3]), .ZN(n56) );
  NAND2_X1 U74 ( .A1(B[3]), .A2(A[3]), .ZN(n57) );
  NAND3_X1 U75 ( .A1(n55), .A2(n56), .A3(n57), .ZN(carry[4]) );
  XNOR2_X1 U76 ( .A(carry[15]), .B(n58), .ZN(SUM[15]) );
  XNOR2_X1 U77 ( .A(B[15]), .B(A[15]), .ZN(n58) );
  CLKBUF_X1 U78 ( .A(n70), .Z(n59) );
  NAND3_X1 U79 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n60) );
  NAND3_X1 U80 ( .A1(n63), .A2(n1), .A3(n65), .ZN(n61) );
  XOR2_X1 U81 ( .A(B[4]), .B(A[4]), .Z(n62) );
  XOR2_X1 U82 ( .A(carry[4]), .B(n62), .Z(SUM[4]) );
  NAND2_X1 U83 ( .A1(n45), .A2(B[4]), .ZN(n63) );
  NAND2_X1 U84 ( .A1(carry[4]), .A2(A[4]), .ZN(n64) );
  NAND2_X1 U85 ( .A1(B[4]), .A2(A[4]), .ZN(n65) );
  NAND3_X1 U86 ( .A1(n63), .A2(n64), .A3(n65), .ZN(carry[5]) );
  NAND3_X1 U87 ( .A1(n69), .A2(n70), .A3(n71), .ZN(n66) );
  NAND3_X1 U88 ( .A1(n69), .A2(n59), .A3(n4), .ZN(n67) );
  XOR2_X1 U89 ( .A(A[5]), .B(B[5]), .Z(n68) );
  XOR2_X1 U90 ( .A(n68), .B(n61), .Z(SUM[5]) );
  NAND2_X1 U91 ( .A1(B[5]), .A2(A[5]), .ZN(n69) );
  NAND2_X1 U92 ( .A1(A[5]), .A2(n60), .ZN(n70) );
  NAND2_X1 U93 ( .A1(B[5]), .A2(carry[5]), .ZN(n71) );
  NAND3_X1 U94 ( .A1(n69), .A2(n70), .A3(n71), .ZN(carry[6]) );
  XOR2_X1 U95 ( .A(A[6]), .B(B[6]), .Z(n72) );
  XOR2_X1 U96 ( .A(n72), .B(n67), .Z(SUM[6]) );
  NAND2_X1 U97 ( .A1(A[6]), .A2(B[6]), .ZN(n73) );
  NAND2_X1 U98 ( .A1(A[6]), .A2(n66), .ZN(n74) );
  NAND2_X1 U99 ( .A1(B[6]), .A2(carry[6]), .ZN(n75) );
  NAND3_X1 U100 ( .A1(n73), .A2(n74), .A3(n75), .ZN(carry[7]) );
  XOR2_X1 U101 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U102 ( .A1(B[0]), .A2(A[0]), .ZN(n77) );
endmodule


module datapath_DW_mult_tc_27 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74,
         n75, n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92,
         n93, n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346;

  FA_X1 U12 ( .A(n54), .B(n55), .CI(n12), .CO(n11), .S(product[4]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n289), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n288), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n292), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n291), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n294), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n88), .B(n101), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  AND3_X1 U157 ( .A1(n210), .A2(n211), .A3(n212), .ZN(product[15]) );
  XOR2_X2 U158 ( .A(a[6]), .B(n290), .Z(n323) );
  XNOR2_X1 U159 ( .A(n11), .B(n207), .ZN(product[5]) );
  XNOR2_X1 U160 ( .A(n50), .B(n53), .ZN(n207) );
  XNOR2_X1 U161 ( .A(n208), .B(n236), .ZN(product[3]) );
  XNOR2_X1 U162 ( .A(n56), .B(n71), .ZN(n208) );
  XOR2_X1 U163 ( .A(n286), .B(n15), .Z(n209) );
  XOR2_X1 U164 ( .A(n2), .B(n209), .Z(product[14]) );
  NAND2_X1 U165 ( .A1(n2), .A2(n286), .ZN(n210) );
  NAND2_X1 U166 ( .A1(n2), .A2(n15), .ZN(n211) );
  NAND2_X1 U167 ( .A1(n286), .A2(n15), .ZN(n212) );
  NAND3_X1 U168 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n213) );
  NAND3_X1 U169 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n214) );
  NAND3_X1 U170 ( .A1(n221), .A2(n222), .A3(n223), .ZN(n215) );
  NAND3_X1 U171 ( .A1(n270), .A2(n271), .A3(n272), .ZN(n216) );
  NAND3_X1 U172 ( .A1(n270), .A2(n271), .A3(n272), .ZN(n217) );
  NAND3_X1 U173 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n218) );
  NAND3_X1 U174 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n219) );
  XOR2_X1 U175 ( .A(n33), .B(n28), .Z(n220) );
  XOR2_X1 U176 ( .A(n214), .B(n220), .Z(product[9]) );
  NAND2_X1 U177 ( .A1(n213), .A2(n33), .ZN(n221) );
  NAND2_X1 U178 ( .A1(n7), .A2(n28), .ZN(n222) );
  NAND2_X1 U179 ( .A1(n33), .A2(n28), .ZN(n223) );
  NAND3_X1 U180 ( .A1(n221), .A2(n222), .A3(n223), .ZN(n6) );
  XOR2_X1 U181 ( .A(n95), .B(n102), .Z(n224) );
  NAND3_X1 U182 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n225) );
  NAND3_X1 U183 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n226) );
  CLKBUF_X1 U184 ( .A(b[3]), .Z(n227) );
  XOR2_X1 U185 ( .A(n17), .B(n285), .Z(n228) );
  XOR2_X1 U186 ( .A(n217), .B(n228), .Z(product[13]) );
  NAND2_X1 U187 ( .A1(n216), .A2(n17), .ZN(n229) );
  NAND2_X1 U188 ( .A1(n3), .A2(n285), .ZN(n230) );
  NAND2_X1 U189 ( .A1(n17), .A2(n285), .ZN(n231) );
  NAND3_X1 U190 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n2) );
  NAND2_X1 U191 ( .A1(n11), .A2(n50), .ZN(n232) );
  NAND2_X1 U192 ( .A1(n11), .A2(n53), .ZN(n233) );
  NAND2_X1 U193 ( .A1(n50), .A2(n53), .ZN(n234) );
  NAND3_X1 U194 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n10) );
  NAND3_X1 U195 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n235) );
  NAND3_X1 U196 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n236) );
  NAND3_X1 U197 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n237) );
  XOR2_X1 U198 ( .A(n46), .B(n49), .Z(n238) );
  XOR2_X1 U199 ( .A(n226), .B(n238), .Z(product[6]) );
  NAND2_X1 U200 ( .A1(n225), .A2(n46), .ZN(n239) );
  NAND2_X1 U201 ( .A1(n10), .A2(n49), .ZN(n240) );
  NAND2_X1 U202 ( .A1(n46), .A2(n49), .ZN(n241) );
  NAND3_X1 U203 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n9) );
  XOR2_X1 U204 ( .A(n27), .B(n24), .Z(n242) );
  XOR2_X1 U205 ( .A(n215), .B(n242), .Z(product[10]) );
  NAND2_X1 U206 ( .A1(n215), .A2(n27), .ZN(n243) );
  NAND2_X1 U207 ( .A1(n6), .A2(n24), .ZN(n244) );
  NAND2_X1 U208 ( .A1(n27), .A2(n24), .ZN(n245) );
  NAND3_X1 U209 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n5) );
  NAND3_X1 U210 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n246) );
  NAND3_X1 U211 ( .A1(n252), .A2(n251), .A3(n250), .ZN(n247) );
  NAND3_X1 U212 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n248) );
  XOR2_X1 U213 ( .A(n40), .B(n45), .Z(n249) );
  XOR2_X1 U214 ( .A(n249), .B(n237), .Z(product[7]) );
  NAND2_X1 U215 ( .A1(n40), .A2(n45), .ZN(n250) );
  NAND2_X1 U216 ( .A1(n40), .A2(n9), .ZN(n251) );
  NAND2_X1 U217 ( .A1(n45), .A2(n9), .ZN(n252) );
  NAND3_X1 U218 ( .A1(n251), .A2(n250), .A3(n252), .ZN(n8) );
  XOR2_X1 U219 ( .A(n34), .B(n39), .Z(n253) );
  XOR2_X1 U220 ( .A(n253), .B(n248), .Z(product[8]) );
  NAND2_X1 U221 ( .A1(n34), .A2(n39), .ZN(n254) );
  NAND2_X1 U222 ( .A1(n34), .A2(n247), .ZN(n255) );
  NAND2_X1 U223 ( .A1(n39), .A2(n8), .ZN(n256) );
  NAND3_X1 U224 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n7) );
  XOR2_X1 U225 ( .A(n103), .B(n96), .Z(n257) );
  XOR2_X1 U226 ( .A(n257), .B(n14), .Z(product[2]) );
  NAND2_X1 U227 ( .A1(n103), .A2(n96), .ZN(n258) );
  NAND2_X1 U228 ( .A1(n103), .A2(n14), .ZN(n259) );
  NAND2_X1 U229 ( .A1(n96), .A2(n14), .ZN(n260) );
  NAND3_X1 U230 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n13) );
  NAND2_X1 U231 ( .A1(n224), .A2(n71), .ZN(n261) );
  NAND2_X1 U232 ( .A1(n224), .A2(n235), .ZN(n262) );
  NAND2_X1 U233 ( .A1(n71), .A2(n13), .ZN(n263) );
  NAND3_X1 U234 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n12) );
  INV_X1 U235 ( .A(b[0]), .ZN(n264) );
  NAND2_X2 U236 ( .A1(n302), .A2(n340), .ZN(n304) );
  XOR2_X1 U237 ( .A(n20), .B(n23), .Z(n265) );
  XOR2_X1 U238 ( .A(n265), .B(n219), .Z(product[11]) );
  NAND2_X1 U239 ( .A1(n20), .A2(n23), .ZN(n266) );
  NAND2_X1 U240 ( .A1(n20), .A2(n5), .ZN(n267) );
  NAND2_X1 U241 ( .A1(n23), .A2(n218), .ZN(n268) );
  NAND3_X1 U242 ( .A1(n268), .A2(n267), .A3(n266), .ZN(n4) );
  XOR2_X1 U243 ( .A(n19), .B(n18), .Z(n269) );
  XOR2_X1 U244 ( .A(n269), .B(n246), .Z(product[12]) );
  NAND2_X1 U245 ( .A1(n19), .A2(n18), .ZN(n270) );
  NAND2_X1 U246 ( .A1(n19), .A2(n4), .ZN(n271) );
  NAND2_X1 U247 ( .A1(n4), .A2(n18), .ZN(n272) );
  NAND3_X1 U248 ( .A1(n270), .A2(n271), .A3(n272), .ZN(n3) );
  INV_X2 U249 ( .A(n284), .ZN(n283) );
  NAND2_X1 U250 ( .A1(a[4]), .A2(a[3]), .ZN(n275) );
  NAND2_X1 U251 ( .A1(n273), .A2(n274), .ZN(n276) );
  NAND2_X2 U252 ( .A1(n275), .A2(n276), .ZN(n312) );
  INV_X1 U253 ( .A(a[4]), .ZN(n273) );
  INV_X1 U254 ( .A(a[3]), .ZN(n274) );
  NAND2_X2 U255 ( .A1(n312), .A2(n341), .ZN(n314) );
  INV_X1 U256 ( .A(n302), .ZN(n277) );
  INV_X1 U257 ( .A(n277), .ZN(n278) );
  NAND2_X1 U258 ( .A1(n281), .A2(n282), .ZN(n302) );
  NAND2_X1 U259 ( .A1(a[2]), .A2(a[1]), .ZN(n281) );
  NAND2_X1 U260 ( .A1(n279), .A2(n280), .ZN(n282) );
  INV_X1 U261 ( .A(a[2]), .ZN(n279) );
  INV_X1 U262 ( .A(a[1]), .ZN(n280) );
  INV_X1 U263 ( .A(a[0]), .ZN(n296) );
  INV_X1 U264 ( .A(n15), .ZN(n285) );
  INV_X1 U265 ( .A(n21), .ZN(n288) );
  INV_X1 U266 ( .A(n321), .ZN(n289) );
  INV_X1 U267 ( .A(n332), .ZN(n286) );
  INV_X1 U268 ( .A(b[0]), .ZN(n284) );
  INV_X1 U269 ( .A(n301), .ZN(n294) );
  INV_X1 U270 ( .A(n310), .ZN(n292) );
  INV_X1 U271 ( .A(n31), .ZN(n291) );
  INV_X1 U272 ( .A(a[5]), .ZN(n290) );
  INV_X1 U273 ( .A(a[7]), .ZN(n287) );
  INV_X1 U274 ( .A(a[3]), .ZN(n293) );
  INV_X1 U275 ( .A(a[1]), .ZN(n295) );
  NOR2_X1 U276 ( .A1(n296), .A2(n264), .ZN(product[0]) );
  OAI22_X1 U277 ( .A1(n297), .A2(n298), .B1(n299), .B2(n296), .ZN(n99) );
  OAI22_X1 U278 ( .A1(n299), .A2(n298), .B1(n300), .B2(n296), .ZN(n98) );
  XNOR2_X1 U279 ( .A(b[6]), .B(a[1]), .ZN(n299) );
  OAI22_X1 U280 ( .A1(n296), .A2(n300), .B1(n298), .B2(n300), .ZN(n301) );
  XNOR2_X1 U281 ( .A(b[7]), .B(a[1]), .ZN(n300) );
  NOR2_X1 U282 ( .A1(n302), .A2(n264), .ZN(n96) );
  OAI22_X1 U283 ( .A1(n303), .A2(n304), .B1(n302), .B2(n305), .ZN(n95) );
  XNOR2_X1 U284 ( .A(a[3]), .B(n283), .ZN(n303) );
  OAI22_X1 U285 ( .A1(n305), .A2(n304), .B1(n278), .B2(n306), .ZN(n94) );
  XNOR2_X1 U286 ( .A(b[1]), .B(a[3]), .ZN(n305) );
  OAI22_X1 U287 ( .A1(n306), .A2(n304), .B1(n278), .B2(n307), .ZN(n93) );
  XNOR2_X1 U288 ( .A(b[2]), .B(a[3]), .ZN(n306) );
  OAI22_X1 U289 ( .A1(n307), .A2(n304), .B1(n278), .B2(n308), .ZN(n92) );
  XNOR2_X1 U290 ( .A(b[3]), .B(a[3]), .ZN(n307) );
  OAI22_X1 U291 ( .A1(n308), .A2(n304), .B1(n278), .B2(n309), .ZN(n91) );
  XNOR2_X1 U292 ( .A(b[4]), .B(a[3]), .ZN(n308) );
  OAI22_X1 U293 ( .A1(n311), .A2(n278), .B1(n304), .B2(n311), .ZN(n310) );
  NOR2_X1 U294 ( .A1(n312), .A2(n264), .ZN(n88) );
  OAI22_X1 U295 ( .A1(n313), .A2(n314), .B1(n312), .B2(n315), .ZN(n87) );
  XNOR2_X1 U296 ( .A(a[5]), .B(n283), .ZN(n313) );
  OAI22_X1 U297 ( .A1(n315), .A2(n314), .B1(n312), .B2(n316), .ZN(n86) );
  XNOR2_X1 U298 ( .A(b[1]), .B(a[5]), .ZN(n315) );
  OAI22_X1 U299 ( .A1(n316), .A2(n314), .B1(n312), .B2(n317), .ZN(n85) );
  XNOR2_X1 U300 ( .A(b[2]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U301 ( .A1(n317), .A2(n314), .B1(n312), .B2(n318), .ZN(n84) );
  XNOR2_X1 U302 ( .A(n227), .B(a[5]), .ZN(n317) );
  OAI22_X1 U303 ( .A1(n318), .A2(n314), .B1(n312), .B2(n319), .ZN(n83) );
  XNOR2_X1 U304 ( .A(b[4]), .B(a[5]), .ZN(n318) );
  OAI22_X1 U305 ( .A1(n319), .A2(n314), .B1(n312), .B2(n320), .ZN(n82) );
  XNOR2_X1 U306 ( .A(b[5]), .B(a[5]), .ZN(n319) );
  OAI22_X1 U307 ( .A1(n322), .A2(n312), .B1(n314), .B2(n322), .ZN(n321) );
  NOR2_X1 U308 ( .A1(n323), .A2(n264), .ZN(n80) );
  OAI22_X1 U309 ( .A1(n324), .A2(n325), .B1(n323), .B2(n326), .ZN(n79) );
  XNOR2_X1 U310 ( .A(a[7]), .B(n283), .ZN(n324) );
  OAI22_X1 U311 ( .A1(n327), .A2(n325), .B1(n323), .B2(n328), .ZN(n77) );
  OAI22_X1 U312 ( .A1(n328), .A2(n325), .B1(n323), .B2(n329), .ZN(n76) );
  XNOR2_X1 U313 ( .A(n227), .B(a[7]), .ZN(n328) );
  OAI22_X1 U314 ( .A1(n329), .A2(n325), .B1(n323), .B2(n330), .ZN(n75) );
  XNOR2_X1 U315 ( .A(b[4]), .B(a[7]), .ZN(n329) );
  OAI22_X1 U316 ( .A1(n330), .A2(n325), .B1(n323), .B2(n331), .ZN(n74) );
  XNOR2_X1 U317 ( .A(b[5]), .B(a[7]), .ZN(n330) );
  OAI22_X1 U318 ( .A1(n333), .A2(n323), .B1(n325), .B2(n333), .ZN(n332) );
  OAI21_X1 U319 ( .B1(n283), .B2(n295), .A(n298), .ZN(n72) );
  OAI21_X1 U320 ( .B1(n293), .B2(n304), .A(n334), .ZN(n71) );
  OR3_X1 U321 ( .A1(n302), .A2(n283), .A3(n293), .ZN(n334) );
  OAI21_X1 U322 ( .B1(n290), .B2(n314), .A(n335), .ZN(n70) );
  OR3_X1 U323 ( .A1(n312), .A2(n283), .A3(n290), .ZN(n335) );
  OAI21_X1 U324 ( .B1(n287), .B2(n325), .A(n336), .ZN(n69) );
  OR3_X1 U325 ( .A1(n323), .A2(n283), .A3(n287), .ZN(n336) );
  XNOR2_X1 U326 ( .A(n337), .B(n338), .ZN(n38) );
  OR2_X1 U327 ( .A1(n337), .A2(n338), .ZN(n37) );
  OAI22_X1 U328 ( .A1(n309), .A2(n304), .B1(n278), .B2(n339), .ZN(n338) );
  XNOR2_X1 U329 ( .A(b[5]), .B(a[3]), .ZN(n309) );
  OAI22_X1 U330 ( .A1(n326), .A2(n325), .B1(n323), .B2(n327), .ZN(n337) );
  XNOR2_X1 U331 ( .A(b[2]), .B(a[7]), .ZN(n327) );
  XNOR2_X1 U332 ( .A(b[1]), .B(a[7]), .ZN(n326) );
  OAI22_X1 U333 ( .A1(n339), .A2(n304), .B1(n278), .B2(n311), .ZN(n31) );
  XNOR2_X1 U334 ( .A(b[7]), .B(a[3]), .ZN(n311) );
  XNOR2_X1 U335 ( .A(n293), .B(a[2]), .ZN(n340) );
  XNOR2_X1 U336 ( .A(b[6]), .B(a[3]), .ZN(n339) );
  OAI22_X1 U337 ( .A1(n320), .A2(n314), .B1(n312), .B2(n322), .ZN(n21) );
  XNOR2_X1 U338 ( .A(b[7]), .B(a[5]), .ZN(n322) );
  XNOR2_X1 U339 ( .A(n290), .B(a[4]), .ZN(n341) );
  XNOR2_X1 U340 ( .A(b[6]), .B(a[5]), .ZN(n320) );
  OAI22_X1 U341 ( .A1(n331), .A2(n325), .B1(n323), .B2(n333), .ZN(n15) );
  XNOR2_X1 U342 ( .A(b[7]), .B(a[7]), .ZN(n333) );
  NAND2_X1 U343 ( .A1(n323), .A2(n342), .ZN(n325) );
  XNOR2_X1 U344 ( .A(n287), .B(a[6]), .ZN(n342) );
  XNOR2_X1 U345 ( .A(b[6]), .B(a[7]), .ZN(n331) );
  OAI22_X1 U346 ( .A1(n283), .A2(n298), .B1(n343), .B2(n296), .ZN(n104) );
  OAI22_X1 U347 ( .A1(n343), .A2(n298), .B1(n344), .B2(n296), .ZN(n103) );
  XNOR2_X1 U348 ( .A(b[1]), .B(a[1]), .ZN(n343) );
  OAI22_X1 U349 ( .A1(n344), .A2(n298), .B1(n345), .B2(n296), .ZN(n102) );
  XNOR2_X1 U350 ( .A(b[2]), .B(a[1]), .ZN(n344) );
  OAI22_X1 U351 ( .A1(n345), .A2(n298), .B1(n346), .B2(n296), .ZN(n101) );
  XNOR2_X1 U352 ( .A(b[3]), .B(a[1]), .ZN(n345) );
  OAI22_X1 U353 ( .A1(n346), .A2(n298), .B1(n297), .B2(n296), .ZN(n100) );
  XNOR2_X1 U354 ( .A(b[5]), .B(a[1]), .ZN(n297) );
  NAND2_X1 U355 ( .A1(a[1]), .A2(n296), .ZN(n298) );
  XNOR2_X1 U356 ( .A(b[4]), .B(a[1]), .ZN(n346) );
endmodule


module datapath_DW01_add_27 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n68;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n68), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND3_X1 U1 ( .A1(n23), .A2(n24), .A3(n25), .ZN(n1) );
  NAND3_X1 U2 ( .A1(n23), .A2(n24), .A3(n25), .ZN(n2) );
  CLKBUF_X1 U3 ( .A(carry[10]), .Z(n3) );
  CLKBUF_X1 U4 ( .A(n58), .Z(n4) );
  XOR2_X1 U5 ( .A(B[11]), .B(A[11]), .Z(n5) );
  XOR2_X1 U6 ( .A(n2), .B(n5), .Z(SUM[11]) );
  NAND2_X1 U7 ( .A1(n1), .A2(B[11]), .ZN(n6) );
  NAND2_X1 U8 ( .A1(carry[11]), .A2(A[11]), .ZN(n7) );
  NAND2_X1 U9 ( .A1(B[11]), .A2(A[11]), .ZN(n8) );
  NAND3_X1 U10 ( .A1(n6), .A2(n7), .A3(n8), .ZN(carry[12]) );
  XOR2_X1 U11 ( .A(B[9]), .B(A[9]), .Z(n9) );
  XOR2_X1 U12 ( .A(carry[9]), .B(n9), .Z(SUM[9]) );
  NAND2_X1 U13 ( .A1(carry[9]), .A2(B[9]), .ZN(n10) );
  NAND2_X1 U14 ( .A1(carry[9]), .A2(A[9]), .ZN(n11) );
  NAND2_X1 U15 ( .A1(B[9]), .A2(A[9]), .ZN(n12) );
  NAND3_X1 U16 ( .A1(n10), .A2(n11), .A3(n12), .ZN(carry[10]) );
  CLKBUF_X1 U17 ( .A(n16), .Z(n13) );
  NAND3_X1 U18 ( .A1(n35), .A2(n36), .A3(n37), .ZN(n14) );
  NAND3_X1 U19 ( .A1(n35), .A2(n36), .A3(n37), .ZN(n15) );
  NAND3_X1 U20 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n16) );
  NAND3_X1 U21 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n17) );
  NAND3_X1 U22 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n18) );
  NAND3_X1 U23 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n19) );
  NAND3_X1 U24 ( .A1(n60), .A2(n61), .A3(n62), .ZN(n20) );
  NAND3_X1 U25 ( .A1(n60), .A2(n61), .A3(n62), .ZN(n21) );
  XOR2_X1 U26 ( .A(B[10]), .B(A[10]), .Z(n22) );
  XOR2_X1 U27 ( .A(n3), .B(n22), .Z(SUM[10]) );
  NAND2_X1 U28 ( .A1(carry[10]), .A2(B[10]), .ZN(n23) );
  NAND2_X1 U29 ( .A1(carry[10]), .A2(A[10]), .ZN(n24) );
  NAND2_X1 U30 ( .A1(B[10]), .A2(A[10]), .ZN(n25) );
  NAND3_X1 U31 ( .A1(n23), .A2(n24), .A3(n25), .ZN(carry[11]) );
  NAND3_X1 U32 ( .A1(n58), .A2(n57), .A3(n56), .ZN(n26) );
  NAND3_X1 U33 ( .A1(n56), .A2(n57), .A3(n4), .ZN(n27) );
  NAND3_X1 U34 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n28) );
  NAND3_X1 U35 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n29) );
  XOR2_X1 U36 ( .A(B[8]), .B(A[8]), .Z(n30) );
  XOR2_X1 U37 ( .A(n27), .B(n30), .Z(SUM[8]) );
  NAND2_X1 U38 ( .A1(n26), .A2(B[8]), .ZN(n31) );
  NAND2_X1 U39 ( .A1(carry[8]), .A2(A[8]), .ZN(n32) );
  NAND2_X1 U40 ( .A1(B[8]), .A2(A[8]), .ZN(n33) );
  NAND3_X1 U41 ( .A1(n31), .A2(n32), .A3(n33), .ZN(carry[9]) );
  XOR2_X1 U42 ( .A(n29), .B(A[4]), .Z(n34) );
  XOR2_X1 U43 ( .A(B[4]), .B(n34), .Z(SUM[4]) );
  NAND2_X1 U44 ( .A1(B[4]), .A2(n28), .ZN(n35) );
  NAND2_X1 U45 ( .A1(B[4]), .A2(A[4]), .ZN(n36) );
  NAND2_X1 U46 ( .A1(carry[4]), .A2(A[4]), .ZN(n37) );
  NAND3_X1 U47 ( .A1(n35), .A2(n36), .A3(n37), .ZN(carry[5]) );
  XOR2_X1 U48 ( .A(B[12]), .B(A[12]), .Z(n38) );
  XOR2_X1 U49 ( .A(carry[12]), .B(n38), .Z(SUM[12]) );
  NAND2_X1 U50 ( .A1(carry[12]), .A2(B[12]), .ZN(n39) );
  NAND2_X1 U51 ( .A1(carry[12]), .A2(A[12]), .ZN(n40) );
  NAND2_X1 U52 ( .A1(B[12]), .A2(A[12]), .ZN(n41) );
  NAND3_X1 U53 ( .A1(n39), .A2(n40), .A3(n41), .ZN(carry[13]) );
  XOR2_X1 U54 ( .A(B[13]), .B(A[13]), .Z(n42) );
  XOR2_X1 U55 ( .A(n13), .B(n42), .Z(SUM[13]) );
  NAND2_X1 U56 ( .A1(n16), .A2(B[13]), .ZN(n43) );
  NAND2_X1 U57 ( .A1(carry[13]), .A2(A[13]), .ZN(n44) );
  NAND2_X1 U58 ( .A1(B[13]), .A2(A[13]), .ZN(n45) );
  NAND3_X1 U59 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[14]) );
  XNOR2_X1 U60 ( .A(carry[15]), .B(n46), .ZN(SUM[15]) );
  XNOR2_X1 U61 ( .A(B[15]), .B(A[15]), .ZN(n46) );
  XOR2_X1 U62 ( .A(B[5]), .B(A[5]), .Z(n47) );
  XOR2_X1 U63 ( .A(n15), .B(n47), .Z(SUM[5]) );
  NAND2_X1 U64 ( .A1(B[5]), .A2(n14), .ZN(n48) );
  NAND2_X1 U65 ( .A1(carry[5]), .A2(A[5]), .ZN(n49) );
  NAND2_X1 U66 ( .A1(B[5]), .A2(A[5]), .ZN(n50) );
  NAND3_X1 U67 ( .A1(n48), .A2(n49), .A3(n50), .ZN(carry[6]) );
  XOR2_X1 U68 ( .A(A[6]), .B(B[6]), .Z(n51) );
  XOR2_X1 U69 ( .A(n51), .B(n18), .Z(SUM[6]) );
  NAND2_X1 U70 ( .A1(A[6]), .A2(B[6]), .ZN(n52) );
  NAND2_X1 U71 ( .A1(A[6]), .A2(n17), .ZN(n53) );
  NAND2_X1 U72 ( .A1(B[6]), .A2(carry[6]), .ZN(n54) );
  NAND3_X1 U73 ( .A1(n52), .A2(n53), .A3(n54), .ZN(carry[7]) );
  XOR2_X1 U74 ( .A(A[7]), .B(B[7]), .Z(n55) );
  XOR2_X1 U75 ( .A(n55), .B(carry[7]), .Z(SUM[7]) );
  NAND2_X1 U76 ( .A1(A[7]), .A2(B[7]), .ZN(n56) );
  NAND2_X1 U77 ( .A1(A[7]), .A2(n19), .ZN(n57) );
  NAND2_X1 U78 ( .A1(B[7]), .A2(carry[7]), .ZN(n58) );
  NAND3_X1 U79 ( .A1(n56), .A2(n57), .A3(n58), .ZN(carry[8]) );
  XOR2_X1 U80 ( .A(A[2]), .B(B[2]), .Z(n59) );
  XOR2_X1 U81 ( .A(n59), .B(carry[2]), .Z(SUM[2]) );
  NAND2_X1 U82 ( .A1(A[2]), .A2(B[2]), .ZN(n60) );
  NAND2_X1 U83 ( .A1(A[2]), .A2(carry[2]), .ZN(n61) );
  NAND2_X1 U84 ( .A1(B[2]), .A2(carry[2]), .ZN(n62) );
  NAND3_X1 U85 ( .A1(n60), .A2(n61), .A3(n62), .ZN(carry[3]) );
  XOR2_X1 U86 ( .A(A[3]), .B(B[3]), .Z(n63) );
  XOR2_X1 U87 ( .A(n63), .B(n21), .Z(SUM[3]) );
  NAND2_X1 U88 ( .A1(A[3]), .A2(B[3]), .ZN(n64) );
  NAND2_X1 U89 ( .A1(A[3]), .A2(n20), .ZN(n65) );
  NAND2_X1 U90 ( .A1(B[3]), .A2(carry[3]), .ZN(n66) );
  NAND3_X1 U91 ( .A1(n64), .A2(n65), .A3(n66), .ZN(carry[4]) );
  XOR2_X1 U92 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U93 ( .A1(B[0]), .A2(A[0]), .ZN(n68) );
endmodule


module datapath_DW_mult_tc_26 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74,
         n75, n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92,
         n93, n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343;

  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n288), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n287), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n291), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n290), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n292), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  INV_X1 U157 ( .A(n15), .ZN(n284) );
  XNOR2_X1 U158 ( .A(n285), .B(n15), .ZN(n206) );
  AND3_X1 U159 ( .A1(n267), .A2(n268), .A3(n269), .ZN(product[15]) );
  XNOR2_X1 U160 ( .A(n208), .B(n241), .ZN(product[6]) );
  XNOR2_X1 U161 ( .A(n46), .B(n49), .ZN(n208) );
  NAND2_X1 U162 ( .A1(n216), .A2(n27), .ZN(n209) );
  NAND3_X1 U163 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n210) );
  NAND3_X1 U164 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n211) );
  NAND2_X2 U165 ( .A1(n320), .A2(n339), .ZN(n322) );
  XOR2_X2 U166 ( .A(a[6]), .B(n289), .Z(n320) );
  XOR2_X1 U167 ( .A(n34), .B(n39), .Z(n212) );
  XOR2_X1 U168 ( .A(n211), .B(n212), .Z(product[8]) );
  NAND2_X1 U169 ( .A1(n210), .A2(n34), .ZN(n213) );
  NAND2_X1 U170 ( .A1(n8), .A2(n39), .ZN(n214) );
  NAND2_X1 U171 ( .A1(n34), .A2(n39), .ZN(n215) );
  NAND3_X1 U172 ( .A1(n213), .A2(n214), .A3(n215), .ZN(n7) );
  NAND3_X1 U173 ( .A1(n218), .A2(n219), .A3(n220), .ZN(n216) );
  XOR2_X1 U174 ( .A(n33), .B(n28), .Z(n217) );
  XOR2_X1 U175 ( .A(n7), .B(n217), .Z(product[9]) );
  NAND2_X1 U176 ( .A1(n7), .A2(n33), .ZN(n218) );
  NAND2_X1 U177 ( .A1(n7), .A2(n28), .ZN(n219) );
  NAND2_X1 U178 ( .A1(n33), .A2(n28), .ZN(n220) );
  NAND3_X1 U179 ( .A1(n218), .A2(n219), .A3(n220), .ZN(n6) );
  NAND3_X1 U180 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n221) );
  NAND3_X1 U181 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n222) );
  CLKBUF_X1 U182 ( .A(n12), .Z(n223) );
  NAND3_X1 U183 ( .A1(n209), .A2(n234), .A3(n235), .ZN(n224) );
  NAND3_X1 U184 ( .A1(n209), .A2(n234), .A3(n235), .ZN(n225) );
  NAND3_X1 U185 ( .A1(n245), .A2(n244), .A3(n243), .ZN(n226) );
  XNOR2_X1 U186 ( .A(n2), .B(n206), .ZN(product[14]) );
  CLKBUF_X1 U187 ( .A(b[1]), .Z(n227) );
  XOR2_X1 U188 ( .A(n17), .B(n284), .Z(n228) );
  XOR2_X1 U189 ( .A(n222), .B(n228), .Z(product[13]) );
  NAND2_X1 U190 ( .A1(n221), .A2(n17), .ZN(n229) );
  NAND2_X1 U191 ( .A1(n3), .A2(n284), .ZN(n230) );
  NAND2_X1 U192 ( .A1(n17), .A2(n284), .ZN(n231) );
  NAND3_X1 U193 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n2) );
  XOR2_X1 U194 ( .A(n27), .B(n24), .Z(n232) );
  XOR2_X1 U195 ( .A(n216), .B(n232), .Z(product[10]) );
  NAND2_X1 U196 ( .A1(n216), .A2(n27), .ZN(n233) );
  NAND2_X1 U197 ( .A1(n6), .A2(n24), .ZN(n234) );
  NAND2_X1 U198 ( .A1(n27), .A2(n24), .ZN(n235) );
  NAND3_X1 U199 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n5) );
  CLKBUF_X1 U200 ( .A(n257), .Z(n236) );
  NAND3_X1 U201 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n237) );
  NAND3_X1 U202 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n238) );
  CLKBUF_X1 U203 ( .A(b[1]), .Z(n239) );
  NAND3_X1 U204 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n240) );
  NAND3_X1 U205 ( .A1(n256), .A2(n236), .A3(n258), .ZN(n241) );
  XOR2_X1 U206 ( .A(n20), .B(n23), .Z(n242) );
  XOR2_X1 U207 ( .A(n242), .B(n225), .Z(product[11]) );
  NAND2_X1 U208 ( .A1(n20), .A2(n23), .ZN(n243) );
  NAND2_X1 U209 ( .A1(n20), .A2(n5), .ZN(n244) );
  NAND2_X1 U210 ( .A1(n23), .A2(n224), .ZN(n245) );
  NAND3_X1 U211 ( .A1(n245), .A2(n244), .A3(n243), .ZN(n4) );
  XOR2_X1 U212 ( .A(n19), .B(n18), .Z(n246) );
  XOR2_X1 U213 ( .A(n246), .B(n226), .Z(product[12]) );
  NAND2_X1 U214 ( .A1(n19), .A2(n18), .ZN(n247) );
  NAND2_X1 U215 ( .A1(n19), .A2(n4), .ZN(n248) );
  NAND2_X1 U216 ( .A1(n18), .A2(n4), .ZN(n249) );
  NAND3_X1 U217 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n3) );
  XOR2_X1 U218 ( .A(n54), .B(n55), .Z(n250) );
  XOR2_X1 U219 ( .A(n223), .B(n250), .Z(product[4]) );
  NAND2_X1 U220 ( .A1(n12), .A2(n54), .ZN(n251) );
  NAND2_X1 U221 ( .A1(n12), .A2(n55), .ZN(n252) );
  NAND2_X1 U222 ( .A1(n54), .A2(n55), .ZN(n253) );
  NAND3_X1 U223 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n11) );
  NAND3_X1 U224 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n254) );
  XOR2_X1 U225 ( .A(n50), .B(n53), .Z(n255) );
  XOR2_X1 U226 ( .A(n238), .B(n255), .Z(product[5]) );
  NAND2_X1 U227 ( .A1(n237), .A2(n50), .ZN(n256) );
  NAND2_X1 U228 ( .A1(n11), .A2(n53), .ZN(n257) );
  NAND2_X1 U229 ( .A1(n50), .A2(n53), .ZN(n258) );
  NAND3_X1 U230 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n10) );
  INV_X1 U231 ( .A(n283), .ZN(n259) );
  INV_X1 U232 ( .A(n283), .ZN(n282) );
  NAND2_X2 U233 ( .A1(n299), .A2(n337), .ZN(n301) );
  NAND2_X1 U234 ( .A1(n46), .A2(n49), .ZN(n260) );
  NAND2_X1 U235 ( .A1(n46), .A2(n240), .ZN(n261) );
  NAND2_X1 U236 ( .A1(n49), .A2(n10), .ZN(n262) );
  NAND3_X1 U237 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n9) );
  XOR2_X1 U238 ( .A(n40), .B(n45), .Z(n263) );
  XOR2_X1 U239 ( .A(n263), .B(n254), .Z(product[7]) );
  NAND2_X1 U240 ( .A1(n40), .A2(n45), .ZN(n264) );
  NAND2_X1 U241 ( .A1(n40), .A2(n9), .ZN(n265) );
  NAND2_X1 U242 ( .A1(n45), .A2(n9), .ZN(n266) );
  NAND3_X1 U243 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n8) );
  NAND2_X1 U244 ( .A1(n2), .A2(n285), .ZN(n267) );
  NAND2_X1 U245 ( .A1(n2), .A2(n15), .ZN(n268) );
  NAND2_X1 U246 ( .A1(n285), .A2(n15), .ZN(n269) );
  NAND2_X1 U247 ( .A1(a[4]), .A2(a[3]), .ZN(n272) );
  NAND2_X1 U248 ( .A1(n270), .A2(n271), .ZN(n273) );
  NAND2_X2 U249 ( .A1(n272), .A2(n273), .ZN(n309) );
  INV_X1 U250 ( .A(a[4]), .ZN(n270) );
  INV_X1 U251 ( .A(a[3]), .ZN(n271) );
  NAND2_X2 U252 ( .A1(n309), .A2(n338), .ZN(n311) );
  INV_X1 U253 ( .A(a[0]), .ZN(n293) );
  OR2_X1 U254 ( .A1(n295), .A2(n340), .ZN(n274) );
  OR2_X1 U255 ( .A1(n341), .A2(n293), .ZN(n275) );
  NAND2_X1 U256 ( .A1(n274), .A2(n275), .ZN(n103) );
  INV_X1 U257 ( .A(n299), .ZN(n276) );
  INV_X1 U258 ( .A(n276), .ZN(n277) );
  NAND2_X1 U259 ( .A1(n280), .A2(n281), .ZN(n299) );
  NAND2_X1 U260 ( .A1(a[2]), .A2(a[1]), .ZN(n280) );
  NAND2_X1 U261 ( .A1(n278), .A2(n279), .ZN(n281) );
  INV_X1 U262 ( .A(a[2]), .ZN(n278) );
  INV_X1 U263 ( .A(a[1]), .ZN(n279) );
  INV_X1 U264 ( .A(n21), .ZN(n287) );
  INV_X1 U265 ( .A(n318), .ZN(n288) );
  INV_X1 U266 ( .A(n329), .ZN(n285) );
  INV_X1 U267 ( .A(b[0]), .ZN(n283) );
  INV_X1 U268 ( .A(n298), .ZN(n292) );
  INV_X1 U269 ( .A(n307), .ZN(n291) );
  INV_X1 U270 ( .A(n31), .ZN(n290) );
  INV_X1 U271 ( .A(a[5]), .ZN(n289) );
  INV_X1 U272 ( .A(a[7]), .ZN(n286) );
  NOR2_X1 U273 ( .A1(n293), .A2(n283), .ZN(product[0]) );
  OAI22_X1 U274 ( .A1(n294), .A2(n295), .B1(n296), .B2(n293), .ZN(n99) );
  OAI22_X1 U275 ( .A1(n296), .A2(n295), .B1(n297), .B2(n293), .ZN(n98) );
  XNOR2_X1 U276 ( .A(b[6]), .B(a[1]), .ZN(n296) );
  OAI22_X1 U277 ( .A1(n293), .A2(n297), .B1(n295), .B2(n297), .ZN(n298) );
  XNOR2_X1 U278 ( .A(b[7]), .B(a[1]), .ZN(n297) );
  NOR2_X1 U279 ( .A1(n299), .A2(n283), .ZN(n96) );
  OAI22_X1 U280 ( .A1(n300), .A2(n301), .B1(n299), .B2(n302), .ZN(n95) );
  XNOR2_X1 U281 ( .A(a[3]), .B(n282), .ZN(n300) );
  OAI22_X1 U282 ( .A1(n302), .A2(n301), .B1(n277), .B2(n303), .ZN(n94) );
  XNOR2_X1 U283 ( .A(n227), .B(a[3]), .ZN(n302) );
  OAI22_X1 U284 ( .A1(n303), .A2(n301), .B1(n277), .B2(n304), .ZN(n93) );
  XNOR2_X1 U285 ( .A(b[2]), .B(a[3]), .ZN(n303) );
  OAI22_X1 U286 ( .A1(n304), .A2(n301), .B1(n277), .B2(n305), .ZN(n92) );
  XNOR2_X1 U287 ( .A(b[3]), .B(a[3]), .ZN(n304) );
  OAI22_X1 U288 ( .A1(n305), .A2(n301), .B1(n277), .B2(n306), .ZN(n91) );
  XNOR2_X1 U289 ( .A(b[4]), .B(a[3]), .ZN(n305) );
  OAI22_X1 U290 ( .A1(n308), .A2(n277), .B1(n301), .B2(n308), .ZN(n307) );
  NOR2_X1 U291 ( .A1(n309), .A2(n283), .ZN(n88) );
  OAI22_X1 U292 ( .A1(n310), .A2(n311), .B1(n309), .B2(n312), .ZN(n87) );
  XNOR2_X1 U293 ( .A(a[5]), .B(n259), .ZN(n310) );
  OAI22_X1 U294 ( .A1(n312), .A2(n311), .B1(n309), .B2(n313), .ZN(n86) );
  XNOR2_X1 U295 ( .A(n239), .B(a[5]), .ZN(n312) );
  OAI22_X1 U296 ( .A1(n313), .A2(n311), .B1(n309), .B2(n314), .ZN(n85) );
  XNOR2_X1 U297 ( .A(b[2]), .B(a[5]), .ZN(n313) );
  OAI22_X1 U298 ( .A1(n314), .A2(n311), .B1(n309), .B2(n315), .ZN(n84) );
  XNOR2_X1 U299 ( .A(b[3]), .B(a[5]), .ZN(n314) );
  OAI22_X1 U300 ( .A1(n315), .A2(n311), .B1(n309), .B2(n316), .ZN(n83) );
  XNOR2_X1 U301 ( .A(b[4]), .B(a[5]), .ZN(n315) );
  OAI22_X1 U302 ( .A1(n316), .A2(n311), .B1(n309), .B2(n317), .ZN(n82) );
  XNOR2_X1 U303 ( .A(b[5]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U304 ( .A1(n319), .A2(n309), .B1(n311), .B2(n319), .ZN(n318) );
  NOR2_X1 U305 ( .A1(n320), .A2(n283), .ZN(n80) );
  OAI22_X1 U306 ( .A1(n321), .A2(n322), .B1(n320), .B2(n323), .ZN(n79) );
  XNOR2_X1 U307 ( .A(a[7]), .B(n259), .ZN(n321) );
  OAI22_X1 U308 ( .A1(n324), .A2(n322), .B1(n320), .B2(n325), .ZN(n77) );
  OAI22_X1 U309 ( .A1(n325), .A2(n322), .B1(n320), .B2(n326), .ZN(n76) );
  XNOR2_X1 U310 ( .A(b[3]), .B(a[7]), .ZN(n325) );
  OAI22_X1 U311 ( .A1(n326), .A2(n322), .B1(n320), .B2(n327), .ZN(n75) );
  XNOR2_X1 U312 ( .A(b[4]), .B(a[7]), .ZN(n326) );
  OAI22_X1 U313 ( .A1(n327), .A2(n322), .B1(n320), .B2(n328), .ZN(n74) );
  XNOR2_X1 U314 ( .A(b[5]), .B(a[7]), .ZN(n327) );
  OAI22_X1 U315 ( .A1(n330), .A2(n320), .B1(n322), .B2(n330), .ZN(n329) );
  OAI21_X1 U316 ( .B1(n282), .B2(n279), .A(n295), .ZN(n72) );
  OAI21_X1 U317 ( .B1(n271), .B2(n301), .A(n331), .ZN(n71) );
  OR3_X1 U318 ( .A1(n299), .A2(n259), .A3(n271), .ZN(n331) );
  OAI21_X1 U319 ( .B1(n289), .B2(n311), .A(n332), .ZN(n70) );
  OR3_X1 U320 ( .A1(n309), .A2(n282), .A3(n289), .ZN(n332) );
  OAI21_X1 U321 ( .B1(n286), .B2(n322), .A(n333), .ZN(n69) );
  OR3_X1 U322 ( .A1(n320), .A2(n259), .A3(n286), .ZN(n333) );
  XNOR2_X1 U323 ( .A(n334), .B(n335), .ZN(n38) );
  OR2_X1 U324 ( .A1(n334), .A2(n335), .ZN(n37) );
  OAI22_X1 U325 ( .A1(n306), .A2(n301), .B1(n277), .B2(n336), .ZN(n335) );
  XNOR2_X1 U326 ( .A(b[5]), .B(a[3]), .ZN(n306) );
  OAI22_X1 U327 ( .A1(n323), .A2(n322), .B1(n320), .B2(n324), .ZN(n334) );
  XNOR2_X1 U328 ( .A(b[2]), .B(a[7]), .ZN(n324) );
  XNOR2_X1 U329 ( .A(n239), .B(a[7]), .ZN(n323) );
  OAI22_X1 U330 ( .A1(n336), .A2(n301), .B1(n277), .B2(n308), .ZN(n31) );
  XNOR2_X1 U331 ( .A(b[7]), .B(a[3]), .ZN(n308) );
  XNOR2_X1 U332 ( .A(n271), .B(a[2]), .ZN(n337) );
  XNOR2_X1 U333 ( .A(b[6]), .B(a[3]), .ZN(n336) );
  OAI22_X1 U334 ( .A1(n317), .A2(n311), .B1(n309), .B2(n319), .ZN(n21) );
  XNOR2_X1 U335 ( .A(b[7]), .B(a[5]), .ZN(n319) );
  XNOR2_X1 U336 ( .A(n289), .B(a[4]), .ZN(n338) );
  XNOR2_X1 U337 ( .A(b[6]), .B(a[5]), .ZN(n317) );
  OAI22_X1 U338 ( .A1(n328), .A2(n322), .B1(n320), .B2(n330), .ZN(n15) );
  XNOR2_X1 U339 ( .A(b[7]), .B(a[7]), .ZN(n330) );
  XNOR2_X1 U340 ( .A(n286), .B(a[6]), .ZN(n339) );
  XNOR2_X1 U341 ( .A(b[6]), .B(a[7]), .ZN(n328) );
  OAI22_X1 U342 ( .A1(n282), .A2(n295), .B1(n340), .B2(n293), .ZN(n104) );
  XNOR2_X1 U343 ( .A(b[1]), .B(a[1]), .ZN(n340) );
  OAI22_X1 U344 ( .A1(n341), .A2(n295), .B1(n342), .B2(n293), .ZN(n102) );
  XNOR2_X1 U345 ( .A(b[2]), .B(a[1]), .ZN(n341) );
  OAI22_X1 U346 ( .A1(n342), .A2(n295), .B1(n343), .B2(n293), .ZN(n101) );
  XNOR2_X1 U347 ( .A(b[3]), .B(a[1]), .ZN(n342) );
  OAI22_X1 U348 ( .A1(n343), .A2(n295), .B1(n294), .B2(n293), .ZN(n100) );
  XNOR2_X1 U349 ( .A(b[5]), .B(a[1]), .ZN(n294) );
  NAND2_X1 U350 ( .A1(a[1]), .A2(n293), .ZN(n295) );
  XNOR2_X1 U351 ( .A(b[4]), .B(a[1]), .ZN(n343) );
endmodule


module datapath_DW01_add_26 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n79;
  wire   [15:1] carry;

  FA_X1 U1_1 ( .A(A[1]), .B(n79), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[14]), .ZN(n30) );
  XNOR2_X1 U2 ( .A(n53), .B(n1), .ZN(SUM[14]) );
  AND3_X1 U3 ( .A1(n50), .A2(n51), .A3(n52), .ZN(n1) );
  CLKBUF_X1 U4 ( .A(B[4]), .Z(n2) );
  CLKBUF_X1 U5 ( .A(n77), .Z(n3) );
  XOR2_X1 U6 ( .A(carry[2]), .B(A[2]), .Z(n4) );
  XOR2_X1 U7 ( .A(B[2]), .B(n4), .Z(SUM[2]) );
  NAND2_X1 U8 ( .A1(B[2]), .A2(carry[2]), .ZN(n5) );
  NAND2_X1 U9 ( .A1(B[2]), .A2(A[2]), .ZN(n6) );
  NAND2_X1 U10 ( .A1(carry[2]), .A2(A[2]), .ZN(n7) );
  NAND3_X1 U11 ( .A1(n5), .A2(n6), .A3(n7), .ZN(carry[3]) );
  NAND3_X1 U12 ( .A1(n76), .A2(n77), .A3(n75), .ZN(n8) );
  CLKBUF_X1 U13 ( .A(n72), .Z(n9) );
  NAND3_X1 U14 ( .A1(n32), .A2(n33), .A3(n34), .ZN(n10) );
  NAND3_X1 U15 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n11) );
  NAND3_X1 U16 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n12) );
  CLKBUF_X1 U17 ( .A(n22), .Z(n13) );
  CLKBUF_X1 U18 ( .A(n10), .Z(n14) );
  NAND3_X1 U19 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n15) );
  CLKBUF_X1 U20 ( .A(n11), .Z(n16) );
  NAND3_X1 U21 ( .A1(n39), .A2(n38), .A3(n40), .ZN(n17) );
  NAND3_X1 U22 ( .A1(n66), .A2(n67), .A3(n68), .ZN(n18) );
  NAND3_X1 U23 ( .A1(n66), .A2(n67), .A3(n68), .ZN(n19) );
  XOR2_X1 U24 ( .A(B[11]), .B(A[11]), .Z(n20) );
  XOR2_X1 U25 ( .A(n14), .B(n20), .Z(SUM[11]) );
  NAND2_X1 U26 ( .A1(carry[11]), .A2(B[11]), .ZN(n21) );
  NAND2_X1 U27 ( .A1(n10), .A2(A[11]), .ZN(n22) );
  NAND2_X1 U28 ( .A1(B[11]), .A2(A[11]), .ZN(n23) );
  NAND3_X1 U29 ( .A1(n21), .A2(n13), .A3(n23), .ZN(carry[12]) );
  XOR2_X1 U30 ( .A(n19), .B(A[9]), .Z(n24) );
  XOR2_X1 U31 ( .A(B[9]), .B(n24), .Z(SUM[9]) );
  NAND2_X1 U32 ( .A1(B[9]), .A2(n18), .ZN(n25) );
  NAND2_X1 U33 ( .A1(B[9]), .A2(A[9]), .ZN(n26) );
  NAND2_X1 U34 ( .A1(carry[9]), .A2(A[9]), .ZN(n27) );
  NAND3_X1 U35 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[10]) );
  NAND3_X1 U36 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n28) );
  NAND3_X1 U37 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n29) );
  XNOR2_X1 U38 ( .A(B[14]), .B(n30), .ZN(n53) );
  XOR2_X1 U39 ( .A(B[10]), .B(A[10]), .Z(n31) );
  XOR2_X1 U40 ( .A(n16), .B(n31), .Z(SUM[10]) );
  NAND2_X1 U41 ( .A1(n11), .A2(B[10]), .ZN(n32) );
  NAND2_X1 U42 ( .A1(carry[10]), .A2(A[10]), .ZN(n33) );
  NAND2_X1 U43 ( .A1(B[10]), .A2(A[10]), .ZN(n34) );
  NAND3_X1 U44 ( .A1(n32), .A2(n33), .A3(n34), .ZN(carry[11]) );
  NAND3_X1 U45 ( .A1(n50), .A2(n51), .A3(n52), .ZN(n35) );
  NAND3_X1 U46 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n36) );
  XOR2_X1 U47 ( .A(B[3]), .B(A[3]), .Z(n37) );
  XOR2_X1 U48 ( .A(carry[3]), .B(n37), .Z(SUM[3]) );
  NAND2_X1 U49 ( .A1(carry[3]), .A2(B[3]), .ZN(n38) );
  NAND2_X1 U50 ( .A1(carry[3]), .A2(A[3]), .ZN(n39) );
  NAND2_X1 U51 ( .A1(B[3]), .A2(A[3]), .ZN(n40) );
  NAND3_X1 U52 ( .A1(n38), .A2(n39), .A3(n40), .ZN(carry[4]) );
  XOR2_X1 U53 ( .A(n2), .B(A[4]), .Z(n41) );
  XOR2_X1 U54 ( .A(carry[4]), .B(n41), .Z(SUM[4]) );
  NAND2_X1 U55 ( .A1(n17), .A2(B[4]), .ZN(n42) );
  NAND2_X1 U56 ( .A1(carry[4]), .A2(A[4]), .ZN(n43) );
  NAND2_X1 U57 ( .A1(B[4]), .A2(A[4]), .ZN(n44) );
  NAND3_X1 U58 ( .A1(n42), .A2(n43), .A3(n44), .ZN(carry[5]) );
  XOR2_X1 U59 ( .A(B[12]), .B(A[12]), .Z(n45) );
  XOR2_X1 U60 ( .A(carry[12]), .B(n45), .Z(SUM[12]) );
  NAND2_X1 U61 ( .A1(n15), .A2(B[12]), .ZN(n46) );
  NAND2_X1 U62 ( .A1(n15), .A2(A[12]), .ZN(n47) );
  NAND2_X1 U63 ( .A1(B[12]), .A2(A[12]), .ZN(n48) );
  NAND3_X1 U64 ( .A1(n46), .A2(n47), .A3(n48), .ZN(carry[13]) );
  XOR2_X1 U65 ( .A(B[13]), .B(A[13]), .Z(n49) );
  XOR2_X1 U66 ( .A(n49), .B(n29), .Z(SUM[13]) );
  NAND2_X1 U67 ( .A1(B[13]), .A2(A[13]), .ZN(n50) );
  NAND2_X1 U68 ( .A1(B[13]), .A2(n28), .ZN(n51) );
  NAND2_X1 U69 ( .A1(A[13]), .A2(carry[13]), .ZN(n52) );
  NAND3_X1 U70 ( .A1(n50), .A2(n51), .A3(n52), .ZN(carry[14]) );
  NAND2_X1 U71 ( .A1(B[14]), .A2(A[14]), .ZN(n54) );
  NAND2_X1 U72 ( .A1(A[14]), .A2(carry[14]), .ZN(n55) );
  NAND2_X1 U73 ( .A1(n35), .A2(B[14]), .ZN(n56) );
  NAND3_X1 U74 ( .A1(n55), .A2(n54), .A3(n56), .ZN(carry[15]) );
  XOR2_X1 U75 ( .A(B[5]), .B(A[5]), .Z(n57) );
  XOR2_X1 U76 ( .A(n12), .B(n57), .Z(SUM[5]) );
  NAND2_X1 U77 ( .A1(n12), .A2(B[5]), .ZN(n58) );
  NAND2_X1 U78 ( .A1(carry[5]), .A2(A[5]), .ZN(n59) );
  NAND2_X1 U79 ( .A1(B[5]), .A2(A[5]), .ZN(n60) );
  NAND3_X1 U80 ( .A1(n59), .A2(n58), .A3(n60), .ZN(carry[6]) );
  XNOR2_X1 U81 ( .A(carry[15]), .B(n61), .ZN(SUM[15]) );
  XNOR2_X1 U82 ( .A(B[15]), .B(A[15]), .ZN(n61) );
  NAND3_X1 U83 ( .A1(n76), .A2(n77), .A3(n75), .ZN(n62) );
  NAND3_X1 U84 ( .A1(n71), .A2(n72), .A3(n73), .ZN(n63) );
  NAND3_X1 U85 ( .A1(n71), .A2(n9), .A3(n73), .ZN(n64) );
  XOR2_X1 U86 ( .A(B[8]), .B(A[8]), .Z(n65) );
  XOR2_X1 U87 ( .A(carry[8]), .B(n65), .Z(SUM[8]) );
  NAND2_X1 U88 ( .A1(n8), .A2(B[8]), .ZN(n66) );
  NAND2_X1 U89 ( .A1(n62), .A2(A[8]), .ZN(n67) );
  NAND2_X1 U90 ( .A1(B[8]), .A2(A[8]), .ZN(n68) );
  NAND3_X1 U91 ( .A1(n66), .A2(n67), .A3(n68), .ZN(carry[9]) );
  CLKBUF_X1 U92 ( .A(n36), .Z(n69) );
  XOR2_X1 U93 ( .A(A[6]), .B(B[6]), .Z(n70) );
  XOR2_X1 U94 ( .A(n70), .B(n69), .Z(SUM[6]) );
  NAND2_X1 U95 ( .A1(A[6]), .A2(B[6]), .ZN(n71) );
  NAND2_X1 U96 ( .A1(A[6]), .A2(n36), .ZN(n72) );
  NAND2_X1 U97 ( .A1(B[6]), .A2(carry[6]), .ZN(n73) );
  NAND3_X1 U98 ( .A1(n71), .A2(n72), .A3(n73), .ZN(carry[7]) );
  XOR2_X1 U99 ( .A(A[7]), .B(B[7]), .Z(n74) );
  XOR2_X1 U100 ( .A(n74), .B(n64), .Z(SUM[7]) );
  NAND2_X1 U101 ( .A1(A[7]), .A2(B[7]), .ZN(n75) );
  NAND2_X1 U102 ( .A1(A[7]), .A2(n63), .ZN(n76) );
  NAND2_X1 U103 ( .A1(B[7]), .A2(carry[7]), .ZN(n77) );
  NAND3_X1 U104 ( .A1(n75), .A2(n76), .A3(n3), .ZN(carry[8]) );
  XOR2_X1 U105 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U106 ( .A1(B[0]), .A2(A[0]), .ZN(n79) );
endmodule


module datapath_DW_mult_tc_25 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345;

  FA_X1 U13 ( .A(n13), .B(n71), .CI(n56), .CO(n12), .S(product[3]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n288), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n287), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n291), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n290), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n293), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  NAND2_X1 U157 ( .A1(n17), .A2(n284), .ZN(n211) );
  AND3_X1 U158 ( .A1(n215), .A2(n216), .A3(n217), .ZN(product[15]) );
  CLKBUF_X1 U159 ( .A(n7), .Z(n207) );
  NAND3_X1 U160 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n208) );
  NAND3_X1 U161 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n209) );
  XOR2_X1 U162 ( .A(n17), .B(n284), .Z(n210) );
  XOR2_X1 U163 ( .A(n210), .B(n209), .Z(product[13]) );
  NAND2_X1 U164 ( .A1(n17), .A2(n208), .ZN(n212) );
  NAND2_X1 U165 ( .A1(n284), .A2(n3), .ZN(n213) );
  NAND3_X1 U166 ( .A1(n211), .A2(n212), .A3(n213), .ZN(n2) );
  XOR2_X1 U167 ( .A(n285), .B(n15), .Z(n214) );
  XOR2_X1 U168 ( .A(n214), .B(n2), .Z(product[14]) );
  NAND2_X1 U169 ( .A1(n285), .A2(n15), .ZN(n215) );
  NAND2_X1 U170 ( .A1(n285), .A2(n2), .ZN(n216) );
  NAND2_X1 U171 ( .A1(n15), .A2(n2), .ZN(n217) );
  NAND3_X1 U172 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n218) );
  XOR2_X2 U173 ( .A(a[6]), .B(n289), .Z(n322) );
  NAND3_X1 U174 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n219) );
  CLKBUF_X1 U175 ( .A(n223), .Z(n220) );
  INV_X1 U176 ( .A(n283), .ZN(n221) );
  CLKBUF_X1 U177 ( .A(n12), .Z(n222) );
  NAND3_X1 U178 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n223) );
  XOR2_X1 U179 ( .A(n54), .B(n55), .Z(n224) );
  XOR2_X1 U180 ( .A(n222), .B(n224), .Z(product[4]) );
  NAND2_X1 U181 ( .A1(n12), .A2(n54), .ZN(n225) );
  NAND2_X1 U182 ( .A1(n12), .A2(n55), .ZN(n226) );
  NAND2_X1 U183 ( .A1(n54), .A2(n55), .ZN(n227) );
  NAND3_X1 U184 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n11) );
  NAND3_X1 U185 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n228) );
  NAND3_X1 U186 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n229) );
  CLKBUF_X1 U187 ( .A(n303), .Z(n230) );
  NAND2_X1 U188 ( .A1(n301), .A2(n339), .ZN(n303) );
  NAND3_X1 U189 ( .A1(n251), .A2(n252), .A3(n250), .ZN(n231) );
  NAND3_X1 U190 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n232) );
  NAND3_X1 U191 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n233) );
  INV_X1 U192 ( .A(n283), .ZN(n234) );
  XOR2_X1 U193 ( .A(n33), .B(n28), .Z(n235) );
  XOR2_X1 U194 ( .A(n207), .B(n235), .Z(product[9]) );
  NAND2_X1 U195 ( .A1(n7), .A2(n33), .ZN(n236) );
  NAND2_X1 U196 ( .A1(n7), .A2(n28), .ZN(n237) );
  NAND2_X1 U197 ( .A1(n33), .A2(n28), .ZN(n238) );
  NAND3_X1 U198 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n6) );
  XOR2_X1 U199 ( .A(n50), .B(n53), .Z(n239) );
  XOR2_X1 U200 ( .A(n220), .B(n239), .Z(product[5]) );
  NAND2_X1 U201 ( .A1(n223), .A2(n50), .ZN(n240) );
  NAND2_X1 U202 ( .A1(n11), .A2(n53), .ZN(n241) );
  NAND2_X1 U203 ( .A1(n50), .A2(n53), .ZN(n242) );
  NAND3_X1 U204 ( .A1(n246), .A2(n245), .A3(n247), .ZN(n243) );
  XOR2_X1 U205 ( .A(n27), .B(n24), .Z(n244) );
  XOR2_X1 U206 ( .A(n229), .B(n244), .Z(product[10]) );
  NAND2_X1 U207 ( .A1(n228), .A2(n27), .ZN(n245) );
  NAND2_X1 U208 ( .A1(n6), .A2(n24), .ZN(n246) );
  NAND2_X1 U209 ( .A1(n27), .A2(n24), .ZN(n247) );
  NAND3_X1 U210 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n5) );
  NAND3_X1 U211 ( .A1(n252), .A2(n251), .A3(n250), .ZN(n248) );
  XOR2_X1 U212 ( .A(n20), .B(n23), .Z(n249) );
  XOR2_X1 U213 ( .A(n249), .B(n219), .Z(product[11]) );
  NAND2_X1 U214 ( .A1(n20), .A2(n23), .ZN(n250) );
  NAND2_X1 U215 ( .A1(n20), .A2(n5), .ZN(n251) );
  NAND2_X1 U216 ( .A1(n23), .A2(n243), .ZN(n252) );
  NAND3_X1 U217 ( .A1(n251), .A2(n250), .A3(n252), .ZN(n4) );
  XOR2_X1 U218 ( .A(n19), .B(n18), .Z(n253) );
  XOR2_X1 U219 ( .A(n253), .B(n231), .Z(product[12]) );
  NAND2_X1 U220 ( .A1(n19), .A2(n18), .ZN(n254) );
  NAND2_X1 U221 ( .A1(n19), .A2(n248), .ZN(n255) );
  NAND2_X1 U222 ( .A1(n18), .A2(n4), .ZN(n256) );
  NAND3_X1 U223 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n3) );
  NAND3_X1 U224 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n257) );
  XOR2_X1 U225 ( .A(n34), .B(n39), .Z(n258) );
  XOR2_X1 U226 ( .A(n257), .B(n258), .Z(product[8]) );
  NAND2_X1 U227 ( .A1(n257), .A2(n34), .ZN(n259) );
  NAND2_X1 U228 ( .A1(n8), .A2(n39), .ZN(n260) );
  NAND2_X1 U229 ( .A1(n34), .A2(n39), .ZN(n261) );
  NAND3_X1 U230 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n7) );
  NAND3_X1 U231 ( .A1(n267), .A2(n266), .A3(n265), .ZN(n262) );
  NAND3_X1 U232 ( .A1(n267), .A2(n266), .A3(n265), .ZN(n263) );
  XOR2_X1 U233 ( .A(n46), .B(n49), .Z(n264) );
  XOR2_X1 U234 ( .A(n264), .B(n218), .Z(product[6]) );
  NAND2_X1 U235 ( .A1(n46), .A2(n49), .ZN(n265) );
  NAND2_X1 U236 ( .A1(n46), .A2(n232), .ZN(n266) );
  NAND2_X1 U237 ( .A1(n49), .A2(n233), .ZN(n267) );
  NAND3_X1 U238 ( .A1(n266), .A2(n265), .A3(n267), .ZN(n9) );
  XOR2_X1 U239 ( .A(n40), .B(n45), .Z(n268) );
  XOR2_X1 U240 ( .A(n268), .B(n263), .Z(product[7]) );
  NAND2_X1 U241 ( .A1(n40), .A2(n45), .ZN(n269) );
  NAND2_X1 U242 ( .A1(n40), .A2(n262), .ZN(n270) );
  NAND2_X1 U243 ( .A1(n45), .A2(n9), .ZN(n271) );
  NAND3_X1 U244 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n8) );
  XOR2_X1 U245 ( .A(n103), .B(n96), .Z(n272) );
  XOR2_X1 U246 ( .A(n272), .B(n14), .Z(product[2]) );
  NAND2_X1 U247 ( .A1(n14), .A2(n103), .ZN(n273) );
  NAND2_X1 U248 ( .A1(n14), .A2(n96), .ZN(n274) );
  NAND2_X1 U249 ( .A1(n103), .A2(n96), .ZN(n275) );
  NAND3_X1 U250 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n13) );
  NAND2_X1 U251 ( .A1(a[4]), .A2(a[3]), .ZN(n278) );
  NAND2_X1 U252 ( .A1(n276), .A2(n277), .ZN(n279) );
  NAND2_X2 U253 ( .A1(n278), .A2(n279), .ZN(n311) );
  INV_X1 U254 ( .A(a[4]), .ZN(n276) );
  INV_X1 U255 ( .A(a[3]), .ZN(n277) );
  NAND2_X2 U256 ( .A1(n311), .A2(n340), .ZN(n313) );
  BUF_X1 U257 ( .A(n301), .Z(n281) );
  CLKBUF_X1 U258 ( .A(n301), .Z(n280) );
  XNOR2_X1 U259 ( .A(a[2]), .B(a[1]), .ZN(n301) );
  INV_X1 U260 ( .A(n15), .ZN(n284) );
  INV_X1 U261 ( .A(n21), .ZN(n287) );
  INV_X1 U262 ( .A(n320), .ZN(n288) );
  INV_X1 U263 ( .A(n331), .ZN(n285) );
  INV_X1 U264 ( .A(b[0]), .ZN(n283) );
  INV_X1 U265 ( .A(n300), .ZN(n293) );
  INV_X1 U266 ( .A(n309), .ZN(n291) );
  INV_X1 U267 ( .A(n31), .ZN(n290) );
  INV_X1 U268 ( .A(a[0]), .ZN(n295) );
  INV_X1 U269 ( .A(a[5]), .ZN(n289) );
  INV_X1 U270 ( .A(a[7]), .ZN(n286) );
  XNOR2_X1 U271 ( .A(a[1]), .B(b[1]), .ZN(n282) );
  INV_X1 U272 ( .A(a[3]), .ZN(n292) );
  INV_X1 U273 ( .A(a[1]), .ZN(n294) );
  NOR2_X1 U274 ( .A1(n295), .A2(n283), .ZN(product[0]) );
  OAI22_X1 U275 ( .A1(n296), .A2(n297), .B1(n298), .B2(n295), .ZN(n99) );
  OAI22_X1 U276 ( .A1(n298), .A2(n297), .B1(n299), .B2(n295), .ZN(n98) );
  XNOR2_X1 U277 ( .A(b[6]), .B(a[1]), .ZN(n298) );
  OAI22_X1 U278 ( .A1(n295), .A2(n299), .B1(n297), .B2(n299), .ZN(n300) );
  XNOR2_X1 U279 ( .A(b[7]), .B(a[1]), .ZN(n299) );
  NOR2_X1 U280 ( .A1(n281), .A2(n283), .ZN(n96) );
  OAI22_X1 U281 ( .A1(n302), .A2(n303), .B1(n280), .B2(n304), .ZN(n95) );
  XNOR2_X1 U282 ( .A(a[3]), .B(n234), .ZN(n302) );
  OAI22_X1 U283 ( .A1(n304), .A2(n303), .B1(n281), .B2(n305), .ZN(n94) );
  XNOR2_X1 U284 ( .A(b[1]), .B(a[3]), .ZN(n304) );
  OAI22_X1 U285 ( .A1(n305), .A2(n303), .B1(n281), .B2(n306), .ZN(n93) );
  XNOR2_X1 U286 ( .A(b[2]), .B(a[3]), .ZN(n305) );
  OAI22_X1 U287 ( .A1(n306), .A2(n303), .B1(n280), .B2(n307), .ZN(n92) );
  XNOR2_X1 U288 ( .A(b[3]), .B(a[3]), .ZN(n306) );
  OAI22_X1 U289 ( .A1(n307), .A2(n230), .B1(n280), .B2(n308), .ZN(n91) );
  XNOR2_X1 U290 ( .A(b[4]), .B(a[3]), .ZN(n307) );
  OAI22_X1 U291 ( .A1(n310), .A2(n281), .B1(n230), .B2(n310), .ZN(n309) );
  NOR2_X1 U292 ( .A1(n311), .A2(n283), .ZN(n88) );
  OAI22_X1 U293 ( .A1(n312), .A2(n313), .B1(n311), .B2(n314), .ZN(n87) );
  XNOR2_X1 U294 ( .A(a[5]), .B(n234), .ZN(n312) );
  OAI22_X1 U295 ( .A1(n314), .A2(n313), .B1(n311), .B2(n315), .ZN(n86) );
  XNOR2_X1 U296 ( .A(b[1]), .B(a[5]), .ZN(n314) );
  OAI22_X1 U297 ( .A1(n315), .A2(n313), .B1(n311), .B2(n316), .ZN(n85) );
  XNOR2_X1 U298 ( .A(b[2]), .B(a[5]), .ZN(n315) );
  OAI22_X1 U299 ( .A1(n316), .A2(n313), .B1(n311), .B2(n317), .ZN(n84) );
  XNOR2_X1 U300 ( .A(b[3]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U301 ( .A1(n317), .A2(n313), .B1(n311), .B2(n318), .ZN(n83) );
  XNOR2_X1 U302 ( .A(b[4]), .B(a[5]), .ZN(n317) );
  OAI22_X1 U303 ( .A1(n318), .A2(n313), .B1(n311), .B2(n319), .ZN(n82) );
  XNOR2_X1 U304 ( .A(b[5]), .B(a[5]), .ZN(n318) );
  OAI22_X1 U305 ( .A1(n321), .A2(n311), .B1(n313), .B2(n321), .ZN(n320) );
  NOR2_X1 U306 ( .A1(n322), .A2(n283), .ZN(n80) );
  OAI22_X1 U307 ( .A1(n323), .A2(n324), .B1(n322), .B2(n325), .ZN(n79) );
  XNOR2_X1 U308 ( .A(a[7]), .B(n234), .ZN(n323) );
  OAI22_X1 U309 ( .A1(n326), .A2(n324), .B1(n322), .B2(n327), .ZN(n77) );
  OAI22_X1 U310 ( .A1(n327), .A2(n324), .B1(n322), .B2(n328), .ZN(n76) );
  XNOR2_X1 U311 ( .A(b[3]), .B(a[7]), .ZN(n327) );
  OAI22_X1 U312 ( .A1(n328), .A2(n324), .B1(n322), .B2(n329), .ZN(n75) );
  XNOR2_X1 U313 ( .A(b[4]), .B(a[7]), .ZN(n328) );
  OAI22_X1 U314 ( .A1(n329), .A2(n324), .B1(n322), .B2(n330), .ZN(n74) );
  XNOR2_X1 U315 ( .A(b[5]), .B(a[7]), .ZN(n329) );
  OAI22_X1 U316 ( .A1(n332), .A2(n322), .B1(n324), .B2(n332), .ZN(n331) );
  OAI21_X1 U317 ( .B1(n221), .B2(n294), .A(n297), .ZN(n72) );
  OAI21_X1 U318 ( .B1(n292), .B2(n303), .A(n333), .ZN(n71) );
  OR3_X1 U319 ( .A1(n280), .A2(n234), .A3(n292), .ZN(n333) );
  OAI21_X1 U320 ( .B1(n289), .B2(n313), .A(n334), .ZN(n70) );
  OR3_X1 U321 ( .A1(n311), .A2(n221), .A3(n289), .ZN(n334) );
  OAI21_X1 U322 ( .B1(n286), .B2(n324), .A(n335), .ZN(n69) );
  OR3_X1 U323 ( .A1(n322), .A2(n234), .A3(n286), .ZN(n335) );
  XNOR2_X1 U324 ( .A(n336), .B(n337), .ZN(n38) );
  OR2_X1 U325 ( .A1(n336), .A2(n337), .ZN(n37) );
  OAI22_X1 U326 ( .A1(n308), .A2(n230), .B1(n281), .B2(n338), .ZN(n337) );
  XNOR2_X1 U327 ( .A(b[5]), .B(a[3]), .ZN(n308) );
  OAI22_X1 U328 ( .A1(n325), .A2(n324), .B1(n322), .B2(n326), .ZN(n336) );
  XNOR2_X1 U329 ( .A(b[2]), .B(a[7]), .ZN(n326) );
  XNOR2_X1 U330 ( .A(b[1]), .B(a[7]), .ZN(n325) );
  OAI22_X1 U331 ( .A1(n338), .A2(n230), .B1(n280), .B2(n310), .ZN(n31) );
  XNOR2_X1 U332 ( .A(b[7]), .B(a[3]), .ZN(n310) );
  XNOR2_X1 U333 ( .A(n292), .B(a[2]), .ZN(n339) );
  XNOR2_X1 U334 ( .A(b[6]), .B(a[3]), .ZN(n338) );
  OAI22_X1 U335 ( .A1(n319), .A2(n313), .B1(n311), .B2(n321), .ZN(n21) );
  XNOR2_X1 U336 ( .A(b[7]), .B(a[5]), .ZN(n321) );
  XNOR2_X1 U337 ( .A(n289), .B(a[4]), .ZN(n340) );
  XNOR2_X1 U338 ( .A(b[6]), .B(a[5]), .ZN(n319) );
  OAI22_X1 U339 ( .A1(n330), .A2(n324), .B1(n322), .B2(n332), .ZN(n15) );
  XNOR2_X1 U340 ( .A(b[7]), .B(a[7]), .ZN(n332) );
  NAND2_X1 U341 ( .A1(n322), .A2(n341), .ZN(n324) );
  XNOR2_X1 U342 ( .A(n286), .B(a[6]), .ZN(n341) );
  XNOR2_X1 U343 ( .A(b[6]), .B(a[7]), .ZN(n330) );
  OAI22_X1 U344 ( .A1(n221), .A2(n297), .B1(n342), .B2(n295), .ZN(n104) );
  OAI22_X1 U345 ( .A1(n282), .A2(n297), .B1(n343), .B2(n295), .ZN(n103) );
  XNOR2_X1 U346 ( .A(b[1]), .B(a[1]), .ZN(n342) );
  OAI22_X1 U347 ( .A1(n343), .A2(n297), .B1(n344), .B2(n295), .ZN(n102) );
  XNOR2_X1 U348 ( .A(b[2]), .B(a[1]), .ZN(n343) );
  OAI22_X1 U349 ( .A1(n344), .A2(n297), .B1(n345), .B2(n295), .ZN(n101) );
  XNOR2_X1 U350 ( .A(b[3]), .B(a[1]), .ZN(n344) );
  OAI22_X1 U351 ( .A1(n345), .A2(n297), .B1(n296), .B2(n295), .ZN(n100) );
  XNOR2_X1 U352 ( .A(b[5]), .B(a[1]), .ZN(n296) );
  NAND2_X1 U353 ( .A1(a[1]), .A2(n295), .ZN(n297) );
  XNOR2_X1 U354 ( .A(b[4]), .B(a[1]), .ZN(n345) );
endmodule


module datapath_DW01_add_25 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n69;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_2 ( .A(A[2]), .B(carry[2]), .CI(B[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n69), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  XNOR2_X1 U1 ( .A(B[15]), .B(A[15]), .ZN(n46) );
  CLKBUF_X1 U2 ( .A(B[5]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(carry[3]), .Z(n2) );
  NAND3_X1 U4 ( .A1(n5), .A2(n6), .A3(n7), .ZN(n3) );
  XOR2_X1 U5 ( .A(B[3]), .B(A[3]), .Z(n4) );
  XOR2_X1 U6 ( .A(n2), .B(n4), .Z(SUM[3]) );
  NAND2_X1 U7 ( .A1(carry[3]), .A2(B[3]), .ZN(n5) );
  NAND2_X1 U8 ( .A1(carry[3]), .A2(A[3]), .ZN(n6) );
  NAND2_X1 U9 ( .A1(B[3]), .A2(A[3]), .ZN(n7) );
  NAND3_X1 U10 ( .A1(n5), .A2(n6), .A3(n7), .ZN(carry[4]) );
  NAND3_X1 U11 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n8) );
  NAND3_X1 U12 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n9) );
  CLKBUF_X1 U13 ( .A(n67), .Z(n10) );
  CLKBUF_X1 U14 ( .A(carry[12]), .Z(n11) );
  CLKBUF_X1 U15 ( .A(n66), .Z(n12) );
  XOR2_X1 U16 ( .A(B[11]), .B(A[11]), .Z(n13) );
  XOR2_X1 U17 ( .A(n9), .B(n13), .Z(SUM[11]) );
  NAND2_X1 U18 ( .A1(n8), .A2(B[11]), .ZN(n14) );
  NAND2_X1 U19 ( .A1(carry[11]), .A2(A[11]), .ZN(n15) );
  NAND2_X1 U20 ( .A1(B[11]), .A2(A[11]), .ZN(n16) );
  NAND3_X1 U21 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[12]) );
  NAND3_X1 U22 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n17) );
  NAND3_X1 U23 ( .A1(n22), .A2(n23), .A3(n24), .ZN(n18) );
  NAND3_X1 U24 ( .A1(n22), .A2(n23), .A3(n24), .ZN(n19) );
  NAND3_X1 U25 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n20) );
  XOR2_X1 U26 ( .A(n3), .B(A[4]), .Z(n21) );
  XOR2_X1 U27 ( .A(B[4]), .B(n21), .Z(SUM[4]) );
  NAND2_X1 U28 ( .A1(n3), .A2(B[4]), .ZN(n22) );
  NAND2_X1 U29 ( .A1(B[4]), .A2(A[4]), .ZN(n23) );
  NAND2_X1 U30 ( .A1(carry[4]), .A2(A[4]), .ZN(n24) );
  NAND3_X1 U31 ( .A1(n22), .A2(n23), .A3(n24), .ZN(carry[5]) );
  XOR2_X1 U32 ( .A(n1), .B(A[5]), .Z(n25) );
  XOR2_X1 U33 ( .A(n19), .B(n25), .Z(SUM[5]) );
  NAND2_X1 U34 ( .A1(n18), .A2(B[5]), .ZN(n26) );
  NAND2_X1 U35 ( .A1(carry[5]), .A2(A[5]), .ZN(n27) );
  NAND2_X1 U36 ( .A1(B[5]), .A2(A[5]), .ZN(n28) );
  NAND3_X1 U37 ( .A1(n26), .A2(n27), .A3(n28), .ZN(carry[6]) );
  CLKBUF_X1 U38 ( .A(n20), .Z(n29) );
  NAND3_X1 U39 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n30) );
  NAND3_X1 U40 ( .A1(n65), .A2(n12), .A3(n10), .ZN(n31) );
  XOR2_X1 U41 ( .A(B[10]), .B(A[10]), .Z(n32) );
  XOR2_X1 U42 ( .A(n31), .B(n32), .Z(SUM[10]) );
  NAND2_X1 U43 ( .A1(n30), .A2(B[10]), .ZN(n33) );
  NAND2_X1 U44 ( .A1(carry[10]), .A2(A[10]), .ZN(n34) );
  NAND2_X1 U45 ( .A1(B[10]), .A2(A[10]), .ZN(n35) );
  NAND3_X1 U46 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[11]) );
  CLKBUF_X1 U47 ( .A(n55), .Z(n36) );
  XOR2_X1 U48 ( .A(B[12]), .B(A[12]), .Z(n37) );
  XOR2_X1 U49 ( .A(n11), .B(n37), .Z(SUM[12]) );
  NAND2_X1 U50 ( .A1(carry[12]), .A2(B[12]), .ZN(n38) );
  NAND2_X1 U51 ( .A1(carry[12]), .A2(A[12]), .ZN(n39) );
  NAND2_X1 U52 ( .A1(B[12]), .A2(A[12]), .ZN(n40) );
  NAND3_X1 U53 ( .A1(n38), .A2(n39), .A3(n40), .ZN(carry[13]) );
  NAND3_X1 U54 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n41) );
  XOR2_X1 U55 ( .A(B[13]), .B(A[13]), .Z(n42) );
  XOR2_X1 U56 ( .A(n29), .B(n42), .Z(SUM[13]) );
  NAND2_X1 U57 ( .A1(n20), .A2(B[13]), .ZN(n43) );
  NAND2_X1 U58 ( .A1(carry[13]), .A2(A[13]), .ZN(n44) );
  NAND2_X1 U59 ( .A1(B[13]), .A2(A[13]), .ZN(n45) );
  NAND3_X1 U60 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[14]) );
  XNOR2_X1 U61 ( .A(carry[15]), .B(n46), .ZN(SUM[15]) );
  CLKBUF_X1 U62 ( .A(n62), .Z(n47) );
  XOR2_X1 U63 ( .A(B[6]), .B(A[6]), .Z(n48) );
  XOR2_X1 U64 ( .A(carry[6]), .B(n48), .Z(SUM[6]) );
  NAND2_X1 U65 ( .A1(n17), .A2(B[6]), .ZN(n49) );
  NAND2_X1 U66 ( .A1(carry[6]), .A2(A[6]), .ZN(n50) );
  NAND2_X1 U67 ( .A1(B[6]), .A2(A[6]), .ZN(n51) );
  NAND3_X1 U68 ( .A1(n49), .A2(n50), .A3(n51), .ZN(carry[7]) );
  NAND3_X1 U69 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n52) );
  NAND3_X1 U70 ( .A1(n36), .A2(n56), .A3(n57), .ZN(n53) );
  XOR2_X1 U71 ( .A(B[7]), .B(A[7]), .Z(n54) );
  XOR2_X1 U72 ( .A(n41), .B(n54), .Z(SUM[7]) );
  NAND2_X1 U73 ( .A1(n41), .A2(B[7]), .ZN(n55) );
  NAND2_X1 U74 ( .A1(carry[7]), .A2(A[7]), .ZN(n56) );
  NAND2_X1 U75 ( .A1(B[7]), .A2(A[7]), .ZN(n57) );
  NAND3_X1 U76 ( .A1(n55), .A2(n56), .A3(n57), .ZN(carry[8]) );
  NAND3_X1 U77 ( .A1(n63), .A2(n62), .A3(n61), .ZN(n58) );
  NAND3_X1 U78 ( .A1(n61), .A2(n47), .A3(n63), .ZN(n59) );
  XOR2_X1 U79 ( .A(A[8]), .B(B[8]), .Z(n60) );
  XOR2_X1 U80 ( .A(n60), .B(n53), .Z(SUM[8]) );
  NAND2_X1 U81 ( .A1(A[8]), .A2(B[8]), .ZN(n61) );
  NAND2_X1 U82 ( .A1(A[8]), .A2(n52), .ZN(n62) );
  NAND2_X1 U83 ( .A1(carry[8]), .A2(B[8]), .ZN(n63) );
  NAND3_X1 U84 ( .A1(n62), .A2(n63), .A3(n61), .ZN(carry[9]) );
  XOR2_X1 U85 ( .A(A[9]), .B(B[9]), .Z(n64) );
  XOR2_X1 U86 ( .A(n64), .B(n59), .Z(SUM[9]) );
  NAND2_X1 U87 ( .A1(A[9]), .A2(B[9]), .ZN(n65) );
  NAND2_X1 U88 ( .A1(A[9]), .A2(n58), .ZN(n66) );
  NAND2_X1 U89 ( .A1(B[9]), .A2(carry[9]), .ZN(n67) );
  NAND3_X1 U90 ( .A1(n65), .A2(n66), .A3(n67), .ZN(carry[10]) );
  XOR2_X1 U91 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U92 ( .A1(B[0]), .A2(A[0]), .ZN(n69) );
endmodule


module datapath_DW_mult_tc_24 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323;

  FA_X1 U6 ( .A(n24), .B(n27), .CI(n6), .CO(n5), .S(product[10]) );
  FA_X1 U7 ( .A(n28), .B(n33), .CI(n7), .CO(n6), .S(product[9]) );
  FA_X1 U8 ( .A(n34), .B(n39), .CI(n8), .CO(n7), .S(product[8]) );
  FA_X1 U9 ( .A(n40), .B(n45), .CI(n9), .CO(n8), .S(product[7]) );
  FA_X1 U11 ( .A(n50), .B(n53), .CI(n11), .CO(n10), .S(product[5]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n266), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n265), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n269), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n268), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n271), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  NAND2_X1 U157 ( .A1(n289), .A2(n318), .ZN(n291) );
  AND2_X1 U158 ( .A1(n104), .A2(n72), .ZN(n206) );
  AND3_X1 U159 ( .A1(n252), .A2(n253), .A3(n254), .ZN(product[15]) );
  INV_X1 U160 ( .A(n237), .ZN(n208) );
  NAND2_X2 U161 ( .A1(n257), .A2(n258), .ZN(n209) );
  NAND2_X1 U162 ( .A1(n257), .A2(n258), .ZN(n289) );
  NAND3_X1 U163 ( .A1(n214), .A2(n215), .A3(n216), .ZN(n210) );
  NAND3_X1 U164 ( .A1(n214), .A2(n215), .A3(n216), .ZN(n211) );
  XOR2_X1 U165 ( .A(n95), .B(n102), .Z(n212) );
  XOR2_X1 U166 ( .A(n23), .B(n20), .Z(n213) );
  XOR2_X1 U167 ( .A(n5), .B(n213), .Z(product[11]) );
  NAND2_X1 U168 ( .A1(n5), .A2(n23), .ZN(n214) );
  NAND2_X1 U169 ( .A1(n5), .A2(n20), .ZN(n215) );
  NAND2_X1 U170 ( .A1(n23), .A2(n20), .ZN(n216) );
  NAND3_X1 U171 ( .A1(n214), .A2(n215), .A3(n216), .ZN(n4) );
  CLKBUF_X1 U172 ( .A(n10), .Z(n217) );
  NAND3_X1 U173 ( .A1(n249), .A2(n250), .A3(n251), .ZN(n218) );
  NAND3_X1 U174 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n219) );
  NAND3_X1 U175 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n220) );
  NAND3_X1 U176 ( .A1(n235), .A2(n234), .A3(n236), .ZN(n221) );
  NAND3_X1 U177 ( .A1(n234), .A2(n235), .A3(n236), .ZN(n222) );
  OAI22_X1 U178 ( .A1(n260), .A2(n275), .B1(n320), .B2(n273), .ZN(n223) );
  XNOR2_X1 U179 ( .A(n206), .B(n224), .ZN(product[2]) );
  XNOR2_X1 U180 ( .A(n103), .B(n96), .ZN(n224) );
  NAND2_X1 U181 ( .A1(n206), .A2(n103), .ZN(n225) );
  NAND2_X1 U182 ( .A1(n206), .A2(n96), .ZN(n226) );
  NAND2_X1 U183 ( .A1(n103), .A2(n96), .ZN(n227) );
  NAND3_X1 U184 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n13) );
  NAND2_X2 U185 ( .A1(n279), .A2(n317), .ZN(n281) );
  CLKBUF_X3 U186 ( .A(a[1]), .Z(n228) );
  XOR2_X1 U187 ( .A(n223), .B(n72), .Z(product[1]) );
  XNOR2_X1 U188 ( .A(a[2]), .B(a[1]), .ZN(n279) );
  XOR2_X1 U189 ( .A(n46), .B(n49), .Z(n229) );
  XOR2_X1 U190 ( .A(n217), .B(n229), .Z(product[6]) );
  NAND2_X1 U191 ( .A1(n10), .A2(n46), .ZN(n230) );
  NAND2_X1 U192 ( .A1(n10), .A2(n49), .ZN(n231) );
  NAND2_X1 U193 ( .A1(n46), .A2(n49), .ZN(n232) );
  NAND3_X1 U194 ( .A1(n230), .A2(n231), .A3(n232), .ZN(n9) );
  XOR2_X1 U195 ( .A(n18), .B(n19), .Z(n233) );
  XOR2_X1 U196 ( .A(n211), .B(n233), .Z(product[12]) );
  NAND2_X1 U197 ( .A1(n210), .A2(n18), .ZN(n234) );
  NAND2_X1 U198 ( .A1(n4), .A2(n19), .ZN(n235) );
  NAND2_X1 U199 ( .A1(n18), .A2(n19), .ZN(n236) );
  NAND3_X1 U200 ( .A1(n234), .A2(n235), .A3(n236), .ZN(n3) );
  INV_X1 U201 ( .A(n261), .ZN(n237) );
  NAND3_X1 U202 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n238) );
  INV_X1 U203 ( .A(n261), .ZN(n260) );
  XNOR2_X1 U204 ( .A(n239), .B(n220), .ZN(product[3]) );
  XNOR2_X1 U205 ( .A(n212), .B(n71), .ZN(n239) );
  NAND2_X1 U206 ( .A1(n56), .A2(n71), .ZN(n240) );
  NAND2_X1 U207 ( .A1(n13), .A2(n212), .ZN(n241) );
  NAND2_X1 U208 ( .A1(n71), .A2(n219), .ZN(n242) );
  NAND3_X1 U209 ( .A1(n242), .A2(n241), .A3(n240), .ZN(n12) );
  XOR2_X1 U210 ( .A(n54), .B(n55), .Z(n243) );
  XOR2_X1 U211 ( .A(n243), .B(n238), .Z(product[4]) );
  NAND2_X1 U212 ( .A1(n54), .A2(n55), .ZN(n244) );
  NAND2_X1 U213 ( .A1(n54), .A2(n12), .ZN(n245) );
  NAND2_X1 U214 ( .A1(n12), .A2(n55), .ZN(n246) );
  NAND3_X1 U215 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n11) );
  XNOR2_X1 U216 ( .A(n247), .B(n218), .ZN(product[14]) );
  XNOR2_X1 U217 ( .A(n263), .B(n15), .ZN(n247) );
  XNOR2_X1 U218 ( .A(n248), .B(n222), .ZN(product[13]) );
  XNOR2_X1 U219 ( .A(n17), .B(n262), .ZN(n248) );
  NAND2_X1 U220 ( .A1(n17), .A2(n262), .ZN(n249) );
  NAND2_X1 U221 ( .A1(n17), .A2(n221), .ZN(n250) );
  NAND2_X1 U222 ( .A1(n262), .A2(n3), .ZN(n251) );
  NAND3_X1 U223 ( .A1(n249), .A2(n250), .A3(n251), .ZN(n2) );
  NAND2_X1 U224 ( .A1(n263), .A2(n15), .ZN(n252) );
  NAND2_X1 U225 ( .A1(n263), .A2(n2), .ZN(n253) );
  NAND2_X1 U226 ( .A1(n15), .A2(n2), .ZN(n254) );
  NAND2_X1 U227 ( .A1(a[4]), .A2(a[3]), .ZN(n257) );
  NAND2_X1 U228 ( .A1(n255), .A2(n256), .ZN(n258) );
  INV_X1 U229 ( .A(a[4]), .ZN(n255) );
  INV_X1 U230 ( .A(a[3]), .ZN(n256) );
  BUF_X1 U231 ( .A(n279), .Z(n259) );
  INV_X1 U232 ( .A(n15), .ZN(n262) );
  INV_X1 U233 ( .A(n21), .ZN(n265) );
  INV_X1 U234 ( .A(n298), .ZN(n266) );
  INV_X1 U235 ( .A(n309), .ZN(n263) );
  INV_X1 U236 ( .A(b[0]), .ZN(n261) );
  INV_X1 U237 ( .A(n278), .ZN(n271) );
  INV_X1 U238 ( .A(n287), .ZN(n269) );
  INV_X1 U239 ( .A(n31), .ZN(n268) );
  XOR2_X1 U240 ( .A(a[6]), .B(n267), .Z(n300) );
  INV_X1 U241 ( .A(a[0]), .ZN(n273) );
  INV_X1 U242 ( .A(a[5]), .ZN(n267) );
  INV_X1 U243 ( .A(a[7]), .ZN(n264) );
  INV_X1 U244 ( .A(a[3]), .ZN(n270) );
  INV_X1 U245 ( .A(a[1]), .ZN(n272) );
  NOR2_X1 U246 ( .A1(n273), .A2(n208), .ZN(product[0]) );
  OAI22_X1 U247 ( .A1(n274), .A2(n275), .B1(n276), .B2(n273), .ZN(n99) );
  OAI22_X1 U248 ( .A1(n276), .A2(n275), .B1(n277), .B2(n273), .ZN(n98) );
  XNOR2_X1 U249 ( .A(b[6]), .B(n228), .ZN(n276) );
  OAI22_X1 U250 ( .A1(n273), .A2(n277), .B1(n275), .B2(n277), .ZN(n278) );
  XNOR2_X1 U251 ( .A(b[7]), .B(n228), .ZN(n277) );
  NOR2_X1 U252 ( .A1(n279), .A2(n261), .ZN(n96) );
  OAI22_X1 U253 ( .A1(n280), .A2(n281), .B1(n279), .B2(n282), .ZN(n95) );
  XNOR2_X1 U254 ( .A(a[3]), .B(n260), .ZN(n280) );
  OAI22_X1 U255 ( .A1(n282), .A2(n281), .B1(n259), .B2(n283), .ZN(n94) );
  XNOR2_X1 U256 ( .A(b[1]), .B(a[3]), .ZN(n282) );
  OAI22_X1 U257 ( .A1(n283), .A2(n281), .B1(n259), .B2(n284), .ZN(n93) );
  XNOR2_X1 U258 ( .A(b[2]), .B(a[3]), .ZN(n283) );
  OAI22_X1 U259 ( .A1(n284), .A2(n281), .B1(n259), .B2(n285), .ZN(n92) );
  XNOR2_X1 U260 ( .A(b[3]), .B(a[3]), .ZN(n284) );
  OAI22_X1 U261 ( .A1(n285), .A2(n281), .B1(n259), .B2(n286), .ZN(n91) );
  XNOR2_X1 U262 ( .A(b[4]), .B(a[3]), .ZN(n285) );
  OAI22_X1 U263 ( .A1(n288), .A2(n259), .B1(n281), .B2(n288), .ZN(n287) );
  NOR2_X1 U264 ( .A1(n209), .A2(n208), .ZN(n88) );
  OAI22_X1 U265 ( .A1(n290), .A2(n291), .B1(n209), .B2(n292), .ZN(n87) );
  XNOR2_X1 U266 ( .A(a[5]), .B(n237), .ZN(n290) );
  OAI22_X1 U267 ( .A1(n292), .A2(n291), .B1(n209), .B2(n293), .ZN(n86) );
  XNOR2_X1 U268 ( .A(b[1]), .B(a[5]), .ZN(n292) );
  OAI22_X1 U269 ( .A1(n293), .A2(n291), .B1(n209), .B2(n294), .ZN(n85) );
  XNOR2_X1 U270 ( .A(b[2]), .B(a[5]), .ZN(n293) );
  OAI22_X1 U271 ( .A1(n294), .A2(n291), .B1(n209), .B2(n295), .ZN(n84) );
  XNOR2_X1 U272 ( .A(b[3]), .B(a[5]), .ZN(n294) );
  OAI22_X1 U273 ( .A1(n295), .A2(n291), .B1(n209), .B2(n296), .ZN(n83) );
  XNOR2_X1 U274 ( .A(b[4]), .B(a[5]), .ZN(n295) );
  OAI22_X1 U275 ( .A1(n296), .A2(n291), .B1(n209), .B2(n297), .ZN(n82) );
  XNOR2_X1 U276 ( .A(b[5]), .B(a[5]), .ZN(n296) );
  OAI22_X1 U277 ( .A1(n299), .A2(n209), .B1(n291), .B2(n299), .ZN(n298) );
  NOR2_X1 U278 ( .A1(n300), .A2(n208), .ZN(n80) );
  OAI22_X1 U279 ( .A1(n301), .A2(n302), .B1(n300), .B2(n303), .ZN(n79) );
  XNOR2_X1 U280 ( .A(a[7]), .B(n237), .ZN(n301) );
  OAI22_X1 U281 ( .A1(n304), .A2(n302), .B1(n300), .B2(n305), .ZN(n77) );
  OAI22_X1 U282 ( .A1(n305), .A2(n302), .B1(n300), .B2(n306), .ZN(n76) );
  XNOR2_X1 U283 ( .A(b[3]), .B(a[7]), .ZN(n305) );
  OAI22_X1 U284 ( .A1(n306), .A2(n302), .B1(n300), .B2(n307), .ZN(n75) );
  XNOR2_X1 U285 ( .A(b[4]), .B(a[7]), .ZN(n306) );
  OAI22_X1 U286 ( .A1(n307), .A2(n302), .B1(n300), .B2(n308), .ZN(n74) );
  XNOR2_X1 U287 ( .A(b[5]), .B(a[7]), .ZN(n307) );
  OAI22_X1 U288 ( .A1(n310), .A2(n300), .B1(n302), .B2(n310), .ZN(n309) );
  OAI21_X1 U289 ( .B1(n260), .B2(n272), .A(n275), .ZN(n72) );
  OAI21_X1 U290 ( .B1(n270), .B2(n281), .A(n311), .ZN(n71) );
  OR3_X1 U291 ( .A1(n259), .A2(n237), .A3(n270), .ZN(n311) );
  OAI21_X1 U292 ( .B1(n267), .B2(n291), .A(n312), .ZN(n70) );
  OR3_X1 U293 ( .A1(n289), .A2(n237), .A3(n267), .ZN(n312) );
  OAI21_X1 U294 ( .B1(n264), .B2(n302), .A(n313), .ZN(n69) );
  OR3_X1 U295 ( .A1(n300), .A2(n237), .A3(n264), .ZN(n313) );
  XNOR2_X1 U296 ( .A(n314), .B(n315), .ZN(n38) );
  OR2_X1 U297 ( .A1(n314), .A2(n315), .ZN(n37) );
  OAI22_X1 U298 ( .A1(n286), .A2(n281), .B1(n259), .B2(n316), .ZN(n315) );
  XNOR2_X1 U299 ( .A(b[5]), .B(a[3]), .ZN(n286) );
  OAI22_X1 U300 ( .A1(n303), .A2(n302), .B1(n300), .B2(n304), .ZN(n314) );
  XNOR2_X1 U301 ( .A(b[2]), .B(a[7]), .ZN(n304) );
  XNOR2_X1 U302 ( .A(b[1]), .B(a[7]), .ZN(n303) );
  OAI22_X1 U303 ( .A1(n316), .A2(n281), .B1(n259), .B2(n288), .ZN(n31) );
  XNOR2_X1 U304 ( .A(b[7]), .B(a[3]), .ZN(n288) );
  XNOR2_X1 U305 ( .A(n270), .B(a[2]), .ZN(n317) );
  XNOR2_X1 U306 ( .A(b[6]), .B(a[3]), .ZN(n316) );
  OAI22_X1 U307 ( .A1(n297), .A2(n291), .B1(n209), .B2(n299), .ZN(n21) );
  XNOR2_X1 U308 ( .A(b[7]), .B(a[5]), .ZN(n299) );
  XNOR2_X1 U309 ( .A(n267), .B(a[4]), .ZN(n318) );
  XNOR2_X1 U310 ( .A(b[6]), .B(a[5]), .ZN(n297) );
  OAI22_X1 U311 ( .A1(n308), .A2(n302), .B1(n300), .B2(n310), .ZN(n15) );
  XNOR2_X1 U312 ( .A(b[7]), .B(a[7]), .ZN(n310) );
  NAND2_X1 U313 ( .A1(n300), .A2(n319), .ZN(n302) );
  XNOR2_X1 U314 ( .A(n264), .B(a[6]), .ZN(n319) );
  XNOR2_X1 U315 ( .A(b[6]), .B(a[7]), .ZN(n308) );
  OAI22_X1 U316 ( .A1(n260), .A2(n275), .B1(n320), .B2(n273), .ZN(n104) );
  OAI22_X1 U317 ( .A1(n275), .A2(n320), .B1(n321), .B2(n273), .ZN(n103) );
  XNOR2_X1 U318 ( .A(b[1]), .B(n228), .ZN(n320) );
  OAI22_X1 U319 ( .A1(n321), .A2(n275), .B1(n322), .B2(n273), .ZN(n102) );
  XNOR2_X1 U320 ( .A(b[2]), .B(n228), .ZN(n321) );
  OAI22_X1 U321 ( .A1(n322), .A2(n275), .B1(n323), .B2(n273), .ZN(n101) );
  XNOR2_X1 U322 ( .A(b[3]), .B(n228), .ZN(n322) );
  OAI22_X1 U323 ( .A1(n323), .A2(n275), .B1(n274), .B2(n273), .ZN(n100) );
  XNOR2_X1 U324 ( .A(b[5]), .B(n228), .ZN(n274) );
  NAND2_X1 U325 ( .A1(a[1]), .A2(n273), .ZN(n275) );
  XNOR2_X1 U326 ( .A(b[4]), .B(n228), .ZN(n323) );
endmodule


module datapath_DW01_add_24 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n62;
  wire   [15:1] carry;

  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n62), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(n7), .Z(n1) );
  CLKBUF_X1 U2 ( .A(n8), .Z(n2) );
  NAND3_X1 U3 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n3) );
  NAND3_X1 U4 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n4) );
  NAND3_X1 U5 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n5) );
  NAND3_X1 U6 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n6) );
  NAND3_X1 U7 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n7) );
  NAND3_X1 U8 ( .A1(n23), .A2(n24), .A3(n25), .ZN(n8) );
  CLKBUF_X1 U9 ( .A(carry[12]), .Z(n9) );
  NAND3_X1 U10 ( .A1(n19), .A2(n20), .A3(n21), .ZN(n10) );
  CLKBUF_X1 U11 ( .A(n3), .Z(n11) );
  NAND3_X1 U12 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n12) );
  XOR2_X1 U13 ( .A(B[8]), .B(A[8]), .Z(n13) );
  XOR2_X1 U14 ( .A(n11), .B(n13), .Z(SUM[8]) );
  NAND2_X1 U15 ( .A1(n3), .A2(B[8]), .ZN(n14) );
  NAND2_X1 U16 ( .A1(carry[8]), .A2(A[8]), .ZN(n15) );
  NAND2_X1 U17 ( .A1(B[8]), .A2(A[8]), .ZN(n16) );
  NAND3_X1 U18 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[9]) );
  NAND3_X1 U19 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n17) );
  XNOR2_X1 U20 ( .A(B[14]), .B(A[14]), .ZN(n26) );
  XOR2_X1 U21 ( .A(B[13]), .B(A[13]), .Z(n18) );
  XOR2_X1 U22 ( .A(n1), .B(n18), .Z(SUM[13]) );
  NAND2_X1 U23 ( .A1(n7), .A2(B[13]), .ZN(n19) );
  NAND2_X1 U24 ( .A1(carry[13]), .A2(A[13]), .ZN(n20) );
  NAND2_X1 U25 ( .A1(B[13]), .A2(A[13]), .ZN(n21) );
  NAND3_X1 U26 ( .A1(n20), .A2(n19), .A3(n21), .ZN(carry[14]) );
  XOR2_X1 U27 ( .A(B[9]), .B(A[9]), .Z(n22) );
  XOR2_X1 U28 ( .A(carry[9]), .B(n22), .Z(SUM[9]) );
  NAND2_X1 U29 ( .A1(n12), .A2(B[9]), .ZN(n23) );
  NAND2_X1 U30 ( .A1(carry[9]), .A2(A[9]), .ZN(n24) );
  NAND2_X1 U31 ( .A1(B[9]), .A2(A[9]), .ZN(n25) );
  NAND3_X1 U32 ( .A1(n23), .A2(n24), .A3(n25), .ZN(carry[10]) );
  CLKBUF_X1 U33 ( .A(n10), .Z(n36) );
  XNOR2_X1 U34 ( .A(n26), .B(n36), .ZN(SUM[14]) );
  XOR2_X1 U35 ( .A(B[7]), .B(A[7]), .Z(n27) );
  XOR2_X1 U36 ( .A(carry[7]), .B(n27), .Z(SUM[7]) );
  NAND2_X1 U37 ( .A1(carry[7]), .A2(B[7]), .ZN(n28) );
  NAND2_X1 U38 ( .A1(carry[7]), .A2(A[7]), .ZN(n29) );
  NAND2_X1 U39 ( .A1(B[7]), .A2(A[7]), .ZN(n30) );
  NAND3_X1 U40 ( .A1(n28), .A2(n29), .A3(n30), .ZN(carry[8]) );
  CLKBUF_X1 U41 ( .A(B[4]), .Z(n31) );
  XOR2_X1 U42 ( .A(B[10]), .B(A[10]), .Z(n32) );
  XOR2_X1 U43 ( .A(n2), .B(n32), .Z(SUM[10]) );
  NAND2_X1 U44 ( .A1(n8), .A2(B[10]), .ZN(n33) );
  NAND2_X1 U45 ( .A1(carry[10]), .A2(A[10]), .ZN(n34) );
  NAND2_X1 U46 ( .A1(B[10]), .A2(A[10]), .ZN(n35) );
  NAND3_X1 U47 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[11]) );
  XNOR2_X1 U48 ( .A(n37), .B(carry[15]), .ZN(SUM[15]) );
  XNOR2_X1 U49 ( .A(B[15]), .B(A[15]), .ZN(n37) );
  XOR2_X1 U50 ( .A(B[11]), .B(A[11]), .Z(n38) );
  XOR2_X1 U51 ( .A(carry[11]), .B(n38), .Z(SUM[11]) );
  NAND2_X1 U52 ( .A1(n17), .A2(B[11]), .ZN(n39) );
  NAND2_X1 U53 ( .A1(n17), .A2(A[11]), .ZN(n40) );
  NAND2_X1 U54 ( .A1(B[11]), .A2(A[11]), .ZN(n41) );
  NAND3_X1 U55 ( .A1(n39), .A2(n40), .A3(n41), .ZN(carry[12]) );
  XOR2_X1 U56 ( .A(B[12]), .B(A[12]), .Z(n42) );
  XOR2_X1 U57 ( .A(n9), .B(n42), .Z(SUM[12]) );
  NAND2_X1 U58 ( .A1(B[12]), .A2(n4), .ZN(n43) );
  NAND2_X1 U59 ( .A1(carry[12]), .A2(A[12]), .ZN(n44) );
  NAND2_X1 U60 ( .A1(B[12]), .A2(A[12]), .ZN(n45) );
  NAND3_X1 U61 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[13]) );
  XOR2_X1 U62 ( .A(A[3]), .B(B[3]), .Z(n46) );
  XOR2_X1 U63 ( .A(n46), .B(n6), .Z(SUM[3]) );
  NAND2_X1 U64 ( .A1(A[3]), .A2(B[3]), .ZN(n47) );
  NAND2_X1 U65 ( .A1(A[3]), .A2(n5), .ZN(n48) );
  NAND2_X1 U66 ( .A1(B[3]), .A2(carry[3]), .ZN(n49) );
  NAND3_X1 U67 ( .A1(n47), .A2(n48), .A3(n49), .ZN(carry[4]) );
  XOR2_X1 U68 ( .A(A[4]), .B(n31), .Z(n50) );
  XOR2_X1 U69 ( .A(n50), .B(carry[4]), .Z(SUM[4]) );
  NAND2_X1 U70 ( .A1(A[4]), .A2(B[4]), .ZN(n51) );
  NAND2_X1 U71 ( .A1(A[4]), .A2(carry[4]), .ZN(n52) );
  NAND2_X1 U72 ( .A1(B[4]), .A2(carry[4]), .ZN(n53) );
  NAND3_X1 U73 ( .A1(n51), .A2(n52), .A3(n53), .ZN(carry[5]) );
  XOR2_X1 U74 ( .A(carry[2]), .B(A[2]), .Z(n54) );
  XOR2_X1 U75 ( .A(B[2]), .B(n54), .Z(SUM[2]) );
  NAND2_X1 U76 ( .A1(B[2]), .A2(carry[2]), .ZN(n55) );
  NAND2_X1 U77 ( .A1(B[2]), .A2(A[2]), .ZN(n56) );
  NAND2_X1 U78 ( .A1(carry[2]), .A2(A[2]), .ZN(n57) );
  NAND3_X1 U79 ( .A1(n55), .A2(n56), .A3(n57), .ZN(carry[3]) );
  NAND2_X1 U80 ( .A1(carry[14]), .A2(B[14]), .ZN(n58) );
  NAND2_X1 U81 ( .A1(n10), .A2(A[14]), .ZN(n59) );
  NAND2_X1 U82 ( .A1(B[14]), .A2(A[14]), .ZN(n60) );
  NAND3_X1 U83 ( .A1(n59), .A2(n58), .A3(n60), .ZN(carry[15]) );
  XOR2_X1 U84 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U85 ( .A1(B[0]), .A2(A[0]), .ZN(n62) );
endmodule


module datapath_DW_mult_tc_23 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74,
         n75, n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92,
         n93, n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342;

  FA_X1 U4 ( .A(n19), .B(n18), .CI(n4), .CO(n3), .S(product[12]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n285), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n284), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n288), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n287), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n290), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n94), .B(n88), .CI(n101), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  NAND2_X1 U157 ( .A1(n308), .A2(n337), .ZN(n310) );
  INV_X1 U158 ( .A(n15), .ZN(n281) );
  INV_X1 U159 ( .A(a[0]), .ZN(n292) );
  XNOR2_X1 U160 ( .A(n282), .B(n15), .ZN(n206) );
  AND3_X1 U161 ( .A1(n260), .A2(n261), .A3(n262), .ZN(product[15]) );
  XNOR2_X1 U162 ( .A(n224), .B(n208), .ZN(product[5]) );
  XNOR2_X1 U163 ( .A(n50), .B(n53), .ZN(n208) );
  XOR2_X1 U164 ( .A(n23), .B(n20), .Z(n209) );
  XOR2_X1 U165 ( .A(n5), .B(n209), .Z(product[11]) );
  NAND2_X1 U166 ( .A1(n5), .A2(n23), .ZN(n210) );
  NAND2_X1 U167 ( .A1(n5), .A2(n20), .ZN(n211) );
  NAND2_X1 U168 ( .A1(n23), .A2(n20), .ZN(n212) );
  NAND3_X1 U169 ( .A1(n210), .A2(n211), .A3(n212), .ZN(n4) );
  XOR2_X1 U170 ( .A(n54), .B(n55), .Z(n213) );
  XOR2_X1 U171 ( .A(n12), .B(n213), .Z(product[4]) );
  NAND2_X1 U172 ( .A1(n12), .A2(n54), .ZN(n214) );
  NAND2_X1 U173 ( .A1(n12), .A2(n55), .ZN(n215) );
  NAND2_X1 U174 ( .A1(n54), .A2(n55), .ZN(n216) );
  NAND3_X1 U175 ( .A1(n214), .A2(n215), .A3(n216), .ZN(n11) );
  CLKBUF_X1 U176 ( .A(b[1]), .Z(n217) );
  NAND3_X1 U177 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n218) );
  CLKBUF_X1 U178 ( .A(n267), .Z(n219) );
  NAND3_X1 U179 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n220) );
  CLKBUF_X1 U180 ( .A(n225), .Z(n221) );
  CLKBUF_X1 U181 ( .A(n272), .Z(n222) );
  BUF_X2 U182 ( .A(n308), .Z(n223) );
  XNOR2_X1 U183 ( .A(a[4]), .B(a[3]), .ZN(n308) );
  CLKBUF_X1 U184 ( .A(n11), .Z(n224) );
  NAND3_X1 U185 ( .A1(n227), .A2(n226), .A3(n228), .ZN(n225) );
  NAND2_X1 U186 ( .A1(n11), .A2(n50), .ZN(n226) );
  NAND2_X1 U187 ( .A1(n11), .A2(n53), .ZN(n227) );
  NAND2_X1 U188 ( .A1(n50), .A2(n53), .ZN(n228) );
  NAND3_X1 U189 ( .A1(n226), .A2(n227), .A3(n228), .ZN(n10) );
  XNOR2_X1 U190 ( .A(n2), .B(n206), .ZN(product[14]) );
  XNOR2_X1 U191 ( .A(n229), .B(n242), .ZN(product[3]) );
  XNOR2_X1 U192 ( .A(n56), .B(n71), .ZN(n229) );
  AND2_X1 U193 ( .A1(n104), .A2(n72), .ZN(n230) );
  NAND3_X1 U194 ( .A1(n272), .A2(n271), .A3(n270), .ZN(n231) );
  NAND3_X1 U195 ( .A1(n270), .A2(n271), .A3(n222), .ZN(n232) );
  NAND3_X1 U196 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n233) );
  XOR2_X1 U197 ( .A(n28), .B(n33), .Z(n234) );
  XOR2_X1 U198 ( .A(n234), .B(n232), .Z(product[9]) );
  NAND2_X1 U199 ( .A1(n28), .A2(n33), .ZN(n235) );
  NAND2_X1 U200 ( .A1(n28), .A2(n231), .ZN(n236) );
  NAND2_X1 U201 ( .A1(n33), .A2(n7), .ZN(n237) );
  NAND3_X1 U202 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n6) );
  XOR2_X1 U203 ( .A(n24), .B(n27), .Z(n238) );
  XOR2_X1 U204 ( .A(n238), .B(n220), .Z(product[10]) );
  NAND2_X1 U205 ( .A1(n24), .A2(n27), .ZN(n239) );
  NAND2_X1 U206 ( .A1(n24), .A2(n233), .ZN(n240) );
  NAND2_X1 U207 ( .A1(n27), .A2(n6), .ZN(n241) );
  NAND3_X1 U208 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n5) );
  NAND3_X1 U209 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n242) );
  NAND3_X1 U210 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n243) );
  NAND3_X1 U211 ( .A1(n219), .A2(n266), .A3(n268), .ZN(n244) );
  XOR2_X1 U212 ( .A(n46), .B(n49), .Z(n245) );
  XOR2_X1 U213 ( .A(n221), .B(n245), .Z(product[6]) );
  NAND2_X1 U214 ( .A1(n225), .A2(n46), .ZN(n246) );
  NAND2_X1 U215 ( .A1(n10), .A2(n49), .ZN(n247) );
  NAND2_X1 U216 ( .A1(n46), .A2(n49), .ZN(n248) );
  NAND3_X1 U217 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n9) );
  XOR2_X1 U218 ( .A(n17), .B(n281), .Z(n249) );
  XOR2_X1 U219 ( .A(n3), .B(n249), .Z(product[13]) );
  NAND2_X1 U220 ( .A1(n3), .A2(n17), .ZN(n250) );
  NAND2_X1 U221 ( .A1(n3), .A2(n281), .ZN(n251) );
  NAND2_X1 U222 ( .A1(n17), .A2(n281), .ZN(n252) );
  NAND3_X1 U223 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n2) );
  NAND3_X1 U224 ( .A1(n268), .A2(n267), .A3(n266), .ZN(n253) );
  INV_X2 U225 ( .A(n280), .ZN(n279) );
  XNOR2_X1 U226 ( .A(n254), .B(n230), .ZN(product[2]) );
  XNOR2_X1 U227 ( .A(n103), .B(n96), .ZN(n254) );
  XOR2_X1 U228 ( .A(n95), .B(n102), .Z(n255) );
  NAND2_X1 U229 ( .A1(a[2]), .A2(a[1]), .ZN(n258) );
  NAND2_X1 U230 ( .A1(n256), .A2(n257), .ZN(n259) );
  NAND2_X2 U231 ( .A1(n258), .A2(n259), .ZN(n298) );
  INV_X1 U232 ( .A(a[2]), .ZN(n256) );
  INV_X1 U233 ( .A(a[1]), .ZN(n257) );
  NAND2_X1 U234 ( .A1(n2), .A2(n282), .ZN(n260) );
  NAND2_X1 U235 ( .A1(n2), .A2(n15), .ZN(n261) );
  NAND2_X1 U236 ( .A1(n282), .A2(n15), .ZN(n262) );
  CLKBUF_X1 U237 ( .A(b[1]), .Z(n263) );
  CLKBUF_X1 U238 ( .A(b[2]), .Z(n264) );
  XOR2_X1 U239 ( .A(n40), .B(n45), .Z(n265) );
  XOR2_X1 U240 ( .A(n265), .B(n218), .Z(product[7]) );
  NAND2_X1 U241 ( .A1(n40), .A2(n45), .ZN(n266) );
  NAND2_X1 U242 ( .A1(n40), .A2(n243), .ZN(n267) );
  NAND2_X1 U243 ( .A1(n45), .A2(n9), .ZN(n268) );
  NAND3_X1 U244 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n8) );
  XOR2_X1 U245 ( .A(n34), .B(n39), .Z(n269) );
  XOR2_X1 U246 ( .A(n269), .B(n244), .Z(product[8]) );
  NAND2_X1 U247 ( .A1(n34), .A2(n39), .ZN(n270) );
  NAND2_X1 U248 ( .A1(n34), .A2(n253), .ZN(n271) );
  NAND2_X1 U249 ( .A1(n39), .A2(n8), .ZN(n272) );
  NAND3_X1 U250 ( .A1(n270), .A2(n271), .A3(n272), .ZN(n7) );
  NAND2_X1 U251 ( .A1(n103), .A2(n96), .ZN(n273) );
  NAND2_X1 U252 ( .A1(n230), .A2(n103), .ZN(n274) );
  NAND2_X1 U253 ( .A1(n96), .A2(n14), .ZN(n275) );
  NAND3_X1 U254 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n13) );
  NAND2_X1 U255 ( .A1(n255), .A2(n71), .ZN(n276) );
  NAND2_X1 U256 ( .A1(n255), .A2(n242), .ZN(n277) );
  NAND2_X1 U257 ( .A1(n71), .A2(n13), .ZN(n278) );
  NAND3_X1 U258 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n12) );
  INV_X1 U259 ( .A(n21), .ZN(n284) );
  INV_X1 U260 ( .A(n317), .ZN(n285) );
  INV_X1 U261 ( .A(n328), .ZN(n282) );
  INV_X1 U262 ( .A(n297), .ZN(n290) );
  INV_X1 U263 ( .A(n306), .ZN(n288) );
  INV_X1 U264 ( .A(n31), .ZN(n287) );
  INV_X1 U265 ( .A(b[0]), .ZN(n280) );
  INV_X1 U266 ( .A(a[5]), .ZN(n286) );
  INV_X1 U267 ( .A(a[7]), .ZN(n283) );
  INV_X1 U268 ( .A(a[3]), .ZN(n289) );
  NAND2_X2 U269 ( .A1(n298), .A2(n336), .ZN(n300) );
  INV_X1 U270 ( .A(a[1]), .ZN(n291) );
  XOR2_X2 U271 ( .A(a[6]), .B(n286), .Z(n319) );
  NOR2_X1 U272 ( .A1(n292), .A2(n280), .ZN(product[0]) );
  OAI22_X1 U273 ( .A1(n293), .A2(n294), .B1(n295), .B2(n292), .ZN(n99) );
  OAI22_X1 U274 ( .A1(n295), .A2(n294), .B1(n296), .B2(n292), .ZN(n98) );
  XNOR2_X1 U275 ( .A(b[6]), .B(a[1]), .ZN(n295) );
  OAI22_X1 U276 ( .A1(n292), .A2(n296), .B1(n294), .B2(n296), .ZN(n297) );
  XNOR2_X1 U277 ( .A(b[7]), .B(a[1]), .ZN(n296) );
  NOR2_X1 U278 ( .A1(n298), .A2(n280), .ZN(n96) );
  OAI22_X1 U279 ( .A1(n299), .A2(n300), .B1(n298), .B2(n301), .ZN(n95) );
  XNOR2_X1 U280 ( .A(a[3]), .B(n279), .ZN(n299) );
  OAI22_X1 U281 ( .A1(n301), .A2(n300), .B1(n298), .B2(n302), .ZN(n94) );
  XNOR2_X1 U282 ( .A(n217), .B(a[3]), .ZN(n301) );
  OAI22_X1 U283 ( .A1(n302), .A2(n300), .B1(n298), .B2(n303), .ZN(n93) );
  XNOR2_X1 U284 ( .A(b[2]), .B(a[3]), .ZN(n302) );
  OAI22_X1 U285 ( .A1(n303), .A2(n300), .B1(n298), .B2(n304), .ZN(n92) );
  XNOR2_X1 U286 ( .A(b[3]), .B(a[3]), .ZN(n303) );
  OAI22_X1 U287 ( .A1(n304), .A2(n300), .B1(n298), .B2(n305), .ZN(n91) );
  XNOR2_X1 U288 ( .A(b[4]), .B(a[3]), .ZN(n304) );
  OAI22_X1 U289 ( .A1(n307), .A2(n298), .B1(n300), .B2(n307), .ZN(n306) );
  NOR2_X1 U290 ( .A1(n223), .A2(n280), .ZN(n88) );
  OAI22_X1 U291 ( .A1(n309), .A2(n310), .B1(n223), .B2(n311), .ZN(n87) );
  XNOR2_X1 U292 ( .A(a[5]), .B(n279), .ZN(n309) );
  OAI22_X1 U293 ( .A1(n311), .A2(n310), .B1(n223), .B2(n312), .ZN(n86) );
  XNOR2_X1 U294 ( .A(n263), .B(a[5]), .ZN(n311) );
  OAI22_X1 U295 ( .A1(n312), .A2(n310), .B1(n223), .B2(n313), .ZN(n85) );
  XNOR2_X1 U296 ( .A(n264), .B(a[5]), .ZN(n312) );
  OAI22_X1 U297 ( .A1(n313), .A2(n310), .B1(n223), .B2(n314), .ZN(n84) );
  XNOR2_X1 U298 ( .A(b[3]), .B(a[5]), .ZN(n313) );
  OAI22_X1 U299 ( .A1(n314), .A2(n310), .B1(n223), .B2(n315), .ZN(n83) );
  XNOR2_X1 U300 ( .A(b[4]), .B(a[5]), .ZN(n314) );
  OAI22_X1 U301 ( .A1(n315), .A2(n310), .B1(n223), .B2(n316), .ZN(n82) );
  XNOR2_X1 U302 ( .A(b[5]), .B(a[5]), .ZN(n315) );
  OAI22_X1 U303 ( .A1(n318), .A2(n223), .B1(n310), .B2(n318), .ZN(n317) );
  NOR2_X1 U304 ( .A1(n319), .A2(n280), .ZN(n80) );
  OAI22_X1 U305 ( .A1(n320), .A2(n321), .B1(n319), .B2(n322), .ZN(n79) );
  XNOR2_X1 U306 ( .A(a[7]), .B(n279), .ZN(n320) );
  OAI22_X1 U307 ( .A1(n323), .A2(n321), .B1(n319), .B2(n324), .ZN(n77) );
  OAI22_X1 U308 ( .A1(n324), .A2(n321), .B1(n319), .B2(n325), .ZN(n76) );
  XNOR2_X1 U309 ( .A(b[3]), .B(a[7]), .ZN(n324) );
  OAI22_X1 U310 ( .A1(n325), .A2(n321), .B1(n319), .B2(n326), .ZN(n75) );
  XNOR2_X1 U311 ( .A(b[4]), .B(a[7]), .ZN(n325) );
  OAI22_X1 U312 ( .A1(n326), .A2(n321), .B1(n319), .B2(n327), .ZN(n74) );
  XNOR2_X1 U313 ( .A(b[5]), .B(a[7]), .ZN(n326) );
  OAI22_X1 U314 ( .A1(n329), .A2(n319), .B1(n321), .B2(n329), .ZN(n328) );
  OAI21_X1 U315 ( .B1(n279), .B2(n291), .A(n294), .ZN(n72) );
  OAI21_X1 U316 ( .B1(n289), .B2(n300), .A(n330), .ZN(n71) );
  OR3_X1 U317 ( .A1(n298), .A2(n279), .A3(n289), .ZN(n330) );
  OAI21_X1 U318 ( .B1(n286), .B2(n310), .A(n331), .ZN(n70) );
  OR3_X1 U319 ( .A1(n223), .A2(n279), .A3(n286), .ZN(n331) );
  OAI21_X1 U320 ( .B1(n283), .B2(n321), .A(n332), .ZN(n69) );
  OR3_X1 U321 ( .A1(n319), .A2(n279), .A3(n283), .ZN(n332) );
  XNOR2_X1 U322 ( .A(n333), .B(n334), .ZN(n38) );
  OR2_X1 U323 ( .A1(n333), .A2(n334), .ZN(n37) );
  OAI22_X1 U324 ( .A1(n305), .A2(n300), .B1(n298), .B2(n335), .ZN(n334) );
  XNOR2_X1 U325 ( .A(b[5]), .B(a[3]), .ZN(n305) );
  OAI22_X1 U326 ( .A1(n322), .A2(n321), .B1(n319), .B2(n323), .ZN(n333) );
  XNOR2_X1 U327 ( .A(n264), .B(a[7]), .ZN(n323) );
  XNOR2_X1 U328 ( .A(n263), .B(a[7]), .ZN(n322) );
  OAI22_X1 U329 ( .A1(n335), .A2(n300), .B1(n298), .B2(n307), .ZN(n31) );
  XNOR2_X1 U330 ( .A(b[7]), .B(a[3]), .ZN(n307) );
  XNOR2_X1 U331 ( .A(n289), .B(a[2]), .ZN(n336) );
  XNOR2_X1 U332 ( .A(b[6]), .B(a[3]), .ZN(n335) );
  OAI22_X1 U333 ( .A1(n316), .A2(n310), .B1(n223), .B2(n318), .ZN(n21) );
  XNOR2_X1 U334 ( .A(b[7]), .B(a[5]), .ZN(n318) );
  XNOR2_X1 U335 ( .A(n286), .B(a[4]), .ZN(n337) );
  XNOR2_X1 U336 ( .A(b[6]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U337 ( .A1(n327), .A2(n321), .B1(n319), .B2(n329), .ZN(n15) );
  XNOR2_X1 U338 ( .A(b[7]), .B(a[7]), .ZN(n329) );
  NAND2_X1 U339 ( .A1(n319), .A2(n338), .ZN(n321) );
  XNOR2_X1 U340 ( .A(n283), .B(a[6]), .ZN(n338) );
  XNOR2_X1 U341 ( .A(b[6]), .B(a[7]), .ZN(n327) );
  OAI22_X1 U342 ( .A1(n279), .A2(n294), .B1(n339), .B2(n292), .ZN(n104) );
  OAI22_X1 U343 ( .A1(n339), .A2(n294), .B1(n340), .B2(n292), .ZN(n103) );
  XNOR2_X1 U344 ( .A(b[1]), .B(a[1]), .ZN(n339) );
  OAI22_X1 U345 ( .A1(n340), .A2(n294), .B1(n341), .B2(n292), .ZN(n102) );
  XNOR2_X1 U346 ( .A(b[2]), .B(a[1]), .ZN(n340) );
  OAI22_X1 U347 ( .A1(n341), .A2(n294), .B1(n342), .B2(n292), .ZN(n101) );
  XNOR2_X1 U348 ( .A(b[3]), .B(a[1]), .ZN(n341) );
  OAI22_X1 U349 ( .A1(n342), .A2(n294), .B1(n293), .B2(n292), .ZN(n100) );
  XNOR2_X1 U350 ( .A(b[5]), .B(a[1]), .ZN(n293) );
  NAND2_X1 U351 ( .A1(a[1]), .A2(n292), .ZN(n294) );
  XNOR2_X1 U352 ( .A(b[4]), .B(a[1]), .ZN(n342) );
endmodule


module datapath_DW01_add_23 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n75;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n75), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(B[9]), .Z(n1) );
  CLKBUF_X1 U2 ( .A(n23), .Z(n2) );
  NAND3_X1 U3 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n3) );
  CLKBUF_X1 U4 ( .A(carry[12]), .Z(n4) );
  CLKBUF_X1 U5 ( .A(n42), .Z(n5) );
  CLKBUF_X1 U6 ( .A(n63), .Z(n6) );
  NAND3_X1 U7 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n7) );
  NAND3_X1 U8 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n8) );
  NAND3_X1 U9 ( .A1(n62), .A2(n6), .A3(n64), .ZN(n9) );
  NAND3_X1 U10 ( .A1(n42), .A2(n41), .A3(n43), .ZN(n10) );
  NAND3_X1 U11 ( .A1(n41), .A2(n5), .A3(n43), .ZN(n11) );
  NAND3_X1 U12 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n12) );
  NAND3_X1 U13 ( .A1(n21), .A2(n22), .A3(n2), .ZN(n13) );
  NAND3_X1 U14 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n14) );
  NAND3_X1 U15 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n15) );
  XOR2_X1 U16 ( .A(n1), .B(A[9]), .Z(n16) );
  XOR2_X1 U17 ( .A(n9), .B(n16), .Z(SUM[9]) );
  NAND2_X1 U18 ( .A1(n8), .A2(B[9]), .ZN(n17) );
  NAND2_X1 U19 ( .A1(carry[9]), .A2(A[9]), .ZN(n18) );
  NAND2_X1 U20 ( .A1(B[9]), .A2(A[9]), .ZN(n19) );
  NAND3_X1 U21 ( .A1(n17), .A2(n18), .A3(n19), .ZN(carry[10]) );
  XOR2_X1 U22 ( .A(n15), .B(A[5]), .Z(n20) );
  XOR2_X1 U23 ( .A(B[5]), .B(n20), .Z(SUM[5]) );
  NAND2_X1 U24 ( .A1(B[5]), .A2(n14), .ZN(n21) );
  NAND2_X1 U25 ( .A1(B[5]), .A2(A[5]), .ZN(n22) );
  NAND2_X1 U26 ( .A1(carry[5]), .A2(A[5]), .ZN(n23) );
  NAND3_X1 U27 ( .A1(n21), .A2(n22), .A3(n23), .ZN(carry[6]) );
  XOR2_X1 U28 ( .A(B[2]), .B(A[2]), .Z(n24) );
  XOR2_X1 U29 ( .A(carry[2]), .B(n24), .Z(SUM[2]) );
  NAND2_X1 U30 ( .A1(carry[2]), .A2(B[2]), .ZN(n25) );
  NAND2_X1 U31 ( .A1(carry[2]), .A2(A[2]), .ZN(n26) );
  NAND2_X1 U32 ( .A1(B[2]), .A2(A[2]), .ZN(n27) );
  NAND3_X1 U33 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[3]) );
  CLKBUF_X1 U34 ( .A(n52), .Z(n28) );
  CLKBUF_X1 U35 ( .A(n55), .Z(n29) );
  CLKBUF_X1 U36 ( .A(carry[10]), .Z(n30) );
  CLKBUF_X1 U37 ( .A(B[12]), .Z(n31) );
  XOR2_X1 U38 ( .A(B[3]), .B(A[3]), .Z(n32) );
  XOR2_X1 U39 ( .A(carry[3]), .B(n32), .Z(SUM[3]) );
  NAND2_X1 U40 ( .A1(carry[3]), .A2(B[3]), .ZN(n33) );
  NAND2_X1 U41 ( .A1(carry[3]), .A2(A[3]), .ZN(n34) );
  NAND2_X1 U42 ( .A1(B[3]), .A2(A[3]), .ZN(n35) );
  NAND3_X1 U43 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[4]) );
  XOR2_X1 U44 ( .A(B[4]), .B(A[4]), .Z(n36) );
  XOR2_X1 U45 ( .A(n3), .B(n36), .Z(SUM[4]) );
  NAND2_X1 U46 ( .A1(n3), .A2(B[4]), .ZN(n37) );
  NAND2_X1 U47 ( .A1(carry[4]), .A2(A[4]), .ZN(n38) );
  NAND2_X1 U48 ( .A1(B[4]), .A2(A[4]), .ZN(n39) );
  NAND3_X1 U49 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[5]) );
  XOR2_X1 U50 ( .A(B[10]), .B(A[10]), .Z(n40) );
  XOR2_X1 U51 ( .A(n30), .B(n40), .Z(SUM[10]) );
  NAND2_X1 U52 ( .A1(n7), .A2(B[10]), .ZN(n41) );
  NAND2_X1 U53 ( .A1(carry[10]), .A2(A[10]), .ZN(n42) );
  NAND2_X1 U54 ( .A1(B[10]), .A2(A[10]), .ZN(n43) );
  NAND3_X1 U55 ( .A1(n41), .A2(n42), .A3(n43), .ZN(carry[11]) );
  NAND3_X1 U56 ( .A1(n47), .A2(n46), .A3(n48), .ZN(n44) );
  XOR2_X1 U57 ( .A(B[11]), .B(A[11]), .Z(n45) );
  XOR2_X1 U58 ( .A(n11), .B(n45), .Z(SUM[11]) );
  NAND2_X1 U59 ( .A1(n10), .A2(B[11]), .ZN(n46) );
  NAND2_X1 U60 ( .A1(carry[11]), .A2(A[11]), .ZN(n47) );
  NAND2_X1 U61 ( .A1(B[11]), .A2(A[11]), .ZN(n48) );
  NAND3_X1 U62 ( .A1(n46), .A2(n47), .A3(n48), .ZN(carry[12]) );
  NAND3_X1 U63 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n49) );
  NAND3_X1 U64 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n50) );
  NAND3_X1 U65 ( .A1(n54), .A2(n29), .A3(n56), .ZN(n51) );
  NAND3_X1 U66 ( .A1(n69), .A2(n67), .A3(n68), .ZN(n52) );
  XOR2_X1 U67 ( .A(B[6]), .B(A[6]), .Z(n53) );
  XOR2_X1 U68 ( .A(n13), .B(n53), .Z(SUM[6]) );
  NAND2_X1 U69 ( .A1(n12), .A2(B[6]), .ZN(n54) );
  NAND2_X1 U70 ( .A1(carry[6]), .A2(A[6]), .ZN(n55) );
  NAND2_X1 U71 ( .A1(B[6]), .A2(A[6]), .ZN(n56) );
  NAND3_X1 U72 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[7]) );
  XOR2_X1 U73 ( .A(B[7]), .B(A[7]), .Z(n57) );
  XOR2_X1 U74 ( .A(n51), .B(n57), .Z(SUM[7]) );
  NAND2_X1 U75 ( .A1(n50), .A2(B[7]), .ZN(n58) );
  NAND2_X1 U76 ( .A1(carry[7]), .A2(A[7]), .ZN(n59) );
  NAND2_X1 U77 ( .A1(B[7]), .A2(A[7]), .ZN(n60) );
  NAND3_X1 U78 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[8]) );
  XOR2_X1 U79 ( .A(B[8]), .B(A[8]), .Z(n61) );
  XOR2_X1 U80 ( .A(carry[8]), .B(n61), .Z(SUM[8]) );
  NAND2_X1 U81 ( .A1(n49), .A2(B[8]), .ZN(n62) );
  NAND2_X1 U82 ( .A1(carry[8]), .A2(A[8]), .ZN(n63) );
  NAND2_X1 U83 ( .A1(B[8]), .A2(A[8]), .ZN(n64) );
  NAND3_X1 U84 ( .A1(n62), .A2(n63), .A3(n64), .ZN(carry[9]) );
  NAND2_X1 U85 ( .A1(B[12]), .A2(A[12]), .ZN(n67) );
  XNOR2_X1 U86 ( .A(carry[15]), .B(n65), .ZN(SUM[15]) );
  XNOR2_X1 U87 ( .A(B[15]), .B(A[15]), .ZN(n65) );
  XOR2_X1 U88 ( .A(A[12]), .B(n31), .Z(n66) );
  XOR2_X1 U89 ( .A(n66), .B(n4), .Z(SUM[12]) );
  NAND2_X1 U90 ( .A1(A[12]), .A2(n44), .ZN(n68) );
  NAND2_X1 U91 ( .A1(carry[12]), .A2(B[12]), .ZN(n69) );
  NAND3_X1 U92 ( .A1(n67), .A2(n68), .A3(n69), .ZN(carry[13]) );
  XOR2_X1 U93 ( .A(A[13]), .B(B[13]), .Z(n70) );
  XOR2_X1 U94 ( .A(n70), .B(n28), .Z(SUM[13]) );
  NAND2_X1 U95 ( .A1(A[13]), .A2(B[13]), .ZN(n71) );
  NAND2_X1 U96 ( .A1(n52), .A2(A[13]), .ZN(n72) );
  NAND2_X1 U97 ( .A1(B[13]), .A2(carry[13]), .ZN(n73) );
  NAND3_X1 U98 ( .A1(n71), .A2(n72), .A3(n73), .ZN(carry[14]) );
  XOR2_X1 U99 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U100 ( .A1(B[0]), .A2(A[0]), .ZN(n75) );
endmodule


module datapath_DW_mult_tc_22 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n17, n18, n19,
         n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345;

  FA_X1 U4 ( .A(n19), .B(n18), .CI(n4), .CO(n3), .S(product[12]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n288), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n287), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n291), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n290), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n293), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  INV_X1 U157 ( .A(n256), .ZN(n257) );
  NAND2_X1 U158 ( .A1(n24), .A2(n27), .ZN(n222) );
  INV_X1 U159 ( .A(n15), .ZN(n284) );
  AND3_X1 U160 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n211) );
  AND3_X1 U161 ( .A1(n260), .A2(n261), .A3(n262), .ZN(product[15]) );
  NAND3_X1 U162 ( .A1(n222), .A2(n223), .A3(n224), .ZN(n207) );
  NAND3_X1 U163 ( .A1(n222), .A2(n223), .A3(n224), .ZN(n208) );
  CLKBUF_X1 U164 ( .A(n240), .Z(n209) );
  NAND3_X1 U165 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n210) );
  XNOR2_X1 U166 ( .A(n211), .B(n259), .ZN(product[14]) );
  CLKBUF_X1 U167 ( .A(n301), .Z(n212) );
  XOR2_X1 U168 ( .A(n104), .B(n72), .Z(product[1]) );
  CLKBUF_X1 U169 ( .A(n13), .Z(n213) );
  AND2_X1 U170 ( .A1(n104), .A2(n72), .ZN(n214) );
  INV_X1 U171 ( .A(n289), .ZN(n215) );
  XNOR2_X1 U172 ( .A(n216), .B(n218), .ZN(product[4]) );
  XNOR2_X1 U173 ( .A(n54), .B(n55), .ZN(n216) );
  NAND3_X1 U174 ( .A1(n281), .A2(n280), .A3(n279), .ZN(n217) );
  NAND3_X1 U175 ( .A1(n219), .A2(n280), .A3(n279), .ZN(n218) );
  CLKBUF_X1 U176 ( .A(n281), .Z(n219) );
  NAND3_X1 U177 ( .A1(n281), .A2(n280), .A3(n279), .ZN(n12) );
  XNOR2_X1 U178 ( .A(n220), .B(n214), .ZN(product[2]) );
  XNOR2_X1 U179 ( .A(n103), .B(n96), .ZN(n220) );
  XOR2_X1 U180 ( .A(n24), .B(n27), .Z(n221) );
  XOR2_X1 U181 ( .A(n221), .B(n6), .Z(product[10]) );
  NAND2_X1 U182 ( .A1(n24), .A2(n6), .ZN(n223) );
  NAND2_X1 U183 ( .A1(n27), .A2(n6), .ZN(n224) );
  NAND3_X1 U184 ( .A1(n222), .A2(n223), .A3(n224), .ZN(n5) );
  XOR2_X1 U185 ( .A(n20), .B(n23), .Z(n225) );
  XOR2_X1 U186 ( .A(n225), .B(n208), .Z(product[11]) );
  NAND2_X1 U187 ( .A1(n20), .A2(n23), .ZN(n226) );
  NAND2_X1 U188 ( .A1(n20), .A2(n207), .ZN(n227) );
  NAND2_X1 U189 ( .A1(n23), .A2(n5), .ZN(n228) );
  NAND3_X1 U190 ( .A1(n226), .A2(n227), .A3(n228), .ZN(n4) );
  NAND3_X1 U191 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n229) );
  NAND3_X1 U192 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n230) );
  NAND3_X1 U193 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n231) );
  XOR2_X1 U194 ( .A(n46), .B(n49), .Z(n232) );
  XOR2_X1 U195 ( .A(n10), .B(n232), .Z(product[6]) );
  NAND2_X1 U196 ( .A1(n10), .A2(n46), .ZN(n233) );
  NAND2_X1 U197 ( .A1(n10), .A2(n49), .ZN(n234) );
  NAND2_X1 U198 ( .A1(n46), .A2(n49), .ZN(n235) );
  NAND3_X1 U199 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n9) );
  XOR2_X1 U200 ( .A(n17), .B(n284), .Z(n236) );
  XOR2_X1 U201 ( .A(n3), .B(n236), .Z(product[13]) );
  NAND2_X1 U202 ( .A1(n3), .A2(n17), .ZN(n237) );
  NAND2_X1 U203 ( .A1(n3), .A2(n284), .ZN(n238) );
  NAND2_X1 U204 ( .A1(n17), .A2(n284), .ZN(n239) );
  NAND3_X1 U205 ( .A1(n275), .A2(n274), .A3(n273), .ZN(n240) );
  NAND2_X1 U206 ( .A1(n54), .A2(n55), .ZN(n241) );
  NAND2_X1 U207 ( .A1(n54), .A2(n217), .ZN(n242) );
  NAND2_X1 U208 ( .A1(n55), .A2(n12), .ZN(n243) );
  NAND3_X1 U209 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n11) );
  XOR2_X1 U210 ( .A(n50), .B(n53), .Z(n244) );
  XOR2_X1 U211 ( .A(n244), .B(n230), .Z(product[5]) );
  NAND2_X1 U212 ( .A1(n50), .A2(n53), .ZN(n245) );
  NAND2_X1 U213 ( .A1(n50), .A2(n229), .ZN(n246) );
  NAND2_X1 U214 ( .A1(n53), .A2(n11), .ZN(n247) );
  NAND3_X1 U215 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n10) );
  XOR2_X1 U216 ( .A(n33), .B(n28), .Z(n248) );
  XOR2_X1 U217 ( .A(n209), .B(n248), .Z(product[9]) );
  NAND2_X1 U218 ( .A1(n240), .A2(n33), .ZN(n249) );
  NAND2_X1 U219 ( .A1(n7), .A2(n28), .ZN(n250) );
  NAND2_X1 U220 ( .A1(n33), .A2(n28), .ZN(n251) );
  NAND3_X1 U221 ( .A1(n249), .A2(n250), .A3(n251), .ZN(n6) );
  XNOR2_X1 U222 ( .A(n252), .B(n213), .ZN(product[3]) );
  XNOR2_X1 U223 ( .A(n56), .B(n71), .ZN(n252) );
  NAND3_X1 U224 ( .A1(n276), .A2(n277), .A3(n278), .ZN(n253) );
  NAND3_X1 U225 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n254) );
  CLKBUF_X1 U226 ( .A(b[1]), .Z(n255) );
  INV_X1 U227 ( .A(n311), .ZN(n256) );
  CLKBUF_X3 U228 ( .A(a[3]), .Z(n258) );
  XNOR2_X1 U229 ( .A(a[4]), .B(a[3]), .ZN(n311) );
  INV_X2 U230 ( .A(n283), .ZN(n282) );
  XOR2_X1 U231 ( .A(n285), .B(n15), .Z(n259) );
  NAND2_X1 U232 ( .A1(n210), .A2(n285), .ZN(n260) );
  NAND2_X1 U233 ( .A1(n210), .A2(n15), .ZN(n261) );
  NAND2_X1 U234 ( .A1(n285), .A2(n15), .ZN(n262) );
  OAI22_X1 U235 ( .A1(n302), .A2(n303), .B1(n301), .B2(n304), .ZN(n263) );
  XOR2_X1 U236 ( .A(n263), .B(n102), .Z(n264) );
  NAND2_X1 U237 ( .A1(a[2]), .A2(a[1]), .ZN(n266) );
  NAND2_X1 U238 ( .A1(n265), .A2(n294), .ZN(n267) );
  NAND2_X2 U239 ( .A1(n266), .A2(n267), .ZN(n301) );
  INV_X1 U240 ( .A(a[2]), .ZN(n265) );
  XOR2_X1 U241 ( .A(n40), .B(n45), .Z(n268) );
  XOR2_X1 U242 ( .A(n268), .B(n9), .Z(product[7]) );
  NAND2_X1 U243 ( .A1(n40), .A2(n45), .ZN(n269) );
  NAND2_X1 U244 ( .A1(n40), .A2(n231), .ZN(n270) );
  NAND2_X1 U245 ( .A1(n231), .A2(n45), .ZN(n271) );
  NAND3_X1 U246 ( .A1(n270), .A2(n269), .A3(n271), .ZN(n8) );
  XOR2_X1 U247 ( .A(n34), .B(n39), .Z(n272) );
  XOR2_X1 U248 ( .A(n272), .B(n254), .Z(product[8]) );
  NAND2_X1 U249 ( .A1(n34), .A2(n39), .ZN(n273) );
  NAND2_X1 U250 ( .A1(n34), .A2(n8), .ZN(n274) );
  NAND2_X1 U251 ( .A1(n39), .A2(n8), .ZN(n275) );
  NAND3_X1 U252 ( .A1(n274), .A2(n273), .A3(n275), .ZN(n7) );
  NAND2_X1 U253 ( .A1(n103), .A2(n96), .ZN(n276) );
  NAND2_X1 U254 ( .A1(n103), .A2(n214), .ZN(n277) );
  NAND2_X1 U255 ( .A1(n96), .A2(n214), .ZN(n278) );
  NAND3_X1 U256 ( .A1(n278), .A2(n277), .A3(n276), .ZN(n13) );
  NAND2_X1 U257 ( .A1(n264), .A2(n71), .ZN(n279) );
  NAND2_X1 U258 ( .A1(n264), .A2(n253), .ZN(n280) );
  NAND2_X1 U259 ( .A1(n71), .A2(n13), .ZN(n281) );
  INV_X1 U260 ( .A(n21), .ZN(n287) );
  INV_X1 U261 ( .A(n320), .ZN(n288) );
  INV_X1 U262 ( .A(n331), .ZN(n285) );
  INV_X1 U263 ( .A(n300), .ZN(n293) );
  INV_X1 U264 ( .A(n309), .ZN(n291) );
  INV_X1 U265 ( .A(n31), .ZN(n290) );
  INV_X1 U266 ( .A(b[0]), .ZN(n283) );
  INV_X1 U267 ( .A(a[5]), .ZN(n289) );
  INV_X1 U268 ( .A(a[7]), .ZN(n286) );
  INV_X1 U269 ( .A(a[3]), .ZN(n292) );
  NAND2_X2 U270 ( .A1(n311), .A2(n340), .ZN(n313) );
  INV_X1 U271 ( .A(a[1]), .ZN(n294) );
  NAND2_X2 U272 ( .A1(n301), .A2(n339), .ZN(n303) );
  XOR2_X2 U273 ( .A(a[6]), .B(n289), .Z(n322) );
  INV_X2 U274 ( .A(a[0]), .ZN(n295) );
  NOR2_X1 U275 ( .A1(n295), .A2(n283), .ZN(product[0]) );
  OAI22_X1 U276 ( .A1(n296), .A2(n297), .B1(n298), .B2(n295), .ZN(n99) );
  OAI22_X1 U277 ( .A1(n298), .A2(n297), .B1(n299), .B2(n295), .ZN(n98) );
  XNOR2_X1 U278 ( .A(b[6]), .B(a[1]), .ZN(n298) );
  OAI22_X1 U279 ( .A1(n295), .A2(n299), .B1(n297), .B2(n299), .ZN(n300) );
  XNOR2_X1 U280 ( .A(b[7]), .B(a[1]), .ZN(n299) );
  NOR2_X1 U281 ( .A1(n301), .A2(n283), .ZN(n96) );
  OAI22_X1 U282 ( .A1(n302), .A2(n303), .B1(n301), .B2(n304), .ZN(n95) );
  XNOR2_X1 U283 ( .A(n258), .B(n282), .ZN(n302) );
  OAI22_X1 U284 ( .A1(n304), .A2(n303), .B1(n301), .B2(n305), .ZN(n94) );
  XNOR2_X1 U285 ( .A(b[1]), .B(n258), .ZN(n304) );
  OAI22_X1 U286 ( .A1(n305), .A2(n303), .B1(n301), .B2(n306), .ZN(n93) );
  XNOR2_X1 U287 ( .A(b[2]), .B(n258), .ZN(n305) );
  OAI22_X1 U288 ( .A1(n306), .A2(n303), .B1(n301), .B2(n307), .ZN(n92) );
  XNOR2_X1 U289 ( .A(b[3]), .B(n258), .ZN(n306) );
  OAI22_X1 U290 ( .A1(n307), .A2(n303), .B1(n301), .B2(n308), .ZN(n91) );
  XNOR2_X1 U291 ( .A(b[4]), .B(n258), .ZN(n307) );
  OAI22_X1 U292 ( .A1(n310), .A2(n212), .B1(n303), .B2(n310), .ZN(n309) );
  NOR2_X1 U293 ( .A1(n311), .A2(n283), .ZN(n88) );
  OAI22_X1 U294 ( .A1(n312), .A2(n313), .B1(n311), .B2(n314), .ZN(n87) );
  XNOR2_X1 U295 ( .A(a[5]), .B(n282), .ZN(n312) );
  OAI22_X1 U296 ( .A1(n314), .A2(n313), .B1(n257), .B2(n315), .ZN(n86) );
  XNOR2_X1 U297 ( .A(b[1]), .B(a[5]), .ZN(n314) );
  OAI22_X1 U298 ( .A1(n315), .A2(n313), .B1(n257), .B2(n316), .ZN(n85) );
  XNOR2_X1 U299 ( .A(b[2]), .B(n215), .ZN(n315) );
  OAI22_X1 U300 ( .A1(n316), .A2(n313), .B1(n257), .B2(n317), .ZN(n84) );
  XNOR2_X1 U301 ( .A(b[3]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U302 ( .A1(n317), .A2(n313), .B1(n257), .B2(n318), .ZN(n83) );
  XNOR2_X1 U303 ( .A(b[4]), .B(n215), .ZN(n317) );
  OAI22_X1 U304 ( .A1(n318), .A2(n313), .B1(n257), .B2(n319), .ZN(n82) );
  XNOR2_X1 U305 ( .A(b[5]), .B(n215), .ZN(n318) );
  OAI22_X1 U306 ( .A1(n321), .A2(n257), .B1(n313), .B2(n321), .ZN(n320) );
  NOR2_X1 U307 ( .A1(n322), .A2(n283), .ZN(n80) );
  OAI22_X1 U308 ( .A1(n323), .A2(n324), .B1(n322), .B2(n325), .ZN(n79) );
  XNOR2_X1 U309 ( .A(a[7]), .B(n282), .ZN(n323) );
  OAI22_X1 U310 ( .A1(n326), .A2(n324), .B1(n322), .B2(n327), .ZN(n77) );
  OAI22_X1 U311 ( .A1(n327), .A2(n324), .B1(n322), .B2(n328), .ZN(n76) );
  XNOR2_X1 U312 ( .A(b[3]), .B(a[7]), .ZN(n327) );
  OAI22_X1 U313 ( .A1(n328), .A2(n324), .B1(n322), .B2(n329), .ZN(n75) );
  XNOR2_X1 U314 ( .A(b[4]), .B(a[7]), .ZN(n328) );
  OAI22_X1 U315 ( .A1(n329), .A2(n324), .B1(n322), .B2(n330), .ZN(n74) );
  XNOR2_X1 U316 ( .A(b[5]), .B(a[7]), .ZN(n329) );
  OAI22_X1 U317 ( .A1(n332), .A2(n322), .B1(n324), .B2(n332), .ZN(n331) );
  OAI21_X1 U318 ( .B1(n282), .B2(n294), .A(n297), .ZN(n72) );
  OAI21_X1 U319 ( .B1(n292), .B2(n303), .A(n333), .ZN(n71) );
  OR3_X1 U320 ( .A1(n301), .A2(n282), .A3(n292), .ZN(n333) );
  OAI21_X1 U321 ( .B1(n289), .B2(n313), .A(n334), .ZN(n70) );
  OR3_X1 U322 ( .A1(n311), .A2(n282), .A3(n289), .ZN(n334) );
  OAI21_X1 U323 ( .B1(n286), .B2(n324), .A(n335), .ZN(n69) );
  OR3_X1 U324 ( .A1(n322), .A2(n282), .A3(n286), .ZN(n335) );
  XNOR2_X1 U325 ( .A(n336), .B(n337), .ZN(n38) );
  OR2_X1 U326 ( .A1(n336), .A2(n337), .ZN(n37) );
  OAI22_X1 U327 ( .A1(n308), .A2(n303), .B1(n212), .B2(n338), .ZN(n337) );
  XNOR2_X1 U328 ( .A(b[5]), .B(n258), .ZN(n308) );
  OAI22_X1 U329 ( .A1(n325), .A2(n324), .B1(n322), .B2(n326), .ZN(n336) );
  XNOR2_X1 U330 ( .A(b[2]), .B(a[7]), .ZN(n326) );
  XNOR2_X1 U331 ( .A(n255), .B(a[7]), .ZN(n325) );
  OAI22_X1 U332 ( .A1(n338), .A2(n303), .B1(n212), .B2(n310), .ZN(n31) );
  XNOR2_X1 U333 ( .A(b[7]), .B(n258), .ZN(n310) );
  XNOR2_X1 U334 ( .A(n292), .B(a[2]), .ZN(n339) );
  XNOR2_X1 U335 ( .A(b[6]), .B(n258), .ZN(n338) );
  OAI22_X1 U336 ( .A1(n319), .A2(n313), .B1(n257), .B2(n321), .ZN(n21) );
  XNOR2_X1 U337 ( .A(b[7]), .B(n215), .ZN(n321) );
  XNOR2_X1 U338 ( .A(n289), .B(a[4]), .ZN(n340) );
  XNOR2_X1 U339 ( .A(b[6]), .B(n215), .ZN(n319) );
  OAI22_X1 U340 ( .A1(n330), .A2(n324), .B1(n322), .B2(n332), .ZN(n15) );
  XNOR2_X1 U341 ( .A(b[7]), .B(a[7]), .ZN(n332) );
  NAND2_X1 U342 ( .A1(n322), .A2(n341), .ZN(n324) );
  XNOR2_X1 U343 ( .A(n286), .B(a[6]), .ZN(n341) );
  XNOR2_X1 U344 ( .A(b[6]), .B(a[7]), .ZN(n330) );
  OAI22_X1 U345 ( .A1(n282), .A2(n297), .B1(n342), .B2(n295), .ZN(n104) );
  OAI22_X1 U346 ( .A1(n297), .A2(n342), .B1(n343), .B2(n295), .ZN(n103) );
  XNOR2_X1 U347 ( .A(b[1]), .B(a[1]), .ZN(n342) );
  OAI22_X1 U348 ( .A1(n343), .A2(n297), .B1(n344), .B2(n295), .ZN(n102) );
  XNOR2_X1 U349 ( .A(b[2]), .B(a[1]), .ZN(n343) );
  OAI22_X1 U350 ( .A1(n344), .A2(n297), .B1(n345), .B2(n295), .ZN(n101) );
  XNOR2_X1 U351 ( .A(b[3]), .B(a[1]), .ZN(n344) );
  OAI22_X1 U352 ( .A1(n345), .A2(n297), .B1(n296), .B2(n295), .ZN(n100) );
  XNOR2_X1 U353 ( .A(b[5]), .B(a[1]), .ZN(n296) );
  NAND2_X1 U354 ( .A1(a[1]), .A2(n295), .ZN(n297) );
  XNOR2_X1 U355 ( .A(b[4]), .B(a[1]), .ZN(n345) );
endmodule


module datapath_DW01_add_22 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n73;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n73), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(B[9]), .Z(n1) );
  NAND3_X1 U2 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n2) );
  NAND3_X1 U3 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n3) );
  CLKBUF_X1 U4 ( .A(n33), .Z(n4) );
  NAND3_X1 U5 ( .A1(n60), .A2(n61), .A3(n62), .ZN(n5) );
  NAND3_X1 U6 ( .A1(n60), .A2(n61), .A3(n62), .ZN(n6) );
  NAND3_X1 U7 ( .A1(n19), .A2(n18), .A3(n20), .ZN(n7) );
  CLKBUF_X1 U8 ( .A(n25), .Z(n8) );
  CLKBUF_X1 U9 ( .A(n42), .Z(n9) );
  CLKBUF_X1 U10 ( .A(B[5]), .Z(n10) );
  NAND3_X1 U11 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n11) );
  NAND3_X1 U12 ( .A1(n41), .A2(n9), .A3(n43), .ZN(n12) );
  XOR2_X1 U13 ( .A(B[2]), .B(A[2]), .Z(n13) );
  XOR2_X1 U14 ( .A(carry[2]), .B(n13), .Z(SUM[2]) );
  NAND2_X1 U15 ( .A1(carry[2]), .A2(B[2]), .ZN(n14) );
  NAND2_X1 U16 ( .A1(carry[2]), .A2(A[2]), .ZN(n15) );
  NAND2_X1 U17 ( .A1(B[2]), .A2(A[2]), .ZN(n16) );
  NAND3_X1 U18 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[3]) );
  XOR2_X1 U19 ( .A(n1), .B(A[9]), .Z(n17) );
  XOR2_X1 U20 ( .A(n6), .B(n17), .Z(SUM[9]) );
  NAND2_X1 U21 ( .A1(n5), .A2(B[9]), .ZN(n18) );
  NAND2_X1 U22 ( .A1(carry[9]), .A2(A[9]), .ZN(n19) );
  NAND2_X1 U23 ( .A1(B[9]), .A2(A[9]), .ZN(n20) );
  NAND3_X1 U24 ( .A1(n18), .A2(n19), .A3(n20), .ZN(carry[10]) );
  NAND3_X1 U25 ( .A1(n41), .A2(n42), .A3(n43), .ZN(carry[12]) );
  CLKBUF_X1 U26 ( .A(n50), .Z(n21) );
  NAND3_X1 U27 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n22) );
  NAND3_X1 U28 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n23) );
  NAND3_X1 U29 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n24) );
  NAND3_X1 U30 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n25) );
  NAND3_X1 U31 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n26) );
  CLKBUF_X1 U32 ( .A(B[12]), .Z(n27) );
  XOR2_X1 U33 ( .A(n3), .B(A[3]), .Z(n28) );
  XOR2_X1 U34 ( .A(B[3]), .B(n28), .Z(SUM[3]) );
  NAND2_X1 U35 ( .A1(n2), .A2(B[3]), .ZN(n29) );
  NAND2_X1 U36 ( .A1(B[3]), .A2(A[3]), .ZN(n30) );
  NAND2_X1 U37 ( .A1(carry[3]), .A2(A[3]), .ZN(n31) );
  NAND3_X1 U38 ( .A1(n29), .A2(n30), .A3(n31), .ZN(carry[4]) );
  XOR2_X1 U39 ( .A(n7), .B(A[10]), .Z(n32) );
  XOR2_X1 U40 ( .A(B[10]), .B(n32), .Z(SUM[10]) );
  NAND2_X1 U41 ( .A1(B[10]), .A2(n7), .ZN(n33) );
  NAND2_X1 U42 ( .A1(B[10]), .A2(A[10]), .ZN(n34) );
  NAND2_X1 U43 ( .A1(carry[10]), .A2(A[10]), .ZN(n35) );
  NAND3_X1 U44 ( .A1(n4), .A2(n34), .A3(n35), .ZN(carry[11]) );
  XOR2_X1 U45 ( .A(n10), .B(A[5]), .Z(n36) );
  XOR2_X1 U46 ( .A(n22), .B(n36), .Z(SUM[5]) );
  NAND2_X1 U47 ( .A1(n22), .A2(B[5]), .ZN(n37) );
  NAND2_X1 U48 ( .A1(carry[5]), .A2(A[5]), .ZN(n38) );
  NAND2_X1 U49 ( .A1(B[5]), .A2(A[5]), .ZN(n39) );
  NAND3_X1 U50 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[6]) );
  XOR2_X1 U51 ( .A(B[11]), .B(A[11]), .Z(n40) );
  XOR2_X1 U52 ( .A(carry[11]), .B(n40), .Z(SUM[11]) );
  NAND2_X1 U53 ( .A1(n24), .A2(B[11]), .ZN(n41) );
  NAND2_X1 U54 ( .A1(n24), .A2(A[11]), .ZN(n42) );
  NAND2_X1 U55 ( .A1(B[11]), .A2(A[11]), .ZN(n43) );
  XOR2_X1 U56 ( .A(B[4]), .B(A[4]), .Z(n44) );
  XOR2_X1 U57 ( .A(carry[4]), .B(n44), .Z(SUM[4]) );
  NAND2_X1 U58 ( .A1(n26), .A2(B[4]), .ZN(n45) );
  NAND2_X1 U59 ( .A1(n26), .A2(A[4]), .ZN(n46) );
  NAND2_X1 U60 ( .A1(B[4]), .A2(A[4]), .ZN(n47) );
  NAND3_X1 U61 ( .A1(n45), .A2(n46), .A3(n47), .ZN(carry[5]) );
  NAND3_X1 U62 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n48) );
  NAND3_X1 U63 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n49) );
  NAND3_X1 U64 ( .A1(n67), .A2(n65), .A3(n66), .ZN(n50) );
  XOR2_X1 U65 ( .A(B[6]), .B(A[6]), .Z(n51) );
  XOR2_X1 U66 ( .A(n23), .B(n51), .Z(SUM[6]) );
  NAND2_X1 U67 ( .A1(n23), .A2(B[6]), .ZN(n52) );
  NAND2_X1 U68 ( .A1(carry[6]), .A2(A[6]), .ZN(n53) );
  NAND2_X1 U69 ( .A1(B[6]), .A2(A[6]), .ZN(n54) );
  NAND3_X1 U70 ( .A1(n52), .A2(n53), .A3(n54), .ZN(carry[7]) );
  XOR2_X1 U71 ( .A(B[7]), .B(A[7]), .Z(n55) );
  XOR2_X1 U72 ( .A(n49), .B(n55), .Z(SUM[7]) );
  NAND2_X1 U73 ( .A1(n49), .A2(B[7]), .ZN(n56) );
  NAND2_X1 U74 ( .A1(carry[7]), .A2(A[7]), .ZN(n57) );
  NAND2_X1 U75 ( .A1(B[7]), .A2(A[7]), .ZN(n58) );
  XOR2_X1 U76 ( .A(B[8]), .B(A[8]), .Z(n59) );
  XOR2_X1 U77 ( .A(n8), .B(n59), .Z(SUM[8]) );
  NAND2_X1 U78 ( .A1(n25), .A2(B[8]), .ZN(n60) );
  NAND2_X1 U79 ( .A1(n48), .A2(A[8]), .ZN(n61) );
  NAND2_X1 U80 ( .A1(B[8]), .A2(A[8]), .ZN(n62) );
  NAND3_X1 U81 ( .A1(n60), .A2(n61), .A3(n62), .ZN(carry[9]) );
  NAND2_X1 U82 ( .A1(A[12]), .A2(B[12]), .ZN(n65) );
  XNOR2_X1 U83 ( .A(carry[15]), .B(n63), .ZN(SUM[15]) );
  XNOR2_X1 U84 ( .A(B[15]), .B(A[15]), .ZN(n63) );
  XOR2_X1 U85 ( .A(A[12]), .B(n27), .Z(n64) );
  XOR2_X1 U86 ( .A(n64), .B(n12), .Z(SUM[12]) );
  NAND2_X1 U87 ( .A1(carry[12]), .A2(A[12]), .ZN(n66) );
  NAND2_X1 U88 ( .A1(B[12]), .A2(n11), .ZN(n67) );
  NAND3_X1 U89 ( .A1(n65), .A2(n66), .A3(n67), .ZN(carry[13]) );
  XOR2_X1 U90 ( .A(A[13]), .B(B[13]), .Z(n68) );
  XOR2_X1 U91 ( .A(n68), .B(n21), .Z(SUM[13]) );
  NAND2_X1 U92 ( .A1(A[13]), .A2(B[13]), .ZN(n69) );
  NAND2_X1 U93 ( .A1(n50), .A2(A[13]), .ZN(n70) );
  NAND2_X1 U94 ( .A1(B[13]), .A2(carry[13]), .ZN(n71) );
  NAND3_X1 U95 ( .A1(n69), .A2(n70), .A3(n71), .ZN(carry[14]) );
  XOR2_X1 U96 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U97 ( .A1(B[0]), .A2(A[0]), .ZN(n73) );
endmodule


module datapath_DW_mult_tc_21 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347;

  FA_X1 U11 ( .A(n50), .B(n53), .CI(n11), .CO(n10), .S(product[5]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n290), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n289), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n293), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n292), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n295), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  INV_X1 U157 ( .A(n285), .ZN(n284) );
  INV_X1 U158 ( .A(n15), .ZN(n286) );
  CLKBUF_X1 U159 ( .A(n2), .Z(n206) );
  AND2_X1 U160 ( .A1(n225), .A2(n102), .ZN(n207) );
  AND3_X1 U161 ( .A1(n227), .A2(n228), .A3(n229), .ZN(product[15]) );
  NAND3_X1 U162 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n209) );
  NAND3_X1 U163 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n210) );
  NAND3_X1 U164 ( .A1(n231), .A2(n232), .A3(n233), .ZN(n211) );
  NAND3_X1 U165 ( .A1(n231), .A2(n232), .A3(n233), .ZN(n212) );
  NAND3_X1 U166 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n213) );
  NAND3_X1 U167 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n214) );
  BUF_X1 U168 ( .A(n10), .Z(n217) );
  NAND3_X1 U169 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n215) );
  BUF_X1 U170 ( .A(n344), .Z(n236) );
  XOR2_X2 U171 ( .A(a[6]), .B(n291), .Z(n324) );
  NAND3_X1 U172 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n216) );
  XOR2_X1 U173 ( .A(n17), .B(n286), .Z(n218) );
  XOR2_X1 U174 ( .A(n210), .B(n218), .Z(product[13]) );
  NAND2_X1 U175 ( .A1(n209), .A2(n17), .ZN(n219) );
  NAND2_X1 U176 ( .A1(n3), .A2(n286), .ZN(n220) );
  NAND2_X1 U177 ( .A1(n17), .A2(n286), .ZN(n221) );
  NAND3_X1 U178 ( .A1(n219), .A2(n220), .A3(n221), .ZN(n2) );
  NAND3_X1 U179 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n222) );
  XOR2_X1 U180 ( .A(n95), .B(n102), .Z(n223) );
  OAI22_X1 U181 ( .A1(n236), .A2(n299), .B1(n345), .B2(n297), .ZN(n224) );
  BUF_X1 U182 ( .A(n14), .Z(n247) );
  OAI22_X1 U183 ( .A1(n304), .A2(n305), .B1(n282), .B2(n306), .ZN(n225) );
  XOR2_X1 U184 ( .A(n287), .B(n15), .Z(n226) );
  XOR2_X1 U185 ( .A(n2), .B(n226), .Z(product[14]) );
  NAND2_X1 U186 ( .A1(n206), .A2(n287), .ZN(n227) );
  NAND2_X1 U187 ( .A1(n2), .A2(n15), .ZN(n228) );
  NAND2_X1 U188 ( .A1(n287), .A2(n15), .ZN(n229) );
  XOR2_X1 U189 ( .A(n34), .B(n39), .Z(n230) );
  XOR2_X1 U190 ( .A(n215), .B(n230), .Z(product[8]) );
  NAND2_X1 U191 ( .A1(n222), .A2(n34), .ZN(n231) );
  NAND2_X1 U192 ( .A1(n8), .A2(n39), .ZN(n232) );
  NAND2_X1 U193 ( .A1(n34), .A2(n39), .ZN(n233) );
  NAND3_X1 U194 ( .A1(n231), .A2(n232), .A3(n233), .ZN(n7) );
  NAND3_X1 U195 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n234) );
  NAND3_X1 U196 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n235) );
  XNOR2_X1 U197 ( .A(n238), .B(n237), .ZN(product[4]) );
  XNOR2_X1 U198 ( .A(n54), .B(n207), .ZN(n237) );
  CLKBUF_X1 U199 ( .A(n12), .Z(n238) );
  XOR2_X1 U200 ( .A(n225), .B(n102), .Z(n239) );
  XOR2_X1 U201 ( .A(n18), .B(n19), .Z(n240) );
  XOR2_X1 U202 ( .A(n235), .B(n240), .Z(product[12]) );
  NAND2_X1 U203 ( .A1(n234), .A2(n18), .ZN(n241) );
  NAND2_X1 U204 ( .A1(n4), .A2(n19), .ZN(n242) );
  NAND2_X1 U205 ( .A1(n18), .A2(n19), .ZN(n243) );
  NAND3_X1 U206 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n3) );
  NAND2_X1 U207 ( .A1(n12), .A2(n54), .ZN(n244) );
  NAND2_X1 U208 ( .A1(n12), .A2(n207), .ZN(n245) );
  NAND2_X1 U209 ( .A1(n54), .A2(n207), .ZN(n246) );
  NAND3_X1 U210 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n11) );
  XNOR2_X1 U211 ( .A(n248), .B(n247), .ZN(product[2]) );
  XNOR2_X1 U212 ( .A(n103), .B(n96), .ZN(n248) );
  XNOR2_X1 U213 ( .A(n249), .B(n214), .ZN(product[3]) );
  XNOR2_X1 U214 ( .A(n239), .B(n71), .ZN(n249) );
  XOR2_X1 U215 ( .A(n46), .B(n49), .Z(n250) );
  XOR2_X1 U216 ( .A(n217), .B(n250), .Z(product[6]) );
  NAND2_X1 U217 ( .A1(n10), .A2(n46), .ZN(n251) );
  NAND2_X1 U218 ( .A1(n10), .A2(n49), .ZN(n252) );
  NAND2_X1 U219 ( .A1(n46), .A2(n49), .ZN(n253) );
  NAND3_X1 U220 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n9) );
  XOR2_X1 U221 ( .A(n40), .B(n45), .Z(n254) );
  XOR2_X1 U222 ( .A(n9), .B(n254), .Z(product[7]) );
  NAND2_X1 U223 ( .A1(n216), .A2(n40), .ZN(n255) );
  NAND2_X1 U224 ( .A1(n9), .A2(n45), .ZN(n256) );
  NAND2_X1 U225 ( .A1(n40), .A2(n45), .ZN(n257) );
  NAND3_X1 U226 ( .A1(n256), .A2(n255), .A3(n257), .ZN(n8) );
  NAND2_X1 U227 ( .A1(n224), .A2(n96), .ZN(n258) );
  NAND2_X1 U228 ( .A1(n224), .A2(n14), .ZN(n259) );
  NAND2_X1 U229 ( .A1(n96), .A2(n14), .ZN(n260) );
  NAND3_X1 U230 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n13) );
  NAND2_X1 U231 ( .A1(n223), .A2(n71), .ZN(n261) );
  NAND2_X1 U232 ( .A1(n223), .A2(n213), .ZN(n262) );
  NAND2_X1 U233 ( .A1(n71), .A2(n13), .ZN(n263) );
  NAND3_X1 U234 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n12) );
  BUF_X1 U235 ( .A(b[1]), .Z(n271) );
  NAND3_X1 U236 ( .A1(n279), .A2(n278), .A3(n277), .ZN(n264) );
  XOR2_X1 U237 ( .A(n23), .B(n20), .Z(n265) );
  XOR2_X1 U238 ( .A(n264), .B(n265), .Z(product[11]) );
  NAND2_X1 U239 ( .A1(n264), .A2(n23), .ZN(n266) );
  NAND2_X1 U240 ( .A1(n5), .A2(n20), .ZN(n267) );
  NAND2_X1 U241 ( .A1(n23), .A2(n20), .ZN(n268) );
  NAND3_X1 U242 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n4) );
  NAND3_X1 U243 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n269) );
  NAND3_X1 U244 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n270) );
  XOR2_X1 U245 ( .A(n28), .B(n33), .Z(n272) );
  XOR2_X1 U246 ( .A(n272), .B(n212), .Z(product[9]) );
  NAND2_X1 U247 ( .A1(n28), .A2(n33), .ZN(n273) );
  NAND2_X1 U248 ( .A1(n28), .A2(n211), .ZN(n274) );
  NAND2_X1 U249 ( .A1(n33), .A2(n7), .ZN(n275) );
  NAND3_X1 U250 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n6) );
  XOR2_X1 U251 ( .A(n24), .B(n27), .Z(n276) );
  XOR2_X1 U252 ( .A(n276), .B(n270), .Z(product[10]) );
  NAND2_X1 U253 ( .A1(n24), .A2(n27), .ZN(n277) );
  NAND2_X1 U254 ( .A1(n24), .A2(n269), .ZN(n278) );
  NAND2_X1 U255 ( .A1(n27), .A2(n6), .ZN(n279) );
  NAND3_X1 U256 ( .A1(n277), .A2(n278), .A3(n279), .ZN(n5) );
  INV_X1 U257 ( .A(n280), .ZN(n281) );
  INV_X1 U258 ( .A(n313), .ZN(n280) );
  XNOR2_X2 U259 ( .A(a[2]), .B(a[1]), .ZN(n282) );
  XOR2_X1 U260 ( .A(a[4]), .B(n294), .Z(n313) );
  INV_X1 U261 ( .A(n21), .ZN(n289) );
  INV_X1 U262 ( .A(n322), .ZN(n290) );
  INV_X1 U263 ( .A(n333), .ZN(n287) );
  INV_X1 U264 ( .A(n302), .ZN(n295) );
  INV_X1 U265 ( .A(n311), .ZN(n293) );
  INV_X1 U266 ( .A(n31), .ZN(n292) );
  INV_X1 U267 ( .A(b[0]), .ZN(n285) );
  XNOR2_X1 U268 ( .A(a[2]), .B(a[1]), .ZN(n303) );
  NAND2_X1 U269 ( .A1(n313), .A2(n342), .ZN(n315) );
  INV_X1 U270 ( .A(n294), .ZN(n283) );
  NAND2_X1 U271 ( .A1(n303), .A2(n341), .ZN(n305) );
  INV_X1 U272 ( .A(a[0]), .ZN(n297) );
  INV_X1 U273 ( .A(a[5]), .ZN(n291) );
  INV_X1 U274 ( .A(a[7]), .ZN(n288) );
  INV_X1 U275 ( .A(a[3]), .ZN(n294) );
  INV_X1 U276 ( .A(a[1]), .ZN(n296) );
  NOR2_X1 U277 ( .A1(n297), .A2(n285), .ZN(product[0]) );
  OAI22_X1 U278 ( .A1(n298), .A2(n299), .B1(n300), .B2(n297), .ZN(n99) );
  OAI22_X1 U279 ( .A1(n300), .A2(n299), .B1(n301), .B2(n297), .ZN(n98) );
  XNOR2_X1 U280 ( .A(b[6]), .B(a[1]), .ZN(n300) );
  OAI22_X1 U281 ( .A1(n297), .A2(n301), .B1(n299), .B2(n301), .ZN(n302) );
  XNOR2_X1 U282 ( .A(b[7]), .B(a[1]), .ZN(n301) );
  NOR2_X1 U283 ( .A1(n282), .A2(n285), .ZN(n96) );
  OAI22_X1 U284 ( .A1(n304), .A2(n305), .B1(n282), .B2(n306), .ZN(n95) );
  XNOR2_X1 U285 ( .A(n283), .B(n284), .ZN(n304) );
  OAI22_X1 U286 ( .A1(n306), .A2(n305), .B1(n282), .B2(n307), .ZN(n94) );
  XNOR2_X1 U287 ( .A(n271), .B(n283), .ZN(n306) );
  OAI22_X1 U288 ( .A1(n307), .A2(n305), .B1(n282), .B2(n308), .ZN(n93) );
  XNOR2_X1 U289 ( .A(b[2]), .B(n283), .ZN(n307) );
  OAI22_X1 U290 ( .A1(n308), .A2(n305), .B1(n282), .B2(n309), .ZN(n92) );
  XNOR2_X1 U291 ( .A(b[3]), .B(n283), .ZN(n308) );
  OAI22_X1 U292 ( .A1(n309), .A2(n305), .B1(n282), .B2(n310), .ZN(n91) );
  XNOR2_X1 U293 ( .A(b[4]), .B(n283), .ZN(n309) );
  OAI22_X1 U294 ( .A1(n312), .A2(n282), .B1(n305), .B2(n312), .ZN(n311) );
  NOR2_X1 U295 ( .A1(n313), .A2(n285), .ZN(n88) );
  OAI22_X1 U296 ( .A1(n314), .A2(n315), .B1(n281), .B2(n316), .ZN(n87) );
  XNOR2_X1 U297 ( .A(a[5]), .B(n284), .ZN(n314) );
  OAI22_X1 U298 ( .A1(n316), .A2(n315), .B1(n281), .B2(n317), .ZN(n86) );
  XNOR2_X1 U299 ( .A(n271), .B(a[5]), .ZN(n316) );
  OAI22_X1 U300 ( .A1(n317), .A2(n315), .B1(n281), .B2(n318), .ZN(n85) );
  XNOR2_X1 U301 ( .A(b[2]), .B(a[5]), .ZN(n317) );
  OAI22_X1 U302 ( .A1(n318), .A2(n315), .B1(n281), .B2(n319), .ZN(n84) );
  XNOR2_X1 U303 ( .A(b[3]), .B(a[5]), .ZN(n318) );
  OAI22_X1 U304 ( .A1(n319), .A2(n315), .B1(n281), .B2(n320), .ZN(n83) );
  XNOR2_X1 U305 ( .A(b[4]), .B(a[5]), .ZN(n319) );
  OAI22_X1 U306 ( .A1(n320), .A2(n315), .B1(n281), .B2(n321), .ZN(n82) );
  XNOR2_X1 U307 ( .A(b[5]), .B(a[5]), .ZN(n320) );
  OAI22_X1 U308 ( .A1(n323), .A2(n281), .B1(n315), .B2(n323), .ZN(n322) );
  NOR2_X1 U309 ( .A1(n324), .A2(n285), .ZN(n80) );
  OAI22_X1 U310 ( .A1(n325), .A2(n326), .B1(n324), .B2(n327), .ZN(n79) );
  XNOR2_X1 U311 ( .A(a[7]), .B(n284), .ZN(n325) );
  OAI22_X1 U312 ( .A1(n328), .A2(n326), .B1(n324), .B2(n329), .ZN(n77) );
  OAI22_X1 U313 ( .A1(n329), .A2(n326), .B1(n324), .B2(n330), .ZN(n76) );
  XNOR2_X1 U314 ( .A(b[3]), .B(a[7]), .ZN(n329) );
  OAI22_X1 U315 ( .A1(n330), .A2(n326), .B1(n324), .B2(n331), .ZN(n75) );
  XNOR2_X1 U316 ( .A(b[4]), .B(a[7]), .ZN(n330) );
  OAI22_X1 U317 ( .A1(n331), .A2(n326), .B1(n324), .B2(n332), .ZN(n74) );
  XNOR2_X1 U318 ( .A(b[5]), .B(a[7]), .ZN(n331) );
  OAI22_X1 U319 ( .A1(n334), .A2(n324), .B1(n326), .B2(n334), .ZN(n333) );
  OAI21_X1 U320 ( .B1(n284), .B2(n296), .A(n299), .ZN(n72) );
  OAI21_X1 U321 ( .B1(n294), .B2(n305), .A(n335), .ZN(n71) );
  OR3_X1 U322 ( .A1(n282), .A2(n284), .A3(n294), .ZN(n335) );
  OAI21_X1 U323 ( .B1(n291), .B2(n315), .A(n336), .ZN(n70) );
  OR3_X1 U324 ( .A1(n313), .A2(n284), .A3(n291), .ZN(n336) );
  OAI21_X1 U325 ( .B1(n288), .B2(n326), .A(n337), .ZN(n69) );
  OR3_X1 U326 ( .A1(n324), .A2(n284), .A3(n288), .ZN(n337) );
  XNOR2_X1 U327 ( .A(n338), .B(n339), .ZN(n38) );
  OR2_X1 U328 ( .A1(n338), .A2(n339), .ZN(n37) );
  OAI22_X1 U329 ( .A1(n310), .A2(n305), .B1(n282), .B2(n340), .ZN(n339) );
  XNOR2_X1 U330 ( .A(b[5]), .B(n283), .ZN(n310) );
  OAI22_X1 U331 ( .A1(n327), .A2(n326), .B1(n324), .B2(n328), .ZN(n338) );
  XNOR2_X1 U332 ( .A(b[2]), .B(a[7]), .ZN(n328) );
  XNOR2_X1 U333 ( .A(n271), .B(a[7]), .ZN(n327) );
  OAI22_X1 U334 ( .A1(n340), .A2(n305), .B1(n282), .B2(n312), .ZN(n31) );
  XNOR2_X1 U335 ( .A(b[7]), .B(n283), .ZN(n312) );
  XNOR2_X1 U336 ( .A(n294), .B(a[2]), .ZN(n341) );
  XNOR2_X1 U337 ( .A(b[6]), .B(n283), .ZN(n340) );
  OAI22_X1 U338 ( .A1(n321), .A2(n315), .B1(n281), .B2(n323), .ZN(n21) );
  XNOR2_X1 U339 ( .A(b[7]), .B(a[5]), .ZN(n323) );
  XNOR2_X1 U340 ( .A(n291), .B(a[4]), .ZN(n342) );
  XNOR2_X1 U341 ( .A(b[6]), .B(a[5]), .ZN(n321) );
  OAI22_X1 U342 ( .A1(n332), .A2(n326), .B1(n324), .B2(n334), .ZN(n15) );
  XNOR2_X1 U343 ( .A(b[7]), .B(a[7]), .ZN(n334) );
  NAND2_X1 U344 ( .A1(n324), .A2(n343), .ZN(n326) );
  XNOR2_X1 U345 ( .A(n288), .B(a[6]), .ZN(n343) );
  XNOR2_X1 U346 ( .A(b[6]), .B(a[7]), .ZN(n332) );
  OAI22_X1 U347 ( .A1(n284), .A2(n299), .B1(n344), .B2(n297), .ZN(n104) );
  OAI22_X1 U348 ( .A1(n236), .A2(n299), .B1(n345), .B2(n297), .ZN(n103) );
  XNOR2_X1 U349 ( .A(b[1]), .B(a[1]), .ZN(n344) );
  OAI22_X1 U350 ( .A1(n345), .A2(n299), .B1(n346), .B2(n297), .ZN(n102) );
  XNOR2_X1 U351 ( .A(b[2]), .B(a[1]), .ZN(n345) );
  OAI22_X1 U352 ( .A1(n346), .A2(n299), .B1(n347), .B2(n297), .ZN(n101) );
  XNOR2_X1 U353 ( .A(b[3]), .B(a[1]), .ZN(n346) );
  OAI22_X1 U354 ( .A1(n347), .A2(n299), .B1(n298), .B2(n297), .ZN(n100) );
  XNOR2_X1 U355 ( .A(b[5]), .B(a[1]), .ZN(n298) );
  NAND2_X1 U356 ( .A1(a[1]), .A2(n297), .ZN(n299) );
  XNOR2_X1 U357 ( .A(b[4]), .B(a[1]), .ZN(n347) );
endmodule


module datapath_DW01_add_21 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n65;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n65), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND3_X1 U1 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n1) );
  NAND3_X1 U2 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n2) );
  NAND3_X1 U3 ( .A1(n8), .A2(n9), .A3(n10), .ZN(n3) );
  CLKBUF_X1 U4 ( .A(B[6]), .Z(n4) );
  CLKBUF_X1 U5 ( .A(n1), .Z(n5) );
  NAND3_X1 U6 ( .A1(n62), .A2(n61), .A3(n63), .ZN(n6) );
  XOR2_X1 U7 ( .A(B[5]), .B(A[5]), .Z(n7) );
  XOR2_X1 U8 ( .A(n5), .B(n7), .Z(SUM[5]) );
  NAND2_X1 U9 ( .A1(n1), .A2(B[5]), .ZN(n8) );
  NAND2_X1 U10 ( .A1(carry[5]), .A2(A[5]), .ZN(n9) );
  NAND2_X1 U11 ( .A1(B[5]), .A2(A[5]), .ZN(n10) );
  NAND3_X1 U12 ( .A1(n8), .A2(n9), .A3(n10), .ZN(carry[6]) );
  CLKBUF_X1 U13 ( .A(carry[4]), .Z(n11) );
  CLKBUF_X1 U14 ( .A(n2), .Z(n12) );
  XOR2_X1 U15 ( .A(B[10]), .B(A[10]), .Z(n13) );
  XOR2_X1 U16 ( .A(n6), .B(n13), .Z(SUM[10]) );
  NAND2_X1 U17 ( .A1(n6), .A2(B[10]), .ZN(n14) );
  NAND2_X1 U18 ( .A1(carry[10]), .A2(A[10]), .ZN(n15) );
  NAND2_X1 U19 ( .A1(B[10]), .A2(A[10]), .ZN(n16) );
  NAND3_X1 U20 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[11]) );
  NAND3_X1 U21 ( .A1(n21), .A2(n20), .A3(n22), .ZN(n17) );
  CLKBUF_X1 U22 ( .A(n25), .Z(n18) );
  XOR2_X1 U23 ( .A(B[11]), .B(A[11]), .Z(n19) );
  XOR2_X1 U24 ( .A(n12), .B(n19), .Z(SUM[11]) );
  NAND2_X1 U25 ( .A1(n2), .A2(B[11]), .ZN(n20) );
  NAND2_X1 U26 ( .A1(carry[11]), .A2(A[11]), .ZN(n21) );
  NAND2_X1 U27 ( .A1(B[11]), .A2(A[11]), .ZN(n22) );
  NAND3_X1 U28 ( .A1(n20), .A2(n21), .A3(n22), .ZN(carry[12]) );
  CLKBUF_X1 U29 ( .A(carry[6]), .Z(n23) );
  CLKBUF_X1 U30 ( .A(n53), .Z(n24) );
  NAND3_X1 U31 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n25) );
  NAND3_X1 U32 ( .A1(n40), .A2(n42), .A3(n41), .ZN(n26) );
  CLKBUF_X1 U33 ( .A(n55), .Z(n27) );
  XOR2_X1 U34 ( .A(B[12]), .B(A[12]), .Z(n28) );
  XOR2_X1 U35 ( .A(carry[12]), .B(n28), .Z(SUM[12]) );
  NAND2_X1 U36 ( .A1(n17), .A2(B[12]), .ZN(n29) );
  NAND2_X1 U37 ( .A1(carry[12]), .A2(A[12]), .ZN(n30) );
  NAND2_X1 U38 ( .A1(B[12]), .A2(A[12]), .ZN(n31) );
  NAND3_X1 U39 ( .A1(n29), .A2(n30), .A3(n31), .ZN(carry[13]) );
  NAND3_X1 U40 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n32) );
  NAND3_X1 U41 ( .A1(n52), .A2(n24), .A3(n54), .ZN(n33) );
  XNOR2_X1 U42 ( .A(carry[15]), .B(n34), .ZN(SUM[15]) );
  XNOR2_X1 U43 ( .A(B[15]), .B(A[15]), .ZN(n34) );
  XOR2_X1 U44 ( .A(B[13]), .B(A[13]), .Z(n35) );
  XOR2_X1 U45 ( .A(n18), .B(n35), .Z(SUM[13]) );
  NAND2_X1 U46 ( .A1(n25), .A2(B[13]), .ZN(n36) );
  NAND2_X1 U47 ( .A1(carry[13]), .A2(A[13]), .ZN(n37) );
  NAND2_X1 U48 ( .A1(B[13]), .A2(A[13]), .ZN(n38) );
  NAND3_X1 U49 ( .A1(n36), .A2(n37), .A3(n38), .ZN(carry[14]) );
  XOR2_X1 U50 ( .A(n23), .B(A[6]), .Z(n39) );
  XOR2_X1 U51 ( .A(n4), .B(n39), .Z(SUM[6]) );
  NAND2_X1 U52 ( .A1(B[6]), .A2(n3), .ZN(n40) );
  NAND2_X1 U53 ( .A1(B[6]), .A2(A[6]), .ZN(n41) );
  NAND2_X1 U54 ( .A1(carry[6]), .A2(A[6]), .ZN(n42) );
  NAND3_X1 U55 ( .A1(n40), .A2(n42), .A3(n41), .ZN(carry[7]) );
  XOR2_X1 U56 ( .A(B[3]), .B(A[3]), .Z(n43) );
  XOR2_X1 U57 ( .A(carry[3]), .B(n43), .Z(SUM[3]) );
  NAND2_X1 U58 ( .A1(carry[3]), .A2(B[3]), .ZN(n44) );
  NAND2_X1 U59 ( .A1(carry[3]), .A2(A[3]), .ZN(n45) );
  NAND2_X1 U60 ( .A1(B[3]), .A2(A[3]), .ZN(n46) );
  NAND3_X1 U61 ( .A1(n44), .A2(n45), .A3(n46), .ZN(carry[4]) );
  XOR2_X1 U62 ( .A(B[4]), .B(A[4]), .Z(n47) );
  XOR2_X1 U63 ( .A(n11), .B(n47), .Z(SUM[4]) );
  NAND2_X1 U64 ( .A1(carry[4]), .A2(B[4]), .ZN(n48) );
  NAND2_X1 U65 ( .A1(carry[4]), .A2(A[4]), .ZN(n49) );
  NAND2_X1 U66 ( .A1(B[4]), .A2(A[4]), .ZN(n50) );
  NAND3_X1 U67 ( .A1(n48), .A2(n49), .A3(n50), .ZN(carry[5]) );
  XOR2_X1 U68 ( .A(B[7]), .B(A[7]), .Z(n51) );
  XOR2_X1 U69 ( .A(n26), .B(n51), .Z(SUM[7]) );
  NAND2_X1 U70 ( .A1(carry[7]), .A2(B[7]), .ZN(n52) );
  NAND2_X1 U71 ( .A1(carry[7]), .A2(A[7]), .ZN(n53) );
  NAND2_X1 U72 ( .A1(B[7]), .A2(A[7]), .ZN(n54) );
  NAND3_X1 U73 ( .A1(n52), .A2(n53), .A3(n54), .ZN(carry[8]) );
  NAND3_X1 U74 ( .A1(n59), .A2(n58), .A3(n57), .ZN(n55) );
  XOR2_X1 U75 ( .A(A[8]), .B(B[8]), .Z(n56) );
  XOR2_X1 U76 ( .A(n56), .B(n33), .Z(SUM[8]) );
  NAND2_X1 U77 ( .A1(A[8]), .A2(B[8]), .ZN(n57) );
  NAND2_X1 U78 ( .A1(A[8]), .A2(carry[8]), .ZN(n58) );
  NAND2_X1 U79 ( .A1(B[8]), .A2(n32), .ZN(n59) );
  NAND3_X1 U80 ( .A1(n58), .A2(n59), .A3(n57), .ZN(carry[9]) );
  XOR2_X1 U81 ( .A(A[9]), .B(B[9]), .Z(n60) );
  XOR2_X1 U82 ( .A(n60), .B(n27), .Z(SUM[9]) );
  NAND2_X1 U83 ( .A1(A[9]), .A2(B[9]), .ZN(n61) );
  NAND2_X1 U84 ( .A1(n55), .A2(A[9]), .ZN(n62) );
  NAND2_X1 U85 ( .A1(B[9]), .A2(carry[9]), .ZN(n63) );
  NAND3_X1 U86 ( .A1(n62), .A2(n61), .A3(n63), .ZN(carry[10]) );
  XOR2_X1 U87 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U88 ( .A1(B[0]), .A2(A[0]), .ZN(n65) );
endmodule


module datapath_DW_mult_tc_20 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74,
         n75, n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92,
         n93, n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330;

  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n274), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n273), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n277), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n276), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n279), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  NAND2_X1 U157 ( .A1(n296), .A2(n325), .ZN(n298) );
  INV_X1 U158 ( .A(n15), .ZN(n270) );
  INV_X1 U159 ( .A(n269), .ZN(n268) );
  XNOR2_X1 U160 ( .A(n271), .B(n15), .ZN(n206) );
  AND3_X1 U161 ( .A1(n262), .A2(n263), .A3(n264), .ZN(product[15]) );
  NAND3_X1 U162 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n208) );
  NAND3_X1 U163 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n209) );
  XNOR2_X1 U164 ( .A(n2), .B(n206), .ZN(product[14]) );
  BUF_X2 U165 ( .A(n296), .Z(n210) );
  XNOR2_X1 U166 ( .A(a[4]), .B(a[3]), .ZN(n296) );
  XOR2_X2 U167 ( .A(a[6]), .B(n275), .Z(n307) );
  XOR2_X1 U168 ( .A(n18), .B(n19), .Z(n211) );
  XOR2_X1 U169 ( .A(n209), .B(n211), .Z(product[12]) );
  NAND2_X1 U170 ( .A1(n208), .A2(n18), .ZN(n212) );
  NAND2_X1 U171 ( .A1(n4), .A2(n19), .ZN(n213) );
  NAND2_X1 U172 ( .A1(n18), .A2(n19), .ZN(n214) );
  NAND3_X1 U173 ( .A1(n212), .A2(n213), .A3(n214), .ZN(n3) );
  NAND3_X1 U174 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n215) );
  NAND3_X1 U175 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n216) );
  NAND3_X1 U176 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n217) );
  NAND3_X1 U177 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n218) );
  NAND3_X1 U178 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n219) );
  NAND3_X1 U179 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n220) );
  NAND3_X1 U180 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n221) );
  NAND3_X1 U181 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n222) );
  CLKBUF_X1 U182 ( .A(n327), .Z(n235) );
  XOR2_X1 U183 ( .A(n17), .B(n270), .Z(n223) );
  XOR2_X1 U184 ( .A(n3), .B(n223), .Z(product[13]) );
  NAND2_X1 U185 ( .A1(n3), .A2(n17), .ZN(n224) );
  NAND2_X1 U186 ( .A1(n3), .A2(n270), .ZN(n225) );
  NAND2_X1 U187 ( .A1(n17), .A2(n270), .ZN(n226) );
  NAND3_X1 U188 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n2) );
  XOR2_X1 U189 ( .A(n50), .B(n53), .Z(n227) );
  XOR2_X1 U190 ( .A(n220), .B(n227), .Z(product[5]) );
  NAND2_X1 U191 ( .A1(n220), .A2(n50), .ZN(n228) );
  NAND2_X1 U192 ( .A1(n11), .A2(n53), .ZN(n229) );
  NAND2_X1 U193 ( .A1(n50), .A2(n53), .ZN(n230) );
  NAND3_X1 U194 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n10) );
  XOR2_X1 U195 ( .A(n33), .B(n28), .Z(n231) );
  XOR2_X1 U196 ( .A(n7), .B(n231), .Z(product[9]) );
  NAND2_X1 U197 ( .A1(n7), .A2(n33), .ZN(n232) );
  NAND2_X1 U198 ( .A1(n7), .A2(n28), .ZN(n233) );
  NAND2_X1 U199 ( .A1(n33), .A2(n28), .ZN(n234) );
  NAND3_X1 U200 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n6) );
  NAND3_X1 U201 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n236) );
  XOR2_X1 U202 ( .A(n27), .B(n24), .Z(n237) );
  XOR2_X1 U203 ( .A(n218), .B(n237), .Z(product[10]) );
  NAND2_X1 U204 ( .A1(n218), .A2(n27), .ZN(n238) );
  NAND2_X1 U205 ( .A1(n6), .A2(n24), .ZN(n239) );
  NAND2_X1 U206 ( .A1(n27), .A2(n24), .ZN(n240) );
  NAND3_X1 U207 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n5) );
  XOR2_X1 U208 ( .A(n40), .B(n45), .Z(n241) );
  XOR2_X1 U209 ( .A(n217), .B(n241), .Z(product[7]) );
  NAND2_X1 U210 ( .A1(n217), .A2(n40), .ZN(n242) );
  NAND2_X1 U211 ( .A1(n9), .A2(n45), .ZN(n243) );
  NAND2_X1 U212 ( .A1(n40), .A2(n45), .ZN(n244) );
  NAND3_X1 U213 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n8) );
  CLKBUF_X1 U214 ( .A(b[1]), .Z(n245) );
  XOR2_X1 U215 ( .A(n54), .B(n55), .Z(n246) );
  XOR2_X1 U216 ( .A(n246), .B(n12), .Z(product[4]) );
  NAND2_X1 U217 ( .A1(n12), .A2(n54), .ZN(n247) );
  NAND2_X1 U218 ( .A1(n12), .A2(n55), .ZN(n248) );
  NAND2_X1 U219 ( .A1(n54), .A2(n55), .ZN(n249) );
  NAND3_X1 U220 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n11) );
  XOR2_X1 U221 ( .A(n46), .B(n49), .Z(n250) );
  XOR2_X1 U222 ( .A(n216), .B(n250), .Z(product[6]) );
  NAND2_X1 U223 ( .A1(n215), .A2(n46), .ZN(n251) );
  NAND2_X1 U224 ( .A1(n10), .A2(n49), .ZN(n252) );
  NAND2_X1 U225 ( .A1(n46), .A2(n49), .ZN(n253) );
  NAND3_X1 U226 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n9) );
  XOR2_X1 U227 ( .A(n34), .B(n39), .Z(n254) );
  XOR2_X1 U228 ( .A(n222), .B(n254), .Z(product[8]) );
  NAND2_X1 U229 ( .A1(n221), .A2(n34), .ZN(n255) );
  NAND2_X1 U230 ( .A1(n8), .A2(n39), .ZN(n256) );
  NAND2_X1 U231 ( .A1(n34), .A2(n39), .ZN(n257) );
  NAND3_X1 U232 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n7) );
  XOR2_X1 U233 ( .A(n23), .B(n20), .Z(n258) );
  XOR2_X1 U234 ( .A(n236), .B(n258), .Z(product[11]) );
  NAND2_X1 U235 ( .A1(n236), .A2(n23), .ZN(n259) );
  NAND2_X1 U236 ( .A1(n5), .A2(n20), .ZN(n260) );
  NAND2_X1 U237 ( .A1(n23), .A2(n20), .ZN(n261) );
  NAND3_X1 U238 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n4) );
  NAND2_X1 U239 ( .A1(n219), .A2(n271), .ZN(n262) );
  NAND2_X1 U240 ( .A1(n219), .A2(n15), .ZN(n263) );
  NAND2_X1 U241 ( .A1(n271), .A2(n15), .ZN(n264) );
  CLKBUF_X1 U242 ( .A(n286), .Z(n265) );
  XOR2_X1 U243 ( .A(a[2]), .B(n266), .Z(n286) );
  INV_X1 U244 ( .A(n21), .ZN(n273) );
  INV_X1 U245 ( .A(n305), .ZN(n274) );
  INV_X1 U246 ( .A(n316), .ZN(n271) );
  INV_X1 U247 ( .A(n285), .ZN(n279) );
  INV_X1 U248 ( .A(n294), .ZN(n277) );
  INV_X1 U249 ( .A(n31), .ZN(n276) );
  INV_X1 U250 ( .A(b[0]), .ZN(n269) );
  NAND2_X1 U251 ( .A1(n286), .A2(n324), .ZN(n288) );
  INV_X1 U252 ( .A(n266), .ZN(n267) );
  INV_X1 U253 ( .A(a[0]), .ZN(n280) );
  INV_X1 U254 ( .A(a[5]), .ZN(n275) );
  INV_X1 U255 ( .A(a[7]), .ZN(n272) );
  INV_X1 U256 ( .A(a[3]), .ZN(n278) );
  INV_X1 U257 ( .A(a[1]), .ZN(n266) );
  NOR2_X1 U258 ( .A1(n280), .A2(n269), .ZN(product[0]) );
  OAI22_X1 U259 ( .A1(n281), .A2(n282), .B1(n283), .B2(n280), .ZN(n99) );
  OAI22_X1 U260 ( .A1(n283), .A2(n282), .B1(n284), .B2(n280), .ZN(n98) );
  XNOR2_X1 U261 ( .A(b[6]), .B(n267), .ZN(n283) );
  OAI22_X1 U262 ( .A1(n280), .A2(n284), .B1(n282), .B2(n284), .ZN(n285) );
  XNOR2_X1 U263 ( .A(b[7]), .B(n267), .ZN(n284) );
  NOR2_X1 U264 ( .A1(n286), .A2(n269), .ZN(n96) );
  OAI22_X1 U265 ( .A1(n287), .A2(n288), .B1(n286), .B2(n289), .ZN(n95) );
  XNOR2_X1 U266 ( .A(a[3]), .B(n268), .ZN(n287) );
  OAI22_X1 U267 ( .A1(n289), .A2(n288), .B1(n265), .B2(n290), .ZN(n94) );
  XNOR2_X1 U268 ( .A(b[1]), .B(a[3]), .ZN(n289) );
  OAI22_X1 U269 ( .A1(n290), .A2(n288), .B1(n265), .B2(n291), .ZN(n93) );
  XNOR2_X1 U270 ( .A(b[2]), .B(a[3]), .ZN(n290) );
  OAI22_X1 U271 ( .A1(n291), .A2(n288), .B1(n265), .B2(n292), .ZN(n92) );
  XNOR2_X1 U272 ( .A(b[3]), .B(a[3]), .ZN(n291) );
  OAI22_X1 U273 ( .A1(n292), .A2(n288), .B1(n265), .B2(n293), .ZN(n91) );
  XNOR2_X1 U274 ( .A(b[4]), .B(a[3]), .ZN(n292) );
  OAI22_X1 U275 ( .A1(n295), .A2(n265), .B1(n288), .B2(n295), .ZN(n294) );
  NOR2_X1 U276 ( .A1(n210), .A2(n269), .ZN(n88) );
  OAI22_X1 U277 ( .A1(n297), .A2(n298), .B1(n210), .B2(n299), .ZN(n87) );
  XNOR2_X1 U278 ( .A(a[5]), .B(n268), .ZN(n297) );
  OAI22_X1 U279 ( .A1(n299), .A2(n298), .B1(n210), .B2(n300), .ZN(n86) );
  XNOR2_X1 U280 ( .A(n245), .B(a[5]), .ZN(n299) );
  OAI22_X1 U281 ( .A1(n300), .A2(n298), .B1(n210), .B2(n301), .ZN(n85) );
  XNOR2_X1 U282 ( .A(b[2]), .B(a[5]), .ZN(n300) );
  OAI22_X1 U283 ( .A1(n301), .A2(n298), .B1(n210), .B2(n302), .ZN(n84) );
  XNOR2_X1 U284 ( .A(b[3]), .B(a[5]), .ZN(n301) );
  OAI22_X1 U285 ( .A1(n302), .A2(n298), .B1(n210), .B2(n303), .ZN(n83) );
  XNOR2_X1 U286 ( .A(b[4]), .B(a[5]), .ZN(n302) );
  OAI22_X1 U287 ( .A1(n303), .A2(n298), .B1(n210), .B2(n304), .ZN(n82) );
  XNOR2_X1 U288 ( .A(b[5]), .B(a[5]), .ZN(n303) );
  OAI22_X1 U289 ( .A1(n306), .A2(n210), .B1(n298), .B2(n306), .ZN(n305) );
  NOR2_X1 U290 ( .A1(n307), .A2(n269), .ZN(n80) );
  OAI22_X1 U291 ( .A1(n308), .A2(n309), .B1(n307), .B2(n310), .ZN(n79) );
  XNOR2_X1 U292 ( .A(a[7]), .B(n268), .ZN(n308) );
  OAI22_X1 U293 ( .A1(n311), .A2(n309), .B1(n307), .B2(n312), .ZN(n77) );
  OAI22_X1 U294 ( .A1(n312), .A2(n309), .B1(n307), .B2(n313), .ZN(n76) );
  XNOR2_X1 U295 ( .A(b[3]), .B(a[7]), .ZN(n312) );
  OAI22_X1 U296 ( .A1(n313), .A2(n309), .B1(n307), .B2(n314), .ZN(n75) );
  XNOR2_X1 U297 ( .A(b[4]), .B(a[7]), .ZN(n313) );
  OAI22_X1 U298 ( .A1(n314), .A2(n309), .B1(n307), .B2(n315), .ZN(n74) );
  XNOR2_X1 U299 ( .A(b[5]), .B(a[7]), .ZN(n314) );
  OAI22_X1 U300 ( .A1(n317), .A2(n307), .B1(n309), .B2(n317), .ZN(n316) );
  OAI21_X1 U301 ( .B1(n268), .B2(n266), .A(n282), .ZN(n72) );
  OAI21_X1 U302 ( .B1(n278), .B2(n288), .A(n318), .ZN(n71) );
  OR3_X1 U303 ( .A1(n286), .A2(n268), .A3(n278), .ZN(n318) );
  OAI21_X1 U304 ( .B1(n275), .B2(n298), .A(n319), .ZN(n70) );
  OR3_X1 U305 ( .A1(n210), .A2(n268), .A3(n275), .ZN(n319) );
  OAI21_X1 U306 ( .B1(n272), .B2(n309), .A(n320), .ZN(n69) );
  OR3_X1 U307 ( .A1(n307), .A2(n268), .A3(n272), .ZN(n320) );
  XNOR2_X1 U308 ( .A(n321), .B(n322), .ZN(n38) );
  OR2_X1 U309 ( .A1(n321), .A2(n322), .ZN(n37) );
  OAI22_X1 U310 ( .A1(n293), .A2(n288), .B1(n265), .B2(n323), .ZN(n322) );
  XNOR2_X1 U311 ( .A(b[5]), .B(a[3]), .ZN(n293) );
  OAI22_X1 U312 ( .A1(n310), .A2(n309), .B1(n307), .B2(n311), .ZN(n321) );
  XNOR2_X1 U313 ( .A(b[2]), .B(a[7]), .ZN(n311) );
  XNOR2_X1 U314 ( .A(n245), .B(a[7]), .ZN(n310) );
  OAI22_X1 U315 ( .A1(n323), .A2(n288), .B1(n265), .B2(n295), .ZN(n31) );
  XNOR2_X1 U316 ( .A(b[7]), .B(a[3]), .ZN(n295) );
  XNOR2_X1 U317 ( .A(n278), .B(a[2]), .ZN(n324) );
  XNOR2_X1 U318 ( .A(b[6]), .B(a[3]), .ZN(n323) );
  OAI22_X1 U319 ( .A1(n304), .A2(n298), .B1(n210), .B2(n306), .ZN(n21) );
  XNOR2_X1 U320 ( .A(b[7]), .B(a[5]), .ZN(n306) );
  XNOR2_X1 U321 ( .A(n275), .B(a[4]), .ZN(n325) );
  XNOR2_X1 U322 ( .A(b[6]), .B(a[5]), .ZN(n304) );
  OAI22_X1 U323 ( .A1(n315), .A2(n309), .B1(n307), .B2(n317), .ZN(n15) );
  XNOR2_X1 U324 ( .A(b[7]), .B(a[7]), .ZN(n317) );
  NAND2_X1 U325 ( .A1(n307), .A2(n326), .ZN(n309) );
  XNOR2_X1 U326 ( .A(n272), .B(a[6]), .ZN(n326) );
  XNOR2_X1 U327 ( .A(b[6]), .B(a[7]), .ZN(n315) );
  OAI22_X1 U328 ( .A1(n268), .A2(n282), .B1(n327), .B2(n280), .ZN(n104) );
  OAI22_X1 U329 ( .A1(n235), .A2(n282), .B1(n328), .B2(n280), .ZN(n103) );
  XNOR2_X1 U330 ( .A(b[1]), .B(n267), .ZN(n327) );
  OAI22_X1 U331 ( .A1(n328), .A2(n282), .B1(n329), .B2(n280), .ZN(n102) );
  XNOR2_X1 U332 ( .A(b[2]), .B(n267), .ZN(n328) );
  OAI22_X1 U333 ( .A1(n329), .A2(n282), .B1(n330), .B2(n280), .ZN(n101) );
  XNOR2_X1 U334 ( .A(b[3]), .B(n267), .ZN(n329) );
  OAI22_X1 U335 ( .A1(n330), .A2(n282), .B1(n281), .B2(n280), .ZN(n100) );
  XNOR2_X1 U336 ( .A(b[5]), .B(n267), .ZN(n281) );
  NAND2_X1 U337 ( .A1(a[1]), .A2(n280), .ZN(n282) );
  XNOR2_X1 U338 ( .A(b[4]), .B(n267), .ZN(n330) );
endmodule


module datapath_DW01_add_20 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n77;
  wire   [15:1] carry;

  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n77), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(B[13]), .Z(n1) );
  CLKBUF_X1 U2 ( .A(n42), .Z(n2) );
  NAND3_X1 U3 ( .A1(n61), .A2(n60), .A3(n62), .ZN(n3) );
  NAND3_X1 U4 ( .A1(n61), .A2(n60), .A3(n62), .ZN(n4) );
  NAND3_X1 U5 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n5) );
  CLKBUF_X1 U6 ( .A(n70), .Z(n6) );
  CLKBUF_X1 U7 ( .A(n13), .Z(n7) );
  NAND3_X1 U8 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n8) );
  XOR2_X1 U9 ( .A(carry[2]), .B(A[2]), .Z(n9) );
  XOR2_X1 U10 ( .A(B[2]), .B(n9), .Z(SUM[2]) );
  NAND2_X1 U11 ( .A1(B[2]), .A2(carry[2]), .ZN(n10) );
  NAND2_X1 U12 ( .A1(B[2]), .A2(A[2]), .ZN(n11) );
  NAND2_X1 U13 ( .A1(carry[2]), .A2(A[2]), .ZN(n12) );
  NAND3_X1 U14 ( .A1(n10), .A2(n11), .A3(n12), .ZN(carry[3]) );
  NAND3_X1 U15 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n13) );
  CLKBUF_X1 U16 ( .A(n28), .Z(n14) );
  CLKBUF_X1 U17 ( .A(n32), .Z(n15) );
  XOR2_X1 U18 ( .A(B[8]), .B(A[8]), .Z(n16) );
  XOR2_X1 U19 ( .A(n4), .B(n16), .Z(SUM[8]) );
  NAND2_X1 U20 ( .A1(n3), .A2(B[8]), .ZN(n17) );
  NAND2_X1 U21 ( .A1(carry[8]), .A2(A[8]), .ZN(n18) );
  NAND2_X1 U22 ( .A1(B[8]), .A2(A[8]), .ZN(n19) );
  NAND3_X1 U23 ( .A1(n17), .A2(n18), .A3(n19), .ZN(carry[9]) );
  NAND3_X1 U24 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n20) );
  NAND3_X1 U25 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n21) );
  XOR2_X1 U26 ( .A(B[11]), .B(A[11]), .Z(n22) );
  XOR2_X1 U27 ( .A(n21), .B(n22), .Z(SUM[11]) );
  NAND2_X1 U28 ( .A1(n20), .A2(B[11]), .ZN(n23) );
  NAND2_X1 U29 ( .A1(carry[11]), .A2(A[11]), .ZN(n24) );
  NAND2_X1 U30 ( .A1(B[11]), .A2(A[11]), .ZN(n25) );
  NAND3_X1 U31 ( .A1(n23), .A2(n24), .A3(n25), .ZN(carry[12]) );
  NAND3_X1 U32 ( .A1(n31), .A2(n32), .A3(n33), .ZN(n26) );
  NAND3_X1 U33 ( .A1(n31), .A2(n15), .A3(n33), .ZN(n27) );
  NAND3_X1 U34 ( .A1(n35), .A2(n37), .A3(n36), .ZN(n28) );
  XNOR2_X1 U35 ( .A(n2), .B(n29), .ZN(SUM[14]) );
  XNOR2_X1 U36 ( .A(B[14]), .B(A[14]), .ZN(n29) );
  XOR2_X1 U37 ( .A(B[9]), .B(A[9]), .Z(n30) );
  XOR2_X1 U38 ( .A(carry[9]), .B(n30), .Z(SUM[9]) );
  NAND2_X1 U39 ( .A1(n5), .A2(B[9]), .ZN(n31) );
  NAND2_X1 U40 ( .A1(carry[9]), .A2(A[9]), .ZN(n32) );
  NAND2_X1 U41 ( .A1(B[9]), .A2(A[9]), .ZN(n33) );
  NAND3_X1 U42 ( .A1(n31), .A2(n32), .A3(n33), .ZN(carry[10]) );
  XOR2_X1 U43 ( .A(B[5]), .B(A[5]), .Z(n34) );
  XOR2_X1 U44 ( .A(carry[5]), .B(n34), .Z(SUM[5]) );
  NAND2_X1 U45 ( .A1(carry[5]), .A2(B[5]), .ZN(n35) );
  NAND2_X1 U46 ( .A1(carry[5]), .A2(A[5]), .ZN(n36) );
  NAND2_X1 U47 ( .A1(B[5]), .A2(A[5]), .ZN(n37) );
  NAND3_X1 U48 ( .A1(n36), .A2(n35), .A3(n37), .ZN(carry[6]) );
  XNOR2_X1 U49 ( .A(n38), .B(carry[15]), .ZN(SUM[15]) );
  XNOR2_X1 U50 ( .A(B[15]), .B(A[15]), .ZN(n38) );
  CLKBUF_X1 U51 ( .A(carry[12]), .Z(n39) );
  NAND3_X1 U52 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n40) );
  NAND3_X1 U53 ( .A1(n74), .A2(n75), .A3(n73), .ZN(n41) );
  NAND3_X1 U54 ( .A1(n75), .A2(n74), .A3(n73), .ZN(n42) );
  NAND2_X1 U55 ( .A1(n42), .A2(B[14]), .ZN(n43) );
  NAND2_X1 U56 ( .A1(n41), .A2(A[14]), .ZN(n44) );
  NAND2_X1 U57 ( .A1(B[14]), .A2(A[14]), .ZN(n45) );
  NAND3_X1 U58 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[15]) );
  XOR2_X1 U59 ( .A(B[6]), .B(A[6]), .Z(n46) );
  XOR2_X1 U60 ( .A(n14), .B(n46), .Z(SUM[6]) );
  NAND2_X1 U61 ( .A1(n28), .A2(B[6]), .ZN(n47) );
  NAND2_X1 U62 ( .A1(carry[6]), .A2(A[6]), .ZN(n48) );
  NAND2_X1 U63 ( .A1(B[6]), .A2(A[6]), .ZN(n49) );
  CLKBUF_X1 U64 ( .A(carry[4]), .Z(n50) );
  XOR2_X1 U65 ( .A(B[3]), .B(A[3]), .Z(n51) );
  XOR2_X1 U66 ( .A(carry[3]), .B(n51), .Z(SUM[3]) );
  NAND2_X1 U67 ( .A1(carry[3]), .A2(B[3]), .ZN(n52) );
  NAND2_X1 U68 ( .A1(carry[3]), .A2(A[3]), .ZN(n53) );
  NAND2_X1 U69 ( .A1(B[3]), .A2(A[3]), .ZN(n54) );
  NAND3_X1 U70 ( .A1(n52), .A2(n53), .A3(n54), .ZN(carry[4]) );
  XOR2_X1 U71 ( .A(B[4]), .B(A[4]), .Z(n55) );
  XOR2_X1 U72 ( .A(n50), .B(n55), .Z(SUM[4]) );
  NAND2_X1 U73 ( .A1(n8), .A2(B[4]), .ZN(n56) );
  NAND2_X1 U74 ( .A1(carry[4]), .A2(A[4]), .ZN(n57) );
  NAND2_X1 U75 ( .A1(B[4]), .A2(A[4]), .ZN(n58) );
  NAND3_X1 U76 ( .A1(n56), .A2(n57), .A3(n58), .ZN(carry[5]) );
  XOR2_X1 U77 ( .A(B[7]), .B(A[7]), .Z(n59) );
  XOR2_X1 U78 ( .A(n7), .B(n59), .Z(SUM[7]) );
  NAND2_X1 U79 ( .A1(n40), .A2(B[7]), .ZN(n60) );
  NAND2_X1 U80 ( .A1(n13), .A2(A[7]), .ZN(n61) );
  NAND2_X1 U81 ( .A1(B[7]), .A2(A[7]), .ZN(n62) );
  NAND3_X1 U82 ( .A1(n61), .A2(n60), .A3(n62), .ZN(carry[8]) );
  XOR2_X1 U83 ( .A(B[10]), .B(A[10]), .Z(n63) );
  XOR2_X1 U84 ( .A(n27), .B(n63), .Z(SUM[10]) );
  NAND2_X1 U85 ( .A1(n26), .A2(B[10]), .ZN(n64) );
  NAND2_X1 U86 ( .A1(carry[10]), .A2(A[10]), .ZN(n65) );
  NAND2_X1 U87 ( .A1(B[10]), .A2(A[10]), .ZN(n66) );
  NAND3_X1 U88 ( .A1(n64), .A2(n65), .A3(n66), .ZN(carry[11]) );
  NAND3_X1 U89 ( .A1(n71), .A2(n70), .A3(n69), .ZN(n67) );
  XOR2_X1 U90 ( .A(A[12]), .B(B[12]), .Z(n68) );
  XOR2_X1 U91 ( .A(n68), .B(n39), .Z(SUM[12]) );
  NAND2_X1 U92 ( .A1(A[12]), .A2(B[12]), .ZN(n69) );
  NAND2_X1 U93 ( .A1(A[12]), .A2(carry[12]), .ZN(n70) );
  NAND2_X1 U94 ( .A1(B[12]), .A2(carry[12]), .ZN(n71) );
  NAND3_X1 U95 ( .A1(n69), .A2(n6), .A3(n71), .ZN(carry[13]) );
  XOR2_X1 U96 ( .A(A[13]), .B(n1), .Z(n72) );
  XOR2_X1 U97 ( .A(n72), .B(carry[13]), .Z(SUM[13]) );
  NAND2_X1 U98 ( .A1(A[13]), .A2(B[13]), .ZN(n73) );
  NAND2_X1 U99 ( .A1(n67), .A2(A[13]), .ZN(n74) );
  NAND2_X1 U100 ( .A1(B[13]), .A2(n67), .ZN(n75) );
  XOR2_X1 U101 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U102 ( .A1(B[0]), .A2(A[0]), .ZN(n77) );
endmodule


module datapath_DW_mult_tc_19 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336;

  FA_X1 U12 ( .A(n54), .B(n206), .CI(n12), .CO(n11), .S(product[4]) );
  FA_X1 U13 ( .A(n13), .B(n71), .CI(n56), .CO(n12), .S(product[3]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n279), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n278), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n282), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n281), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n284), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  INV_X1 U157 ( .A(n274), .ZN(n273) );
  BUF_X1 U158 ( .A(n274), .Z(n224) );
  INV_X1 U159 ( .A(n15), .ZN(n275) );
  AND2_X1 U160 ( .A1(n95), .A2(n102), .ZN(n206) );
  XNOR2_X1 U161 ( .A(n276), .B(n15), .ZN(n207) );
  AND3_X1 U162 ( .A1(n265), .A2(n266), .A3(n267), .ZN(product[15]) );
  CLKBUF_X1 U163 ( .A(n14), .Z(n209) );
  NAND3_X1 U164 ( .A1(n213), .A2(n214), .A3(n215), .ZN(n210) );
  XNOR2_X1 U165 ( .A(n11), .B(n211), .ZN(product[5]) );
  XNOR2_X1 U166 ( .A(n50), .B(n53), .ZN(n211) );
  XNOR2_X1 U167 ( .A(n2), .B(n207), .ZN(product[14]) );
  XOR2_X1 U168 ( .A(n17), .B(n275), .Z(n212) );
  XOR2_X1 U169 ( .A(n3), .B(n212), .Z(product[13]) );
  NAND2_X1 U170 ( .A1(n3), .A2(n17), .ZN(n213) );
  NAND2_X1 U171 ( .A1(n3), .A2(n275), .ZN(n214) );
  NAND2_X1 U172 ( .A1(n17), .A2(n275), .ZN(n215) );
  NAND3_X1 U173 ( .A1(n213), .A2(n214), .A3(n215), .ZN(n2) );
  XOR2_X1 U174 ( .A(n216), .B(n217), .Z(product[7]) );
  XNOR2_X1 U175 ( .A(n40), .B(n45), .ZN(n216) );
  AND3_X1 U176 ( .A1(n261), .A2(n260), .A3(n259), .ZN(n217) );
  NAND3_X1 U177 ( .A1(n219), .A2(n220), .A3(n221), .ZN(n218) );
  NAND2_X1 U178 ( .A1(n11), .A2(n50), .ZN(n219) );
  NAND2_X1 U179 ( .A1(n11), .A2(n53), .ZN(n220) );
  NAND2_X1 U180 ( .A1(n50), .A2(n53), .ZN(n221) );
  NAND3_X1 U181 ( .A1(n219), .A2(n220), .A3(n221), .ZN(n10) );
  NAND3_X1 U182 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n222) );
  NAND3_X1 U183 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n223) );
  XOR2_X1 U184 ( .A(n19), .B(n18), .Z(n225) );
  XOR2_X1 U185 ( .A(n223), .B(n225), .Z(product[12]) );
  NAND2_X1 U186 ( .A1(n222), .A2(n19), .ZN(n226) );
  NAND2_X1 U187 ( .A1(n4), .A2(n18), .ZN(n227) );
  NAND2_X1 U188 ( .A1(n19), .A2(n18), .ZN(n228) );
  NAND3_X1 U189 ( .A1(n226), .A2(n227), .A3(n228), .ZN(n3) );
  XNOR2_X1 U190 ( .A(n229), .B(n218), .ZN(product[6]) );
  XNOR2_X1 U191 ( .A(n46), .B(n49), .ZN(n229) );
  NAND3_X1 U192 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n230) );
  XOR2_X1 U193 ( .A(n231), .B(n232), .Z(product[10]) );
  XNOR2_X1 U194 ( .A(n24), .B(n27), .ZN(n231) );
  AND3_X1 U195 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n232) );
  NAND3_X1 U196 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n233) );
  NAND3_X1 U197 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n234) );
  NAND3_X1 U198 ( .A1(n239), .A2(n240), .A3(n238), .ZN(n235) );
  NAND3_X1 U199 ( .A1(n239), .A2(n238), .A3(n240), .ZN(n236) );
  XOR2_X1 U200 ( .A(n34), .B(n39), .Z(n237) );
  XOR2_X1 U201 ( .A(n230), .B(n237), .Z(product[8]) );
  NAND2_X1 U202 ( .A1(n8), .A2(n34), .ZN(n238) );
  NAND2_X1 U203 ( .A1(n8), .A2(n39), .ZN(n239) );
  NAND2_X1 U204 ( .A1(n34), .A2(n39), .ZN(n240) );
  NAND3_X1 U205 ( .A1(n238), .A2(n240), .A3(n239), .ZN(n7) );
  XOR2_X1 U206 ( .A(n23), .B(n20), .Z(n241) );
  XOR2_X1 U207 ( .A(n234), .B(n241), .Z(product[11]) );
  NAND2_X1 U208 ( .A1(n233), .A2(n23), .ZN(n242) );
  NAND2_X1 U209 ( .A1(n5), .A2(n20), .ZN(n243) );
  NAND2_X1 U210 ( .A1(n23), .A2(n20), .ZN(n244) );
  NAND3_X1 U211 ( .A1(n243), .A2(n242), .A3(n244), .ZN(n4) );
  NAND3_X1 U212 ( .A1(n255), .A2(n254), .A3(n253), .ZN(n245) );
  XOR2_X1 U213 ( .A(n103), .B(n96), .Z(n246) );
  XOR2_X1 U214 ( .A(n246), .B(n209), .Z(product[2]) );
  NAND2_X1 U215 ( .A1(n14), .A2(n103), .ZN(n247) );
  NAND2_X1 U216 ( .A1(n14), .A2(n96), .ZN(n248) );
  NAND2_X1 U217 ( .A1(n103), .A2(n96), .ZN(n249) );
  NAND3_X1 U218 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n13) );
  NAND3_X1 U219 ( .A1(n261), .A2(n259), .A3(n260), .ZN(n250) );
  XOR2_X1 U220 ( .A(n95), .B(n102), .Z(n56) );
  BUF_X1 U221 ( .A(n333), .Z(n251) );
  XOR2_X1 U222 ( .A(n28), .B(n33), .Z(n252) );
  XOR2_X1 U223 ( .A(n252), .B(n236), .Z(product[9]) );
  NAND2_X1 U224 ( .A1(n28), .A2(n33), .ZN(n253) );
  NAND2_X1 U225 ( .A1(n28), .A2(n7), .ZN(n254) );
  NAND2_X1 U226 ( .A1(n235), .A2(n33), .ZN(n255) );
  NAND3_X1 U227 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n6) );
  NAND2_X1 U228 ( .A1(n24), .A2(n27), .ZN(n256) );
  NAND2_X1 U229 ( .A1(n24), .A2(n245), .ZN(n257) );
  NAND2_X1 U230 ( .A1(n27), .A2(n6), .ZN(n258) );
  NAND3_X1 U231 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n5) );
  XNOR2_X2 U232 ( .A(a[4]), .B(a[3]), .ZN(n302) );
  CLKBUF_X1 U233 ( .A(n304), .Z(n272) );
  XOR2_X1 U234 ( .A(a[3]), .B(n274), .Z(n293) );
  NAND2_X1 U235 ( .A1(n46), .A2(n49), .ZN(n259) );
  NAND2_X1 U236 ( .A1(n46), .A2(n10), .ZN(n260) );
  NAND2_X1 U237 ( .A1(n49), .A2(n10), .ZN(n261) );
  NAND3_X1 U238 ( .A1(n260), .A2(n261), .A3(n259), .ZN(n9) );
  NAND2_X1 U239 ( .A1(n40), .A2(n45), .ZN(n262) );
  NAND2_X1 U240 ( .A1(n40), .A2(n250), .ZN(n263) );
  NAND2_X1 U241 ( .A1(n45), .A2(n9), .ZN(n264) );
  NAND3_X1 U242 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n8) );
  NAND2_X1 U243 ( .A1(n210), .A2(n276), .ZN(n265) );
  NAND2_X1 U244 ( .A1(n210), .A2(n15), .ZN(n266) );
  NAND2_X1 U245 ( .A1(n276), .A2(n15), .ZN(n267) );
  CLKBUF_X1 U246 ( .A(n294), .Z(n268) );
  NAND2_X2 U247 ( .A1(a[1]), .A2(n286), .ZN(n288) );
  NAND2_X1 U248 ( .A1(a[2]), .A2(a[1]), .ZN(n270) );
  NAND2_X1 U249 ( .A1(n269), .A2(n285), .ZN(n271) );
  NAND2_X2 U250 ( .A1(n270), .A2(n271), .ZN(n292) );
  INV_X1 U251 ( .A(a[2]), .ZN(n269) );
  NAND2_X1 U252 ( .A1(n302), .A2(n331), .ZN(n304) );
  INV_X1 U253 ( .A(n21), .ZN(n278) );
  INV_X1 U254 ( .A(n311), .ZN(n279) );
  INV_X1 U255 ( .A(n322), .ZN(n276) );
  INV_X1 U256 ( .A(n291), .ZN(n284) );
  INV_X1 U257 ( .A(n300), .ZN(n282) );
  INV_X1 U258 ( .A(n31), .ZN(n281) );
  INV_X1 U259 ( .A(b[0]), .ZN(n274) );
  INV_X1 U260 ( .A(a[5]), .ZN(n280) );
  INV_X1 U261 ( .A(a[7]), .ZN(n277) );
  INV_X1 U262 ( .A(a[3]), .ZN(n283) );
  NAND2_X2 U263 ( .A1(n292), .A2(n330), .ZN(n294) );
  INV_X1 U264 ( .A(a[1]), .ZN(n285) );
  XOR2_X2 U265 ( .A(a[6]), .B(n280), .Z(n313) );
  INV_X2 U266 ( .A(a[0]), .ZN(n286) );
  NOR2_X1 U267 ( .A1(n286), .A2(n224), .ZN(product[0]) );
  OAI22_X1 U268 ( .A1(n287), .A2(n288), .B1(n289), .B2(n286), .ZN(n99) );
  OAI22_X1 U269 ( .A1(n289), .A2(n288), .B1(n290), .B2(n286), .ZN(n98) );
  XNOR2_X1 U270 ( .A(b[6]), .B(a[1]), .ZN(n289) );
  OAI22_X1 U271 ( .A1(n286), .A2(n290), .B1(n288), .B2(n290), .ZN(n291) );
  XNOR2_X1 U272 ( .A(b[7]), .B(a[1]), .ZN(n290) );
  NOR2_X1 U273 ( .A1(n292), .A2(n224), .ZN(n96) );
  OAI22_X1 U274 ( .A1(n293), .A2(n294), .B1(n292), .B2(n295), .ZN(n95) );
  OAI22_X1 U275 ( .A1(n295), .A2(n294), .B1(n292), .B2(n296), .ZN(n94) );
  XNOR2_X1 U276 ( .A(b[1]), .B(a[3]), .ZN(n295) );
  OAI22_X1 U277 ( .A1(n296), .A2(n294), .B1(n292), .B2(n297), .ZN(n93) );
  XNOR2_X1 U278 ( .A(b[2]), .B(a[3]), .ZN(n296) );
  OAI22_X1 U279 ( .A1(n297), .A2(n294), .B1(n292), .B2(n298), .ZN(n92) );
  XNOR2_X1 U280 ( .A(b[3]), .B(a[3]), .ZN(n297) );
  OAI22_X1 U281 ( .A1(n298), .A2(n294), .B1(n292), .B2(n299), .ZN(n91) );
  XNOR2_X1 U282 ( .A(b[4]), .B(a[3]), .ZN(n298) );
  OAI22_X1 U283 ( .A1(n301), .A2(n292), .B1(n268), .B2(n301), .ZN(n300) );
  NOR2_X1 U284 ( .A1(n302), .A2(n224), .ZN(n88) );
  OAI22_X1 U285 ( .A1(n303), .A2(n304), .B1(n302), .B2(n305), .ZN(n87) );
  XNOR2_X1 U286 ( .A(a[5]), .B(n273), .ZN(n303) );
  OAI22_X1 U287 ( .A1(n305), .A2(n272), .B1(n302), .B2(n306), .ZN(n86) );
  XNOR2_X1 U288 ( .A(b[1]), .B(a[5]), .ZN(n305) );
  OAI22_X1 U289 ( .A1(n306), .A2(n304), .B1(n302), .B2(n307), .ZN(n85) );
  XNOR2_X1 U290 ( .A(b[2]), .B(a[5]), .ZN(n306) );
  OAI22_X1 U291 ( .A1(n307), .A2(n272), .B1(n302), .B2(n308), .ZN(n84) );
  XNOR2_X1 U292 ( .A(b[3]), .B(a[5]), .ZN(n307) );
  OAI22_X1 U293 ( .A1(n308), .A2(n272), .B1(n302), .B2(n309), .ZN(n83) );
  XNOR2_X1 U294 ( .A(b[4]), .B(a[5]), .ZN(n308) );
  OAI22_X1 U295 ( .A1(n309), .A2(n272), .B1(n302), .B2(n310), .ZN(n82) );
  XNOR2_X1 U296 ( .A(b[5]), .B(a[5]), .ZN(n309) );
  OAI22_X1 U297 ( .A1(n312), .A2(n302), .B1(n272), .B2(n312), .ZN(n311) );
  NOR2_X1 U298 ( .A1(n313), .A2(n224), .ZN(n80) );
  OAI22_X1 U299 ( .A1(n314), .A2(n315), .B1(n313), .B2(n316), .ZN(n79) );
  XNOR2_X1 U300 ( .A(a[7]), .B(n273), .ZN(n314) );
  OAI22_X1 U301 ( .A1(n317), .A2(n315), .B1(n313), .B2(n318), .ZN(n77) );
  OAI22_X1 U302 ( .A1(n318), .A2(n315), .B1(n313), .B2(n319), .ZN(n76) );
  XNOR2_X1 U303 ( .A(b[3]), .B(a[7]), .ZN(n318) );
  OAI22_X1 U304 ( .A1(n319), .A2(n315), .B1(n313), .B2(n320), .ZN(n75) );
  XNOR2_X1 U305 ( .A(b[4]), .B(a[7]), .ZN(n319) );
  OAI22_X1 U306 ( .A1(n320), .A2(n315), .B1(n313), .B2(n321), .ZN(n74) );
  XNOR2_X1 U307 ( .A(b[5]), .B(a[7]), .ZN(n320) );
  OAI22_X1 U308 ( .A1(n323), .A2(n313), .B1(n315), .B2(n323), .ZN(n322) );
  OAI21_X1 U309 ( .B1(n273), .B2(n285), .A(n288), .ZN(n72) );
  OAI21_X1 U310 ( .B1(n283), .B2(n294), .A(n324), .ZN(n71) );
  OR3_X1 U311 ( .A1(n292), .A2(n273), .A3(n283), .ZN(n324) );
  OAI21_X1 U312 ( .B1(n280), .B2(n304), .A(n325), .ZN(n70) );
  OR3_X1 U313 ( .A1(n302), .A2(n273), .A3(n280), .ZN(n325) );
  OAI21_X1 U314 ( .B1(n277), .B2(n315), .A(n326), .ZN(n69) );
  OR3_X1 U315 ( .A1(n313), .A2(n273), .A3(n277), .ZN(n326) );
  XNOR2_X1 U316 ( .A(n327), .B(n328), .ZN(n38) );
  OR2_X1 U317 ( .A1(n327), .A2(n328), .ZN(n37) );
  OAI22_X1 U318 ( .A1(n299), .A2(n268), .B1(n292), .B2(n329), .ZN(n328) );
  XNOR2_X1 U319 ( .A(b[5]), .B(a[3]), .ZN(n299) );
  OAI22_X1 U320 ( .A1(n316), .A2(n315), .B1(n313), .B2(n317), .ZN(n327) );
  XNOR2_X1 U321 ( .A(b[2]), .B(a[7]), .ZN(n317) );
  XNOR2_X1 U322 ( .A(b[1]), .B(a[7]), .ZN(n316) );
  OAI22_X1 U323 ( .A1(n329), .A2(n268), .B1(n292), .B2(n301), .ZN(n31) );
  XNOR2_X1 U324 ( .A(b[7]), .B(a[3]), .ZN(n301) );
  XNOR2_X1 U325 ( .A(n283), .B(a[2]), .ZN(n330) );
  XNOR2_X1 U326 ( .A(b[6]), .B(a[3]), .ZN(n329) );
  OAI22_X1 U327 ( .A1(n310), .A2(n272), .B1(n302), .B2(n312), .ZN(n21) );
  XNOR2_X1 U328 ( .A(b[7]), .B(a[5]), .ZN(n312) );
  XNOR2_X1 U329 ( .A(n280), .B(a[4]), .ZN(n331) );
  XNOR2_X1 U330 ( .A(b[6]), .B(a[5]), .ZN(n310) );
  OAI22_X1 U331 ( .A1(n321), .A2(n315), .B1(n313), .B2(n323), .ZN(n15) );
  XNOR2_X1 U332 ( .A(b[7]), .B(a[7]), .ZN(n323) );
  NAND2_X1 U333 ( .A1(n313), .A2(n332), .ZN(n315) );
  XNOR2_X1 U334 ( .A(n277), .B(a[6]), .ZN(n332) );
  XNOR2_X1 U335 ( .A(b[6]), .B(a[7]), .ZN(n321) );
  OAI22_X1 U336 ( .A1(n273), .A2(n288), .B1(n333), .B2(n286), .ZN(n104) );
  OAI22_X1 U337 ( .A1(n251), .A2(n288), .B1(n334), .B2(n286), .ZN(n103) );
  XNOR2_X1 U338 ( .A(b[1]), .B(a[1]), .ZN(n333) );
  OAI22_X1 U339 ( .A1(n334), .A2(n288), .B1(n335), .B2(n286), .ZN(n102) );
  XNOR2_X1 U340 ( .A(b[2]), .B(a[1]), .ZN(n334) );
  OAI22_X1 U341 ( .A1(n335), .A2(n288), .B1(n336), .B2(n286), .ZN(n101) );
  XNOR2_X1 U342 ( .A(b[3]), .B(a[1]), .ZN(n335) );
  OAI22_X1 U343 ( .A1(n336), .A2(n288), .B1(n287), .B2(n286), .ZN(n100) );
  XNOR2_X1 U344 ( .A(b[5]), .B(a[1]), .ZN(n287) );
  XNOR2_X1 U345 ( .A(b[4]), .B(a[1]), .ZN(n336) );
endmodule


module datapath_DW01_add_19 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n68;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n68), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(B[2]), .Z(n1) );
  CLKBUF_X1 U2 ( .A(carry[7]), .Z(n2) );
  NAND3_X1 U3 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n3) );
  NAND3_X1 U4 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n4) );
  CLKBUF_X1 U5 ( .A(n38), .Z(n5) );
  CLKBUF_X1 U6 ( .A(n40), .Z(n6) );
  CLKBUF_X1 U7 ( .A(B[3]), .Z(n7) );
  CLKBUF_X1 U8 ( .A(n15), .Z(n8) );
  CLKBUF_X1 U9 ( .A(n42), .Z(n9) );
  CLKBUF_X1 U10 ( .A(B[4]), .Z(n10) );
  XOR2_X1 U11 ( .A(n1), .B(A[2]), .Z(n11) );
  XOR2_X1 U12 ( .A(carry[2]), .B(n11), .Z(SUM[2]) );
  NAND2_X1 U13 ( .A1(carry[2]), .A2(B[2]), .ZN(n12) );
  NAND2_X1 U14 ( .A1(carry[2]), .A2(A[2]), .ZN(n13) );
  NAND2_X1 U15 ( .A1(B[2]), .A2(A[2]), .ZN(n14) );
  NAND3_X1 U16 ( .A1(n12), .A2(n13), .A3(n14), .ZN(carry[3]) );
  NAND3_X1 U17 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n15) );
  CLKBUF_X1 U18 ( .A(n49), .Z(n16) );
  CLKBUF_X1 U19 ( .A(n27), .Z(n17) );
  NAND3_X1 U20 ( .A1(n38), .A2(n40), .A3(n39), .ZN(n18) );
  NAND3_X1 U21 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n19) );
  NAND3_X1 U22 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n20) );
  NAND3_X1 U23 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n21) );
  NAND3_X1 U24 ( .A1(n9), .A2(n43), .A3(n44), .ZN(n22) );
  NAND3_X1 U25 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n23) );
  NAND3_X1 U26 ( .A1(n26), .A2(n17), .A3(n28), .ZN(n24) );
  XOR2_X1 U27 ( .A(n7), .B(A[3]), .Z(n25) );
  XOR2_X1 U28 ( .A(carry[3]), .B(n25), .Z(SUM[3]) );
  NAND2_X1 U29 ( .A1(carry[3]), .A2(B[3]), .ZN(n26) );
  NAND2_X1 U30 ( .A1(carry[3]), .A2(A[3]), .ZN(n27) );
  NAND2_X1 U31 ( .A1(B[3]), .A2(A[3]), .ZN(n28) );
  NAND3_X1 U32 ( .A1(n26), .A2(n27), .A3(n28), .ZN(carry[4]) );
  XOR2_X1 U33 ( .A(A[4]), .B(n10), .Z(n29) );
  XOR2_X1 U34 ( .A(n29), .B(n24), .Z(SUM[4]) );
  NAND2_X1 U35 ( .A1(A[4]), .A2(B[4]), .ZN(n30) );
  NAND2_X1 U36 ( .A1(A[4]), .A2(n23), .ZN(n31) );
  NAND2_X1 U37 ( .A1(B[4]), .A2(carry[4]), .ZN(n32) );
  NAND3_X1 U38 ( .A1(n30), .A2(n31), .A3(n32), .ZN(carry[5]) );
  XOR2_X1 U39 ( .A(A[5]), .B(B[5]), .Z(n33) );
  XOR2_X1 U40 ( .A(n33), .B(n20), .Z(SUM[5]) );
  NAND2_X1 U41 ( .A1(A[5]), .A2(B[5]), .ZN(n34) );
  NAND2_X1 U42 ( .A1(n19), .A2(A[5]), .ZN(n35) );
  NAND2_X1 U43 ( .A1(B[5]), .A2(carry[5]), .ZN(n36) );
  NAND3_X1 U44 ( .A1(n36), .A2(n35), .A3(n34), .ZN(carry[6]) );
  XOR2_X1 U45 ( .A(n22), .B(A[11]), .Z(n37) );
  XOR2_X1 U46 ( .A(B[11]), .B(n37), .Z(SUM[11]) );
  NAND2_X1 U47 ( .A1(B[11]), .A2(carry[11]), .ZN(n38) );
  NAND2_X1 U48 ( .A1(B[11]), .A2(A[11]), .ZN(n39) );
  NAND2_X1 U49 ( .A1(carry[11]), .A2(A[11]), .ZN(n40) );
  NAND3_X1 U50 ( .A1(n5), .A2(n6), .A3(n39), .ZN(carry[12]) );
  XOR2_X1 U51 ( .A(B[10]), .B(A[10]), .Z(n41) );
  XOR2_X1 U52 ( .A(n8), .B(n41), .Z(SUM[10]) );
  NAND2_X1 U53 ( .A1(B[10]), .A2(n15), .ZN(n42) );
  NAND2_X1 U54 ( .A1(carry[10]), .A2(A[10]), .ZN(n43) );
  NAND2_X1 U55 ( .A1(B[10]), .A2(A[10]), .ZN(n44) );
  NAND3_X1 U56 ( .A1(n42), .A2(n44), .A3(n43), .ZN(carry[11]) );
  XOR2_X1 U57 ( .A(B[7]), .B(A[7]), .Z(n45) );
  XOR2_X1 U58 ( .A(n2), .B(n45), .Z(SUM[7]) );
  NAND2_X1 U59 ( .A1(carry[7]), .A2(B[7]), .ZN(n46) );
  NAND2_X1 U60 ( .A1(carry[7]), .A2(A[7]), .ZN(n47) );
  NAND2_X1 U61 ( .A1(B[7]), .A2(A[7]), .ZN(n48) );
  NAND3_X1 U62 ( .A1(n46), .A2(n47), .A3(n48), .ZN(carry[8]) );
  NAND3_X1 U63 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n49) );
  XOR2_X1 U64 ( .A(B[12]), .B(A[12]), .Z(n50) );
  XOR2_X1 U65 ( .A(carry[12]), .B(n50), .Z(SUM[12]) );
  NAND2_X1 U66 ( .A1(n18), .A2(B[12]), .ZN(n51) );
  NAND2_X1 U67 ( .A1(n18), .A2(A[12]), .ZN(n52) );
  NAND2_X1 U68 ( .A1(B[12]), .A2(A[12]), .ZN(n53) );
  NAND3_X1 U69 ( .A1(n52), .A2(n51), .A3(n53), .ZN(carry[13]) );
  XOR2_X1 U70 ( .A(B[13]), .B(A[13]), .Z(n54) );
  XOR2_X1 U71 ( .A(n21), .B(n54), .Z(SUM[13]) );
  NAND2_X1 U72 ( .A1(B[13]), .A2(n21), .ZN(n55) );
  NAND2_X1 U73 ( .A1(carry[13]), .A2(A[13]), .ZN(n56) );
  NAND2_X1 U74 ( .A1(B[13]), .A2(A[13]), .ZN(n57) );
  NAND3_X1 U75 ( .A1(n55), .A2(n56), .A3(n57), .ZN(carry[14]) );
  XOR2_X1 U76 ( .A(B[9]), .B(A[9]), .Z(n58) );
  XOR2_X1 U77 ( .A(n16), .B(n58), .Z(SUM[9]) );
  NAND2_X1 U78 ( .A1(n49), .A2(B[9]), .ZN(n59) );
  NAND2_X1 U79 ( .A1(carry[9]), .A2(A[9]), .ZN(n60) );
  NAND2_X1 U80 ( .A1(B[9]), .A2(A[9]), .ZN(n61) );
  NAND3_X1 U81 ( .A1(n59), .A2(n60), .A3(n61), .ZN(carry[10]) );
  XNOR2_X1 U82 ( .A(carry[15]), .B(n62), .ZN(SUM[15]) );
  XNOR2_X1 U83 ( .A(B[15]), .B(A[15]), .ZN(n62) );
  XOR2_X1 U84 ( .A(B[8]), .B(A[8]), .Z(n63) );
  XOR2_X1 U85 ( .A(n4), .B(n63), .Z(SUM[8]) );
  NAND2_X1 U86 ( .A1(n3), .A2(B[8]), .ZN(n64) );
  NAND2_X1 U87 ( .A1(carry[8]), .A2(A[8]), .ZN(n65) );
  NAND2_X1 U88 ( .A1(B[8]), .A2(A[8]), .ZN(n66) );
  NAND3_X1 U89 ( .A1(n65), .A2(n64), .A3(n66), .ZN(carry[9]) );
  XOR2_X1 U90 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U91 ( .A1(B[0]), .A2(A[0]), .ZN(n68) );
endmodule


module datapath_DW_mult_tc_18 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n6, n7, n8, n9, n12, n13, n14, n15, n17, n18, n19, n20,
         n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75, n76, n77,
         n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94, n95,
         n96, n98, n99, n100, n101, n102, n103, n104, n206, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342;

  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n285), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n284), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n288), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n287), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n290), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n88), .B(n94), .CI(n101), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  XNOR2_X1 U157 ( .A(n282), .B(n15), .ZN(n206) );
  AND3_X1 U158 ( .A1(n217), .A2(n218), .A3(n219), .ZN(product[15]) );
  XNOR2_X1 U159 ( .A(n233), .B(n208), .ZN(product[7]) );
  XNOR2_X1 U160 ( .A(n40), .B(n45), .ZN(n208) );
  NAND3_X1 U161 ( .A1(n260), .A2(n259), .A3(n258), .ZN(n209) );
  NAND3_X1 U162 ( .A1(n260), .A2(n259), .A3(n258), .ZN(n210) );
  XOR2_X1 U163 ( .A(n34), .B(n39), .Z(n211) );
  XOR2_X1 U164 ( .A(n210), .B(n211), .Z(product[8]) );
  NAND2_X1 U165 ( .A1(n209), .A2(n34), .ZN(n212) );
  NAND2_X1 U166 ( .A1(n8), .A2(n39), .ZN(n213) );
  NAND2_X1 U167 ( .A1(n34), .A2(n39), .ZN(n214) );
  NAND3_X1 U168 ( .A1(n212), .A2(n213), .A3(n214), .ZN(n7) );
  XNOR2_X1 U169 ( .A(n2), .B(n206), .ZN(product[14]) );
  NAND2_X1 U170 ( .A1(n221), .A2(n27), .ZN(n215) );
  NAND3_X1 U171 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n216) );
  NAND2_X1 U172 ( .A1(n2), .A2(n282), .ZN(n217) );
  NAND2_X1 U173 ( .A1(n2), .A2(n15), .ZN(n218) );
  NAND2_X1 U174 ( .A1(n282), .A2(n15), .ZN(n219) );
  NAND3_X1 U175 ( .A1(n215), .A2(n247), .A3(n248), .ZN(n220) );
  NAND3_X1 U176 ( .A1(n236), .A2(n235), .A3(n237), .ZN(n221) );
  XOR2_X1 U177 ( .A(n222), .B(n223), .Z(product[11]) );
  XNOR2_X1 U178 ( .A(n20), .B(n23), .ZN(n222) );
  AND3_X1 U179 ( .A1(n215), .A2(n247), .A3(n248), .ZN(n223) );
  XOR2_X1 U180 ( .A(n17), .B(n281), .Z(n224) );
  XOR2_X1 U181 ( .A(n3), .B(n224), .Z(product[13]) );
  NAND2_X1 U182 ( .A1(n3), .A2(n17), .ZN(n225) );
  NAND2_X1 U183 ( .A1(n3), .A2(n281), .ZN(n226) );
  NAND2_X1 U184 ( .A1(n17), .A2(n281), .ZN(n227) );
  NAND3_X1 U185 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n2) );
  CLKBUF_X1 U186 ( .A(n14), .Z(n228) );
  CLKBUF_X1 U187 ( .A(n339), .Z(n269) );
  XNOR2_X1 U188 ( .A(n228), .B(n229), .ZN(product[2]) );
  XNOR2_X1 U189 ( .A(n103), .B(n96), .ZN(n229) );
  NAND3_X1 U190 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n230) );
  NAND3_X1 U191 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n231) );
  NAND3_X1 U192 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n232) );
  NAND3_X1 U193 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n233) );
  XOR2_X1 U194 ( .A(n33), .B(n28), .Z(n234) );
  XOR2_X1 U195 ( .A(n7), .B(n234), .Z(product[9]) );
  NAND2_X1 U196 ( .A1(n7), .A2(n33), .ZN(n235) );
  NAND2_X1 U197 ( .A1(n7), .A2(n28), .ZN(n236) );
  NAND2_X1 U198 ( .A1(n33), .A2(n28), .ZN(n237) );
  NAND3_X1 U199 ( .A1(n235), .A2(n236), .A3(n237), .ZN(n6) );
  NAND3_X1 U200 ( .A1(n267), .A2(n266), .A3(n268), .ZN(n238) );
  NAND3_X1 U201 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n239) );
  OAI22_X1 U202 ( .A1(n269), .A2(n294), .B1(n340), .B2(n292), .ZN(n240) );
  NAND2_X1 U203 ( .A1(a[4]), .A2(a[3]), .ZN(n243) );
  NAND2_X1 U204 ( .A1(n241), .A2(n242), .ZN(n244) );
  NAND2_X2 U205 ( .A1(n243), .A2(n244), .ZN(n308) );
  INV_X1 U206 ( .A(a[4]), .ZN(n241) );
  INV_X1 U207 ( .A(a[3]), .ZN(n242) );
  XOR2_X1 U208 ( .A(n27), .B(n24), .Z(n245) );
  XOR2_X1 U209 ( .A(n221), .B(n245), .Z(product[10]) );
  NAND2_X1 U210 ( .A1(n221), .A2(n27), .ZN(n246) );
  NAND2_X1 U211 ( .A1(n6), .A2(n24), .ZN(n247) );
  NAND2_X1 U212 ( .A1(n27), .A2(n24), .ZN(n248) );
  NAND3_X1 U213 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n249) );
  INV_X1 U214 ( .A(n280), .ZN(n250) );
  NAND2_X1 U215 ( .A1(n14), .A2(n240), .ZN(n251) );
  NAND2_X1 U216 ( .A1(n14), .A2(n96), .ZN(n252) );
  NAND2_X1 U217 ( .A1(n240), .A2(n96), .ZN(n253) );
  NAND3_X1 U218 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n13) );
  XOR2_X1 U219 ( .A(n46), .B(n49), .Z(n254) );
  XOR2_X1 U220 ( .A(n254), .B(n239), .Z(product[6]) );
  NAND2_X1 U221 ( .A1(n46), .A2(n49), .ZN(n255) );
  NAND2_X1 U222 ( .A1(n46), .A2(n238), .ZN(n256) );
  NAND2_X1 U223 ( .A1(n238), .A2(n49), .ZN(n257) );
  NAND3_X1 U224 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n9) );
  NAND2_X1 U225 ( .A1(n40), .A2(n45), .ZN(n258) );
  NAND2_X1 U226 ( .A1(n249), .A2(n40), .ZN(n259) );
  NAND2_X1 U227 ( .A1(n9), .A2(n45), .ZN(n260) );
  NAND3_X1 U228 ( .A1(n260), .A2(n259), .A3(n258), .ZN(n8) );
  XOR2_X1 U229 ( .A(n54), .B(n55), .Z(n261) );
  XOR2_X1 U230 ( .A(n12), .B(n261), .Z(product[4]) );
  NAND2_X1 U231 ( .A1(n12), .A2(n54), .ZN(n262) );
  NAND2_X1 U232 ( .A1(n12), .A2(n55), .ZN(n263) );
  NAND2_X1 U233 ( .A1(n54), .A2(n55), .ZN(n264) );
  XOR2_X1 U234 ( .A(n50), .B(n53), .Z(n265) );
  XOR2_X1 U235 ( .A(n216), .B(n265), .Z(product[5]) );
  NAND2_X1 U236 ( .A1(n230), .A2(n50), .ZN(n266) );
  NAND2_X1 U237 ( .A1(n231), .A2(n53), .ZN(n267) );
  NAND2_X1 U238 ( .A1(n50), .A2(n53), .ZN(n268) );
  NAND3_X1 U239 ( .A1(n272), .A2(n273), .A3(n274), .ZN(n270) );
  XNOR2_X2 U240 ( .A(a[2]), .B(a[1]), .ZN(n271) );
  XNOR2_X1 U241 ( .A(a[2]), .B(a[1]), .ZN(n298) );
  NAND2_X1 U242 ( .A1(n20), .A2(n23), .ZN(n272) );
  NAND2_X1 U243 ( .A1(n232), .A2(n20), .ZN(n273) );
  NAND2_X1 U244 ( .A1(n220), .A2(n23), .ZN(n274) );
  NAND3_X1 U245 ( .A1(n274), .A2(n273), .A3(n272), .ZN(n4) );
  XOR2_X1 U246 ( .A(n19), .B(n18), .Z(n275) );
  XOR2_X1 U247 ( .A(n275), .B(n270), .Z(product[12]) );
  NAND2_X1 U248 ( .A1(n19), .A2(n18), .ZN(n276) );
  NAND2_X1 U249 ( .A1(n4), .A2(n19), .ZN(n277) );
  NAND2_X1 U250 ( .A1(n4), .A2(n18), .ZN(n278) );
  NAND3_X1 U251 ( .A1(n278), .A2(n277), .A3(n276), .ZN(n3) );
  INV_X1 U252 ( .A(n15), .ZN(n281) );
  INV_X1 U253 ( .A(n21), .ZN(n284) );
  INV_X1 U254 ( .A(n317), .ZN(n285) );
  INV_X1 U255 ( .A(n328), .ZN(n282) );
  INV_X1 U256 ( .A(n297), .ZN(n290) );
  INV_X1 U257 ( .A(n306), .ZN(n288) );
  INV_X1 U258 ( .A(n31), .ZN(n287) );
  INV_X1 U259 ( .A(b[0]), .ZN(n280) );
  INV_X1 U260 ( .A(a[5]), .ZN(n286) );
  INV_X1 U261 ( .A(a[7]), .ZN(n283) );
  INV_X1 U262 ( .A(a[3]), .ZN(n289) );
  NAND2_X2 U263 ( .A1(n308), .A2(n337), .ZN(n310) );
  INV_X1 U264 ( .A(a[1]), .ZN(n291) );
  NAND2_X2 U265 ( .A1(n298), .A2(n336), .ZN(n300) );
  XOR2_X2 U266 ( .A(a[6]), .B(n286), .Z(n319) );
  INV_X1 U267 ( .A(n280), .ZN(n279) );
  INV_X2 U268 ( .A(a[0]), .ZN(n292) );
  NOR2_X1 U269 ( .A1(n292), .A2(n280), .ZN(product[0]) );
  OAI22_X1 U270 ( .A1(n293), .A2(n294), .B1(n295), .B2(n292), .ZN(n99) );
  OAI22_X1 U271 ( .A1(n295), .A2(n294), .B1(n296), .B2(n292), .ZN(n98) );
  XNOR2_X1 U272 ( .A(b[6]), .B(a[1]), .ZN(n295) );
  OAI22_X1 U273 ( .A1(n292), .A2(n296), .B1(n294), .B2(n296), .ZN(n297) );
  XNOR2_X1 U274 ( .A(b[7]), .B(a[1]), .ZN(n296) );
  NOR2_X1 U275 ( .A1(n271), .A2(n280), .ZN(n96) );
  OAI22_X1 U276 ( .A1(n299), .A2(n300), .B1(n271), .B2(n301), .ZN(n95) );
  XNOR2_X1 U277 ( .A(a[3]), .B(n250), .ZN(n299) );
  OAI22_X1 U278 ( .A1(n301), .A2(n300), .B1(n271), .B2(n302), .ZN(n94) );
  XNOR2_X1 U279 ( .A(b[1]), .B(a[3]), .ZN(n301) );
  OAI22_X1 U280 ( .A1(n302), .A2(n300), .B1(n271), .B2(n303), .ZN(n93) );
  XNOR2_X1 U281 ( .A(b[2]), .B(a[3]), .ZN(n302) );
  OAI22_X1 U282 ( .A1(n303), .A2(n300), .B1(n271), .B2(n304), .ZN(n92) );
  XNOR2_X1 U283 ( .A(b[3]), .B(a[3]), .ZN(n303) );
  OAI22_X1 U284 ( .A1(n304), .A2(n300), .B1(n271), .B2(n305), .ZN(n91) );
  XNOR2_X1 U285 ( .A(b[4]), .B(a[3]), .ZN(n304) );
  OAI22_X1 U286 ( .A1(n307), .A2(n271), .B1(n300), .B2(n307), .ZN(n306) );
  NOR2_X1 U287 ( .A1(n308), .A2(n280), .ZN(n88) );
  OAI22_X1 U288 ( .A1(n309), .A2(n310), .B1(n308), .B2(n311), .ZN(n87) );
  XNOR2_X1 U289 ( .A(a[5]), .B(n279), .ZN(n309) );
  OAI22_X1 U290 ( .A1(n311), .A2(n310), .B1(n308), .B2(n312), .ZN(n86) );
  XNOR2_X1 U291 ( .A(b[1]), .B(a[5]), .ZN(n311) );
  OAI22_X1 U292 ( .A1(n312), .A2(n310), .B1(n308), .B2(n313), .ZN(n85) );
  XNOR2_X1 U293 ( .A(b[2]), .B(a[5]), .ZN(n312) );
  OAI22_X1 U294 ( .A1(n313), .A2(n310), .B1(n308), .B2(n314), .ZN(n84) );
  XNOR2_X1 U295 ( .A(b[3]), .B(a[5]), .ZN(n313) );
  OAI22_X1 U296 ( .A1(n314), .A2(n310), .B1(n308), .B2(n315), .ZN(n83) );
  XNOR2_X1 U297 ( .A(b[4]), .B(a[5]), .ZN(n314) );
  OAI22_X1 U298 ( .A1(n315), .A2(n310), .B1(n308), .B2(n316), .ZN(n82) );
  XNOR2_X1 U299 ( .A(b[5]), .B(a[5]), .ZN(n315) );
  OAI22_X1 U300 ( .A1(n318), .A2(n308), .B1(n310), .B2(n318), .ZN(n317) );
  NOR2_X1 U301 ( .A1(n319), .A2(n280), .ZN(n80) );
  OAI22_X1 U302 ( .A1(n320), .A2(n321), .B1(n319), .B2(n322), .ZN(n79) );
  XNOR2_X1 U303 ( .A(a[7]), .B(n250), .ZN(n320) );
  OAI22_X1 U304 ( .A1(n323), .A2(n321), .B1(n319), .B2(n324), .ZN(n77) );
  OAI22_X1 U305 ( .A1(n324), .A2(n321), .B1(n319), .B2(n325), .ZN(n76) );
  XNOR2_X1 U306 ( .A(b[3]), .B(a[7]), .ZN(n324) );
  OAI22_X1 U307 ( .A1(n325), .A2(n321), .B1(n319), .B2(n326), .ZN(n75) );
  XNOR2_X1 U308 ( .A(b[4]), .B(a[7]), .ZN(n325) );
  OAI22_X1 U309 ( .A1(n326), .A2(n321), .B1(n319), .B2(n327), .ZN(n74) );
  XNOR2_X1 U310 ( .A(b[5]), .B(a[7]), .ZN(n326) );
  OAI22_X1 U311 ( .A1(n329), .A2(n319), .B1(n321), .B2(n329), .ZN(n328) );
  OAI21_X1 U312 ( .B1(n279), .B2(n291), .A(n294), .ZN(n72) );
  OAI21_X1 U313 ( .B1(n289), .B2(n300), .A(n330), .ZN(n71) );
  OR3_X1 U314 ( .A1(n271), .A2(n250), .A3(n289), .ZN(n330) );
  OAI21_X1 U315 ( .B1(n286), .B2(n310), .A(n331), .ZN(n70) );
  OR3_X1 U316 ( .A1(n308), .A2(n279), .A3(n286), .ZN(n331) );
  OAI21_X1 U317 ( .B1(n283), .B2(n321), .A(n332), .ZN(n69) );
  OR3_X1 U318 ( .A1(n319), .A2(n279), .A3(n283), .ZN(n332) );
  XNOR2_X1 U319 ( .A(n333), .B(n334), .ZN(n38) );
  OR2_X1 U320 ( .A1(n333), .A2(n334), .ZN(n37) );
  OAI22_X1 U321 ( .A1(n305), .A2(n300), .B1(n271), .B2(n335), .ZN(n334) );
  XNOR2_X1 U322 ( .A(b[5]), .B(a[3]), .ZN(n305) );
  OAI22_X1 U323 ( .A1(n322), .A2(n321), .B1(n319), .B2(n323), .ZN(n333) );
  XNOR2_X1 U324 ( .A(b[2]), .B(a[7]), .ZN(n323) );
  XNOR2_X1 U325 ( .A(b[1]), .B(a[7]), .ZN(n322) );
  OAI22_X1 U326 ( .A1(n335), .A2(n300), .B1(n271), .B2(n307), .ZN(n31) );
  XNOR2_X1 U327 ( .A(b[7]), .B(a[3]), .ZN(n307) );
  XNOR2_X1 U328 ( .A(n289), .B(a[2]), .ZN(n336) );
  XNOR2_X1 U329 ( .A(b[6]), .B(a[3]), .ZN(n335) );
  OAI22_X1 U330 ( .A1(n316), .A2(n310), .B1(n308), .B2(n318), .ZN(n21) );
  XNOR2_X1 U331 ( .A(b[7]), .B(a[5]), .ZN(n318) );
  XNOR2_X1 U332 ( .A(n286), .B(a[4]), .ZN(n337) );
  XNOR2_X1 U333 ( .A(b[6]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U334 ( .A1(n327), .A2(n321), .B1(n319), .B2(n329), .ZN(n15) );
  XNOR2_X1 U335 ( .A(b[7]), .B(a[7]), .ZN(n329) );
  NAND2_X1 U336 ( .A1(n319), .A2(n338), .ZN(n321) );
  XNOR2_X1 U337 ( .A(n283), .B(a[6]), .ZN(n338) );
  XNOR2_X1 U338 ( .A(b[6]), .B(a[7]), .ZN(n327) );
  OAI22_X1 U339 ( .A1(n250), .A2(n294), .B1(n339), .B2(n292), .ZN(n104) );
  OAI22_X1 U340 ( .A1(n269), .A2(n294), .B1(n340), .B2(n292), .ZN(n103) );
  XNOR2_X1 U341 ( .A(b[1]), .B(a[1]), .ZN(n339) );
  OAI22_X1 U342 ( .A1(n340), .A2(n294), .B1(n341), .B2(n292), .ZN(n102) );
  XNOR2_X1 U343 ( .A(b[2]), .B(a[1]), .ZN(n340) );
  OAI22_X1 U344 ( .A1(n341), .A2(n294), .B1(n342), .B2(n292), .ZN(n101) );
  XNOR2_X1 U345 ( .A(b[3]), .B(a[1]), .ZN(n341) );
  OAI22_X1 U346 ( .A1(n342), .A2(n294), .B1(n293), .B2(n292), .ZN(n100) );
  XNOR2_X1 U347 ( .A(b[5]), .B(a[1]), .ZN(n293) );
  NAND2_X1 U348 ( .A1(a[1]), .A2(n292), .ZN(n294) );
  XNOR2_X1 U349 ( .A(b[4]), .B(a[1]), .ZN(n342) );
endmodule


module datapath_DW01_add_18 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n71;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  CLKBUF_X1 U1 ( .A(carry[5]), .Z(n1) );
  CLKBUF_X1 U2 ( .A(carry[6]), .Z(n2) );
  NAND3_X1 U3 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n3) );
  NAND3_X1 U4 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n4) );
  XOR2_X1 U5 ( .A(B[4]), .B(A[4]), .Z(n5) );
  XOR2_X1 U6 ( .A(n4), .B(n5), .Z(SUM[4]) );
  NAND2_X1 U7 ( .A1(n3), .A2(B[4]), .ZN(n6) );
  NAND2_X1 U8 ( .A1(carry[4]), .A2(A[4]), .ZN(n7) );
  NAND2_X1 U9 ( .A1(B[4]), .A2(A[4]), .ZN(n8) );
  NAND3_X1 U10 ( .A1(n6), .A2(n7), .A3(n8), .ZN(carry[5]) );
  CLKBUF_X1 U11 ( .A(n56), .Z(n9) );
  NAND3_X1 U12 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n10) );
  NAND2_X1 U13 ( .A1(B[12]), .A2(A[12]), .ZN(n63) );
  CLKBUF_X1 U14 ( .A(n10), .Z(n11) );
  NAND3_X1 U15 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n12) );
  XOR2_X1 U16 ( .A(B[6]), .B(A[6]), .Z(n13) );
  XOR2_X1 U17 ( .A(n2), .B(n13), .Z(SUM[6]) );
  NAND2_X1 U18 ( .A1(carry[6]), .A2(B[6]), .ZN(n14) );
  NAND2_X1 U19 ( .A1(carry[6]), .A2(A[6]), .ZN(n15) );
  NAND2_X1 U20 ( .A1(B[6]), .A2(A[6]), .ZN(n16) );
  NAND3_X1 U21 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[7]) );
  CLKBUF_X1 U22 ( .A(n37), .Z(n17) );
  XOR2_X1 U23 ( .A(n71), .B(A[1]), .Z(n18) );
  XOR2_X1 U24 ( .A(B[1]), .B(n18), .Z(SUM[1]) );
  NAND2_X1 U25 ( .A1(B[1]), .A2(n71), .ZN(n19) );
  NAND2_X1 U26 ( .A1(B[1]), .A2(A[1]), .ZN(n20) );
  NAND2_X1 U27 ( .A1(n71), .A2(A[1]), .ZN(n21) );
  NAND3_X1 U28 ( .A1(n19), .A2(n20), .A3(n21), .ZN(carry[2]) );
  XOR2_X1 U29 ( .A(B[5]), .B(A[5]), .Z(n22) );
  XOR2_X1 U30 ( .A(n1), .B(n22), .Z(SUM[5]) );
  NAND2_X1 U31 ( .A1(carry[5]), .A2(B[5]), .ZN(n23) );
  NAND2_X1 U32 ( .A1(carry[5]), .A2(A[5]), .ZN(n24) );
  NAND2_X1 U33 ( .A1(B[5]), .A2(A[5]), .ZN(n25) );
  NAND3_X1 U34 ( .A1(n23), .A2(n24), .A3(n25), .ZN(carry[6]) );
  XOR2_X1 U35 ( .A(B[7]), .B(A[7]), .Z(n26) );
  XOR2_X1 U36 ( .A(n11), .B(n26), .Z(SUM[7]) );
  NAND2_X1 U37 ( .A1(n10), .A2(B[7]), .ZN(n27) );
  NAND2_X1 U38 ( .A1(carry[7]), .A2(A[7]), .ZN(n28) );
  NAND2_X1 U39 ( .A1(B[7]), .A2(A[7]), .ZN(n29) );
  NAND3_X1 U40 ( .A1(n27), .A2(n28), .A3(n29), .ZN(carry[8]) );
  NAND3_X1 U41 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n30) );
  NAND3_X1 U42 ( .A1(n35), .A2(n34), .A3(n36), .ZN(n31) );
  NAND3_X1 U43 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n32) );
  XOR2_X1 U44 ( .A(B[8]), .B(A[8]), .Z(n33) );
  XOR2_X1 U45 ( .A(carry[8]), .B(n33), .Z(SUM[8]) );
  NAND2_X1 U46 ( .A1(n12), .A2(B[8]), .ZN(n34) );
  NAND2_X1 U47 ( .A1(carry[8]), .A2(A[8]), .ZN(n35) );
  NAND2_X1 U48 ( .A1(B[8]), .A2(A[8]), .ZN(n36) );
  NAND3_X1 U49 ( .A1(n34), .A2(n35), .A3(n36), .ZN(carry[9]) );
  NAND3_X1 U50 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n37) );
  XOR2_X1 U51 ( .A(A[2]), .B(B[2]), .Z(n38) );
  XOR2_X1 U52 ( .A(n38), .B(carry[2]), .Z(SUM[2]) );
  NAND2_X1 U53 ( .A1(A[2]), .A2(B[2]), .ZN(n39) );
  NAND2_X1 U54 ( .A1(A[2]), .A2(carry[2]), .ZN(n40) );
  NAND2_X1 U55 ( .A1(B[2]), .A2(carry[2]), .ZN(n41) );
  NAND3_X1 U56 ( .A1(n39), .A2(n40), .A3(n41), .ZN(carry[3]) );
  XOR2_X1 U57 ( .A(A[3]), .B(B[3]), .Z(n42) );
  XOR2_X1 U58 ( .A(n42), .B(carry[3]), .Z(SUM[3]) );
  NAND2_X1 U59 ( .A1(A[3]), .A2(B[3]), .ZN(n43) );
  NAND2_X1 U60 ( .A1(A[3]), .A2(n30), .ZN(n44) );
  NAND2_X1 U61 ( .A1(B[3]), .A2(carry[3]), .ZN(n45) );
  NAND3_X1 U62 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[4]) );
  XOR2_X1 U63 ( .A(B[9]), .B(A[9]), .Z(n46) );
  XOR2_X1 U64 ( .A(n31), .B(n46), .Z(SUM[9]) );
  NAND2_X1 U65 ( .A1(n31), .A2(B[9]), .ZN(n47) );
  NAND2_X1 U66 ( .A1(carry[9]), .A2(A[9]), .ZN(n48) );
  NAND2_X1 U67 ( .A1(B[9]), .A2(A[9]), .ZN(n49) );
  NAND3_X1 U68 ( .A1(n47), .A2(n48), .A3(n49), .ZN(carry[10]) );
  CLKBUF_X1 U69 ( .A(n32), .Z(n50) );
  XOR2_X1 U70 ( .A(B[10]), .B(A[10]), .Z(n51) );
  XOR2_X1 U71 ( .A(n17), .B(n51), .Z(SUM[10]) );
  NAND2_X1 U72 ( .A1(n37), .A2(B[10]), .ZN(n52) );
  NAND2_X1 U73 ( .A1(carry[10]), .A2(A[10]), .ZN(n53) );
  NAND2_X1 U74 ( .A1(B[10]), .A2(A[10]), .ZN(n54) );
  NAND3_X1 U75 ( .A1(n52), .A2(n53), .A3(n54), .ZN(carry[11]) );
  NAND3_X1 U76 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n55) );
  NAND3_X1 U77 ( .A1(n63), .A2(n65), .A3(n64), .ZN(n56) );
  XOR2_X1 U78 ( .A(B[11]), .B(A[11]), .Z(n57) );
  XOR2_X1 U79 ( .A(n50), .B(n57), .Z(SUM[11]) );
  NAND2_X1 U80 ( .A1(n32), .A2(B[11]), .ZN(n58) );
  NAND2_X1 U81 ( .A1(carry[11]), .A2(A[11]), .ZN(n59) );
  NAND2_X1 U82 ( .A1(B[11]), .A2(A[11]), .ZN(n60) );
  NAND3_X1 U83 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[12]) );
  XNOR2_X1 U84 ( .A(carry[15]), .B(n61), .ZN(SUM[15]) );
  XNOR2_X1 U85 ( .A(B[15]), .B(A[15]), .ZN(n61) );
  XOR2_X1 U86 ( .A(A[12]), .B(B[12]), .Z(n62) );
  XOR2_X1 U87 ( .A(n62), .B(n55), .Z(SUM[12]) );
  NAND2_X1 U88 ( .A1(carry[12]), .A2(A[12]), .ZN(n64) );
  NAND2_X1 U89 ( .A1(B[12]), .A2(carry[12]), .ZN(n65) );
  NAND3_X1 U90 ( .A1(n63), .A2(n65), .A3(n64), .ZN(carry[13]) );
  XOR2_X1 U91 ( .A(A[13]), .B(B[13]), .Z(n66) );
  XOR2_X1 U92 ( .A(n66), .B(n9), .Z(SUM[13]) );
  NAND2_X1 U93 ( .A1(A[13]), .A2(B[13]), .ZN(n67) );
  NAND2_X1 U94 ( .A1(A[13]), .A2(n56), .ZN(n68) );
  NAND2_X1 U95 ( .A1(B[13]), .A2(carry[13]), .ZN(n69) );
  NAND3_X1 U96 ( .A1(n67), .A2(n68), .A3(n69), .ZN(carry[14]) );
  XOR2_X1 U97 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U98 ( .A1(B[0]), .A2(A[0]), .ZN(n71) );
endmodule


module datapath_DW_mult_tc_17 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347;

  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n291), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n290), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n294), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n293), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n295), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n88), .B(n94), .CI(n101), .CO(n53), .S(n54) );
  INV_X2 U157 ( .A(n286), .ZN(n285) );
  BUF_X1 U158 ( .A(n303), .Z(n259) );
  NAND2_X1 U159 ( .A1(n303), .A2(n341), .ZN(n305) );
  INV_X1 U160 ( .A(n15), .ZN(n287) );
  INV_X1 U161 ( .A(a[0]), .ZN(n297) );
  AND2_X1 U162 ( .A1(n95), .A2(n102), .ZN(n206) );
  XNOR2_X1 U163 ( .A(n288), .B(n15), .ZN(n207) );
  AND3_X1 U164 ( .A1(n260), .A2(n261), .A3(n262), .ZN(product[15]) );
  NAND3_X1 U165 ( .A1(n271), .A2(n270), .A3(n272), .ZN(n209) );
  XNOR2_X1 U166 ( .A(n226), .B(n210), .ZN(product[5]) );
  XNOR2_X1 U167 ( .A(n50), .B(n53), .ZN(n210) );
  XOR2_X1 U168 ( .A(n33), .B(n28), .Z(n211) );
  XOR2_X1 U169 ( .A(n7), .B(n211), .Z(product[9]) );
  NAND2_X1 U170 ( .A1(n7), .A2(n33), .ZN(n212) );
  NAND2_X1 U171 ( .A1(n7), .A2(n28), .ZN(n213) );
  NAND2_X1 U172 ( .A1(n33), .A2(n28), .ZN(n214) );
  NAND3_X1 U173 ( .A1(n212), .A2(n213), .A3(n214), .ZN(n6) );
  NAND3_X1 U174 ( .A1(n283), .A2(n282), .A3(n281), .ZN(n215) );
  NAND3_X1 U175 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n216) );
  NAND3_X1 U176 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n217) );
  NAND2_X1 U177 ( .A1(n11), .A2(n50), .ZN(n218) );
  NAND3_X1 U178 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n219) );
  NAND3_X1 U179 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n220) );
  XNOR2_X1 U180 ( .A(n221), .B(n248), .ZN(product[3]) );
  XNOR2_X1 U181 ( .A(n56), .B(n71), .ZN(n221) );
  NAND3_X1 U182 ( .A1(n218), .A2(n250), .A3(n251), .ZN(n222) );
  NAND3_X1 U183 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n223) );
  NAND3_X1 U184 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n224) );
  NAND3_X1 U185 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n225) );
  NAND3_X1 U186 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n226) );
  XOR2_X1 U187 ( .A(n18), .B(n19), .Z(n227) );
  XOR2_X1 U188 ( .A(n4), .B(n227), .Z(product[12]) );
  NAND2_X1 U189 ( .A1(n4), .A2(n18), .ZN(n228) );
  NAND2_X1 U190 ( .A1(n4), .A2(n19), .ZN(n229) );
  NAND2_X1 U191 ( .A1(n18), .A2(n19), .ZN(n230) );
  NAND3_X1 U192 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n3) );
  XOR2_X1 U193 ( .A(n27), .B(n24), .Z(n231) );
  XOR2_X1 U194 ( .A(n6), .B(n231), .Z(product[10]) );
  NAND2_X1 U195 ( .A1(n6), .A2(n27), .ZN(n232) );
  NAND2_X1 U196 ( .A1(n6), .A2(n24), .ZN(n233) );
  NAND2_X1 U197 ( .A1(n27), .A2(n24), .ZN(n234) );
  NAND3_X1 U198 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n5) );
  XOR2_X1 U199 ( .A(n54), .B(n206), .Z(n235) );
  XOR2_X1 U200 ( .A(n12), .B(n235), .Z(product[4]) );
  NAND2_X1 U201 ( .A1(n215), .A2(n54), .ZN(n236) );
  NAND2_X1 U202 ( .A1(n215), .A2(n206), .ZN(n237) );
  NAND2_X1 U203 ( .A1(n54), .A2(n206), .ZN(n238) );
  NAND3_X1 U204 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n11) );
  NAND2_X1 U205 ( .A1(a[4]), .A2(a[3]), .ZN(n241) );
  NAND2_X1 U206 ( .A1(n239), .A2(n240), .ZN(n242) );
  NAND2_X2 U207 ( .A1(n241), .A2(n242), .ZN(n313) );
  INV_X1 U208 ( .A(a[4]), .ZN(n239) );
  INV_X1 U209 ( .A(a[3]), .ZN(n240) );
  XOR2_X1 U210 ( .A(n23), .B(n20), .Z(n243) );
  XOR2_X1 U211 ( .A(n224), .B(n243), .Z(product[11]) );
  NAND2_X1 U212 ( .A1(n5), .A2(n23), .ZN(n244) );
  NAND2_X1 U213 ( .A1(n223), .A2(n20), .ZN(n245) );
  NAND2_X1 U214 ( .A1(n23), .A2(n20), .ZN(n246) );
  NAND3_X1 U215 ( .A1(n245), .A2(n244), .A3(n246), .ZN(n4) );
  NAND3_X1 U216 ( .A1(n218), .A2(n250), .A3(n251), .ZN(n247) );
  NAND3_X1 U217 ( .A1(n278), .A2(n279), .A3(n280), .ZN(n248) );
  XNOR2_X1 U218 ( .A(n2), .B(n207), .ZN(product[14]) );
  NAND2_X1 U219 ( .A1(n11), .A2(n50), .ZN(n249) );
  NAND2_X1 U220 ( .A1(n225), .A2(n53), .ZN(n250) );
  NAND2_X1 U221 ( .A1(n50), .A2(n53), .ZN(n251) );
  NAND3_X1 U222 ( .A1(n250), .A2(n249), .A3(n251), .ZN(n10) );
  XOR2_X1 U223 ( .A(n95), .B(n102), .Z(n56) );
  OAI22_X1 U224 ( .A1(n304), .A2(n305), .B1(n259), .B2(n306), .ZN(n252) );
  XOR2_X1 U225 ( .A(n17), .B(n287), .Z(n253) );
  XOR2_X1 U226 ( .A(n220), .B(n253), .Z(product[13]) );
  NAND2_X1 U227 ( .A1(n219), .A2(n17), .ZN(n254) );
  NAND2_X1 U228 ( .A1(n3), .A2(n287), .ZN(n255) );
  NAND2_X1 U229 ( .A1(n17), .A2(n287), .ZN(n256) );
  NAND3_X1 U230 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n2) );
  NAND3_X1 U231 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n257) );
  XOR2_X1 U232 ( .A(n252), .B(n102), .Z(n258) );
  XNOR2_X1 U233 ( .A(a[2]), .B(a[1]), .ZN(n303) );
  NAND2_X1 U234 ( .A1(n217), .A2(n288), .ZN(n260) );
  NAND2_X1 U235 ( .A1(n216), .A2(n15), .ZN(n261) );
  NAND2_X1 U236 ( .A1(n288), .A2(n15), .ZN(n262) );
  XOR2_X1 U237 ( .A(n46), .B(n49), .Z(n263) );
  XOR2_X1 U238 ( .A(n222), .B(n263), .Z(product[6]) );
  NAND2_X1 U239 ( .A1(n247), .A2(n46), .ZN(n264) );
  NAND2_X1 U240 ( .A1(n10), .A2(n49), .ZN(n265) );
  NAND2_X1 U241 ( .A1(n46), .A2(n49), .ZN(n266) );
  NAND3_X1 U242 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n9) );
  NAND3_X1 U243 ( .A1(n270), .A2(n271), .A3(n272), .ZN(n267) );
  XNOR2_X1 U244 ( .A(b[1]), .B(a[1]), .ZN(n268) );
  XOR2_X1 U245 ( .A(n40), .B(n45), .Z(n269) );
  XOR2_X1 U246 ( .A(n269), .B(n257), .Z(product[7]) );
  NAND2_X1 U247 ( .A1(n40), .A2(n45), .ZN(n270) );
  NAND2_X1 U248 ( .A1(n40), .A2(n9), .ZN(n271) );
  NAND2_X1 U249 ( .A1(n9), .A2(n45), .ZN(n272) );
  NAND3_X1 U250 ( .A1(n271), .A2(n270), .A3(n272), .ZN(n8) );
  XOR2_X1 U251 ( .A(n34), .B(n39), .Z(n273) );
  XOR2_X1 U252 ( .A(n273), .B(n267), .Z(product[8]) );
  NAND2_X1 U253 ( .A1(n34), .A2(n39), .ZN(n274) );
  NAND2_X1 U254 ( .A1(n34), .A2(n8), .ZN(n275) );
  NAND2_X1 U255 ( .A1(n209), .A2(n39), .ZN(n276) );
  NAND3_X1 U256 ( .A1(n274), .A2(n275), .A3(n276), .ZN(n7) );
  XOR2_X1 U257 ( .A(n103), .B(n96), .Z(n277) );
  XOR2_X1 U258 ( .A(n277), .B(n14), .Z(product[2]) );
  NAND2_X1 U259 ( .A1(n103), .A2(n96), .ZN(n278) );
  NAND2_X1 U260 ( .A1(n103), .A2(n14), .ZN(n279) );
  NAND2_X1 U261 ( .A1(n96), .A2(n14), .ZN(n280) );
  NAND3_X1 U262 ( .A1(n278), .A2(n279), .A3(n280), .ZN(n13) );
  NAND2_X1 U263 ( .A1(n258), .A2(n71), .ZN(n281) );
  NAND2_X1 U264 ( .A1(n258), .A2(n13), .ZN(n282) );
  NAND2_X1 U265 ( .A1(n71), .A2(n13), .ZN(n283) );
  NAND3_X1 U266 ( .A1(n281), .A2(n282), .A3(n283), .ZN(n12) );
  CLKBUF_X1 U267 ( .A(b[1]), .Z(n284) );
  INV_X1 U268 ( .A(n21), .ZN(n290) );
  INV_X1 U269 ( .A(n322), .ZN(n291) );
  INV_X1 U270 ( .A(n333), .ZN(n288) );
  INV_X1 U271 ( .A(n302), .ZN(n295) );
  INV_X1 U272 ( .A(n311), .ZN(n294) );
  INV_X1 U273 ( .A(n31), .ZN(n293) );
  INV_X1 U274 ( .A(b[0]), .ZN(n286) );
  INV_X1 U275 ( .A(a[5]), .ZN(n292) );
  INV_X1 U276 ( .A(a[7]), .ZN(n289) );
  NAND2_X2 U277 ( .A1(n313), .A2(n342), .ZN(n315) );
  INV_X1 U278 ( .A(a[1]), .ZN(n296) );
  XOR2_X2 U279 ( .A(a[6]), .B(n292), .Z(n324) );
  NOR2_X1 U280 ( .A1(n297), .A2(n286), .ZN(product[0]) );
  OAI22_X1 U281 ( .A1(n298), .A2(n299), .B1(n300), .B2(n297), .ZN(n99) );
  OAI22_X1 U282 ( .A1(n300), .A2(n299), .B1(n301), .B2(n297), .ZN(n98) );
  XNOR2_X1 U283 ( .A(b[6]), .B(a[1]), .ZN(n300) );
  OAI22_X1 U284 ( .A1(n297), .A2(n301), .B1(n299), .B2(n301), .ZN(n302) );
  XNOR2_X1 U285 ( .A(b[7]), .B(a[1]), .ZN(n301) );
  NOR2_X1 U286 ( .A1(n259), .A2(n286), .ZN(n96) );
  OAI22_X1 U287 ( .A1(n304), .A2(n305), .B1(n259), .B2(n306), .ZN(n95) );
  XNOR2_X1 U288 ( .A(a[3]), .B(n285), .ZN(n304) );
  OAI22_X1 U289 ( .A1(n306), .A2(n305), .B1(n259), .B2(n307), .ZN(n94) );
  XNOR2_X1 U290 ( .A(b[1]), .B(a[3]), .ZN(n306) );
  OAI22_X1 U291 ( .A1(n307), .A2(n305), .B1(n259), .B2(n308), .ZN(n93) );
  XNOR2_X1 U292 ( .A(b[2]), .B(a[3]), .ZN(n307) );
  OAI22_X1 U293 ( .A1(n308), .A2(n305), .B1(n259), .B2(n309), .ZN(n92) );
  XNOR2_X1 U294 ( .A(b[3]), .B(a[3]), .ZN(n308) );
  OAI22_X1 U295 ( .A1(n309), .A2(n305), .B1(n259), .B2(n310), .ZN(n91) );
  XNOR2_X1 U296 ( .A(b[4]), .B(a[3]), .ZN(n309) );
  OAI22_X1 U297 ( .A1(n312), .A2(n259), .B1(n305), .B2(n312), .ZN(n311) );
  NOR2_X1 U298 ( .A1(n313), .A2(n286), .ZN(n88) );
  OAI22_X1 U299 ( .A1(n314), .A2(n315), .B1(n313), .B2(n316), .ZN(n87) );
  XNOR2_X1 U300 ( .A(a[5]), .B(n285), .ZN(n314) );
  OAI22_X1 U301 ( .A1(n316), .A2(n315), .B1(n313), .B2(n317), .ZN(n86) );
  XNOR2_X1 U302 ( .A(b[1]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U303 ( .A1(n317), .A2(n315), .B1(n313), .B2(n318), .ZN(n85) );
  XNOR2_X1 U304 ( .A(b[2]), .B(a[5]), .ZN(n317) );
  OAI22_X1 U305 ( .A1(n318), .A2(n315), .B1(n313), .B2(n319), .ZN(n84) );
  XNOR2_X1 U306 ( .A(b[3]), .B(a[5]), .ZN(n318) );
  OAI22_X1 U307 ( .A1(n319), .A2(n315), .B1(n313), .B2(n320), .ZN(n83) );
  XNOR2_X1 U308 ( .A(b[4]), .B(a[5]), .ZN(n319) );
  OAI22_X1 U309 ( .A1(n320), .A2(n315), .B1(n313), .B2(n321), .ZN(n82) );
  XNOR2_X1 U310 ( .A(b[5]), .B(a[5]), .ZN(n320) );
  OAI22_X1 U311 ( .A1(n323), .A2(n313), .B1(n315), .B2(n323), .ZN(n322) );
  NOR2_X1 U312 ( .A1(n324), .A2(n286), .ZN(n80) );
  OAI22_X1 U313 ( .A1(n325), .A2(n326), .B1(n324), .B2(n327), .ZN(n79) );
  XNOR2_X1 U314 ( .A(a[7]), .B(n285), .ZN(n325) );
  OAI22_X1 U315 ( .A1(n328), .A2(n326), .B1(n324), .B2(n329), .ZN(n77) );
  OAI22_X1 U316 ( .A1(n329), .A2(n326), .B1(n324), .B2(n330), .ZN(n76) );
  XNOR2_X1 U317 ( .A(b[3]), .B(a[7]), .ZN(n329) );
  OAI22_X1 U318 ( .A1(n330), .A2(n326), .B1(n324), .B2(n331), .ZN(n75) );
  XNOR2_X1 U319 ( .A(b[4]), .B(a[7]), .ZN(n330) );
  OAI22_X1 U320 ( .A1(n331), .A2(n326), .B1(n324), .B2(n332), .ZN(n74) );
  XNOR2_X1 U321 ( .A(b[5]), .B(a[7]), .ZN(n331) );
  OAI22_X1 U322 ( .A1(n334), .A2(n324), .B1(n326), .B2(n334), .ZN(n333) );
  OAI21_X1 U323 ( .B1(n285), .B2(n296), .A(n299), .ZN(n72) );
  OAI21_X1 U324 ( .B1(n240), .B2(n305), .A(n335), .ZN(n71) );
  OR3_X1 U325 ( .A1(n259), .A2(n285), .A3(n240), .ZN(n335) );
  OAI21_X1 U326 ( .B1(n292), .B2(n315), .A(n336), .ZN(n70) );
  OR3_X1 U327 ( .A1(n313), .A2(n285), .A3(n292), .ZN(n336) );
  OAI21_X1 U328 ( .B1(n289), .B2(n326), .A(n337), .ZN(n69) );
  OR3_X1 U329 ( .A1(n324), .A2(n285), .A3(n289), .ZN(n337) );
  XNOR2_X1 U330 ( .A(n338), .B(n339), .ZN(n38) );
  OR2_X1 U331 ( .A1(n338), .A2(n339), .ZN(n37) );
  OAI22_X1 U332 ( .A1(n310), .A2(n305), .B1(n259), .B2(n340), .ZN(n339) );
  XNOR2_X1 U333 ( .A(b[5]), .B(a[3]), .ZN(n310) );
  OAI22_X1 U334 ( .A1(n327), .A2(n326), .B1(n324), .B2(n328), .ZN(n338) );
  XNOR2_X1 U335 ( .A(b[2]), .B(a[7]), .ZN(n328) );
  XNOR2_X1 U336 ( .A(n284), .B(a[7]), .ZN(n327) );
  OAI22_X1 U337 ( .A1(n340), .A2(n305), .B1(n259), .B2(n312), .ZN(n31) );
  XNOR2_X1 U338 ( .A(b[7]), .B(a[3]), .ZN(n312) );
  XNOR2_X1 U339 ( .A(n240), .B(a[2]), .ZN(n341) );
  XNOR2_X1 U340 ( .A(b[6]), .B(a[3]), .ZN(n340) );
  OAI22_X1 U341 ( .A1(n321), .A2(n315), .B1(n313), .B2(n323), .ZN(n21) );
  XNOR2_X1 U342 ( .A(b[7]), .B(a[5]), .ZN(n323) );
  XNOR2_X1 U343 ( .A(n292), .B(a[4]), .ZN(n342) );
  XNOR2_X1 U344 ( .A(b[6]), .B(a[5]), .ZN(n321) );
  OAI22_X1 U345 ( .A1(n332), .A2(n326), .B1(n324), .B2(n334), .ZN(n15) );
  XNOR2_X1 U346 ( .A(b[7]), .B(a[7]), .ZN(n334) );
  NAND2_X1 U347 ( .A1(n324), .A2(n343), .ZN(n326) );
  XNOR2_X1 U348 ( .A(n289), .B(a[6]), .ZN(n343) );
  XNOR2_X1 U349 ( .A(b[6]), .B(a[7]), .ZN(n332) );
  OAI22_X1 U350 ( .A1(n285), .A2(n299), .B1(n344), .B2(n297), .ZN(n104) );
  OAI22_X1 U351 ( .A1(n268), .A2(n299), .B1(n345), .B2(n297), .ZN(n103) );
  XNOR2_X1 U352 ( .A(b[1]), .B(a[1]), .ZN(n344) );
  OAI22_X1 U353 ( .A1(n345), .A2(n299), .B1(n346), .B2(n297), .ZN(n102) );
  XNOR2_X1 U354 ( .A(b[2]), .B(a[1]), .ZN(n345) );
  OAI22_X1 U355 ( .A1(n346), .A2(n299), .B1(n347), .B2(n297), .ZN(n101) );
  XNOR2_X1 U356 ( .A(b[3]), .B(a[1]), .ZN(n346) );
  OAI22_X1 U357 ( .A1(n347), .A2(n299), .B1(n298), .B2(n297), .ZN(n100) );
  XNOR2_X1 U358 ( .A(b[5]), .B(a[1]), .ZN(n298) );
  NAND2_X1 U359 ( .A1(a[1]), .A2(n297), .ZN(n299) );
  XNOR2_X1 U360 ( .A(b[4]), .B(a[1]), .ZN(n347) );
endmodule


module datapath_DW01_add_17 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n74;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  CLKBUF_X1 U1 ( .A(carry[7]), .Z(n1) );
  CLKBUF_X1 U2 ( .A(n49), .Z(n2) );
  NAND3_X1 U3 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n3) );
  NAND3_X1 U4 ( .A1(n2), .A2(n50), .A3(n51), .ZN(n4) );
  CLKBUF_X1 U5 ( .A(n34), .Z(n5) );
  XOR2_X1 U6 ( .A(n74), .B(A[1]), .Z(n6) );
  XOR2_X1 U7 ( .A(B[1]), .B(n6), .Z(SUM[1]) );
  NAND2_X1 U8 ( .A1(B[1]), .A2(n74), .ZN(n7) );
  NAND2_X1 U9 ( .A1(B[1]), .A2(A[1]), .ZN(n8) );
  NAND2_X1 U10 ( .A1(n74), .A2(A[1]), .ZN(n9) );
  NAND3_X1 U11 ( .A1(n7), .A2(n8), .A3(n9), .ZN(carry[2]) );
  NAND3_X1 U12 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n10) );
  NAND3_X1 U13 ( .A1(n36), .A2(n37), .A3(n38), .ZN(n11) );
  XOR2_X1 U14 ( .A(B[2]), .B(A[2]), .Z(n12) );
  XOR2_X1 U15 ( .A(carry[2]), .B(n12), .Z(SUM[2]) );
  NAND2_X1 U16 ( .A1(carry[2]), .A2(B[2]), .ZN(n13) );
  NAND2_X1 U17 ( .A1(carry[2]), .A2(A[2]), .ZN(n14) );
  NAND2_X1 U18 ( .A1(B[2]), .A2(A[2]), .ZN(n15) );
  NAND3_X1 U19 ( .A1(n13), .A2(n14), .A3(n15), .ZN(carry[3]) );
  XOR2_X1 U20 ( .A(B[5]), .B(A[5]), .Z(n16) );
  XOR2_X1 U21 ( .A(carry[5]), .B(n16), .Z(SUM[5]) );
  NAND2_X1 U22 ( .A1(n11), .A2(B[5]), .ZN(n17) );
  NAND2_X1 U23 ( .A1(n11), .A2(A[5]), .ZN(n18) );
  NAND2_X1 U24 ( .A1(B[5]), .A2(A[5]), .ZN(n19) );
  NAND3_X1 U25 ( .A1(n17), .A2(n18), .A3(n19), .ZN(carry[6]) );
  CLKBUF_X1 U26 ( .A(n68), .Z(n20) );
  CLKBUF_X1 U27 ( .A(n67), .Z(n21) );
  NAND3_X1 U28 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n22) );
  NAND3_X1 U29 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n23) );
  XOR2_X1 U30 ( .A(B[8]), .B(A[8]), .Z(n24) );
  XOR2_X1 U31 ( .A(n22), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U32 ( .A1(n22), .A2(B[8]), .ZN(n25) );
  NAND2_X1 U33 ( .A1(carry[8]), .A2(A[8]), .ZN(n26) );
  NAND2_X1 U34 ( .A1(B[8]), .A2(A[8]), .ZN(n27) );
  NAND3_X1 U35 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[9]) );
  NAND3_X1 U36 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n28) );
  NAND3_X1 U37 ( .A1(n31), .A2(n32), .A3(n33), .ZN(n29) );
  XOR2_X1 U38 ( .A(B[3]), .B(A[3]), .Z(n30) );
  XOR2_X1 U39 ( .A(carry[3]), .B(n30), .Z(SUM[3]) );
  NAND2_X1 U40 ( .A1(carry[3]), .A2(B[3]), .ZN(n31) );
  NAND2_X1 U41 ( .A1(carry[3]), .A2(A[3]), .ZN(n32) );
  NAND2_X1 U42 ( .A1(B[3]), .A2(A[3]), .ZN(n33) );
  NAND3_X1 U43 ( .A1(n31), .A2(n32), .A3(n33), .ZN(carry[4]) );
  NAND3_X1 U44 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n34) );
  XOR2_X1 U45 ( .A(n29), .B(A[4]), .Z(n35) );
  XOR2_X1 U46 ( .A(B[4]), .B(n35), .Z(SUM[4]) );
  NAND2_X1 U47 ( .A1(n29), .A2(B[4]), .ZN(n36) );
  NAND2_X1 U48 ( .A1(B[4]), .A2(A[4]), .ZN(n37) );
  NAND2_X1 U49 ( .A1(carry[4]), .A2(A[4]), .ZN(n38) );
  NAND3_X1 U50 ( .A1(n36), .A2(n37), .A3(n38), .ZN(carry[5]) );
  CLKBUF_X1 U51 ( .A(n56), .Z(n39) );
  XOR2_X1 U52 ( .A(B[9]), .B(A[9]), .Z(n40) );
  XOR2_X1 U53 ( .A(n23), .B(n40), .Z(SUM[9]) );
  NAND2_X1 U54 ( .A1(n23), .A2(B[9]), .ZN(n41) );
  NAND2_X1 U55 ( .A1(carry[9]), .A2(A[9]), .ZN(n42) );
  NAND2_X1 U56 ( .A1(B[9]), .A2(A[9]), .ZN(n43) );
  NAND3_X1 U57 ( .A1(n41), .A2(n42), .A3(n43), .ZN(carry[10]) );
  XOR2_X1 U58 ( .A(B[6]), .B(A[6]), .Z(n44) );
  XOR2_X1 U59 ( .A(carry[6]), .B(n44), .Z(SUM[6]) );
  NAND2_X1 U60 ( .A1(n10), .A2(B[6]), .ZN(n45) );
  NAND2_X1 U61 ( .A1(n10), .A2(A[6]), .ZN(n46) );
  NAND2_X1 U62 ( .A1(B[6]), .A2(A[6]), .ZN(n47) );
  NAND3_X1 U63 ( .A1(n45), .A2(n46), .A3(n47), .ZN(carry[7]) );
  XOR2_X1 U64 ( .A(B[10]), .B(A[10]), .Z(n48) );
  XOR2_X1 U65 ( .A(n5), .B(n48), .Z(SUM[10]) );
  NAND2_X1 U66 ( .A1(n34), .A2(B[10]), .ZN(n49) );
  NAND2_X1 U67 ( .A1(carry[10]), .A2(A[10]), .ZN(n50) );
  NAND2_X1 U68 ( .A1(B[10]), .A2(A[10]), .ZN(n51) );
  NAND3_X1 U69 ( .A1(n49), .A2(n50), .A3(n51), .ZN(carry[11]) );
  NAND3_X1 U70 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n52) );
  NAND3_X1 U71 ( .A1(n55), .A2(n39), .A3(n57), .ZN(n53) );
  XOR2_X1 U72 ( .A(B[11]), .B(A[11]), .Z(n54) );
  XOR2_X1 U73 ( .A(n4), .B(n54), .Z(SUM[11]) );
  NAND2_X1 U74 ( .A1(n3), .A2(B[11]), .ZN(n55) );
  NAND2_X1 U75 ( .A1(carry[11]), .A2(A[11]), .ZN(n56) );
  NAND2_X1 U76 ( .A1(B[11]), .A2(A[11]), .ZN(n57) );
  XOR2_X1 U77 ( .A(B[7]), .B(A[7]), .Z(n58) );
  XOR2_X1 U78 ( .A(n1), .B(n58), .Z(SUM[7]) );
  NAND2_X1 U79 ( .A1(carry[7]), .A2(B[7]), .ZN(n59) );
  NAND2_X1 U80 ( .A1(n28), .A2(A[7]), .ZN(n60) );
  NAND2_X1 U81 ( .A1(B[7]), .A2(A[7]), .ZN(n61) );
  NAND3_X1 U82 ( .A1(n59), .A2(n61), .A3(n60), .ZN(carry[8]) );
  NAND3_X1 U83 ( .A1(n68), .A2(n67), .A3(n66), .ZN(n62) );
  NAND3_X1 U84 ( .A1(n66), .A2(n21), .A3(n20), .ZN(n63) );
  XNOR2_X1 U85 ( .A(carry[15]), .B(n64), .ZN(SUM[15]) );
  XNOR2_X1 U86 ( .A(B[15]), .B(A[15]), .ZN(n64) );
  NAND2_X1 U87 ( .A1(B[12]), .A2(A[12]), .ZN(n66) );
  XOR2_X1 U88 ( .A(A[12]), .B(B[12]), .Z(n65) );
  XOR2_X1 U89 ( .A(n65), .B(n53), .Z(SUM[12]) );
  NAND2_X1 U90 ( .A1(A[12]), .A2(n52), .ZN(n67) );
  NAND2_X1 U91 ( .A1(B[12]), .A2(n52), .ZN(n68) );
  NAND3_X1 U92 ( .A1(n67), .A2(n66), .A3(n68), .ZN(carry[13]) );
  XOR2_X1 U93 ( .A(A[13]), .B(B[13]), .Z(n69) );
  XOR2_X1 U94 ( .A(n69), .B(n63), .Z(SUM[13]) );
  NAND2_X1 U95 ( .A1(A[13]), .A2(B[13]), .ZN(n70) );
  NAND2_X1 U96 ( .A1(A[13]), .A2(n62), .ZN(n71) );
  NAND2_X1 U97 ( .A1(B[13]), .A2(carry[13]), .ZN(n72) );
  NAND3_X1 U98 ( .A1(n72), .A2(n71), .A3(n70), .ZN(carry[14]) );
  XOR2_X1 U99 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U100 ( .A1(B[0]), .A2(A[0]), .ZN(n74) );
endmodule


module datapath_DW_mult_tc_16 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325;

  FA_X1 U8 ( .A(n34), .B(n39), .CI(n8), .CO(n7), .S(product[8]) );
  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n269), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n268), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n272), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n271), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n274), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  INV_X1 U157 ( .A(n15), .ZN(n265) );
  XOR2_X1 U158 ( .A(a[2]), .B(n261), .Z(n281) );
  AND2_X1 U159 ( .A1(n95), .A2(n102), .ZN(n206) );
  AND3_X1 U160 ( .A1(n232), .A2(n233), .A3(n234), .ZN(product[15]) );
  CLKBUF_X1 U161 ( .A(n254), .Z(n208) );
  NAND3_X1 U162 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n209) );
  NAND3_X1 U163 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n210) );
  XOR2_X1 U164 ( .A(n17), .B(n265), .Z(n211) );
  XOR2_X1 U165 ( .A(n3), .B(n211), .Z(product[13]) );
  NAND2_X1 U166 ( .A1(n3), .A2(n17), .ZN(n212) );
  NAND2_X1 U167 ( .A1(n3), .A2(n265), .ZN(n213) );
  NAND2_X1 U168 ( .A1(n17), .A2(n265), .ZN(n214) );
  NAND3_X1 U169 ( .A1(n212), .A2(n213), .A3(n214), .ZN(n2) );
  NAND3_X1 U170 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n215) );
  NAND3_X1 U171 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n216) );
  NAND3_X1 U172 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n217) );
  NAND3_X1 U173 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n218) );
  XNOR2_X1 U174 ( .A(n12), .B(n219), .ZN(product[4]) );
  XNOR2_X1 U175 ( .A(n54), .B(n206), .ZN(n219) );
  XOR2_X1 U176 ( .A(n18), .B(n19), .Z(n220) );
  XOR2_X1 U177 ( .A(n218), .B(n220), .Z(product[12]) );
  NAND2_X1 U178 ( .A1(n217), .A2(n18), .ZN(n221) );
  NAND2_X1 U179 ( .A1(n4), .A2(n19), .ZN(n222) );
  NAND2_X1 U180 ( .A1(n18), .A2(n19), .ZN(n223) );
  NAND3_X1 U181 ( .A1(n221), .A2(n222), .A3(n223), .ZN(n3) );
  XOR2_X1 U182 ( .A(n102), .B(n95), .Z(n56) );
  INV_X2 U183 ( .A(n261), .ZN(n262) );
  NAND2_X2 U184 ( .A1(n281), .A2(n319), .ZN(n283) );
  XOR2_X1 U185 ( .A(n23), .B(n20), .Z(n224) );
  XOR2_X1 U186 ( .A(n216), .B(n224), .Z(product[11]) );
  NAND2_X1 U187 ( .A1(n215), .A2(n23), .ZN(n225) );
  NAND2_X1 U188 ( .A1(n5), .A2(n20), .ZN(n226) );
  NAND2_X1 U189 ( .A1(n23), .A2(n20), .ZN(n227) );
  NAND3_X1 U190 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n4) );
  NAND2_X1 U191 ( .A1(n12), .A2(n54), .ZN(n228) );
  NAND2_X1 U192 ( .A1(n12), .A2(n206), .ZN(n229) );
  NAND2_X1 U193 ( .A1(n54), .A2(n206), .ZN(n230) );
  NAND3_X1 U194 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n11) );
  XOR2_X1 U195 ( .A(n266), .B(n15), .Z(n231) );
  XOR2_X1 U196 ( .A(n2), .B(n231), .Z(product[14]) );
  NAND2_X1 U197 ( .A1(n2), .A2(n266), .ZN(n232) );
  NAND2_X1 U198 ( .A1(n2), .A2(n15), .ZN(n233) );
  NAND2_X1 U199 ( .A1(n266), .A2(n15), .ZN(n234) );
  NAND3_X1 U200 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n235) );
  XOR2_X1 U201 ( .A(n50), .B(n53), .Z(n236) );
  XOR2_X1 U202 ( .A(n210), .B(n236), .Z(product[5]) );
  NAND2_X1 U203 ( .A1(n209), .A2(n50), .ZN(n237) );
  NAND2_X1 U204 ( .A1(n11), .A2(n53), .ZN(n238) );
  NAND2_X1 U205 ( .A1(n50), .A2(n53), .ZN(n239) );
  NAND3_X1 U206 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n10) );
  NAND3_X1 U207 ( .A1(n244), .A2(n243), .A3(n242), .ZN(n240) );
  XOR2_X1 U208 ( .A(n28), .B(n33), .Z(n241) );
  XOR2_X1 U209 ( .A(n241), .B(n7), .Z(product[9]) );
  NAND2_X1 U210 ( .A1(n28), .A2(n33), .ZN(n242) );
  NAND2_X1 U211 ( .A1(n28), .A2(n7), .ZN(n243) );
  NAND2_X1 U212 ( .A1(n33), .A2(n7), .ZN(n244) );
  NAND3_X1 U213 ( .A1(n244), .A2(n243), .A3(n242), .ZN(n6) );
  XOR2_X1 U214 ( .A(n24), .B(n27), .Z(n245) );
  XOR2_X1 U215 ( .A(n245), .B(n240), .Z(product[10]) );
  NAND2_X1 U216 ( .A1(n24), .A2(n27), .ZN(n246) );
  NAND2_X1 U217 ( .A1(n6), .A2(n24), .ZN(n247) );
  NAND2_X1 U218 ( .A1(n6), .A2(n27), .ZN(n248) );
  NAND3_X1 U219 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n5) );
  NAND3_X1 U220 ( .A1(n255), .A2(n254), .A3(n253), .ZN(n249) );
  NAND3_X1 U221 ( .A1(n255), .A2(n208), .A3(n253), .ZN(n250) );
  INV_X1 U222 ( .A(n264), .ZN(n251) );
  XOR2_X1 U223 ( .A(n46), .B(n49), .Z(n252) );
  XOR2_X1 U224 ( .A(n252), .B(n10), .Z(product[6]) );
  NAND2_X1 U225 ( .A1(n46), .A2(n49), .ZN(n253) );
  NAND2_X1 U226 ( .A1(n46), .A2(n235), .ZN(n254) );
  NAND2_X1 U227 ( .A1(n49), .A2(n235), .ZN(n255) );
  NAND3_X1 U228 ( .A1(n255), .A2(n254), .A3(n253), .ZN(n9) );
  XOR2_X1 U229 ( .A(n40), .B(n45), .Z(n256) );
  XOR2_X1 U230 ( .A(n256), .B(n250), .Z(product[7]) );
  NAND2_X1 U231 ( .A1(n40), .A2(n45), .ZN(n257) );
  NAND2_X1 U232 ( .A1(n40), .A2(n9), .ZN(n258) );
  NAND2_X1 U233 ( .A1(n45), .A2(n249), .ZN(n259) );
  NAND3_X1 U234 ( .A1(n259), .A2(n258), .A3(n257), .ZN(n8) );
  NAND2_X2 U235 ( .A1(n291), .A2(n320), .ZN(n293) );
  XNOR2_X2 U236 ( .A(a[4]), .B(a[3]), .ZN(n291) );
  CLKBUF_X1 U237 ( .A(n281), .Z(n260) );
  INV_X1 U238 ( .A(n21), .ZN(n268) );
  INV_X1 U239 ( .A(n300), .ZN(n269) );
  INV_X1 U240 ( .A(n311), .ZN(n266) );
  INV_X1 U241 ( .A(n280), .ZN(n274) );
  INV_X1 U242 ( .A(n289), .ZN(n272) );
  INV_X1 U243 ( .A(n31), .ZN(n271) );
  INV_X1 U244 ( .A(b[0]), .ZN(n264) );
  XOR2_X1 U245 ( .A(a[6]), .B(n270), .Z(n302) );
  INV_X1 U246 ( .A(a[0]), .ZN(n275) );
  INV_X1 U247 ( .A(a[5]), .ZN(n270) );
  INV_X1 U248 ( .A(a[7]), .ZN(n267) );
  INV_X1 U249 ( .A(a[3]), .ZN(n273) );
  INV_X1 U250 ( .A(a[1]), .ZN(n261) );
  INV_X1 U251 ( .A(n264), .ZN(n263) );
  NOR2_X1 U252 ( .A1(n275), .A2(n264), .ZN(product[0]) );
  OAI22_X1 U253 ( .A1(n276), .A2(n277), .B1(n278), .B2(n275), .ZN(n99) );
  OAI22_X1 U254 ( .A1(n278), .A2(n277), .B1(n279), .B2(n275), .ZN(n98) );
  XNOR2_X1 U255 ( .A(b[6]), .B(n262), .ZN(n278) );
  OAI22_X1 U256 ( .A1(n275), .A2(n279), .B1(n277), .B2(n279), .ZN(n280) );
  XNOR2_X1 U257 ( .A(b[7]), .B(n262), .ZN(n279) );
  NOR2_X1 U258 ( .A1(n281), .A2(n264), .ZN(n96) );
  OAI22_X1 U259 ( .A1(n282), .A2(n283), .B1(n281), .B2(n284), .ZN(n95) );
  XNOR2_X1 U260 ( .A(a[3]), .B(n251), .ZN(n282) );
  OAI22_X1 U261 ( .A1(n284), .A2(n283), .B1(n260), .B2(n285), .ZN(n94) );
  XNOR2_X1 U262 ( .A(b[1]), .B(a[3]), .ZN(n284) );
  OAI22_X1 U263 ( .A1(n285), .A2(n283), .B1(n260), .B2(n286), .ZN(n93) );
  XNOR2_X1 U264 ( .A(b[2]), .B(a[3]), .ZN(n285) );
  OAI22_X1 U265 ( .A1(n286), .A2(n283), .B1(n260), .B2(n287), .ZN(n92) );
  XNOR2_X1 U266 ( .A(b[3]), .B(a[3]), .ZN(n286) );
  OAI22_X1 U267 ( .A1(n287), .A2(n283), .B1(n260), .B2(n288), .ZN(n91) );
  XNOR2_X1 U268 ( .A(b[4]), .B(a[3]), .ZN(n287) );
  OAI22_X1 U269 ( .A1(n290), .A2(n260), .B1(n283), .B2(n290), .ZN(n289) );
  NOR2_X1 U270 ( .A1(n291), .A2(n264), .ZN(n88) );
  OAI22_X1 U271 ( .A1(n292), .A2(n293), .B1(n291), .B2(n294), .ZN(n87) );
  XNOR2_X1 U272 ( .A(a[5]), .B(n263), .ZN(n292) );
  OAI22_X1 U273 ( .A1(n294), .A2(n293), .B1(n291), .B2(n295), .ZN(n86) );
  XNOR2_X1 U274 ( .A(b[1]), .B(a[5]), .ZN(n294) );
  OAI22_X1 U275 ( .A1(n295), .A2(n293), .B1(n291), .B2(n296), .ZN(n85) );
  XNOR2_X1 U276 ( .A(b[2]), .B(a[5]), .ZN(n295) );
  OAI22_X1 U277 ( .A1(n296), .A2(n293), .B1(n291), .B2(n297), .ZN(n84) );
  XNOR2_X1 U278 ( .A(b[3]), .B(a[5]), .ZN(n296) );
  OAI22_X1 U279 ( .A1(n297), .A2(n293), .B1(n291), .B2(n298), .ZN(n83) );
  XNOR2_X1 U280 ( .A(b[4]), .B(a[5]), .ZN(n297) );
  OAI22_X1 U281 ( .A1(n298), .A2(n293), .B1(n291), .B2(n299), .ZN(n82) );
  XNOR2_X1 U282 ( .A(b[5]), .B(a[5]), .ZN(n298) );
  OAI22_X1 U283 ( .A1(n301), .A2(n291), .B1(n293), .B2(n301), .ZN(n300) );
  NOR2_X1 U284 ( .A1(n302), .A2(n264), .ZN(n80) );
  OAI22_X1 U285 ( .A1(n303), .A2(n304), .B1(n302), .B2(n305), .ZN(n79) );
  XNOR2_X1 U286 ( .A(a[7]), .B(n251), .ZN(n303) );
  OAI22_X1 U287 ( .A1(n306), .A2(n304), .B1(n302), .B2(n307), .ZN(n77) );
  OAI22_X1 U288 ( .A1(n307), .A2(n304), .B1(n302), .B2(n308), .ZN(n76) );
  XNOR2_X1 U289 ( .A(b[3]), .B(a[7]), .ZN(n307) );
  OAI22_X1 U290 ( .A1(n308), .A2(n304), .B1(n302), .B2(n309), .ZN(n75) );
  XNOR2_X1 U291 ( .A(b[4]), .B(a[7]), .ZN(n308) );
  OAI22_X1 U292 ( .A1(n309), .A2(n304), .B1(n302), .B2(n310), .ZN(n74) );
  XNOR2_X1 U293 ( .A(b[5]), .B(a[7]), .ZN(n309) );
  OAI22_X1 U294 ( .A1(n312), .A2(n302), .B1(n304), .B2(n312), .ZN(n311) );
  OAI21_X1 U295 ( .B1(n263), .B2(n261), .A(n277), .ZN(n72) );
  OAI21_X1 U296 ( .B1(n273), .B2(n283), .A(n313), .ZN(n71) );
  OR3_X1 U297 ( .A1(n281), .A2(n251), .A3(n273), .ZN(n313) );
  OAI21_X1 U298 ( .B1(n270), .B2(n293), .A(n314), .ZN(n70) );
  OR3_X1 U299 ( .A1(n291), .A2(n251), .A3(n270), .ZN(n314) );
  OAI21_X1 U300 ( .B1(n267), .B2(n304), .A(n315), .ZN(n69) );
  OR3_X1 U301 ( .A1(n302), .A2(n263), .A3(n267), .ZN(n315) );
  XNOR2_X1 U302 ( .A(n316), .B(n317), .ZN(n38) );
  OR2_X1 U303 ( .A1(n316), .A2(n317), .ZN(n37) );
  OAI22_X1 U304 ( .A1(n288), .A2(n283), .B1(n260), .B2(n318), .ZN(n317) );
  XNOR2_X1 U305 ( .A(b[5]), .B(a[3]), .ZN(n288) );
  OAI22_X1 U306 ( .A1(n305), .A2(n304), .B1(n302), .B2(n306), .ZN(n316) );
  XNOR2_X1 U307 ( .A(b[2]), .B(a[7]), .ZN(n306) );
  XNOR2_X1 U308 ( .A(b[1]), .B(a[7]), .ZN(n305) );
  OAI22_X1 U309 ( .A1(n318), .A2(n283), .B1(n260), .B2(n290), .ZN(n31) );
  XNOR2_X1 U310 ( .A(b[7]), .B(a[3]), .ZN(n290) );
  XNOR2_X1 U311 ( .A(n273), .B(a[2]), .ZN(n319) );
  XNOR2_X1 U312 ( .A(b[6]), .B(a[3]), .ZN(n318) );
  OAI22_X1 U313 ( .A1(n299), .A2(n293), .B1(n291), .B2(n301), .ZN(n21) );
  XNOR2_X1 U314 ( .A(b[7]), .B(a[5]), .ZN(n301) );
  XNOR2_X1 U315 ( .A(n270), .B(a[4]), .ZN(n320) );
  XNOR2_X1 U316 ( .A(b[6]), .B(a[5]), .ZN(n299) );
  OAI22_X1 U317 ( .A1(n310), .A2(n304), .B1(n302), .B2(n312), .ZN(n15) );
  XNOR2_X1 U318 ( .A(b[7]), .B(a[7]), .ZN(n312) );
  NAND2_X1 U319 ( .A1(n302), .A2(n321), .ZN(n304) );
  XNOR2_X1 U320 ( .A(n267), .B(a[6]), .ZN(n321) );
  XNOR2_X1 U321 ( .A(b[6]), .B(a[7]), .ZN(n310) );
  OAI22_X1 U322 ( .A1(n263), .A2(n277), .B1(n322), .B2(n275), .ZN(n104) );
  OAI22_X1 U323 ( .A1(n322), .A2(n277), .B1(n323), .B2(n275), .ZN(n103) );
  XNOR2_X1 U324 ( .A(b[1]), .B(n262), .ZN(n322) );
  OAI22_X1 U325 ( .A1(n323), .A2(n277), .B1(n324), .B2(n275), .ZN(n102) );
  XNOR2_X1 U326 ( .A(b[2]), .B(n262), .ZN(n323) );
  OAI22_X1 U327 ( .A1(n324), .A2(n277), .B1(n325), .B2(n275), .ZN(n101) );
  XNOR2_X1 U328 ( .A(b[3]), .B(n262), .ZN(n324) );
  OAI22_X1 U329 ( .A1(n325), .A2(n277), .B1(n276), .B2(n275), .ZN(n100) );
  XNOR2_X1 U330 ( .A(b[5]), .B(n262), .ZN(n276) );
  NAND2_X1 U331 ( .A1(a[1]), .A2(n275), .ZN(n277) );
  XNOR2_X1 U332 ( .A(b[4]), .B(n262), .ZN(n325) );
endmodule


module datapath_DW01_add_16 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n71;
  wire   [15:1] carry;

  FA_X1 U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n71), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[14]), .ZN(n65) );
  CLKBUF_X1 U2 ( .A(n13), .Z(n1) );
  XOR2_X1 U3 ( .A(B[3]), .B(A[3]), .Z(n2) );
  XOR2_X1 U4 ( .A(carry[3]), .B(n2), .Z(SUM[3]) );
  NAND2_X1 U5 ( .A1(carry[3]), .A2(B[3]), .ZN(n3) );
  NAND2_X1 U6 ( .A1(carry[3]), .A2(A[3]), .ZN(n4) );
  NAND2_X1 U7 ( .A1(B[3]), .A2(A[3]), .ZN(n5) );
  NAND3_X1 U8 ( .A1(n3), .A2(n4), .A3(n5), .ZN(carry[4]) );
  CLKBUF_X1 U9 ( .A(n21), .Z(n6) );
  NAND2_X1 U10 ( .A1(n21), .A2(B[13]), .ZN(n7) );
  XOR2_X1 U11 ( .A(B[4]), .B(A[4]), .Z(n8) );
  XOR2_X1 U12 ( .A(carry[4]), .B(n8), .Z(SUM[4]) );
  NAND2_X1 U13 ( .A1(carry[4]), .A2(B[4]), .ZN(n9) );
  NAND2_X1 U14 ( .A1(carry[4]), .A2(A[4]), .ZN(n10) );
  NAND2_X1 U15 ( .A1(B[4]), .A2(A[4]), .ZN(n11) );
  NAND3_X1 U16 ( .A1(n9), .A2(n10), .A3(n11), .ZN(carry[5]) );
  NAND3_X1 U17 ( .A1(n16), .A2(n17), .A3(n18), .ZN(n12) );
  NAND3_X1 U18 ( .A1(n64), .A2(n63), .A3(n62), .ZN(n13) );
  CLKBUF_X1 U19 ( .A(carry[7]), .Z(n14) );
  XOR2_X1 U20 ( .A(B[11]), .B(A[11]), .Z(n15) );
  XOR2_X1 U21 ( .A(n1), .B(n15), .Z(SUM[11]) );
  NAND2_X1 U22 ( .A1(n13), .A2(B[11]), .ZN(n16) );
  NAND2_X1 U23 ( .A1(carry[11]), .A2(A[11]), .ZN(n17) );
  NAND2_X1 U24 ( .A1(B[11]), .A2(A[11]), .ZN(n18) );
  NAND3_X1 U25 ( .A1(n16), .A2(n17), .A3(n18), .ZN(carry[12]) );
  NAND3_X1 U26 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n19) );
  NAND3_X1 U27 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n20) );
  NAND3_X1 U28 ( .A1(n23), .A2(n24), .A3(n25), .ZN(n21) );
  XOR2_X1 U29 ( .A(B[12]), .B(A[12]), .Z(n22) );
  XOR2_X1 U30 ( .A(n12), .B(n22), .Z(SUM[12]) );
  NAND2_X1 U31 ( .A1(n12), .A2(B[12]), .ZN(n23) );
  NAND2_X1 U32 ( .A1(carry[12]), .A2(A[12]), .ZN(n24) );
  NAND2_X1 U33 ( .A1(B[12]), .A2(A[12]), .ZN(n25) );
  NAND3_X1 U34 ( .A1(n23), .A2(n24), .A3(n25), .ZN(carry[13]) );
  XOR2_X1 U35 ( .A(B[5]), .B(A[5]), .Z(n26) );
  XOR2_X1 U36 ( .A(carry[5]), .B(n26), .Z(SUM[5]) );
  NAND2_X1 U37 ( .A1(carry[5]), .A2(B[5]), .ZN(n27) );
  NAND2_X1 U38 ( .A1(carry[5]), .A2(A[5]), .ZN(n28) );
  NAND2_X1 U39 ( .A1(B[5]), .A2(A[5]), .ZN(n29) );
  NAND3_X1 U40 ( .A1(n27), .A2(n28), .A3(n29), .ZN(carry[6]) );
  NAND3_X1 U41 ( .A1(n34), .A2(n33), .A3(n35), .ZN(n30) );
  CLKBUF_X1 U42 ( .A(n49), .Z(n31) );
  XOR2_X1 U43 ( .A(B[6]), .B(A[6]), .Z(n32) );
  XOR2_X1 U44 ( .A(n20), .B(n32), .Z(SUM[6]) );
  NAND2_X1 U45 ( .A1(n19), .A2(B[6]), .ZN(n33) );
  NAND2_X1 U46 ( .A1(carry[6]), .A2(A[6]), .ZN(n34) );
  NAND2_X1 U47 ( .A1(B[6]), .A2(A[6]), .ZN(n35) );
  NAND3_X1 U48 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[7]) );
  CLKBUF_X1 U49 ( .A(n60), .Z(n36) );
  NAND3_X1 U50 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n37) );
  NAND3_X1 U51 ( .A1(n48), .A2(n31), .A3(n50), .ZN(n38) );
  NAND3_X1 U52 ( .A1(n7), .A2(n43), .A3(n44), .ZN(n39) );
  NAND3_X1 U53 ( .A1(n7), .A2(n43), .A3(n44), .ZN(n40) );
  XOR2_X1 U54 ( .A(B[13]), .B(A[13]), .Z(n41) );
  XOR2_X1 U55 ( .A(n6), .B(n41), .Z(SUM[13]) );
  NAND2_X1 U56 ( .A1(n21), .A2(B[13]), .ZN(n42) );
  NAND2_X1 U57 ( .A1(carry[13]), .A2(A[13]), .ZN(n43) );
  NAND2_X1 U58 ( .A1(B[13]), .A2(A[13]), .ZN(n44) );
  NAND3_X1 U59 ( .A1(n42), .A2(n43), .A3(n44), .ZN(carry[14]) );
  NAND3_X1 U60 ( .A1(n60), .A2(n59), .A3(n58), .ZN(n45) );
  NAND3_X1 U61 ( .A1(n58), .A2(n59), .A3(n36), .ZN(n46) );
  XOR2_X1 U62 ( .A(B[7]), .B(A[7]), .Z(n47) );
  XOR2_X1 U63 ( .A(n14), .B(n47), .Z(SUM[7]) );
  NAND2_X1 U64 ( .A1(n30), .A2(B[7]), .ZN(n48) );
  NAND2_X1 U65 ( .A1(carry[7]), .A2(A[7]), .ZN(n49) );
  NAND2_X1 U66 ( .A1(B[7]), .A2(A[7]), .ZN(n50) );
  NAND3_X1 U67 ( .A1(n49), .A2(n48), .A3(n50), .ZN(carry[8]) );
  NAND3_X1 U68 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n51) );
  XOR2_X1 U69 ( .A(B[8]), .B(A[8]), .Z(n52) );
  XOR2_X1 U70 ( .A(n38), .B(n52), .Z(SUM[8]) );
  NAND2_X1 U71 ( .A1(n37), .A2(B[8]), .ZN(n53) );
  NAND2_X1 U72 ( .A1(carry[8]), .A2(A[8]), .ZN(n54) );
  NAND2_X1 U73 ( .A1(B[8]), .A2(A[8]), .ZN(n55) );
  NAND3_X1 U74 ( .A1(n53), .A2(n54), .A3(n55), .ZN(carry[9]) );
  XNOR2_X1 U75 ( .A(carry[15]), .B(n56), .ZN(SUM[15]) );
  XNOR2_X1 U76 ( .A(B[15]), .B(A[15]), .ZN(n56) );
  XOR2_X1 U77 ( .A(A[9]), .B(B[9]), .Z(n57) );
  XOR2_X1 U78 ( .A(carry[9]), .B(n57), .Z(SUM[9]) );
  NAND2_X1 U79 ( .A1(A[9]), .A2(B[9]), .ZN(n58) );
  NAND2_X1 U80 ( .A1(A[9]), .A2(n51), .ZN(n59) );
  NAND2_X1 U81 ( .A1(carry[9]), .A2(B[9]), .ZN(n60) );
  NAND3_X1 U82 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[10]) );
  XOR2_X1 U83 ( .A(A[10]), .B(B[10]), .Z(n61) );
  XOR2_X1 U84 ( .A(n61), .B(n46), .Z(SUM[10]) );
  NAND2_X1 U85 ( .A1(A[10]), .A2(B[10]), .ZN(n62) );
  NAND2_X1 U86 ( .A1(carry[10]), .A2(A[10]), .ZN(n63) );
  NAND2_X1 U87 ( .A1(B[10]), .A2(n45), .ZN(n64) );
  NAND3_X1 U88 ( .A1(n64), .A2(n63), .A3(n62), .ZN(carry[11]) );
  XNOR2_X1 U89 ( .A(B[14]), .B(n65), .ZN(n66) );
  XOR2_X1 U90 ( .A(n66), .B(n40), .Z(SUM[14]) );
  NAND2_X1 U91 ( .A1(B[14]), .A2(n39), .ZN(n67) );
  NAND2_X1 U92 ( .A1(carry[14]), .A2(A[14]), .ZN(n68) );
  NAND2_X1 U93 ( .A1(B[14]), .A2(A[14]), .ZN(n69) );
  NAND3_X1 U94 ( .A1(n67), .A2(n68), .A3(n69), .ZN(carry[15]) );
  XOR2_X1 U95 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U96 ( .A1(B[0]), .A2(A[0]), .ZN(n71) );
endmodule


module datapath_DW_mult_tc_15 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326;

  FA_X1 U10 ( .A(n46), .B(n49), .CI(n10), .CO(n9), .S(product[6]) );
  FA_X1 U11 ( .A(n50), .B(n53), .CI(n11), .CO(n10), .S(product[5]) );
  FA_X1 U12 ( .A(n54), .B(n206), .CI(n12), .CO(n11), .S(product[4]) );
  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n269), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n268), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n272), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n271), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n274), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  INV_X1 U157 ( .A(n15), .ZN(n265) );
  AND2_X1 U158 ( .A1(n213), .A2(n102), .ZN(n206) );
  XNOR2_X1 U159 ( .A(n266), .B(n15), .ZN(n207) );
  AND3_X1 U160 ( .A1(n249), .A2(n250), .A3(n251), .ZN(product[15]) );
  NAND3_X1 U161 ( .A1(n215), .A2(n216), .A3(n217), .ZN(n209) );
  NAND3_X1 U162 ( .A1(n221), .A2(n222), .A3(n223), .ZN(n210) );
  NAND3_X1 U163 ( .A1(n221), .A2(n222), .A3(n223), .ZN(n211) );
  XOR2_X1 U164 ( .A(a[3]), .B(n264), .Z(n283) );
  CLKBUF_X1 U165 ( .A(b[1]), .Z(n212) );
  XNOR2_X1 U166 ( .A(n209), .B(n207), .ZN(product[14]) );
  OAI22_X1 U167 ( .A1(n283), .A2(n284), .B1(n261), .B2(n285), .ZN(n213) );
  XOR2_X1 U168 ( .A(n17), .B(n265), .Z(n214) );
  XOR2_X1 U169 ( .A(n211), .B(n214), .Z(product[13]) );
  NAND2_X1 U170 ( .A1(n210), .A2(n17), .ZN(n215) );
  NAND2_X1 U171 ( .A1(n3), .A2(n265), .ZN(n216) );
  NAND2_X1 U172 ( .A1(n17), .A2(n265), .ZN(n217) );
  NAND3_X1 U173 ( .A1(n215), .A2(n216), .A3(n217), .ZN(n2) );
  NAND3_X1 U174 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n218) );
  NAND3_X1 U175 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n219) );
  XOR2_X1 U176 ( .A(n18), .B(n19), .Z(n220) );
  XOR2_X1 U177 ( .A(n219), .B(n220), .Z(product[12]) );
  NAND2_X1 U178 ( .A1(n218), .A2(n18), .ZN(n221) );
  NAND2_X1 U179 ( .A1(n4), .A2(n19), .ZN(n222) );
  NAND2_X1 U180 ( .A1(n18), .A2(n19), .ZN(n223) );
  NAND3_X1 U181 ( .A1(n221), .A2(n222), .A3(n223), .ZN(n3) );
  NAND3_X1 U182 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n224) );
  CLKBUF_X1 U183 ( .A(n14), .Z(n225) );
  NAND3_X1 U184 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n226) );
  NAND3_X1 U185 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n227) );
  XOR2_X1 U186 ( .A(n102), .B(n95), .Z(n56) );
  XOR2_X1 U187 ( .A(n40), .B(n45), .Z(n228) );
  XOR2_X1 U188 ( .A(n9), .B(n228), .Z(product[7]) );
  NAND2_X1 U189 ( .A1(n9), .A2(n40), .ZN(n229) );
  NAND2_X1 U190 ( .A1(n9), .A2(n45), .ZN(n230) );
  NAND2_X1 U191 ( .A1(n40), .A2(n45), .ZN(n231) );
  NAND3_X1 U192 ( .A1(n229), .A2(n230), .A3(n231), .ZN(n8) );
  NAND2_X2 U193 ( .A1(n282), .A2(n320), .ZN(n284) );
  XOR2_X1 U194 ( .A(n103), .B(n96), .Z(n232) );
  XOR2_X1 U195 ( .A(n225), .B(n232), .Z(product[2]) );
  NAND2_X1 U196 ( .A1(n14), .A2(n103), .ZN(n233) );
  NAND2_X1 U197 ( .A1(n14), .A2(n96), .ZN(n234) );
  NAND2_X1 U198 ( .A1(n103), .A2(n96), .ZN(n235) );
  NAND3_X1 U199 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n13) );
  NAND3_X1 U200 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n236) );
  XOR2_X1 U201 ( .A(n34), .B(n39), .Z(n237) );
  XOR2_X1 U202 ( .A(n8), .B(n237), .Z(product[8]) );
  NAND2_X1 U203 ( .A1(n226), .A2(n34), .ZN(n238) );
  NAND2_X1 U204 ( .A1(n226), .A2(n39), .ZN(n239) );
  NAND2_X1 U205 ( .A1(n34), .A2(n39), .ZN(n240) );
  NAND3_X1 U206 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n7) );
  INV_X1 U207 ( .A(n264), .ZN(n241) );
  NAND3_X1 U208 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n242) );
  NAND3_X1 U209 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n243) );
  XNOR2_X1 U210 ( .A(b[1]), .B(a[1]), .ZN(n244) );
  XOR2_X1 U211 ( .A(n33), .B(n28), .Z(n245) );
  XOR2_X1 U212 ( .A(n224), .B(n245), .Z(product[9]) );
  NAND2_X1 U213 ( .A1(n227), .A2(n33), .ZN(n246) );
  NAND2_X1 U214 ( .A1(n7), .A2(n28), .ZN(n247) );
  NAND2_X1 U215 ( .A1(n33), .A2(n28), .ZN(n248) );
  NAND3_X1 U216 ( .A1(n247), .A2(n246), .A3(n248), .ZN(n6) );
  NAND2_X1 U217 ( .A1(n2), .A2(n266), .ZN(n249) );
  NAND2_X1 U218 ( .A1(n2), .A2(n15), .ZN(n250) );
  NAND2_X1 U219 ( .A1(n266), .A2(n15), .ZN(n251) );
  NAND3_X1 U220 ( .A1(n256), .A2(n255), .A3(n254), .ZN(n252) );
  XOR2_X1 U221 ( .A(n24), .B(n27), .Z(n253) );
  XOR2_X1 U222 ( .A(n253), .B(n236), .Z(product[10]) );
  NAND2_X1 U223 ( .A1(n24), .A2(n27), .ZN(n254) );
  NAND2_X1 U224 ( .A1(n24), .A2(n6), .ZN(n255) );
  NAND2_X1 U225 ( .A1(n27), .A2(n243), .ZN(n256) );
  NAND3_X1 U226 ( .A1(n255), .A2(n254), .A3(n256), .ZN(n5) );
  XOR2_X1 U227 ( .A(n20), .B(n23), .Z(n257) );
  XOR2_X1 U228 ( .A(n257), .B(n242), .Z(product[11]) );
  NAND2_X1 U229 ( .A1(n20), .A2(n23), .ZN(n258) );
  NAND2_X1 U230 ( .A1(n20), .A2(n252), .ZN(n259) );
  NAND2_X1 U231 ( .A1(n23), .A2(n5), .ZN(n260) );
  NAND3_X1 U232 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n4) );
  XNOR2_X2 U233 ( .A(a[4]), .B(a[3]), .ZN(n292) );
  INV_X1 U234 ( .A(n21), .ZN(n268) );
  INV_X1 U235 ( .A(n301), .ZN(n269) );
  INV_X1 U236 ( .A(n312), .ZN(n266) );
  INV_X1 U237 ( .A(n281), .ZN(n274) );
  INV_X1 U238 ( .A(n290), .ZN(n272) );
  INV_X1 U239 ( .A(n31), .ZN(n271) );
  INV_X1 U240 ( .A(b[0]), .ZN(n264) );
  INV_X1 U241 ( .A(a[5]), .ZN(n270) );
  INV_X1 U242 ( .A(a[7]), .ZN(n267) );
  BUF_X1 U243 ( .A(n282), .Z(n261) );
  BUF_X1 U244 ( .A(n282), .Z(n262) );
  XNOR2_X1 U245 ( .A(a[2]), .B(a[1]), .ZN(n282) );
  INV_X1 U246 ( .A(a[3]), .ZN(n273) );
  NAND2_X2 U247 ( .A1(n292), .A2(n321), .ZN(n294) );
  INV_X1 U248 ( .A(a[1]), .ZN(n275) );
  XOR2_X2 U249 ( .A(a[6]), .B(n270), .Z(n303) );
  INV_X1 U250 ( .A(n264), .ZN(n263) );
  INV_X2 U251 ( .A(a[0]), .ZN(n276) );
  NOR2_X1 U252 ( .A1(n276), .A2(n264), .ZN(product[0]) );
  OAI22_X1 U253 ( .A1(n277), .A2(n278), .B1(n279), .B2(n276), .ZN(n99) );
  OAI22_X1 U254 ( .A1(n279), .A2(n278), .B1(n280), .B2(n276), .ZN(n98) );
  XNOR2_X1 U255 ( .A(b[6]), .B(a[1]), .ZN(n279) );
  OAI22_X1 U256 ( .A1(n276), .A2(n280), .B1(n278), .B2(n280), .ZN(n281) );
  XNOR2_X1 U257 ( .A(b[7]), .B(a[1]), .ZN(n280) );
  NOR2_X1 U258 ( .A1(n262), .A2(n264), .ZN(n96) );
  OAI22_X1 U259 ( .A1(n283), .A2(n284), .B1(n261), .B2(n285), .ZN(n95) );
  OAI22_X1 U260 ( .A1(n285), .A2(n284), .B1(n261), .B2(n286), .ZN(n94) );
  XNOR2_X1 U261 ( .A(b[1]), .B(a[3]), .ZN(n285) );
  OAI22_X1 U262 ( .A1(n286), .A2(n284), .B1(n261), .B2(n287), .ZN(n93) );
  XNOR2_X1 U263 ( .A(b[2]), .B(a[3]), .ZN(n286) );
  OAI22_X1 U264 ( .A1(n287), .A2(n284), .B1(n262), .B2(n288), .ZN(n92) );
  XNOR2_X1 U265 ( .A(a[3]), .B(b[3]), .ZN(n287) );
  OAI22_X1 U266 ( .A1(n288), .A2(n284), .B1(n262), .B2(n289), .ZN(n91) );
  XNOR2_X1 U267 ( .A(b[4]), .B(a[3]), .ZN(n288) );
  OAI22_X1 U268 ( .A1(n291), .A2(n261), .B1(n284), .B2(n291), .ZN(n290) );
  NOR2_X1 U269 ( .A1(n292), .A2(n264), .ZN(n88) );
  OAI22_X1 U270 ( .A1(n293), .A2(n294), .B1(n292), .B2(n295), .ZN(n87) );
  XNOR2_X1 U271 ( .A(a[5]), .B(n263), .ZN(n293) );
  OAI22_X1 U272 ( .A1(n295), .A2(n294), .B1(n292), .B2(n296), .ZN(n86) );
  XNOR2_X1 U273 ( .A(n212), .B(a[5]), .ZN(n295) );
  OAI22_X1 U274 ( .A1(n296), .A2(n294), .B1(n292), .B2(n297), .ZN(n85) );
  XNOR2_X1 U275 ( .A(b[2]), .B(a[5]), .ZN(n296) );
  OAI22_X1 U276 ( .A1(n297), .A2(n294), .B1(n292), .B2(n298), .ZN(n84) );
  XNOR2_X1 U277 ( .A(b[3]), .B(a[5]), .ZN(n297) );
  OAI22_X1 U278 ( .A1(n298), .A2(n294), .B1(n292), .B2(n299), .ZN(n83) );
  XNOR2_X1 U279 ( .A(b[4]), .B(a[5]), .ZN(n298) );
  OAI22_X1 U280 ( .A1(n299), .A2(n294), .B1(n292), .B2(n300), .ZN(n82) );
  XNOR2_X1 U281 ( .A(b[5]), .B(a[5]), .ZN(n299) );
  OAI22_X1 U282 ( .A1(n302), .A2(n292), .B1(n294), .B2(n302), .ZN(n301) );
  NOR2_X1 U283 ( .A1(n303), .A2(n264), .ZN(n80) );
  OAI22_X1 U284 ( .A1(n304), .A2(n305), .B1(n303), .B2(n306), .ZN(n79) );
  XNOR2_X1 U285 ( .A(a[7]), .B(n241), .ZN(n304) );
  OAI22_X1 U286 ( .A1(n307), .A2(n305), .B1(n303), .B2(n308), .ZN(n77) );
  OAI22_X1 U287 ( .A1(n308), .A2(n305), .B1(n303), .B2(n309), .ZN(n76) );
  XNOR2_X1 U288 ( .A(b[3]), .B(a[7]), .ZN(n308) );
  OAI22_X1 U289 ( .A1(n309), .A2(n305), .B1(n303), .B2(n310), .ZN(n75) );
  XNOR2_X1 U290 ( .A(b[4]), .B(a[7]), .ZN(n309) );
  OAI22_X1 U291 ( .A1(n310), .A2(n305), .B1(n303), .B2(n311), .ZN(n74) );
  XNOR2_X1 U292 ( .A(b[5]), .B(a[7]), .ZN(n310) );
  OAI22_X1 U293 ( .A1(n313), .A2(n303), .B1(n305), .B2(n313), .ZN(n312) );
  OAI21_X1 U294 ( .B1(n241), .B2(n275), .A(n278), .ZN(n72) );
  OAI21_X1 U295 ( .B1(n273), .B2(n284), .A(n314), .ZN(n71) );
  OR3_X1 U296 ( .A1(n262), .A2(n241), .A3(n273), .ZN(n314) );
  OAI21_X1 U297 ( .B1(n270), .B2(n294), .A(n315), .ZN(n70) );
  OR3_X1 U298 ( .A1(n292), .A2(n241), .A3(n270), .ZN(n315) );
  OAI21_X1 U299 ( .B1(n267), .B2(n305), .A(n316), .ZN(n69) );
  OR3_X1 U300 ( .A1(n303), .A2(n263), .A3(n267), .ZN(n316) );
  XNOR2_X1 U301 ( .A(n317), .B(n318), .ZN(n38) );
  OR2_X1 U302 ( .A1(n317), .A2(n318), .ZN(n37) );
  OAI22_X1 U303 ( .A1(n289), .A2(n284), .B1(n262), .B2(n319), .ZN(n318) );
  XNOR2_X1 U304 ( .A(b[5]), .B(a[3]), .ZN(n289) );
  OAI22_X1 U305 ( .A1(n306), .A2(n305), .B1(n303), .B2(n307), .ZN(n317) );
  XNOR2_X1 U306 ( .A(b[2]), .B(a[7]), .ZN(n307) );
  XNOR2_X1 U307 ( .A(n212), .B(a[7]), .ZN(n306) );
  OAI22_X1 U308 ( .A1(n319), .A2(n284), .B1(n261), .B2(n291), .ZN(n31) );
  XNOR2_X1 U309 ( .A(b[7]), .B(a[3]), .ZN(n291) );
  XNOR2_X1 U310 ( .A(n273), .B(a[2]), .ZN(n320) );
  XNOR2_X1 U311 ( .A(b[6]), .B(a[3]), .ZN(n319) );
  OAI22_X1 U312 ( .A1(n300), .A2(n294), .B1(n292), .B2(n302), .ZN(n21) );
  XNOR2_X1 U313 ( .A(b[7]), .B(a[5]), .ZN(n302) );
  XNOR2_X1 U314 ( .A(n270), .B(a[4]), .ZN(n321) );
  XNOR2_X1 U315 ( .A(b[6]), .B(a[5]), .ZN(n300) );
  OAI22_X1 U316 ( .A1(n311), .A2(n305), .B1(n303), .B2(n313), .ZN(n15) );
  XNOR2_X1 U317 ( .A(b[7]), .B(a[7]), .ZN(n313) );
  NAND2_X1 U318 ( .A1(n303), .A2(n322), .ZN(n305) );
  XNOR2_X1 U319 ( .A(n267), .B(a[6]), .ZN(n322) );
  XNOR2_X1 U320 ( .A(b[6]), .B(a[7]), .ZN(n311) );
  OAI22_X1 U321 ( .A1(n263), .A2(n278), .B1(n323), .B2(n276), .ZN(n104) );
  OAI22_X1 U322 ( .A1(n244), .A2(n278), .B1(n324), .B2(n276), .ZN(n103) );
  XNOR2_X1 U323 ( .A(b[1]), .B(a[1]), .ZN(n323) );
  OAI22_X1 U324 ( .A1(n324), .A2(n278), .B1(n325), .B2(n276), .ZN(n102) );
  XNOR2_X1 U325 ( .A(b[2]), .B(a[1]), .ZN(n324) );
  OAI22_X1 U326 ( .A1(n325), .A2(n278), .B1(n326), .B2(n276), .ZN(n101) );
  XNOR2_X1 U327 ( .A(b[3]), .B(a[1]), .ZN(n325) );
  OAI22_X1 U328 ( .A1(n326), .A2(n278), .B1(n277), .B2(n276), .ZN(n100) );
  XNOR2_X1 U329 ( .A(b[5]), .B(a[1]), .ZN(n277) );
  NAND2_X1 U330 ( .A1(a[1]), .A2(n276), .ZN(n278) );
  XNOR2_X1 U331 ( .A(b[4]), .B(a[1]), .ZN(n326) );
endmodule


module datapath_DW01_add_15 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n77;
  wire   [15:1] carry;

  FA_X1 U1_1 ( .A(A[1]), .B(n77), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[14]), .ZN(n71) );
  CLKBUF_X1 U2 ( .A(n46), .Z(n1) );
  CLKBUF_X1 U3 ( .A(B[13]), .Z(n2) );
  CLKBUF_X1 U4 ( .A(B[11]), .Z(n3) );
  XOR2_X1 U5 ( .A(carry[3]), .B(A[3]), .Z(n4) );
  XOR2_X1 U6 ( .A(B[3]), .B(n4), .Z(SUM[3]) );
  NAND2_X1 U7 ( .A1(B[3]), .A2(carry[3]), .ZN(n5) );
  NAND2_X1 U8 ( .A1(B[3]), .A2(A[3]), .ZN(n6) );
  NAND2_X1 U9 ( .A1(carry[3]), .A2(A[3]), .ZN(n7) );
  NAND3_X1 U10 ( .A1(n5), .A2(n6), .A3(n7), .ZN(carry[4]) );
  NAND3_X1 U11 ( .A1(n19), .A2(n20), .A3(n21), .ZN(n8) );
  NAND3_X1 U12 ( .A1(n19), .A2(n20), .A3(n21), .ZN(n9) );
  CLKBUF_X1 U13 ( .A(n44), .Z(n10) );
  CLKBUF_X1 U14 ( .A(n68), .Z(n11) );
  NAND3_X1 U15 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n12) );
  NAND3_X1 U16 ( .A1(n44), .A2(n45), .A3(n46), .ZN(n13) );
  NAND3_X1 U17 ( .A1(n10), .A2(n45), .A3(n1), .ZN(n14) );
  NAND3_X1 U18 ( .A1(n69), .A2(n68), .A3(n67), .ZN(n15) );
  NAND3_X1 U19 ( .A1(n69), .A2(n11), .A3(n67), .ZN(n16) );
  NAND2_X1 U20 ( .A1(B[8]), .A2(carry[8]), .ZN(n17) );
  XOR2_X1 U21 ( .A(carry[6]), .B(A[6]), .Z(n18) );
  XOR2_X1 U22 ( .A(B[6]), .B(n18), .Z(SUM[6]) );
  NAND2_X1 U23 ( .A1(B[6]), .A2(n12), .ZN(n19) );
  NAND2_X1 U24 ( .A1(B[6]), .A2(A[6]), .ZN(n20) );
  NAND2_X1 U25 ( .A1(carry[6]), .A2(A[6]), .ZN(n21) );
  NAND3_X1 U26 ( .A1(n19), .A2(n20), .A3(n21), .ZN(carry[7]) );
  CLKBUF_X1 U27 ( .A(n37), .Z(n22) );
  NAND3_X1 U28 ( .A1(n40), .A2(n41), .A3(n42), .ZN(n23) );
  XOR2_X1 U29 ( .A(B[4]), .B(A[4]), .Z(n24) );
  XOR2_X1 U30 ( .A(carry[4]), .B(n24), .Z(SUM[4]) );
  NAND2_X1 U31 ( .A1(carry[4]), .A2(B[4]), .ZN(n25) );
  NAND2_X1 U32 ( .A1(carry[4]), .A2(A[4]), .ZN(n26) );
  NAND2_X1 U33 ( .A1(B[4]), .A2(A[4]), .ZN(n27) );
  NAND3_X1 U34 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[5]) );
  XOR2_X1 U35 ( .A(B[5]), .B(A[5]), .Z(n28) );
  XOR2_X1 U36 ( .A(carry[5]), .B(n28), .Z(SUM[5]) );
  NAND2_X1 U37 ( .A1(carry[5]), .A2(B[5]), .ZN(n29) );
  NAND2_X1 U38 ( .A1(carry[5]), .A2(A[5]), .ZN(n30) );
  NAND2_X1 U39 ( .A1(B[5]), .A2(A[5]), .ZN(n31) );
  NAND3_X1 U40 ( .A1(n29), .A2(n30), .A3(n31), .ZN(carry[6]) );
  XOR2_X1 U41 ( .A(carry[2]), .B(A[2]), .Z(n32) );
  XOR2_X1 U42 ( .A(B[2]), .B(n32), .Z(SUM[2]) );
  NAND2_X1 U43 ( .A1(B[2]), .A2(carry[2]), .ZN(n33) );
  NAND2_X1 U44 ( .A1(B[2]), .A2(A[2]), .ZN(n34) );
  NAND2_X1 U45 ( .A1(carry[2]), .A2(A[2]), .ZN(n35) );
  NAND3_X1 U46 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[3]) );
  CLKBUF_X1 U47 ( .A(n23), .Z(n36) );
  NAND3_X1 U48 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n37) );
  NAND3_X1 U49 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n38) );
  XOR2_X1 U50 ( .A(B[10]), .B(A[10]), .Z(n39) );
  XOR2_X1 U51 ( .A(n16), .B(n39), .Z(SUM[10]) );
  NAND2_X1 U52 ( .A1(n15), .A2(B[10]), .ZN(n40) );
  NAND2_X1 U53 ( .A1(carry[10]), .A2(A[10]), .ZN(n41) );
  NAND2_X1 U54 ( .A1(B[10]), .A2(A[10]), .ZN(n42) );
  NAND3_X1 U55 ( .A1(n40), .A2(n41), .A3(n42), .ZN(carry[11]) );
  XOR2_X1 U56 ( .A(n3), .B(A[11]), .Z(n43) );
  XOR2_X1 U57 ( .A(n36), .B(n43), .Z(SUM[11]) );
  NAND2_X1 U58 ( .A1(n23), .A2(B[11]), .ZN(n44) );
  NAND2_X1 U59 ( .A1(carry[11]), .A2(A[11]), .ZN(n45) );
  NAND2_X1 U60 ( .A1(B[11]), .A2(A[11]), .ZN(n46) );
  NAND3_X1 U61 ( .A1(n44), .A2(n45), .A3(n46), .ZN(carry[12]) );
  XOR2_X1 U62 ( .A(B[12]), .B(A[12]), .Z(n47) );
  XOR2_X1 U63 ( .A(n14), .B(n47), .Z(SUM[12]) );
  NAND2_X1 U64 ( .A1(n13), .A2(B[12]), .ZN(n48) );
  NAND2_X1 U65 ( .A1(carry[12]), .A2(A[12]), .ZN(n49) );
  NAND2_X1 U66 ( .A1(B[12]), .A2(A[12]), .ZN(n50) );
  NAND3_X1 U67 ( .A1(n49), .A2(n48), .A3(n50), .ZN(carry[13]) );
  XOR2_X1 U68 ( .A(B[7]), .B(A[7]), .Z(n51) );
  XOR2_X1 U69 ( .A(n9), .B(n51), .Z(SUM[7]) );
  NAND2_X1 U70 ( .A1(n8), .A2(B[7]), .ZN(n52) );
  NAND2_X1 U71 ( .A1(carry[7]), .A2(A[7]), .ZN(n53) );
  NAND2_X1 U72 ( .A1(B[7]), .A2(A[7]), .ZN(n54) );
  NAND3_X1 U73 ( .A1(n52), .A2(n53), .A3(n54), .ZN(carry[8]) );
  NAND3_X1 U74 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n55) );
  NAND3_X1 U75 ( .A1(n65), .A2(n64), .A3(n63), .ZN(n56) );
  NAND3_X1 U76 ( .A1(n63), .A2(n64), .A3(n17), .ZN(n57) );
  XOR2_X1 U77 ( .A(n2), .B(A[13]), .Z(n58) );
  XOR2_X1 U78 ( .A(n22), .B(n58), .Z(SUM[13]) );
  NAND2_X1 U79 ( .A1(n37), .A2(B[13]), .ZN(n59) );
  NAND2_X1 U80 ( .A1(carry[13]), .A2(A[13]), .ZN(n60) );
  NAND2_X1 U81 ( .A1(B[13]), .A2(A[13]), .ZN(n61) );
  NAND3_X1 U82 ( .A1(n59), .A2(n60), .A3(n61), .ZN(carry[14]) );
  XOR2_X1 U83 ( .A(A[8]), .B(B[8]), .Z(n62) );
  XOR2_X1 U84 ( .A(n62), .B(n38), .Z(SUM[8]) );
  NAND2_X1 U85 ( .A1(A[8]), .A2(B[8]), .ZN(n63) );
  NAND2_X1 U86 ( .A1(carry[8]), .A2(A[8]), .ZN(n64) );
  NAND2_X1 U87 ( .A1(B[8]), .A2(n38), .ZN(n65) );
  NAND3_X1 U88 ( .A1(n17), .A2(n64), .A3(n63), .ZN(carry[9]) );
  XOR2_X1 U89 ( .A(A[9]), .B(B[9]), .Z(n66) );
  XOR2_X1 U90 ( .A(n66), .B(n57), .Z(SUM[9]) );
  NAND2_X1 U91 ( .A1(A[9]), .A2(B[9]), .ZN(n67) );
  NAND2_X1 U92 ( .A1(A[9]), .A2(n56), .ZN(n68) );
  NAND2_X1 U93 ( .A1(B[9]), .A2(carry[9]), .ZN(n69) );
  NAND3_X1 U94 ( .A1(n69), .A2(n68), .A3(n67), .ZN(carry[10]) );
  XNOR2_X1 U95 ( .A(carry[15]), .B(n70), .ZN(SUM[15]) );
  XNOR2_X1 U96 ( .A(B[15]), .B(A[15]), .ZN(n70) );
  XNOR2_X1 U97 ( .A(B[14]), .B(n71), .ZN(n72) );
  XOR2_X1 U98 ( .A(n72), .B(carry[14]), .Z(SUM[14]) );
  NAND2_X1 U99 ( .A1(n55), .A2(B[14]), .ZN(n73) );
  NAND2_X1 U100 ( .A1(n55), .A2(A[14]), .ZN(n74) );
  NAND2_X1 U101 ( .A1(B[14]), .A2(A[14]), .ZN(n75) );
  NAND3_X1 U102 ( .A1(n74), .A2(n73), .A3(n75), .ZN(carry[15]) );
  XOR2_X1 U103 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U104 ( .A1(B[0]), .A2(A[0]), .ZN(n77) );
endmodule


module datapath_DW_mult_tc_14 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340;

  FA_X1 U11 ( .A(n50), .B(n53), .CI(n11), .CO(n10), .S(product[5]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n284), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n283), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n287), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n286), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n289), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n207), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  CLKBUF_X3 U157 ( .A(a[1]), .Z(n206) );
  INV_X1 U158 ( .A(n279), .ZN(n278) );
  NAND2_X1 U159 ( .A1(n297), .A2(n335), .ZN(n299) );
  INV_X1 U160 ( .A(n15), .ZN(n280) );
  AND2_X1 U161 ( .A1(n70), .A2(n87), .ZN(n207) );
  XNOR2_X1 U162 ( .A(n281), .B(n15), .ZN(n208) );
  AND3_X1 U163 ( .A1(n216), .A2(n217), .A3(n218), .ZN(product[15]) );
  NAND3_X1 U164 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n210) );
  NAND3_X1 U165 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n211) );
  NAND3_X1 U166 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n212) );
  XOR2_X1 U167 ( .A(a[3]), .B(n279), .Z(n298) );
  CLKBUF_X1 U168 ( .A(n10), .Z(n222) );
  XNOR2_X1 U169 ( .A(n222), .B(n213), .ZN(product[6]) );
  XNOR2_X1 U170 ( .A(n46), .B(n49), .ZN(n213) );
  XNOR2_X1 U171 ( .A(a[4]), .B(a[3]), .ZN(n307) );
  XNOR2_X1 U172 ( .A(n2), .B(n208), .ZN(product[14]) );
  NAND3_X1 U173 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n214) );
  NAND3_X1 U174 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n215) );
  NAND2_X1 U175 ( .A1(n2), .A2(n281), .ZN(n216) );
  NAND2_X1 U176 ( .A1(n210), .A2(n15), .ZN(n217) );
  NAND2_X1 U177 ( .A1(n281), .A2(n15), .ZN(n218) );
  NAND3_X1 U178 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n219) );
  NAND3_X1 U179 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n220) );
  NAND3_X1 U180 ( .A1(n226), .A2(n227), .A3(n228), .ZN(n221) );
  NAND3_X1 U181 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n223) );
  NAND3_X1 U182 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n224) );
  XOR2_X1 U183 ( .A(n33), .B(n28), .Z(n225) );
  XOR2_X1 U184 ( .A(n220), .B(n225), .Z(product[9]) );
  NAND2_X1 U185 ( .A1(n219), .A2(n33), .ZN(n226) );
  NAND2_X1 U186 ( .A1(n7), .A2(n28), .ZN(n227) );
  NAND2_X1 U187 ( .A1(n33), .A2(n28), .ZN(n228) );
  NAND3_X1 U188 ( .A1(n226), .A2(n227), .A3(n228), .ZN(n6) );
  NAND3_X1 U189 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n229) );
  NAND3_X1 U190 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n230) );
  XOR2_X1 U191 ( .A(n27), .B(n24), .Z(n231) );
  XOR2_X1 U192 ( .A(n221), .B(n231), .Z(product[10]) );
  NAND2_X1 U193 ( .A1(n221), .A2(n27), .ZN(n232) );
  NAND2_X1 U194 ( .A1(n6), .A2(n24), .ZN(n233) );
  NAND2_X1 U195 ( .A1(n27), .A2(n24), .ZN(n234) );
  NAND3_X1 U196 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n5) );
  NAND3_X1 U197 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n235) );
  NAND2_X1 U198 ( .A1(n266), .A2(n267), .ZN(n236) );
  NAND2_X1 U199 ( .A1(n266), .A2(n267), .ZN(n237) );
  NAND2_X1 U200 ( .A1(n266), .A2(n267), .ZN(n297) );
  NAND2_X2 U201 ( .A1(n206), .A2(n291), .ZN(n293) );
  XNOR2_X1 U202 ( .A(n238), .B(n212), .ZN(product[3]) );
  XNOR2_X1 U203 ( .A(n56), .B(n71), .ZN(n238) );
  XOR2_X1 U204 ( .A(n23), .B(n20), .Z(n239) );
  XOR2_X1 U205 ( .A(n223), .B(n239), .Z(product[11]) );
  NAND2_X1 U206 ( .A1(n223), .A2(n23), .ZN(n240) );
  NAND2_X1 U207 ( .A1(n5), .A2(n20), .ZN(n241) );
  NAND2_X1 U208 ( .A1(n23), .A2(n20), .ZN(n242) );
  NAND3_X1 U209 ( .A1(n240), .A2(n241), .A3(n242), .ZN(n4) );
  NAND2_X1 U210 ( .A1(n10), .A2(n46), .ZN(n243) );
  NAND2_X1 U211 ( .A1(n10), .A2(n49), .ZN(n244) );
  NAND2_X1 U212 ( .A1(n46), .A2(n49), .ZN(n245) );
  NAND3_X1 U213 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n9) );
  XOR2_X1 U214 ( .A(n70), .B(n87), .Z(n52) );
  XOR2_X1 U215 ( .A(n40), .B(n45), .Z(n246) );
  XOR2_X1 U216 ( .A(n246), .B(n230), .Z(product[7]) );
  NAND2_X1 U217 ( .A1(n40), .A2(n45), .ZN(n247) );
  NAND2_X1 U218 ( .A1(n40), .A2(n9), .ZN(n248) );
  NAND2_X1 U219 ( .A1(n45), .A2(n9), .ZN(n249) );
  NAND3_X1 U220 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n8) );
  XOR2_X1 U221 ( .A(n34), .B(n39), .Z(n250) );
  XOR2_X1 U222 ( .A(n250), .B(n224), .Z(product[8]) );
  NAND2_X1 U223 ( .A1(n34), .A2(n39), .ZN(n251) );
  NAND2_X1 U224 ( .A1(n34), .A2(n8), .ZN(n252) );
  NAND2_X1 U225 ( .A1(n39), .A2(n8), .ZN(n253) );
  NAND3_X1 U226 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n7) );
  XOR2_X1 U227 ( .A(n103), .B(n96), .Z(n254) );
  XOR2_X1 U228 ( .A(n254), .B(n14), .Z(product[2]) );
  NAND2_X1 U229 ( .A1(n14), .A2(n103), .ZN(n255) );
  NAND2_X1 U230 ( .A1(n14), .A2(n96), .ZN(n256) );
  NAND2_X1 U231 ( .A1(n103), .A2(n96), .ZN(n257) );
  NAND3_X1 U232 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n13) );
  NAND2_X1 U233 ( .A1(n56), .A2(n71), .ZN(n258) );
  NAND2_X1 U234 ( .A1(n56), .A2(n211), .ZN(n259) );
  NAND2_X1 U235 ( .A1(n71), .A2(n13), .ZN(n260) );
  NAND3_X1 U236 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n12) );
  XOR2_X1 U237 ( .A(n54), .B(n55), .Z(n261) );
  XOR2_X1 U238 ( .A(n261), .B(n215), .Z(product[4]) );
  NAND2_X1 U239 ( .A1(n54), .A2(n55), .ZN(n262) );
  NAND2_X1 U240 ( .A1(n54), .A2(n214), .ZN(n263) );
  NAND2_X1 U241 ( .A1(n55), .A2(n12), .ZN(n264) );
  NAND3_X1 U242 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n11) );
  NAND2_X1 U243 ( .A1(a[2]), .A2(n206), .ZN(n266) );
  NAND2_X1 U244 ( .A1(n265), .A2(n290), .ZN(n267) );
  INV_X1 U245 ( .A(a[2]), .ZN(n265) );
  XOR2_X1 U246 ( .A(n18), .B(n19), .Z(n268) );
  XOR2_X1 U247 ( .A(n235), .B(n268), .Z(product[12]) );
  NAND2_X1 U248 ( .A1(n235), .A2(n18), .ZN(n269) );
  NAND2_X1 U249 ( .A1(n4), .A2(n19), .ZN(n270) );
  NAND2_X1 U250 ( .A1(n18), .A2(n19), .ZN(n271) );
  NAND3_X1 U251 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n3) );
  XOR2_X1 U252 ( .A(n17), .B(n280), .Z(n272) );
  XOR2_X1 U253 ( .A(n3), .B(n272), .Z(product[13]) );
  NAND2_X1 U254 ( .A1(n229), .A2(n17), .ZN(n273) );
  NAND2_X1 U255 ( .A1(n3), .A2(n280), .ZN(n274) );
  NAND2_X1 U256 ( .A1(n17), .A2(n280), .ZN(n275) );
  NAND3_X1 U257 ( .A1(n273), .A2(n274), .A3(n275), .ZN(n2) );
  NAND2_X1 U258 ( .A1(n307), .A2(n276), .ZN(n309) );
  XNOR2_X1 U259 ( .A(n285), .B(a[4]), .ZN(n276) );
  INV_X1 U260 ( .A(n21), .ZN(n283) );
  INV_X1 U261 ( .A(n316), .ZN(n284) );
  INV_X1 U262 ( .A(n327), .ZN(n281) );
  INV_X1 U263 ( .A(n296), .ZN(n289) );
  INV_X1 U264 ( .A(n305), .ZN(n287) );
  INV_X1 U265 ( .A(n31), .ZN(n286) );
  INV_X1 U266 ( .A(b[0]), .ZN(n279) );
  INV_X1 U267 ( .A(a[5]), .ZN(n285) );
  INV_X1 U268 ( .A(a[7]), .ZN(n282) );
  BUF_X2 U269 ( .A(n307), .Z(n277) );
  INV_X1 U270 ( .A(a[3]), .ZN(n288) );
  INV_X1 U271 ( .A(a[1]), .ZN(n290) );
  XOR2_X2 U272 ( .A(a[6]), .B(n285), .Z(n318) );
  INV_X2 U273 ( .A(a[0]), .ZN(n291) );
  NOR2_X1 U274 ( .A1(n291), .A2(n279), .ZN(product[0]) );
  OAI22_X1 U275 ( .A1(n292), .A2(n293), .B1(n294), .B2(n291), .ZN(n99) );
  OAI22_X1 U276 ( .A1(n294), .A2(n293), .B1(n295), .B2(n291), .ZN(n98) );
  XNOR2_X1 U277 ( .A(b[6]), .B(n206), .ZN(n294) );
  OAI22_X1 U278 ( .A1(n291), .A2(n295), .B1(n293), .B2(n295), .ZN(n296) );
  XNOR2_X1 U279 ( .A(b[7]), .B(n206), .ZN(n295) );
  NOR2_X1 U280 ( .A1(n237), .A2(n279), .ZN(n96) );
  OAI22_X1 U281 ( .A1(n298), .A2(n299), .B1(n236), .B2(n300), .ZN(n95) );
  OAI22_X1 U282 ( .A1(n300), .A2(n299), .B1(n237), .B2(n301), .ZN(n94) );
  XNOR2_X1 U283 ( .A(b[1]), .B(a[3]), .ZN(n300) );
  OAI22_X1 U284 ( .A1(n301), .A2(n299), .B1(n236), .B2(n302), .ZN(n93) );
  XNOR2_X1 U285 ( .A(b[2]), .B(a[3]), .ZN(n301) );
  OAI22_X1 U286 ( .A1(n302), .A2(n299), .B1(n237), .B2(n303), .ZN(n92) );
  XNOR2_X1 U287 ( .A(b[3]), .B(a[3]), .ZN(n302) );
  OAI22_X1 U288 ( .A1(n303), .A2(n299), .B1(n237), .B2(n304), .ZN(n91) );
  XNOR2_X1 U289 ( .A(b[4]), .B(a[3]), .ZN(n303) );
  OAI22_X1 U290 ( .A1(n306), .A2(n236), .B1(n299), .B2(n306), .ZN(n305) );
  NOR2_X1 U291 ( .A1(n277), .A2(n279), .ZN(n88) );
  OAI22_X1 U292 ( .A1(n308), .A2(n309), .B1(n277), .B2(n310), .ZN(n87) );
  XNOR2_X1 U293 ( .A(a[5]), .B(n278), .ZN(n308) );
  OAI22_X1 U294 ( .A1(n310), .A2(n309), .B1(n277), .B2(n311), .ZN(n86) );
  XNOR2_X1 U295 ( .A(b[1]), .B(a[5]), .ZN(n310) );
  OAI22_X1 U296 ( .A1(n311), .A2(n309), .B1(n277), .B2(n312), .ZN(n85) );
  XNOR2_X1 U297 ( .A(b[2]), .B(a[5]), .ZN(n311) );
  OAI22_X1 U298 ( .A1(n312), .A2(n309), .B1(n277), .B2(n313), .ZN(n84) );
  XNOR2_X1 U299 ( .A(b[3]), .B(a[5]), .ZN(n312) );
  OAI22_X1 U300 ( .A1(n313), .A2(n309), .B1(n277), .B2(n314), .ZN(n83) );
  XNOR2_X1 U301 ( .A(b[4]), .B(a[5]), .ZN(n313) );
  OAI22_X1 U302 ( .A1(n314), .A2(n309), .B1(n277), .B2(n315), .ZN(n82) );
  XNOR2_X1 U303 ( .A(b[5]), .B(a[5]), .ZN(n314) );
  OAI22_X1 U304 ( .A1(n317), .A2(n277), .B1(n309), .B2(n317), .ZN(n316) );
  NOR2_X1 U305 ( .A1(n318), .A2(n279), .ZN(n80) );
  OAI22_X1 U306 ( .A1(n319), .A2(n320), .B1(n318), .B2(n321), .ZN(n79) );
  XNOR2_X1 U307 ( .A(a[7]), .B(n278), .ZN(n319) );
  OAI22_X1 U308 ( .A1(n322), .A2(n320), .B1(n318), .B2(n323), .ZN(n77) );
  OAI22_X1 U309 ( .A1(n323), .A2(n320), .B1(n318), .B2(n324), .ZN(n76) );
  XNOR2_X1 U310 ( .A(b[3]), .B(a[7]), .ZN(n323) );
  OAI22_X1 U311 ( .A1(n324), .A2(n320), .B1(n318), .B2(n325), .ZN(n75) );
  XNOR2_X1 U312 ( .A(b[4]), .B(a[7]), .ZN(n324) );
  OAI22_X1 U313 ( .A1(n325), .A2(n320), .B1(n318), .B2(n326), .ZN(n74) );
  XNOR2_X1 U314 ( .A(b[5]), .B(a[7]), .ZN(n325) );
  OAI22_X1 U315 ( .A1(n328), .A2(n318), .B1(n320), .B2(n328), .ZN(n327) );
  OAI21_X1 U316 ( .B1(n278), .B2(n290), .A(n293), .ZN(n72) );
  OAI21_X1 U317 ( .B1(n288), .B2(n299), .A(n329), .ZN(n71) );
  OR3_X1 U318 ( .A1(n236), .A2(n278), .A3(n288), .ZN(n329) );
  OAI21_X1 U319 ( .B1(n285), .B2(n309), .A(n330), .ZN(n70) );
  OR3_X1 U320 ( .A1(n277), .A2(n278), .A3(n285), .ZN(n330) );
  OAI21_X1 U321 ( .B1(n282), .B2(n320), .A(n331), .ZN(n69) );
  OR3_X1 U322 ( .A1(n318), .A2(n278), .A3(n282), .ZN(n331) );
  XNOR2_X1 U323 ( .A(n332), .B(n333), .ZN(n38) );
  OR2_X1 U324 ( .A1(n332), .A2(n333), .ZN(n37) );
  OAI22_X1 U325 ( .A1(n304), .A2(n299), .B1(n237), .B2(n334), .ZN(n333) );
  XNOR2_X1 U326 ( .A(b[5]), .B(a[3]), .ZN(n304) );
  OAI22_X1 U327 ( .A1(n321), .A2(n320), .B1(n318), .B2(n322), .ZN(n332) );
  XNOR2_X1 U328 ( .A(b[2]), .B(a[7]), .ZN(n322) );
  XNOR2_X1 U329 ( .A(b[1]), .B(a[7]), .ZN(n321) );
  OAI22_X1 U330 ( .A1(n334), .A2(n299), .B1(n236), .B2(n306), .ZN(n31) );
  XNOR2_X1 U331 ( .A(b[7]), .B(a[3]), .ZN(n306) );
  XNOR2_X1 U332 ( .A(n288), .B(a[2]), .ZN(n335) );
  XNOR2_X1 U333 ( .A(b[6]), .B(a[3]), .ZN(n334) );
  OAI22_X1 U334 ( .A1(n315), .A2(n309), .B1(n277), .B2(n317), .ZN(n21) );
  XNOR2_X1 U335 ( .A(b[7]), .B(a[5]), .ZN(n317) );
  XNOR2_X1 U336 ( .A(b[6]), .B(a[5]), .ZN(n315) );
  OAI22_X1 U337 ( .A1(n326), .A2(n320), .B1(n318), .B2(n328), .ZN(n15) );
  XNOR2_X1 U338 ( .A(b[7]), .B(a[7]), .ZN(n328) );
  NAND2_X1 U339 ( .A1(n318), .A2(n336), .ZN(n320) );
  XNOR2_X1 U340 ( .A(n282), .B(a[6]), .ZN(n336) );
  XNOR2_X1 U341 ( .A(b[6]), .B(a[7]), .ZN(n326) );
  OAI22_X1 U342 ( .A1(n278), .A2(n293), .B1(n337), .B2(n291), .ZN(n104) );
  OAI22_X1 U343 ( .A1(n293), .A2(n337), .B1(n338), .B2(n291), .ZN(n103) );
  XNOR2_X1 U344 ( .A(b[1]), .B(n206), .ZN(n337) );
  OAI22_X1 U345 ( .A1(n338), .A2(n293), .B1(n339), .B2(n291), .ZN(n102) );
  XNOR2_X1 U346 ( .A(b[2]), .B(n206), .ZN(n338) );
  OAI22_X1 U347 ( .A1(n339), .A2(n293), .B1(n340), .B2(n291), .ZN(n101) );
  XNOR2_X1 U348 ( .A(b[3]), .B(n206), .ZN(n339) );
  OAI22_X1 U349 ( .A1(n340), .A2(n293), .B1(n292), .B2(n291), .ZN(n100) );
  XNOR2_X1 U350 ( .A(b[5]), .B(n206), .ZN(n292) );
  XNOR2_X1 U351 ( .A(b[4]), .B(n206), .ZN(n340) );
endmodule


module datapath_DW01_add_14 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n72;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n72), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(carry[4]), .Z(n1) );
  NAND3_X1 U2 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n2) );
  NAND3_X1 U3 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n3) );
  XOR2_X1 U4 ( .A(B[2]), .B(A[2]), .Z(n4) );
  XOR2_X1 U5 ( .A(carry[2]), .B(n4), .Z(SUM[2]) );
  NAND2_X1 U6 ( .A1(carry[2]), .A2(B[2]), .ZN(n5) );
  NAND2_X1 U7 ( .A1(carry[2]), .A2(A[2]), .ZN(n6) );
  NAND2_X1 U8 ( .A1(B[2]), .A2(A[2]), .ZN(n7) );
  NAND3_X1 U9 ( .A1(n5), .A2(n6), .A3(n7), .ZN(carry[3]) );
  CLKBUF_X1 U10 ( .A(n33), .Z(n8) );
  XOR2_X1 U11 ( .A(B[3]), .B(A[3]), .Z(n9) );
  XOR2_X1 U12 ( .A(carry[3]), .B(n9), .Z(SUM[3]) );
  NAND2_X1 U13 ( .A1(carry[3]), .A2(B[3]), .ZN(n10) );
  NAND2_X1 U14 ( .A1(carry[3]), .A2(A[3]), .ZN(n11) );
  NAND2_X1 U15 ( .A1(B[3]), .A2(A[3]), .ZN(n12) );
  NAND3_X1 U16 ( .A1(n10), .A2(n11), .A3(n12), .ZN(carry[4]) );
  XOR2_X1 U17 ( .A(B[4]), .B(A[4]), .Z(n13) );
  XOR2_X1 U18 ( .A(n1), .B(n13), .Z(SUM[4]) );
  NAND2_X1 U19 ( .A1(carry[4]), .A2(B[4]), .ZN(n14) );
  NAND2_X1 U20 ( .A1(carry[4]), .A2(A[4]), .ZN(n15) );
  NAND2_X1 U21 ( .A1(B[4]), .A2(A[4]), .ZN(n16) );
  NAND3_X1 U22 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[5]) );
  NAND2_X1 U23 ( .A1(carry[10]), .A2(A[10]), .ZN(n17) );
  NAND3_X1 U24 ( .A1(n32), .A2(n33), .A3(n34), .ZN(n18) );
  NAND3_X1 U25 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n19) );
  NAND2_X1 U26 ( .A1(n50), .A2(A[11]), .ZN(n20) );
  CLKBUF_X1 U27 ( .A(n44), .Z(n21) );
  NAND2_X1 U28 ( .A1(n44), .A2(B[10]), .ZN(n22) );
  CLKBUF_X1 U29 ( .A(n22), .Z(n23) );
  XOR2_X1 U30 ( .A(n3), .B(A[5]), .Z(n24) );
  XOR2_X1 U31 ( .A(B[5]), .B(n24), .Z(SUM[5]) );
  NAND2_X1 U32 ( .A1(B[5]), .A2(n2), .ZN(n25) );
  NAND2_X1 U33 ( .A1(B[5]), .A2(A[5]), .ZN(n26) );
  NAND2_X1 U34 ( .A1(carry[5]), .A2(A[5]), .ZN(n27) );
  NAND3_X1 U35 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[6]) );
  NAND3_X1 U36 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n28) );
  NAND3_X1 U37 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n29) );
  NAND3_X1 U38 ( .A1(n23), .A2(n17), .A3(n56), .ZN(n30) );
  XOR2_X1 U39 ( .A(B[6]), .B(A[6]), .Z(n31) );
  XOR2_X1 U40 ( .A(carry[6]), .B(n31), .Z(SUM[6]) );
  NAND2_X1 U41 ( .A1(n19), .A2(B[6]), .ZN(n32) );
  NAND2_X1 U42 ( .A1(n19), .A2(A[6]), .ZN(n33) );
  NAND2_X1 U43 ( .A1(B[6]), .A2(A[6]), .ZN(n34) );
  NAND3_X1 U44 ( .A1(n32), .A2(n8), .A3(n34), .ZN(carry[7]) );
  NAND3_X1 U45 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n35) );
  XOR2_X1 U46 ( .A(B[7]), .B(A[7]), .Z(n36) );
  XOR2_X1 U47 ( .A(carry[7]), .B(n36), .Z(SUM[7]) );
  NAND2_X1 U48 ( .A1(n18), .A2(B[7]), .ZN(n37) );
  NAND2_X1 U49 ( .A1(n18), .A2(A[7]), .ZN(n38) );
  NAND2_X1 U50 ( .A1(B[7]), .A2(A[7]), .ZN(n39) );
  NAND3_X1 U51 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[8]) );
  XOR2_X1 U52 ( .A(B[8]), .B(A[8]), .Z(n40) );
  XOR2_X1 U53 ( .A(n35), .B(n40), .Z(SUM[8]) );
  NAND2_X1 U54 ( .A1(n35), .A2(B[8]), .ZN(n41) );
  NAND2_X1 U55 ( .A1(carry[8]), .A2(A[8]), .ZN(n42) );
  NAND2_X1 U56 ( .A1(B[8]), .A2(A[8]), .ZN(n43) );
  NAND3_X1 U57 ( .A1(n41), .A2(n42), .A3(n43), .ZN(carry[9]) );
  NAND3_X1 U58 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n44) );
  XOR2_X1 U59 ( .A(B[9]), .B(A[9]), .Z(n45) );
  XOR2_X1 U60 ( .A(n29), .B(n45), .Z(SUM[9]) );
  NAND2_X1 U61 ( .A1(n28), .A2(B[9]), .ZN(n46) );
  NAND2_X1 U62 ( .A1(carry[9]), .A2(A[9]), .ZN(n47) );
  NAND2_X1 U63 ( .A1(B[9]), .A2(A[9]), .ZN(n48) );
  NAND3_X1 U64 ( .A1(n47), .A2(n46), .A3(n48), .ZN(carry[10]) );
  XNOR2_X1 U65 ( .A(carry[15]), .B(n49), .ZN(SUM[15]) );
  XNOR2_X1 U66 ( .A(B[15]), .B(A[15]), .ZN(n49) );
  NAND3_X1 U67 ( .A1(n22), .A2(n17), .A3(n56), .ZN(n50) );
  NAND3_X1 U68 ( .A1(n66), .A2(n65), .A3(n64), .ZN(n51) );
  CLKBUF_X1 U69 ( .A(n20), .Z(n52) );
  XOR2_X1 U70 ( .A(B[10]), .B(A[10]), .Z(n53) );
  XOR2_X1 U71 ( .A(n21), .B(n53), .Z(SUM[10]) );
  NAND2_X1 U72 ( .A1(n44), .A2(B[10]), .ZN(n54) );
  NAND2_X1 U73 ( .A1(carry[10]), .A2(A[10]), .ZN(n55) );
  NAND2_X1 U74 ( .A1(B[10]), .A2(A[10]), .ZN(n56) );
  NAND3_X1 U75 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[11]) );
  NAND3_X1 U76 ( .A1(n61), .A2(n60), .A3(n62), .ZN(n57) );
  NAND3_X1 U77 ( .A1(n60), .A2(n52), .A3(n62), .ZN(n58) );
  XOR2_X1 U78 ( .A(B[11]), .B(A[11]), .Z(n59) );
  XOR2_X1 U79 ( .A(n30), .B(n59), .Z(SUM[11]) );
  NAND2_X1 U80 ( .A1(carry[11]), .A2(B[11]), .ZN(n60) );
  NAND2_X1 U81 ( .A1(n50), .A2(A[11]), .ZN(n61) );
  NAND2_X1 U82 ( .A1(B[11]), .A2(A[11]), .ZN(n62) );
  NAND3_X1 U83 ( .A1(n20), .A2(n60), .A3(n62), .ZN(carry[12]) );
  NAND2_X1 U84 ( .A1(A[12]), .A2(B[12]), .ZN(n64) );
  XOR2_X1 U85 ( .A(A[12]), .B(B[12]), .Z(n63) );
  XOR2_X1 U86 ( .A(n63), .B(n58), .Z(SUM[12]) );
  NAND2_X1 U87 ( .A1(A[12]), .A2(n57), .ZN(n65) );
  NAND2_X1 U88 ( .A1(carry[12]), .A2(B[12]), .ZN(n66) );
  NAND3_X1 U89 ( .A1(n66), .A2(n65), .A3(n64), .ZN(carry[13]) );
  XOR2_X1 U90 ( .A(A[13]), .B(B[13]), .Z(n67) );
  XOR2_X1 U91 ( .A(n67), .B(carry[13]), .Z(SUM[13]) );
  NAND2_X1 U92 ( .A1(A[13]), .A2(B[13]), .ZN(n68) );
  NAND2_X1 U93 ( .A1(n51), .A2(A[13]), .ZN(n69) );
  NAND2_X1 U94 ( .A1(B[13]), .A2(carry[13]), .ZN(n70) );
  NAND3_X1 U95 ( .A1(n70), .A2(n69), .A3(n68), .ZN(carry[14]) );
  XOR2_X1 U96 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U97 ( .A1(B[0]), .A2(A[0]), .ZN(n72) );
endmodule


module datapath_DW_mult_tc_13 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74,
         n75, n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92,
         n93, n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332;

  FA_X1 U11 ( .A(n50), .B(n53), .CI(n11), .CO(n10), .S(product[5]) );
  FA_X1 U12 ( .A(n54), .B(n55), .CI(n12), .CO(n11), .S(product[4]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n275), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n274), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n278), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n277), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n280), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  INV_X1 U157 ( .A(n15), .ZN(n271) );
  AND3_X1 U158 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n229) );
  XNOR2_X1 U159 ( .A(n272), .B(n15), .ZN(n206) );
  AND3_X1 U160 ( .A1(n232), .A2(n233), .A3(n234), .ZN(product[15]) );
  XOR2_X1 U161 ( .A(n229), .B(n230), .Z(product[10]) );
  NAND3_X1 U162 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n208) );
  XOR2_X1 U163 ( .A(n209), .B(n210), .Z(product[3]) );
  XNOR2_X1 U164 ( .A(n56), .B(n71), .ZN(n209) );
  AND3_X1 U165 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n210) );
  NAND3_X1 U166 ( .A1(n214), .A2(n215), .A3(n216), .ZN(n211) );
  NAND3_X1 U167 ( .A1(n214), .A2(n215), .A3(n216), .ZN(n212) );
  XOR2_X1 U168 ( .A(n46), .B(n49), .Z(n213) );
  XOR2_X1 U169 ( .A(n10), .B(n213), .Z(product[6]) );
  NAND2_X1 U170 ( .A1(n10), .A2(n46), .ZN(n214) );
  NAND2_X1 U171 ( .A1(n10), .A2(n49), .ZN(n215) );
  NAND2_X1 U172 ( .A1(n46), .A2(n49), .ZN(n216) );
  NAND3_X1 U173 ( .A1(n214), .A2(n215), .A3(n216), .ZN(n9) );
  NAND3_X1 U174 ( .A1(n219), .A2(n220), .A3(n221), .ZN(n217) );
  XNOR2_X1 U175 ( .A(n2), .B(n206), .ZN(product[14]) );
  XOR2_X1 U176 ( .A(n40), .B(n45), .Z(n218) );
  XOR2_X1 U177 ( .A(n212), .B(n218), .Z(product[7]) );
  NAND2_X1 U178 ( .A1(n211), .A2(n40), .ZN(n219) );
  NAND2_X1 U179 ( .A1(n9), .A2(n45), .ZN(n220) );
  NAND2_X1 U180 ( .A1(n40), .A2(n45), .ZN(n221) );
  NAND3_X1 U181 ( .A1(n219), .A2(n220), .A3(n221), .ZN(n8) );
  NAND3_X1 U182 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n222) );
  NAND3_X1 U183 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n223) );
  XOR2_X1 U184 ( .A(n17), .B(n271), .Z(n224) );
  XOR2_X1 U185 ( .A(n223), .B(n224), .Z(product[13]) );
  NAND2_X1 U186 ( .A1(n222), .A2(n17), .ZN(n225) );
  NAND2_X1 U187 ( .A1(n3), .A2(n271), .ZN(n226) );
  NAND2_X1 U188 ( .A1(n17), .A2(n271), .ZN(n227) );
  NAND3_X1 U189 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n2) );
  NAND2_X1 U190 ( .A1(n298), .A2(n327), .ZN(n228) );
  NAND2_X1 U191 ( .A1(n298), .A2(n327), .ZN(n300) );
  XNOR2_X1 U192 ( .A(n27), .B(n24), .ZN(n230) );
  CLKBUF_X1 U193 ( .A(b[1]), .Z(n231) );
  NAND2_X1 U194 ( .A1(n208), .A2(n272), .ZN(n232) );
  NAND2_X1 U195 ( .A1(n208), .A2(n15), .ZN(n233) );
  NAND2_X1 U196 ( .A1(n272), .A2(n15), .ZN(n234) );
  XNOR2_X2 U197 ( .A(a[2]), .B(a[1]), .ZN(n235) );
  XNOR2_X1 U198 ( .A(a[2]), .B(a[1]), .ZN(n288) );
  INV_X2 U199 ( .A(n270), .ZN(n269) );
  NAND3_X1 U200 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n236) );
  XOR2_X1 U201 ( .A(n34), .B(n39), .Z(n237) );
  XOR2_X1 U202 ( .A(n217), .B(n237), .Z(product[8]) );
  NAND2_X1 U203 ( .A1(n217), .A2(n34), .ZN(n238) );
  NAND2_X1 U204 ( .A1(n8), .A2(n39), .ZN(n239) );
  NAND2_X1 U205 ( .A1(n34), .A2(n39), .ZN(n240) );
  NAND3_X1 U206 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n7) );
  AND2_X1 U207 ( .A1(n104), .A2(n72), .ZN(n241) );
  NAND3_X1 U208 ( .A1(n259), .A2(n258), .A3(n260), .ZN(n242) );
  NAND3_X1 U209 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n243) );
  NAND3_X1 U210 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n244) );
  XOR2_X1 U211 ( .A(n95), .B(n102), .Z(n245) );
  XOR2_X1 U212 ( .A(n33), .B(n28), .Z(n246) );
  XOR2_X1 U213 ( .A(n236), .B(n246), .Z(product[9]) );
  NAND2_X1 U214 ( .A1(n236), .A2(n33), .ZN(n247) );
  NAND2_X1 U215 ( .A1(n7), .A2(n28), .ZN(n248) );
  NAND2_X1 U216 ( .A1(n33), .A2(n28), .ZN(n249) );
  NAND3_X1 U217 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n6) );
  NAND3_X1 U218 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n250) );
  XOR2_X1 U219 ( .A(n103), .B(n96), .Z(n251) );
  XOR2_X1 U220 ( .A(n251), .B(n241), .Z(product[2]) );
  NAND2_X1 U221 ( .A1(n103), .A2(n96), .ZN(n252) );
  NAND2_X1 U222 ( .A1(n103), .A2(n241), .ZN(n253) );
  NAND2_X1 U223 ( .A1(n96), .A2(n14), .ZN(n254) );
  NAND3_X1 U224 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n13) );
  NAND2_X1 U225 ( .A1(n245), .A2(n71), .ZN(n255) );
  NAND2_X1 U226 ( .A1(n245), .A2(n250), .ZN(n256) );
  NAND2_X1 U227 ( .A1(n71), .A2(n13), .ZN(n257) );
  NAND3_X1 U228 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n12) );
  NAND2_X1 U229 ( .A1(n6), .A2(n27), .ZN(n258) );
  NAND2_X1 U230 ( .A1(n244), .A2(n24), .ZN(n259) );
  NAND2_X1 U231 ( .A1(n27), .A2(n24), .ZN(n260) );
  NAND3_X1 U232 ( .A1(n258), .A2(n259), .A3(n260), .ZN(n5) );
  XNOR2_X2 U233 ( .A(a[4]), .B(a[3]), .ZN(n298) );
  XOR2_X1 U234 ( .A(n20), .B(n23), .Z(n261) );
  XOR2_X1 U235 ( .A(n261), .B(n242), .Z(product[11]) );
  NAND2_X1 U236 ( .A1(n20), .A2(n23), .ZN(n262) );
  NAND2_X1 U237 ( .A1(n20), .A2(n5), .ZN(n263) );
  NAND2_X1 U238 ( .A1(n23), .A2(n5), .ZN(n264) );
  NAND3_X1 U239 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n4) );
  XOR2_X1 U240 ( .A(n19), .B(n18), .Z(n265) );
  XOR2_X1 U241 ( .A(n265), .B(n243), .Z(product[12]) );
  NAND2_X1 U242 ( .A1(n19), .A2(n18), .ZN(n266) );
  NAND2_X1 U243 ( .A1(n19), .A2(n4), .ZN(n267) );
  NAND2_X1 U244 ( .A1(n18), .A2(n4), .ZN(n268) );
  NAND3_X1 U245 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n3) );
  INV_X1 U246 ( .A(n21), .ZN(n274) );
  INV_X1 U247 ( .A(n307), .ZN(n275) );
  INV_X1 U248 ( .A(n318), .ZN(n272) );
  INV_X1 U249 ( .A(n287), .ZN(n280) );
  INV_X1 U250 ( .A(n296), .ZN(n278) );
  INV_X1 U251 ( .A(n31), .ZN(n277) );
  INV_X1 U252 ( .A(b[0]), .ZN(n270) );
  INV_X1 U253 ( .A(a[5]), .ZN(n276) );
  INV_X1 U254 ( .A(a[7]), .ZN(n273) );
  INV_X1 U255 ( .A(a[3]), .ZN(n279) );
  NAND2_X2 U256 ( .A1(n288), .A2(n326), .ZN(n290) );
  INV_X1 U257 ( .A(a[1]), .ZN(n281) );
  XOR2_X2 U258 ( .A(a[6]), .B(n276), .Z(n309) );
  INV_X2 U259 ( .A(a[0]), .ZN(n282) );
  NOR2_X1 U260 ( .A1(n282), .A2(n270), .ZN(product[0]) );
  OAI22_X1 U261 ( .A1(n283), .A2(n284), .B1(n285), .B2(n282), .ZN(n99) );
  OAI22_X1 U262 ( .A1(n285), .A2(n284), .B1(n286), .B2(n282), .ZN(n98) );
  XNOR2_X1 U263 ( .A(b[6]), .B(a[1]), .ZN(n285) );
  OAI22_X1 U264 ( .A1(n282), .A2(n286), .B1(n284), .B2(n286), .ZN(n287) );
  XNOR2_X1 U265 ( .A(b[7]), .B(a[1]), .ZN(n286) );
  NOR2_X1 U266 ( .A1(n235), .A2(n270), .ZN(n96) );
  OAI22_X1 U267 ( .A1(n289), .A2(n290), .B1(n235), .B2(n291), .ZN(n95) );
  XNOR2_X1 U268 ( .A(a[3]), .B(n269), .ZN(n289) );
  OAI22_X1 U269 ( .A1(n291), .A2(n290), .B1(n235), .B2(n292), .ZN(n94) );
  XNOR2_X1 U270 ( .A(b[1]), .B(a[3]), .ZN(n291) );
  OAI22_X1 U271 ( .A1(n292), .A2(n290), .B1(n235), .B2(n293), .ZN(n93) );
  XNOR2_X1 U272 ( .A(b[2]), .B(a[3]), .ZN(n292) );
  OAI22_X1 U273 ( .A1(n293), .A2(n290), .B1(n235), .B2(n294), .ZN(n92) );
  XNOR2_X1 U274 ( .A(b[3]), .B(a[3]), .ZN(n293) );
  OAI22_X1 U275 ( .A1(n294), .A2(n290), .B1(n235), .B2(n295), .ZN(n91) );
  XNOR2_X1 U276 ( .A(b[4]), .B(a[3]), .ZN(n294) );
  OAI22_X1 U277 ( .A1(n297), .A2(n235), .B1(n290), .B2(n297), .ZN(n296) );
  NOR2_X1 U278 ( .A1(n298), .A2(n270), .ZN(n88) );
  OAI22_X1 U279 ( .A1(n299), .A2(n300), .B1(n298), .B2(n301), .ZN(n87) );
  XNOR2_X1 U280 ( .A(a[5]), .B(n269), .ZN(n299) );
  OAI22_X1 U281 ( .A1(n301), .A2(n228), .B1(n298), .B2(n302), .ZN(n86) );
  XNOR2_X1 U282 ( .A(b[1]), .B(a[5]), .ZN(n301) );
  OAI22_X1 U283 ( .A1(n302), .A2(n228), .B1(n298), .B2(n303), .ZN(n85) );
  XNOR2_X1 U284 ( .A(b[2]), .B(a[5]), .ZN(n302) );
  OAI22_X1 U285 ( .A1(n303), .A2(n228), .B1(n298), .B2(n304), .ZN(n84) );
  XNOR2_X1 U286 ( .A(b[3]), .B(a[5]), .ZN(n303) );
  OAI22_X1 U287 ( .A1(n304), .A2(n228), .B1(n298), .B2(n305), .ZN(n83) );
  XNOR2_X1 U288 ( .A(b[4]), .B(a[5]), .ZN(n304) );
  OAI22_X1 U289 ( .A1(n305), .A2(n228), .B1(n298), .B2(n306), .ZN(n82) );
  XNOR2_X1 U290 ( .A(b[5]), .B(a[5]), .ZN(n305) );
  OAI22_X1 U291 ( .A1(n308), .A2(n298), .B1(n228), .B2(n308), .ZN(n307) );
  NOR2_X1 U292 ( .A1(n309), .A2(n270), .ZN(n80) );
  OAI22_X1 U293 ( .A1(n310), .A2(n311), .B1(n309), .B2(n312), .ZN(n79) );
  XNOR2_X1 U294 ( .A(a[7]), .B(n269), .ZN(n310) );
  OAI22_X1 U295 ( .A1(n313), .A2(n311), .B1(n309), .B2(n314), .ZN(n77) );
  OAI22_X1 U296 ( .A1(n314), .A2(n311), .B1(n309), .B2(n315), .ZN(n76) );
  XNOR2_X1 U297 ( .A(b[3]), .B(a[7]), .ZN(n314) );
  OAI22_X1 U298 ( .A1(n315), .A2(n311), .B1(n309), .B2(n316), .ZN(n75) );
  XNOR2_X1 U299 ( .A(b[4]), .B(a[7]), .ZN(n315) );
  OAI22_X1 U300 ( .A1(n316), .A2(n311), .B1(n309), .B2(n317), .ZN(n74) );
  XNOR2_X1 U301 ( .A(b[5]), .B(a[7]), .ZN(n316) );
  OAI22_X1 U302 ( .A1(n319), .A2(n309), .B1(n311), .B2(n319), .ZN(n318) );
  OAI21_X1 U303 ( .B1(n269), .B2(n281), .A(n284), .ZN(n72) );
  OAI21_X1 U304 ( .B1(n279), .B2(n290), .A(n320), .ZN(n71) );
  OR3_X1 U305 ( .A1(n235), .A2(n269), .A3(n279), .ZN(n320) );
  OAI21_X1 U306 ( .B1(n276), .B2(n300), .A(n321), .ZN(n70) );
  OR3_X1 U307 ( .A1(n298), .A2(n269), .A3(n276), .ZN(n321) );
  OAI21_X1 U308 ( .B1(n273), .B2(n311), .A(n322), .ZN(n69) );
  OR3_X1 U309 ( .A1(n309), .A2(n269), .A3(n273), .ZN(n322) );
  XNOR2_X1 U310 ( .A(n323), .B(n324), .ZN(n38) );
  OR2_X1 U311 ( .A1(n323), .A2(n324), .ZN(n37) );
  OAI22_X1 U312 ( .A1(n295), .A2(n290), .B1(n235), .B2(n325), .ZN(n324) );
  XNOR2_X1 U313 ( .A(b[5]), .B(a[3]), .ZN(n295) );
  OAI22_X1 U314 ( .A1(n312), .A2(n311), .B1(n309), .B2(n313), .ZN(n323) );
  XNOR2_X1 U315 ( .A(b[2]), .B(a[7]), .ZN(n313) );
  XNOR2_X1 U316 ( .A(n231), .B(a[7]), .ZN(n312) );
  OAI22_X1 U317 ( .A1(n325), .A2(n290), .B1(n235), .B2(n297), .ZN(n31) );
  XNOR2_X1 U318 ( .A(b[7]), .B(a[3]), .ZN(n297) );
  XNOR2_X1 U319 ( .A(n279), .B(a[2]), .ZN(n326) );
  XNOR2_X1 U320 ( .A(b[6]), .B(a[3]), .ZN(n325) );
  OAI22_X1 U321 ( .A1(n306), .A2(n228), .B1(n298), .B2(n308), .ZN(n21) );
  XNOR2_X1 U322 ( .A(b[7]), .B(a[5]), .ZN(n308) );
  XNOR2_X1 U323 ( .A(n276), .B(a[4]), .ZN(n327) );
  XNOR2_X1 U324 ( .A(b[6]), .B(a[5]), .ZN(n306) );
  OAI22_X1 U325 ( .A1(n317), .A2(n311), .B1(n309), .B2(n319), .ZN(n15) );
  XNOR2_X1 U326 ( .A(b[7]), .B(a[7]), .ZN(n319) );
  NAND2_X1 U327 ( .A1(n309), .A2(n328), .ZN(n311) );
  XNOR2_X1 U328 ( .A(n273), .B(a[6]), .ZN(n328) );
  XNOR2_X1 U329 ( .A(b[6]), .B(a[7]), .ZN(n317) );
  OAI22_X1 U330 ( .A1(n269), .A2(n284), .B1(n329), .B2(n282), .ZN(n104) );
  OAI22_X1 U331 ( .A1(n284), .A2(n329), .B1(n330), .B2(n282), .ZN(n103) );
  XNOR2_X1 U332 ( .A(b[1]), .B(a[1]), .ZN(n329) );
  OAI22_X1 U333 ( .A1(n330), .A2(n284), .B1(n331), .B2(n282), .ZN(n102) );
  XNOR2_X1 U334 ( .A(b[2]), .B(a[1]), .ZN(n330) );
  OAI22_X1 U335 ( .A1(n331), .A2(n284), .B1(n332), .B2(n282), .ZN(n101) );
  XNOR2_X1 U336 ( .A(b[3]), .B(a[1]), .ZN(n331) );
  OAI22_X1 U337 ( .A1(n332), .A2(n284), .B1(n283), .B2(n282), .ZN(n100) );
  XNOR2_X1 U338 ( .A(b[5]), .B(a[1]), .ZN(n283) );
  NAND2_X1 U339 ( .A1(a[1]), .A2(n282), .ZN(n284) );
  XNOR2_X1 U340 ( .A(b[4]), .B(a[1]), .ZN(n332) );
endmodule


module datapath_DW01_add_13 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n70;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n70), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND3_X1 U1 ( .A1(n6), .A2(n7), .A3(n8), .ZN(n1) );
  NAND3_X1 U2 ( .A1(n6), .A2(n7), .A3(n8), .ZN(n2) );
  CLKBUF_X1 U3 ( .A(n59), .Z(n3) );
  CLKBUF_X1 U4 ( .A(n64), .Z(n4) );
  XOR2_X1 U5 ( .A(B[3]), .B(A[3]), .Z(n5) );
  XOR2_X1 U6 ( .A(carry[3]), .B(n5), .Z(SUM[3]) );
  NAND2_X1 U7 ( .A1(carry[3]), .A2(B[3]), .ZN(n6) );
  NAND2_X1 U8 ( .A1(carry[3]), .A2(A[3]), .ZN(n7) );
  NAND2_X1 U9 ( .A1(B[3]), .A2(A[3]), .ZN(n8) );
  NAND3_X1 U10 ( .A1(n6), .A2(n7), .A3(n8), .ZN(carry[4]) );
  NAND3_X1 U11 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n9) );
  NAND3_X1 U12 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n10) );
  NAND3_X1 U13 ( .A1(n58), .A2(n3), .A3(n60), .ZN(n11) );
  NAND3_X1 U14 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n12) );
  XOR2_X1 U15 ( .A(B[11]), .B(A[11]), .Z(n13) );
  XOR2_X1 U16 ( .A(n11), .B(n13), .Z(SUM[11]) );
  NAND2_X1 U17 ( .A1(n10), .A2(B[11]), .ZN(n14) );
  NAND2_X1 U18 ( .A1(carry[11]), .A2(A[11]), .ZN(n15) );
  NAND2_X1 U19 ( .A1(B[11]), .A2(A[11]), .ZN(n16) );
  NAND3_X1 U20 ( .A1(n15), .A2(n14), .A3(n16), .ZN(carry[12]) );
  NAND3_X1 U21 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n17) );
  CLKBUF_X1 U22 ( .A(n31), .Z(n18) );
  NAND3_X1 U23 ( .A1(n36), .A2(n37), .A3(n38), .ZN(n19) );
  XOR2_X1 U24 ( .A(B[4]), .B(A[4]), .Z(n20) );
  XOR2_X1 U25 ( .A(n2), .B(n20), .Z(SUM[4]) );
  NAND2_X1 U26 ( .A1(n1), .A2(B[4]), .ZN(n21) );
  NAND2_X1 U27 ( .A1(carry[4]), .A2(A[4]), .ZN(n22) );
  NAND2_X1 U28 ( .A1(B[4]), .A2(A[4]), .ZN(n23) );
  NAND3_X1 U29 ( .A1(n21), .A2(n22), .A3(n23), .ZN(carry[5]) );
  NAND3_X1 U30 ( .A1(n50), .A2(n51), .A3(n52), .ZN(n24) );
  CLKBUF_X1 U31 ( .A(carry[6]), .Z(n25) );
  CLKBUF_X1 U32 ( .A(n63), .Z(n26) );
  CLKBUF_X1 U33 ( .A(n17), .Z(n27) );
  NAND3_X1 U34 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n28) );
  CLKBUF_X1 U35 ( .A(n24), .Z(n29) );
  XNOR2_X1 U36 ( .A(carry[15]), .B(n30), .ZN(SUM[15]) );
  XNOR2_X1 U37 ( .A(B[15]), .B(A[15]), .ZN(n30) );
  NAND3_X1 U38 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n31) );
  CLKBUF_X1 U39 ( .A(carry[9]), .Z(n32) );
  NAND3_X1 U40 ( .A1(n64), .A2(n63), .A3(n62), .ZN(n33) );
  NAND3_X1 U41 ( .A1(n4), .A2(n26), .A3(n62), .ZN(n34) );
  XOR2_X1 U42 ( .A(B[5]), .B(A[5]), .Z(n35) );
  XOR2_X1 U43 ( .A(n12), .B(n35), .Z(SUM[5]) );
  NAND2_X1 U44 ( .A1(n12), .A2(B[5]), .ZN(n36) );
  NAND2_X1 U45 ( .A1(carry[5]), .A2(A[5]), .ZN(n37) );
  NAND2_X1 U46 ( .A1(B[5]), .A2(A[5]), .ZN(n38) );
  NAND3_X1 U47 ( .A1(n36), .A2(n37), .A3(n38), .ZN(carry[6]) );
  NAND3_X1 U48 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n39) );
  XOR2_X1 U49 ( .A(B[8]), .B(A[8]), .Z(n40) );
  XOR2_X1 U50 ( .A(n29), .B(n40), .Z(SUM[8]) );
  NAND2_X1 U51 ( .A1(n24), .A2(B[8]), .ZN(n41) );
  NAND2_X1 U52 ( .A1(carry[8]), .A2(A[8]), .ZN(n42) );
  NAND2_X1 U53 ( .A1(B[8]), .A2(A[8]), .ZN(n43) );
  NAND3_X1 U54 ( .A1(n41), .A2(n42), .A3(n43), .ZN(carry[9]) );
  XOR2_X1 U55 ( .A(B[6]), .B(A[6]), .Z(n44) );
  XOR2_X1 U56 ( .A(n25), .B(n44), .Z(SUM[6]) );
  NAND2_X1 U57 ( .A1(n19), .A2(B[6]), .ZN(n45) );
  NAND2_X1 U58 ( .A1(carry[6]), .A2(A[6]), .ZN(n46) );
  NAND2_X1 U59 ( .A1(B[6]), .A2(A[6]), .ZN(n47) );
  CLKBUF_X1 U60 ( .A(n9), .Z(n48) );
  NAND2_X1 U61 ( .A1(A[12]), .A2(B[12]), .ZN(n62) );
  XOR2_X1 U62 ( .A(B[7]), .B(A[7]), .Z(n49) );
  XOR2_X1 U63 ( .A(n27), .B(n49), .Z(SUM[7]) );
  NAND2_X1 U64 ( .A1(n17), .A2(B[7]), .ZN(n50) );
  NAND2_X1 U65 ( .A1(n39), .A2(A[7]), .ZN(n51) );
  NAND2_X1 U66 ( .A1(B[7]), .A2(A[7]), .ZN(n52) );
  NAND3_X1 U67 ( .A1(n50), .A2(n51), .A3(n52), .ZN(carry[8]) );
  XOR2_X1 U68 ( .A(B[9]), .B(A[9]), .Z(n53) );
  XOR2_X1 U69 ( .A(n32), .B(n53), .Z(SUM[9]) );
  NAND2_X1 U70 ( .A1(n28), .A2(B[9]), .ZN(n54) );
  NAND2_X1 U71 ( .A1(carry[9]), .A2(A[9]), .ZN(n55) );
  NAND2_X1 U72 ( .A1(B[9]), .A2(A[9]), .ZN(n56) );
  NAND3_X1 U73 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[10]) );
  XOR2_X1 U74 ( .A(B[10]), .B(A[10]), .Z(n57) );
  XOR2_X1 U75 ( .A(n18), .B(n57), .Z(SUM[10]) );
  NAND2_X1 U76 ( .A1(carry[10]), .A2(B[10]), .ZN(n58) );
  NAND2_X1 U77 ( .A1(n31), .A2(A[10]), .ZN(n59) );
  NAND2_X1 U78 ( .A1(B[10]), .A2(A[10]), .ZN(n60) );
  NAND3_X1 U79 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[11]) );
  XOR2_X1 U80 ( .A(A[12]), .B(B[12]), .Z(n61) );
  XOR2_X1 U81 ( .A(n61), .B(n48), .Z(SUM[12]) );
  NAND2_X1 U82 ( .A1(A[12]), .A2(carry[12]), .ZN(n63) );
  NAND2_X1 U83 ( .A1(n9), .A2(B[12]), .ZN(n64) );
  NAND3_X1 U84 ( .A1(n64), .A2(n63), .A3(n62), .ZN(carry[13]) );
  XOR2_X1 U85 ( .A(A[13]), .B(B[13]), .Z(n65) );
  XOR2_X1 U86 ( .A(n65), .B(n34), .Z(SUM[13]) );
  NAND2_X1 U87 ( .A1(A[13]), .A2(B[13]), .ZN(n66) );
  NAND2_X1 U88 ( .A1(A[13]), .A2(n33), .ZN(n67) );
  NAND2_X1 U89 ( .A1(B[13]), .A2(carry[13]), .ZN(n68) );
  NAND3_X1 U90 ( .A1(n66), .A2(n67), .A3(n68), .ZN(carry[14]) );
  XOR2_X1 U91 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U92 ( .A1(B[0]), .A2(A[0]), .ZN(n70) );
endmodule


module datapath_DW_mult_tc_12 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333;

  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n277), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n276), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n280), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n279), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n282), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  INV_X1 U157 ( .A(n15), .ZN(n273) );
  XNOR2_X1 U158 ( .A(n274), .B(n15), .ZN(n206) );
  AND3_X1 U159 ( .A1(n266), .A2(n265), .A3(n267), .ZN(product[15]) );
  NAND3_X1 U160 ( .A1(n227), .A2(n228), .A3(n229), .ZN(n208) );
  NAND3_X1 U161 ( .A1(n227), .A2(n228), .A3(n229), .ZN(n209) );
  NAND3_X1 U162 ( .A1(n223), .A2(n224), .A3(n225), .ZN(n210) );
  NAND3_X1 U163 ( .A1(n216), .A2(n217), .A3(n218), .ZN(n211) );
  NAND3_X1 U164 ( .A1(n216), .A2(n217), .A3(n218), .ZN(n212) );
  NAND3_X1 U165 ( .A1(n246), .A2(n245), .A3(n244), .ZN(n213) );
  NAND3_X1 U166 ( .A1(n246), .A2(n245), .A3(n244), .ZN(n214) );
  XOR2_X1 U167 ( .A(n34), .B(n39), .Z(n215) );
  XOR2_X1 U168 ( .A(n209), .B(n215), .Z(product[8]) );
  NAND2_X1 U169 ( .A1(n8), .A2(n34), .ZN(n216) );
  NAND2_X1 U170 ( .A1(n208), .A2(n39), .ZN(n217) );
  NAND2_X1 U171 ( .A1(n34), .A2(n39), .ZN(n218) );
  NAND3_X1 U172 ( .A1(n217), .A2(n216), .A3(n218), .ZN(n7) );
  NAND3_X1 U173 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n219) );
  XNOR2_X1 U174 ( .A(n220), .B(n252), .ZN(product[11]) );
  XNOR2_X1 U175 ( .A(n20), .B(n23), .ZN(n220) );
  NAND3_X1 U176 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n221) );
  XOR2_X1 U177 ( .A(n54), .B(n55), .Z(n222) );
  XOR2_X1 U178 ( .A(n12), .B(n222), .Z(product[4]) );
  NAND2_X1 U179 ( .A1(n12), .A2(n54), .ZN(n223) );
  NAND2_X1 U180 ( .A1(n12), .A2(n55), .ZN(n224) );
  NAND2_X1 U181 ( .A1(n54), .A2(n55), .ZN(n225) );
  NAND3_X1 U182 ( .A1(n223), .A2(n224), .A3(n225), .ZN(n11) );
  XOR2_X1 U183 ( .A(n40), .B(n45), .Z(n226) );
  XOR2_X1 U184 ( .A(n219), .B(n226), .Z(product[7]) );
  NAND2_X1 U185 ( .A1(n219), .A2(n40), .ZN(n227) );
  NAND2_X1 U186 ( .A1(n9), .A2(n45), .ZN(n228) );
  NAND2_X1 U187 ( .A1(n40), .A2(n45), .ZN(n229) );
  NAND3_X1 U188 ( .A1(n227), .A2(n228), .A3(n229), .ZN(n8) );
  XNOR2_X1 U189 ( .A(n2), .B(n206), .ZN(product[14]) );
  NAND3_X1 U190 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n230) );
  NAND3_X1 U191 ( .A1(n234), .A2(n235), .A3(n236), .ZN(n231) );
  NAND3_X1 U192 ( .A1(n234), .A2(n235), .A3(n236), .ZN(n232) );
  XOR2_X1 U193 ( .A(n18), .B(n19), .Z(n233) );
  XOR2_X1 U194 ( .A(n230), .B(n233), .Z(product[12]) );
  NAND2_X1 U195 ( .A1(n230), .A2(n18), .ZN(n234) );
  NAND2_X1 U196 ( .A1(n4), .A2(n19), .ZN(n235) );
  NAND2_X1 U197 ( .A1(n18), .A2(n19), .ZN(n236) );
  NAND3_X1 U198 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n237) );
  CLKBUF_X1 U199 ( .A(n330), .Z(n242) );
  XOR2_X1 U200 ( .A(n33), .B(n28), .Z(n238) );
  XOR2_X1 U201 ( .A(n212), .B(n238), .Z(product[9]) );
  NAND2_X1 U202 ( .A1(n211), .A2(n33), .ZN(n239) );
  NAND2_X1 U203 ( .A1(n7), .A2(n28), .ZN(n240) );
  NAND2_X1 U204 ( .A1(n33), .A2(n28), .ZN(n241) );
  NAND3_X1 U205 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n6) );
  XOR2_X1 U206 ( .A(n50), .B(n53), .Z(n243) );
  XOR2_X1 U207 ( .A(n243), .B(n210), .Z(product[5]) );
  NAND2_X1 U208 ( .A1(n50), .A2(n53), .ZN(n244) );
  NAND2_X1 U209 ( .A1(n50), .A2(n11), .ZN(n245) );
  NAND2_X1 U210 ( .A1(n53), .A2(n210), .ZN(n246) );
  NAND3_X1 U211 ( .A1(n246), .A2(n245), .A3(n244), .ZN(n10) );
  XOR2_X1 U212 ( .A(n46), .B(n49), .Z(n247) );
  XOR2_X1 U213 ( .A(n247), .B(n214), .Z(product[6]) );
  NAND2_X1 U214 ( .A1(n46), .A2(n49), .ZN(n248) );
  NAND2_X1 U215 ( .A1(n46), .A2(n213), .ZN(n249) );
  NAND2_X1 U216 ( .A1(n49), .A2(n10), .ZN(n250) );
  NAND3_X1 U217 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n9) );
  NAND3_X1 U218 ( .A1(n255), .A2(n256), .A3(n254), .ZN(n251) );
  NAND3_X1 U219 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n252) );
  XOR2_X1 U220 ( .A(n24), .B(n27), .Z(n253) );
  XOR2_X1 U221 ( .A(n253), .B(n6), .Z(product[10]) );
  NAND2_X1 U222 ( .A1(n24), .A2(n27), .ZN(n254) );
  NAND2_X1 U223 ( .A1(n24), .A2(n6), .ZN(n255) );
  NAND2_X1 U224 ( .A1(n27), .A2(n237), .ZN(n256) );
  NAND3_X1 U225 ( .A1(n255), .A2(n254), .A3(n256), .ZN(n5) );
  NAND2_X1 U226 ( .A1(n20), .A2(n23), .ZN(n257) );
  NAND2_X1 U227 ( .A1(n20), .A2(n251), .ZN(n258) );
  NAND2_X1 U228 ( .A1(n23), .A2(n5), .ZN(n259) );
  NAND3_X1 U229 ( .A1(n257), .A2(n258), .A3(n259), .ZN(n4) );
  XOR2_X1 U230 ( .A(n17), .B(n273), .Z(n260) );
  XOR2_X1 U231 ( .A(n232), .B(n260), .Z(product[13]) );
  NAND2_X1 U232 ( .A1(n231), .A2(n17), .ZN(n261) );
  NAND2_X1 U233 ( .A1(n231), .A2(n273), .ZN(n262) );
  NAND2_X1 U234 ( .A1(n17), .A2(n273), .ZN(n263) );
  NAND3_X1 U235 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n2) );
  INV_X1 U236 ( .A(n272), .ZN(n264) );
  NAND2_X1 U237 ( .A1(n221), .A2(n274), .ZN(n265) );
  NAND2_X1 U238 ( .A1(n221), .A2(n15), .ZN(n266) );
  NAND2_X1 U239 ( .A1(n274), .A2(n15), .ZN(n267) );
  XNOR2_X2 U240 ( .A(a[4]), .B(a[3]), .ZN(n299) );
  BUF_X2 U241 ( .A(n289), .Z(n268) );
  XOR2_X1 U242 ( .A(a[2]), .B(n269), .Z(n289) );
  INV_X1 U243 ( .A(n21), .ZN(n276) );
  INV_X1 U244 ( .A(n308), .ZN(n277) );
  INV_X1 U245 ( .A(n319), .ZN(n274) );
  INV_X1 U246 ( .A(n288), .ZN(n282) );
  INV_X1 U247 ( .A(n297), .ZN(n280) );
  INV_X1 U248 ( .A(n31), .ZN(n279) );
  INV_X1 U249 ( .A(b[0]), .ZN(n272) );
  INV_X1 U250 ( .A(a[5]), .ZN(n278) );
  INV_X1 U251 ( .A(a[7]), .ZN(n275) );
  INV_X1 U252 ( .A(a[3]), .ZN(n281) );
  NAND2_X2 U253 ( .A1(n299), .A2(n328), .ZN(n301) );
  INV_X1 U254 ( .A(a[1]), .ZN(n269) );
  INV_X2 U255 ( .A(n269), .ZN(n270) );
  NAND2_X2 U256 ( .A1(n289), .A2(n327), .ZN(n291) );
  XOR2_X2 U257 ( .A(a[6]), .B(n278), .Z(n310) );
  INV_X1 U258 ( .A(n272), .ZN(n271) );
  INV_X2 U259 ( .A(a[0]), .ZN(n283) );
  NOR2_X1 U260 ( .A1(n283), .A2(n272), .ZN(product[0]) );
  OAI22_X1 U261 ( .A1(n284), .A2(n285), .B1(n286), .B2(n283), .ZN(n99) );
  OAI22_X1 U262 ( .A1(n286), .A2(n285), .B1(n287), .B2(n283), .ZN(n98) );
  XNOR2_X1 U263 ( .A(b[6]), .B(n270), .ZN(n286) );
  OAI22_X1 U264 ( .A1(n283), .A2(n287), .B1(n285), .B2(n287), .ZN(n288) );
  XNOR2_X1 U265 ( .A(b[7]), .B(n270), .ZN(n287) );
  NOR2_X1 U266 ( .A1(n289), .A2(n272), .ZN(n96) );
  OAI22_X1 U267 ( .A1(n290), .A2(n291), .B1(n289), .B2(n292), .ZN(n95) );
  XNOR2_X1 U268 ( .A(a[3]), .B(n271), .ZN(n290) );
  OAI22_X1 U269 ( .A1(n292), .A2(n291), .B1(n268), .B2(n293), .ZN(n94) );
  XNOR2_X1 U270 ( .A(b[1]), .B(a[3]), .ZN(n292) );
  OAI22_X1 U271 ( .A1(n293), .A2(n291), .B1(n268), .B2(n294), .ZN(n93) );
  XNOR2_X1 U272 ( .A(b[2]), .B(a[3]), .ZN(n293) );
  OAI22_X1 U273 ( .A1(n294), .A2(n291), .B1(n268), .B2(n295), .ZN(n92) );
  XNOR2_X1 U274 ( .A(b[3]), .B(a[3]), .ZN(n294) );
  OAI22_X1 U275 ( .A1(n295), .A2(n291), .B1(n268), .B2(n296), .ZN(n91) );
  XNOR2_X1 U276 ( .A(b[4]), .B(a[3]), .ZN(n295) );
  OAI22_X1 U277 ( .A1(n298), .A2(n268), .B1(n291), .B2(n298), .ZN(n297) );
  NOR2_X1 U278 ( .A1(n299), .A2(n272), .ZN(n88) );
  OAI22_X1 U279 ( .A1(n300), .A2(n301), .B1(n299), .B2(n302), .ZN(n87) );
  XNOR2_X1 U280 ( .A(a[5]), .B(n271), .ZN(n300) );
  OAI22_X1 U281 ( .A1(n302), .A2(n301), .B1(n299), .B2(n303), .ZN(n86) );
  XNOR2_X1 U282 ( .A(b[1]), .B(a[5]), .ZN(n302) );
  OAI22_X1 U283 ( .A1(n303), .A2(n301), .B1(n299), .B2(n304), .ZN(n85) );
  XNOR2_X1 U284 ( .A(b[2]), .B(a[5]), .ZN(n303) );
  OAI22_X1 U285 ( .A1(n304), .A2(n301), .B1(n299), .B2(n305), .ZN(n84) );
  XNOR2_X1 U286 ( .A(b[3]), .B(a[5]), .ZN(n304) );
  OAI22_X1 U287 ( .A1(n305), .A2(n301), .B1(n299), .B2(n306), .ZN(n83) );
  XNOR2_X1 U288 ( .A(b[4]), .B(a[5]), .ZN(n305) );
  OAI22_X1 U289 ( .A1(n306), .A2(n301), .B1(n299), .B2(n307), .ZN(n82) );
  XNOR2_X1 U290 ( .A(b[5]), .B(a[5]), .ZN(n306) );
  OAI22_X1 U291 ( .A1(n309), .A2(n299), .B1(n301), .B2(n309), .ZN(n308) );
  NOR2_X1 U292 ( .A1(n310), .A2(n272), .ZN(n80) );
  OAI22_X1 U293 ( .A1(n311), .A2(n312), .B1(n310), .B2(n313), .ZN(n79) );
  XNOR2_X1 U294 ( .A(a[7]), .B(n264), .ZN(n311) );
  OAI22_X1 U295 ( .A1(n314), .A2(n312), .B1(n310), .B2(n315), .ZN(n77) );
  OAI22_X1 U296 ( .A1(n315), .A2(n312), .B1(n310), .B2(n316), .ZN(n76) );
  XNOR2_X1 U297 ( .A(b[3]), .B(a[7]), .ZN(n315) );
  OAI22_X1 U298 ( .A1(n316), .A2(n312), .B1(n310), .B2(n317), .ZN(n75) );
  XNOR2_X1 U299 ( .A(b[4]), .B(a[7]), .ZN(n316) );
  OAI22_X1 U300 ( .A1(n317), .A2(n312), .B1(n310), .B2(n318), .ZN(n74) );
  XNOR2_X1 U301 ( .A(b[5]), .B(a[7]), .ZN(n317) );
  OAI22_X1 U302 ( .A1(n320), .A2(n310), .B1(n312), .B2(n320), .ZN(n319) );
  OAI21_X1 U303 ( .B1(n264), .B2(n269), .A(n285), .ZN(n72) );
  OAI21_X1 U304 ( .B1(n281), .B2(n291), .A(n321), .ZN(n71) );
  OR3_X1 U305 ( .A1(n268), .A2(n264), .A3(n281), .ZN(n321) );
  OAI21_X1 U306 ( .B1(n278), .B2(n301), .A(n322), .ZN(n70) );
  OR3_X1 U307 ( .A1(n299), .A2(n264), .A3(n278), .ZN(n322) );
  OAI21_X1 U308 ( .B1(n275), .B2(n312), .A(n323), .ZN(n69) );
  OR3_X1 U309 ( .A1(n310), .A2(n271), .A3(n275), .ZN(n323) );
  XNOR2_X1 U310 ( .A(n324), .B(n325), .ZN(n38) );
  OR2_X1 U311 ( .A1(n324), .A2(n325), .ZN(n37) );
  OAI22_X1 U312 ( .A1(n296), .A2(n291), .B1(n268), .B2(n326), .ZN(n325) );
  XNOR2_X1 U313 ( .A(b[5]), .B(a[3]), .ZN(n296) );
  OAI22_X1 U314 ( .A1(n313), .A2(n312), .B1(n310), .B2(n314), .ZN(n324) );
  XNOR2_X1 U315 ( .A(b[2]), .B(a[7]), .ZN(n314) );
  XNOR2_X1 U316 ( .A(b[1]), .B(a[7]), .ZN(n313) );
  OAI22_X1 U317 ( .A1(n326), .A2(n291), .B1(n268), .B2(n298), .ZN(n31) );
  XNOR2_X1 U318 ( .A(b[7]), .B(a[3]), .ZN(n298) );
  XNOR2_X1 U319 ( .A(n281), .B(a[2]), .ZN(n327) );
  XNOR2_X1 U320 ( .A(b[6]), .B(a[3]), .ZN(n326) );
  OAI22_X1 U321 ( .A1(n307), .A2(n301), .B1(n299), .B2(n309), .ZN(n21) );
  XNOR2_X1 U322 ( .A(b[7]), .B(a[5]), .ZN(n309) );
  XNOR2_X1 U323 ( .A(n278), .B(a[4]), .ZN(n328) );
  XNOR2_X1 U324 ( .A(b[6]), .B(a[5]), .ZN(n307) );
  OAI22_X1 U325 ( .A1(n318), .A2(n312), .B1(n310), .B2(n320), .ZN(n15) );
  XNOR2_X1 U326 ( .A(b[7]), .B(a[7]), .ZN(n320) );
  NAND2_X1 U327 ( .A1(n310), .A2(n329), .ZN(n312) );
  XNOR2_X1 U328 ( .A(n275), .B(a[6]), .ZN(n329) );
  XNOR2_X1 U329 ( .A(b[6]), .B(a[7]), .ZN(n318) );
  OAI22_X1 U330 ( .A1(n271), .A2(n285), .B1(n330), .B2(n283), .ZN(n104) );
  OAI22_X1 U331 ( .A1(n242), .A2(n285), .B1(n331), .B2(n283), .ZN(n103) );
  XNOR2_X1 U332 ( .A(b[1]), .B(n270), .ZN(n330) );
  OAI22_X1 U333 ( .A1(n331), .A2(n285), .B1(n332), .B2(n283), .ZN(n102) );
  XNOR2_X1 U334 ( .A(b[2]), .B(n270), .ZN(n331) );
  OAI22_X1 U335 ( .A1(n332), .A2(n285), .B1(n333), .B2(n283), .ZN(n101) );
  XNOR2_X1 U336 ( .A(b[3]), .B(n270), .ZN(n332) );
  OAI22_X1 U337 ( .A1(n333), .A2(n285), .B1(n284), .B2(n283), .ZN(n100) );
  XNOR2_X1 U338 ( .A(b[5]), .B(n270), .ZN(n284) );
  NAND2_X1 U339 ( .A1(a[1]), .A2(n283), .ZN(n285) );
  XNOR2_X1 U340 ( .A(b[4]), .B(n270), .ZN(n333) );
endmodule


module datapath_DW01_add_12 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n77;
  wire   [15:1] carry;

  FA_X1 U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n77), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[14]), .ZN(n37) );
  CLKBUF_X1 U2 ( .A(carry[3]), .Z(n1) );
  NAND3_X1 U3 ( .A1(n8), .A2(n9), .A3(n10), .ZN(n2) );
  NAND3_X1 U4 ( .A1(n8), .A2(n9), .A3(n10), .ZN(n3) );
  NAND3_X1 U5 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n4) );
  CLKBUF_X1 U6 ( .A(n29), .Z(n5) );
  NAND3_X1 U7 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n6) );
  XOR2_X1 U8 ( .A(B[3]), .B(A[3]), .Z(n7) );
  XOR2_X1 U9 ( .A(n1), .B(n7), .Z(SUM[3]) );
  NAND2_X1 U10 ( .A1(carry[3]), .A2(B[3]), .ZN(n8) );
  NAND2_X1 U11 ( .A1(carry[3]), .A2(A[3]), .ZN(n9) );
  NAND2_X1 U12 ( .A1(B[3]), .A2(A[3]), .ZN(n10) );
  NAND3_X1 U13 ( .A1(n8), .A2(n9), .A3(n10), .ZN(carry[4]) );
  CLKBUF_X1 U14 ( .A(n39), .Z(n11) );
  NAND3_X1 U15 ( .A1(n75), .A2(n74), .A3(n73), .ZN(n12) );
  CLKBUF_X1 U16 ( .A(n23), .Z(n13) );
  NAND3_X1 U17 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n14) );
  CLKBUF_X1 U18 ( .A(n4), .Z(n15) );
  XOR2_X1 U19 ( .A(B[4]), .B(A[4]), .Z(n16) );
  XOR2_X1 U20 ( .A(n3), .B(n16), .Z(SUM[4]) );
  NAND2_X1 U21 ( .A1(n2), .A2(B[4]), .ZN(n17) );
  NAND2_X1 U22 ( .A1(carry[4]), .A2(A[4]), .ZN(n18) );
  NAND2_X1 U23 ( .A1(B[4]), .A2(A[4]), .ZN(n19) );
  NAND3_X1 U24 ( .A1(n17), .A2(n18), .A3(n19), .ZN(carry[5]) );
  CLKBUF_X1 U25 ( .A(n6), .Z(n20) );
  NAND3_X1 U26 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n21) );
  NAND3_X1 U27 ( .A1(n5), .A2(n30), .A3(n31), .ZN(n22) );
  NAND3_X1 U28 ( .A1(n44), .A2(n43), .A3(n45), .ZN(n23) );
  NAND3_X1 U29 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n24) );
  NAND3_X1 U30 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n25) );
  NAND3_X1 U31 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n26) );
  NAND3_X1 U32 ( .A1(n11), .A2(n40), .A3(n41), .ZN(n27) );
  XOR2_X1 U33 ( .A(n12), .B(A[10]), .Z(n28) );
  XOR2_X1 U34 ( .A(B[10]), .B(n28), .Z(SUM[10]) );
  NAND2_X1 U35 ( .A1(n12), .A2(B[10]), .ZN(n29) );
  NAND2_X1 U36 ( .A1(B[10]), .A2(A[10]), .ZN(n30) );
  NAND2_X1 U37 ( .A1(carry[10]), .A2(A[10]), .ZN(n31) );
  NAND3_X1 U38 ( .A1(n29), .A2(n30), .A3(n31), .ZN(carry[11]) );
  CLKBUF_X1 U39 ( .A(n71), .Z(n32) );
  XOR2_X1 U40 ( .A(B[5]), .B(A[5]), .Z(n33) );
  XOR2_X1 U41 ( .A(n15), .B(n33), .Z(SUM[5]) );
  NAND2_X1 U42 ( .A1(n4), .A2(B[5]), .ZN(n34) );
  NAND2_X1 U43 ( .A1(carry[5]), .A2(A[5]), .ZN(n35) );
  NAND2_X1 U44 ( .A1(B[5]), .A2(A[5]), .ZN(n36) );
  NAND3_X1 U45 ( .A1(n34), .A2(n35), .A3(n36), .ZN(carry[6]) );
  XNOR2_X1 U46 ( .A(B[14]), .B(n37), .ZN(n57) );
  XOR2_X1 U47 ( .A(n13), .B(A[12]), .Z(n38) );
  XOR2_X1 U48 ( .A(B[12]), .B(n38), .Z(SUM[12]) );
  NAND2_X1 U49 ( .A1(n23), .A2(B[12]), .ZN(n39) );
  NAND2_X1 U50 ( .A1(B[12]), .A2(A[12]), .ZN(n40) );
  NAND2_X1 U51 ( .A1(carry[12]), .A2(A[12]), .ZN(n41) );
  NAND3_X1 U52 ( .A1(n39), .A2(n40), .A3(n41), .ZN(carry[13]) );
  XOR2_X1 U53 ( .A(B[11]), .B(A[11]), .Z(n42) );
  XOR2_X1 U54 ( .A(n22), .B(n42), .Z(SUM[11]) );
  NAND2_X1 U55 ( .A1(n21), .A2(B[11]), .ZN(n43) );
  NAND2_X1 U56 ( .A1(carry[11]), .A2(A[11]), .ZN(n44) );
  NAND2_X1 U57 ( .A1(B[11]), .A2(A[11]), .ZN(n45) );
  NAND3_X1 U58 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[12]) );
  CLKBUF_X1 U59 ( .A(n14), .Z(n46) );
  XOR2_X1 U60 ( .A(B[6]), .B(A[6]), .Z(n47) );
  XOR2_X1 U61 ( .A(n20), .B(n47), .Z(SUM[6]) );
  NAND2_X1 U62 ( .A1(n6), .A2(B[6]), .ZN(n48) );
  NAND2_X1 U63 ( .A1(carry[6]), .A2(A[6]), .ZN(n49) );
  NAND2_X1 U64 ( .A1(B[6]), .A2(A[6]), .ZN(n50) );
  NAND3_X1 U65 ( .A1(n48), .A2(n49), .A3(n50), .ZN(carry[7]) );
  NAND3_X1 U66 ( .A1(n56), .A2(n55), .A3(n54), .ZN(n51) );
  NAND3_X1 U67 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n52) );
  XOR2_X1 U68 ( .A(A[13]), .B(B[13]), .Z(n53) );
  XOR2_X1 U69 ( .A(n53), .B(n27), .Z(SUM[13]) );
  NAND2_X1 U70 ( .A1(A[13]), .A2(B[13]), .ZN(n54) );
  NAND2_X1 U71 ( .A1(carry[13]), .A2(A[13]), .ZN(n55) );
  NAND2_X1 U72 ( .A1(n26), .A2(B[13]), .ZN(n56) );
  NAND3_X1 U73 ( .A1(n56), .A2(n55), .A3(n54), .ZN(carry[14]) );
  XOR2_X1 U74 ( .A(n57), .B(n52), .Z(SUM[14]) );
  NAND2_X1 U75 ( .A1(A[14]), .A2(B[14]), .ZN(n58) );
  NAND2_X1 U76 ( .A1(A[14]), .A2(n51), .ZN(n59) );
  NAND2_X1 U77 ( .A1(B[14]), .A2(carry[14]), .ZN(n60) );
  NAND3_X1 U78 ( .A1(n59), .A2(n60), .A3(n58), .ZN(carry[15]) );
  XOR2_X1 U79 ( .A(B[7]), .B(A[7]), .Z(n61) );
  XOR2_X1 U80 ( .A(n46), .B(n61), .Z(SUM[7]) );
  NAND2_X1 U81 ( .A1(n14), .A2(B[7]), .ZN(n62) );
  NAND2_X1 U82 ( .A1(carry[7]), .A2(A[7]), .ZN(n63) );
  NAND2_X1 U83 ( .A1(B[7]), .A2(A[7]), .ZN(n64) );
  NAND3_X1 U84 ( .A1(n62), .A2(n63), .A3(n64), .ZN(carry[8]) );
  NAND3_X1 U85 ( .A1(n71), .A2(n70), .A3(n69), .ZN(n65) );
  NAND3_X1 U86 ( .A1(n69), .A2(n70), .A3(n32), .ZN(n66) );
  XNOR2_X1 U87 ( .A(carry[15]), .B(n67), .ZN(SUM[15]) );
  XNOR2_X1 U88 ( .A(B[15]), .B(A[15]), .ZN(n67) );
  XOR2_X1 U89 ( .A(A[8]), .B(B[8]), .Z(n68) );
  XOR2_X1 U90 ( .A(n68), .B(n25), .Z(SUM[8]) );
  NAND2_X1 U91 ( .A1(A[8]), .A2(B[8]), .ZN(n69) );
  NAND2_X1 U92 ( .A1(carry[8]), .A2(A[8]), .ZN(n70) );
  NAND2_X1 U93 ( .A1(B[8]), .A2(n24), .ZN(n71) );
  NAND3_X1 U94 ( .A1(n69), .A2(n70), .A3(n71), .ZN(carry[9]) );
  XOR2_X1 U95 ( .A(A[9]), .B(B[9]), .Z(n72) );
  XOR2_X1 U96 ( .A(n72), .B(n66), .Z(SUM[9]) );
  NAND2_X1 U97 ( .A1(A[9]), .A2(B[9]), .ZN(n73) );
  NAND2_X1 U98 ( .A1(n65), .A2(A[9]), .ZN(n74) );
  NAND2_X1 U99 ( .A1(B[9]), .A2(carry[9]), .ZN(n75) );
  NAND3_X1 U100 ( .A1(n75), .A2(n74), .A3(n73), .ZN(carry[10]) );
  XOR2_X1 U101 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U102 ( .A1(B[0]), .A2(A[0]), .ZN(n77) );
endmodule


module datapath_DW_mult_tc_11 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74,
         n75, n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92,
         n93, n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206,
         n207, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337;

  FA_X1 U12 ( .A(n54), .B(n55), .CI(n12), .CO(n11), .S(product[4]) );
  FA_X1 U13 ( .A(n71), .B(n13), .CI(n56), .CO(n12), .S(product[3]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n280), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n279), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n283), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n282), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n285), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  BUF_X2 U157 ( .A(a[1]), .Z(n206) );
  NAND2_X1 U158 ( .A1(n303), .A2(n332), .ZN(n305) );
  CLKBUF_X1 U159 ( .A(n275), .Z(n223) );
  NOR2_X1 U160 ( .A1(n270), .A2(n223), .ZN(n96) );
  INV_X1 U161 ( .A(n15), .ZN(n276) );
  CLKBUF_X1 U162 ( .A(n334), .Z(n207) );
  AND3_X1 U163 ( .A1(n224), .A2(n225), .A3(n226), .ZN(product[15]) );
  XNOR2_X1 U164 ( .A(n277), .B(n15), .ZN(n209) );
  XOR2_X1 U165 ( .A(n50), .B(n53), .Z(n210) );
  XOR2_X1 U166 ( .A(n11), .B(n210), .Z(product[5]) );
  NAND2_X1 U167 ( .A1(n11), .A2(n50), .ZN(n211) );
  NAND2_X1 U168 ( .A1(n11), .A2(n53), .ZN(n212) );
  NAND2_X1 U169 ( .A1(n50), .A2(n53), .ZN(n213) );
  NAND3_X1 U170 ( .A1(n211), .A2(n212), .A3(n213), .ZN(n10) );
  XOR2_X2 U171 ( .A(a[6]), .B(n281), .Z(n314) );
  XOR2_X1 U172 ( .A(n103), .B(n96), .Z(n214) );
  XOR2_X1 U173 ( .A(n14), .B(n214), .Z(product[2]) );
  NAND2_X1 U174 ( .A1(n14), .A2(n103), .ZN(n215) );
  NAND2_X1 U175 ( .A1(n14), .A2(n96), .ZN(n216) );
  NAND2_X1 U176 ( .A1(n103), .A2(n96), .ZN(n217) );
  NAND3_X1 U177 ( .A1(n215), .A2(n216), .A3(n217), .ZN(n13) );
  XOR2_X1 U178 ( .A(n46), .B(n49), .Z(n218) );
  XOR2_X1 U179 ( .A(n10), .B(n218), .Z(product[6]) );
  NAND2_X1 U180 ( .A1(n10), .A2(n46), .ZN(n219) );
  NAND2_X1 U181 ( .A1(n10), .A2(n49), .ZN(n220) );
  NAND2_X1 U182 ( .A1(n46), .A2(n49), .ZN(n221) );
  NAND3_X1 U183 ( .A1(n219), .A2(n220), .A3(n221), .ZN(n9) );
  NAND3_X1 U184 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n222) );
  XNOR2_X1 U185 ( .A(n2), .B(n209), .ZN(product[14]) );
  NAND2_X1 U186 ( .A1(n2), .A2(n277), .ZN(n224) );
  NAND2_X1 U187 ( .A1(n2), .A2(n15), .ZN(n225) );
  NAND2_X1 U188 ( .A1(n277), .A2(n15), .ZN(n226) );
  NAND3_X1 U189 ( .A1(n252), .A2(n251), .A3(n253), .ZN(n227) );
  NAND3_X1 U190 ( .A1(n252), .A2(n251), .A3(n253), .ZN(n228) );
  NAND3_X1 U191 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n229) );
  NAND3_X1 U192 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n230) );
  INV_X2 U193 ( .A(a[0]), .ZN(n287) );
  XOR2_X1 U194 ( .A(n40), .B(n45), .Z(n231) );
  XOR2_X1 U195 ( .A(n9), .B(n231), .Z(product[7]) );
  NAND2_X1 U196 ( .A1(n9), .A2(n40), .ZN(n232) );
  NAND2_X1 U197 ( .A1(n9), .A2(n45), .ZN(n233) );
  NAND2_X1 U198 ( .A1(n40), .A2(n45), .ZN(n234) );
  NAND3_X1 U199 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n8) );
  NAND3_X1 U200 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n235) );
  NAND3_X1 U201 ( .A1(n258), .A2(n257), .A3(n259), .ZN(n236) );
  XOR2_X1 U202 ( .A(n34), .B(n39), .Z(n237) );
  XOR2_X1 U203 ( .A(n222), .B(n237), .Z(product[8]) );
  NAND2_X1 U204 ( .A1(n222), .A2(n34), .ZN(n238) );
  NAND2_X1 U205 ( .A1(n8), .A2(n39), .ZN(n239) );
  NAND2_X1 U206 ( .A1(n34), .A2(n39), .ZN(n240) );
  NAND3_X1 U207 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n7) );
  XOR2_X1 U208 ( .A(n18), .B(n19), .Z(n241) );
  XOR2_X1 U209 ( .A(n228), .B(n241), .Z(product[12]) );
  NAND2_X1 U210 ( .A1(n227), .A2(n18), .ZN(n242) );
  NAND2_X1 U211 ( .A1(n4), .A2(n19), .ZN(n243) );
  NAND2_X1 U212 ( .A1(n18), .A2(n19), .ZN(n244) );
  NAND3_X1 U213 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n3) );
  NAND3_X1 U214 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n245) );
  XOR2_X1 U215 ( .A(n17), .B(n276), .Z(n246) );
  XOR2_X1 U216 ( .A(n230), .B(n246), .Z(product[13]) );
  NAND2_X1 U217 ( .A1(n229), .A2(n17), .ZN(n247) );
  NAND2_X1 U218 ( .A1(n3), .A2(n276), .ZN(n248) );
  NAND2_X1 U219 ( .A1(n17), .A2(n276), .ZN(n249) );
  NAND3_X1 U220 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n2) );
  NAND2_X2 U221 ( .A1(n293), .A2(n331), .ZN(n295) );
  XOR2_X1 U222 ( .A(n23), .B(n20), .Z(n250) );
  XOR2_X1 U223 ( .A(n245), .B(n250), .Z(product[11]) );
  NAND2_X1 U224 ( .A1(n5), .A2(n23), .ZN(n251) );
  NAND2_X1 U225 ( .A1(n245), .A2(n20), .ZN(n252) );
  NAND2_X1 U226 ( .A1(n23), .A2(n20), .ZN(n253) );
  NAND3_X1 U227 ( .A1(n252), .A2(n251), .A3(n253), .ZN(n4) );
  NAND3_X1 U228 ( .A1(n259), .A2(n258), .A3(n257), .ZN(n254) );
  CLKBUF_X1 U229 ( .A(b[1]), .Z(n255) );
  XOR2_X1 U230 ( .A(n28), .B(n33), .Z(n256) );
  XOR2_X1 U231 ( .A(n256), .B(n235), .Z(product[9]) );
  NAND2_X1 U232 ( .A1(n28), .A2(n33), .ZN(n257) );
  NAND2_X1 U233 ( .A1(n28), .A2(n7), .ZN(n258) );
  NAND2_X1 U234 ( .A1(n33), .A2(n7), .ZN(n259) );
  NAND3_X1 U235 ( .A1(n259), .A2(n258), .A3(n257), .ZN(n6) );
  XOR2_X1 U236 ( .A(n24), .B(n27), .Z(n260) );
  XOR2_X1 U237 ( .A(n260), .B(n236), .Z(product[10]) );
  NAND2_X1 U238 ( .A1(n24), .A2(n27), .ZN(n261) );
  NAND2_X1 U239 ( .A1(n24), .A2(n254), .ZN(n262) );
  NAND2_X1 U240 ( .A1(n27), .A2(n6), .ZN(n263) );
  NAND3_X1 U241 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n5) );
  INV_X1 U242 ( .A(n275), .ZN(n264) );
  NAND2_X1 U243 ( .A1(a[4]), .A2(a[3]), .ZN(n267) );
  NAND2_X1 U244 ( .A1(n265), .A2(n266), .ZN(n268) );
  NAND2_X2 U245 ( .A1(n267), .A2(n268), .ZN(n303) );
  INV_X1 U246 ( .A(a[4]), .ZN(n265) );
  INV_X1 U247 ( .A(a[3]), .ZN(n266) );
  NAND2_X1 U248 ( .A1(n272), .A2(n273), .ZN(n269) );
  NAND2_X1 U249 ( .A1(n272), .A2(n273), .ZN(n270) );
  NAND2_X1 U250 ( .A1(n272), .A2(n273), .ZN(n293) );
  NAND2_X1 U251 ( .A1(a[2]), .A2(n206), .ZN(n272) );
  NAND2_X1 U252 ( .A1(n271), .A2(n286), .ZN(n273) );
  INV_X1 U253 ( .A(a[2]), .ZN(n271) );
  INV_X1 U254 ( .A(n21), .ZN(n279) );
  INV_X1 U255 ( .A(n312), .ZN(n280) );
  INV_X1 U256 ( .A(n323), .ZN(n277) );
  INV_X1 U257 ( .A(n292), .ZN(n285) );
  INV_X1 U258 ( .A(n301), .ZN(n283) );
  INV_X1 U259 ( .A(n31), .ZN(n282) );
  INV_X1 U260 ( .A(b[0]), .ZN(n275) );
  INV_X1 U261 ( .A(a[5]), .ZN(n281) );
  INV_X1 U262 ( .A(a[7]), .ZN(n278) );
  INV_X1 U263 ( .A(a[3]), .ZN(n284) );
  INV_X1 U264 ( .A(a[1]), .ZN(n286) );
  INV_X1 U265 ( .A(n275), .ZN(n274) );
  NOR2_X1 U266 ( .A1(n287), .A2(n223), .ZN(product[0]) );
  OAI22_X1 U267 ( .A1(n288), .A2(n289), .B1(n290), .B2(n287), .ZN(n99) );
  OAI22_X1 U268 ( .A1(n290), .A2(n289), .B1(n291), .B2(n287), .ZN(n98) );
  XNOR2_X1 U269 ( .A(b[6]), .B(n206), .ZN(n290) );
  OAI22_X1 U270 ( .A1(n287), .A2(n291), .B1(n289), .B2(n291), .ZN(n292) );
  XNOR2_X1 U271 ( .A(b[7]), .B(n206), .ZN(n291) );
  OAI22_X1 U272 ( .A1(n294), .A2(n295), .B1(n269), .B2(n296), .ZN(n95) );
  XNOR2_X1 U273 ( .A(a[3]), .B(n274), .ZN(n294) );
  OAI22_X1 U274 ( .A1(n296), .A2(n295), .B1(n269), .B2(n297), .ZN(n94) );
  XNOR2_X1 U275 ( .A(n255), .B(a[3]), .ZN(n296) );
  OAI22_X1 U276 ( .A1(n297), .A2(n295), .B1(n269), .B2(n298), .ZN(n93) );
  XNOR2_X1 U277 ( .A(b[2]), .B(a[3]), .ZN(n297) );
  OAI22_X1 U278 ( .A1(n298), .A2(n295), .B1(n270), .B2(n299), .ZN(n92) );
  XNOR2_X1 U279 ( .A(b[3]), .B(a[3]), .ZN(n298) );
  OAI22_X1 U280 ( .A1(n299), .A2(n295), .B1(n270), .B2(n300), .ZN(n91) );
  XNOR2_X1 U281 ( .A(b[4]), .B(a[3]), .ZN(n299) );
  OAI22_X1 U282 ( .A1(n302), .A2(n269), .B1(n295), .B2(n302), .ZN(n301) );
  NOR2_X1 U283 ( .A1(n303), .A2(n223), .ZN(n88) );
  OAI22_X1 U284 ( .A1(n304), .A2(n305), .B1(n303), .B2(n306), .ZN(n87) );
  XNOR2_X1 U285 ( .A(a[5]), .B(n274), .ZN(n304) );
  OAI22_X1 U286 ( .A1(n306), .A2(n305), .B1(n303), .B2(n307), .ZN(n86) );
  XNOR2_X1 U287 ( .A(n255), .B(a[5]), .ZN(n306) );
  OAI22_X1 U288 ( .A1(n307), .A2(n305), .B1(n303), .B2(n308), .ZN(n85) );
  XNOR2_X1 U289 ( .A(b[2]), .B(a[5]), .ZN(n307) );
  OAI22_X1 U290 ( .A1(n308), .A2(n305), .B1(n303), .B2(n309), .ZN(n84) );
  XNOR2_X1 U291 ( .A(b[3]), .B(a[5]), .ZN(n308) );
  OAI22_X1 U292 ( .A1(n309), .A2(n305), .B1(n303), .B2(n310), .ZN(n83) );
  XNOR2_X1 U293 ( .A(b[4]), .B(a[5]), .ZN(n309) );
  OAI22_X1 U294 ( .A1(n310), .A2(n305), .B1(n303), .B2(n311), .ZN(n82) );
  XNOR2_X1 U295 ( .A(b[5]), .B(a[5]), .ZN(n310) );
  OAI22_X1 U296 ( .A1(n313), .A2(n303), .B1(n305), .B2(n313), .ZN(n312) );
  NOR2_X1 U297 ( .A1(n314), .A2(n223), .ZN(n80) );
  OAI22_X1 U298 ( .A1(n315), .A2(n316), .B1(n314), .B2(n317), .ZN(n79) );
  XNOR2_X1 U299 ( .A(a[7]), .B(n264), .ZN(n315) );
  OAI22_X1 U300 ( .A1(n318), .A2(n316), .B1(n314), .B2(n319), .ZN(n77) );
  OAI22_X1 U301 ( .A1(n319), .A2(n316), .B1(n314), .B2(n320), .ZN(n76) );
  XNOR2_X1 U302 ( .A(b[3]), .B(a[7]), .ZN(n319) );
  OAI22_X1 U303 ( .A1(n320), .A2(n316), .B1(n314), .B2(n321), .ZN(n75) );
  XNOR2_X1 U304 ( .A(b[4]), .B(a[7]), .ZN(n320) );
  OAI22_X1 U305 ( .A1(n321), .A2(n316), .B1(n314), .B2(n322), .ZN(n74) );
  XNOR2_X1 U306 ( .A(b[5]), .B(a[7]), .ZN(n321) );
  OAI22_X1 U307 ( .A1(n324), .A2(n314), .B1(n316), .B2(n324), .ZN(n323) );
  OAI21_X1 U308 ( .B1(n264), .B2(n286), .A(n289), .ZN(n72) );
  OAI21_X1 U309 ( .B1(n284), .B2(n295), .A(n325), .ZN(n71) );
  OR3_X1 U310 ( .A1(n270), .A2(n264), .A3(n284), .ZN(n325) );
  OAI21_X1 U311 ( .B1(n281), .B2(n305), .A(n326), .ZN(n70) );
  OR3_X1 U312 ( .A1(n303), .A2(n264), .A3(n281), .ZN(n326) );
  OAI21_X1 U313 ( .B1(n278), .B2(n316), .A(n327), .ZN(n69) );
  OR3_X1 U314 ( .A1(n314), .A2(n274), .A3(n278), .ZN(n327) );
  XNOR2_X1 U315 ( .A(n328), .B(n329), .ZN(n38) );
  OR2_X1 U316 ( .A1(n328), .A2(n329), .ZN(n37) );
  OAI22_X1 U317 ( .A1(n300), .A2(n295), .B1(n269), .B2(n330), .ZN(n329) );
  XNOR2_X1 U318 ( .A(b[5]), .B(a[3]), .ZN(n300) );
  OAI22_X1 U319 ( .A1(n317), .A2(n316), .B1(n314), .B2(n318), .ZN(n328) );
  XNOR2_X1 U320 ( .A(b[2]), .B(a[7]), .ZN(n318) );
  XNOR2_X1 U321 ( .A(n255), .B(a[7]), .ZN(n317) );
  OAI22_X1 U322 ( .A1(n330), .A2(n295), .B1(n270), .B2(n302), .ZN(n31) );
  XNOR2_X1 U323 ( .A(b[7]), .B(a[3]), .ZN(n302) );
  XNOR2_X1 U324 ( .A(n284), .B(a[2]), .ZN(n331) );
  XNOR2_X1 U325 ( .A(b[6]), .B(a[3]), .ZN(n330) );
  OAI22_X1 U326 ( .A1(n311), .A2(n305), .B1(n303), .B2(n313), .ZN(n21) );
  XNOR2_X1 U327 ( .A(b[7]), .B(a[5]), .ZN(n313) );
  XNOR2_X1 U328 ( .A(n281), .B(a[4]), .ZN(n332) );
  XNOR2_X1 U329 ( .A(b[6]), .B(a[5]), .ZN(n311) );
  OAI22_X1 U330 ( .A1(n322), .A2(n316), .B1(n314), .B2(n324), .ZN(n15) );
  XNOR2_X1 U331 ( .A(b[7]), .B(a[7]), .ZN(n324) );
  NAND2_X1 U332 ( .A1(n314), .A2(n333), .ZN(n316) );
  XNOR2_X1 U333 ( .A(n278), .B(a[6]), .ZN(n333) );
  XNOR2_X1 U334 ( .A(b[6]), .B(a[7]), .ZN(n322) );
  OAI22_X1 U335 ( .A1(n274), .A2(n289), .B1(n334), .B2(n287), .ZN(n104) );
  OAI22_X1 U336 ( .A1(n207), .A2(n289), .B1(n335), .B2(n287), .ZN(n103) );
  XNOR2_X1 U337 ( .A(b[1]), .B(n206), .ZN(n334) );
  OAI22_X1 U338 ( .A1(n335), .A2(n289), .B1(n336), .B2(n287), .ZN(n102) );
  XNOR2_X1 U339 ( .A(b[2]), .B(n206), .ZN(n335) );
  OAI22_X1 U340 ( .A1(n336), .A2(n289), .B1(n337), .B2(n287), .ZN(n101) );
  XNOR2_X1 U341 ( .A(b[3]), .B(n206), .ZN(n336) );
  OAI22_X1 U342 ( .A1(n337), .A2(n289), .B1(n288), .B2(n287), .ZN(n100) );
  XNOR2_X1 U343 ( .A(b[5]), .B(n206), .ZN(n288) );
  NAND2_X1 U344 ( .A1(n206), .A2(n287), .ZN(n289) );
  XNOR2_X1 U345 ( .A(b[4]), .B(n206), .ZN(n337) );
endmodule


module datapath_DW01_add_11 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n67;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n67), .CO(carry[2]), .S(SUM[1]) );
  XNOR2_X1 U1 ( .A(B[15]), .B(A[15]), .ZN(n52) );
  NAND3_X1 U2 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n1) );
  NAND3_X1 U3 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n2) );
  NAND3_X1 U4 ( .A1(n6), .A2(n7), .A3(n8), .ZN(n3) );
  CLKBUF_X1 U5 ( .A(B[2]), .Z(n4) );
  XOR2_X1 U6 ( .A(n4), .B(A[2]), .Z(n5) );
  XOR2_X1 U7 ( .A(n5), .B(carry[2]), .Z(SUM[2]) );
  NAND2_X1 U8 ( .A1(B[2]), .A2(A[2]), .ZN(n6) );
  NAND2_X1 U9 ( .A1(B[2]), .A2(carry[2]), .ZN(n7) );
  NAND2_X1 U10 ( .A1(A[2]), .A2(carry[2]), .ZN(n8) );
  NAND3_X1 U11 ( .A1(n6), .A2(n7), .A3(n8), .ZN(carry[3]) );
  XOR2_X1 U12 ( .A(A[3]), .B(B[3]), .Z(n9) );
  XOR2_X1 U13 ( .A(n9), .B(carry[3]), .Z(SUM[3]) );
  NAND2_X1 U14 ( .A1(A[3]), .A2(B[3]), .ZN(n10) );
  NAND2_X1 U15 ( .A1(A[3]), .A2(n3), .ZN(n11) );
  NAND2_X1 U16 ( .A1(B[3]), .A2(carry[3]), .ZN(n12) );
  NAND3_X1 U17 ( .A1(n10), .A2(n11), .A3(n12), .ZN(carry[4]) );
  CLKBUF_X1 U18 ( .A(n64), .Z(n13) );
  CLKBUF_X1 U19 ( .A(n47), .Z(n14) );
  CLKBUF_X1 U20 ( .A(carry[12]), .Z(n15) );
  NAND3_X1 U21 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n16) );
  XOR2_X1 U22 ( .A(B[5]), .B(A[5]), .Z(n17) );
  XOR2_X1 U23 ( .A(carry[5]), .B(n17), .Z(SUM[5]) );
  NAND2_X1 U24 ( .A1(carry[5]), .A2(B[5]), .ZN(n18) );
  NAND2_X1 U25 ( .A1(carry[5]), .A2(A[5]), .ZN(n19) );
  NAND2_X1 U26 ( .A1(B[5]), .A2(A[5]), .ZN(n20) );
  NAND3_X1 U27 ( .A1(n18), .A2(n19), .A3(n20), .ZN(carry[6]) );
  NAND3_X1 U28 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n21) );
  NAND3_X1 U29 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n22) );
  NAND3_X1 U30 ( .A1(n45), .A2(n46), .A3(n14), .ZN(n23) );
  NAND3_X1 U31 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n24) );
  XOR2_X1 U32 ( .A(B[13]), .B(A[13]), .Z(n25) );
  XOR2_X1 U33 ( .A(n23), .B(n25), .Z(SUM[13]) );
  NAND2_X1 U34 ( .A1(n22), .A2(B[13]), .ZN(n26) );
  NAND2_X1 U35 ( .A1(carry[13]), .A2(A[13]), .ZN(n27) );
  NAND2_X1 U36 ( .A1(B[13]), .A2(A[13]), .ZN(n28) );
  NAND3_X1 U37 ( .A1(n26), .A2(n27), .A3(n28), .ZN(carry[14]) );
  CLKBUF_X1 U38 ( .A(carry[8]), .Z(n29) );
  CLKBUF_X1 U39 ( .A(n21), .Z(n30) );
  CLKBUF_X1 U40 ( .A(carry[10]), .Z(n31) );
  CLKBUF_X1 U41 ( .A(n65), .Z(n32) );
  XOR2_X1 U42 ( .A(B[6]), .B(A[6]), .Z(n33) );
  XOR2_X1 U43 ( .A(n2), .B(n33), .Z(SUM[6]) );
  NAND2_X1 U44 ( .A1(n1), .A2(B[6]), .ZN(n34) );
  NAND2_X1 U45 ( .A1(carry[6]), .A2(A[6]), .ZN(n35) );
  NAND2_X1 U46 ( .A1(B[6]), .A2(A[6]), .ZN(n36) );
  NAND3_X1 U47 ( .A1(n35), .A2(n34), .A3(n36), .ZN(carry[7]) );
  NAND3_X1 U48 ( .A1(n65), .A2(n64), .A3(n63), .ZN(n37) );
  NAND3_X1 U49 ( .A1(n63), .A2(n13), .A3(n32), .ZN(n38) );
  NAND3_X1 U50 ( .A1(n42), .A2(n41), .A3(n43), .ZN(n39) );
  XOR2_X1 U51 ( .A(A[11]), .B(B[11]), .Z(n40) );
  XOR2_X1 U52 ( .A(n40), .B(n38), .Z(SUM[11]) );
  NAND2_X1 U53 ( .A1(A[11]), .A2(B[11]), .ZN(n41) );
  NAND2_X1 U54 ( .A1(A[11]), .A2(n37), .ZN(n42) );
  NAND2_X1 U55 ( .A1(B[11]), .A2(carry[11]), .ZN(n43) );
  NAND3_X1 U56 ( .A1(n43), .A2(n42), .A3(n41), .ZN(carry[12]) );
  XOR2_X1 U57 ( .A(A[12]), .B(B[12]), .Z(n44) );
  XOR2_X1 U58 ( .A(n44), .B(n15), .Z(SUM[12]) );
  NAND2_X1 U59 ( .A1(A[12]), .A2(B[12]), .ZN(n45) );
  NAND2_X1 U60 ( .A1(A[12]), .A2(n39), .ZN(n46) );
  NAND2_X1 U61 ( .A1(B[12]), .A2(carry[12]), .ZN(n47) );
  NAND3_X1 U62 ( .A1(n45), .A2(n46), .A3(n47), .ZN(carry[13]) );
  XOR2_X1 U63 ( .A(B[7]), .B(A[7]), .Z(n48) );
  XOR2_X1 U64 ( .A(n30), .B(n48), .Z(SUM[7]) );
  NAND2_X1 U65 ( .A1(n21), .A2(B[7]), .ZN(n49) );
  NAND2_X1 U66 ( .A1(carry[7]), .A2(A[7]), .ZN(n50) );
  NAND2_X1 U67 ( .A1(B[7]), .A2(A[7]), .ZN(n51) );
  NAND3_X1 U68 ( .A1(n49), .A2(n50), .A3(n51), .ZN(carry[8]) );
  XNOR2_X1 U69 ( .A(carry[15]), .B(n52), .ZN(SUM[15]) );
  XOR2_X1 U70 ( .A(B[8]), .B(A[8]), .Z(n53) );
  XOR2_X1 U71 ( .A(n29), .B(n53), .Z(SUM[8]) );
  NAND2_X1 U72 ( .A1(carry[8]), .A2(B[8]), .ZN(n54) );
  NAND2_X1 U73 ( .A1(n16), .A2(A[8]), .ZN(n55) );
  NAND2_X1 U74 ( .A1(B[8]), .A2(A[8]), .ZN(n56) );
  NAND3_X1 U75 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[9]) );
  NAND3_X1 U76 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n57) );
  XOR2_X1 U77 ( .A(A[9]), .B(B[9]), .Z(n58) );
  XOR2_X1 U78 ( .A(n58), .B(carry[9]), .Z(SUM[9]) );
  NAND2_X1 U79 ( .A1(A[9]), .A2(B[9]), .ZN(n59) );
  NAND2_X1 U80 ( .A1(n24), .A2(A[9]), .ZN(n60) );
  NAND2_X1 U81 ( .A1(B[9]), .A2(n24), .ZN(n61) );
  NAND3_X1 U82 ( .A1(n61), .A2(n60), .A3(n59), .ZN(carry[10]) );
  XOR2_X1 U83 ( .A(A[10]), .B(B[10]), .Z(n62) );
  XOR2_X1 U84 ( .A(n62), .B(n31), .Z(SUM[10]) );
  NAND2_X1 U85 ( .A1(B[10]), .A2(A[10]), .ZN(n63) );
  NAND2_X1 U86 ( .A1(A[10]), .A2(n57), .ZN(n64) );
  NAND2_X1 U87 ( .A1(carry[10]), .A2(B[10]), .ZN(n65) );
  NAND3_X1 U88 ( .A1(n65), .A2(n64), .A3(n63), .ZN(carry[11]) );
  XOR2_X1 U89 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U90 ( .A1(B[0]), .A2(A[0]), .ZN(n67) );
endmodule


module datapath_DW_mult_tc_10 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334;

  FA_X1 U5 ( .A(n20), .B(n23), .CI(n5), .CO(n4), .S(product[11]) );
  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n277), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n276), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n280), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n279), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n282), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n206), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  OR3_X1 U157 ( .A1(n300), .A2(n265), .A3(n278), .ZN(n323) );
  INV_X1 U158 ( .A(n15), .ZN(n273) );
  AND2_X1 U159 ( .A1(n223), .A2(n87), .ZN(n206) );
  XNOR2_X1 U160 ( .A(n274), .B(n15), .ZN(n207) );
  AND3_X1 U161 ( .A1(n236), .A2(n237), .A3(n238), .ZN(product[15]) );
  XNOR2_X1 U162 ( .A(n2), .B(n207), .ZN(product[14]) );
  XOR2_X1 U163 ( .A(n95), .B(n102), .Z(n209) );
  NAND3_X1 U164 ( .A1(n218), .A2(n219), .A3(n220), .ZN(n210) );
  NAND3_X1 U165 ( .A1(n218), .A2(n219), .A3(n220), .ZN(n211) );
  NAND3_X1 U166 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n212) );
  NAND3_X1 U167 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n213) );
  NAND3_X1 U168 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n214) );
  XOR2_X1 U169 ( .A(a[4]), .B(a[3]), .Z(n215) );
  INV_X2 U170 ( .A(n215), .ZN(n300) );
  XNOR2_X1 U171 ( .A(n216), .B(n12), .ZN(product[4]) );
  XNOR2_X1 U172 ( .A(n54), .B(n55), .ZN(n216) );
  XOR2_X1 U173 ( .A(n19), .B(n18), .Z(n217) );
  XOR2_X1 U174 ( .A(n4), .B(n217), .Z(product[12]) );
  NAND2_X1 U175 ( .A1(n4), .A2(n19), .ZN(n218) );
  NAND2_X1 U176 ( .A1(n4), .A2(n18), .ZN(n219) );
  NAND2_X1 U177 ( .A1(n19), .A2(n18), .ZN(n220) );
  NAND3_X1 U178 ( .A1(n218), .A2(n219), .A3(n220), .ZN(n3) );
  NAND3_X1 U179 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n221) );
  NAND3_X1 U180 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n222) );
  OAI21_X1 U181 ( .B1(n278), .B2(n302), .A(n323), .ZN(n223) );
  XOR2_X2 U182 ( .A(a[6]), .B(n278), .Z(n311) );
  XOR2_X1 U183 ( .A(n34), .B(n39), .Z(n224) );
  XOR2_X1 U184 ( .A(n8), .B(n224), .Z(product[8]) );
  NAND2_X1 U185 ( .A1(n8), .A2(n34), .ZN(n225) );
  NAND2_X1 U186 ( .A1(n8), .A2(n39), .ZN(n226) );
  NAND2_X1 U187 ( .A1(n34), .A2(n39), .ZN(n227) );
  NAND3_X1 U188 ( .A1(n225), .A2(n226), .A3(n227), .ZN(n7) );
  NAND3_X1 U189 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n228) );
  NAND3_X1 U190 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n229) );
  XOR2_X1 U191 ( .A(n40), .B(n45), .Z(n230) );
  XOR2_X1 U192 ( .A(n229), .B(n230), .Z(product[7]) );
  NAND2_X1 U193 ( .A1(n228), .A2(n40), .ZN(n231) );
  NAND2_X1 U194 ( .A1(n9), .A2(n45), .ZN(n232) );
  NAND2_X1 U195 ( .A1(n40), .A2(n45), .ZN(n233) );
  NAND3_X1 U196 ( .A1(n231), .A2(n232), .A3(n233), .ZN(n8) );
  NAND3_X1 U197 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n234) );
  XNOR2_X1 U198 ( .A(n13), .B(n235), .ZN(product[3]) );
  XNOR2_X1 U199 ( .A(n56), .B(n71), .ZN(n235) );
  NAND2_X2 U200 ( .A1(n300), .A2(n329), .ZN(n302) );
  NAND2_X1 U201 ( .A1(n2), .A2(n274), .ZN(n236) );
  NAND2_X1 U202 ( .A1(n2), .A2(n15), .ZN(n237) );
  NAND2_X1 U203 ( .A1(n274), .A2(n15), .ZN(n238) );
  XOR2_X1 U204 ( .A(n70), .B(n87), .Z(n52) );
  XNOR2_X1 U205 ( .A(n239), .B(n214), .ZN(product[5]) );
  XNOR2_X1 U206 ( .A(n50), .B(n53), .ZN(n239) );
  XOR2_X1 U207 ( .A(n28), .B(n33), .Z(n240) );
  XOR2_X1 U208 ( .A(n240), .B(n7), .Z(product[9]) );
  NAND2_X1 U209 ( .A1(n28), .A2(n33), .ZN(n241) );
  NAND2_X1 U210 ( .A1(n28), .A2(n212), .ZN(n242) );
  NAND2_X1 U211 ( .A1(n33), .A2(n7), .ZN(n243) );
  NAND3_X1 U212 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n6) );
  XOR2_X1 U213 ( .A(n24), .B(n27), .Z(n244) );
  XOR2_X1 U214 ( .A(n244), .B(n222), .Z(product[10]) );
  NAND2_X1 U215 ( .A1(n24), .A2(n27), .ZN(n245) );
  NAND2_X1 U216 ( .A1(n24), .A2(n221), .ZN(n246) );
  NAND2_X1 U217 ( .A1(n27), .A2(n6), .ZN(n247) );
  NAND3_X1 U218 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n5) );
  NAND2_X1 U219 ( .A1(n13), .A2(n209), .ZN(n248) );
  NAND2_X1 U220 ( .A1(n13), .A2(n71), .ZN(n249) );
  NAND2_X1 U221 ( .A1(n209), .A2(n71), .ZN(n250) );
  NAND3_X1 U222 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n12) );
  NAND2_X2 U223 ( .A1(n290), .A2(n328), .ZN(n292) );
  XOR2_X1 U224 ( .A(n46), .B(n49), .Z(n251) );
  XOR2_X1 U225 ( .A(n234), .B(n251), .Z(product[6]) );
  NAND2_X1 U226 ( .A1(n234), .A2(n46), .ZN(n252) );
  NAND2_X1 U227 ( .A1(n10), .A2(n49), .ZN(n253) );
  NAND2_X1 U228 ( .A1(n46), .A2(n49), .ZN(n254) );
  NAND3_X1 U229 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n9) );
  XOR2_X1 U230 ( .A(n17), .B(n273), .Z(n255) );
  XOR2_X1 U231 ( .A(n211), .B(n255), .Z(product[13]) );
  NAND2_X1 U232 ( .A1(n210), .A2(n17), .ZN(n256) );
  NAND2_X1 U233 ( .A1(n3), .A2(n273), .ZN(n257) );
  NAND2_X1 U234 ( .A1(n17), .A2(n273), .ZN(n258) );
  NAND3_X1 U235 ( .A1(n256), .A2(n257), .A3(n258), .ZN(n2) );
  NAND2_X1 U236 ( .A1(n54), .A2(n55), .ZN(n259) );
  NAND2_X1 U237 ( .A1(n54), .A2(n12), .ZN(n260) );
  NAND2_X1 U238 ( .A1(n55), .A2(n12), .ZN(n261) );
  NAND3_X1 U239 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n11) );
  NAND2_X1 U240 ( .A1(n50), .A2(n53), .ZN(n262) );
  NAND2_X1 U241 ( .A1(n50), .A2(n213), .ZN(n263) );
  NAND2_X1 U242 ( .A1(n53), .A2(n11), .ZN(n264) );
  NAND3_X1 U243 ( .A1(n262), .A2(n263), .A3(n264), .ZN(n10) );
  INV_X1 U244 ( .A(n272), .ZN(n265) );
  NAND2_X1 U245 ( .A1(n269), .A2(n270), .ZN(n266) );
  NAND2_X1 U246 ( .A1(n269), .A2(n270), .ZN(n267) );
  NAND2_X1 U247 ( .A1(n269), .A2(n270), .ZN(n290) );
  INV_X1 U248 ( .A(a[0]), .ZN(n284) );
  NAND2_X1 U249 ( .A1(a[2]), .A2(a[1]), .ZN(n269) );
  NAND2_X1 U250 ( .A1(n268), .A2(n283), .ZN(n270) );
  INV_X1 U251 ( .A(a[2]), .ZN(n268) );
  INV_X1 U252 ( .A(n21), .ZN(n276) );
  INV_X1 U253 ( .A(n309), .ZN(n277) );
  INV_X1 U254 ( .A(n320), .ZN(n274) );
  INV_X1 U255 ( .A(n289), .ZN(n282) );
  INV_X1 U256 ( .A(n298), .ZN(n280) );
  INV_X1 U257 ( .A(n31), .ZN(n279) );
  INV_X1 U258 ( .A(b[0]), .ZN(n272) );
  INV_X1 U259 ( .A(a[5]), .ZN(n278) );
  INV_X1 U260 ( .A(a[7]), .ZN(n275) );
  INV_X1 U261 ( .A(a[3]), .ZN(n281) );
  INV_X1 U262 ( .A(a[1]), .ZN(n283) );
  INV_X1 U263 ( .A(n272), .ZN(n271) );
  NOR2_X1 U264 ( .A1(n284), .A2(n272), .ZN(product[0]) );
  OAI22_X1 U265 ( .A1(n285), .A2(n286), .B1(n287), .B2(n284), .ZN(n99) );
  OAI22_X1 U266 ( .A1(n287), .A2(n286), .B1(n288), .B2(n284), .ZN(n98) );
  XNOR2_X1 U267 ( .A(b[6]), .B(a[1]), .ZN(n287) );
  OAI22_X1 U268 ( .A1(n284), .A2(n288), .B1(n286), .B2(n288), .ZN(n289) );
  XNOR2_X1 U269 ( .A(b[7]), .B(a[1]), .ZN(n288) );
  NOR2_X1 U270 ( .A1(n267), .A2(n272), .ZN(n96) );
  OAI22_X1 U271 ( .A1(n291), .A2(n292), .B1(n266), .B2(n293), .ZN(n95) );
  XNOR2_X1 U272 ( .A(a[3]), .B(n271), .ZN(n291) );
  OAI22_X1 U273 ( .A1(n293), .A2(n292), .B1(n266), .B2(n294), .ZN(n94) );
  XNOR2_X1 U274 ( .A(b[1]), .B(a[3]), .ZN(n293) );
  OAI22_X1 U275 ( .A1(n294), .A2(n292), .B1(n266), .B2(n295), .ZN(n93) );
  XNOR2_X1 U276 ( .A(b[2]), .B(a[3]), .ZN(n294) );
  OAI22_X1 U277 ( .A1(n295), .A2(n292), .B1(n267), .B2(n296), .ZN(n92) );
  XNOR2_X1 U278 ( .A(b[3]), .B(a[3]), .ZN(n295) );
  OAI22_X1 U279 ( .A1(n296), .A2(n292), .B1(n267), .B2(n297), .ZN(n91) );
  XNOR2_X1 U280 ( .A(b[4]), .B(a[3]), .ZN(n296) );
  OAI22_X1 U281 ( .A1(n299), .A2(n266), .B1(n292), .B2(n299), .ZN(n298) );
  NOR2_X1 U282 ( .A1(n300), .A2(n272), .ZN(n88) );
  OAI22_X1 U283 ( .A1(n301), .A2(n302), .B1(n300), .B2(n303), .ZN(n87) );
  XNOR2_X1 U284 ( .A(a[5]), .B(n271), .ZN(n301) );
  OAI22_X1 U285 ( .A1(n303), .A2(n302), .B1(n300), .B2(n304), .ZN(n86) );
  XNOR2_X1 U286 ( .A(b[1]), .B(a[5]), .ZN(n303) );
  OAI22_X1 U287 ( .A1(n304), .A2(n302), .B1(n300), .B2(n305), .ZN(n85) );
  XNOR2_X1 U288 ( .A(b[2]), .B(a[5]), .ZN(n304) );
  OAI22_X1 U289 ( .A1(n305), .A2(n302), .B1(n300), .B2(n306), .ZN(n84) );
  XNOR2_X1 U290 ( .A(b[3]), .B(a[5]), .ZN(n305) );
  OAI22_X1 U291 ( .A1(n306), .A2(n302), .B1(n300), .B2(n307), .ZN(n83) );
  XNOR2_X1 U292 ( .A(b[4]), .B(a[5]), .ZN(n306) );
  OAI22_X1 U293 ( .A1(n307), .A2(n302), .B1(n300), .B2(n308), .ZN(n82) );
  XNOR2_X1 U294 ( .A(b[5]), .B(a[5]), .ZN(n307) );
  OAI22_X1 U295 ( .A1(n310), .A2(n300), .B1(n302), .B2(n310), .ZN(n309) );
  NOR2_X1 U296 ( .A1(n311), .A2(n272), .ZN(n80) );
  OAI22_X1 U297 ( .A1(n312), .A2(n313), .B1(n311), .B2(n314), .ZN(n79) );
  XNOR2_X1 U298 ( .A(a[7]), .B(n265), .ZN(n312) );
  OAI22_X1 U299 ( .A1(n315), .A2(n313), .B1(n311), .B2(n316), .ZN(n77) );
  OAI22_X1 U300 ( .A1(n316), .A2(n313), .B1(n311), .B2(n317), .ZN(n76) );
  XNOR2_X1 U301 ( .A(b[3]), .B(a[7]), .ZN(n316) );
  OAI22_X1 U302 ( .A1(n317), .A2(n313), .B1(n311), .B2(n318), .ZN(n75) );
  XNOR2_X1 U303 ( .A(b[4]), .B(a[7]), .ZN(n317) );
  OAI22_X1 U304 ( .A1(n318), .A2(n313), .B1(n311), .B2(n319), .ZN(n74) );
  XNOR2_X1 U305 ( .A(b[5]), .B(a[7]), .ZN(n318) );
  OAI22_X1 U306 ( .A1(n321), .A2(n311), .B1(n313), .B2(n321), .ZN(n320) );
  OAI21_X1 U307 ( .B1(n265), .B2(n283), .A(n286), .ZN(n72) );
  OAI21_X1 U308 ( .B1(n281), .B2(n292), .A(n322), .ZN(n71) );
  OR3_X1 U309 ( .A1(n267), .A2(n265), .A3(n281), .ZN(n322) );
  OAI21_X1 U310 ( .B1(n278), .B2(n302), .A(n323), .ZN(n70) );
  OAI21_X1 U311 ( .B1(n275), .B2(n313), .A(n324), .ZN(n69) );
  OR3_X1 U312 ( .A1(n311), .A2(n271), .A3(n275), .ZN(n324) );
  XNOR2_X1 U313 ( .A(n325), .B(n326), .ZN(n38) );
  OR2_X1 U314 ( .A1(n325), .A2(n326), .ZN(n37) );
  OAI22_X1 U315 ( .A1(n297), .A2(n292), .B1(n266), .B2(n327), .ZN(n326) );
  XNOR2_X1 U316 ( .A(b[5]), .B(a[3]), .ZN(n297) );
  OAI22_X1 U317 ( .A1(n314), .A2(n313), .B1(n311), .B2(n315), .ZN(n325) );
  XNOR2_X1 U318 ( .A(b[2]), .B(a[7]), .ZN(n315) );
  XNOR2_X1 U319 ( .A(b[1]), .B(a[7]), .ZN(n314) );
  OAI22_X1 U320 ( .A1(n327), .A2(n292), .B1(n267), .B2(n299), .ZN(n31) );
  XNOR2_X1 U321 ( .A(b[7]), .B(a[3]), .ZN(n299) );
  XNOR2_X1 U322 ( .A(n281), .B(a[2]), .ZN(n328) );
  XNOR2_X1 U323 ( .A(b[6]), .B(a[3]), .ZN(n327) );
  OAI22_X1 U324 ( .A1(n308), .A2(n302), .B1(n300), .B2(n310), .ZN(n21) );
  XNOR2_X1 U325 ( .A(b[7]), .B(a[5]), .ZN(n310) );
  XNOR2_X1 U326 ( .A(n278), .B(a[4]), .ZN(n329) );
  XNOR2_X1 U327 ( .A(b[6]), .B(a[5]), .ZN(n308) );
  OAI22_X1 U328 ( .A1(n319), .A2(n313), .B1(n311), .B2(n321), .ZN(n15) );
  XNOR2_X1 U329 ( .A(b[7]), .B(a[7]), .ZN(n321) );
  NAND2_X1 U330 ( .A1(n311), .A2(n330), .ZN(n313) );
  XNOR2_X1 U331 ( .A(n275), .B(a[6]), .ZN(n330) );
  XNOR2_X1 U332 ( .A(b[6]), .B(a[7]), .ZN(n319) );
  OAI22_X1 U333 ( .A1(n271), .A2(n286), .B1(n331), .B2(n284), .ZN(n104) );
  OAI22_X1 U334 ( .A1(n331), .A2(n286), .B1(n332), .B2(n284), .ZN(n103) );
  XNOR2_X1 U335 ( .A(b[1]), .B(a[1]), .ZN(n331) );
  OAI22_X1 U336 ( .A1(n332), .A2(n286), .B1(n333), .B2(n284), .ZN(n102) );
  XNOR2_X1 U337 ( .A(b[2]), .B(a[1]), .ZN(n332) );
  OAI22_X1 U338 ( .A1(n333), .A2(n286), .B1(n334), .B2(n284), .ZN(n101) );
  XNOR2_X1 U339 ( .A(b[3]), .B(a[1]), .ZN(n333) );
  OAI22_X1 U340 ( .A1(n334), .A2(n286), .B1(n285), .B2(n284), .ZN(n100) );
  XNOR2_X1 U341 ( .A(b[5]), .B(a[1]), .ZN(n285) );
  NAND2_X1 U342 ( .A1(a[1]), .A2(n284), .ZN(n286) );
  XNOR2_X1 U343 ( .A(b[4]), .B(a[1]), .ZN(n334) );
endmodule


module datapath_DW01_add_10 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n69;
  wire   [15:1] carry;

  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n69), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[14]), .ZN(n18) );
  XOR2_X1 U2 ( .A(B[9]), .B(A[9]), .Z(n1) );
  XOR2_X1 U3 ( .A(carry[9]), .B(n1), .Z(SUM[9]) );
  NAND2_X1 U4 ( .A1(carry[9]), .A2(B[9]), .ZN(n2) );
  NAND2_X1 U5 ( .A1(carry[9]), .A2(A[9]), .ZN(n3) );
  NAND2_X1 U6 ( .A1(B[9]), .A2(A[9]), .ZN(n4) );
  NAND3_X1 U7 ( .A1(n2), .A2(n3), .A3(n4), .ZN(carry[10]) );
  CLKBUF_X1 U8 ( .A(n17), .Z(n5) );
  NAND3_X1 U9 ( .A1(n8), .A2(n9), .A3(n10), .ZN(n6) );
  XOR2_X1 U10 ( .A(B[10]), .B(A[10]), .Z(n7) );
  XOR2_X1 U11 ( .A(carry[10]), .B(n7), .Z(SUM[10]) );
  NAND2_X1 U12 ( .A1(carry[10]), .A2(B[10]), .ZN(n8) );
  NAND2_X1 U13 ( .A1(carry[10]), .A2(A[10]), .ZN(n9) );
  NAND2_X1 U14 ( .A1(B[10]), .A2(A[10]), .ZN(n10) );
  NAND3_X1 U15 ( .A1(n8), .A2(n9), .A3(n10), .ZN(carry[11]) );
  NAND3_X1 U16 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n11) );
  NAND3_X1 U17 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n12) );
  XOR2_X1 U18 ( .A(carry[2]), .B(A[2]), .Z(n13) );
  XOR2_X1 U19 ( .A(B[2]), .B(n13), .Z(SUM[2]) );
  NAND2_X1 U20 ( .A1(B[2]), .A2(carry[2]), .ZN(n14) );
  NAND2_X1 U21 ( .A1(B[2]), .A2(A[2]), .ZN(n15) );
  NAND2_X1 U22 ( .A1(carry[2]), .A2(A[2]), .ZN(n16) );
  NAND3_X1 U23 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[3]) );
  NAND3_X1 U24 ( .A1(n20), .A2(n21), .A3(n22), .ZN(n17) );
  XNOR2_X1 U25 ( .A(B[14]), .B(n18), .ZN(n28) );
  XOR2_X1 U26 ( .A(B[11]), .B(A[11]), .Z(n19) );
  XOR2_X1 U27 ( .A(n6), .B(n19), .Z(SUM[11]) );
  NAND2_X1 U28 ( .A1(n6), .A2(B[11]), .ZN(n20) );
  NAND2_X1 U29 ( .A1(carry[11]), .A2(A[11]), .ZN(n21) );
  NAND2_X1 U30 ( .A1(B[11]), .A2(A[11]), .ZN(n22) );
  NAND3_X1 U31 ( .A1(n20), .A2(n21), .A3(n22), .ZN(carry[12]) );
  NAND3_X1 U32 ( .A1(n48), .A2(n49), .A3(n50), .ZN(n23) );
  NAND3_X1 U33 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n24) );
  CLKBUF_X1 U34 ( .A(carry[13]), .Z(n25) );
  NAND3_X1 U35 ( .A1(n57), .A2(n58), .A3(n59), .ZN(n26) );
  NAND3_X1 U36 ( .A1(n57), .A2(n58), .A3(n59), .ZN(n27) );
  XOR2_X1 U37 ( .A(n28), .B(carry[14]), .Z(SUM[14]) );
  NAND2_X1 U38 ( .A1(B[14]), .A2(n23), .ZN(n29) );
  NAND2_X1 U39 ( .A1(carry[14]), .A2(A[14]), .ZN(n30) );
  NAND2_X1 U40 ( .A1(B[14]), .A2(A[14]), .ZN(n31) );
  NAND3_X1 U41 ( .A1(n30), .A2(n29), .A3(n31), .ZN(carry[15]) );
  XNOR2_X1 U42 ( .A(carry[15]), .B(n32), .ZN(SUM[15]) );
  XNOR2_X1 U43 ( .A(B[15]), .B(A[15]), .ZN(n32) );
  XOR2_X1 U44 ( .A(B[3]), .B(A[3]), .Z(n33) );
  XOR2_X1 U45 ( .A(carry[3]), .B(n33), .Z(SUM[3]) );
  NAND2_X1 U46 ( .A1(carry[3]), .A2(B[3]), .ZN(n34) );
  NAND2_X1 U47 ( .A1(carry[3]), .A2(A[3]), .ZN(n35) );
  NAND2_X1 U48 ( .A1(B[3]), .A2(A[3]), .ZN(n36) );
  NAND3_X1 U49 ( .A1(n34), .A2(n35), .A3(n36), .ZN(carry[4]) );
  XOR2_X1 U50 ( .A(B[12]), .B(A[12]), .Z(n37) );
  XOR2_X1 U51 ( .A(n5), .B(n37), .Z(SUM[12]) );
  NAND2_X1 U52 ( .A1(n17), .A2(B[12]), .ZN(n38) );
  NAND2_X1 U53 ( .A1(carry[12]), .A2(A[12]), .ZN(n39) );
  NAND2_X1 U54 ( .A1(B[12]), .A2(A[12]), .ZN(n40) );
  NAND3_X1 U55 ( .A1(n38), .A2(n39), .A3(n40), .ZN(carry[13]) );
  XOR2_X1 U56 ( .A(B[7]), .B(A[7]), .Z(n41) );
  XOR2_X1 U57 ( .A(n11), .B(n41), .Z(SUM[7]) );
  NAND2_X1 U58 ( .A1(n11), .A2(B[7]), .ZN(n42) );
  NAND2_X1 U59 ( .A1(carry[7]), .A2(A[7]), .ZN(n43) );
  NAND2_X1 U60 ( .A1(B[7]), .A2(A[7]), .ZN(n44) );
  NAND3_X1 U61 ( .A1(n42), .A2(n43), .A3(n44), .ZN(carry[8]) );
  NAND3_X1 U62 ( .A1(n63), .A2(n62), .A3(n61), .ZN(n45) );
  NAND3_X1 U63 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n46) );
  XOR2_X1 U64 ( .A(B[13]), .B(A[13]), .Z(n47) );
  XOR2_X1 U65 ( .A(n25), .B(n47), .Z(SUM[13]) );
  NAND2_X1 U66 ( .A1(carry[13]), .A2(B[13]), .ZN(n48) );
  NAND2_X1 U67 ( .A1(carry[13]), .A2(A[13]), .ZN(n49) );
  NAND2_X1 U68 ( .A1(B[13]), .A2(A[13]), .ZN(n50) );
  NAND3_X1 U69 ( .A1(n48), .A2(n49), .A3(n50), .ZN(carry[14]) );
  XOR2_X1 U70 ( .A(B[8]), .B(A[8]), .Z(n51) );
  XOR2_X1 U71 ( .A(carry[8]), .B(n51), .Z(SUM[8]) );
  NAND2_X1 U72 ( .A1(n24), .A2(B[8]), .ZN(n52) );
  NAND2_X1 U73 ( .A1(carry[8]), .A2(A[8]), .ZN(n53) );
  NAND2_X1 U74 ( .A1(B[8]), .A2(A[8]), .ZN(n54) );
  NAND3_X1 U75 ( .A1(n52), .A2(n53), .A3(n54), .ZN(carry[9]) );
  CLKBUF_X1 U76 ( .A(n12), .Z(n55) );
  XOR2_X1 U77 ( .A(B[4]), .B(A[4]), .Z(n56) );
  XOR2_X1 U78 ( .A(n55), .B(n56), .Z(SUM[4]) );
  NAND2_X1 U79 ( .A1(n12), .A2(B[4]), .ZN(n57) );
  NAND2_X1 U80 ( .A1(carry[4]), .A2(A[4]), .ZN(n58) );
  NAND2_X1 U81 ( .A1(B[4]), .A2(A[4]), .ZN(n59) );
  NAND3_X1 U82 ( .A1(n57), .A2(n58), .A3(n59), .ZN(carry[5]) );
  XOR2_X1 U83 ( .A(A[5]), .B(B[5]), .Z(n60) );
  XOR2_X1 U84 ( .A(n60), .B(n27), .Z(SUM[5]) );
  NAND2_X1 U85 ( .A1(B[5]), .A2(A[5]), .ZN(n61) );
  NAND2_X1 U86 ( .A1(A[5]), .A2(carry[5]), .ZN(n62) );
  NAND2_X1 U87 ( .A1(B[5]), .A2(n26), .ZN(n63) );
  NAND3_X1 U88 ( .A1(n61), .A2(n62), .A3(n63), .ZN(carry[6]) );
  XOR2_X1 U89 ( .A(A[6]), .B(B[6]), .Z(n64) );
  XOR2_X1 U90 ( .A(n64), .B(n46), .Z(SUM[6]) );
  NAND2_X1 U91 ( .A1(A[6]), .A2(B[6]), .ZN(n65) );
  NAND2_X1 U92 ( .A1(A[6]), .A2(n45), .ZN(n66) );
  NAND2_X1 U93 ( .A1(B[6]), .A2(carry[6]), .ZN(n67) );
  NAND3_X1 U94 ( .A1(n65), .A2(n66), .A3(n67), .ZN(carry[7]) );
  XOR2_X1 U95 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U96 ( .A1(B[0]), .A2(A[0]), .ZN(n69) );
endmodule


module datapath_DW_mult_tc_9 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331;

  FA_X1 U11 ( .A(n50), .B(n53), .CI(n11), .CO(n10), .S(product[5]) );
  FA_X1 U12 ( .A(n54), .B(n206), .CI(n12), .CO(n11), .S(product[4]) );
  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  FA_X1 U14 ( .A(n103), .B(n96), .CI(n14), .CO(n13), .S(product[2]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n274), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n273), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n277), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n276), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n279), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  AND2_X1 U157 ( .A1(n95), .A2(n102), .ZN(n206) );
  XNOR2_X1 U158 ( .A(n271), .B(n15), .ZN(n207) );
  AND3_X1 U159 ( .A1(n246), .A2(n247), .A3(n248), .ZN(product[15]) );
  NAND3_X1 U160 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n209) );
  NAND3_X1 U161 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n210) );
  NAND3_X1 U162 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n211) );
  NAND3_X1 U163 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n212) );
  NAND3_X1 U164 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n213) );
  NAND3_X1 U165 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n214) );
  INV_X2 U166 ( .A(a[0]), .ZN(n281) );
  NAND3_X1 U167 ( .A1(n220), .A2(n221), .A3(n222), .ZN(n215) );
  NAND3_X1 U168 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n216) );
  NAND3_X1 U169 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n217) );
  CLKBUF_X1 U170 ( .A(b[3]), .Z(n218) );
  XOR2_X1 U171 ( .A(n19), .B(n18), .Z(n219) );
  XOR2_X1 U172 ( .A(n219), .B(n214), .Z(product[12]) );
  NAND2_X1 U173 ( .A1(n19), .A2(n18), .ZN(n220) );
  NAND2_X1 U174 ( .A1(n19), .A2(n213), .ZN(n221) );
  NAND2_X1 U175 ( .A1(n18), .A2(n4), .ZN(n222) );
  NAND3_X1 U176 ( .A1(n220), .A2(n221), .A3(n222), .ZN(n3) );
  XOR2_X1 U177 ( .A(n17), .B(n270), .Z(n223) );
  XOR2_X1 U178 ( .A(n223), .B(n215), .Z(product[13]) );
  NAND2_X1 U179 ( .A1(n17), .A2(n270), .ZN(n224) );
  NAND2_X1 U180 ( .A1(n17), .A2(n3), .ZN(n225) );
  NAND2_X1 U181 ( .A1(n270), .A2(n3), .ZN(n226) );
  NAND3_X1 U182 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n2) );
  XOR2_X1 U183 ( .A(n33), .B(n28), .Z(n227) );
  XOR2_X1 U184 ( .A(n7), .B(n227), .Z(product[9]) );
  NAND2_X1 U185 ( .A1(n7), .A2(n33), .ZN(n228) );
  NAND2_X1 U186 ( .A1(n7), .A2(n28), .ZN(n229) );
  NAND2_X1 U187 ( .A1(n33), .A2(n28), .ZN(n230) );
  NAND3_X1 U188 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n6) );
  XOR2_X1 U189 ( .A(n46), .B(n49), .Z(n231) );
  XOR2_X1 U190 ( .A(n231), .B(n10), .Z(product[6]) );
  NAND2_X1 U191 ( .A1(n46), .A2(n49), .ZN(n232) );
  NAND2_X1 U192 ( .A1(n46), .A2(n10), .ZN(n233) );
  NAND2_X1 U193 ( .A1(n49), .A2(n10), .ZN(n234) );
  NAND3_X1 U194 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n9) );
  XOR2_X1 U195 ( .A(n40), .B(n45), .Z(n235) );
  XOR2_X1 U196 ( .A(n235), .B(n217), .Z(product[7]) );
  NAND2_X1 U197 ( .A1(n40), .A2(n45), .ZN(n236) );
  NAND2_X1 U198 ( .A1(n40), .A2(n216), .ZN(n237) );
  NAND2_X1 U199 ( .A1(n45), .A2(n9), .ZN(n238) );
  NAND3_X1 U200 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n8) );
  NAND2_X2 U201 ( .A1(n287), .A2(n325), .ZN(n289) );
  INV_X1 U202 ( .A(n269), .ZN(n239) );
  INV_X1 U203 ( .A(n269), .ZN(n268) );
  XOR2_X1 U204 ( .A(n34), .B(n39), .Z(n240) );
  XOR2_X1 U205 ( .A(n210), .B(n240), .Z(product[8]) );
  NAND2_X1 U206 ( .A1(n209), .A2(n34), .ZN(n241) );
  NAND2_X1 U207 ( .A1(n8), .A2(n39), .ZN(n242) );
  NAND2_X1 U208 ( .A1(n34), .A2(n39), .ZN(n243) );
  NAND3_X1 U209 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n7) );
  XOR2_X1 U210 ( .A(a[3]), .B(n269), .Z(n288) );
  XNOR2_X1 U211 ( .A(n2), .B(n207), .ZN(product[14]) );
  NAND3_X1 U212 ( .A1(n252), .A2(n251), .A3(n250), .ZN(n244) );
  NAND3_X1 U213 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n245) );
  XOR2_X1 U214 ( .A(n95), .B(n102), .Z(n56) );
  NAND2_X1 U215 ( .A1(n2), .A2(n271), .ZN(n246) );
  NAND2_X1 U216 ( .A1(n2), .A2(n15), .ZN(n247) );
  NAND2_X1 U217 ( .A1(n271), .A2(n15), .ZN(n248) );
  XOR2_X1 U218 ( .A(n24), .B(n27), .Z(n249) );
  XOR2_X1 U219 ( .A(n249), .B(n212), .Z(product[10]) );
  NAND2_X1 U220 ( .A1(n24), .A2(n27), .ZN(n250) );
  NAND2_X1 U221 ( .A1(n24), .A2(n6), .ZN(n251) );
  NAND2_X1 U222 ( .A1(n27), .A2(n211), .ZN(n252) );
  NAND3_X1 U223 ( .A1(n250), .A2(n251), .A3(n252), .ZN(n5) );
  XOR2_X1 U224 ( .A(n20), .B(n23), .Z(n253) );
  XOR2_X1 U225 ( .A(n253), .B(n245), .Z(product[11]) );
  NAND2_X1 U226 ( .A1(n20), .A2(n23), .ZN(n254) );
  NAND2_X1 U227 ( .A1(n20), .A2(n244), .ZN(n255) );
  NAND2_X1 U228 ( .A1(n23), .A2(n5), .ZN(n256) );
  NAND3_X1 U229 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n4) );
  NAND2_X1 U230 ( .A1(a[4]), .A2(a[3]), .ZN(n259) );
  NAND2_X1 U231 ( .A1(n257), .A2(n258), .ZN(n260) );
  NAND2_X2 U232 ( .A1(n259), .A2(n260), .ZN(n297) );
  INV_X1 U233 ( .A(a[4]), .ZN(n257) );
  INV_X1 U234 ( .A(a[3]), .ZN(n258) );
  NAND2_X2 U235 ( .A1(n297), .A2(n326), .ZN(n299) );
  NAND2_X1 U236 ( .A1(n265), .A2(n266), .ZN(n261) );
  NAND2_X1 U237 ( .A1(n265), .A2(n266), .ZN(n262) );
  NAND2_X1 U238 ( .A1(n265), .A2(n266), .ZN(n287) );
  NAND2_X1 U239 ( .A1(a[2]), .A2(a[1]), .ZN(n265) );
  NAND2_X1 U240 ( .A1(n263), .A2(n264), .ZN(n266) );
  INV_X1 U241 ( .A(a[2]), .ZN(n263) );
  INV_X1 U242 ( .A(a[1]), .ZN(n264) );
  INV_X1 U243 ( .A(n15), .ZN(n270) );
  INV_X1 U244 ( .A(n295), .ZN(n277) );
  INV_X1 U245 ( .A(n21), .ZN(n273) );
  INV_X1 U246 ( .A(n306), .ZN(n274) );
  INV_X1 U247 ( .A(n317), .ZN(n271) );
  INV_X1 U248 ( .A(n286), .ZN(n279) );
  INV_X1 U249 ( .A(n31), .ZN(n276) );
  INV_X1 U250 ( .A(b[0]), .ZN(n269) );
  XOR2_X1 U251 ( .A(a[6]), .B(n275), .Z(n308) );
  INV_X1 U252 ( .A(a[5]), .ZN(n275) );
  INV_X1 U253 ( .A(a[7]), .ZN(n272) );
  CLKBUF_X1 U254 ( .A(b[1]), .Z(n267) );
  INV_X1 U255 ( .A(a[3]), .ZN(n278) );
  INV_X1 U256 ( .A(a[1]), .ZN(n280) );
  NOR2_X1 U257 ( .A1(n281), .A2(n269), .ZN(product[0]) );
  OAI22_X1 U258 ( .A1(n282), .A2(n283), .B1(n284), .B2(n281), .ZN(n99) );
  OAI22_X1 U259 ( .A1(n284), .A2(n283), .B1(n285), .B2(n281), .ZN(n98) );
  XNOR2_X1 U260 ( .A(b[6]), .B(a[1]), .ZN(n284) );
  OAI22_X1 U261 ( .A1(n281), .A2(n285), .B1(n283), .B2(n285), .ZN(n286) );
  XNOR2_X1 U262 ( .A(b[7]), .B(a[1]), .ZN(n285) );
  NOR2_X1 U263 ( .A1(n262), .A2(n269), .ZN(n96) );
  OAI22_X1 U264 ( .A1(n288), .A2(n289), .B1(n261), .B2(n290), .ZN(n95) );
  OAI22_X1 U265 ( .A1(n290), .A2(n289), .B1(n261), .B2(n291), .ZN(n94) );
  XNOR2_X1 U266 ( .A(n267), .B(a[3]), .ZN(n290) );
  OAI22_X1 U267 ( .A1(n291), .A2(n289), .B1(n261), .B2(n292), .ZN(n93) );
  XNOR2_X1 U268 ( .A(b[2]), .B(a[3]), .ZN(n291) );
  OAI22_X1 U269 ( .A1(n292), .A2(n289), .B1(n262), .B2(n293), .ZN(n92) );
  XNOR2_X1 U270 ( .A(n218), .B(a[3]), .ZN(n292) );
  OAI22_X1 U271 ( .A1(n293), .A2(n289), .B1(n262), .B2(n294), .ZN(n91) );
  XNOR2_X1 U272 ( .A(b[4]), .B(a[3]), .ZN(n293) );
  OAI22_X1 U273 ( .A1(n296), .A2(n261), .B1(n289), .B2(n296), .ZN(n295) );
  NOR2_X1 U274 ( .A1(n297), .A2(n269), .ZN(n88) );
  OAI22_X1 U275 ( .A1(n298), .A2(n299), .B1(n297), .B2(n300), .ZN(n87) );
  XNOR2_X1 U276 ( .A(a[5]), .B(n239), .ZN(n298) );
  OAI22_X1 U277 ( .A1(n300), .A2(n299), .B1(n297), .B2(n301), .ZN(n86) );
  XNOR2_X1 U278 ( .A(n267), .B(a[5]), .ZN(n300) );
  OAI22_X1 U279 ( .A1(n301), .A2(n299), .B1(n297), .B2(n302), .ZN(n85) );
  XNOR2_X1 U280 ( .A(b[2]), .B(a[5]), .ZN(n301) );
  OAI22_X1 U281 ( .A1(n302), .A2(n299), .B1(n297), .B2(n303), .ZN(n84) );
  XNOR2_X1 U282 ( .A(n218), .B(a[5]), .ZN(n302) );
  OAI22_X1 U283 ( .A1(n303), .A2(n299), .B1(n297), .B2(n304), .ZN(n83) );
  XNOR2_X1 U284 ( .A(b[4]), .B(a[5]), .ZN(n303) );
  OAI22_X1 U285 ( .A1(n304), .A2(n299), .B1(n297), .B2(n305), .ZN(n82) );
  XNOR2_X1 U286 ( .A(b[5]), .B(a[5]), .ZN(n304) );
  OAI22_X1 U287 ( .A1(n307), .A2(n297), .B1(n299), .B2(n307), .ZN(n306) );
  NOR2_X1 U288 ( .A1(n308), .A2(n269), .ZN(n80) );
  OAI22_X1 U289 ( .A1(n309), .A2(n310), .B1(n308), .B2(n311), .ZN(n79) );
  XNOR2_X1 U290 ( .A(a[7]), .B(n239), .ZN(n309) );
  OAI22_X1 U291 ( .A1(n312), .A2(n310), .B1(n308), .B2(n313), .ZN(n77) );
  OAI22_X1 U292 ( .A1(n313), .A2(n310), .B1(n308), .B2(n314), .ZN(n76) );
  XNOR2_X1 U293 ( .A(n218), .B(a[7]), .ZN(n313) );
  OAI22_X1 U294 ( .A1(n314), .A2(n310), .B1(n308), .B2(n315), .ZN(n75) );
  XNOR2_X1 U295 ( .A(b[4]), .B(a[7]), .ZN(n314) );
  OAI22_X1 U296 ( .A1(n315), .A2(n310), .B1(n308), .B2(n316), .ZN(n74) );
  XNOR2_X1 U297 ( .A(b[5]), .B(a[7]), .ZN(n315) );
  OAI22_X1 U298 ( .A1(n318), .A2(n308), .B1(n310), .B2(n318), .ZN(n317) );
  OAI21_X1 U299 ( .B1(n268), .B2(n280), .A(n283), .ZN(n72) );
  OAI21_X1 U300 ( .B1(n278), .B2(n289), .A(n319), .ZN(n71) );
  OR3_X1 U301 ( .A1(n262), .A2(n239), .A3(n278), .ZN(n319) );
  OAI21_X1 U302 ( .B1(n275), .B2(n299), .A(n320), .ZN(n70) );
  OR3_X1 U303 ( .A1(n297), .A2(n268), .A3(n275), .ZN(n320) );
  OAI21_X1 U304 ( .B1(n272), .B2(n310), .A(n321), .ZN(n69) );
  OR3_X1 U305 ( .A1(n308), .A2(n239), .A3(n272), .ZN(n321) );
  XNOR2_X1 U306 ( .A(n322), .B(n323), .ZN(n38) );
  OR2_X1 U307 ( .A1(n322), .A2(n323), .ZN(n37) );
  OAI22_X1 U308 ( .A1(n294), .A2(n289), .B1(n261), .B2(n324), .ZN(n323) );
  XNOR2_X1 U309 ( .A(b[5]), .B(a[3]), .ZN(n294) );
  OAI22_X1 U310 ( .A1(n311), .A2(n310), .B1(n308), .B2(n312), .ZN(n322) );
  XNOR2_X1 U311 ( .A(b[2]), .B(a[7]), .ZN(n312) );
  XNOR2_X1 U312 ( .A(n267), .B(a[7]), .ZN(n311) );
  OAI22_X1 U313 ( .A1(n324), .A2(n289), .B1(n262), .B2(n296), .ZN(n31) );
  XNOR2_X1 U314 ( .A(b[7]), .B(a[3]), .ZN(n296) );
  XNOR2_X1 U315 ( .A(n278), .B(a[2]), .ZN(n325) );
  XNOR2_X1 U316 ( .A(b[6]), .B(a[3]), .ZN(n324) );
  OAI22_X1 U317 ( .A1(n305), .A2(n299), .B1(n297), .B2(n307), .ZN(n21) );
  XNOR2_X1 U318 ( .A(b[7]), .B(a[5]), .ZN(n307) );
  XNOR2_X1 U319 ( .A(n275), .B(a[4]), .ZN(n326) );
  XNOR2_X1 U320 ( .A(b[6]), .B(a[5]), .ZN(n305) );
  OAI22_X1 U321 ( .A1(n316), .A2(n310), .B1(n308), .B2(n318), .ZN(n15) );
  XNOR2_X1 U322 ( .A(b[7]), .B(a[7]), .ZN(n318) );
  NAND2_X1 U323 ( .A1(n327), .A2(n308), .ZN(n310) );
  XNOR2_X1 U324 ( .A(n272), .B(a[6]), .ZN(n327) );
  XNOR2_X1 U325 ( .A(b[6]), .B(a[7]), .ZN(n316) );
  OAI22_X1 U326 ( .A1(n268), .A2(n283), .B1(n328), .B2(n281), .ZN(n104) );
  OAI22_X1 U327 ( .A1(n328), .A2(n283), .B1(n329), .B2(n281), .ZN(n103) );
  XNOR2_X1 U328 ( .A(b[1]), .B(a[1]), .ZN(n328) );
  OAI22_X1 U329 ( .A1(n283), .A2(n329), .B1(n330), .B2(n281), .ZN(n102) );
  XNOR2_X1 U330 ( .A(b[2]), .B(a[1]), .ZN(n329) );
  OAI22_X1 U331 ( .A1(n330), .A2(n283), .B1(n331), .B2(n281), .ZN(n101) );
  XNOR2_X1 U332 ( .A(b[3]), .B(a[1]), .ZN(n330) );
  OAI22_X1 U333 ( .A1(n331), .A2(n283), .B1(n282), .B2(n281), .ZN(n100) );
  XNOR2_X1 U334 ( .A(b[5]), .B(a[1]), .ZN(n282) );
  NAND2_X1 U335 ( .A1(a[1]), .A2(n281), .ZN(n283) );
  XNOR2_X1 U336 ( .A(b[4]), .B(a[1]), .ZN(n331) );
endmodule


module datapath_DW01_add_9 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n68;
  wire   [15:1] carry;

  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n68), .CO(carry[2]), .S(SUM[1]) );
  CLKBUF_X1 U1 ( .A(carry[6]), .Z(n1) );
  XOR2_X1 U2 ( .A(carry[2]), .B(A[2]), .Z(n2) );
  XOR2_X1 U3 ( .A(B[2]), .B(n2), .Z(SUM[2]) );
  NAND2_X1 U4 ( .A1(B[2]), .A2(carry[2]), .ZN(n3) );
  NAND2_X1 U5 ( .A1(B[2]), .A2(A[2]), .ZN(n4) );
  NAND2_X1 U6 ( .A1(carry[2]), .A2(A[2]), .ZN(n5) );
  NAND3_X1 U7 ( .A1(n3), .A2(n4), .A3(n5), .ZN(carry[3]) );
  CLKBUF_X1 U8 ( .A(n33), .Z(n6) );
  CLKBUF_X1 U9 ( .A(n53), .Z(n7) );
  NAND3_X1 U10 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n8) );
  NAND3_X1 U11 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n9) );
  NAND3_X1 U12 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n10) );
  XOR2_X1 U13 ( .A(B[3]), .B(A[3]), .Z(n11) );
  XOR2_X1 U14 ( .A(n11), .B(carry[3]), .Z(SUM[3]) );
  NAND2_X1 U15 ( .A1(B[3]), .A2(A[3]), .ZN(n12) );
  NAND2_X1 U16 ( .A1(B[3]), .A2(carry[3]), .ZN(n13) );
  NAND2_X1 U17 ( .A1(A[3]), .A2(carry[3]), .ZN(n14) );
  NAND3_X1 U18 ( .A1(n12), .A2(n13), .A3(n14), .ZN(carry[4]) );
  XOR2_X1 U19 ( .A(A[4]), .B(B[4]), .Z(n15) );
  XOR2_X1 U20 ( .A(n15), .B(carry[4]), .Z(SUM[4]) );
  NAND2_X1 U21 ( .A1(A[4]), .A2(B[4]), .ZN(n16) );
  NAND2_X1 U22 ( .A1(A[4]), .A2(carry[4]), .ZN(n17) );
  NAND2_X1 U23 ( .A1(B[4]), .A2(carry[4]), .ZN(n18) );
  NAND3_X1 U24 ( .A1(n16), .A2(n17), .A3(n18), .ZN(carry[5]) );
  CLKBUF_X1 U25 ( .A(n26), .Z(n19) );
  XOR2_X1 U26 ( .A(B[6]), .B(A[6]), .Z(n20) );
  XOR2_X1 U27 ( .A(n1), .B(n20), .Z(SUM[6]) );
  NAND2_X1 U28 ( .A1(carry[6]), .A2(B[6]), .ZN(n21) );
  NAND2_X1 U29 ( .A1(carry[6]), .A2(A[6]), .ZN(n22) );
  NAND2_X1 U30 ( .A1(B[6]), .A2(A[6]), .ZN(n23) );
  NAND3_X1 U31 ( .A1(n21), .A2(n22), .A3(n23), .ZN(carry[7]) );
  NAND3_X1 U32 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n24) );
  NAND3_X1 U33 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n25) );
  NAND3_X1 U34 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n26) );
  NAND3_X1 U35 ( .A1(n30), .A2(n31), .A3(n32), .ZN(n27) );
  XNOR2_X1 U36 ( .A(n49), .B(n28), .ZN(SUM[14]) );
  XNOR2_X1 U37 ( .A(B[14]), .B(A[14]), .ZN(n28) );
  XOR2_X1 U38 ( .A(B[12]), .B(A[12]), .Z(n29) );
  XOR2_X1 U39 ( .A(n25), .B(n29), .Z(SUM[12]) );
  NAND2_X1 U40 ( .A1(n24), .A2(B[12]), .ZN(n30) );
  NAND2_X1 U41 ( .A1(carry[12]), .A2(A[12]), .ZN(n31) );
  NAND2_X1 U42 ( .A1(B[12]), .A2(A[12]), .ZN(n32) );
  NAND3_X1 U43 ( .A1(n31), .A2(n30), .A3(n32), .ZN(carry[13]) );
  NAND3_X1 U44 ( .A1(n41), .A2(n42), .A3(n43), .ZN(n33) );
  NAND3_X1 U45 ( .A1(n54), .A2(n53), .A3(n52), .ZN(n34) );
  NAND3_X1 U46 ( .A1(n52), .A2(n7), .A3(n54), .ZN(n35) );
  XOR2_X1 U47 ( .A(B[9]), .B(A[9]), .Z(n36) );
  XOR2_X1 U48 ( .A(n19), .B(n36), .Z(SUM[9]) );
  NAND2_X1 U49 ( .A1(n26), .A2(B[9]), .ZN(n37) );
  NAND2_X1 U50 ( .A1(carry[9]), .A2(A[9]), .ZN(n38) );
  NAND2_X1 U51 ( .A1(B[9]), .A2(A[9]), .ZN(n39) );
  NAND3_X1 U52 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[10]) );
  XOR2_X1 U53 ( .A(B[7]), .B(A[7]), .Z(n40) );
  XOR2_X1 U54 ( .A(n10), .B(n40), .Z(SUM[7]) );
  NAND2_X1 U55 ( .A1(n9), .A2(B[7]), .ZN(n41) );
  NAND2_X1 U56 ( .A1(carry[7]), .A2(A[7]), .ZN(n42) );
  NAND2_X1 U57 ( .A1(B[7]), .A2(A[7]), .ZN(n43) );
  NAND3_X1 U58 ( .A1(n42), .A2(n41), .A3(n43), .ZN(carry[8]) );
  XNOR2_X1 U59 ( .A(carry[15]), .B(n44), .ZN(SUM[15]) );
  XNOR2_X1 U60 ( .A(B[15]), .B(A[15]), .ZN(n44) );
  XOR2_X1 U61 ( .A(B[8]), .B(A[8]), .Z(n45) );
  XOR2_X1 U62 ( .A(n6), .B(n45), .Z(SUM[8]) );
  NAND2_X1 U63 ( .A1(n33), .A2(B[8]), .ZN(n46) );
  NAND2_X1 U64 ( .A1(carry[8]), .A2(A[8]), .ZN(n47) );
  NAND2_X1 U65 ( .A1(B[8]), .A2(A[8]), .ZN(n48) );
  NAND3_X1 U66 ( .A1(n46), .A2(n47), .A3(n48), .ZN(carry[9]) );
  CLKBUF_X1 U67 ( .A(n59), .Z(n49) );
  CLKBUF_X1 U68 ( .A(n8), .Z(n50) );
  XOR2_X1 U69 ( .A(A[10]), .B(B[10]), .Z(n51) );
  XOR2_X1 U70 ( .A(n51), .B(n50), .Z(SUM[10]) );
  NAND2_X1 U71 ( .A1(A[10]), .A2(B[10]), .ZN(n52) );
  NAND2_X1 U72 ( .A1(A[10]), .A2(n8), .ZN(n53) );
  NAND2_X1 U73 ( .A1(B[10]), .A2(carry[10]), .ZN(n54) );
  NAND3_X1 U74 ( .A1(n52), .A2(n53), .A3(n54), .ZN(carry[11]) );
  XOR2_X1 U75 ( .A(A[11]), .B(B[11]), .Z(n55) );
  XOR2_X1 U76 ( .A(n55), .B(n35), .Z(SUM[11]) );
  NAND2_X1 U77 ( .A1(A[11]), .A2(B[11]), .ZN(n56) );
  NAND2_X1 U78 ( .A1(A[11]), .A2(n34), .ZN(n57) );
  NAND2_X1 U79 ( .A1(B[11]), .A2(carry[11]), .ZN(n58) );
  NAND3_X1 U80 ( .A1(n56), .A2(n57), .A3(n58), .ZN(carry[12]) );
  NAND3_X1 U81 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n59) );
  XOR2_X1 U82 ( .A(B[13]), .B(A[13]), .Z(n60) );
  XOR2_X1 U83 ( .A(n27), .B(n60), .Z(SUM[13]) );
  NAND2_X1 U84 ( .A1(n27), .A2(B[13]), .ZN(n61) );
  NAND2_X1 U85 ( .A1(carry[13]), .A2(A[13]), .ZN(n62) );
  NAND2_X1 U86 ( .A1(B[13]), .A2(A[13]), .ZN(n63) );
  NAND3_X1 U87 ( .A1(n61), .A2(n62), .A3(n63), .ZN(carry[14]) );
  NAND2_X1 U88 ( .A1(n59), .A2(B[14]), .ZN(n64) );
  NAND2_X1 U89 ( .A1(carry[14]), .A2(A[14]), .ZN(n65) );
  NAND2_X1 U90 ( .A1(B[14]), .A2(A[14]), .ZN(n66) );
  NAND3_X1 U91 ( .A1(n64), .A2(n65), .A3(n66), .ZN(carry[15]) );
  XOR2_X1 U92 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U93 ( .A1(B[0]), .A2(A[0]), .ZN(n68) );
endmodule


module datapath_DW_mult_tc_8 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340;

  FA_X1 U7 ( .A(n28), .B(n33), .CI(n7), .CO(n6), .S(product[9]) );
  FA_X1 U11 ( .A(n50), .B(n53), .CI(n11), .CO(n10), .S(product[5]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n284), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n283), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n287), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n286), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n288), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n94), .B(n88), .CI(n101), .CO(n53), .S(n54) );
  BUF_X2 U157 ( .A(n308), .Z(n206) );
  NAND2_X1 U158 ( .A1(n306), .A2(n335), .ZN(n308) );
  INV_X1 U159 ( .A(n15), .ZN(n280) );
  AND2_X1 U160 ( .A1(n211), .A2(n102), .ZN(n207) );
  XNOR2_X1 U161 ( .A(n281), .B(n15), .ZN(n208) );
  AND3_X1 U162 ( .A1(n250), .A2(n251), .A3(n252), .ZN(product[15]) );
  NAND2_X2 U163 ( .A1(n259), .A2(n260), .ZN(n210) );
  NAND2_X1 U164 ( .A1(n259), .A2(n260), .ZN(n306) );
  OAI22_X1 U165 ( .A1(n297), .A2(n298), .B1(n296), .B2(n299), .ZN(n211) );
  CLKBUF_X1 U166 ( .A(b[1]), .Z(n275) );
  CLKBUF_X1 U167 ( .A(n264), .Z(n212) );
  NAND2_X1 U168 ( .A1(n296), .A2(n334), .ZN(n213) );
  NAND2_X1 U169 ( .A1(n296), .A2(n334), .ZN(n298) );
  XOR2_X2 U170 ( .A(a[2]), .B(n289), .Z(n296) );
  XOR2_X1 U171 ( .A(n34), .B(n39), .Z(n214) );
  XOR2_X1 U172 ( .A(n8), .B(n214), .Z(product[8]) );
  NAND2_X1 U173 ( .A1(n8), .A2(n34), .ZN(n215) );
  NAND2_X1 U174 ( .A1(n8), .A2(n39), .ZN(n216) );
  NAND2_X1 U175 ( .A1(n34), .A2(n39), .ZN(n217) );
  NAND3_X1 U176 ( .A1(n215), .A2(n216), .A3(n217), .ZN(n7) );
  XOR2_X1 U177 ( .A(n19), .B(n18), .Z(n218) );
  XOR2_X1 U178 ( .A(n4), .B(n218), .Z(product[12]) );
  NAND2_X1 U179 ( .A1(n4), .A2(n19), .ZN(n219) );
  NAND2_X1 U180 ( .A1(n4), .A2(n18), .ZN(n220) );
  NAND2_X1 U181 ( .A1(n19), .A2(n18), .ZN(n221) );
  NAND3_X1 U182 ( .A1(n219), .A2(n220), .A3(n221), .ZN(n3) );
  XNOR2_X1 U183 ( .A(n2), .B(n208), .ZN(product[14]) );
  XOR2_X1 U184 ( .A(n17), .B(n280), .Z(n222) );
  XOR2_X1 U185 ( .A(n3), .B(n222), .Z(product[13]) );
  NAND2_X1 U186 ( .A1(n3), .A2(n17), .ZN(n223) );
  NAND2_X1 U187 ( .A1(n3), .A2(n280), .ZN(n224) );
  NAND2_X1 U188 ( .A1(n17), .A2(n280), .ZN(n225) );
  NAND3_X1 U189 ( .A1(n223), .A2(n224), .A3(n225), .ZN(n2) );
  NAND3_X1 U190 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n226) );
  NAND3_X1 U191 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n227) );
  NAND3_X1 U192 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n228) );
  NAND3_X1 U193 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n229) );
  CLKBUF_X1 U194 ( .A(b[3]), .Z(n230) );
  XOR2_X1 U195 ( .A(n27), .B(n24), .Z(n231) );
  XOR2_X1 U196 ( .A(n6), .B(n231), .Z(product[10]) );
  NAND2_X1 U197 ( .A1(n6), .A2(n27), .ZN(n232) );
  NAND2_X1 U198 ( .A1(n6), .A2(n24), .ZN(n233) );
  NAND2_X1 U199 ( .A1(n27), .A2(n24), .ZN(n234) );
  NAND3_X1 U200 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n5) );
  OAI22_X1 U201 ( .A1(n253), .A2(n292), .B1(n338), .B2(n290), .ZN(n235) );
  XOR2_X1 U202 ( .A(n23), .B(n20), .Z(n236) );
  XOR2_X1 U203 ( .A(n227), .B(n236), .Z(product[11]) );
  NAND2_X1 U204 ( .A1(n226), .A2(n23), .ZN(n237) );
  NAND2_X1 U205 ( .A1(n5), .A2(n20), .ZN(n238) );
  NAND2_X1 U206 ( .A1(n23), .A2(n20), .ZN(n239) );
  NAND3_X1 U207 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n4) );
  CLKBUF_X1 U208 ( .A(b[4]), .Z(n240) );
  XOR2_X1 U209 ( .A(n95), .B(n102), .Z(n241) );
  XOR2_X1 U210 ( .A(n46), .B(n49), .Z(n242) );
  XOR2_X1 U211 ( .A(n242), .B(n10), .Z(product[6]) );
  NAND2_X1 U212 ( .A1(n46), .A2(n49), .ZN(n243) );
  NAND2_X1 U213 ( .A1(n46), .A2(n10), .ZN(n244) );
  NAND2_X1 U214 ( .A1(n49), .A2(n10), .ZN(n245) );
  NAND3_X1 U215 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n9) );
  XOR2_X1 U216 ( .A(n40), .B(n45), .Z(n246) );
  XOR2_X1 U217 ( .A(n246), .B(n229), .Z(product[7]) );
  NAND2_X1 U218 ( .A1(n40), .A2(n45), .ZN(n247) );
  NAND2_X1 U219 ( .A1(n40), .A2(n228), .ZN(n248) );
  NAND2_X1 U220 ( .A1(n45), .A2(n9), .ZN(n249) );
  NAND3_X1 U221 ( .A1(n247), .A2(n248), .A3(n249), .ZN(n8) );
  NAND2_X1 U222 ( .A1(n2), .A2(n281), .ZN(n250) );
  NAND2_X1 U223 ( .A1(n2), .A2(n15), .ZN(n251) );
  NAND2_X1 U224 ( .A1(n281), .A2(n15), .ZN(n252) );
  BUF_X1 U225 ( .A(n337), .Z(n253) );
  NAND3_X1 U226 ( .A1(n265), .A2(n264), .A3(n263), .ZN(n254) );
  NAND3_X1 U227 ( .A1(n263), .A2(n212), .A3(n265), .ZN(n255) );
  CLKBUF_X1 U228 ( .A(n13), .Z(n256) );
  NAND2_X1 U229 ( .A1(a[4]), .A2(a[3]), .ZN(n259) );
  NAND2_X1 U230 ( .A1(n257), .A2(n258), .ZN(n260) );
  INV_X1 U231 ( .A(a[4]), .ZN(n257) );
  INV_X1 U232 ( .A(a[3]), .ZN(n258) );
  XNOR2_X1 U233 ( .A(n14), .B(n261), .ZN(product[2]) );
  XNOR2_X1 U234 ( .A(n103), .B(n96), .ZN(n261) );
  XNOR2_X1 U235 ( .A(n262), .B(n256), .ZN(product[3]) );
  XNOR2_X1 U236 ( .A(n241), .B(n71), .ZN(n262) );
  NAND2_X1 U237 ( .A1(n56), .A2(n71), .ZN(n263) );
  NAND2_X1 U238 ( .A1(n13), .A2(n241), .ZN(n264) );
  NAND2_X1 U239 ( .A1(n71), .A2(n13), .ZN(n265) );
  NAND3_X1 U240 ( .A1(n263), .A2(n264), .A3(n265), .ZN(n12) );
  XOR2_X1 U241 ( .A(n54), .B(n207), .Z(n266) );
  XOR2_X1 U242 ( .A(n266), .B(n255), .Z(product[4]) );
  NAND2_X1 U243 ( .A1(n54), .A2(n207), .ZN(n267) );
  NAND2_X1 U244 ( .A1(n54), .A2(n254), .ZN(n268) );
  NAND2_X1 U245 ( .A1(n207), .A2(n12), .ZN(n269) );
  NAND3_X1 U246 ( .A1(n267), .A2(n268), .A3(n269), .ZN(n11) );
  NAND2_X1 U247 ( .A1(n14), .A2(n235), .ZN(n270) );
  NAND2_X1 U248 ( .A1(n14), .A2(n96), .ZN(n271) );
  NAND2_X1 U249 ( .A1(n235), .A2(n96), .ZN(n272) );
  NAND3_X1 U250 ( .A1(n270), .A2(n271), .A3(n272), .ZN(n13) );
  XOR2_X1 U251 ( .A(n211), .B(n102), .Z(n56) );
  INV_X1 U252 ( .A(n279), .ZN(n273) );
  BUF_X2 U253 ( .A(n296), .Z(n274) );
  INV_X1 U254 ( .A(n21), .ZN(n283) );
  INV_X1 U255 ( .A(n315), .ZN(n284) );
  INV_X1 U256 ( .A(n326), .ZN(n281) );
  INV_X1 U257 ( .A(n295), .ZN(n288) );
  INV_X1 U258 ( .A(n304), .ZN(n287) );
  INV_X1 U259 ( .A(n31), .ZN(n286) );
  INV_X1 U260 ( .A(b[0]), .ZN(n279) );
  INV_X1 U261 ( .A(a[5]), .ZN(n285) );
  INV_X1 U262 ( .A(a[7]), .ZN(n282) );
  INV_X1 U263 ( .A(a[1]), .ZN(n276) );
  INV_X2 U264 ( .A(n276), .ZN(n277) );
  INV_X1 U265 ( .A(a[1]), .ZN(n289) );
  XOR2_X2 U266 ( .A(a[6]), .B(n285), .Z(n317) );
  INV_X1 U267 ( .A(n279), .ZN(n278) );
  INV_X2 U268 ( .A(a[0]), .ZN(n290) );
  NOR2_X1 U269 ( .A1(n290), .A2(n279), .ZN(product[0]) );
  OAI22_X1 U270 ( .A1(n291), .A2(n292), .B1(n293), .B2(n290), .ZN(n99) );
  OAI22_X1 U271 ( .A1(n293), .A2(n292), .B1(n294), .B2(n290), .ZN(n98) );
  XNOR2_X1 U272 ( .A(b[6]), .B(n277), .ZN(n293) );
  OAI22_X1 U273 ( .A1(n290), .A2(n294), .B1(n292), .B2(n294), .ZN(n295) );
  XNOR2_X1 U274 ( .A(b[7]), .B(n277), .ZN(n294) );
  NOR2_X1 U275 ( .A1(n296), .A2(n279), .ZN(n96) );
  OAI22_X1 U276 ( .A1(n297), .A2(n298), .B1(n296), .B2(n299), .ZN(n95) );
  XNOR2_X1 U277 ( .A(a[3]), .B(n278), .ZN(n297) );
  OAI22_X1 U278 ( .A1(n299), .A2(n298), .B1(n274), .B2(n300), .ZN(n94) );
  XNOR2_X1 U279 ( .A(n275), .B(a[3]), .ZN(n299) );
  OAI22_X1 U280 ( .A1(n300), .A2(n213), .B1(n274), .B2(n301), .ZN(n93) );
  XNOR2_X1 U281 ( .A(b[2]), .B(a[3]), .ZN(n300) );
  OAI22_X1 U282 ( .A1(n301), .A2(n213), .B1(n274), .B2(n302), .ZN(n92) );
  XNOR2_X1 U283 ( .A(n230), .B(a[3]), .ZN(n301) );
  OAI22_X1 U284 ( .A1(n302), .A2(n213), .B1(n274), .B2(n303), .ZN(n91) );
  XNOR2_X1 U285 ( .A(b[4]), .B(a[3]), .ZN(n302) );
  OAI22_X1 U286 ( .A1(n305), .A2(n274), .B1(n213), .B2(n305), .ZN(n304) );
  NOR2_X1 U287 ( .A1(n210), .A2(n279), .ZN(n88) );
  OAI22_X1 U288 ( .A1(n307), .A2(n308), .B1(n210), .B2(n309), .ZN(n87) );
  XNOR2_X1 U289 ( .A(a[5]), .B(n278), .ZN(n307) );
  OAI22_X1 U290 ( .A1(n309), .A2(n206), .B1(n210), .B2(n310), .ZN(n86) );
  XNOR2_X1 U291 ( .A(n275), .B(a[5]), .ZN(n309) );
  OAI22_X1 U292 ( .A1(n310), .A2(n206), .B1(n210), .B2(n311), .ZN(n85) );
  XNOR2_X1 U293 ( .A(b[2]), .B(a[5]), .ZN(n310) );
  OAI22_X1 U294 ( .A1(n311), .A2(n206), .B1(n210), .B2(n312), .ZN(n84) );
  XNOR2_X1 U295 ( .A(n230), .B(a[5]), .ZN(n311) );
  OAI22_X1 U296 ( .A1(n312), .A2(n206), .B1(n210), .B2(n313), .ZN(n83) );
  XNOR2_X1 U297 ( .A(n240), .B(a[5]), .ZN(n312) );
  OAI22_X1 U298 ( .A1(n313), .A2(n206), .B1(n210), .B2(n314), .ZN(n82) );
  XNOR2_X1 U299 ( .A(b[5]), .B(a[5]), .ZN(n313) );
  OAI22_X1 U300 ( .A1(n316), .A2(n210), .B1(n206), .B2(n316), .ZN(n315) );
  NOR2_X1 U301 ( .A1(n317), .A2(n279), .ZN(n80) );
  OAI22_X1 U302 ( .A1(n318), .A2(n319), .B1(n317), .B2(n320), .ZN(n79) );
  XNOR2_X1 U303 ( .A(a[7]), .B(n273), .ZN(n318) );
  OAI22_X1 U304 ( .A1(n321), .A2(n319), .B1(n317), .B2(n322), .ZN(n77) );
  OAI22_X1 U305 ( .A1(n322), .A2(n319), .B1(n317), .B2(n323), .ZN(n76) );
  XNOR2_X1 U306 ( .A(n230), .B(a[7]), .ZN(n322) );
  OAI22_X1 U307 ( .A1(n323), .A2(n319), .B1(n317), .B2(n324), .ZN(n75) );
  XNOR2_X1 U308 ( .A(n240), .B(a[7]), .ZN(n323) );
  OAI22_X1 U309 ( .A1(n324), .A2(n319), .B1(n317), .B2(n325), .ZN(n74) );
  XNOR2_X1 U310 ( .A(b[5]), .B(a[7]), .ZN(n324) );
  OAI22_X1 U311 ( .A1(n327), .A2(n317), .B1(n319), .B2(n327), .ZN(n326) );
  OAI21_X1 U312 ( .B1(n273), .B2(n289), .A(n292), .ZN(n72) );
  OAI21_X1 U313 ( .B1(n258), .B2(n213), .A(n328), .ZN(n71) );
  OR3_X1 U314 ( .A1(n274), .A2(n273), .A3(n258), .ZN(n328) );
  OAI21_X1 U315 ( .B1(n285), .B2(n308), .A(n329), .ZN(n70) );
  OR3_X1 U316 ( .A1(n306), .A2(n273), .A3(n285), .ZN(n329) );
  OAI21_X1 U317 ( .B1(n282), .B2(n319), .A(n330), .ZN(n69) );
  OR3_X1 U318 ( .A1(n317), .A2(n278), .A3(n282), .ZN(n330) );
  XNOR2_X1 U319 ( .A(n331), .B(n332), .ZN(n38) );
  OR2_X1 U320 ( .A1(n331), .A2(n332), .ZN(n37) );
  OAI22_X1 U321 ( .A1(n303), .A2(n213), .B1(n274), .B2(n333), .ZN(n332) );
  XNOR2_X1 U322 ( .A(b[5]), .B(a[3]), .ZN(n303) );
  OAI22_X1 U323 ( .A1(n320), .A2(n319), .B1(n317), .B2(n321), .ZN(n331) );
  XNOR2_X1 U324 ( .A(b[2]), .B(a[7]), .ZN(n321) );
  XNOR2_X1 U325 ( .A(n275), .B(a[7]), .ZN(n320) );
  OAI22_X1 U326 ( .A1(n333), .A2(n213), .B1(n274), .B2(n305), .ZN(n31) );
  XNOR2_X1 U327 ( .A(b[7]), .B(a[3]), .ZN(n305) );
  XNOR2_X1 U328 ( .A(n258), .B(a[2]), .ZN(n334) );
  XNOR2_X1 U329 ( .A(b[6]), .B(a[3]), .ZN(n333) );
  OAI22_X1 U330 ( .A1(n314), .A2(n206), .B1(n210), .B2(n316), .ZN(n21) );
  XNOR2_X1 U331 ( .A(b[7]), .B(a[5]), .ZN(n316) );
  XNOR2_X1 U332 ( .A(n285), .B(a[4]), .ZN(n335) );
  XNOR2_X1 U333 ( .A(b[6]), .B(a[5]), .ZN(n314) );
  OAI22_X1 U334 ( .A1(n325), .A2(n319), .B1(n317), .B2(n327), .ZN(n15) );
  XNOR2_X1 U335 ( .A(b[7]), .B(a[7]), .ZN(n327) );
  NAND2_X1 U336 ( .A1(n317), .A2(n336), .ZN(n319) );
  XNOR2_X1 U337 ( .A(n282), .B(a[6]), .ZN(n336) );
  XNOR2_X1 U338 ( .A(b[6]), .B(a[7]), .ZN(n325) );
  OAI22_X1 U339 ( .A1(n278), .A2(n292), .B1(n337), .B2(n290), .ZN(n104) );
  OAI22_X1 U340 ( .A1(n253), .A2(n292), .B1(n338), .B2(n290), .ZN(n103) );
  XNOR2_X1 U341 ( .A(b[1]), .B(n277), .ZN(n337) );
  OAI22_X1 U342 ( .A1(n338), .A2(n292), .B1(n339), .B2(n290), .ZN(n102) );
  XNOR2_X1 U343 ( .A(b[2]), .B(n277), .ZN(n338) );
  OAI22_X1 U344 ( .A1(n339), .A2(n292), .B1(n340), .B2(n290), .ZN(n101) );
  XNOR2_X1 U345 ( .A(b[3]), .B(n277), .ZN(n339) );
  OAI22_X1 U346 ( .A1(n340), .A2(n292), .B1(n291), .B2(n290), .ZN(n100) );
  XNOR2_X1 U347 ( .A(b[5]), .B(n277), .ZN(n291) );
  NAND2_X1 U348 ( .A1(a[1]), .A2(n290), .ZN(n292) );
  XNOR2_X1 U349 ( .A(b[4]), .B(n277), .ZN(n340) );
endmodule


module datapath_DW01_add_8 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n65;
  wire   [15:1] carry;

  FA_X1 U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n65), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[14]), .ZN(n8) );
  NAND3_X1 U2 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n1) );
  NAND3_X1 U3 ( .A1(n21), .A2(n22), .A3(n23), .ZN(n2) );
  NAND2_X1 U4 ( .A1(n46), .A2(B[8]), .ZN(n3) );
  XOR2_X1 U5 ( .A(n2), .B(A[5]), .Z(n4) );
  XOR2_X1 U6 ( .A(B[5]), .B(n4), .Z(SUM[5]) );
  NAND2_X1 U7 ( .A1(B[5]), .A2(n1), .ZN(n5) );
  NAND2_X1 U8 ( .A1(B[5]), .A2(A[5]), .ZN(n6) );
  NAND2_X1 U9 ( .A1(carry[5]), .A2(A[5]), .ZN(n7) );
  NAND3_X1 U10 ( .A1(n5), .A2(n6), .A3(n7), .ZN(carry[6]) );
  XNOR2_X1 U11 ( .A(B[14]), .B(n8), .ZN(n9) );
  XOR2_X1 U12 ( .A(n14), .B(n9), .Z(SUM[14]) );
  NAND2_X1 U13 ( .A1(n13), .A2(B[14]), .ZN(n10) );
  NAND2_X1 U14 ( .A1(carry[14]), .A2(A[14]), .ZN(n11) );
  NAND2_X1 U15 ( .A1(B[14]), .A2(A[14]), .ZN(n12) );
  NAND3_X1 U16 ( .A1(n10), .A2(n11), .A3(n12), .ZN(carry[15]) );
  NAND3_X1 U17 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n13) );
  NAND3_X1 U18 ( .A1(n52), .A2(n53), .A3(n54), .ZN(n14) );
  NAND3_X1 U19 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n15) );
  XOR2_X1 U20 ( .A(carry[3]), .B(A[3]), .Z(n16) );
  XOR2_X1 U21 ( .A(B[3]), .B(n16), .Z(SUM[3]) );
  NAND2_X1 U22 ( .A1(carry[3]), .A2(B[3]), .ZN(n17) );
  NAND2_X1 U23 ( .A1(B[3]), .A2(A[3]), .ZN(n18) );
  NAND2_X1 U24 ( .A1(carry[3]), .A2(A[3]), .ZN(n19) );
  NAND3_X1 U25 ( .A1(n17), .A2(n18), .A3(n19), .ZN(carry[4]) );
  XOR2_X1 U26 ( .A(B[4]), .B(A[4]), .Z(n20) );
  XOR2_X1 U27 ( .A(carry[4]), .B(n20), .Z(SUM[4]) );
  NAND2_X1 U28 ( .A1(carry[4]), .A2(B[4]), .ZN(n21) );
  NAND2_X1 U29 ( .A1(carry[4]), .A2(A[4]), .ZN(n22) );
  NAND2_X1 U30 ( .A1(B[4]), .A2(A[4]), .ZN(n23) );
  NAND3_X1 U31 ( .A1(n21), .A2(n22), .A3(n23), .ZN(carry[5]) );
  NAND3_X1 U32 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n24) );
  NAND3_X1 U33 ( .A1(n3), .A2(n49), .A3(n50), .ZN(n25) );
  NAND3_X1 U34 ( .A1(n3), .A2(n49), .A3(n50), .ZN(n26) );
  XOR2_X1 U35 ( .A(B[9]), .B(A[9]), .Z(n27) );
  XOR2_X1 U36 ( .A(n26), .B(n27), .Z(SUM[9]) );
  NAND2_X1 U37 ( .A1(n25), .A2(B[9]), .ZN(n28) );
  NAND2_X1 U38 ( .A1(carry[9]), .A2(A[9]), .ZN(n29) );
  NAND2_X1 U39 ( .A1(B[9]), .A2(A[9]), .ZN(n30) );
  NAND3_X1 U40 ( .A1(n28), .A2(n29), .A3(n30), .ZN(carry[10]) );
  NAND3_X1 U41 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n31) );
  NAND3_X1 U42 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n32) );
  XOR2_X1 U43 ( .A(B[10]), .B(A[10]), .Z(n33) );
  XOR2_X1 U44 ( .A(n15), .B(n33), .Z(SUM[10]) );
  NAND2_X1 U45 ( .A1(n15), .A2(B[10]), .ZN(n34) );
  NAND2_X1 U46 ( .A1(carry[10]), .A2(A[10]), .ZN(n35) );
  NAND2_X1 U47 ( .A1(B[10]), .A2(A[10]), .ZN(n36) );
  NAND3_X1 U48 ( .A1(n35), .A2(n34), .A3(n36), .ZN(carry[11]) );
  XOR2_X1 U49 ( .A(B[12]), .B(A[12]), .Z(n37) );
  XOR2_X1 U50 ( .A(carry[12]), .B(n37), .Z(SUM[12]) );
  NAND2_X1 U51 ( .A1(n31), .A2(B[12]), .ZN(n38) );
  NAND2_X1 U52 ( .A1(carry[12]), .A2(A[12]), .ZN(n39) );
  NAND2_X1 U53 ( .A1(B[12]), .A2(A[12]), .ZN(n40) );
  NAND3_X1 U54 ( .A1(n38), .A2(n39), .A3(n40), .ZN(carry[13]) );
  NAND3_X1 U55 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n41) );
  XOR2_X1 U56 ( .A(B[11]), .B(A[11]), .Z(n42) );
  XOR2_X1 U57 ( .A(n24), .B(n42), .Z(SUM[11]) );
  NAND2_X1 U58 ( .A1(n24), .A2(B[11]), .ZN(n43) );
  NAND2_X1 U59 ( .A1(carry[11]), .A2(A[11]), .ZN(n44) );
  NAND2_X1 U60 ( .A1(B[11]), .A2(A[11]), .ZN(n45) );
  NAND3_X1 U61 ( .A1(n43), .A2(n44), .A3(n45), .ZN(carry[12]) );
  NAND3_X1 U62 ( .A1(n60), .A2(n61), .A3(n62), .ZN(n46) );
  XOR2_X1 U63 ( .A(B[8]), .B(A[8]), .Z(n47) );
  XOR2_X1 U64 ( .A(n46), .B(n47), .Z(SUM[8]) );
  NAND2_X1 U65 ( .A1(n46), .A2(B[8]), .ZN(n48) );
  NAND2_X1 U66 ( .A1(carry[8]), .A2(A[8]), .ZN(n49) );
  NAND2_X1 U67 ( .A1(B[8]), .A2(A[8]), .ZN(n50) );
  NAND3_X1 U68 ( .A1(n48), .A2(n49), .A3(n50), .ZN(carry[9]) );
  XOR2_X1 U69 ( .A(B[13]), .B(A[13]), .Z(n51) );
  XOR2_X1 U70 ( .A(carry[13]), .B(n51), .Z(SUM[13]) );
  NAND2_X1 U71 ( .A1(B[13]), .A2(carry[13]), .ZN(n52) );
  NAND2_X1 U72 ( .A1(n32), .A2(A[13]), .ZN(n53) );
  NAND2_X1 U73 ( .A1(B[13]), .A2(A[13]), .ZN(n54) );
  NAND3_X1 U74 ( .A1(n52), .A2(n53), .A3(n54), .ZN(carry[14]) );
  XOR2_X1 U75 ( .A(B[6]), .B(A[6]), .Z(n55) );
  XOR2_X1 U76 ( .A(carry[6]), .B(n55), .Z(SUM[6]) );
  NAND2_X1 U77 ( .A1(carry[6]), .A2(B[6]), .ZN(n56) );
  NAND2_X1 U78 ( .A1(carry[6]), .A2(A[6]), .ZN(n57) );
  NAND2_X1 U79 ( .A1(B[6]), .A2(A[6]), .ZN(n58) );
  NAND3_X1 U80 ( .A1(n56), .A2(n57), .A3(n58), .ZN(carry[7]) );
  XOR2_X1 U81 ( .A(B[7]), .B(A[7]), .Z(n59) );
  XOR2_X1 U82 ( .A(carry[7]), .B(n59), .Z(SUM[7]) );
  NAND2_X1 U83 ( .A1(n41), .A2(B[7]), .ZN(n60) );
  NAND2_X1 U84 ( .A1(n41), .A2(A[7]), .ZN(n61) );
  NAND2_X1 U85 ( .A1(B[7]), .A2(A[7]), .ZN(n62) );
  NAND3_X1 U86 ( .A1(n60), .A2(n61), .A3(n62), .ZN(carry[8]) );
  XNOR2_X1 U87 ( .A(carry[15]), .B(n63), .ZN(SUM[15]) );
  XNOR2_X1 U88 ( .A(B[15]), .B(A[15]), .ZN(n63) );
  XOR2_X1 U89 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U90 ( .A1(B[0]), .A2(A[0]), .ZN(n65) );
endmodule


module datapath_DW_mult_tc_7 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74,
         n75, n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92,
         n93, n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330;

  FA_X1 U10 ( .A(n46), .B(n49), .CI(n10), .CO(n9), .S(product[6]) );
  FA_X1 U13 ( .A(n13), .B(n71), .CI(n56), .CO(n12), .S(product[3]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n273), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n272), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n276), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n275), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n278), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  NAND2_X1 U157 ( .A1(n19), .A2(n18), .ZN(n216) );
  NAND2_X2 U158 ( .A1(n286), .A2(n324), .ZN(n288) );
  XNOR2_X1 U159 ( .A(n270), .B(n15), .ZN(n206) );
  AND3_X1 U160 ( .A1(n256), .A2(n257), .A3(n258), .ZN(product[15]) );
  NAND3_X1 U161 ( .A1(n238), .A2(n237), .A3(n239), .ZN(n208) );
  NAND3_X1 U162 ( .A1(n238), .A2(n237), .A3(n239), .ZN(n209) );
  NAND3_X1 U163 ( .A1(n216), .A2(n217), .A3(n218), .ZN(n210) );
  NAND3_X1 U164 ( .A1(n216), .A2(n217), .A3(n218), .ZN(n211) );
  INV_X1 U165 ( .A(n268), .ZN(n212) );
  XOR2_X2 U166 ( .A(a[6]), .B(n274), .Z(n307) );
  XNOR2_X1 U167 ( .A(n2), .B(n206), .ZN(product[14]) );
  XNOR2_X1 U168 ( .A(n213), .B(n11), .ZN(product[5]) );
  XNOR2_X1 U169 ( .A(n50), .B(n53), .ZN(n213) );
  XNOR2_X1 U170 ( .A(n214), .B(n12), .ZN(product[4]) );
  XNOR2_X1 U171 ( .A(n54), .B(n55), .ZN(n214) );
  XOR2_X1 U172 ( .A(a[3]), .B(n268), .Z(n287) );
  INV_X1 U173 ( .A(n268), .ZN(n267) );
  XOR2_X1 U174 ( .A(n19), .B(n18), .Z(n215) );
  XOR2_X1 U175 ( .A(n215), .B(n209), .Z(product[12]) );
  NAND2_X1 U176 ( .A1(n19), .A2(n208), .ZN(n217) );
  NAND2_X1 U177 ( .A1(n18), .A2(n4), .ZN(n218) );
  NAND3_X1 U178 ( .A1(n216), .A2(n217), .A3(n218), .ZN(n3) );
  XOR2_X1 U179 ( .A(n17), .B(n269), .Z(n219) );
  XOR2_X1 U180 ( .A(n219), .B(n211), .Z(product[13]) );
  NAND2_X1 U181 ( .A1(n17), .A2(n269), .ZN(n220) );
  NAND2_X1 U182 ( .A1(n17), .A2(n210), .ZN(n221) );
  NAND2_X1 U183 ( .A1(n269), .A2(n3), .ZN(n222) );
  NAND3_X1 U184 ( .A1(n220), .A2(n221), .A3(n222), .ZN(n2) );
  NAND3_X1 U185 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n223) );
  NAND3_X1 U186 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n224) );
  NAND3_X1 U187 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n225) );
  NAND3_X1 U188 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n226) );
  XOR2_X1 U189 ( .A(n40), .B(n45), .Z(n227) );
  XOR2_X1 U190 ( .A(n227), .B(n9), .Z(product[7]) );
  NAND2_X1 U191 ( .A1(n40), .A2(n45), .ZN(n228) );
  NAND2_X1 U192 ( .A1(n40), .A2(n9), .ZN(n229) );
  NAND2_X1 U193 ( .A1(n45), .A2(n9), .ZN(n230) );
  NAND3_X1 U194 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n8) );
  XOR2_X1 U195 ( .A(n34), .B(n39), .Z(n231) );
  XOR2_X1 U196 ( .A(n231), .B(n226), .Z(product[8]) );
  NAND2_X1 U197 ( .A1(n34), .A2(n39), .ZN(n232) );
  NAND2_X1 U198 ( .A1(n34), .A2(n225), .ZN(n233) );
  NAND2_X1 U199 ( .A1(n39), .A2(n8), .ZN(n234) );
  NAND3_X1 U200 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n7) );
  NAND3_X1 U201 ( .A1(n246), .A2(n247), .A3(n248), .ZN(n235) );
  XOR2_X1 U202 ( .A(n23), .B(n20), .Z(n236) );
  XOR2_X1 U203 ( .A(n235), .B(n236), .Z(product[11]) );
  NAND2_X1 U204 ( .A1(n5), .A2(n23), .ZN(n237) );
  NAND2_X1 U205 ( .A1(n5), .A2(n20), .ZN(n238) );
  NAND2_X1 U206 ( .A1(n23), .A2(n20), .ZN(n239) );
  NAND3_X1 U207 ( .A1(n238), .A2(n237), .A3(n239), .ZN(n4) );
  XOR2_X1 U208 ( .A(n33), .B(n28), .Z(n240) );
  XOR2_X1 U209 ( .A(n224), .B(n240), .Z(product[9]) );
  NAND2_X1 U210 ( .A1(n223), .A2(n33), .ZN(n241) );
  NAND2_X1 U211 ( .A1(n7), .A2(n28), .ZN(n242) );
  NAND2_X1 U212 ( .A1(n33), .A2(n28), .ZN(n243) );
  NAND3_X1 U213 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n6) );
  NAND3_X1 U214 ( .A1(n250), .A2(n249), .A3(n251), .ZN(n244) );
  XOR2_X1 U215 ( .A(n27), .B(n24), .Z(n245) );
  XOR2_X1 U216 ( .A(n6), .B(n245), .Z(product[10]) );
  NAND2_X1 U217 ( .A1(n6), .A2(n27), .ZN(n246) );
  NAND2_X1 U218 ( .A1(n6), .A2(n24), .ZN(n247) );
  NAND2_X1 U219 ( .A1(n27), .A2(n24), .ZN(n248) );
  NAND3_X1 U220 ( .A1(n247), .A2(n246), .A3(n248), .ZN(n5) );
  NAND2_X1 U221 ( .A1(n54), .A2(n55), .ZN(n249) );
  NAND2_X1 U222 ( .A1(n12), .A2(n54), .ZN(n250) );
  NAND2_X1 U223 ( .A1(n55), .A2(n12), .ZN(n251) );
  NAND3_X1 U224 ( .A1(n251), .A2(n250), .A3(n249), .ZN(n11) );
  NAND2_X1 U225 ( .A1(n50), .A2(n53), .ZN(n252) );
  NAND2_X1 U226 ( .A1(n50), .A2(n244), .ZN(n253) );
  NAND2_X1 U227 ( .A1(n53), .A2(n11), .ZN(n254) );
  NAND3_X1 U228 ( .A1(n254), .A2(n253), .A3(n252), .ZN(n10) );
  CLKBUF_X1 U229 ( .A(n14), .Z(n255) );
  NAND2_X1 U230 ( .A1(n2), .A2(n270), .ZN(n256) );
  NAND2_X1 U231 ( .A1(n2), .A2(n15), .ZN(n257) );
  NAND2_X1 U232 ( .A1(n270), .A2(n15), .ZN(n258) );
  NAND2_X1 U233 ( .A1(a[4]), .A2(a[3]), .ZN(n260) );
  NAND2_X1 U234 ( .A1(n259), .A2(n277), .ZN(n261) );
  NAND2_X2 U235 ( .A1(n260), .A2(n261), .ZN(n296) );
  INV_X1 U236 ( .A(a[4]), .ZN(n259) );
  NAND2_X2 U237 ( .A1(n296), .A2(n325), .ZN(n298) );
  XNOR2_X1 U238 ( .A(a[2]), .B(a[1]), .ZN(n262) );
  INV_X1 U239 ( .A(n15), .ZN(n269) );
  INV_X1 U240 ( .A(n21), .ZN(n272) );
  INV_X1 U241 ( .A(n305), .ZN(n273) );
  INV_X1 U242 ( .A(n316), .ZN(n270) );
  INV_X1 U243 ( .A(n285), .ZN(n278) );
  INV_X1 U244 ( .A(n294), .ZN(n276) );
  INV_X1 U245 ( .A(n31), .ZN(n275) );
  INV_X1 U246 ( .A(b[0]), .ZN(n268) );
  XNOR2_X1 U247 ( .A(a[2]), .B(a[1]), .ZN(n286) );
  INV_X1 U248 ( .A(a[0]), .ZN(n280) );
  INV_X1 U249 ( .A(a[5]), .ZN(n274) );
  INV_X1 U250 ( .A(a[7]), .ZN(n271) );
  XNOR2_X1 U251 ( .A(n255), .B(n263), .ZN(product[2]) );
  XNOR2_X1 U252 ( .A(n103), .B(n96), .ZN(n263) );
  NAND2_X1 U253 ( .A1(n14), .A2(n103), .ZN(n264) );
  NAND2_X1 U254 ( .A1(n14), .A2(n96), .ZN(n265) );
  NAND2_X1 U255 ( .A1(n103), .A2(n96), .ZN(n266) );
  NAND3_X1 U256 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n13) );
  INV_X1 U257 ( .A(a[3]), .ZN(n277) );
  INV_X1 U258 ( .A(a[1]), .ZN(n279) );
  NOR2_X1 U259 ( .A1(n280), .A2(n268), .ZN(product[0]) );
  OAI22_X1 U260 ( .A1(n281), .A2(n282), .B1(n283), .B2(n280), .ZN(n99) );
  OAI22_X1 U261 ( .A1(n283), .A2(n282), .B1(n284), .B2(n280), .ZN(n98) );
  XNOR2_X1 U262 ( .A(b[6]), .B(a[1]), .ZN(n283) );
  OAI22_X1 U263 ( .A1(n280), .A2(n284), .B1(n282), .B2(n284), .ZN(n285) );
  XNOR2_X1 U264 ( .A(b[7]), .B(a[1]), .ZN(n284) );
  NOR2_X1 U265 ( .A1(n262), .A2(n268), .ZN(n96) );
  OAI22_X1 U266 ( .A1(n287), .A2(n288), .B1(n262), .B2(n289), .ZN(n95) );
  OAI22_X1 U267 ( .A1(n289), .A2(n288), .B1(n262), .B2(n290), .ZN(n94) );
  XNOR2_X1 U268 ( .A(b[1]), .B(a[3]), .ZN(n289) );
  OAI22_X1 U269 ( .A1(n290), .A2(n288), .B1(n262), .B2(n291), .ZN(n93) );
  XNOR2_X1 U270 ( .A(b[2]), .B(a[3]), .ZN(n290) );
  OAI22_X1 U271 ( .A1(n291), .A2(n288), .B1(n262), .B2(n292), .ZN(n92) );
  XNOR2_X1 U272 ( .A(b[3]), .B(a[3]), .ZN(n291) );
  OAI22_X1 U273 ( .A1(n292), .A2(n288), .B1(n262), .B2(n293), .ZN(n91) );
  XNOR2_X1 U274 ( .A(b[4]), .B(a[3]), .ZN(n292) );
  OAI22_X1 U275 ( .A1(n295), .A2(n262), .B1(n288), .B2(n295), .ZN(n294) );
  NOR2_X1 U276 ( .A1(n296), .A2(n268), .ZN(n88) );
  OAI22_X1 U277 ( .A1(n297), .A2(n298), .B1(n296), .B2(n299), .ZN(n87) );
  XNOR2_X1 U278 ( .A(a[5]), .B(n212), .ZN(n297) );
  OAI22_X1 U279 ( .A1(n299), .A2(n298), .B1(n296), .B2(n300), .ZN(n86) );
  XNOR2_X1 U280 ( .A(b[1]), .B(a[5]), .ZN(n299) );
  OAI22_X1 U281 ( .A1(n300), .A2(n298), .B1(n296), .B2(n301), .ZN(n85) );
  XNOR2_X1 U282 ( .A(b[2]), .B(a[5]), .ZN(n300) );
  OAI22_X1 U283 ( .A1(n301), .A2(n298), .B1(n296), .B2(n302), .ZN(n84) );
  XNOR2_X1 U284 ( .A(b[3]), .B(a[5]), .ZN(n301) );
  OAI22_X1 U285 ( .A1(n302), .A2(n298), .B1(n296), .B2(n303), .ZN(n83) );
  XNOR2_X1 U286 ( .A(b[4]), .B(a[5]), .ZN(n302) );
  OAI22_X1 U287 ( .A1(n303), .A2(n298), .B1(n296), .B2(n304), .ZN(n82) );
  XNOR2_X1 U288 ( .A(b[5]), .B(a[5]), .ZN(n303) );
  OAI22_X1 U289 ( .A1(n306), .A2(n296), .B1(n298), .B2(n306), .ZN(n305) );
  NOR2_X1 U290 ( .A1(n307), .A2(n268), .ZN(n80) );
  OAI22_X1 U291 ( .A1(n308), .A2(n309), .B1(n307), .B2(n310), .ZN(n79) );
  XNOR2_X1 U292 ( .A(a[7]), .B(n212), .ZN(n308) );
  OAI22_X1 U293 ( .A1(n311), .A2(n309), .B1(n307), .B2(n312), .ZN(n77) );
  OAI22_X1 U294 ( .A1(n312), .A2(n309), .B1(n307), .B2(n313), .ZN(n76) );
  XNOR2_X1 U295 ( .A(b[3]), .B(a[7]), .ZN(n312) );
  OAI22_X1 U296 ( .A1(n313), .A2(n309), .B1(n307), .B2(n314), .ZN(n75) );
  XNOR2_X1 U297 ( .A(b[4]), .B(a[7]), .ZN(n313) );
  OAI22_X1 U298 ( .A1(n314), .A2(n309), .B1(n307), .B2(n315), .ZN(n74) );
  XNOR2_X1 U299 ( .A(b[5]), .B(a[7]), .ZN(n314) );
  OAI22_X1 U300 ( .A1(n317), .A2(n307), .B1(n309), .B2(n317), .ZN(n316) );
  OAI21_X1 U301 ( .B1(n267), .B2(n279), .A(n282), .ZN(n72) );
  OAI21_X1 U302 ( .B1(n277), .B2(n288), .A(n318), .ZN(n71) );
  OR3_X1 U303 ( .A1(n262), .A2(n212), .A3(n277), .ZN(n318) );
  OAI21_X1 U304 ( .B1(n274), .B2(n298), .A(n319), .ZN(n70) );
  OR3_X1 U305 ( .A1(n296), .A2(n267), .A3(n274), .ZN(n319) );
  OAI21_X1 U306 ( .B1(n271), .B2(n309), .A(n320), .ZN(n69) );
  OR3_X1 U307 ( .A1(n307), .A2(n212), .A3(n271), .ZN(n320) );
  XNOR2_X1 U308 ( .A(n321), .B(n322), .ZN(n38) );
  OR2_X1 U309 ( .A1(n321), .A2(n322), .ZN(n37) );
  OAI22_X1 U310 ( .A1(n293), .A2(n288), .B1(n262), .B2(n323), .ZN(n322) );
  XNOR2_X1 U311 ( .A(b[5]), .B(a[3]), .ZN(n293) );
  OAI22_X1 U312 ( .A1(n310), .A2(n309), .B1(n307), .B2(n311), .ZN(n321) );
  XNOR2_X1 U313 ( .A(b[2]), .B(a[7]), .ZN(n311) );
  XNOR2_X1 U314 ( .A(b[1]), .B(a[7]), .ZN(n310) );
  OAI22_X1 U315 ( .A1(n323), .A2(n288), .B1(n262), .B2(n295), .ZN(n31) );
  XNOR2_X1 U316 ( .A(b[7]), .B(a[3]), .ZN(n295) );
  XNOR2_X1 U317 ( .A(n277), .B(a[2]), .ZN(n324) );
  XNOR2_X1 U318 ( .A(b[6]), .B(a[3]), .ZN(n323) );
  OAI22_X1 U319 ( .A1(n304), .A2(n298), .B1(n296), .B2(n306), .ZN(n21) );
  XNOR2_X1 U320 ( .A(b[7]), .B(a[5]), .ZN(n306) );
  XNOR2_X1 U321 ( .A(n274), .B(a[4]), .ZN(n325) );
  XNOR2_X1 U322 ( .A(b[6]), .B(a[5]), .ZN(n304) );
  OAI22_X1 U323 ( .A1(n315), .A2(n309), .B1(n307), .B2(n317), .ZN(n15) );
  XNOR2_X1 U324 ( .A(b[7]), .B(a[7]), .ZN(n317) );
  NAND2_X1 U325 ( .A1(n307), .A2(n326), .ZN(n309) );
  XNOR2_X1 U326 ( .A(n271), .B(a[6]), .ZN(n326) );
  XNOR2_X1 U327 ( .A(b[6]), .B(a[7]), .ZN(n315) );
  OAI22_X1 U328 ( .A1(n267), .A2(n282), .B1(n327), .B2(n280), .ZN(n104) );
  OAI22_X1 U329 ( .A1(n327), .A2(n282), .B1(n328), .B2(n280), .ZN(n103) );
  XNOR2_X1 U330 ( .A(b[1]), .B(a[1]), .ZN(n327) );
  OAI22_X1 U331 ( .A1(n328), .A2(n282), .B1(n329), .B2(n280), .ZN(n102) );
  XNOR2_X1 U332 ( .A(b[2]), .B(a[1]), .ZN(n328) );
  OAI22_X1 U333 ( .A1(n329), .A2(n282), .B1(n330), .B2(n280), .ZN(n101) );
  XNOR2_X1 U334 ( .A(b[3]), .B(a[1]), .ZN(n329) );
  OAI22_X1 U335 ( .A1(n330), .A2(n282), .B1(n281), .B2(n280), .ZN(n100) );
  XNOR2_X1 U336 ( .A(b[5]), .B(a[1]), .ZN(n281) );
  NAND2_X1 U337 ( .A1(a[1]), .A2(n280), .ZN(n282) );
  XNOR2_X1 U338 ( .A(b[4]), .B(a[1]), .ZN(n330) );
endmodule


module datapath_DW01_add_7 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n64;
  wire   [15:1] carry;

  FA_X1 U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n64), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  NAND3_X1 U1 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n1) );
  NAND3_X1 U2 ( .A1(n53), .A2(n54), .A3(n55), .ZN(n2) );
  NAND3_X1 U3 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n3) );
  XOR2_X1 U4 ( .A(B[3]), .B(A[3]), .Z(n4) );
  XOR2_X1 U5 ( .A(carry[3]), .B(n4), .Z(SUM[3]) );
  NAND2_X1 U6 ( .A1(carry[3]), .A2(B[3]), .ZN(n5) );
  NAND2_X1 U7 ( .A1(carry[3]), .A2(A[3]), .ZN(n6) );
  NAND2_X1 U8 ( .A1(B[3]), .A2(A[3]), .ZN(n7) );
  NAND3_X1 U9 ( .A1(n5), .A2(n6), .A3(n7), .ZN(carry[4]) );
  XNOR2_X1 U10 ( .A(carry[15]), .B(n8), .ZN(SUM[15]) );
  XNOR2_X1 U11 ( .A(B[15]), .B(A[15]), .ZN(n8) );
  XOR2_X1 U12 ( .A(B[11]), .B(A[11]), .Z(n9) );
  XOR2_X1 U13 ( .A(carry[11]), .B(n9), .Z(SUM[11]) );
  NAND2_X1 U14 ( .A1(carry[11]), .A2(B[11]), .ZN(n10) );
  NAND2_X1 U15 ( .A1(carry[11]), .A2(A[11]), .ZN(n11) );
  NAND2_X1 U16 ( .A1(B[11]), .A2(A[11]), .ZN(n12) );
  NAND3_X1 U17 ( .A1(n10), .A2(n11), .A3(n12), .ZN(carry[12]) );
  NAND3_X1 U18 ( .A1(n17), .A2(n18), .A3(n19), .ZN(n13) );
  NAND3_X1 U19 ( .A1(n32), .A2(n33), .A3(n34), .ZN(n14) );
  NAND3_X1 U20 ( .A1(n32), .A2(n33), .A3(n34), .ZN(n15) );
  XOR2_X1 U21 ( .A(B[5]), .B(A[5]), .Z(n16) );
  XOR2_X1 U22 ( .A(n15), .B(n16), .Z(SUM[5]) );
  NAND2_X1 U23 ( .A1(n14), .A2(B[5]), .ZN(n17) );
  NAND2_X1 U24 ( .A1(carry[5]), .A2(A[5]), .ZN(n18) );
  NAND2_X1 U25 ( .A1(B[5]), .A2(A[5]), .ZN(n19) );
  NAND3_X1 U26 ( .A1(n17), .A2(n18), .A3(n19), .ZN(carry[6]) );
  CLKBUF_X1 U27 ( .A(carry[12]), .Z(n20) );
  NAND3_X1 U28 ( .A1(n36), .A2(n37), .A3(n38), .ZN(n21) );
  NAND3_X1 U29 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n22) );
  NAND3_X1 U30 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n23) );
  XNOR2_X1 U31 ( .A(n2), .B(n24), .ZN(SUM[14]) );
  XNOR2_X1 U32 ( .A(B[14]), .B(A[14]), .ZN(n24) );
  CLKBUF_X1 U33 ( .A(n3), .Z(n25) );
  NAND3_X1 U34 ( .A1(n60), .A2(n61), .A3(n62), .ZN(n26) );
  XOR2_X1 U35 ( .A(B[9]), .B(A[9]), .Z(n27) );
  XOR2_X1 U36 ( .A(carry[9]), .B(n27), .Z(SUM[9]) );
  NAND2_X1 U37 ( .A1(n26), .A2(B[9]), .ZN(n28) );
  NAND2_X1 U38 ( .A1(n26), .A2(A[9]), .ZN(n29) );
  NAND2_X1 U39 ( .A1(B[9]), .A2(A[9]), .ZN(n30) );
  NAND3_X1 U40 ( .A1(n28), .A2(n29), .A3(n30), .ZN(carry[10]) );
  XOR2_X1 U41 ( .A(carry[4]), .B(A[4]), .Z(n31) );
  XOR2_X1 U42 ( .A(B[4]), .B(n31), .Z(SUM[4]) );
  NAND2_X1 U43 ( .A1(carry[4]), .A2(B[4]), .ZN(n32) );
  NAND2_X1 U44 ( .A1(B[4]), .A2(A[4]), .ZN(n33) );
  NAND2_X1 U45 ( .A1(carry[4]), .A2(A[4]), .ZN(n34) );
  NAND3_X1 U46 ( .A1(n32), .A2(n33), .A3(n34), .ZN(carry[5]) );
  XOR2_X1 U47 ( .A(B[6]), .B(A[6]), .Z(n35) );
  XOR2_X1 U48 ( .A(n13), .B(n35), .Z(SUM[6]) );
  NAND2_X1 U49 ( .A1(n13), .A2(B[6]), .ZN(n36) );
  NAND2_X1 U50 ( .A1(carry[6]), .A2(A[6]), .ZN(n37) );
  NAND2_X1 U51 ( .A1(B[6]), .A2(A[6]), .ZN(n38) );
  NAND3_X1 U52 ( .A1(n36), .A2(n37), .A3(n38), .ZN(carry[7]) );
  NAND3_X1 U53 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n39) );
  XOR2_X1 U54 ( .A(B[10]), .B(A[10]), .Z(n40) );
  XOR2_X1 U55 ( .A(n25), .B(n40), .Z(SUM[10]) );
  NAND2_X1 U56 ( .A1(n3), .A2(B[10]), .ZN(n41) );
  NAND2_X1 U57 ( .A1(carry[10]), .A2(A[10]), .ZN(n42) );
  NAND2_X1 U58 ( .A1(B[10]), .A2(A[10]), .ZN(n43) );
  NAND3_X1 U59 ( .A1(n41), .A2(n42), .A3(n43), .ZN(carry[11]) );
  XOR2_X1 U60 ( .A(B[7]), .B(A[7]), .Z(n44) );
  XOR2_X1 U61 ( .A(n21), .B(n44), .Z(SUM[7]) );
  NAND2_X1 U62 ( .A1(n21), .A2(B[7]), .ZN(n45) );
  NAND2_X1 U63 ( .A1(carry[7]), .A2(A[7]), .ZN(n46) );
  NAND2_X1 U64 ( .A1(B[7]), .A2(A[7]), .ZN(n47) );
  NAND3_X1 U65 ( .A1(n45), .A2(n46), .A3(n47), .ZN(carry[8]) );
  XOR2_X1 U66 ( .A(A[12]), .B(B[12]), .Z(n48) );
  XOR2_X1 U67 ( .A(n48), .B(n20), .Z(SUM[12]) );
  NAND2_X1 U68 ( .A1(A[12]), .A2(B[12]), .ZN(n49) );
  NAND2_X1 U69 ( .A1(A[12]), .A2(carry[12]), .ZN(n50) );
  NAND2_X1 U70 ( .A1(carry[12]), .A2(B[12]), .ZN(n51) );
  NAND3_X1 U71 ( .A1(n49), .A2(n50), .A3(n51), .ZN(carry[13]) );
  XOR2_X1 U72 ( .A(B[13]), .B(A[13]), .Z(n52) );
  XOR2_X1 U73 ( .A(n52), .B(n23), .Z(SUM[13]) );
  NAND2_X1 U74 ( .A1(B[13]), .A2(A[13]), .ZN(n53) );
  NAND2_X1 U75 ( .A1(B[13]), .A2(n22), .ZN(n54) );
  NAND2_X1 U76 ( .A1(A[13]), .A2(carry[13]), .ZN(n55) );
  NAND3_X1 U77 ( .A1(n53), .A2(n54), .A3(n55), .ZN(carry[14]) );
  NAND2_X1 U78 ( .A1(B[14]), .A2(carry[14]), .ZN(n56) );
  NAND2_X1 U79 ( .A1(n1), .A2(A[14]), .ZN(n57) );
  NAND2_X1 U80 ( .A1(B[14]), .A2(A[14]), .ZN(n58) );
  NAND3_X1 U81 ( .A1(n56), .A2(n57), .A3(n58), .ZN(carry[15]) );
  XOR2_X1 U82 ( .A(B[8]), .B(A[8]), .Z(n59) );
  XOR2_X1 U83 ( .A(carry[8]), .B(n59), .Z(SUM[8]) );
  NAND2_X1 U84 ( .A1(n39), .A2(B[8]), .ZN(n60) );
  NAND2_X1 U85 ( .A1(n39), .A2(A[8]), .ZN(n61) );
  NAND2_X1 U86 ( .A1(B[8]), .A2(A[8]), .ZN(n62) );
  NAND3_X1 U87 ( .A1(n60), .A2(n61), .A3(n62), .ZN(carry[9]) );
  XOR2_X1 U88 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U89 ( .A1(B[0]), .A2(A[0]), .ZN(n64) );
endmodule


module datapath_DW_mult_tc_6 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340;

  FA_X1 U11 ( .A(n50), .B(n53), .CI(n11), .CO(n10), .S(product[5]) );
  FA_X1 U12 ( .A(n54), .B(n206), .CI(n12), .CO(n11), .S(product[4]) );
  FA_X1 U13 ( .A(n56), .B(n71), .CI(n13), .CO(n12), .S(product[3]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n283), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n282), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n286), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n285), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n288), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  NAND3_X1 U157 ( .A1(n264), .A2(n265), .A3(n266), .ZN(n49) );
  INV_X1 U158 ( .A(n15), .ZN(n279) );
  AND2_X1 U159 ( .A1(n95), .A2(n102), .ZN(n206) );
  AND3_X1 U160 ( .A1(n267), .A2(n268), .A3(n269), .ZN(product[15]) );
  XNOR2_X1 U161 ( .A(n280), .B(n15), .ZN(n208) );
  NAND3_X1 U162 ( .A1(n220), .A2(n221), .A3(n222), .ZN(n209) );
  NAND3_X1 U163 ( .A1(n220), .A2(n221), .A3(n222), .ZN(n210) );
  INV_X1 U164 ( .A(n289), .ZN(n211) );
  INV_X1 U165 ( .A(n270), .ZN(n212) );
  OAI22_X1 U166 ( .A1(n231), .A2(n292), .B1(n338), .B2(n290), .ZN(n213) );
  XNOR2_X1 U167 ( .A(n52), .B(n214), .ZN(n50) );
  XNOR2_X1 U168 ( .A(n100), .B(n93), .ZN(n214) );
  NAND3_X1 U169 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n215) );
  NAND3_X1 U170 ( .A1(n227), .A2(n228), .A3(n229), .ZN(n216) );
  NAND3_X1 U171 ( .A1(n227), .A2(n228), .A3(n229), .ZN(n217) );
  NAND3_X1 U172 ( .A1(n249), .A2(n250), .A3(n251), .ZN(n218) );
  XOR2_X1 U173 ( .A(n46), .B(n49), .Z(n219) );
  XOR2_X1 U174 ( .A(n10), .B(n219), .Z(product[6]) );
  NAND2_X1 U175 ( .A1(n10), .A2(n46), .ZN(n220) );
  NAND2_X1 U176 ( .A1(n10), .A2(n49), .ZN(n221) );
  NAND2_X1 U177 ( .A1(n46), .A2(n49), .ZN(n222) );
  NAND3_X1 U178 ( .A1(n220), .A2(n221), .A3(n222), .ZN(n9) );
  XNOR2_X1 U179 ( .A(n218), .B(n223), .ZN(product[10]) );
  XNOR2_X1 U180 ( .A(n27), .B(n24), .ZN(n223) );
  XNOR2_X1 U181 ( .A(n260), .B(n224), .ZN(product[12]) );
  AND3_X1 U182 ( .A1(n259), .A2(n258), .A3(n257), .ZN(n224) );
  XNOR2_X1 U183 ( .A(n256), .B(n225), .ZN(product[11]) );
  AND3_X1 U184 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n225) );
  XNOR2_X1 U185 ( .A(n2), .B(n208), .ZN(product[14]) );
  XOR2_X2 U186 ( .A(a[6]), .B(n284), .Z(n317) );
  XOR2_X1 U187 ( .A(n40), .B(n45), .Z(n226) );
  XOR2_X1 U188 ( .A(n210), .B(n226), .Z(product[7]) );
  NAND2_X1 U189 ( .A1(n209), .A2(n40), .ZN(n227) );
  NAND2_X1 U190 ( .A1(n9), .A2(n45), .ZN(n228) );
  NAND2_X1 U191 ( .A1(n40), .A2(n45), .ZN(n229) );
  NAND3_X1 U192 ( .A1(n227), .A2(n228), .A3(n229), .ZN(n8) );
  NAND3_X1 U193 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n230) );
  BUF_X1 U194 ( .A(n337), .Z(n231) );
  XOR2_X1 U195 ( .A(n17), .B(n279), .Z(n232) );
  XOR2_X1 U196 ( .A(n3), .B(n232), .Z(product[13]) );
  NAND2_X1 U197 ( .A1(n215), .A2(n17), .ZN(n233) );
  NAND2_X1 U198 ( .A1(n3), .A2(n279), .ZN(n234) );
  NAND2_X1 U199 ( .A1(n17), .A2(n279), .ZN(n235) );
  NAND3_X1 U200 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n2) );
  CLKBUF_X1 U201 ( .A(b[3]), .Z(n236) );
  NAND3_X1 U202 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n237) );
  XOR2_X1 U203 ( .A(n34), .B(n39), .Z(n238) );
  XOR2_X1 U204 ( .A(n217), .B(n238), .Z(product[8]) );
  NAND2_X1 U205 ( .A1(n216), .A2(n34), .ZN(n239) );
  NAND2_X1 U206 ( .A1(n8), .A2(n39), .ZN(n240) );
  NAND2_X1 U207 ( .A1(n34), .A2(n39), .ZN(n241) );
  NAND3_X1 U208 ( .A1(n239), .A2(n240), .A3(n241), .ZN(n7) );
  XOR2_X1 U209 ( .A(n95), .B(n102), .Z(n56) );
  XNOR2_X1 U210 ( .A(n14), .B(n242), .ZN(product[2]) );
  XNOR2_X1 U211 ( .A(n103), .B(n96), .ZN(n242) );
  NAND3_X1 U212 ( .A1(n259), .A2(n258), .A3(n257), .ZN(n243) );
  NAND3_X1 U213 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n244) );
  NAND2_X1 U214 ( .A1(n14), .A2(n213), .ZN(n245) );
  NAND2_X1 U215 ( .A1(n14), .A2(n96), .ZN(n246) );
  NAND2_X1 U216 ( .A1(n213), .A2(n96), .ZN(n247) );
  NAND3_X1 U217 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n13) );
  XOR2_X1 U218 ( .A(n33), .B(n28), .Z(n248) );
  XOR2_X1 U219 ( .A(n7), .B(n248), .Z(product[9]) );
  NAND2_X1 U220 ( .A1(n237), .A2(n33), .ZN(n249) );
  NAND2_X1 U221 ( .A1(n7), .A2(n28), .ZN(n250) );
  NAND2_X1 U222 ( .A1(n33), .A2(n28), .ZN(n251) );
  NAND3_X1 U223 ( .A1(n249), .A2(n250), .A3(n251), .ZN(n6) );
  NAND2_X1 U224 ( .A1(n218), .A2(n27), .ZN(n252) );
  NAND2_X1 U225 ( .A1(n6), .A2(n24), .ZN(n253) );
  NAND2_X1 U226 ( .A1(n27), .A2(n24), .ZN(n254) );
  NAND3_X1 U227 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n5) );
  CLKBUF_X1 U228 ( .A(b[1]), .Z(n255) );
  XOR2_X1 U229 ( .A(n20), .B(n23), .Z(n256) );
  NAND2_X1 U230 ( .A1(n20), .A2(n23), .ZN(n257) );
  NAND2_X1 U231 ( .A1(n20), .A2(n5), .ZN(n258) );
  NAND2_X1 U232 ( .A1(n23), .A2(n244), .ZN(n259) );
  NAND3_X1 U233 ( .A1(n258), .A2(n259), .A3(n257), .ZN(n4) );
  XOR2_X1 U234 ( .A(n19), .B(n18), .Z(n260) );
  NAND2_X1 U235 ( .A1(n19), .A2(n18), .ZN(n261) );
  NAND2_X1 U236 ( .A1(n19), .A2(n243), .ZN(n262) );
  NAND2_X1 U237 ( .A1(n18), .A2(n4), .ZN(n263) );
  NAND3_X1 U238 ( .A1(n261), .A2(n262), .A3(n263), .ZN(n3) );
  NAND2_X2 U239 ( .A1(n296), .A2(n334), .ZN(n298) );
  NAND2_X1 U240 ( .A1(n52), .A2(n100), .ZN(n264) );
  NAND2_X1 U241 ( .A1(n52), .A2(n93), .ZN(n265) );
  NAND2_X1 U242 ( .A1(n100), .A2(n93), .ZN(n266) );
  NAND2_X1 U243 ( .A1(n230), .A2(n280), .ZN(n267) );
  NAND2_X1 U244 ( .A1(n230), .A2(n15), .ZN(n268) );
  NAND2_X1 U245 ( .A1(n280), .A2(n15), .ZN(n269) );
  BUF_X2 U246 ( .A(n306), .Z(n276) );
  INV_X1 U247 ( .A(n278), .ZN(n270) );
  INV_X1 U248 ( .A(n296), .ZN(n271) );
  INV_X1 U249 ( .A(n271), .ZN(n272) );
  NAND2_X1 U250 ( .A1(n274), .A2(n275), .ZN(n296) );
  INV_X1 U251 ( .A(a[0]), .ZN(n290) );
  NAND2_X1 U252 ( .A1(a[2]), .A2(a[1]), .ZN(n274) );
  NAND2_X1 U253 ( .A1(n273), .A2(n289), .ZN(n275) );
  INV_X1 U254 ( .A(a[2]), .ZN(n273) );
  INV_X1 U255 ( .A(n21), .ZN(n282) );
  INV_X1 U256 ( .A(n315), .ZN(n283) );
  INV_X1 U257 ( .A(n326), .ZN(n280) );
  INV_X1 U258 ( .A(n295), .ZN(n288) );
  INV_X1 U259 ( .A(n304), .ZN(n286) );
  INV_X1 U260 ( .A(n31), .ZN(n285) );
  INV_X1 U261 ( .A(b[0]), .ZN(n278) );
  NAND2_X1 U262 ( .A1(n306), .A2(n335), .ZN(n308) );
  INV_X1 U263 ( .A(a[5]), .ZN(n284) );
  INV_X1 U264 ( .A(a[7]), .ZN(n281) );
  XOR2_X1 U265 ( .A(a[4]), .B(n287), .Z(n306) );
  INV_X1 U266 ( .A(a[3]), .ZN(n287) );
  INV_X1 U267 ( .A(a[1]), .ZN(n289) );
  INV_X1 U268 ( .A(n278), .ZN(n277) );
  NOR2_X1 U269 ( .A1(n290), .A2(n278), .ZN(product[0]) );
  OAI22_X1 U270 ( .A1(n291), .A2(n292), .B1(n293), .B2(n290), .ZN(n99) );
  OAI22_X1 U271 ( .A1(n293), .A2(n292), .B1(n294), .B2(n290), .ZN(n98) );
  XNOR2_X1 U272 ( .A(b[6]), .B(n211), .ZN(n293) );
  OAI22_X1 U273 ( .A1(n290), .A2(n294), .B1(n292), .B2(n294), .ZN(n295) );
  XNOR2_X1 U274 ( .A(b[7]), .B(n211), .ZN(n294) );
  NOR2_X1 U275 ( .A1(n296), .A2(n278), .ZN(n96) );
  OAI22_X1 U276 ( .A1(n297), .A2(n298), .B1(n296), .B2(n299), .ZN(n95) );
  XNOR2_X1 U277 ( .A(a[3]), .B(n277), .ZN(n297) );
  OAI22_X1 U278 ( .A1(n299), .A2(n298), .B1(n272), .B2(n300), .ZN(n94) );
  XNOR2_X1 U279 ( .A(b[1]), .B(a[3]), .ZN(n299) );
  OAI22_X1 U280 ( .A1(n300), .A2(n298), .B1(n272), .B2(n301), .ZN(n93) );
  XNOR2_X1 U281 ( .A(b[2]), .B(a[3]), .ZN(n300) );
  OAI22_X1 U282 ( .A1(n301), .A2(n298), .B1(n272), .B2(n302), .ZN(n92) );
  XNOR2_X1 U283 ( .A(b[3]), .B(a[3]), .ZN(n301) );
  OAI22_X1 U284 ( .A1(n302), .A2(n298), .B1(n272), .B2(n303), .ZN(n91) );
  XNOR2_X1 U285 ( .A(b[4]), .B(a[3]), .ZN(n302) );
  OAI22_X1 U286 ( .A1(n305), .A2(n272), .B1(n298), .B2(n305), .ZN(n304) );
  NOR2_X1 U287 ( .A1(n276), .A2(n212), .ZN(n88) );
  OAI22_X1 U288 ( .A1(n307), .A2(n308), .B1(n276), .B2(n309), .ZN(n87) );
  XNOR2_X1 U289 ( .A(a[5]), .B(n270), .ZN(n307) );
  OAI22_X1 U290 ( .A1(n309), .A2(n308), .B1(n276), .B2(n310), .ZN(n86) );
  XNOR2_X1 U291 ( .A(n255), .B(a[5]), .ZN(n309) );
  OAI22_X1 U292 ( .A1(n310), .A2(n308), .B1(n276), .B2(n311), .ZN(n85) );
  XNOR2_X1 U293 ( .A(b[2]), .B(a[5]), .ZN(n310) );
  OAI22_X1 U294 ( .A1(n311), .A2(n308), .B1(n276), .B2(n312), .ZN(n84) );
  XNOR2_X1 U295 ( .A(n236), .B(a[5]), .ZN(n311) );
  OAI22_X1 U296 ( .A1(n312), .A2(n308), .B1(n276), .B2(n313), .ZN(n83) );
  XNOR2_X1 U297 ( .A(b[4]), .B(a[5]), .ZN(n312) );
  OAI22_X1 U298 ( .A1(n313), .A2(n308), .B1(n276), .B2(n314), .ZN(n82) );
  XNOR2_X1 U299 ( .A(b[5]), .B(a[5]), .ZN(n313) );
  OAI22_X1 U300 ( .A1(n316), .A2(n276), .B1(n308), .B2(n316), .ZN(n315) );
  NOR2_X1 U301 ( .A1(n317), .A2(n212), .ZN(n80) );
  OAI22_X1 U302 ( .A1(n318), .A2(n319), .B1(n317), .B2(n320), .ZN(n79) );
  XNOR2_X1 U303 ( .A(a[7]), .B(n270), .ZN(n318) );
  OAI22_X1 U304 ( .A1(n321), .A2(n319), .B1(n317), .B2(n322), .ZN(n77) );
  OAI22_X1 U305 ( .A1(n322), .A2(n319), .B1(n317), .B2(n323), .ZN(n76) );
  XNOR2_X1 U306 ( .A(n236), .B(a[7]), .ZN(n322) );
  OAI22_X1 U307 ( .A1(n323), .A2(n319), .B1(n317), .B2(n324), .ZN(n75) );
  XNOR2_X1 U308 ( .A(b[4]), .B(a[7]), .ZN(n323) );
  OAI22_X1 U309 ( .A1(n324), .A2(n319), .B1(n317), .B2(n325), .ZN(n74) );
  XNOR2_X1 U310 ( .A(b[5]), .B(a[7]), .ZN(n324) );
  OAI22_X1 U311 ( .A1(n327), .A2(n317), .B1(n319), .B2(n327), .ZN(n326) );
  OAI21_X1 U312 ( .B1(n277), .B2(n289), .A(n292), .ZN(n72) );
  OAI21_X1 U313 ( .B1(n287), .B2(n298), .A(n328), .ZN(n71) );
  OR3_X1 U314 ( .A1(n296), .A2(n270), .A3(n287), .ZN(n328) );
  OAI21_X1 U315 ( .B1(n284), .B2(n308), .A(n329), .ZN(n70) );
  OR3_X1 U316 ( .A1(n276), .A2(n277), .A3(n284), .ZN(n329) );
  OAI21_X1 U317 ( .B1(n281), .B2(n319), .A(n330), .ZN(n69) );
  OR3_X1 U318 ( .A1(n317), .A2(n277), .A3(n281), .ZN(n330) );
  XNOR2_X1 U319 ( .A(n331), .B(n332), .ZN(n38) );
  OR2_X1 U320 ( .A1(n331), .A2(n332), .ZN(n37) );
  OAI22_X1 U321 ( .A1(n303), .A2(n298), .B1(n272), .B2(n333), .ZN(n332) );
  XNOR2_X1 U322 ( .A(b[5]), .B(a[3]), .ZN(n303) );
  OAI22_X1 U323 ( .A1(n320), .A2(n319), .B1(n317), .B2(n321), .ZN(n331) );
  XNOR2_X1 U324 ( .A(b[2]), .B(a[7]), .ZN(n321) );
  XNOR2_X1 U325 ( .A(n255), .B(a[7]), .ZN(n320) );
  OAI22_X1 U326 ( .A1(n333), .A2(n298), .B1(n272), .B2(n305), .ZN(n31) );
  XNOR2_X1 U327 ( .A(b[7]), .B(a[3]), .ZN(n305) );
  XNOR2_X1 U328 ( .A(n287), .B(a[2]), .ZN(n334) );
  XNOR2_X1 U329 ( .A(b[6]), .B(a[3]), .ZN(n333) );
  OAI22_X1 U330 ( .A1(n314), .A2(n308), .B1(n276), .B2(n316), .ZN(n21) );
  XNOR2_X1 U331 ( .A(b[7]), .B(a[5]), .ZN(n316) );
  XNOR2_X1 U332 ( .A(n284), .B(a[4]), .ZN(n335) );
  XNOR2_X1 U333 ( .A(b[6]), .B(a[5]), .ZN(n314) );
  OAI22_X1 U334 ( .A1(n325), .A2(n319), .B1(n317), .B2(n327), .ZN(n15) );
  XNOR2_X1 U335 ( .A(b[7]), .B(a[7]), .ZN(n327) );
  NAND2_X1 U336 ( .A1(n317), .A2(n336), .ZN(n319) );
  XNOR2_X1 U337 ( .A(n281), .B(a[6]), .ZN(n336) );
  XNOR2_X1 U338 ( .A(b[6]), .B(a[7]), .ZN(n325) );
  OAI22_X1 U339 ( .A1(n270), .A2(n292), .B1(n337), .B2(n290), .ZN(n104) );
  OAI22_X1 U340 ( .A1(n231), .A2(n292), .B1(n338), .B2(n290), .ZN(n103) );
  XNOR2_X1 U341 ( .A(b[1]), .B(a[1]), .ZN(n337) );
  OAI22_X1 U342 ( .A1(n292), .A2(n338), .B1(n339), .B2(n290), .ZN(n102) );
  XNOR2_X1 U343 ( .A(b[2]), .B(a[1]), .ZN(n338) );
  OAI22_X1 U344 ( .A1(n339), .A2(n292), .B1(n340), .B2(n290), .ZN(n101) );
  XNOR2_X1 U345 ( .A(b[3]), .B(a[1]), .ZN(n339) );
  OAI22_X1 U346 ( .A1(n340), .A2(n292), .B1(n291), .B2(n290), .ZN(n100) );
  XNOR2_X1 U347 ( .A(b[5]), .B(n211), .ZN(n291) );
  NAND2_X1 U348 ( .A1(a[1]), .A2(n290), .ZN(n292) );
  XNOR2_X1 U349 ( .A(b[4]), .B(a[1]), .ZN(n340) );
endmodule


module datapath_DW01_add_6 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n71;
  wire   [15:1] carry;

  FA_X1 U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n71), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  XNOR2_X1 U1 ( .A(B[15]), .B(A[15]), .ZN(n57) );
  CLKBUF_X1 U2 ( .A(B[5]), .Z(n1) );
  CLKBUF_X1 U3 ( .A(n37), .Z(n2) );
  XNOR2_X1 U4 ( .A(n3), .B(n2), .ZN(SUM[14]) );
  XNOR2_X1 U5 ( .A(A[14]), .B(B[14]), .ZN(n3) );
  NAND3_X1 U6 ( .A1(n15), .A2(n16), .A3(n17), .ZN(n4) );
  NAND3_X1 U7 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n5) );
  NAND3_X1 U8 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n6) );
  CLKBUF_X1 U9 ( .A(n30), .Z(n7) );
  XOR2_X1 U10 ( .A(carry[3]), .B(A[3]), .Z(n8) );
  XOR2_X1 U11 ( .A(B[3]), .B(n8), .Z(SUM[3]) );
  NAND2_X1 U12 ( .A1(B[3]), .A2(carry[3]), .ZN(n9) );
  NAND2_X1 U13 ( .A1(B[3]), .A2(A[3]), .ZN(n10) );
  NAND2_X1 U14 ( .A1(carry[3]), .A2(A[3]), .ZN(n11) );
  NAND3_X1 U15 ( .A1(n9), .A2(n10), .A3(n11), .ZN(carry[4]) );
  CLKBUF_X1 U16 ( .A(n64), .Z(n12) );
  CLKBUF_X1 U17 ( .A(n60), .Z(n13) );
  XOR2_X1 U18 ( .A(B[10]), .B(A[10]), .Z(n14) );
  XOR2_X1 U19 ( .A(n6), .B(n14), .Z(SUM[10]) );
  NAND2_X1 U20 ( .A1(n5), .A2(B[10]), .ZN(n15) );
  NAND2_X1 U21 ( .A1(carry[10]), .A2(A[10]), .ZN(n16) );
  NAND2_X1 U22 ( .A1(B[10]), .A2(A[10]), .ZN(n17) );
  NAND3_X1 U23 ( .A1(n15), .A2(n16), .A3(n17), .ZN(carry[11]) );
  NAND3_X1 U24 ( .A1(n22), .A2(n23), .A3(n24), .ZN(n18) );
  NAND3_X1 U25 ( .A1(n22), .A2(n23), .A3(n24), .ZN(n19) );
  CLKBUF_X1 U26 ( .A(n65), .Z(n20) );
  XOR2_X1 U27 ( .A(B[4]), .B(A[4]), .Z(n21) );
  XOR2_X1 U28 ( .A(carry[4]), .B(n21), .Z(SUM[4]) );
  NAND2_X1 U29 ( .A1(carry[4]), .A2(B[4]), .ZN(n22) );
  NAND2_X1 U30 ( .A1(carry[4]), .A2(A[4]), .ZN(n23) );
  NAND2_X1 U31 ( .A1(B[4]), .A2(A[4]), .ZN(n24) );
  NAND3_X1 U32 ( .A1(n22), .A2(n23), .A3(n24), .ZN(carry[5]) );
  NAND3_X1 U33 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n25) );
  XOR2_X1 U34 ( .A(B[11]), .B(A[11]), .Z(n26) );
  XOR2_X1 U35 ( .A(n4), .B(n26), .Z(SUM[11]) );
  NAND2_X1 U36 ( .A1(n4), .A2(B[11]), .ZN(n27) );
  NAND2_X1 U37 ( .A1(carry[11]), .A2(A[11]), .ZN(n28) );
  NAND2_X1 U38 ( .A1(B[11]), .A2(A[11]), .ZN(n29) );
  NAND3_X1 U39 ( .A1(n27), .A2(n28), .A3(n29), .ZN(carry[12]) );
  NAND3_X1 U40 ( .A1(n67), .A2(n68), .A3(n69), .ZN(n30) );
  NAND3_X1 U41 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n31) );
  XOR2_X1 U42 ( .A(B[12]), .B(A[12]), .Z(n32) );
  XOR2_X1 U43 ( .A(carry[12]), .B(n32), .Z(SUM[12]) );
  NAND2_X1 U44 ( .A1(n25), .A2(B[12]), .ZN(n33) );
  NAND2_X1 U45 ( .A1(carry[12]), .A2(A[12]), .ZN(n34) );
  NAND2_X1 U46 ( .A1(B[12]), .A2(A[12]), .ZN(n35) );
  NAND3_X1 U47 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[13]) );
  NAND3_X1 U48 ( .A1(n46), .A2(n47), .A3(n48), .ZN(n36) );
  NAND3_X1 U49 ( .A1(n39), .A2(n40), .A3(n41), .ZN(n37) );
  XOR2_X1 U50 ( .A(B[13]), .B(A[13]), .Z(n38) );
  XOR2_X1 U51 ( .A(n38), .B(n31), .Z(SUM[13]) );
  NAND2_X1 U52 ( .A1(B[13]), .A2(A[13]), .ZN(n39) );
  NAND2_X1 U53 ( .A1(B[13]), .A2(n31), .ZN(n40) );
  NAND2_X1 U54 ( .A1(A[13]), .A2(carry[13]), .ZN(n41) );
  NAND3_X1 U55 ( .A1(n39), .A2(n40), .A3(n41), .ZN(carry[14]) );
  NAND2_X1 U56 ( .A1(A[14]), .A2(B[14]), .ZN(n42) );
  NAND2_X1 U57 ( .A1(A[14]), .A2(n37), .ZN(n43) );
  NAND2_X1 U58 ( .A1(B[14]), .A2(carry[14]), .ZN(n44) );
  NAND3_X1 U59 ( .A1(n42), .A2(n43), .A3(n44), .ZN(carry[15]) );
  XOR2_X1 U60 ( .A(B[8]), .B(A[8]), .Z(n45) );
  XOR2_X1 U61 ( .A(n7), .B(n45), .Z(SUM[8]) );
  NAND2_X1 U62 ( .A1(n30), .A2(B[8]), .ZN(n46) );
  NAND2_X1 U63 ( .A1(carry[8]), .A2(A[8]), .ZN(n47) );
  NAND2_X1 U64 ( .A1(B[8]), .A2(A[8]), .ZN(n48) );
  NAND3_X1 U65 ( .A1(n46), .A2(n47), .A3(n48), .ZN(carry[9]) );
  NAND3_X1 U66 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n49) );
  NAND3_X1 U67 ( .A1(n59), .A2(n13), .A3(n61), .ZN(n50) );
  NAND3_X1 U68 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n51) );
  NAND3_X1 U69 ( .A1(n63), .A2(n12), .A3(n20), .ZN(n52) );
  XOR2_X1 U70 ( .A(n36), .B(A[9]), .Z(n53) );
  XOR2_X1 U71 ( .A(B[9]), .B(n53), .Z(SUM[9]) );
  NAND2_X1 U72 ( .A1(B[9]), .A2(n36), .ZN(n54) );
  NAND2_X1 U73 ( .A1(B[9]), .A2(A[9]), .ZN(n55) );
  NAND2_X1 U74 ( .A1(carry[9]), .A2(A[9]), .ZN(n56) );
  NAND3_X1 U75 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[10]) );
  XNOR2_X1 U76 ( .A(carry[15]), .B(n57), .ZN(SUM[15]) );
  XOR2_X1 U77 ( .A(n1), .B(A[5]), .Z(n58) );
  XOR2_X1 U78 ( .A(n19), .B(n58), .Z(SUM[5]) );
  NAND2_X1 U79 ( .A1(carry[5]), .A2(B[5]), .ZN(n59) );
  NAND2_X1 U80 ( .A1(n18), .A2(A[5]), .ZN(n60) );
  NAND2_X1 U81 ( .A1(B[5]), .A2(A[5]), .ZN(n61) );
  NAND3_X1 U82 ( .A1(n59), .A2(n60), .A3(n61), .ZN(carry[6]) );
  XOR2_X1 U83 ( .A(A[6]), .B(B[6]), .Z(n62) );
  XOR2_X1 U84 ( .A(n62), .B(n50), .Z(SUM[6]) );
  NAND2_X1 U85 ( .A1(A[6]), .A2(B[6]), .ZN(n63) );
  NAND2_X1 U86 ( .A1(A[6]), .A2(n49), .ZN(n64) );
  NAND2_X1 U87 ( .A1(B[6]), .A2(carry[6]), .ZN(n65) );
  NAND3_X1 U88 ( .A1(n63), .A2(n64), .A3(n65), .ZN(carry[7]) );
  XOR2_X1 U89 ( .A(A[7]), .B(B[7]), .Z(n66) );
  XOR2_X1 U90 ( .A(n66), .B(n52), .Z(SUM[7]) );
  NAND2_X1 U91 ( .A1(A[7]), .A2(B[7]), .ZN(n67) );
  NAND2_X1 U92 ( .A1(A[7]), .A2(n51), .ZN(n68) );
  NAND2_X1 U93 ( .A1(B[7]), .A2(carry[7]), .ZN(n69) );
  NAND3_X1 U94 ( .A1(n67), .A2(n68), .A3(n69), .ZN(carry[8]) );
  XOR2_X1 U95 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U96 ( .A1(B[0]), .A2(A[0]), .ZN(n71) );
endmodule


module datapath_DW_mult_tc_5 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n10, n11, n12, n13, n15, n17, n18, n19,
         n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76, n77,
         n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94, n95,
         n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339;

  FA_X1 U17 ( .A(n74), .B(n21), .CI(n283), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n282), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n286), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n285), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n287), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  NAND2_X1 U157 ( .A1(n305), .A2(n334), .ZN(n307) );
  XNOR2_X1 U158 ( .A(n207), .B(n251), .ZN(product[2]) );
  AND2_X1 U159 ( .A1(n95), .A2(n102), .ZN(n206) );
  AND2_X1 U160 ( .A1(n104), .A2(n72), .ZN(n207) );
  XNOR2_X1 U161 ( .A(n280), .B(n15), .ZN(n208) );
  AND3_X1 U162 ( .A1(n224), .A2(n225), .A3(n226), .ZN(product[15]) );
  INV_X1 U163 ( .A(n278), .ZN(n210) );
  INV_X1 U164 ( .A(n278), .ZN(n277) );
  NAND3_X1 U165 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n211) );
  NAND3_X1 U166 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n212) );
  NAND3_X1 U167 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n213) );
  NAND3_X1 U168 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n214) );
  NAND3_X1 U169 ( .A1(n221), .A2(n222), .A3(n223), .ZN(n215) );
  NAND3_X1 U170 ( .A1(n221), .A2(n222), .A3(n223), .ZN(n216) );
  XNOR2_X1 U171 ( .A(n217), .B(n13), .ZN(product[3]) );
  XNOR2_X1 U172 ( .A(n56), .B(n71), .ZN(n217) );
  NAND2_X2 U173 ( .A1(n316), .A2(n335), .ZN(n318) );
  XOR2_X2 U174 ( .A(a[6]), .B(n284), .Z(n316) );
  XOR2_X1 U175 ( .A(n218), .B(n219), .Z(product[9]) );
  AND3_X1 U176 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n218) );
  XNOR2_X1 U177 ( .A(n33), .B(n28), .ZN(n219) );
  XNOR2_X1 U178 ( .A(n2), .B(n208), .ZN(product[14]) );
  XOR2_X1 U179 ( .A(n104), .B(n72), .Z(product[1]) );
  XOR2_X1 U180 ( .A(n50), .B(n53), .Z(n220) );
  XOR2_X1 U181 ( .A(n214), .B(n220), .Z(product[5]) );
  NAND2_X1 U182 ( .A1(n213), .A2(n50), .ZN(n221) );
  NAND2_X1 U183 ( .A1(n11), .A2(n53), .ZN(n222) );
  NAND2_X1 U184 ( .A1(n50), .A2(n53), .ZN(n223) );
  NAND3_X1 U185 ( .A1(n221), .A2(n222), .A3(n223), .ZN(n10) );
  NAND2_X1 U186 ( .A1(n2), .A2(n280), .ZN(n224) );
  NAND2_X1 U187 ( .A1(n2), .A2(n15), .ZN(n225) );
  NAND2_X1 U188 ( .A1(n280), .A2(n15), .ZN(n226) );
  XOR2_X1 U189 ( .A(n46), .B(n49), .Z(n227) );
  XOR2_X1 U190 ( .A(n216), .B(n227), .Z(product[6]) );
  NAND2_X1 U191 ( .A1(n215), .A2(n46), .ZN(n228) );
  NAND2_X1 U192 ( .A1(n10), .A2(n49), .ZN(n229) );
  NAND2_X1 U193 ( .A1(n46), .A2(n49), .ZN(n230) );
  XOR2_X1 U194 ( .A(n18), .B(n19), .Z(n231) );
  XOR2_X1 U195 ( .A(n4), .B(n231), .Z(product[12]) );
  NAND2_X1 U196 ( .A1(n4), .A2(n18), .ZN(n232) );
  NAND2_X1 U197 ( .A1(n4), .A2(n19), .ZN(n233) );
  NAND2_X1 U198 ( .A1(n18), .A2(n19), .ZN(n234) );
  NAND3_X1 U199 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n3) );
  NAND3_X1 U200 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n235) );
  XOR2_X1 U201 ( .A(n95), .B(n102), .Z(n236) );
  XOR2_X1 U202 ( .A(n40), .B(n45), .Z(n237) );
  XOR2_X1 U203 ( .A(n212), .B(n237), .Z(product[7]) );
  NAND2_X1 U204 ( .A1(n212), .A2(n40), .ZN(n238) );
  NAND2_X1 U205 ( .A1(n211), .A2(n45), .ZN(n239) );
  NAND2_X1 U206 ( .A1(n40), .A2(n45), .ZN(n240) );
  NAND3_X1 U207 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n8) );
  NAND3_X1 U208 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n241) );
  XOR2_X1 U209 ( .A(n34), .B(n39), .Z(n242) );
  XOR2_X1 U210 ( .A(n8), .B(n242), .Z(product[8]) );
  NAND2_X1 U211 ( .A1(n235), .A2(n34), .ZN(n243) );
  NAND2_X1 U212 ( .A1(n8), .A2(n39), .ZN(n244) );
  NAND2_X1 U213 ( .A1(n34), .A2(n39), .ZN(n245) );
  NAND3_X1 U214 ( .A1(n243), .A2(n244), .A3(n245), .ZN(n7) );
  NAND2_X1 U215 ( .A1(n7), .A2(n33), .ZN(n246) );
  NAND2_X1 U216 ( .A1(n241), .A2(n28), .ZN(n247) );
  NAND2_X1 U217 ( .A1(n33), .A2(n28), .ZN(n248) );
  NAND3_X1 U218 ( .A1(n247), .A2(n246), .A3(n248), .ZN(n6) );
  NAND3_X1 U219 ( .A1(n257), .A2(n256), .A3(n255), .ZN(n249) );
  NAND3_X1 U220 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n250) );
  XNOR2_X2 U221 ( .A(a[4]), .B(a[3]), .ZN(n305) );
  XNOR2_X1 U222 ( .A(n103), .B(n96), .ZN(n251) );
  NAND2_X1 U223 ( .A1(n207), .A2(n103), .ZN(n252) );
  NAND2_X1 U224 ( .A1(n207), .A2(n96), .ZN(n253) );
  NAND2_X1 U225 ( .A1(n103), .A2(n96), .ZN(n254) );
  NAND3_X1 U226 ( .A1(n252), .A2(n253), .A3(n254), .ZN(n13) );
  NAND2_X1 U227 ( .A1(n236), .A2(n71), .ZN(n255) );
  NAND2_X1 U228 ( .A1(n236), .A2(n13), .ZN(n256) );
  NAND2_X1 U229 ( .A1(n71), .A2(n13), .ZN(n257) );
  NAND3_X1 U230 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n12) );
  XOR2_X1 U231 ( .A(n54), .B(n206), .Z(n258) );
  XOR2_X1 U232 ( .A(n258), .B(n250), .Z(product[4]) );
  NAND2_X1 U233 ( .A1(n54), .A2(n206), .ZN(n259) );
  NAND2_X1 U234 ( .A1(n54), .A2(n249), .ZN(n260) );
  NAND2_X1 U235 ( .A1(n206), .A2(n12), .ZN(n261) );
  NAND3_X1 U236 ( .A1(n259), .A2(n260), .A3(n261), .ZN(n11) );
  XOR2_X1 U237 ( .A(n24), .B(n27), .Z(n262) );
  XOR2_X1 U238 ( .A(n262), .B(n6), .Z(product[10]) );
  NAND2_X1 U239 ( .A1(n24), .A2(n27), .ZN(n263) );
  NAND2_X1 U240 ( .A1(n24), .A2(n6), .ZN(n264) );
  NAND2_X1 U241 ( .A1(n27), .A2(n6), .ZN(n265) );
  NAND3_X1 U242 ( .A1(n263), .A2(n264), .A3(n265), .ZN(n5) );
  XOR2_X1 U243 ( .A(n20), .B(n23), .Z(n266) );
  XOR2_X1 U244 ( .A(n266), .B(n5), .Z(product[11]) );
  NAND2_X1 U245 ( .A1(n20), .A2(n23), .ZN(n267) );
  NAND2_X1 U246 ( .A1(n20), .A2(n5), .ZN(n268) );
  NAND2_X1 U247 ( .A1(n23), .A2(n5), .ZN(n269) );
  NAND3_X1 U248 ( .A1(n269), .A2(n268), .A3(n267), .ZN(n4) );
  XOR2_X1 U249 ( .A(n17), .B(n279), .Z(n270) );
  XOR2_X1 U250 ( .A(n3), .B(n270), .Z(product[13]) );
  NAND2_X1 U251 ( .A1(n3), .A2(n17), .ZN(n271) );
  NAND2_X1 U252 ( .A1(n3), .A2(n279), .ZN(n272) );
  NAND2_X1 U253 ( .A1(n17), .A2(n279), .ZN(n273) );
  NAND3_X1 U254 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n2) );
  XOR2_X1 U255 ( .A(n95), .B(n102), .Z(n56) );
  XNOR2_X1 U256 ( .A(a[2]), .B(a[1]), .ZN(n274) );
  INV_X1 U257 ( .A(a[0]), .ZN(n289) );
  INV_X1 U258 ( .A(n15), .ZN(n279) );
  INV_X1 U259 ( .A(n21), .ZN(n282) );
  INV_X1 U260 ( .A(n314), .ZN(n283) );
  INV_X1 U261 ( .A(n325), .ZN(n280) );
  INV_X1 U262 ( .A(n294), .ZN(n287) );
  INV_X1 U263 ( .A(n303), .ZN(n286) );
  INV_X1 U264 ( .A(n31), .ZN(n285) );
  INV_X1 U265 ( .A(b[0]), .ZN(n278) );
  XNOR2_X1 U266 ( .A(a[2]), .B(a[1]), .ZN(n295) );
  INV_X1 U267 ( .A(n275), .ZN(n276) );
  NAND2_X1 U268 ( .A1(n295), .A2(n333), .ZN(n297) );
  INV_X1 U269 ( .A(a[5]), .ZN(n284) );
  INV_X1 U270 ( .A(a[7]), .ZN(n281) );
  INV_X1 U271 ( .A(a[3]), .ZN(n275) );
  INV_X1 U272 ( .A(a[1]), .ZN(n288) );
  NOR2_X1 U273 ( .A1(n289), .A2(n278), .ZN(product[0]) );
  OAI22_X1 U274 ( .A1(n290), .A2(n291), .B1(n292), .B2(n289), .ZN(n99) );
  OAI22_X1 U275 ( .A1(n292), .A2(n291), .B1(n293), .B2(n289), .ZN(n98) );
  XNOR2_X1 U276 ( .A(b[6]), .B(a[1]), .ZN(n292) );
  OAI22_X1 U277 ( .A1(n289), .A2(n293), .B1(n291), .B2(n293), .ZN(n294) );
  XNOR2_X1 U278 ( .A(b[7]), .B(a[1]), .ZN(n293) );
  NOR2_X1 U279 ( .A1(n274), .A2(n278), .ZN(n96) );
  OAI22_X1 U280 ( .A1(n296), .A2(n297), .B1(n274), .B2(n298), .ZN(n95) );
  XNOR2_X1 U281 ( .A(n276), .B(n210), .ZN(n296) );
  OAI22_X1 U282 ( .A1(n298), .A2(n297), .B1(n274), .B2(n299), .ZN(n94) );
  XNOR2_X1 U283 ( .A(b[1]), .B(n276), .ZN(n298) );
  OAI22_X1 U284 ( .A1(n299), .A2(n297), .B1(n274), .B2(n300), .ZN(n93) );
  XNOR2_X1 U285 ( .A(b[2]), .B(n276), .ZN(n299) );
  OAI22_X1 U286 ( .A1(n300), .A2(n297), .B1(n274), .B2(n301), .ZN(n92) );
  XNOR2_X1 U287 ( .A(b[3]), .B(n276), .ZN(n300) );
  OAI22_X1 U288 ( .A1(n301), .A2(n297), .B1(n274), .B2(n302), .ZN(n91) );
  XNOR2_X1 U289 ( .A(b[4]), .B(n276), .ZN(n301) );
  OAI22_X1 U290 ( .A1(n304), .A2(n274), .B1(n297), .B2(n304), .ZN(n303) );
  NOR2_X1 U291 ( .A1(n305), .A2(n278), .ZN(n88) );
  OAI22_X1 U292 ( .A1(n306), .A2(n307), .B1(n305), .B2(n308), .ZN(n87) );
  XNOR2_X1 U293 ( .A(a[5]), .B(n277), .ZN(n306) );
  OAI22_X1 U294 ( .A1(n308), .A2(n307), .B1(n305), .B2(n309), .ZN(n86) );
  XNOR2_X1 U295 ( .A(b[1]), .B(a[5]), .ZN(n308) );
  OAI22_X1 U296 ( .A1(n309), .A2(n307), .B1(n305), .B2(n310), .ZN(n85) );
  XNOR2_X1 U297 ( .A(b[2]), .B(a[5]), .ZN(n309) );
  OAI22_X1 U298 ( .A1(n310), .A2(n307), .B1(n305), .B2(n311), .ZN(n84) );
  XNOR2_X1 U299 ( .A(b[3]), .B(a[5]), .ZN(n310) );
  OAI22_X1 U300 ( .A1(n311), .A2(n307), .B1(n305), .B2(n312), .ZN(n83) );
  XNOR2_X1 U301 ( .A(b[4]), .B(a[5]), .ZN(n311) );
  OAI22_X1 U302 ( .A1(n312), .A2(n307), .B1(n305), .B2(n313), .ZN(n82) );
  XNOR2_X1 U303 ( .A(b[5]), .B(a[5]), .ZN(n312) );
  OAI22_X1 U304 ( .A1(n315), .A2(n305), .B1(n307), .B2(n315), .ZN(n314) );
  NOR2_X1 U305 ( .A1(n316), .A2(n278), .ZN(n80) );
  OAI22_X1 U306 ( .A1(n317), .A2(n318), .B1(n316), .B2(n319), .ZN(n79) );
  XNOR2_X1 U307 ( .A(a[7]), .B(n210), .ZN(n317) );
  OAI22_X1 U308 ( .A1(n320), .A2(n318), .B1(n316), .B2(n321), .ZN(n77) );
  OAI22_X1 U309 ( .A1(n321), .A2(n318), .B1(n316), .B2(n322), .ZN(n76) );
  XNOR2_X1 U310 ( .A(b[3]), .B(a[7]), .ZN(n321) );
  OAI22_X1 U311 ( .A1(n322), .A2(n318), .B1(n316), .B2(n323), .ZN(n75) );
  XNOR2_X1 U312 ( .A(b[4]), .B(a[7]), .ZN(n322) );
  OAI22_X1 U313 ( .A1(n323), .A2(n318), .B1(n316), .B2(n324), .ZN(n74) );
  XNOR2_X1 U314 ( .A(b[5]), .B(a[7]), .ZN(n323) );
  OAI22_X1 U315 ( .A1(n326), .A2(n316), .B1(n318), .B2(n326), .ZN(n325) );
  OAI21_X1 U316 ( .B1(n210), .B2(n288), .A(n291), .ZN(n72) );
  OAI21_X1 U317 ( .B1(n275), .B2(n297), .A(n327), .ZN(n71) );
  OR3_X1 U318 ( .A1(n274), .A2(n210), .A3(n275), .ZN(n327) );
  OAI21_X1 U319 ( .B1(n284), .B2(n307), .A(n328), .ZN(n70) );
  OR3_X1 U320 ( .A1(n305), .A2(n277), .A3(n284), .ZN(n328) );
  OAI21_X1 U321 ( .B1(n281), .B2(n318), .A(n329), .ZN(n69) );
  OR3_X1 U322 ( .A1(n316), .A2(n210), .A3(n281), .ZN(n329) );
  XNOR2_X1 U323 ( .A(n330), .B(n331), .ZN(n38) );
  OR2_X1 U324 ( .A1(n330), .A2(n331), .ZN(n37) );
  OAI22_X1 U325 ( .A1(n302), .A2(n297), .B1(n274), .B2(n332), .ZN(n331) );
  XNOR2_X1 U326 ( .A(b[5]), .B(n276), .ZN(n302) );
  OAI22_X1 U327 ( .A1(n319), .A2(n318), .B1(n316), .B2(n320), .ZN(n330) );
  XNOR2_X1 U328 ( .A(b[2]), .B(a[7]), .ZN(n320) );
  XNOR2_X1 U329 ( .A(b[1]), .B(a[7]), .ZN(n319) );
  OAI22_X1 U330 ( .A1(n332), .A2(n297), .B1(n274), .B2(n304), .ZN(n31) );
  XNOR2_X1 U331 ( .A(b[7]), .B(n276), .ZN(n304) );
  XNOR2_X1 U332 ( .A(n275), .B(a[2]), .ZN(n333) );
  XNOR2_X1 U333 ( .A(b[6]), .B(n276), .ZN(n332) );
  OAI22_X1 U334 ( .A1(n313), .A2(n307), .B1(n305), .B2(n315), .ZN(n21) );
  XNOR2_X1 U335 ( .A(b[7]), .B(a[5]), .ZN(n315) );
  XNOR2_X1 U336 ( .A(n284), .B(a[4]), .ZN(n334) );
  XNOR2_X1 U337 ( .A(b[6]), .B(a[5]), .ZN(n313) );
  OAI22_X1 U338 ( .A1(n324), .A2(n318), .B1(n316), .B2(n326), .ZN(n15) );
  XNOR2_X1 U339 ( .A(b[7]), .B(a[7]), .ZN(n326) );
  XNOR2_X1 U340 ( .A(n281), .B(a[6]), .ZN(n335) );
  XNOR2_X1 U341 ( .A(b[6]), .B(a[7]), .ZN(n324) );
  OAI22_X1 U342 ( .A1(n277), .A2(n291), .B1(n336), .B2(n289), .ZN(n104) );
  OAI22_X1 U343 ( .A1(n336), .A2(n291), .B1(n337), .B2(n289), .ZN(n103) );
  XNOR2_X1 U344 ( .A(b[1]), .B(a[1]), .ZN(n336) );
  OAI22_X1 U345 ( .A1(n337), .A2(n291), .B1(n338), .B2(n289), .ZN(n102) );
  XNOR2_X1 U346 ( .A(b[2]), .B(a[1]), .ZN(n337) );
  OAI22_X1 U347 ( .A1(n338), .A2(n291), .B1(n339), .B2(n289), .ZN(n101) );
  XNOR2_X1 U348 ( .A(b[3]), .B(a[1]), .ZN(n338) );
  OAI22_X1 U349 ( .A1(n339), .A2(n291), .B1(n290), .B2(n289), .ZN(n100) );
  XNOR2_X1 U350 ( .A(b[5]), .B(a[1]), .ZN(n290) );
  NAND2_X1 U351 ( .A1(a[1]), .A2(n289), .ZN(n291) );
  XNOR2_X1 U352 ( .A(b[4]), .B(a[1]), .ZN(n339) );
endmodule


module datapath_DW01_add_5 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n71;
  wire   [15:1] carry;

  FA_X1 U1_1 ( .A(A[1]), .B(n71), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[14]), .ZN(n40) );
  XOR2_X1 U2 ( .A(B[2]), .B(A[2]), .Z(n1) );
  XOR2_X1 U3 ( .A(carry[2]), .B(n1), .Z(SUM[2]) );
  NAND2_X1 U4 ( .A1(carry[2]), .A2(B[2]), .ZN(n2) );
  NAND2_X1 U5 ( .A1(carry[2]), .A2(A[2]), .ZN(n3) );
  NAND2_X1 U6 ( .A1(B[2]), .A2(A[2]), .ZN(n4) );
  NAND3_X1 U7 ( .A1(n2), .A2(n3), .A3(n4), .ZN(carry[3]) );
  NAND3_X1 U8 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n5) );
  NAND3_X1 U9 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n6) );
  CLKBUF_X1 U10 ( .A(n23), .Z(n7) );
  NAND3_X1 U11 ( .A1(n27), .A2(n28), .A3(n29), .ZN(n8) );
  NAND3_X1 U12 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n9) );
  NAND3_X1 U13 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n10) );
  NAND3_X1 U14 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n11) );
  NAND3_X1 U15 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n12) );
  XOR2_X1 U16 ( .A(B[13]), .B(A[13]), .Z(n13) );
  XOR2_X1 U17 ( .A(carry[13]), .B(n13), .Z(SUM[13]) );
  NAND2_X1 U18 ( .A1(carry[13]), .A2(B[13]), .ZN(n14) );
  NAND2_X1 U19 ( .A1(carry[13]), .A2(A[13]), .ZN(n15) );
  NAND2_X1 U20 ( .A1(B[13]), .A2(A[13]), .ZN(n16) );
  NAND3_X1 U21 ( .A1(n15), .A2(n14), .A3(n16), .ZN(carry[14]) );
  XOR2_X1 U22 ( .A(B[5]), .B(A[5]), .Z(n17) );
  XOR2_X1 U23 ( .A(n12), .B(n17), .Z(SUM[5]) );
  NAND2_X1 U24 ( .A1(n12), .A2(B[5]), .ZN(n18) );
  NAND2_X1 U25 ( .A1(carry[5]), .A2(A[5]), .ZN(n19) );
  NAND2_X1 U26 ( .A1(B[5]), .A2(A[5]), .ZN(n20) );
  NAND3_X1 U27 ( .A1(n18), .A2(n19), .A3(n20), .ZN(carry[6]) );
  CLKBUF_X1 U28 ( .A(n8), .Z(n21) );
  NAND3_X1 U29 ( .A1(n42), .A2(n43), .A3(n44), .ZN(n22) );
  NAND3_X1 U30 ( .A1(n52), .A2(n51), .A3(n50), .ZN(n23) );
  NAND3_X1 U31 ( .A1(n31), .A2(n32), .A3(n33), .ZN(n24) );
  NAND3_X1 U32 ( .A1(n31), .A2(n32), .A3(n33), .ZN(n25) );
  XOR2_X1 U33 ( .A(B[9]), .B(A[9]), .Z(n26) );
  XOR2_X1 U34 ( .A(n10), .B(n26), .Z(SUM[9]) );
  NAND2_X1 U35 ( .A1(n9), .A2(B[9]), .ZN(n27) );
  NAND2_X1 U36 ( .A1(carry[9]), .A2(A[9]), .ZN(n28) );
  NAND2_X1 U37 ( .A1(B[9]), .A2(A[9]), .ZN(n29) );
  NAND3_X1 U38 ( .A1(n27), .A2(n28), .A3(n29), .ZN(carry[10]) );
  XOR2_X1 U39 ( .A(B[6]), .B(A[6]), .Z(n30) );
  XOR2_X1 U40 ( .A(n6), .B(n30), .Z(SUM[6]) );
  NAND2_X1 U41 ( .A1(carry[6]), .A2(B[6]), .ZN(n31) );
  NAND2_X1 U42 ( .A1(n5), .A2(A[6]), .ZN(n32) );
  NAND2_X1 U43 ( .A1(B[6]), .A2(A[6]), .ZN(n33) );
  XOR2_X1 U44 ( .A(B[10]), .B(A[10]), .Z(n34) );
  XOR2_X1 U45 ( .A(n21), .B(n34), .Z(SUM[10]) );
  NAND2_X1 U46 ( .A1(n8), .A2(B[10]), .ZN(n35) );
  NAND2_X1 U47 ( .A1(carry[10]), .A2(A[10]), .ZN(n36) );
  NAND2_X1 U48 ( .A1(B[10]), .A2(A[10]), .ZN(n37) );
  NAND3_X1 U49 ( .A1(n35), .A2(n36), .A3(n37), .ZN(carry[11]) );
  NAND3_X1 U50 ( .A1(n58), .A2(n59), .A3(n60), .ZN(n38) );
  XNOR2_X1 U51 ( .A(carry[15]), .B(n39), .ZN(SUM[15]) );
  XNOR2_X1 U52 ( .A(B[15]), .B(A[15]), .ZN(n39) );
  XNOR2_X1 U53 ( .A(B[14]), .B(n40), .ZN(n66) );
  XOR2_X1 U54 ( .A(B[11]), .B(A[11]), .Z(n41) );
  XOR2_X1 U55 ( .A(carry[11]), .B(n41), .Z(SUM[11]) );
  NAND2_X1 U56 ( .A1(carry[11]), .A2(B[11]), .ZN(n42) );
  NAND2_X1 U57 ( .A1(carry[11]), .A2(A[11]), .ZN(n43) );
  NAND2_X1 U58 ( .A1(B[11]), .A2(A[11]), .ZN(n44) );
  NAND3_X1 U59 ( .A1(n42), .A2(n43), .A3(n44), .ZN(carry[12]) );
  XOR2_X1 U60 ( .A(B[12]), .B(A[12]), .Z(n45) );
  XOR2_X1 U61 ( .A(carry[12]), .B(n45), .Z(SUM[12]) );
  NAND2_X1 U62 ( .A1(n22), .A2(B[12]), .ZN(n46) );
  NAND2_X1 U63 ( .A1(n22), .A2(A[12]), .ZN(n47) );
  NAND2_X1 U64 ( .A1(B[12]), .A2(A[12]), .ZN(n48) );
  NAND3_X1 U65 ( .A1(n46), .A2(n47), .A3(n48), .ZN(carry[13]) );
  XOR2_X1 U66 ( .A(A[7]), .B(B[7]), .Z(n49) );
  XOR2_X1 U67 ( .A(n49), .B(n25), .Z(SUM[7]) );
  NAND2_X1 U68 ( .A1(A[7]), .A2(B[7]), .ZN(n50) );
  NAND2_X1 U69 ( .A1(A[7]), .A2(n24), .ZN(n51) );
  NAND2_X1 U70 ( .A1(B[7]), .A2(n24), .ZN(n52) );
  NAND3_X1 U71 ( .A1(n50), .A2(n51), .A3(n52), .ZN(carry[8]) );
  XOR2_X1 U72 ( .A(A[8]), .B(B[8]), .Z(n53) );
  XOR2_X1 U73 ( .A(n53), .B(n7), .Z(SUM[8]) );
  NAND2_X1 U74 ( .A1(A[8]), .A2(B[8]), .ZN(n54) );
  NAND2_X1 U75 ( .A1(A[8]), .A2(n23), .ZN(n55) );
  NAND2_X1 U76 ( .A1(B[8]), .A2(carry[8]), .ZN(n56) );
  NAND3_X1 U77 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[9]) );
  XOR2_X1 U78 ( .A(B[3]), .B(A[3]), .Z(n57) );
  XOR2_X1 U79 ( .A(carry[3]), .B(n57), .Z(SUM[3]) );
  NAND2_X1 U80 ( .A1(carry[3]), .A2(B[3]), .ZN(n58) );
  NAND2_X1 U81 ( .A1(carry[3]), .A2(A[3]), .ZN(n59) );
  NAND2_X1 U82 ( .A1(B[3]), .A2(A[3]), .ZN(n60) );
  NAND3_X1 U83 ( .A1(n58), .A2(n59), .A3(n60), .ZN(carry[4]) );
  XOR2_X1 U84 ( .A(B[4]), .B(A[4]), .Z(n61) );
  XOR2_X1 U85 ( .A(carry[4]), .B(n61), .Z(SUM[4]) );
  NAND2_X1 U86 ( .A1(n38), .A2(B[4]), .ZN(n62) );
  NAND2_X1 U87 ( .A1(carry[4]), .A2(A[4]), .ZN(n63) );
  NAND2_X1 U88 ( .A1(B[4]), .A2(A[4]), .ZN(n64) );
  NAND3_X1 U89 ( .A1(n62), .A2(n63), .A3(n64), .ZN(carry[5]) );
  CLKBUF_X1 U90 ( .A(n11), .Z(n65) );
  XOR2_X1 U91 ( .A(n65), .B(n66), .Z(SUM[14]) );
  NAND2_X1 U92 ( .A1(B[14]), .A2(carry[14]), .ZN(n67) );
  NAND2_X1 U93 ( .A1(n11), .A2(A[14]), .ZN(n68) );
  NAND2_X1 U94 ( .A1(B[14]), .A2(A[14]), .ZN(n69) );
  NAND3_X1 U95 ( .A1(n68), .A2(n67), .A3(n69), .ZN(carry[15]) );
  XOR2_X1 U96 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U97 ( .A1(B[0]), .A2(A[0]), .ZN(n71) );
endmodule


module datapath_DW_mult_tc_4 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339;

  FA_X1 U13 ( .A(n13), .B(n71), .CI(n56), .CO(n12), .S(product[3]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n282), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n281), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n285), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n284), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n287), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  AND2_X1 U157 ( .A1(n211), .A2(n102), .ZN(n206) );
  XNOR2_X1 U158 ( .A(n279), .B(n15), .ZN(n207) );
  XNOR2_X1 U159 ( .A(n17), .B(n278), .ZN(n208) );
  AND3_X1 U160 ( .A1(n259), .A2(n260), .A3(n261), .ZN(product[15]) );
  CLKBUF_X1 U161 ( .A(n305), .Z(n210) );
  XNOR2_X1 U162 ( .A(a[4]), .B(a[3]), .ZN(n305) );
  OAI22_X1 U163 ( .A1(n296), .A2(n297), .B1(n295), .B2(n298), .ZN(n211) );
  XOR2_X1 U164 ( .A(n46), .B(n49), .Z(n212) );
  XOR2_X1 U165 ( .A(n10), .B(n212), .Z(product[6]) );
  NAND2_X1 U166 ( .A1(n10), .A2(n46), .ZN(n213) );
  NAND2_X1 U167 ( .A1(n10), .A2(n49), .ZN(n214) );
  NAND2_X1 U168 ( .A1(n46), .A2(n49), .ZN(n215) );
  NAND3_X1 U169 ( .A1(n213), .A2(n214), .A3(n215), .ZN(n9) );
  NAND3_X1 U170 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n216) );
  NAND3_X1 U171 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n217) );
  NAND3_X1 U172 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n218) );
  NAND3_X1 U173 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n219) );
  NAND3_X1 U174 ( .A1(n268), .A2(n267), .A3(n266), .ZN(n220) );
  NAND3_X1 U175 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n221) );
  NAND3_X1 U176 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n222) );
  XOR2_X1 U177 ( .A(n40), .B(n45), .Z(n223) );
  XOR2_X1 U178 ( .A(n9), .B(n223), .Z(product[7]) );
  NAND2_X1 U179 ( .A1(n9), .A2(n40), .ZN(n224) );
  NAND2_X1 U180 ( .A1(n9), .A2(n45), .ZN(n225) );
  NAND2_X1 U181 ( .A1(n40), .A2(n45), .ZN(n226) );
  NAND3_X1 U182 ( .A1(n224), .A2(n225), .A3(n226), .ZN(n8) );
  XNOR2_X1 U183 ( .A(n220), .B(n207), .ZN(product[14]) );
  XNOR2_X1 U184 ( .A(n208), .B(n242), .ZN(product[13]) );
  XOR2_X1 U185 ( .A(n54), .B(n206), .Z(n227) );
  XOR2_X1 U186 ( .A(n227), .B(n12), .Z(product[4]) );
  NAND2_X1 U187 ( .A1(n54), .A2(n206), .ZN(n228) );
  NAND2_X1 U188 ( .A1(n54), .A2(n12), .ZN(n229) );
  NAND2_X1 U189 ( .A1(n206), .A2(n12), .ZN(n230) );
  NAND3_X1 U190 ( .A1(n228), .A2(n229), .A3(n230), .ZN(n11) );
  XOR2_X1 U191 ( .A(n50), .B(n53), .Z(n231) );
  XOR2_X1 U192 ( .A(n231), .B(n219), .Z(product[5]) );
  NAND2_X1 U193 ( .A1(n50), .A2(n53), .ZN(n232) );
  NAND2_X1 U194 ( .A1(n50), .A2(n218), .ZN(n233) );
  NAND2_X1 U195 ( .A1(n53), .A2(n11), .ZN(n234) );
  NAND3_X1 U196 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n10) );
  XOR2_X1 U197 ( .A(n33), .B(n28), .Z(n235) );
  XOR2_X1 U198 ( .A(n7), .B(n235), .Z(product[9]) );
  NAND2_X1 U199 ( .A1(n7), .A2(n33), .ZN(n236) );
  NAND2_X1 U200 ( .A1(n7), .A2(n28), .ZN(n237) );
  NAND2_X1 U201 ( .A1(n33), .A2(n28), .ZN(n238) );
  NAND3_X1 U202 ( .A1(n236), .A2(n237), .A3(n238), .ZN(n6) );
  BUF_X1 U203 ( .A(n336), .Z(n239) );
  NAND3_X1 U204 ( .A1(n249), .A2(n248), .A3(n250), .ZN(n240) );
  NAND3_X1 U205 ( .A1(n265), .A2(n264), .A3(n263), .ZN(n241) );
  NAND3_X1 U206 ( .A1(n263), .A2(n264), .A3(n265), .ZN(n242) );
  XOR2_X1 U207 ( .A(n34), .B(n39), .Z(n243) );
  XOR2_X1 U208 ( .A(n221), .B(n243), .Z(product[8]) );
  NAND2_X1 U209 ( .A1(n221), .A2(n34), .ZN(n244) );
  NAND2_X1 U210 ( .A1(n8), .A2(n39), .ZN(n245) );
  NAND2_X1 U211 ( .A1(n34), .A2(n39), .ZN(n246) );
  NAND3_X1 U212 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n7) );
  XOR2_X1 U213 ( .A(n27), .B(n24), .Z(n247) );
  XOR2_X1 U214 ( .A(n217), .B(n247), .Z(product[10]) );
  NAND2_X1 U215 ( .A1(n216), .A2(n27), .ZN(n248) );
  NAND2_X1 U216 ( .A1(n6), .A2(n24), .ZN(n249) );
  NAND2_X1 U217 ( .A1(n27), .A2(n24), .ZN(n250) );
  NAND3_X1 U218 ( .A1(n248), .A2(n249), .A3(n250), .ZN(n5) );
  NAND3_X1 U219 ( .A1(n268), .A2(n267), .A3(n266), .ZN(n251) );
  NAND3_X1 U220 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n252) );
  NAND3_X1 U221 ( .A1(n256), .A2(n255), .A3(n257), .ZN(n253) );
  XOR2_X1 U222 ( .A(n23), .B(n20), .Z(n254) );
  XOR2_X1 U223 ( .A(n222), .B(n254), .Z(product[11]) );
  NAND2_X1 U224 ( .A1(n240), .A2(n23), .ZN(n255) );
  NAND2_X1 U225 ( .A1(n5), .A2(n20), .ZN(n256) );
  NAND2_X1 U226 ( .A1(n23), .A2(n20), .ZN(n257) );
  NAND3_X1 U227 ( .A1(n255), .A2(n256), .A3(n257), .ZN(n4) );
  XNOR2_X1 U228 ( .A(n258), .B(n253), .ZN(product[12]) );
  XNOR2_X1 U229 ( .A(n19), .B(n18), .ZN(n258) );
  NAND2_X1 U230 ( .A1(n251), .A2(n279), .ZN(n259) );
  NAND2_X1 U231 ( .A1(n2), .A2(n15), .ZN(n260) );
  NAND2_X1 U232 ( .A1(n279), .A2(n15), .ZN(n261) );
  XOR2_X1 U233 ( .A(n95), .B(n102), .Z(n56) );
  CLKBUF_X1 U234 ( .A(b[1]), .Z(n262) );
  NAND2_X1 U235 ( .A1(n19), .A2(n18), .ZN(n263) );
  NAND2_X1 U236 ( .A1(n19), .A2(n252), .ZN(n264) );
  NAND2_X1 U237 ( .A1(n18), .A2(n4), .ZN(n265) );
  NAND3_X1 U238 ( .A1(n264), .A2(n263), .A3(n265), .ZN(n3) );
  NAND2_X1 U239 ( .A1(n17), .A2(n278), .ZN(n266) );
  NAND2_X1 U240 ( .A1(n17), .A2(n241), .ZN(n267) );
  NAND2_X1 U241 ( .A1(n278), .A2(n3), .ZN(n268) );
  NAND3_X1 U242 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n2) );
  INV_X2 U243 ( .A(n277), .ZN(n276) );
  BUF_X2 U244 ( .A(n295), .Z(n269) );
  XOR2_X1 U245 ( .A(a[2]), .B(n288), .Z(n295) );
  INV_X1 U246 ( .A(n15), .ZN(n278) );
  INV_X1 U247 ( .A(n21), .ZN(n281) );
  INV_X1 U248 ( .A(n314), .ZN(n282) );
  INV_X1 U249 ( .A(n325), .ZN(n279) );
  INV_X1 U250 ( .A(n294), .ZN(n287) );
  INV_X1 U251 ( .A(n303), .ZN(n285) );
  INV_X1 U252 ( .A(n31), .ZN(n284) );
  INV_X1 U253 ( .A(b[0]), .ZN(n277) );
  XNOR2_X1 U254 ( .A(n14), .B(n270), .ZN(product[2]) );
  XNOR2_X1 U255 ( .A(n103), .B(n96), .ZN(n270) );
  INV_X1 U256 ( .A(a[5]), .ZN(n283) );
  INV_X1 U257 ( .A(a[7]), .ZN(n280) );
  NAND2_X1 U258 ( .A1(n14), .A2(n103), .ZN(n271) );
  NAND2_X1 U259 ( .A1(n14), .A2(n96), .ZN(n272) );
  NAND2_X1 U260 ( .A1(n103), .A2(n96), .ZN(n273) );
  NAND3_X1 U261 ( .A1(n271), .A2(n272), .A3(n273), .ZN(n13) );
  INV_X1 U262 ( .A(a[3]), .ZN(n286) );
  NAND2_X2 U263 ( .A1(n305), .A2(n334), .ZN(n307) );
  INV_X1 U264 ( .A(a[1]), .ZN(n274) );
  INV_X2 U265 ( .A(n274), .ZN(n275) );
  NAND2_X2 U266 ( .A1(n295), .A2(n333), .ZN(n297) );
  INV_X1 U267 ( .A(a[1]), .ZN(n288) );
  XOR2_X2 U268 ( .A(a[6]), .B(n283), .Z(n316) );
  INV_X2 U269 ( .A(a[0]), .ZN(n289) );
  NOR2_X1 U270 ( .A1(n289), .A2(n277), .ZN(product[0]) );
  OAI22_X1 U271 ( .A1(n290), .A2(n291), .B1(n292), .B2(n289), .ZN(n99) );
  OAI22_X1 U272 ( .A1(n292), .A2(n291), .B1(n293), .B2(n289), .ZN(n98) );
  XNOR2_X1 U273 ( .A(b[6]), .B(n275), .ZN(n292) );
  OAI22_X1 U274 ( .A1(n289), .A2(n293), .B1(n291), .B2(n293), .ZN(n294) );
  XNOR2_X1 U275 ( .A(b[7]), .B(n275), .ZN(n293) );
  NOR2_X1 U276 ( .A1(n295), .A2(n277), .ZN(n96) );
  OAI22_X1 U277 ( .A1(n296), .A2(n297), .B1(n295), .B2(n298), .ZN(n95) );
  XNOR2_X1 U278 ( .A(a[3]), .B(n276), .ZN(n296) );
  OAI22_X1 U279 ( .A1(n298), .A2(n297), .B1(n269), .B2(n299), .ZN(n94) );
  XNOR2_X1 U280 ( .A(n262), .B(a[3]), .ZN(n298) );
  OAI22_X1 U281 ( .A1(n299), .A2(n297), .B1(n269), .B2(n300), .ZN(n93) );
  XNOR2_X1 U282 ( .A(b[2]), .B(a[3]), .ZN(n299) );
  OAI22_X1 U283 ( .A1(n300), .A2(n297), .B1(n269), .B2(n301), .ZN(n92) );
  XNOR2_X1 U284 ( .A(b[3]), .B(a[3]), .ZN(n300) );
  OAI22_X1 U285 ( .A1(n301), .A2(n297), .B1(n269), .B2(n302), .ZN(n91) );
  XNOR2_X1 U286 ( .A(b[4]), .B(a[3]), .ZN(n301) );
  OAI22_X1 U287 ( .A1(n304), .A2(n269), .B1(n297), .B2(n304), .ZN(n303) );
  NOR2_X1 U288 ( .A1(n305), .A2(n277), .ZN(n88) );
  OAI22_X1 U289 ( .A1(n306), .A2(n307), .B1(n305), .B2(n308), .ZN(n87) );
  XNOR2_X1 U290 ( .A(a[5]), .B(n276), .ZN(n306) );
  OAI22_X1 U291 ( .A1(n308), .A2(n307), .B1(n305), .B2(n309), .ZN(n86) );
  XNOR2_X1 U292 ( .A(n262), .B(a[5]), .ZN(n308) );
  OAI22_X1 U293 ( .A1(n309), .A2(n307), .B1(n305), .B2(n310), .ZN(n85) );
  XNOR2_X1 U294 ( .A(b[2]), .B(a[5]), .ZN(n309) );
  OAI22_X1 U295 ( .A1(n310), .A2(n307), .B1(n210), .B2(n311), .ZN(n84) );
  XNOR2_X1 U296 ( .A(b[3]), .B(a[5]), .ZN(n310) );
  OAI22_X1 U297 ( .A1(n311), .A2(n307), .B1(n210), .B2(n312), .ZN(n83) );
  XNOR2_X1 U298 ( .A(b[4]), .B(a[5]), .ZN(n311) );
  OAI22_X1 U299 ( .A1(n312), .A2(n307), .B1(n210), .B2(n313), .ZN(n82) );
  XNOR2_X1 U300 ( .A(b[5]), .B(a[5]), .ZN(n312) );
  OAI22_X1 U301 ( .A1(n315), .A2(n210), .B1(n307), .B2(n315), .ZN(n314) );
  NOR2_X1 U302 ( .A1(n316), .A2(n277), .ZN(n80) );
  OAI22_X1 U303 ( .A1(n317), .A2(n318), .B1(n316), .B2(n319), .ZN(n79) );
  XNOR2_X1 U304 ( .A(a[7]), .B(n276), .ZN(n317) );
  OAI22_X1 U305 ( .A1(n320), .A2(n318), .B1(n316), .B2(n321), .ZN(n77) );
  OAI22_X1 U306 ( .A1(n321), .A2(n318), .B1(n316), .B2(n322), .ZN(n76) );
  XNOR2_X1 U307 ( .A(b[3]), .B(a[7]), .ZN(n321) );
  OAI22_X1 U308 ( .A1(n322), .A2(n318), .B1(n316), .B2(n323), .ZN(n75) );
  XNOR2_X1 U309 ( .A(b[4]), .B(a[7]), .ZN(n322) );
  OAI22_X1 U310 ( .A1(n323), .A2(n318), .B1(n316), .B2(n324), .ZN(n74) );
  XNOR2_X1 U311 ( .A(b[5]), .B(a[7]), .ZN(n323) );
  OAI22_X1 U312 ( .A1(n326), .A2(n316), .B1(n318), .B2(n326), .ZN(n325) );
  OAI21_X1 U313 ( .B1(n276), .B2(n288), .A(n291), .ZN(n72) );
  OAI21_X1 U314 ( .B1(n286), .B2(n297), .A(n327), .ZN(n71) );
  OR3_X1 U315 ( .A1(n269), .A2(n276), .A3(n286), .ZN(n327) );
  OAI21_X1 U316 ( .B1(n283), .B2(n307), .A(n328), .ZN(n70) );
  OR3_X1 U317 ( .A1(n305), .A2(n276), .A3(n283), .ZN(n328) );
  OAI21_X1 U318 ( .B1(n280), .B2(n318), .A(n329), .ZN(n69) );
  OR3_X1 U319 ( .A1(n316), .A2(n276), .A3(n280), .ZN(n329) );
  XNOR2_X1 U320 ( .A(n330), .B(n331), .ZN(n38) );
  OR2_X1 U321 ( .A1(n330), .A2(n331), .ZN(n37) );
  OAI22_X1 U322 ( .A1(n302), .A2(n297), .B1(n269), .B2(n332), .ZN(n331) );
  XNOR2_X1 U323 ( .A(b[5]), .B(a[3]), .ZN(n302) );
  OAI22_X1 U324 ( .A1(n319), .A2(n318), .B1(n316), .B2(n320), .ZN(n330) );
  XNOR2_X1 U325 ( .A(b[2]), .B(a[7]), .ZN(n320) );
  XNOR2_X1 U326 ( .A(n262), .B(a[7]), .ZN(n319) );
  OAI22_X1 U327 ( .A1(n332), .A2(n297), .B1(n269), .B2(n304), .ZN(n31) );
  XNOR2_X1 U328 ( .A(b[7]), .B(a[3]), .ZN(n304) );
  XNOR2_X1 U329 ( .A(n286), .B(a[2]), .ZN(n333) );
  XNOR2_X1 U330 ( .A(b[6]), .B(a[3]), .ZN(n332) );
  OAI22_X1 U331 ( .A1(n313), .A2(n307), .B1(n210), .B2(n315), .ZN(n21) );
  XNOR2_X1 U332 ( .A(b[7]), .B(a[5]), .ZN(n315) );
  XNOR2_X1 U333 ( .A(n283), .B(a[4]), .ZN(n334) );
  XNOR2_X1 U334 ( .A(b[6]), .B(a[5]), .ZN(n313) );
  OAI22_X1 U335 ( .A1(n324), .A2(n318), .B1(n316), .B2(n326), .ZN(n15) );
  XNOR2_X1 U336 ( .A(b[7]), .B(a[7]), .ZN(n326) );
  NAND2_X1 U337 ( .A1(n316), .A2(n335), .ZN(n318) );
  XNOR2_X1 U338 ( .A(n280), .B(a[6]), .ZN(n335) );
  XNOR2_X1 U339 ( .A(b[6]), .B(a[7]), .ZN(n324) );
  OAI22_X1 U340 ( .A1(n276), .A2(n291), .B1(n336), .B2(n289), .ZN(n104) );
  OAI22_X1 U341 ( .A1(n291), .A2(n239), .B1(n337), .B2(n289), .ZN(n103) );
  XNOR2_X1 U342 ( .A(b[1]), .B(n275), .ZN(n336) );
  OAI22_X1 U343 ( .A1(n337), .A2(n291), .B1(n338), .B2(n289), .ZN(n102) );
  XNOR2_X1 U344 ( .A(b[2]), .B(n275), .ZN(n337) );
  OAI22_X1 U345 ( .A1(n338), .A2(n291), .B1(n339), .B2(n289), .ZN(n101) );
  XNOR2_X1 U346 ( .A(b[3]), .B(n275), .ZN(n338) );
  OAI22_X1 U347 ( .A1(n339), .A2(n291), .B1(n290), .B2(n289), .ZN(n100) );
  XNOR2_X1 U348 ( .A(b[5]), .B(n275), .ZN(n290) );
  NAND2_X1 U349 ( .A1(a[1]), .A2(n289), .ZN(n291) );
  XNOR2_X1 U350 ( .A(b[4]), .B(n275), .ZN(n339) );
endmodule


module datapath_DW01_add_4 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n73;
  wire   [15:1] carry;

  FA_X1 U1_3 ( .A(B[3]), .B(A[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n73), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[14]), .ZN(n44) );
  CLKBUF_X1 U2 ( .A(n58), .Z(n1) );
  CLKBUF_X1 U3 ( .A(carry[4]), .Z(n2) );
  NAND3_X1 U4 ( .A1(n58), .A2(n57), .A3(n56), .ZN(n3) );
  NAND3_X1 U5 ( .A1(n12), .A2(n13), .A3(n14), .ZN(n4) );
  CLKBUF_X1 U6 ( .A(n37), .Z(n5) );
  NAND3_X1 U7 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n6) );
  NAND3_X1 U8 ( .A1(n18), .A2(n19), .A3(n20), .ZN(n7) );
  CLKBUF_X1 U9 ( .A(carry[12]), .Z(n8) );
  NAND3_X1 U10 ( .A1(n31), .A2(n32), .A3(n33), .ZN(n9) );
  XNOR2_X1 U11 ( .A(n68), .B(n10), .ZN(SUM[14]) );
  AND3_X1 U12 ( .A1(n65), .A2(n66), .A3(n67), .ZN(n10) );
  XOR2_X1 U13 ( .A(B[4]), .B(A[4]), .Z(n11) );
  XOR2_X1 U14 ( .A(n2), .B(n11), .Z(SUM[4]) );
  NAND2_X1 U15 ( .A1(carry[4]), .A2(B[4]), .ZN(n12) );
  NAND2_X1 U16 ( .A1(carry[4]), .A2(A[4]), .ZN(n13) );
  NAND2_X1 U17 ( .A1(B[4]), .A2(A[4]), .ZN(n14) );
  NAND3_X1 U18 ( .A1(n12), .A2(n13), .A3(n14), .ZN(carry[5]) );
  CLKBUF_X1 U19 ( .A(n27), .Z(n15) );
  NAND3_X1 U20 ( .A1(n31), .A2(n32), .A3(n33), .ZN(n16) );
  XOR2_X1 U21 ( .A(B[6]), .B(A[6]), .Z(n17) );
  XOR2_X1 U22 ( .A(n16), .B(n17), .Z(SUM[6]) );
  NAND2_X1 U23 ( .A1(n9), .A2(B[6]), .ZN(n18) );
  NAND2_X1 U24 ( .A1(n16), .A2(A[6]), .ZN(n19) );
  NAND2_X1 U25 ( .A1(B[6]), .A2(A[6]), .ZN(n20) );
  NAND3_X1 U26 ( .A1(n18), .A2(n19), .A3(n20), .ZN(carry[7]) );
  NAND3_X1 U27 ( .A1(n41), .A2(n40), .A3(n42), .ZN(n21) );
  NAND3_X1 U28 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n22) );
  NAND3_X1 U29 ( .A1(n36), .A2(n37), .A3(n38), .ZN(n23) );
  NAND3_X1 U30 ( .A1(n36), .A2(n5), .A3(n38), .ZN(n24) );
  XOR2_X1 U31 ( .A(B[8]), .B(A[8]), .Z(n25) );
  XOR2_X1 U32 ( .A(n24), .B(n25), .Z(SUM[8]) );
  NAND2_X1 U33 ( .A1(n23), .A2(B[8]), .ZN(n26) );
  NAND2_X1 U34 ( .A1(carry[8]), .A2(A[8]), .ZN(n27) );
  NAND2_X1 U35 ( .A1(B[8]), .A2(A[8]), .ZN(n28) );
  NAND3_X1 U36 ( .A1(n26), .A2(n15), .A3(n28), .ZN(carry[9]) );
  NAND3_X1 U37 ( .A1(n61), .A2(n60), .A3(n62), .ZN(n29) );
  XOR2_X1 U38 ( .A(B[5]), .B(A[5]), .Z(n30) );
  XOR2_X1 U39 ( .A(n4), .B(n30), .Z(SUM[5]) );
  NAND2_X1 U40 ( .A1(n4), .A2(B[5]), .ZN(n31) );
  NAND2_X1 U41 ( .A1(carry[5]), .A2(A[5]), .ZN(n32) );
  NAND2_X1 U42 ( .A1(B[5]), .A2(A[5]), .ZN(n33) );
  XNOR2_X1 U43 ( .A(carry[15]), .B(n34), .ZN(SUM[15]) );
  XNOR2_X1 U44 ( .A(B[15]), .B(A[15]), .ZN(n34) );
  XOR2_X1 U45 ( .A(B[7]), .B(A[7]), .Z(n35) );
  XOR2_X1 U46 ( .A(n7), .B(n35), .Z(SUM[7]) );
  NAND2_X1 U47 ( .A1(n6), .A2(B[7]), .ZN(n36) );
  NAND2_X1 U48 ( .A1(carry[7]), .A2(A[7]), .ZN(n37) );
  NAND2_X1 U49 ( .A1(B[7]), .A2(A[7]), .ZN(n38) );
  NAND3_X1 U50 ( .A1(n36), .A2(n37), .A3(n38), .ZN(carry[8]) );
  XOR2_X1 U51 ( .A(B[12]), .B(A[12]), .Z(n39) );
  XOR2_X1 U52 ( .A(n8), .B(n39), .Z(SUM[12]) );
  NAND2_X1 U53 ( .A1(n29), .A2(B[12]), .ZN(n40) );
  NAND2_X1 U54 ( .A1(carry[12]), .A2(A[12]), .ZN(n41) );
  NAND2_X1 U55 ( .A1(B[12]), .A2(A[12]), .ZN(n42) );
  NAND3_X1 U56 ( .A1(n41), .A2(n40), .A3(n42), .ZN(carry[13]) );
  CLKBUF_X1 U57 ( .A(n50), .Z(n43) );
  XNOR2_X1 U58 ( .A(B[14]), .B(n44), .ZN(n68) );
  CLKBUF_X1 U59 ( .A(n57), .Z(n45) );
  NAND3_X1 U60 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n46) );
  NAND3_X1 U61 ( .A1(n49), .A2(n43), .A3(n51), .ZN(n47) );
  XOR2_X1 U62 ( .A(B[9]), .B(A[9]), .Z(n48) );
  XOR2_X1 U63 ( .A(carry[9]), .B(n48), .Z(SUM[9]) );
  NAND2_X1 U64 ( .A1(n22), .A2(B[9]), .ZN(n49) );
  NAND2_X1 U65 ( .A1(n22), .A2(A[9]), .ZN(n50) );
  NAND2_X1 U66 ( .A1(B[9]), .A2(A[9]), .ZN(n51) );
  NAND3_X1 U67 ( .A1(n50), .A2(n49), .A3(n51), .ZN(carry[10]) );
  NAND3_X1 U68 ( .A1(n58), .A2(n57), .A3(n56), .ZN(n52) );
  NAND3_X1 U69 ( .A1(n56), .A2(n45), .A3(n1), .ZN(n53) );
  CLKBUF_X1 U70 ( .A(carry[13]), .Z(n54) );
  XOR2_X1 U71 ( .A(A[10]), .B(B[10]), .Z(n55) );
  XOR2_X1 U72 ( .A(n55), .B(n47), .Z(SUM[10]) );
  NAND2_X1 U73 ( .A1(A[10]), .A2(B[10]), .ZN(n56) );
  NAND2_X1 U74 ( .A1(A[10]), .A2(n46), .ZN(n57) );
  NAND2_X1 U75 ( .A1(B[10]), .A2(carry[10]), .ZN(n58) );
  XOR2_X1 U76 ( .A(A[11]), .B(B[11]), .Z(n59) );
  XOR2_X1 U77 ( .A(n59), .B(n53), .Z(SUM[11]) );
  NAND2_X1 U78 ( .A1(A[11]), .A2(B[11]), .ZN(n60) );
  NAND2_X1 U79 ( .A1(n52), .A2(A[11]), .ZN(n61) );
  NAND2_X1 U80 ( .A1(n3), .A2(B[11]), .ZN(n62) );
  NAND3_X1 U81 ( .A1(n62), .A2(n61), .A3(n60), .ZN(carry[12]) );
  NAND3_X1 U82 ( .A1(n66), .A2(n67), .A3(n65), .ZN(n63) );
  XOR2_X1 U83 ( .A(A[13]), .B(B[13]), .Z(n64) );
  XOR2_X1 U84 ( .A(n64), .B(n54), .Z(SUM[13]) );
  NAND2_X1 U85 ( .A1(A[13]), .A2(B[13]), .ZN(n65) );
  NAND2_X1 U86 ( .A1(carry[13]), .A2(A[13]), .ZN(n66) );
  NAND2_X1 U87 ( .A1(B[13]), .A2(n21), .ZN(n67) );
  NAND3_X1 U88 ( .A1(n67), .A2(n66), .A3(n65), .ZN(carry[14]) );
  NAND2_X1 U89 ( .A1(B[14]), .A2(A[14]), .ZN(n69) );
  NAND2_X1 U90 ( .A1(A[14]), .A2(n63), .ZN(n70) );
  NAND2_X1 U91 ( .A1(carry[14]), .A2(B[14]), .ZN(n71) );
  NAND3_X1 U92 ( .A1(n70), .A2(n69), .A3(n71), .ZN(carry[15]) );
  XOR2_X1 U93 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U94 ( .A1(B[0]), .A2(A[0]), .ZN(n73) );
endmodule


module datapath_DW_mult_tc_3 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75,
         n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93,
         n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207,
         n208, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344;

  FA_X1 U11 ( .A(n50), .B(n53), .CI(n11), .CO(n10), .S(product[5]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n287), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n286), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n290), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n289), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n292), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  INV_X1 U157 ( .A(n15), .ZN(n283) );
  CLKBUF_X1 U158 ( .A(n102), .Z(n206) );
  OAI22_X1 U159 ( .A1(n251), .A2(n296), .B1(n342), .B2(n294), .ZN(n207) );
  XNOR2_X1 U160 ( .A(n284), .B(n15), .ZN(n208) );
  AND3_X1 U161 ( .A1(n243), .A2(n244), .A3(n245), .ZN(product[15]) );
  XOR2_X1 U162 ( .A(n102), .B(n211), .Z(n210) );
  OAI22_X1 U163 ( .A1(n301), .A2(n302), .B1(n276), .B2(n303), .ZN(n211) );
  NAND3_X1 U164 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n212) );
  NAND3_X1 U165 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n213) );
  BUF_X1 U166 ( .A(n341), .Z(n251) );
  XNOR2_X1 U167 ( .A(n2), .B(n208), .ZN(product[14]) );
  XNOR2_X1 U168 ( .A(n54), .B(n242), .ZN(n226) );
  NAND3_X1 U169 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n214) );
  XOR2_X1 U170 ( .A(n46), .B(n49), .Z(n215) );
  XOR2_X1 U171 ( .A(n10), .B(n215), .Z(product[6]) );
  NAND2_X1 U172 ( .A1(n10), .A2(n46), .ZN(n216) );
  NAND2_X1 U173 ( .A1(n10), .A2(n49), .ZN(n217) );
  NAND2_X1 U174 ( .A1(n46), .A2(n49), .ZN(n218) );
  NAND3_X1 U175 ( .A1(n216), .A2(n217), .A3(n218), .ZN(n9) );
  NAND3_X1 U176 ( .A1(n279), .A2(n278), .A3(n280), .ZN(n219) );
  NAND3_X1 U177 ( .A1(n223), .A2(n224), .A3(n225), .ZN(n220) );
  NAND3_X1 U178 ( .A1(n223), .A2(n224), .A3(n225), .ZN(n221) );
  XOR2_X2 U179 ( .A(a[6]), .B(n288), .Z(n321) );
  XOR2_X1 U180 ( .A(n56), .B(n71), .Z(n222) );
  XOR2_X1 U181 ( .A(n222), .B(n13), .Z(product[3]) );
  NAND2_X1 U182 ( .A1(n210), .A2(n71), .ZN(n223) );
  NAND2_X1 U183 ( .A1(n210), .A2(n219), .ZN(n224) );
  NAND2_X1 U184 ( .A1(n71), .A2(n219), .ZN(n225) );
  XOR2_X1 U185 ( .A(n226), .B(n221), .Z(product[4]) );
  NAND2_X1 U186 ( .A1(n54), .A2(n55), .ZN(n227) );
  NAND2_X1 U187 ( .A1(n54), .A2(n220), .ZN(n228) );
  NAND2_X1 U188 ( .A1(n55), .A2(n221), .ZN(n229) );
  NAND3_X1 U189 ( .A1(n229), .A2(n228), .A3(n227), .ZN(n11) );
  XOR2_X1 U190 ( .A(n40), .B(n45), .Z(n230) );
  XOR2_X1 U191 ( .A(n9), .B(n230), .Z(product[7]) );
  NAND2_X1 U192 ( .A1(n9), .A2(n40), .ZN(n231) );
  NAND2_X1 U193 ( .A1(n9), .A2(n45), .ZN(n232) );
  NAND2_X1 U194 ( .A1(n40), .A2(n45), .ZN(n233) );
  NAND3_X1 U195 ( .A1(n231), .A2(n232), .A3(n233), .ZN(n8) );
  NAND3_X1 U196 ( .A1(n248), .A2(n247), .A3(n249), .ZN(n234) );
  NAND3_X1 U197 ( .A1(n248), .A2(n247), .A3(n249), .ZN(n235) );
  XOR2_X1 U198 ( .A(a[3]), .B(a[2]), .Z(n338) );
  XNOR2_X1 U199 ( .A(n214), .B(n236), .ZN(product[11]) );
  XNOR2_X1 U200 ( .A(n23), .B(n20), .ZN(n236) );
  XOR2_X1 U201 ( .A(n34), .B(n39), .Z(n237) );
  XOR2_X1 U202 ( .A(n8), .B(n237), .Z(product[8]) );
  NAND2_X1 U203 ( .A1(n8), .A2(n34), .ZN(n238) );
  NAND2_X1 U204 ( .A1(n8), .A2(n39), .ZN(n239) );
  NAND2_X1 U205 ( .A1(n34), .A2(n39), .ZN(n240) );
  NAND3_X1 U206 ( .A1(n238), .A2(n239), .A3(n240), .ZN(n7) );
  BUF_X1 U207 ( .A(n282), .Z(n241) );
  XOR2_X1 U208 ( .A(n102), .B(n95), .Z(n56) );
  INV_X1 U209 ( .A(n242), .ZN(n55) );
  NAND2_X1 U210 ( .A1(n206), .A2(n95), .ZN(n242) );
  NAND2_X2 U211 ( .A1(n300), .A2(n338), .ZN(n302) );
  NAND2_X1 U212 ( .A1(n2), .A2(n284), .ZN(n243) );
  NAND2_X1 U213 ( .A1(n2), .A2(n15), .ZN(n244) );
  NAND2_X1 U214 ( .A1(n284), .A2(n15), .ZN(n245) );
  XOR2_X1 U215 ( .A(n33), .B(n28), .Z(n246) );
  XOR2_X1 U216 ( .A(n213), .B(n246), .Z(product[9]) );
  NAND2_X1 U217 ( .A1(n7), .A2(n33), .ZN(n247) );
  NAND2_X1 U218 ( .A1(n212), .A2(n28), .ZN(n248) );
  NAND2_X1 U219 ( .A1(n33), .A2(n28), .ZN(n249) );
  NAND3_X1 U220 ( .A1(n248), .A2(n247), .A3(n249), .ZN(n6) );
  NAND3_X1 U221 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n250) );
  XOR2_X1 U222 ( .A(n27), .B(n24), .Z(n252) );
  XOR2_X1 U223 ( .A(n235), .B(n252), .Z(product[10]) );
  NAND2_X1 U224 ( .A1(n234), .A2(n27), .ZN(n253) );
  NAND2_X1 U225 ( .A1(n6), .A2(n24), .ZN(n254) );
  NAND2_X1 U226 ( .A1(n27), .A2(n24), .ZN(n255) );
  NAND3_X1 U227 ( .A1(n253), .A2(n254), .A3(n255), .ZN(n5) );
  NAND3_X1 U228 ( .A1(n265), .A2(n266), .A3(n267), .ZN(n256) );
  NAND3_X1 U229 ( .A1(n265), .A2(n266), .A3(n267), .ZN(n257) );
  NAND3_X1 U230 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n258) );
  XOR2_X1 U231 ( .A(n18), .B(n19), .Z(n259) );
  XOR2_X1 U232 ( .A(n257), .B(n259), .Z(product[12]) );
  NAND2_X1 U233 ( .A1(n256), .A2(n18), .ZN(n260) );
  NAND2_X1 U234 ( .A1(n4), .A2(n19), .ZN(n261) );
  NAND2_X1 U235 ( .A1(n18), .A2(n19), .ZN(n262) );
  NAND3_X1 U236 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n3) );
  AND2_X1 U237 ( .A1(n104), .A2(n72), .ZN(n263) );
  CLKBUF_X1 U238 ( .A(b[1]), .Z(n264) );
  NAND2_X1 U239 ( .A1(n5), .A2(n23), .ZN(n265) );
  NAND2_X1 U240 ( .A1(n250), .A2(n20), .ZN(n266) );
  NAND2_X1 U241 ( .A1(n23), .A2(n20), .ZN(n267) );
  NAND3_X1 U242 ( .A1(n266), .A2(n265), .A3(n267), .ZN(n4) );
  XOR2_X1 U243 ( .A(n17), .B(n283), .Z(n268) );
  XOR2_X1 U244 ( .A(n3), .B(n268), .Z(product[13]) );
  NAND2_X1 U245 ( .A1(n258), .A2(n17), .ZN(n269) );
  NAND2_X1 U246 ( .A1(n258), .A2(n283), .ZN(n270) );
  NAND2_X1 U247 ( .A1(n17), .A2(n283), .ZN(n271) );
  NAND3_X1 U248 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n2) );
  INV_X1 U249 ( .A(n282), .ZN(n272) );
  NAND2_X1 U250 ( .A1(a[4]), .A2(a[3]), .ZN(n274) );
  NAND2_X1 U251 ( .A1(n273), .A2(n291), .ZN(n275) );
  NAND2_X2 U252 ( .A1(n274), .A2(n275), .ZN(n310) );
  INV_X1 U253 ( .A(a[4]), .ZN(n273) );
  NAND2_X2 U254 ( .A1(n310), .A2(n339), .ZN(n312) );
  XNOR2_X1 U255 ( .A(a[2]), .B(a[1]), .ZN(n276) );
  INV_X1 U256 ( .A(n21), .ZN(n286) );
  INV_X1 U257 ( .A(n319), .ZN(n287) );
  INV_X1 U258 ( .A(n330), .ZN(n284) );
  INV_X1 U259 ( .A(n299), .ZN(n292) );
  INV_X1 U260 ( .A(n308), .ZN(n290) );
  INV_X1 U261 ( .A(n31), .ZN(n289) );
  INV_X1 U262 ( .A(b[0]), .ZN(n282) );
  XNOR2_X1 U263 ( .A(a[2]), .B(a[1]), .ZN(n300) );
  INV_X1 U264 ( .A(a[0]), .ZN(n294) );
  INV_X1 U265 ( .A(a[5]), .ZN(n288) );
  INV_X1 U266 ( .A(a[7]), .ZN(n285) );
  XNOR2_X1 U267 ( .A(n263), .B(n277), .ZN(product[2]) );
  XNOR2_X1 U268 ( .A(n103), .B(n96), .ZN(n277) );
  NAND2_X1 U269 ( .A1(n263), .A2(n207), .ZN(n278) );
  NAND2_X1 U270 ( .A1(n14), .A2(n96), .ZN(n279) );
  NAND2_X1 U271 ( .A1(n207), .A2(n96), .ZN(n280) );
  NAND3_X1 U272 ( .A1(n278), .A2(n279), .A3(n280), .ZN(n13) );
  INV_X1 U273 ( .A(a[3]), .ZN(n291) );
  INV_X1 U274 ( .A(a[1]), .ZN(n293) );
  INV_X1 U275 ( .A(n282), .ZN(n281) );
  NOR2_X1 U276 ( .A1(n294), .A2(n241), .ZN(product[0]) );
  OAI22_X1 U277 ( .A1(n295), .A2(n296), .B1(n297), .B2(n294), .ZN(n99) );
  OAI22_X1 U278 ( .A1(n297), .A2(n296), .B1(n298), .B2(n294), .ZN(n98) );
  XNOR2_X1 U279 ( .A(b[6]), .B(a[1]), .ZN(n297) );
  OAI22_X1 U280 ( .A1(n294), .A2(n298), .B1(n296), .B2(n298), .ZN(n299) );
  XNOR2_X1 U281 ( .A(b[7]), .B(a[1]), .ZN(n298) );
  NOR2_X1 U282 ( .A1(n276), .A2(n241), .ZN(n96) );
  OAI22_X1 U283 ( .A1(n301), .A2(n302), .B1(n276), .B2(n303), .ZN(n95) );
  XNOR2_X1 U284 ( .A(a[3]), .B(n281), .ZN(n301) );
  OAI22_X1 U285 ( .A1(n303), .A2(n302), .B1(n276), .B2(n304), .ZN(n94) );
  XNOR2_X1 U286 ( .A(b[1]), .B(a[3]), .ZN(n303) );
  OAI22_X1 U287 ( .A1(n304), .A2(n302), .B1(n276), .B2(n305), .ZN(n93) );
  XNOR2_X1 U288 ( .A(b[2]), .B(a[3]), .ZN(n304) );
  OAI22_X1 U289 ( .A1(n305), .A2(n302), .B1(n276), .B2(n306), .ZN(n92) );
  XNOR2_X1 U290 ( .A(b[3]), .B(a[3]), .ZN(n305) );
  OAI22_X1 U291 ( .A1(n306), .A2(n302), .B1(n276), .B2(n307), .ZN(n91) );
  XNOR2_X1 U292 ( .A(b[4]), .B(a[3]), .ZN(n306) );
  OAI22_X1 U293 ( .A1(n309), .A2(n276), .B1(n302), .B2(n309), .ZN(n308) );
  NOR2_X1 U294 ( .A1(n310), .A2(n241), .ZN(n88) );
  OAI22_X1 U295 ( .A1(n311), .A2(n312), .B1(n310), .B2(n313), .ZN(n87) );
  XNOR2_X1 U296 ( .A(a[5]), .B(n272), .ZN(n311) );
  OAI22_X1 U297 ( .A1(n313), .A2(n312), .B1(n310), .B2(n314), .ZN(n86) );
  XNOR2_X1 U298 ( .A(n264), .B(a[5]), .ZN(n313) );
  OAI22_X1 U299 ( .A1(n314), .A2(n312), .B1(n310), .B2(n315), .ZN(n85) );
  XNOR2_X1 U300 ( .A(b[2]), .B(a[5]), .ZN(n314) );
  OAI22_X1 U301 ( .A1(n315), .A2(n312), .B1(n310), .B2(n316), .ZN(n84) );
  XNOR2_X1 U302 ( .A(b[3]), .B(a[5]), .ZN(n315) );
  OAI22_X1 U303 ( .A1(n316), .A2(n312), .B1(n310), .B2(n317), .ZN(n83) );
  XNOR2_X1 U304 ( .A(b[4]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U305 ( .A1(n317), .A2(n312), .B1(n310), .B2(n318), .ZN(n82) );
  XNOR2_X1 U306 ( .A(b[5]), .B(a[5]), .ZN(n317) );
  OAI22_X1 U307 ( .A1(n320), .A2(n310), .B1(n312), .B2(n320), .ZN(n319) );
  NOR2_X1 U308 ( .A1(n321), .A2(n241), .ZN(n80) );
  OAI22_X1 U309 ( .A1(n322), .A2(n323), .B1(n321), .B2(n324), .ZN(n79) );
  XNOR2_X1 U310 ( .A(a[7]), .B(n272), .ZN(n322) );
  OAI22_X1 U311 ( .A1(n325), .A2(n323), .B1(n321), .B2(n326), .ZN(n77) );
  OAI22_X1 U312 ( .A1(n326), .A2(n323), .B1(n321), .B2(n327), .ZN(n76) );
  XNOR2_X1 U313 ( .A(b[3]), .B(a[7]), .ZN(n326) );
  OAI22_X1 U314 ( .A1(n327), .A2(n323), .B1(n321), .B2(n328), .ZN(n75) );
  XNOR2_X1 U315 ( .A(b[4]), .B(a[7]), .ZN(n327) );
  OAI22_X1 U316 ( .A1(n328), .A2(n323), .B1(n321), .B2(n329), .ZN(n74) );
  XNOR2_X1 U317 ( .A(b[5]), .B(a[7]), .ZN(n328) );
  OAI22_X1 U318 ( .A1(n331), .A2(n321), .B1(n323), .B2(n331), .ZN(n330) );
  OAI21_X1 U319 ( .B1(n281), .B2(n293), .A(n296), .ZN(n72) );
  OAI21_X1 U320 ( .B1(n291), .B2(n302), .A(n332), .ZN(n71) );
  OR3_X1 U321 ( .A1(n276), .A2(n272), .A3(n291), .ZN(n332) );
  OAI21_X1 U322 ( .B1(n288), .B2(n312), .A(n333), .ZN(n70) );
  OR3_X1 U323 ( .A1(n310), .A2(n272), .A3(n288), .ZN(n333) );
  OAI21_X1 U324 ( .B1(n285), .B2(n323), .A(n334), .ZN(n69) );
  OR3_X1 U325 ( .A1(n321), .A2(n272), .A3(n285), .ZN(n334) );
  XNOR2_X1 U326 ( .A(n335), .B(n336), .ZN(n38) );
  OR2_X1 U327 ( .A1(n335), .A2(n336), .ZN(n37) );
  OAI22_X1 U328 ( .A1(n307), .A2(n302), .B1(n276), .B2(n337), .ZN(n336) );
  XNOR2_X1 U329 ( .A(b[5]), .B(a[3]), .ZN(n307) );
  OAI22_X1 U330 ( .A1(n324), .A2(n323), .B1(n321), .B2(n325), .ZN(n335) );
  XNOR2_X1 U331 ( .A(b[2]), .B(a[7]), .ZN(n325) );
  XNOR2_X1 U332 ( .A(n264), .B(a[7]), .ZN(n324) );
  OAI22_X1 U333 ( .A1(n337), .A2(n302), .B1(n276), .B2(n309), .ZN(n31) );
  XNOR2_X1 U334 ( .A(b[7]), .B(a[3]), .ZN(n309) );
  XNOR2_X1 U335 ( .A(b[6]), .B(a[3]), .ZN(n337) );
  OAI22_X1 U336 ( .A1(n318), .A2(n312), .B1(n310), .B2(n320), .ZN(n21) );
  XNOR2_X1 U337 ( .A(b[7]), .B(a[5]), .ZN(n320) );
  XNOR2_X1 U338 ( .A(n288), .B(a[4]), .ZN(n339) );
  XNOR2_X1 U339 ( .A(b[6]), .B(a[5]), .ZN(n318) );
  OAI22_X1 U340 ( .A1(n329), .A2(n323), .B1(n321), .B2(n331), .ZN(n15) );
  XNOR2_X1 U341 ( .A(b[7]), .B(a[7]), .ZN(n331) );
  NAND2_X1 U342 ( .A1(n321), .A2(n340), .ZN(n323) );
  XNOR2_X1 U343 ( .A(n285), .B(a[6]), .ZN(n340) );
  XNOR2_X1 U344 ( .A(b[6]), .B(a[7]), .ZN(n329) );
  OAI22_X1 U345 ( .A1(n281), .A2(n296), .B1(n341), .B2(n294), .ZN(n104) );
  OAI22_X1 U346 ( .A1(n251), .A2(n296), .B1(n342), .B2(n294), .ZN(n103) );
  XNOR2_X1 U347 ( .A(b[1]), .B(a[1]), .ZN(n341) );
  OAI22_X1 U348 ( .A1(n342), .A2(n296), .B1(n343), .B2(n294), .ZN(n102) );
  XNOR2_X1 U349 ( .A(b[2]), .B(a[1]), .ZN(n342) );
  OAI22_X1 U350 ( .A1(n343), .A2(n296), .B1(n344), .B2(n294), .ZN(n101) );
  XNOR2_X1 U351 ( .A(b[3]), .B(a[1]), .ZN(n343) );
  OAI22_X1 U352 ( .A1(n344), .A2(n296), .B1(n295), .B2(n294), .ZN(n100) );
  XNOR2_X1 U353 ( .A(b[5]), .B(a[1]), .ZN(n295) );
  NAND2_X1 U354 ( .A1(a[1]), .A2(n294), .ZN(n296) );
  XNOR2_X1 U355 ( .A(b[4]), .B(a[1]), .ZN(n344) );
endmodule


module datapath_DW01_add_3 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n72;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  NAND3_X1 U1 ( .A1(n13), .A2(n14), .A3(n15), .ZN(n1) );
  CLKBUF_X1 U2 ( .A(B[1]), .Z(n2) );
  CLKBUF_X1 U3 ( .A(carry[12]), .Z(n3) );
  NAND3_X1 U4 ( .A1(n41), .A2(n43), .A3(n42), .ZN(n4) );
  NAND3_X1 U5 ( .A1(n41), .A2(n43), .A3(n42), .ZN(n5) );
  NAND3_X1 U6 ( .A1(n33), .A2(n34), .A3(n35), .ZN(n6) );
  CLKBUF_X1 U7 ( .A(carry[10]), .Z(n7) );
  XOR2_X1 U8 ( .A(n5), .B(A[11]), .Z(n8) );
  XOR2_X1 U9 ( .A(B[11]), .B(n8), .Z(SUM[11]) );
  NAND2_X1 U10 ( .A1(B[11]), .A2(n4), .ZN(n9) );
  NAND2_X1 U11 ( .A1(B[11]), .A2(A[11]), .ZN(n10) );
  NAND2_X1 U12 ( .A1(carry[11]), .A2(A[11]), .ZN(n11) );
  NAND3_X1 U13 ( .A1(n9), .A2(n10), .A3(n11), .ZN(carry[12]) );
  XOR2_X1 U14 ( .A(n72), .B(A[1]), .Z(n12) );
  XOR2_X1 U15 ( .A(n2), .B(n12), .Z(SUM[1]) );
  NAND2_X1 U16 ( .A1(B[1]), .A2(n72), .ZN(n13) );
  NAND2_X1 U17 ( .A1(B[1]), .A2(A[1]), .ZN(n14) );
  NAND2_X1 U18 ( .A1(n72), .A2(A[1]), .ZN(n15) );
  NAND3_X1 U19 ( .A1(n13), .A2(n14), .A3(n15), .ZN(carry[2]) );
  NAND3_X1 U20 ( .A1(n49), .A2(n50), .A3(n51), .ZN(n16) );
  NAND3_X1 U21 ( .A1(n69), .A2(n68), .A3(n70), .ZN(n17) );
  NAND3_X1 U22 ( .A1(n46), .A2(n45), .A3(n47), .ZN(n18) );
  NAND3_X1 U23 ( .A1(n25), .A2(n26), .A3(n27), .ZN(n19) );
  NAND3_X1 U24 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n20) );
  NAND3_X1 U25 ( .A1(n37), .A2(n38), .A3(n39), .ZN(n21) );
  NAND3_X1 U26 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n22) );
  NAND3_X1 U27 ( .A1(n29), .A2(n30), .A3(n31), .ZN(n23) );
  XOR2_X1 U28 ( .A(n21), .B(A[5]), .Z(n24) );
  XOR2_X1 U29 ( .A(B[5]), .B(n24), .Z(SUM[5]) );
  NAND2_X1 U30 ( .A1(B[5]), .A2(n20), .ZN(n25) );
  NAND2_X1 U31 ( .A1(B[5]), .A2(A[5]), .ZN(n26) );
  NAND2_X1 U32 ( .A1(carry[5]), .A2(A[5]), .ZN(n27) );
  NAND3_X1 U33 ( .A1(n25), .A2(n26), .A3(n27), .ZN(carry[6]) );
  XOR2_X1 U34 ( .A(A[2]), .B(B[2]), .Z(n28) );
  XOR2_X1 U35 ( .A(n28), .B(n1), .Z(SUM[2]) );
  NAND2_X1 U36 ( .A1(A[2]), .A2(B[2]), .ZN(n29) );
  NAND2_X1 U37 ( .A1(A[2]), .A2(carry[2]), .ZN(n30) );
  NAND2_X1 U38 ( .A1(n1), .A2(B[2]), .ZN(n31) );
  NAND3_X1 U39 ( .A1(n29), .A2(n30), .A3(n31), .ZN(carry[3]) );
  XOR2_X1 U40 ( .A(B[3]), .B(A[3]), .Z(n32) );
  XOR2_X1 U41 ( .A(n32), .B(n23), .Z(SUM[3]) );
  NAND2_X1 U42 ( .A1(B[3]), .A2(A[3]), .ZN(n33) );
  NAND2_X1 U43 ( .A1(B[3]), .A2(n22), .ZN(n34) );
  NAND2_X1 U44 ( .A1(A[3]), .A2(carry[3]), .ZN(n35) );
  NAND3_X1 U45 ( .A1(n33), .A2(n34), .A3(n35), .ZN(carry[4]) );
  XOR2_X1 U46 ( .A(B[4]), .B(A[4]), .Z(n36) );
  XOR2_X1 U47 ( .A(carry[4]), .B(n36), .Z(SUM[4]) );
  NAND2_X1 U48 ( .A1(n6), .A2(B[4]), .ZN(n37) );
  NAND2_X1 U49 ( .A1(carry[4]), .A2(A[4]), .ZN(n38) );
  NAND2_X1 U50 ( .A1(B[4]), .A2(A[4]), .ZN(n39) );
  NAND3_X1 U51 ( .A1(n37), .A2(n38), .A3(n39), .ZN(carry[5]) );
  XOR2_X1 U52 ( .A(B[10]), .B(A[10]), .Z(n40) );
  XOR2_X1 U53 ( .A(n7), .B(n40), .Z(SUM[10]) );
  NAND2_X1 U54 ( .A1(carry[10]), .A2(B[10]), .ZN(n41) );
  NAND2_X1 U55 ( .A1(n17), .A2(A[10]), .ZN(n42) );
  NAND2_X1 U56 ( .A1(B[10]), .A2(A[10]), .ZN(n43) );
  NAND3_X1 U57 ( .A1(n41), .A2(n43), .A3(n42), .ZN(carry[11]) );
  XOR2_X1 U58 ( .A(B[6]), .B(A[6]), .Z(n44) );
  XOR2_X1 U59 ( .A(carry[6]), .B(n44), .Z(SUM[6]) );
  NAND2_X1 U60 ( .A1(n19), .A2(B[6]), .ZN(n45) );
  NAND2_X1 U61 ( .A1(n19), .A2(A[6]), .ZN(n46) );
  NAND2_X1 U62 ( .A1(B[6]), .A2(A[6]), .ZN(n47) );
  NAND3_X1 U63 ( .A1(n45), .A2(n46), .A3(n47), .ZN(carry[7]) );
  XOR2_X1 U64 ( .A(B[12]), .B(A[12]), .Z(n48) );
  XOR2_X1 U65 ( .A(n3), .B(n48), .Z(SUM[12]) );
  NAND2_X1 U66 ( .A1(carry[12]), .A2(B[12]), .ZN(n49) );
  NAND2_X1 U67 ( .A1(carry[12]), .A2(A[12]), .ZN(n50) );
  NAND2_X1 U68 ( .A1(B[12]), .A2(A[12]), .ZN(n51) );
  NAND3_X1 U69 ( .A1(n50), .A2(n49), .A3(n51), .ZN(carry[13]) );
  NAND3_X1 U70 ( .A1(n63), .A2(n64), .A3(n65), .ZN(n52) );
  NAND3_X1 U71 ( .A1(n59), .A2(n60), .A3(n61), .ZN(n53) );
  XOR2_X1 U72 ( .A(B[13]), .B(A[13]), .Z(n54) );
  XOR2_X1 U73 ( .A(n16), .B(n54), .Z(SUM[13]) );
  NAND2_X1 U74 ( .A1(n16), .A2(B[13]), .ZN(n55) );
  NAND2_X1 U75 ( .A1(carry[13]), .A2(A[13]), .ZN(n56) );
  NAND2_X1 U76 ( .A1(B[13]), .A2(A[13]), .ZN(n57) );
  NAND3_X1 U77 ( .A1(n55), .A2(n56), .A3(n57), .ZN(carry[14]) );
  XOR2_X1 U78 ( .A(B[7]), .B(A[7]), .Z(n58) );
  XOR2_X1 U79 ( .A(carry[7]), .B(n58), .Z(SUM[7]) );
  NAND2_X1 U80 ( .A1(carry[7]), .A2(B[7]), .ZN(n59) );
  NAND2_X1 U81 ( .A1(n18), .A2(A[7]), .ZN(n60) );
  NAND2_X1 U82 ( .A1(B[7]), .A2(A[7]), .ZN(n61) );
  NAND3_X1 U83 ( .A1(n59), .A2(n60), .A3(n61), .ZN(carry[8]) );
  XOR2_X1 U84 ( .A(B[8]), .B(A[8]), .Z(n62) );
  XOR2_X1 U85 ( .A(carry[8]), .B(n62), .Z(SUM[8]) );
  NAND2_X1 U86 ( .A1(n53), .A2(B[8]), .ZN(n63) );
  NAND2_X1 U87 ( .A1(n53), .A2(A[8]), .ZN(n64) );
  NAND2_X1 U88 ( .A1(B[8]), .A2(A[8]), .ZN(n65) );
  NAND3_X1 U89 ( .A1(n63), .A2(n64), .A3(n65), .ZN(carry[9]) );
  XNOR2_X1 U90 ( .A(carry[15]), .B(n66), .ZN(SUM[15]) );
  XNOR2_X1 U91 ( .A(B[15]), .B(A[15]), .ZN(n66) );
  XOR2_X1 U92 ( .A(B[9]), .B(A[9]), .Z(n67) );
  XOR2_X1 U93 ( .A(carry[9]), .B(n67), .Z(SUM[9]) );
  NAND2_X1 U94 ( .A1(n52), .A2(B[9]), .ZN(n68) );
  NAND2_X1 U95 ( .A1(n52), .A2(A[9]), .ZN(n69) );
  NAND2_X1 U96 ( .A1(B[9]), .A2(A[9]), .ZN(n70) );
  NAND3_X1 U97 ( .A1(n68), .A2(n69), .A3(n70), .ZN(carry[10]) );
  XOR2_X1 U98 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U99 ( .A1(B[0]), .A2(A[0]), .ZN(n72) );
endmodule


module datapath_DW_mult_tc_2 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74,
         n75, n76, n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92,
         n93, n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n206,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329;

  FA_X1 U10 ( .A(n46), .B(n49), .CI(n10), .CO(n9), .S(product[6]) );
  FA_X1 U13 ( .A(n13), .B(n71), .CI(n56), .CO(n12), .S(product[3]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n272), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n271), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n275), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n274), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n277), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n87), .B(n70), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n94), .B(n88), .CI(n101), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n95), .B(n102), .CO(n55), .S(n56) );
  XNOR2_X1 U157 ( .A(n269), .B(n15), .ZN(n206) );
  AND3_X1 U158 ( .A1(n240), .A2(n241), .A3(n242), .ZN(product[15]) );
  CLKBUF_X1 U159 ( .A(n287), .Z(n208) );
  INV_X2 U160 ( .A(a[0]), .ZN(n279) );
  XNOR2_X1 U161 ( .A(a[2]), .B(a[1]), .ZN(n261) );
  CLKBUF_X1 U162 ( .A(b[1]), .Z(n209) );
  CLKBUF_X1 U163 ( .A(n326), .Z(n217) );
  XOR2_X1 U164 ( .A(n27), .B(n24), .Z(n210) );
  XOR2_X1 U165 ( .A(n6), .B(n210), .Z(product[10]) );
  NAND2_X1 U166 ( .A1(n6), .A2(n27), .ZN(n211) );
  NAND2_X1 U167 ( .A1(n6), .A2(n24), .ZN(n212) );
  NAND2_X1 U168 ( .A1(n27), .A2(n24), .ZN(n213) );
  NAND3_X1 U169 ( .A1(n211), .A2(n212), .A3(n213), .ZN(n5) );
  NAND3_X1 U170 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n214) );
  NAND3_X1 U171 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n215) );
  NAND3_X1 U172 ( .A1(n233), .A2(n234), .A3(n235), .ZN(n216) );
  XNOR2_X1 U173 ( .A(n12), .B(n218), .ZN(product[4]) );
  XNOR2_X1 U174 ( .A(n54), .B(n55), .ZN(n218) );
  XOR2_X2 U175 ( .A(a[6]), .B(n273), .Z(n306) );
  NAND2_X1 U176 ( .A1(n12), .A2(n54), .ZN(n219) );
  NAND2_X1 U177 ( .A1(n12), .A2(n55), .ZN(n220) );
  NAND2_X1 U178 ( .A1(n54), .A2(n55), .ZN(n221) );
  NAND3_X1 U179 ( .A1(n219), .A2(n220), .A3(n221), .ZN(n11) );
  XOR2_X1 U180 ( .A(n50), .B(n53), .Z(n222) );
  XOR2_X1 U181 ( .A(n11), .B(n222), .Z(product[5]) );
  NAND2_X1 U182 ( .A1(n11), .A2(n50), .ZN(n223) );
  NAND2_X1 U183 ( .A1(n11), .A2(n53), .ZN(n224) );
  NAND2_X1 U184 ( .A1(n50), .A2(n53), .ZN(n225) );
  NAND3_X1 U185 ( .A1(n223), .A2(n224), .A3(n225), .ZN(n10) );
  XOR2_X1 U186 ( .A(n40), .B(n45), .Z(n226) );
  XOR2_X1 U187 ( .A(n9), .B(n226), .Z(product[7]) );
  NAND2_X1 U188 ( .A1(n9), .A2(n40), .ZN(n227) );
  NAND2_X1 U189 ( .A1(n9), .A2(n45), .ZN(n228) );
  NAND2_X1 U190 ( .A1(n40), .A2(n45), .ZN(n229) );
  NAND3_X1 U191 ( .A1(n227), .A2(n228), .A3(n229), .ZN(n8) );
  XNOR2_X1 U192 ( .A(n215), .B(n206), .ZN(product[14]) );
  XNOR2_X1 U193 ( .A(b[2]), .B(a[1]), .ZN(n230) );
  BUF_X1 U194 ( .A(n267), .Z(n231) );
  NAND2_X1 U195 ( .A1(n285), .A2(n323), .ZN(n287) );
  XOR2_X1 U196 ( .A(n34), .B(n39), .Z(n232) );
  XOR2_X1 U197 ( .A(n232), .B(n8), .Z(product[8]) );
  NAND2_X1 U198 ( .A1(n34), .A2(n39), .ZN(n233) );
  NAND2_X1 U199 ( .A1(n34), .A2(n8), .ZN(n234) );
  NAND2_X1 U200 ( .A1(n39), .A2(n8), .ZN(n235) );
  NAND3_X1 U201 ( .A1(n235), .A2(n234), .A3(n233), .ZN(n7) );
  XOR2_X1 U202 ( .A(n28), .B(n33), .Z(n236) );
  XOR2_X1 U203 ( .A(n236), .B(n7), .Z(product[9]) );
  NAND2_X1 U204 ( .A1(n28), .A2(n33), .ZN(n237) );
  NAND2_X1 U205 ( .A1(n28), .A2(n216), .ZN(n238) );
  NAND2_X1 U206 ( .A1(n33), .A2(n7), .ZN(n239) );
  NAND3_X1 U207 ( .A1(n237), .A2(n238), .A3(n239), .ZN(n6) );
  NAND2_X1 U208 ( .A1(n214), .A2(n269), .ZN(n240) );
  NAND2_X1 U209 ( .A1(n2), .A2(n15), .ZN(n241) );
  NAND2_X1 U210 ( .A1(n269), .A2(n15), .ZN(n242) );
  XOR2_X1 U211 ( .A(n23), .B(n20), .Z(n243) );
  XOR2_X1 U212 ( .A(n5), .B(n243), .Z(product[11]) );
  NAND2_X1 U213 ( .A1(n5), .A2(n23), .ZN(n244) );
  NAND2_X1 U214 ( .A1(n5), .A2(n20), .ZN(n245) );
  NAND2_X1 U215 ( .A1(n23), .A2(n20), .ZN(n246) );
  NAND3_X1 U216 ( .A1(n244), .A2(n245), .A3(n246), .ZN(n4) );
  INV_X1 U217 ( .A(n267), .ZN(n247) );
  INV_X1 U218 ( .A(n267), .ZN(n266) );
  XOR2_X1 U219 ( .A(n18), .B(n19), .Z(n248) );
  XOR2_X1 U220 ( .A(n4), .B(n248), .Z(product[12]) );
  NAND2_X1 U221 ( .A1(n4), .A2(n18), .ZN(n249) );
  NAND2_X1 U222 ( .A1(n4), .A2(n19), .ZN(n250) );
  NAND2_X1 U223 ( .A1(n18), .A2(n19), .ZN(n251) );
  NAND3_X1 U224 ( .A1(n249), .A2(n250), .A3(n251), .ZN(n3) );
  AND2_X1 U225 ( .A1(n104), .A2(n72), .ZN(n252) );
  XOR2_X1 U226 ( .A(n17), .B(n268), .Z(n253) );
  XOR2_X1 U227 ( .A(n3), .B(n253), .Z(product[13]) );
  NAND2_X1 U228 ( .A1(n3), .A2(n17), .ZN(n254) );
  NAND2_X1 U229 ( .A1(n3), .A2(n268), .ZN(n255) );
  NAND2_X1 U230 ( .A1(n17), .A2(n268), .ZN(n256) );
  NAND3_X1 U231 ( .A1(n254), .A2(n255), .A3(n256), .ZN(n2) );
  NAND2_X1 U232 ( .A1(a[4]), .A2(a[3]), .ZN(n259) );
  NAND2_X1 U233 ( .A1(n257), .A2(n258), .ZN(n260) );
  NAND2_X2 U234 ( .A1(n259), .A2(n260), .ZN(n295) );
  INV_X1 U235 ( .A(a[4]), .ZN(n257) );
  INV_X1 U236 ( .A(a[3]), .ZN(n258) );
  NAND2_X2 U237 ( .A1(n295), .A2(n324), .ZN(n297) );
  INV_X1 U238 ( .A(n15), .ZN(n268) );
  INV_X1 U239 ( .A(n21), .ZN(n271) );
  INV_X1 U240 ( .A(n304), .ZN(n272) );
  INV_X1 U241 ( .A(n315), .ZN(n269) );
  INV_X1 U242 ( .A(n284), .ZN(n277) );
  INV_X1 U243 ( .A(n293), .ZN(n275) );
  INV_X1 U244 ( .A(n31), .ZN(n274) );
  INV_X1 U245 ( .A(b[0]), .ZN(n267) );
  XNOR2_X1 U246 ( .A(a[2]), .B(a[1]), .ZN(n285) );
  INV_X1 U247 ( .A(a[5]), .ZN(n273) );
  INV_X1 U248 ( .A(a[7]), .ZN(n270) );
  XNOR2_X1 U249 ( .A(n262), .B(n252), .ZN(product[2]) );
  XNOR2_X1 U250 ( .A(n103), .B(n96), .ZN(n262) );
  NAND2_X1 U251 ( .A1(n252), .A2(n103), .ZN(n263) );
  NAND2_X1 U252 ( .A1(n14), .A2(n96), .ZN(n264) );
  NAND2_X1 U253 ( .A1(n103), .A2(n96), .ZN(n265) );
  NAND3_X1 U254 ( .A1(n263), .A2(n264), .A3(n265), .ZN(n13) );
  INV_X1 U255 ( .A(a[3]), .ZN(n276) );
  INV_X1 U256 ( .A(a[1]), .ZN(n278) );
  NOR2_X1 U257 ( .A1(n279), .A2(n231), .ZN(product[0]) );
  OAI22_X1 U258 ( .A1(n280), .A2(n281), .B1(n282), .B2(n279), .ZN(n99) );
  OAI22_X1 U259 ( .A1(n282), .A2(n281), .B1(n283), .B2(n279), .ZN(n98) );
  XNOR2_X1 U260 ( .A(b[6]), .B(a[1]), .ZN(n282) );
  OAI22_X1 U261 ( .A1(n279), .A2(n283), .B1(n281), .B2(n283), .ZN(n284) );
  XNOR2_X1 U262 ( .A(b[7]), .B(a[1]), .ZN(n283) );
  NOR2_X1 U263 ( .A1(n261), .A2(n231), .ZN(n96) );
  OAI22_X1 U264 ( .A1(n286), .A2(n287), .B1(n261), .B2(n288), .ZN(n95) );
  XNOR2_X1 U265 ( .A(a[3]), .B(n266), .ZN(n286) );
  OAI22_X1 U266 ( .A1(n288), .A2(n287), .B1(n261), .B2(n289), .ZN(n94) );
  XNOR2_X1 U267 ( .A(b[1]), .B(a[3]), .ZN(n288) );
  OAI22_X1 U268 ( .A1(n289), .A2(n287), .B1(n261), .B2(n290), .ZN(n93) );
  XNOR2_X1 U269 ( .A(b[2]), .B(a[3]), .ZN(n289) );
  OAI22_X1 U270 ( .A1(n290), .A2(n287), .B1(n261), .B2(n291), .ZN(n92) );
  XNOR2_X1 U271 ( .A(b[3]), .B(a[3]), .ZN(n290) );
  OAI22_X1 U272 ( .A1(n291), .A2(n208), .B1(n261), .B2(n292), .ZN(n91) );
  XNOR2_X1 U273 ( .A(b[4]), .B(a[3]), .ZN(n291) );
  OAI22_X1 U274 ( .A1(n294), .A2(n261), .B1(n208), .B2(n294), .ZN(n293) );
  NOR2_X1 U275 ( .A1(n295), .A2(n231), .ZN(n88) );
  OAI22_X1 U276 ( .A1(n296), .A2(n297), .B1(n295), .B2(n298), .ZN(n87) );
  XNOR2_X1 U277 ( .A(a[5]), .B(n247), .ZN(n296) );
  OAI22_X1 U278 ( .A1(n298), .A2(n297), .B1(n295), .B2(n299), .ZN(n86) );
  XNOR2_X1 U279 ( .A(n209), .B(a[5]), .ZN(n298) );
  OAI22_X1 U280 ( .A1(n299), .A2(n297), .B1(n295), .B2(n300), .ZN(n85) );
  XNOR2_X1 U281 ( .A(b[2]), .B(a[5]), .ZN(n299) );
  OAI22_X1 U282 ( .A1(n300), .A2(n297), .B1(n295), .B2(n301), .ZN(n84) );
  XNOR2_X1 U283 ( .A(b[3]), .B(a[5]), .ZN(n300) );
  OAI22_X1 U284 ( .A1(n301), .A2(n297), .B1(n295), .B2(n302), .ZN(n83) );
  XNOR2_X1 U285 ( .A(b[4]), .B(a[5]), .ZN(n301) );
  OAI22_X1 U286 ( .A1(n302), .A2(n297), .B1(n295), .B2(n303), .ZN(n82) );
  XNOR2_X1 U287 ( .A(b[5]), .B(a[5]), .ZN(n302) );
  OAI22_X1 U288 ( .A1(n305), .A2(n295), .B1(n297), .B2(n305), .ZN(n304) );
  NOR2_X1 U289 ( .A1(n306), .A2(n231), .ZN(n80) );
  OAI22_X1 U290 ( .A1(n307), .A2(n308), .B1(n306), .B2(n309), .ZN(n79) );
  XNOR2_X1 U291 ( .A(a[7]), .B(n247), .ZN(n307) );
  OAI22_X1 U292 ( .A1(n310), .A2(n308), .B1(n306), .B2(n311), .ZN(n77) );
  OAI22_X1 U293 ( .A1(n311), .A2(n308), .B1(n306), .B2(n312), .ZN(n76) );
  XNOR2_X1 U294 ( .A(b[3]), .B(a[7]), .ZN(n311) );
  OAI22_X1 U295 ( .A1(n312), .A2(n308), .B1(n306), .B2(n313), .ZN(n75) );
  XNOR2_X1 U296 ( .A(b[4]), .B(a[7]), .ZN(n312) );
  OAI22_X1 U297 ( .A1(n313), .A2(n308), .B1(n306), .B2(n314), .ZN(n74) );
  XNOR2_X1 U298 ( .A(b[5]), .B(a[7]), .ZN(n313) );
  OAI22_X1 U299 ( .A1(n316), .A2(n306), .B1(n308), .B2(n316), .ZN(n315) );
  OAI21_X1 U300 ( .B1(n266), .B2(n278), .A(n281), .ZN(n72) );
  OAI21_X1 U301 ( .B1(n276), .B2(n287), .A(n317), .ZN(n71) );
  OR3_X1 U302 ( .A1(n261), .A2(n247), .A3(n276), .ZN(n317) );
  OAI21_X1 U303 ( .B1(n273), .B2(n297), .A(n318), .ZN(n70) );
  OR3_X1 U304 ( .A1(n295), .A2(n247), .A3(n273), .ZN(n318) );
  OAI21_X1 U305 ( .B1(n270), .B2(n308), .A(n319), .ZN(n69) );
  OR3_X1 U306 ( .A1(n306), .A2(n247), .A3(n270), .ZN(n319) );
  XNOR2_X1 U307 ( .A(n320), .B(n321), .ZN(n38) );
  OR2_X1 U308 ( .A1(n320), .A2(n321), .ZN(n37) );
  OAI22_X1 U309 ( .A1(n292), .A2(n208), .B1(n261), .B2(n322), .ZN(n321) );
  XNOR2_X1 U310 ( .A(b[5]), .B(a[3]), .ZN(n292) );
  OAI22_X1 U311 ( .A1(n309), .A2(n308), .B1(n306), .B2(n310), .ZN(n320) );
  XNOR2_X1 U312 ( .A(b[2]), .B(a[7]), .ZN(n310) );
  XNOR2_X1 U313 ( .A(n209), .B(a[7]), .ZN(n309) );
  OAI22_X1 U314 ( .A1(n322), .A2(n208), .B1(n261), .B2(n294), .ZN(n31) );
  XNOR2_X1 U315 ( .A(b[7]), .B(a[3]), .ZN(n294) );
  XNOR2_X1 U316 ( .A(n276), .B(a[2]), .ZN(n323) );
  XNOR2_X1 U317 ( .A(b[6]), .B(a[3]), .ZN(n322) );
  OAI22_X1 U318 ( .A1(n303), .A2(n297), .B1(n295), .B2(n305), .ZN(n21) );
  XNOR2_X1 U319 ( .A(b[7]), .B(a[5]), .ZN(n305) );
  XNOR2_X1 U320 ( .A(n273), .B(a[4]), .ZN(n324) );
  XNOR2_X1 U321 ( .A(b[6]), .B(a[5]), .ZN(n303) );
  OAI22_X1 U322 ( .A1(n314), .A2(n308), .B1(n306), .B2(n316), .ZN(n15) );
  XNOR2_X1 U323 ( .A(b[7]), .B(a[7]), .ZN(n316) );
  NAND2_X1 U324 ( .A1(n306), .A2(n325), .ZN(n308) );
  XNOR2_X1 U325 ( .A(n270), .B(a[6]), .ZN(n325) );
  XNOR2_X1 U326 ( .A(b[6]), .B(a[7]), .ZN(n314) );
  OAI22_X1 U327 ( .A1(n266), .A2(n281), .B1(n326), .B2(n279), .ZN(n104) );
  OAI22_X1 U328 ( .A1(n217), .A2(n281), .B1(n327), .B2(n279), .ZN(n103) );
  XNOR2_X1 U329 ( .A(b[1]), .B(a[1]), .ZN(n326) );
  OAI22_X1 U330 ( .A1(n281), .A2(n230), .B1(n328), .B2(n279), .ZN(n102) );
  XNOR2_X1 U331 ( .A(b[2]), .B(a[1]), .ZN(n327) );
  OAI22_X1 U332 ( .A1(n328), .A2(n281), .B1(n329), .B2(n279), .ZN(n101) );
  XNOR2_X1 U333 ( .A(b[3]), .B(a[1]), .ZN(n328) );
  OAI22_X1 U334 ( .A1(n329), .A2(n281), .B1(n280), .B2(n279), .ZN(n100) );
  XNOR2_X1 U335 ( .A(b[5]), .B(a[1]), .ZN(n280) );
  NAND2_X1 U336 ( .A1(a[1]), .A2(n279), .ZN(n281) );
  XNOR2_X1 U337 ( .A(b[4]), .B(a[1]), .ZN(n329) );
endmodule


module datapath_DW01_add_2 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n62;
  wire   [15:1] carry;

  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(B[2]), .B(A[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(n62), .CI(B[1]), .CO(carry[2]), .S(SUM[1]) );
  INV_X1 U1 ( .A(A[14]), .ZN(n48) );
  CLKBUF_X1 U2 ( .A(n33), .Z(n1) );
  CLKBUF_X1 U3 ( .A(n29), .Z(n2) );
  NAND3_X1 U4 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n3) );
  NAND3_X1 U5 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n4) );
  NAND3_X1 U6 ( .A1(n19), .A2(n20), .A3(n21), .ZN(n5) );
  NAND3_X1 U7 ( .A1(n28), .A2(n2), .A3(n30), .ZN(n6) );
  XOR2_X1 U8 ( .A(B[4]), .B(A[4]), .Z(n7) );
  XOR2_X1 U9 ( .A(carry[4]), .B(n7), .Z(SUM[4]) );
  NAND2_X1 U10 ( .A1(carry[4]), .A2(B[4]), .ZN(n8) );
  NAND2_X1 U11 ( .A1(carry[4]), .A2(A[4]), .ZN(n9) );
  NAND2_X1 U12 ( .A1(B[4]), .A2(A[4]), .ZN(n10) );
  NAND3_X1 U13 ( .A1(n8), .A2(n9), .A3(n10), .ZN(carry[5]) );
  XOR2_X1 U14 ( .A(n4), .B(A[8]), .Z(n11) );
  XOR2_X1 U15 ( .A(B[8]), .B(n11), .Z(SUM[8]) );
  NAND2_X1 U16 ( .A1(n3), .A2(B[8]), .ZN(n12) );
  NAND2_X1 U17 ( .A1(B[8]), .A2(A[8]), .ZN(n13) );
  NAND2_X1 U18 ( .A1(carry[8]), .A2(A[8]), .ZN(n14) );
  NAND3_X1 U19 ( .A1(n12), .A2(n13), .A3(n14), .ZN(carry[9]) );
  NAND3_X1 U20 ( .A1(n19), .A2(n20), .A3(n21), .ZN(n15) );
  NAND3_X1 U21 ( .A1(n32), .A2(n33), .A3(n34), .ZN(n16) );
  NAND3_X1 U22 ( .A1(n36), .A2(n37), .A3(n38), .ZN(n17) );
  XOR2_X1 U23 ( .A(carry[11]), .B(A[11]), .Z(n18) );
  XOR2_X1 U24 ( .A(B[11]), .B(n18), .Z(SUM[11]) );
  NAND2_X1 U25 ( .A1(n17), .A2(B[11]), .ZN(n19) );
  NAND2_X1 U26 ( .A1(B[11]), .A2(A[11]), .ZN(n20) );
  NAND2_X1 U27 ( .A1(n17), .A2(A[11]), .ZN(n21) );
  NAND3_X1 U28 ( .A1(n19), .A2(n20), .A3(n21), .ZN(carry[12]) );
  NAND3_X1 U29 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n22) );
  NAND3_X1 U30 ( .A1(n45), .A2(n46), .A3(n47), .ZN(n23) );
  NAND3_X1 U31 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n24) );
  NAND3_X1 U32 ( .A1(n50), .A2(n51), .A3(n52), .ZN(n25) );
  NAND3_X1 U33 ( .A1(n41), .A2(n40), .A3(n42), .ZN(n26) );
  XOR2_X1 U34 ( .A(B[9]), .B(A[9]), .Z(n27) );
  XOR2_X1 U35 ( .A(carry[9]), .B(n27), .Z(SUM[9]) );
  NAND2_X1 U36 ( .A1(carry[9]), .A2(B[9]), .ZN(n28) );
  NAND2_X1 U37 ( .A1(carry[9]), .A2(A[9]), .ZN(n29) );
  NAND2_X1 U38 ( .A1(B[9]), .A2(A[9]), .ZN(n30) );
  NAND3_X1 U39 ( .A1(n28), .A2(n29), .A3(n30), .ZN(carry[10]) );
  XOR2_X1 U40 ( .A(B[5]), .B(A[5]), .Z(n31) );
  XOR2_X1 U41 ( .A(carry[5]), .B(n31), .Z(SUM[5]) );
  NAND2_X1 U42 ( .A1(carry[5]), .A2(B[5]), .ZN(n32) );
  NAND2_X1 U43 ( .A1(carry[5]), .A2(A[5]), .ZN(n33) );
  NAND2_X1 U44 ( .A1(B[5]), .A2(A[5]), .ZN(n34) );
  NAND3_X1 U45 ( .A1(n32), .A2(n1), .A3(n34), .ZN(carry[6]) );
  XOR2_X1 U46 ( .A(B[10]), .B(A[10]), .Z(n35) );
  XOR2_X1 U47 ( .A(n6), .B(n35), .Z(SUM[10]) );
  NAND2_X1 U48 ( .A1(carry[10]), .A2(B[10]), .ZN(n36) );
  NAND2_X1 U49 ( .A1(n24), .A2(A[10]), .ZN(n37) );
  NAND2_X1 U50 ( .A1(B[10]), .A2(A[10]), .ZN(n38) );
  NAND3_X1 U51 ( .A1(n36), .A2(n37), .A3(n38), .ZN(carry[11]) );
  XOR2_X1 U52 ( .A(B[13]), .B(A[13]), .Z(n39) );
  XOR2_X1 U53 ( .A(n23), .B(n39), .Z(SUM[13]) );
  NAND2_X1 U54 ( .A1(n22), .A2(B[13]), .ZN(n40) );
  NAND2_X1 U55 ( .A1(carry[13]), .A2(A[13]), .ZN(n41) );
  NAND2_X1 U56 ( .A1(B[13]), .A2(A[13]), .ZN(n42) );
  NAND3_X1 U57 ( .A1(n40), .A2(n41), .A3(n42), .ZN(carry[14]) );
  XNOR2_X1 U58 ( .A(carry[15]), .B(n43), .ZN(SUM[15]) );
  XNOR2_X1 U59 ( .A(B[15]), .B(A[15]), .ZN(n43) );
  XOR2_X1 U60 ( .A(B[12]), .B(A[12]), .Z(n44) );
  XOR2_X1 U61 ( .A(n5), .B(n44), .Z(SUM[12]) );
  NAND2_X1 U62 ( .A1(carry[12]), .A2(B[12]), .ZN(n45) );
  NAND2_X1 U63 ( .A1(n15), .A2(A[12]), .ZN(n46) );
  NAND2_X1 U64 ( .A1(B[12]), .A2(A[12]), .ZN(n47) );
  NAND3_X1 U65 ( .A1(n45), .A2(n46), .A3(n47), .ZN(carry[13]) );
  XNOR2_X1 U66 ( .A(B[14]), .B(n48), .ZN(n57) );
  XOR2_X1 U67 ( .A(B[6]), .B(A[6]), .Z(n49) );
  XOR2_X1 U68 ( .A(carry[6]), .B(n49), .Z(SUM[6]) );
  NAND2_X1 U69 ( .A1(n16), .A2(B[6]), .ZN(n50) );
  NAND2_X1 U70 ( .A1(n16), .A2(A[6]), .ZN(n51) );
  NAND2_X1 U71 ( .A1(B[6]), .A2(A[6]), .ZN(n52) );
  NAND3_X1 U72 ( .A1(n50), .A2(n51), .A3(n52), .ZN(carry[7]) );
  XOR2_X1 U73 ( .A(B[7]), .B(A[7]), .Z(n53) );
  XOR2_X1 U74 ( .A(n25), .B(n53), .Z(SUM[7]) );
  NAND2_X1 U75 ( .A1(n25), .A2(B[7]), .ZN(n54) );
  NAND2_X1 U76 ( .A1(carry[7]), .A2(A[7]), .ZN(n55) );
  NAND2_X1 U77 ( .A1(B[7]), .A2(A[7]), .ZN(n56) );
  NAND3_X1 U78 ( .A1(n54), .A2(n55), .A3(n56), .ZN(carry[8]) );
  XOR2_X1 U79 ( .A(n57), .B(n26), .Z(SUM[14]) );
  NAND2_X1 U80 ( .A1(carry[14]), .A2(B[14]), .ZN(n58) );
  NAND2_X1 U81 ( .A1(n26), .A2(A[14]), .ZN(n59) );
  NAND2_X1 U82 ( .A1(B[14]), .A2(A[14]), .ZN(n60) );
  NAND3_X1 U83 ( .A1(n59), .A2(n58), .A3(n60), .ZN(carry[15]) );
  XOR2_X1 U84 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U85 ( .A1(B[0]), .A2(A[0]), .ZN(n62) );
endmodule


module datapath_DW_mult_tc_1 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14, n15, n17, n18,
         n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343;

  FA_X1 U2 ( .A(n283), .B(n15), .CI(n2), .CO(n1), .S(product[14]) );
  FA_X1 U10 ( .A(n46), .B(n49), .CI(n10), .CO(n9), .S(product[6]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n286), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n285), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n289), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n288), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n291), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n101), .B(n88), .CI(n94), .CO(n53), .S(n54) );
  CLKBUF_X3 U157 ( .A(a[1]), .Z(n206) );
  NAND2_X1 U158 ( .A1(n309), .A2(n338), .ZN(n311) );
  INV_X1 U159 ( .A(n15), .ZN(n282) );
  BUF_X1 U160 ( .A(n280), .Z(n248) );
  NOR2_X1 U161 ( .A1(n276), .A2(n248), .ZN(n96) );
  CLKBUF_X1 U162 ( .A(n7), .Z(n207) );
  AND2_X1 U163 ( .A1(n209), .A2(n102), .ZN(n208) );
  OAI22_X1 U164 ( .A1(n300), .A2(n301), .B1(n302), .B2(n275), .ZN(n209) );
  OAI22_X1 U165 ( .A1(n277), .A2(n295), .B1(n341), .B2(n293), .ZN(n210) );
  XOR2_X2 U166 ( .A(a[6]), .B(n287), .Z(n320) );
  CLKBUF_X1 U167 ( .A(n249), .Z(n211) );
  NAND3_X1 U168 ( .A1(n246), .A2(n245), .A3(n247), .ZN(n212) );
  NAND3_X1 U169 ( .A1(n222), .A2(n223), .A3(n224), .ZN(n213) );
  XOR2_X1 U170 ( .A(n103), .B(n96), .Z(n214) );
  XOR2_X1 U171 ( .A(n14), .B(n214), .Z(product[2]) );
  NAND2_X1 U172 ( .A1(n14), .A2(n210), .ZN(n215) );
  NAND2_X1 U173 ( .A1(n14), .A2(n96), .ZN(n216) );
  NAND2_X1 U174 ( .A1(n210), .A2(n96), .ZN(n217) );
  NAND3_X1 U175 ( .A1(n215), .A2(n216), .A3(n217), .ZN(n13) );
  CLKBUF_X1 U176 ( .A(b[1]), .Z(n278) );
  XOR2_X1 U177 ( .A(n209), .B(n102), .Z(n218) );
  XNOR2_X1 U178 ( .A(n13), .B(n219), .ZN(product[3]) );
  XNOR2_X1 U179 ( .A(n218), .B(n71), .ZN(n219) );
  CLKBUF_X1 U180 ( .A(n245), .Z(n220) );
  XNOR2_X1 U181 ( .A(n221), .B(n239), .ZN(product[4]) );
  XNOR2_X1 U182 ( .A(n54), .B(n208), .ZN(n221) );
  NAND2_X1 U183 ( .A1(n13), .A2(n56), .ZN(n222) );
  NAND2_X1 U184 ( .A1(n13), .A2(n71), .ZN(n223) );
  NAND2_X1 U185 ( .A1(n56), .A2(n71), .ZN(n224) );
  NAND3_X1 U186 ( .A1(n222), .A2(n223), .A3(n224), .ZN(n12) );
  CLKBUF_X1 U187 ( .A(n213), .Z(n239) );
  CLKBUF_X1 U188 ( .A(n256), .Z(n225) );
  XOR2_X1 U189 ( .A(n40), .B(n45), .Z(n226) );
  XOR2_X1 U190 ( .A(n9), .B(n226), .Z(product[7]) );
  NAND2_X1 U191 ( .A1(n9), .A2(n40), .ZN(n227) );
  NAND2_X1 U192 ( .A1(n9), .A2(n45), .ZN(n228) );
  NAND2_X1 U193 ( .A1(n40), .A2(n45), .ZN(n229) );
  NAND3_X1 U194 ( .A1(n227), .A2(n228), .A3(n229), .ZN(n8) );
  NAND3_X1 U195 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n230) );
  NAND3_X1 U196 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n231) );
  NAND3_X1 U197 ( .A1(n246), .A2(n245), .A3(n247), .ZN(n232) );
  NAND3_X1 U198 ( .A1(n256), .A2(n255), .A3(n257), .ZN(n233) );
  NAND3_X1 U199 ( .A1(n225), .A2(n255), .A3(n257), .ZN(n234) );
  XOR2_X1 U200 ( .A(n34), .B(n39), .Z(n235) );
  XOR2_X1 U201 ( .A(n8), .B(n235), .Z(product[8]) );
  NAND2_X1 U202 ( .A1(n8), .A2(n34), .ZN(n236) );
  NAND2_X1 U203 ( .A1(n8), .A2(n39), .ZN(n237) );
  NAND2_X1 U204 ( .A1(n34), .A2(n39), .ZN(n238) );
  NAND3_X1 U205 ( .A1(n237), .A2(n236), .A3(n238), .ZN(n7) );
  XOR2_X1 U206 ( .A(n33), .B(n28), .Z(n240) );
  XOR2_X1 U207 ( .A(n207), .B(n240), .Z(product[9]) );
  NAND2_X1 U208 ( .A1(n7), .A2(n33), .ZN(n241) );
  NAND2_X1 U209 ( .A1(n7), .A2(n28), .ZN(n242) );
  NAND2_X1 U210 ( .A1(n33), .A2(n28), .ZN(n243) );
  NAND3_X1 U211 ( .A1(n241), .A2(n242), .A3(n243), .ZN(n6) );
  XOR2_X1 U212 ( .A(n18), .B(n19), .Z(n244) );
  XOR2_X1 U213 ( .A(n234), .B(n244), .Z(product[12]) );
  NAND2_X1 U214 ( .A1(n233), .A2(n18), .ZN(n245) );
  NAND2_X1 U215 ( .A1(n4), .A2(n19), .ZN(n246) );
  NAND2_X1 U216 ( .A1(n18), .A2(n19), .ZN(n247) );
  NAND3_X1 U217 ( .A1(n220), .A2(n246), .A3(n247), .ZN(n3) );
  XOR2_X1 U218 ( .A(n95), .B(n102), .Z(n56) );
  NAND3_X1 U219 ( .A1(n252), .A2(n251), .A3(n253), .ZN(n249) );
  XOR2_X1 U220 ( .A(n27), .B(n24), .Z(n250) );
  XOR2_X1 U221 ( .A(n231), .B(n250), .Z(product[10]) );
  NAND2_X1 U222 ( .A1(n230), .A2(n27), .ZN(n251) );
  NAND2_X1 U223 ( .A1(n6), .A2(n24), .ZN(n252) );
  NAND2_X1 U224 ( .A1(n27), .A2(n24), .ZN(n253) );
  NAND3_X1 U225 ( .A1(n251), .A2(n252), .A3(n253), .ZN(n5) );
  XOR2_X1 U226 ( .A(n23), .B(n20), .Z(n254) );
  XOR2_X1 U227 ( .A(n211), .B(n254), .Z(product[11]) );
  NAND2_X1 U228 ( .A1(n5), .A2(n23), .ZN(n255) );
  NAND2_X1 U229 ( .A1(n249), .A2(n20), .ZN(n256) );
  NAND2_X1 U230 ( .A1(n23), .A2(n20), .ZN(n257) );
  NAND3_X1 U231 ( .A1(n256), .A2(n255), .A3(n257), .ZN(n4) );
  NAND3_X1 U232 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n258) );
  NAND3_X1 U233 ( .A1(n260), .A2(n261), .A3(n262), .ZN(n259) );
  NAND2_X1 U234 ( .A1(n54), .A2(n208), .ZN(n260) );
  NAND2_X1 U235 ( .A1(n54), .A2(n213), .ZN(n261) );
  NAND2_X1 U236 ( .A1(n208), .A2(n12), .ZN(n262) );
  XOR2_X1 U237 ( .A(n50), .B(n53), .Z(n263) );
  XOR2_X1 U238 ( .A(n263), .B(n258), .Z(product[5]) );
  NAND2_X1 U239 ( .A1(n50), .A2(n53), .ZN(n264) );
  NAND2_X1 U240 ( .A1(n259), .A2(n50), .ZN(n265) );
  NAND2_X1 U241 ( .A1(n259), .A2(n53), .ZN(n266) );
  NAND3_X1 U242 ( .A1(n265), .A2(n266), .A3(n264), .ZN(n10) );
  XOR2_X1 U243 ( .A(n17), .B(n282), .Z(n267) );
  XOR2_X1 U244 ( .A(n3), .B(n267), .Z(product[13]) );
  NAND2_X1 U245 ( .A1(n212), .A2(n17), .ZN(n268) );
  NAND2_X1 U246 ( .A1(n232), .A2(n282), .ZN(n269) );
  NAND2_X1 U247 ( .A1(n17), .A2(n282), .ZN(n270) );
  NAND3_X1 U248 ( .A1(n268), .A2(n269), .A3(n270), .ZN(n2) );
  INV_X2 U249 ( .A(n280), .ZN(n279) );
  NAND2_X2 U250 ( .A1(n299), .A2(n337), .ZN(n301) );
  NAND2_X1 U251 ( .A1(a[4]), .A2(a[3]), .ZN(n273) );
  NAND2_X1 U252 ( .A1(n271), .A2(n272), .ZN(n274) );
  NAND2_X2 U253 ( .A1(n273), .A2(n274), .ZN(n309) );
  INV_X1 U254 ( .A(a[4]), .ZN(n271) );
  INV_X1 U255 ( .A(a[3]), .ZN(n272) );
  BUF_X1 U256 ( .A(n299), .Z(n276) );
  CLKBUF_X1 U257 ( .A(n299), .Z(n275) );
  XNOR2_X1 U258 ( .A(a[2]), .B(n206), .ZN(n299) );
  INV_X1 U259 ( .A(n21), .ZN(n285) );
  INV_X1 U260 ( .A(n318), .ZN(n286) );
  INV_X1 U261 ( .A(n329), .ZN(n283) );
  INV_X1 U262 ( .A(n298), .ZN(n291) );
  INV_X1 U263 ( .A(n307), .ZN(n289) );
  INV_X1 U264 ( .A(n31), .ZN(n288) );
  INV_X1 U265 ( .A(b[0]), .ZN(n280) );
  INV_X1 U266 ( .A(a[0]), .ZN(n293) );
  INV_X1 U267 ( .A(a[5]), .ZN(n287) );
  INV_X1 U268 ( .A(a[7]), .ZN(n284) );
  INV_X1 U269 ( .A(n1), .ZN(product[15]) );
  INV_X1 U270 ( .A(a[3]), .ZN(n290) );
  XNOR2_X1 U271 ( .A(b[1]), .B(n206), .ZN(n277) );
  INV_X1 U272 ( .A(n206), .ZN(n292) );
  NOR2_X1 U273 ( .A1(n293), .A2(n248), .ZN(product[0]) );
  OAI22_X1 U274 ( .A1(n294), .A2(n295), .B1(n296), .B2(n293), .ZN(n99) );
  OAI22_X1 U275 ( .A1(n296), .A2(n295), .B1(n297), .B2(n293), .ZN(n98) );
  XNOR2_X1 U276 ( .A(b[6]), .B(n206), .ZN(n296) );
  OAI22_X1 U277 ( .A1(n293), .A2(n297), .B1(n295), .B2(n297), .ZN(n298) );
  XNOR2_X1 U278 ( .A(b[7]), .B(n206), .ZN(n297) );
  OAI22_X1 U279 ( .A1(n300), .A2(n301), .B1(n302), .B2(n275), .ZN(n95) );
  XNOR2_X1 U280 ( .A(a[3]), .B(n279), .ZN(n300) );
  OAI22_X1 U281 ( .A1(n302), .A2(n301), .B1(n276), .B2(n303), .ZN(n94) );
  XNOR2_X1 U282 ( .A(n278), .B(a[3]), .ZN(n302) );
  OAI22_X1 U283 ( .A1(n303), .A2(n301), .B1(n276), .B2(n304), .ZN(n93) );
  XNOR2_X1 U284 ( .A(b[2]), .B(a[3]), .ZN(n303) );
  OAI22_X1 U285 ( .A1(n304), .A2(n301), .B1(n275), .B2(n305), .ZN(n92) );
  XNOR2_X1 U286 ( .A(b[3]), .B(a[3]), .ZN(n304) );
  OAI22_X1 U287 ( .A1(n305), .A2(n301), .B1(n275), .B2(n306), .ZN(n91) );
  XNOR2_X1 U288 ( .A(b[4]), .B(a[3]), .ZN(n305) );
  OAI22_X1 U289 ( .A1(n308), .A2(n276), .B1(n301), .B2(n308), .ZN(n307) );
  NOR2_X1 U290 ( .A1(n309), .A2(n248), .ZN(n88) );
  OAI22_X1 U291 ( .A1(n310), .A2(n311), .B1(n309), .B2(n312), .ZN(n87) );
  XNOR2_X1 U292 ( .A(a[5]), .B(n279), .ZN(n310) );
  OAI22_X1 U293 ( .A1(n312), .A2(n311), .B1(n309), .B2(n313), .ZN(n86) );
  XNOR2_X1 U294 ( .A(n278), .B(a[5]), .ZN(n312) );
  OAI22_X1 U295 ( .A1(n313), .A2(n311), .B1(n309), .B2(n314), .ZN(n85) );
  XNOR2_X1 U296 ( .A(b[2]), .B(a[5]), .ZN(n313) );
  OAI22_X1 U297 ( .A1(n314), .A2(n311), .B1(n309), .B2(n315), .ZN(n84) );
  XNOR2_X1 U298 ( .A(b[3]), .B(a[5]), .ZN(n314) );
  OAI22_X1 U299 ( .A1(n315), .A2(n311), .B1(n309), .B2(n316), .ZN(n83) );
  XNOR2_X1 U300 ( .A(b[4]), .B(a[5]), .ZN(n315) );
  OAI22_X1 U301 ( .A1(n316), .A2(n311), .B1(n309), .B2(n317), .ZN(n82) );
  XNOR2_X1 U302 ( .A(b[5]), .B(a[5]), .ZN(n316) );
  OAI22_X1 U303 ( .A1(n319), .A2(n309), .B1(n311), .B2(n319), .ZN(n318) );
  NOR2_X1 U304 ( .A1(n320), .A2(n248), .ZN(n80) );
  OAI22_X1 U305 ( .A1(n321), .A2(n322), .B1(n320), .B2(n323), .ZN(n79) );
  XNOR2_X1 U306 ( .A(a[7]), .B(n279), .ZN(n321) );
  OAI22_X1 U307 ( .A1(n324), .A2(n322), .B1(n320), .B2(n325), .ZN(n77) );
  OAI22_X1 U308 ( .A1(n325), .A2(n322), .B1(n320), .B2(n326), .ZN(n76) );
  XNOR2_X1 U309 ( .A(b[3]), .B(a[7]), .ZN(n325) );
  OAI22_X1 U310 ( .A1(n326), .A2(n322), .B1(n320), .B2(n327), .ZN(n75) );
  XNOR2_X1 U311 ( .A(b[4]), .B(a[7]), .ZN(n326) );
  OAI22_X1 U312 ( .A1(n327), .A2(n322), .B1(n320), .B2(n328), .ZN(n74) );
  XNOR2_X1 U313 ( .A(b[5]), .B(a[7]), .ZN(n327) );
  OAI22_X1 U314 ( .A1(n330), .A2(n320), .B1(n322), .B2(n330), .ZN(n329) );
  OAI21_X1 U315 ( .B1(n279), .B2(n292), .A(n295), .ZN(n72) );
  OAI21_X1 U316 ( .B1(n290), .B2(n301), .A(n331), .ZN(n71) );
  OR3_X1 U317 ( .A1(n275), .A2(n279), .A3(n290), .ZN(n331) );
  OAI21_X1 U318 ( .B1(n287), .B2(n311), .A(n332), .ZN(n70) );
  OR3_X1 U319 ( .A1(n309), .A2(n279), .A3(n287), .ZN(n332) );
  OAI21_X1 U320 ( .B1(n284), .B2(n322), .A(n333), .ZN(n69) );
  OR3_X1 U321 ( .A1(n320), .A2(n279), .A3(n284), .ZN(n333) );
  XNOR2_X1 U322 ( .A(n334), .B(n335), .ZN(n38) );
  OR2_X1 U323 ( .A1(n334), .A2(n335), .ZN(n37) );
  OAI22_X1 U324 ( .A1(n306), .A2(n301), .B1(n276), .B2(n336), .ZN(n335) );
  XNOR2_X1 U325 ( .A(b[5]), .B(a[3]), .ZN(n306) );
  OAI22_X1 U326 ( .A1(n323), .A2(n322), .B1(n320), .B2(n324), .ZN(n334) );
  XNOR2_X1 U327 ( .A(b[2]), .B(a[7]), .ZN(n324) );
  XNOR2_X1 U328 ( .A(n278), .B(a[7]), .ZN(n323) );
  OAI22_X1 U329 ( .A1(n336), .A2(n301), .B1(n275), .B2(n308), .ZN(n31) );
  XNOR2_X1 U330 ( .A(b[7]), .B(a[3]), .ZN(n308) );
  XNOR2_X1 U331 ( .A(n290), .B(a[2]), .ZN(n337) );
  XNOR2_X1 U332 ( .A(b[6]), .B(a[3]), .ZN(n336) );
  OAI22_X1 U333 ( .A1(n317), .A2(n311), .B1(n309), .B2(n319), .ZN(n21) );
  XNOR2_X1 U334 ( .A(b[7]), .B(a[5]), .ZN(n319) );
  XNOR2_X1 U335 ( .A(n287), .B(a[4]), .ZN(n338) );
  XNOR2_X1 U336 ( .A(b[6]), .B(a[5]), .ZN(n317) );
  OAI22_X1 U337 ( .A1(n328), .A2(n322), .B1(n320), .B2(n330), .ZN(n15) );
  XNOR2_X1 U338 ( .A(b[7]), .B(a[7]), .ZN(n330) );
  NAND2_X1 U339 ( .A1(n320), .A2(n339), .ZN(n322) );
  XNOR2_X1 U340 ( .A(n284), .B(a[6]), .ZN(n339) );
  XNOR2_X1 U341 ( .A(b[6]), .B(a[7]), .ZN(n328) );
  OAI22_X1 U342 ( .A1(n279), .A2(n295), .B1(n340), .B2(n293), .ZN(n104) );
  OAI22_X1 U343 ( .A1(n277), .A2(n295), .B1(n341), .B2(n293), .ZN(n103) );
  XNOR2_X1 U344 ( .A(b[1]), .B(n206), .ZN(n340) );
  OAI22_X1 U345 ( .A1(n341), .A2(n295), .B1(n342), .B2(n293), .ZN(n102) );
  XNOR2_X1 U346 ( .A(b[2]), .B(n206), .ZN(n341) );
  OAI22_X1 U347 ( .A1(n342), .A2(n295), .B1(n343), .B2(n293), .ZN(n101) );
  XNOR2_X1 U348 ( .A(b[3]), .B(n206), .ZN(n342) );
  OAI22_X1 U349 ( .A1(n343), .A2(n295), .B1(n294), .B2(n293), .ZN(n100) );
  XNOR2_X1 U350 ( .A(b[5]), .B(n206), .ZN(n294) );
  NAND2_X1 U351 ( .A1(n206), .A2(n293), .ZN(n295) );
  XNOR2_X1 U352 ( .A(b[4]), .B(n206), .ZN(n343) );
endmodule


module datapath_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n74;
  wire   [15:1] carry;

  FA_X1 U1_4 ( .A(B[4]), .B(A[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n74), .CO(carry[2]), .S(SUM[1]) );
  XNOR2_X1 U1 ( .A(B[15]), .B(A[15]), .ZN(n58) );
  INV_X1 U2 ( .A(A[14]), .ZN(n45) );
  NAND3_X1 U3 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n1) );
  NAND3_X1 U4 ( .A1(n14), .A2(n15), .A3(n16), .ZN(n2) );
  NAND3_X1 U5 ( .A1(n72), .A2(n71), .A3(n70), .ZN(n3) );
  NAND3_X1 U6 ( .A1(n72), .A2(n71), .A3(n70), .ZN(n4) );
  NAND3_X1 U7 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n5) );
  NAND3_X1 U8 ( .A1(n60), .A2(n61), .A3(n62), .ZN(n6) );
  XOR2_X1 U9 ( .A(carry[2]), .B(A[2]), .Z(n7) );
  XOR2_X1 U10 ( .A(B[2]), .B(n7), .Z(SUM[2]) );
  NAND2_X1 U11 ( .A1(B[2]), .A2(carry[2]), .ZN(n8) );
  NAND2_X1 U12 ( .A1(B[2]), .A2(A[2]), .ZN(n9) );
  NAND2_X1 U13 ( .A1(carry[2]), .A2(A[2]), .ZN(n10) );
  NAND3_X1 U14 ( .A1(n8), .A2(n9), .A3(n10), .ZN(carry[3]) );
  CLKBUF_X1 U15 ( .A(n39), .Z(n11) );
  CLKBUF_X1 U16 ( .A(n53), .Z(n12) );
  XOR2_X1 U17 ( .A(B[10]), .B(A[10]), .Z(n13) );
  XOR2_X1 U18 ( .A(n4), .B(n13), .Z(SUM[10]) );
  NAND2_X1 U19 ( .A1(n3), .A2(B[10]), .ZN(n14) );
  NAND2_X1 U20 ( .A1(carry[10]), .A2(A[10]), .ZN(n15) );
  NAND2_X1 U21 ( .A1(B[10]), .A2(A[10]), .ZN(n16) );
  NAND3_X1 U22 ( .A1(n14), .A2(n15), .A3(n16), .ZN(carry[11]) );
  CLKBUF_X1 U23 ( .A(n52), .Z(n17) );
  NAND3_X1 U24 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n18) );
  NAND3_X1 U25 ( .A1(n28), .A2(n29), .A3(n30), .ZN(n19) );
  NAND3_X1 U26 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n20) );
  NAND3_X1 U27 ( .A1(n38), .A2(n11), .A3(n40), .ZN(n21) );
  CLKBUF_X1 U28 ( .A(n35), .Z(n22) );
  XOR2_X1 U29 ( .A(B[3]), .B(A[3]), .Z(n23) );
  XOR2_X1 U30 ( .A(carry[3]), .B(n23), .Z(SUM[3]) );
  NAND2_X1 U31 ( .A1(carry[3]), .A2(B[3]), .ZN(n24) );
  NAND2_X1 U32 ( .A1(carry[3]), .A2(A[3]), .ZN(n25) );
  NAND2_X1 U33 ( .A1(B[3]), .A2(A[3]), .ZN(n26) );
  NAND3_X1 U34 ( .A1(n24), .A2(n25), .A3(n26), .ZN(carry[4]) );
  XOR2_X1 U35 ( .A(B[5]), .B(A[5]), .Z(n27) );
  XOR2_X1 U36 ( .A(carry[5]), .B(n27), .Z(SUM[5]) );
  NAND2_X1 U37 ( .A1(carry[5]), .A2(B[5]), .ZN(n28) );
  NAND2_X1 U38 ( .A1(carry[5]), .A2(A[5]), .ZN(n29) );
  NAND2_X1 U39 ( .A1(B[5]), .A2(A[5]), .ZN(n30) );
  NAND3_X1 U40 ( .A1(n28), .A2(n29), .A3(n30), .ZN(carry[6]) );
  NAND3_X1 U41 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n31) );
  CLKBUF_X1 U42 ( .A(n67), .Z(n32) );
  XOR2_X1 U43 ( .A(B[6]), .B(A[6]), .Z(n33) );
  XOR2_X1 U44 ( .A(n19), .B(n33), .Z(SUM[6]) );
  NAND2_X1 U45 ( .A1(n18), .A2(B[6]), .ZN(n34) );
  NAND2_X1 U46 ( .A1(carry[6]), .A2(A[6]), .ZN(n35) );
  NAND2_X1 U47 ( .A1(B[6]), .A2(A[6]), .ZN(n36) );
  NAND3_X1 U48 ( .A1(n34), .A2(n22), .A3(n36), .ZN(carry[7]) );
  XOR2_X1 U49 ( .A(B[11]), .B(A[11]), .Z(n37) );
  XOR2_X1 U50 ( .A(n2), .B(n37), .Z(SUM[11]) );
  NAND2_X1 U51 ( .A1(n1), .A2(B[11]), .ZN(n38) );
  NAND2_X1 U52 ( .A1(carry[11]), .A2(A[11]), .ZN(n39) );
  NAND2_X1 U53 ( .A1(B[11]), .A2(A[11]), .ZN(n40) );
  NAND3_X1 U54 ( .A1(n38), .A2(n39), .A3(n40), .ZN(carry[12]) );
  NAND3_X1 U55 ( .A1(n60), .A2(n61), .A3(n62), .ZN(n41) );
  NAND3_X1 U56 ( .A1(n55), .A2(n56), .A3(n57), .ZN(n42) );
  NAND3_X1 U57 ( .A1(n53), .A2(n52), .A3(n51), .ZN(n43) );
  NAND3_X1 U58 ( .A1(n51), .A2(n17), .A3(n12), .ZN(n44) );
  XNOR2_X1 U59 ( .A(B[14]), .B(n45), .ZN(n46) );
  XOR2_X1 U60 ( .A(n42), .B(n46), .Z(SUM[14]) );
  NAND2_X1 U61 ( .A1(B[14]), .A2(n42), .ZN(n47) );
  NAND2_X1 U62 ( .A1(carry[14]), .A2(A[14]), .ZN(n48) );
  NAND2_X1 U63 ( .A1(B[14]), .A2(A[14]), .ZN(n49) );
  NAND3_X1 U64 ( .A1(n47), .A2(n48), .A3(n49), .ZN(carry[15]) );
  XOR2_X1 U65 ( .A(A[12]), .B(B[12]), .Z(n50) );
  XOR2_X1 U66 ( .A(n50), .B(n21), .Z(SUM[12]) );
  NAND2_X1 U67 ( .A1(A[12]), .A2(B[12]), .ZN(n51) );
  NAND2_X1 U68 ( .A1(A[12]), .A2(n20), .ZN(n52) );
  NAND2_X1 U69 ( .A1(B[12]), .A2(carry[12]), .ZN(n53) );
  NAND3_X1 U70 ( .A1(n53), .A2(n52), .A3(n51), .ZN(carry[13]) );
  XOR2_X1 U71 ( .A(A[13]), .B(B[13]), .Z(n54) );
  XOR2_X1 U72 ( .A(n54), .B(n44), .Z(SUM[13]) );
  NAND2_X1 U73 ( .A1(A[13]), .A2(B[13]), .ZN(n55) );
  NAND2_X1 U74 ( .A1(A[13]), .A2(n43), .ZN(n56) );
  NAND2_X1 U75 ( .A1(B[13]), .A2(carry[13]), .ZN(n57) );
  NAND3_X1 U76 ( .A1(n57), .A2(n56), .A3(n55), .ZN(carry[14]) );
  XNOR2_X1 U77 ( .A(carry[15]), .B(n58), .ZN(SUM[15]) );
  XOR2_X1 U78 ( .A(B[7]), .B(A[7]), .Z(n59) );
  XOR2_X1 U79 ( .A(carry[7]), .B(n59), .Z(SUM[7]) );
  NAND2_X1 U80 ( .A1(n5), .A2(B[7]), .ZN(n60) );
  NAND2_X1 U81 ( .A1(n31), .A2(A[7]), .ZN(n61) );
  NAND2_X1 U82 ( .A1(B[7]), .A2(A[7]), .ZN(n62) );
  NAND3_X1 U83 ( .A1(n60), .A2(n61), .A3(n62), .ZN(carry[8]) );
  NAND3_X1 U84 ( .A1(n68), .A2(n67), .A3(n66), .ZN(n63) );
  NAND3_X1 U85 ( .A1(n66), .A2(n32), .A3(n68), .ZN(n64) );
  XOR2_X1 U86 ( .A(A[8]), .B(B[8]), .Z(n65) );
  XOR2_X1 U87 ( .A(n65), .B(n6), .Z(SUM[8]) );
  NAND2_X1 U88 ( .A1(A[8]), .A2(B[8]), .ZN(n66) );
  NAND2_X1 U89 ( .A1(A[8]), .A2(carry[8]), .ZN(n67) );
  NAND2_X1 U90 ( .A1(B[8]), .A2(n41), .ZN(n68) );
  NAND3_X1 U91 ( .A1(n66), .A2(n67), .A3(n68), .ZN(carry[9]) );
  XOR2_X1 U92 ( .A(A[9]), .B(B[9]), .Z(n69) );
  XOR2_X1 U93 ( .A(n69), .B(n64), .Z(SUM[9]) );
  NAND2_X1 U94 ( .A1(A[9]), .A2(B[9]), .ZN(n70) );
  NAND2_X1 U95 ( .A1(A[9]), .A2(carry[9]), .ZN(n71) );
  NAND2_X1 U96 ( .A1(B[9]), .A2(n63), .ZN(n72) );
  NAND3_X1 U97 ( .A1(n72), .A2(n71), .A3(n70), .ZN(carry[10]) );
  XOR2_X1 U98 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U99 ( .A1(B[0]), .A2(A[0]), .ZN(n74) );
endmodule


module datapath_DW_mult_tc_0 ( a, b, product );
  input [7:0] a;
  input [7:0] b;
  output [15:0] product;
  wire   n2, n3, n4, n5, n7, n8, n10, n11, n12, n13, n14, n15, n17, n18, n19,
         n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n69, n70, n71, n72, n74, n75, n76,
         n77, n79, n80, n82, n83, n84, n85, n86, n87, n88, n91, n92, n93, n94,
         n95, n96, n98, n99, n100, n101, n102, n103, n104, n206, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352;

  FA_X1 U12 ( .A(n54), .B(n55), .CI(n12), .CO(n11), .S(product[4]) );
  HA_X1 U15 ( .A(n104), .B(n72), .CO(n14), .S(product[1]) );
  FA_X1 U17 ( .A(n74), .B(n21), .CI(n295), .CO(n17), .S(n18) );
  FA_X1 U18 ( .A(n294), .B(n75), .CI(n25), .CO(n19), .S(n20) );
  FA_X1 U20 ( .A(n29), .B(n76), .CI(n26), .CO(n23), .S(n24) );
  FA_X1 U21 ( .A(n82), .B(n31), .CI(n298), .CO(n25), .S(n26) );
  FA_X1 U22 ( .A(n35), .B(n37), .CI(n30), .CO(n27), .S(n28) );
  FA_X1 U23 ( .A(n77), .B(n83), .CI(n297), .CO(n29), .S(n30) );
  FA_X1 U25 ( .A(n41), .B(n38), .CI(n36), .CO(n33), .S(n34) );
  FA_X1 U26 ( .A(n300), .B(n84), .CI(n43), .CO(n35), .S(n36) );
  FA_X1 U29 ( .A(n47), .B(n44), .CI(n42), .CO(n39), .S(n40) );
  FA_X1 U30 ( .A(n85), .B(n98), .CI(n91), .CO(n41), .S(n42) );
  HA_X1 U31 ( .A(n69), .B(n79), .CO(n43), .S(n44) );
  FA_X1 U32 ( .A(n51), .B(n86), .CI(n48), .CO(n45), .S(n46) );
  FA_X1 U33 ( .A(n99), .B(n80), .CI(n92), .CO(n47), .S(n48) );
  FA_X1 U34 ( .A(n93), .B(n100), .CI(n52), .CO(n49), .S(n50) );
  HA_X1 U35 ( .A(n70), .B(n87), .CO(n51), .S(n52) );
  FA_X1 U36 ( .A(n88), .B(n94), .CI(n101), .CO(n53), .S(n54) );
  HA_X1 U37 ( .A(n218), .B(n102), .CO(n55), .S(n56) );
  INV_X1 U157 ( .A(n290), .ZN(n289) );
  INV_X1 U158 ( .A(n15), .ZN(n291) );
  XNOR2_X1 U159 ( .A(n292), .B(n15), .ZN(n206) );
  AND3_X1 U160 ( .A1(n262), .A2(n263), .A3(n264), .ZN(product[15]) );
  XNOR2_X1 U161 ( .A(n222), .B(a[3]), .ZN(n208) );
  NAND3_X1 U162 ( .A1(n223), .A2(n224), .A3(n225), .ZN(n209) );
  NAND3_X1 U163 ( .A1(n223), .A2(n224), .A3(n225), .ZN(n210) );
  XNOR2_X1 U164 ( .A(n11), .B(n211), .ZN(product[5]) );
  XNOR2_X1 U165 ( .A(n50), .B(n53), .ZN(n211) );
  XNOR2_X1 U166 ( .A(a[6]), .B(a[5]), .ZN(n329) );
  NAND3_X1 U167 ( .A1(n234), .A2(n235), .A3(n236), .ZN(n212) );
  NAND3_X1 U168 ( .A1(n279), .A2(n278), .A3(n280), .ZN(n213) );
  NAND3_X1 U169 ( .A1(n250), .A2(n249), .A3(n251), .ZN(n214) );
  NAND3_X1 U170 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n215) );
  NAND2_X1 U171 ( .A1(n14), .A2(n96), .ZN(n216) );
  NAND3_X1 U172 ( .A1(n216), .A2(n257), .A3(n256), .ZN(n217) );
  OAI22_X1 U173 ( .A1(n309), .A2(n310), .B1(n284), .B2(n208), .ZN(n218) );
  BUF_X1 U174 ( .A(b[1]), .Z(n222) );
  NAND2_X1 U175 ( .A1(n229), .A2(n34), .ZN(n219) );
  NAND3_X1 U176 ( .A1(n271), .A2(n272), .A3(n270), .ZN(n220) );
  NAND3_X1 U177 ( .A1(n270), .A2(n271), .A3(n272), .ZN(n221) );
  NAND2_X1 U178 ( .A1(n11), .A2(n50), .ZN(n223) );
  NAND2_X1 U179 ( .A1(n11), .A2(n53), .ZN(n224) );
  NAND2_X1 U180 ( .A1(n50), .A2(n53), .ZN(n225) );
  NAND3_X1 U181 ( .A1(n223), .A2(n224), .A3(n225), .ZN(n10) );
  XNOR2_X1 U182 ( .A(n226), .B(n238), .ZN(product[2]) );
  XNOR2_X1 U183 ( .A(n103), .B(n96), .ZN(n226) );
  NAND3_X1 U184 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n227) );
  NAND3_X1 U185 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n228) );
  NAND3_X1 U186 ( .A1(n275), .A2(n274), .A3(n276), .ZN(n229) );
  XNOR2_X1 U187 ( .A(n229), .B(n230), .ZN(product[8]) );
  XNOR2_X1 U188 ( .A(n34), .B(n39), .ZN(n230) );
  XOR2_X1 U189 ( .A(n231), .B(n232), .Z(product[9]) );
  AND3_X1 U190 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n231) );
  XNOR2_X1 U191 ( .A(n33), .B(n28), .ZN(n232) );
  XOR2_X1 U192 ( .A(n17), .B(n291), .Z(n233) );
  XOR2_X1 U193 ( .A(n228), .B(n233), .Z(product[13]) );
  NAND2_X1 U194 ( .A1(n227), .A2(n17), .ZN(n234) );
  NAND2_X1 U195 ( .A1(n3), .A2(n291), .ZN(n235) );
  NAND2_X1 U196 ( .A1(n17), .A2(n291), .ZN(n236) );
  NAND3_X1 U197 ( .A1(n234), .A2(n235), .A3(n236), .ZN(n2) );
  NAND3_X1 U198 ( .A1(n219), .A2(n246), .A3(n247), .ZN(n237) );
  AND2_X1 U199 ( .A1(n104), .A2(n72), .ZN(n238) );
  NAND3_X1 U200 ( .A1(n250), .A2(n249), .A3(n251), .ZN(n239) );
  NAND3_X1 U201 ( .A1(n279), .A2(n278), .A3(n280), .ZN(n240) );
  XOR2_X1 U202 ( .A(n18), .B(n19), .Z(n241) );
  XOR2_X1 U203 ( .A(n4), .B(n241), .Z(product[12]) );
  NAND2_X1 U204 ( .A1(n213), .A2(n18), .ZN(n242) );
  NAND2_X1 U205 ( .A1(n240), .A2(n19), .ZN(n243) );
  NAND2_X1 U206 ( .A1(n18), .A2(n19), .ZN(n244) );
  NAND3_X1 U207 ( .A1(n242), .A2(n243), .A3(n244), .ZN(n3) );
  NAND2_X1 U208 ( .A1(n229), .A2(n34), .ZN(n245) );
  NAND2_X1 U209 ( .A1(n8), .A2(n39), .ZN(n246) );
  NAND2_X1 U210 ( .A1(n34), .A2(n39), .ZN(n247) );
  NAND3_X1 U211 ( .A1(n245), .A2(n246), .A3(n247), .ZN(n7) );
  NAND3_X1 U212 ( .A1(n250), .A2(n249), .A3(n251), .ZN(n248) );
  NAND2_X1 U213 ( .A1(n237), .A2(n33), .ZN(n249) );
  NAND2_X1 U214 ( .A1(n7), .A2(n28), .ZN(n250) );
  NAND2_X1 U215 ( .A1(n33), .A2(n28), .ZN(n251) );
  XNOR2_X1 U216 ( .A(n2), .B(n206), .ZN(product[14]) );
  NAND3_X1 U217 ( .A1(n267), .A2(n266), .A3(n268), .ZN(n252) );
  NAND3_X1 U218 ( .A1(n256), .A2(n257), .A3(n216), .ZN(n253) );
  XNOR2_X1 U219 ( .A(n254), .B(n253), .ZN(product[3]) );
  XNOR2_X1 U220 ( .A(n56), .B(n71), .ZN(n254) );
  XOR2_X1 U221 ( .A(n95), .B(n102), .Z(n255) );
  NAND2_X1 U222 ( .A1(n103), .A2(n96), .ZN(n256) );
  NAND2_X1 U223 ( .A1(n103), .A2(n238), .ZN(n257) );
  NAND2_X1 U224 ( .A1(n14), .A2(n96), .ZN(n258) );
  NAND3_X1 U225 ( .A1(n258), .A2(n257), .A3(n256), .ZN(n13) );
  NAND2_X1 U226 ( .A1(n255), .A2(n71), .ZN(n259) );
  NAND2_X1 U227 ( .A1(n255), .A2(n217), .ZN(n260) );
  NAND2_X1 U228 ( .A1(n13), .A2(n71), .ZN(n261) );
  NAND3_X1 U229 ( .A1(n260), .A2(n261), .A3(n259), .ZN(n12) );
  NAND2_X1 U230 ( .A1(n212), .A2(n292), .ZN(n262) );
  NAND2_X1 U231 ( .A1(n212), .A2(n15), .ZN(n263) );
  NAND2_X1 U232 ( .A1(n292), .A2(n15), .ZN(n264) );
  XOR2_X1 U233 ( .A(n27), .B(n24), .Z(n265) );
  XOR2_X1 U234 ( .A(n214), .B(n265), .Z(product[10]) );
  NAND2_X1 U235 ( .A1(n239), .A2(n27), .ZN(n266) );
  NAND2_X1 U236 ( .A1(n248), .A2(n24), .ZN(n267) );
  NAND2_X1 U237 ( .A1(n27), .A2(n24), .ZN(n268) );
  NAND3_X1 U238 ( .A1(n266), .A2(n267), .A3(n268), .ZN(n5) );
  XOR2_X1 U239 ( .A(n46), .B(n49), .Z(n269) );
  XOR2_X1 U240 ( .A(n210), .B(n269), .Z(product[6]) );
  NAND2_X1 U241 ( .A1(n209), .A2(n46), .ZN(n270) );
  NAND2_X1 U242 ( .A1(n10), .A2(n49), .ZN(n271) );
  NAND2_X1 U243 ( .A1(n46), .A2(n49), .ZN(n272) );
  XOR2_X1 U244 ( .A(n40), .B(n45), .Z(n273) );
  XOR2_X1 U245 ( .A(n221), .B(n273), .Z(product[7]) );
  NAND2_X1 U246 ( .A1(n220), .A2(n40), .ZN(n274) );
  NAND2_X1 U247 ( .A1(n221), .A2(n45), .ZN(n275) );
  NAND2_X1 U248 ( .A1(n40), .A2(n45), .ZN(n276) );
  NAND3_X1 U249 ( .A1(n275), .A2(n274), .A3(n276), .ZN(n8) );
  XOR2_X1 U250 ( .A(n23), .B(n20), .Z(n277) );
  XOR2_X1 U251 ( .A(n215), .B(n277), .Z(product[11]) );
  NAND2_X1 U252 ( .A1(n252), .A2(n23), .ZN(n278) );
  NAND2_X1 U253 ( .A1(n5), .A2(n20), .ZN(n279) );
  NAND2_X1 U254 ( .A1(n23), .A2(n20), .ZN(n280) );
  NAND3_X1 U255 ( .A1(n278), .A2(n279), .A3(n280), .ZN(n4) );
  NAND2_X1 U256 ( .A1(a[4]), .A2(a[3]), .ZN(n282) );
  NAND2_X1 U257 ( .A1(n281), .A2(n299), .ZN(n283) );
  NAND2_X2 U258 ( .A1(n282), .A2(n283), .ZN(n318) );
  INV_X1 U259 ( .A(a[4]), .ZN(n281) );
  NAND2_X2 U260 ( .A1(n318), .A2(n347), .ZN(n320) );
  NAND2_X1 U261 ( .A1(n287), .A2(n288), .ZN(n284) );
  NAND2_X1 U262 ( .A1(n287), .A2(n288), .ZN(n285) );
  NAND2_X1 U263 ( .A1(n308), .A2(n346), .ZN(n310) );
  NAND2_X1 U264 ( .A1(n287), .A2(n288), .ZN(n308) );
  NAND2_X1 U265 ( .A1(a[2]), .A2(a[1]), .ZN(n287) );
  NAND2_X1 U266 ( .A1(n286), .A2(n301), .ZN(n288) );
  INV_X1 U267 ( .A(a[2]), .ZN(n286) );
  INV_X1 U268 ( .A(a[0]), .ZN(n302) );
  INV_X1 U269 ( .A(n21), .ZN(n294) );
  INV_X1 U270 ( .A(n327), .ZN(n295) );
  INV_X1 U271 ( .A(n338), .ZN(n292) );
  INV_X1 U272 ( .A(n307), .ZN(n300) );
  INV_X1 U273 ( .A(n316), .ZN(n298) );
  INV_X1 U274 ( .A(n31), .ZN(n297) );
  INV_X1 U275 ( .A(b[0]), .ZN(n290) );
  INV_X1 U276 ( .A(a[5]), .ZN(n296) );
  INV_X1 U277 ( .A(a[7]), .ZN(n293) );
  INV_X1 U278 ( .A(a[3]), .ZN(n299) );
  INV_X1 U279 ( .A(a[1]), .ZN(n301) );
  NOR2_X1 U280 ( .A1(n302), .A2(n290), .ZN(product[0]) );
  OAI22_X1 U281 ( .A1(n303), .A2(n304), .B1(n305), .B2(n302), .ZN(n99) );
  OAI22_X1 U282 ( .A1(n305), .A2(n304), .B1(n306), .B2(n302), .ZN(n98) );
  XNOR2_X1 U283 ( .A(b[6]), .B(a[1]), .ZN(n305) );
  OAI22_X1 U284 ( .A1(n302), .A2(n306), .B1(n304), .B2(n306), .ZN(n307) );
  XNOR2_X1 U285 ( .A(b[7]), .B(a[1]), .ZN(n306) );
  NOR2_X1 U286 ( .A1(n285), .A2(n290), .ZN(n96) );
  OAI22_X1 U287 ( .A1(n309), .A2(n310), .B1(n284), .B2(n311), .ZN(n95) );
  XNOR2_X1 U288 ( .A(a[3]), .B(n289), .ZN(n309) );
  OAI22_X1 U289 ( .A1(n311), .A2(n310), .B1(n284), .B2(n312), .ZN(n94) );
  XNOR2_X1 U290 ( .A(n222), .B(a[3]), .ZN(n311) );
  OAI22_X1 U291 ( .A1(n312), .A2(n310), .B1(n284), .B2(n313), .ZN(n93) );
  XNOR2_X1 U292 ( .A(b[2]), .B(a[3]), .ZN(n312) );
  OAI22_X1 U293 ( .A1(n313), .A2(n310), .B1(n285), .B2(n314), .ZN(n92) );
  XNOR2_X1 U294 ( .A(b[3]), .B(a[3]), .ZN(n313) );
  OAI22_X1 U295 ( .A1(n314), .A2(n310), .B1(n285), .B2(n315), .ZN(n91) );
  XNOR2_X1 U296 ( .A(b[4]), .B(a[3]), .ZN(n314) );
  OAI22_X1 U297 ( .A1(n317), .A2(n284), .B1(n310), .B2(n317), .ZN(n316) );
  NOR2_X1 U298 ( .A1(n318), .A2(n290), .ZN(n88) );
  OAI22_X1 U299 ( .A1(n319), .A2(n320), .B1(n318), .B2(n321), .ZN(n87) );
  XNOR2_X1 U300 ( .A(a[5]), .B(n289), .ZN(n319) );
  OAI22_X1 U301 ( .A1(n321), .A2(n320), .B1(n318), .B2(n322), .ZN(n86) );
  XNOR2_X1 U302 ( .A(b[1]), .B(a[5]), .ZN(n321) );
  OAI22_X1 U303 ( .A1(n322), .A2(n320), .B1(n318), .B2(n323), .ZN(n85) );
  XNOR2_X1 U304 ( .A(b[2]), .B(a[5]), .ZN(n322) );
  OAI22_X1 U305 ( .A1(n323), .A2(n320), .B1(n318), .B2(n324), .ZN(n84) );
  XNOR2_X1 U306 ( .A(b[3]), .B(a[5]), .ZN(n323) );
  OAI22_X1 U307 ( .A1(n324), .A2(n320), .B1(n318), .B2(n325), .ZN(n83) );
  XNOR2_X1 U308 ( .A(b[4]), .B(a[5]), .ZN(n324) );
  OAI22_X1 U309 ( .A1(n325), .A2(n320), .B1(n318), .B2(n326), .ZN(n82) );
  XNOR2_X1 U310 ( .A(b[5]), .B(a[5]), .ZN(n325) );
  OAI22_X1 U311 ( .A1(n328), .A2(n318), .B1(n320), .B2(n328), .ZN(n327) );
  NOR2_X1 U312 ( .A1(n329), .A2(n290), .ZN(n80) );
  OAI22_X1 U313 ( .A1(n330), .A2(n331), .B1(n329), .B2(n332), .ZN(n79) );
  XNOR2_X1 U314 ( .A(a[7]), .B(n289), .ZN(n330) );
  OAI22_X1 U315 ( .A1(n333), .A2(n331), .B1(n329), .B2(n334), .ZN(n77) );
  OAI22_X1 U316 ( .A1(n334), .A2(n331), .B1(n329), .B2(n335), .ZN(n76) );
  XNOR2_X1 U317 ( .A(b[3]), .B(a[7]), .ZN(n334) );
  OAI22_X1 U318 ( .A1(n335), .A2(n331), .B1(n329), .B2(n336), .ZN(n75) );
  XNOR2_X1 U319 ( .A(b[4]), .B(a[7]), .ZN(n335) );
  OAI22_X1 U320 ( .A1(n336), .A2(n331), .B1(n329), .B2(n337), .ZN(n74) );
  XNOR2_X1 U321 ( .A(b[5]), .B(a[7]), .ZN(n336) );
  OAI22_X1 U322 ( .A1(n339), .A2(n329), .B1(n331), .B2(n339), .ZN(n338) );
  OAI21_X1 U323 ( .B1(n289), .B2(n301), .A(n304), .ZN(n72) );
  OAI21_X1 U324 ( .B1(n299), .B2(n310), .A(n340), .ZN(n71) );
  OR3_X1 U325 ( .A1(n285), .A2(n289), .A3(n299), .ZN(n340) );
  OAI21_X1 U326 ( .B1(n296), .B2(n320), .A(n341), .ZN(n70) );
  OR3_X1 U327 ( .A1(n318), .A2(n289), .A3(n296), .ZN(n341) );
  OAI21_X1 U328 ( .B1(n293), .B2(n331), .A(n342), .ZN(n69) );
  OR3_X1 U329 ( .A1(n329), .A2(n289), .A3(n293), .ZN(n342) );
  XNOR2_X1 U330 ( .A(n343), .B(n344), .ZN(n38) );
  OR2_X1 U331 ( .A1(n343), .A2(n344), .ZN(n37) );
  OAI22_X1 U332 ( .A1(n315), .A2(n310), .B1(n284), .B2(n345), .ZN(n344) );
  XNOR2_X1 U333 ( .A(b[5]), .B(a[3]), .ZN(n315) );
  OAI22_X1 U334 ( .A1(n332), .A2(n331), .B1(n329), .B2(n333), .ZN(n343) );
  XNOR2_X1 U335 ( .A(b[2]), .B(a[7]), .ZN(n333) );
  XNOR2_X1 U336 ( .A(n222), .B(a[7]), .ZN(n332) );
  OAI22_X1 U337 ( .A1(n345), .A2(n310), .B1(n285), .B2(n317), .ZN(n31) );
  XNOR2_X1 U338 ( .A(b[7]), .B(a[3]), .ZN(n317) );
  XNOR2_X1 U339 ( .A(n299), .B(a[2]), .ZN(n346) );
  XNOR2_X1 U340 ( .A(b[6]), .B(a[3]), .ZN(n345) );
  OAI22_X1 U341 ( .A1(n326), .A2(n320), .B1(n318), .B2(n328), .ZN(n21) );
  XNOR2_X1 U342 ( .A(b[7]), .B(a[5]), .ZN(n328) );
  XNOR2_X1 U343 ( .A(n296), .B(a[4]), .ZN(n347) );
  XNOR2_X1 U344 ( .A(b[6]), .B(a[5]), .ZN(n326) );
  OAI22_X1 U345 ( .A1(n337), .A2(n331), .B1(n329), .B2(n339), .ZN(n15) );
  XNOR2_X1 U346 ( .A(b[7]), .B(a[7]), .ZN(n339) );
  NAND2_X1 U347 ( .A1(n329), .A2(n348), .ZN(n331) );
  XNOR2_X1 U348 ( .A(n293), .B(a[6]), .ZN(n348) );
  XNOR2_X1 U349 ( .A(b[6]), .B(a[7]), .ZN(n337) );
  OAI22_X1 U350 ( .A1(n289), .A2(n304), .B1(n349), .B2(n302), .ZN(n104) );
  OAI22_X1 U351 ( .A1(n349), .A2(n304), .B1(n350), .B2(n302), .ZN(n103) );
  XNOR2_X1 U352 ( .A(b[1]), .B(a[1]), .ZN(n349) );
  OAI22_X1 U353 ( .A1(n350), .A2(n304), .B1(n351), .B2(n302), .ZN(n102) );
  XNOR2_X1 U354 ( .A(b[2]), .B(a[1]), .ZN(n350) );
  OAI22_X1 U355 ( .A1(n351), .A2(n304), .B1(n352), .B2(n302), .ZN(n101) );
  XNOR2_X1 U356 ( .A(b[3]), .B(a[1]), .ZN(n351) );
  OAI22_X1 U357 ( .A1(n352), .A2(n304), .B1(n303), .B2(n302), .ZN(n100) );
  XNOR2_X1 U358 ( .A(b[5]), .B(a[1]), .ZN(n303) );
  NAND2_X1 U359 ( .A1(a[1]), .A2(n302), .ZN(n304) );
  XNOR2_X1 U360 ( .A(b[4]), .B(a[1]), .ZN(n352) );
endmodule


module datapath_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n77;
  wire   [15:1] carry;

  FA_X1 U1_14 ( .A(B[14]), .B(A[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  CLKBUF_X1 U1 ( .A(n6), .Z(n1) );
  CLKBUF_X1 U2 ( .A(n11), .Z(n2) );
  NAND3_X1 U3 ( .A1(n73), .A2(n74), .A3(n75), .ZN(n3) );
  NAND3_X1 U4 ( .A1(n47), .A2(n48), .A3(n49), .ZN(n4) );
  NAND3_X1 U5 ( .A1(n34), .A2(n35), .A3(n36), .ZN(n5) );
  NAND3_X1 U6 ( .A1(n38), .A2(n39), .A3(n40), .ZN(n6) );
  NAND3_X1 U7 ( .A1(n19), .A2(n20), .A3(n21), .ZN(n7) );
  NAND3_X1 U8 ( .A1(n19), .A2(n20), .A3(n21), .ZN(n8) );
  NAND3_X1 U9 ( .A1(n15), .A2(n16), .A3(n17), .ZN(n9) );
  NAND3_X1 U10 ( .A1(n15), .A2(n16), .A3(n17), .ZN(n10) );
  NAND3_X1 U11 ( .A1(n43), .A2(n44), .A3(n45), .ZN(n11) );
  CLKBUF_X1 U12 ( .A(n3), .Z(n12) );
  XNOR2_X1 U13 ( .A(carry[15]), .B(n13), .ZN(SUM[15]) );
  XNOR2_X1 U14 ( .A(B[15]), .B(A[15]), .ZN(n13) );
  XOR2_X1 U15 ( .A(A[1]), .B(B[1]), .Z(n14) );
  XOR2_X1 U16 ( .A(n14), .B(n77), .Z(SUM[1]) );
  NAND2_X1 U17 ( .A1(A[1]), .A2(B[1]), .ZN(n15) );
  NAND2_X1 U18 ( .A1(A[1]), .A2(n77), .ZN(n16) );
  NAND2_X1 U19 ( .A1(B[1]), .A2(n77), .ZN(n17) );
  NAND3_X1 U20 ( .A1(n15), .A2(n16), .A3(n17), .ZN(carry[2]) );
  XOR2_X1 U21 ( .A(B[2]), .B(A[2]), .Z(n18) );
  XOR2_X1 U22 ( .A(n18), .B(n10), .Z(SUM[2]) );
  NAND2_X1 U23 ( .A1(B[2]), .A2(A[2]), .ZN(n19) );
  NAND2_X1 U24 ( .A1(B[2]), .A2(n9), .ZN(n20) );
  NAND2_X1 U25 ( .A1(A[2]), .A2(carry[2]), .ZN(n21) );
  NAND3_X1 U26 ( .A1(n19), .A2(n20), .A3(n21), .ZN(carry[3]) );
  NAND3_X1 U27 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n22) );
  NAND3_X1 U28 ( .A1(n26), .A2(n27), .A3(n28), .ZN(n23) );
  NAND3_X1 U29 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n24) );
  XOR2_X1 U30 ( .A(B[3]), .B(A[3]), .Z(n25) );
  XOR2_X1 U31 ( .A(n8), .B(n25), .Z(SUM[3]) );
  NAND2_X1 U32 ( .A1(carry[3]), .A2(B[3]), .ZN(n26) );
  NAND2_X1 U33 ( .A1(n7), .A2(A[3]), .ZN(n27) );
  NAND2_X1 U34 ( .A1(B[3]), .A2(A[3]), .ZN(n28) );
  NAND3_X1 U35 ( .A1(n26), .A2(n27), .A3(n28), .ZN(carry[4]) );
  CLKBUF_X1 U36 ( .A(n64), .Z(n29) );
  CLKBUF_X1 U37 ( .A(carry[9]), .Z(n30) );
  NAND3_X1 U38 ( .A1(n56), .A2(n57), .A3(n58), .ZN(n31) );
  CLKBUF_X1 U39 ( .A(n24), .Z(n32) );
  XOR2_X1 U40 ( .A(B[12]), .B(A[12]), .Z(n33) );
  XOR2_X1 U41 ( .A(n2), .B(n33), .Z(SUM[12]) );
  NAND2_X1 U42 ( .A1(n11), .A2(B[12]), .ZN(n34) );
  NAND2_X1 U43 ( .A1(carry[12]), .A2(A[12]), .ZN(n35) );
  NAND2_X1 U44 ( .A1(B[12]), .A2(A[12]), .ZN(n36) );
  NAND3_X1 U45 ( .A1(n34), .A2(n35), .A3(n36), .ZN(carry[13]) );
  XOR2_X1 U46 ( .A(B[10]), .B(A[10]), .Z(n37) );
  XOR2_X1 U47 ( .A(n12), .B(n37), .Z(SUM[10]) );
  NAND2_X1 U48 ( .A1(n3), .A2(B[10]), .ZN(n38) );
  NAND2_X1 U49 ( .A1(carry[10]), .A2(A[10]), .ZN(n39) );
  NAND2_X1 U50 ( .A1(B[10]), .A2(A[10]), .ZN(n40) );
  NAND3_X1 U51 ( .A1(n38), .A2(n39), .A3(n40), .ZN(carry[11]) );
  NAND3_X1 U52 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n41) );
  XOR2_X1 U53 ( .A(B[11]), .B(A[11]), .Z(n42) );
  XOR2_X1 U54 ( .A(n1), .B(n42), .Z(SUM[11]) );
  NAND2_X1 U55 ( .A1(n6), .A2(B[11]), .ZN(n43) );
  NAND2_X1 U56 ( .A1(carry[11]), .A2(A[11]), .ZN(n44) );
  NAND2_X1 U57 ( .A1(B[11]), .A2(A[11]), .ZN(n45) );
  NAND3_X1 U58 ( .A1(n44), .A2(n43), .A3(n45), .ZN(carry[12]) );
  XOR2_X1 U59 ( .A(B[4]), .B(A[4]), .Z(n46) );
  XOR2_X1 U60 ( .A(carry[4]), .B(n46), .Z(SUM[4]) );
  NAND2_X1 U61 ( .A1(n23), .A2(B[4]), .ZN(n47) );
  NAND2_X1 U62 ( .A1(n23), .A2(A[4]), .ZN(n48) );
  NAND2_X1 U63 ( .A1(B[4]), .A2(A[4]), .ZN(n49) );
  NAND3_X1 U64 ( .A1(n47), .A2(n48), .A3(n49), .ZN(carry[5]) );
  XOR2_X1 U65 ( .A(B[5]), .B(A[5]), .Z(n50) );
  XOR2_X1 U66 ( .A(n4), .B(n50), .Z(SUM[5]) );
  NAND2_X1 U67 ( .A1(n4), .A2(B[5]), .ZN(n51) );
  NAND2_X1 U68 ( .A1(carry[5]), .A2(A[5]), .ZN(n52) );
  NAND2_X1 U69 ( .A1(B[5]), .A2(A[5]), .ZN(n53) );
  NAND3_X1 U70 ( .A1(n52), .A2(n51), .A3(n53), .ZN(carry[6]) );
  CLKBUF_X1 U71 ( .A(n31), .Z(n54) );
  XOR2_X1 U72 ( .A(B[6]), .B(A[6]), .Z(n55) );
  XOR2_X1 U73 ( .A(n32), .B(n55), .Z(SUM[6]) );
  NAND2_X1 U74 ( .A1(n24), .A2(B[6]), .ZN(n56) );
  NAND2_X1 U75 ( .A1(carry[6]), .A2(A[6]), .ZN(n57) );
  NAND2_X1 U76 ( .A1(B[6]), .A2(A[6]), .ZN(n58) );
  NAND3_X1 U77 ( .A1(n56), .A2(n57), .A3(n58), .ZN(carry[7]) );
  XOR2_X1 U78 ( .A(B[13]), .B(A[13]), .Z(n59) );
  XOR2_X1 U79 ( .A(n5), .B(n59), .Z(SUM[13]) );
  NAND2_X1 U80 ( .A1(n5), .A2(B[13]), .ZN(n60) );
  NAND2_X1 U81 ( .A1(carry[13]), .A2(A[13]), .ZN(n61) );
  NAND2_X1 U82 ( .A1(B[13]), .A2(A[13]), .ZN(n62) );
  NAND3_X1 U83 ( .A1(n60), .A2(n61), .A3(n62), .ZN(carry[14]) );
  XOR2_X1 U84 ( .A(B[7]), .B(A[7]), .Z(n63) );
  XOR2_X1 U85 ( .A(n54), .B(n63), .Z(SUM[7]) );
  NAND2_X1 U86 ( .A1(n31), .A2(B[7]), .ZN(n64) );
  NAND2_X1 U87 ( .A1(carry[7]), .A2(A[7]), .ZN(n65) );
  NAND2_X1 U88 ( .A1(B[7]), .A2(A[7]), .ZN(n66) );
  NAND3_X1 U89 ( .A1(n29), .A2(n65), .A3(n66), .ZN(carry[8]) );
  NAND3_X1 U90 ( .A1(n70), .A2(n69), .A3(n71), .ZN(n67) );
  XOR2_X1 U91 ( .A(A[8]), .B(B[8]), .Z(n68) );
  XOR2_X1 U92 ( .A(n68), .B(carry[8]), .Z(SUM[8]) );
  NAND2_X1 U93 ( .A1(A[8]), .A2(B[8]), .ZN(n69) );
  NAND2_X1 U94 ( .A1(A[8]), .A2(n41), .ZN(n70) );
  NAND2_X1 U95 ( .A1(B[8]), .A2(n22), .ZN(n71) );
  NAND3_X1 U96 ( .A1(n71), .A2(n70), .A3(n69), .ZN(carry[9]) );
  XOR2_X1 U97 ( .A(A[9]), .B(B[9]), .Z(n72) );
  XOR2_X1 U98 ( .A(n72), .B(n30), .Z(SUM[9]) );
  NAND2_X1 U99 ( .A1(A[9]), .A2(B[9]), .ZN(n73) );
  NAND2_X1 U100 ( .A1(A[9]), .A2(n67), .ZN(n74) );
  NAND2_X1 U101 ( .A1(carry[9]), .A2(B[9]), .ZN(n75) );
  NAND3_X1 U102 ( .A1(n73), .A2(n74), .A3(n75), .ZN(carry[10]) );
  XOR2_X1 U103 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U104 ( .A1(B[0]), .A2(A[0]), .ZN(n77) );
endmodule


module datapath ( clk, data_in, addr_x, wr_en_x, addr_a1, addr_a2, addr_a3, 
        addr_a4, addr_a5, addr_a6, addr_a7, addr_a8, addr_a9, addr_a10, 
        addr_a11, addr_a12, addr_a13, addr_a14, addr_a15, addr_a16, addr_a17, 
        addr_a18, addr_a19, addr_a20, addr_a21, addr_a22, addr_a23, addr_a24, 
        addr_a25, addr_a26, addr_a27, addr_a28, addr_a29, addr_a30, addr_a31, 
        addr_a32, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6, 
        wr_en_a7, wr_en_a8, wr_en_a9, wr_en_a10, wr_en_a11, wr_en_a12, 
        wr_en_a13, wr_en_a14, wr_en_a15, wr_en_a16, wr_en_a17, wr_en_a18, 
        wr_en_a19, wr_en_a20, wr_en_a21, wr_en_a22, wr_en_a23, wr_en_a24, 
        wr_en_a25, wr_en_a26, wr_en_a27, wr_en_a28, wr_en_a29, wr_en_a30, 
        wr_en_a31, wr_en_a32, addr_y, wr_en_y, clear_acc, clc, clc1, data_out
 );
  input [7:0] data_in;
  input [4:0] addr_x;
  input [4:0] addr_a1;
  input [4:0] addr_a2;
  input [4:0] addr_a3;
  input [4:0] addr_a4;
  input [4:0] addr_a5;
  input [4:0] addr_a6;
  input [4:0] addr_a7;
  input [4:0] addr_a8;
  input [4:0] addr_a9;
  input [4:0] addr_a10;
  input [4:0] addr_a11;
  input [4:0] addr_a12;
  input [4:0] addr_a13;
  input [4:0] addr_a14;
  input [4:0] addr_a15;
  input [4:0] addr_a16;
  input [4:0] addr_a17;
  input [4:0] addr_a18;
  input [4:0] addr_a19;
  input [4:0] addr_a20;
  input [4:0] addr_a21;
  input [4:0] addr_a22;
  input [4:0] addr_a23;
  input [4:0] addr_a24;
  input [4:0] addr_a25;
  input [4:0] addr_a26;
  input [4:0] addr_a27;
  input [4:0] addr_a28;
  input [4:0] addr_a29;
  input [4:0] addr_a30;
  input [4:0] addr_a31;
  input [4:0] addr_a32;
  input [4:0] addr_y;
  output [15:0] data_out;
  input clk, wr_en_x, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5,
         wr_en_a6, wr_en_a7, wr_en_a8, wr_en_a9, wr_en_a10, wr_en_a11,
         wr_en_a12, wr_en_a13, wr_en_a14, wr_en_a15, wr_en_a16, wr_en_a17,
         wr_en_a18, wr_en_a19, wr_en_a20, wr_en_a21, wr_en_a22, wr_en_a23,
         wr_en_a24, wr_en_a25, wr_en_a26, wr_en_a27, wr_en_a28, wr_en_a29,
         wr_en_a30, wr_en_a31, wr_en_a32, wr_en_y, clear_acc, clc, clc1;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         \mul_out1[9] , \mul_out1[8] , \mul_out1[7] , \mul_out1[6] ,
         \mul_out1[5] , \mul_out1[4] , \mul_out1[3] , \mul_out1[2] ,
         \mul_out1[1] , \mul_out1[15] , \mul_out1[14] , \mul_out1[13] ,
         \mul_out1[12] , \mul_out1[11] , \mul_out1[10] , \mul_out1[0] ,
         \mul_out2[9] , \mul_out2[8] , \mul_out2[7] , \mul_out2[6] ,
         \mul_out2[5] , \mul_out2[4] , \mul_out2[3] , \mul_out2[2] ,
         \mul_out2[1] , \mul_out2[15] , \mul_out2[14] , \mul_out2[13] ,
         \mul_out2[12] , \mul_out2[11] , \mul_out2[10] , \mul_out2[0] ,
         \mul_out3[9] , \mul_out3[8] , \mul_out3[7] , \mul_out3[6] ,
         \mul_out3[5] , \mul_out3[4] , \mul_out3[3] , \mul_out3[2] ,
         \mul_out3[1] , \mul_out3[15] , \mul_out3[14] , \mul_out3[13] ,
         \mul_out3[12] , \mul_out3[11] , \mul_out3[10] , \mul_out3[0] ,
         \mul_out4[9] , \mul_out4[8] , \mul_out4[7] , \mul_out4[6] ,
         \mul_out4[5] , \mul_out4[4] , \mul_out4[3] , \mul_out4[2] ,
         \mul_out4[1] , \mul_out4[15] , \mul_out4[14] , \mul_out4[13] ,
         \mul_out4[12] , \mul_out4[11] , \mul_out4[10] , \mul_out4[0] ,
         \mul_out5[9] , \mul_out5[8] , \mul_out5[7] , \mul_out5[6] ,
         \mul_out5[5] , \mul_out5[4] , \mul_out5[3] , \mul_out5[2] ,
         \mul_out5[1] , \mul_out5[15] , \mul_out5[14] , \mul_out5[13] ,
         \mul_out5[12] , \mul_out5[11] , \mul_out5[10] , \mul_out5[0] ,
         \mul_out6[9] , \mul_out6[8] , \mul_out6[7] , \mul_out6[6] ,
         \mul_out6[5] , \mul_out6[4] , \mul_out6[3] , \mul_out6[2] ,
         \mul_out6[1] , \mul_out6[15] , \mul_out6[14] , \mul_out6[13] ,
         \mul_out6[12] , \mul_out6[11] , \mul_out6[10] , \mul_out6[0] ,
         \mul_out7[9] , \mul_out7[8] , \mul_out7[7] , \mul_out7[6] ,
         \mul_out7[5] , \mul_out7[4] , \mul_out7[3] , \mul_out7[2] ,
         \mul_out7[1] , \mul_out7[15] , \mul_out7[14] , \mul_out7[13] ,
         \mul_out7[12] , \mul_out7[11] , \mul_out7[10] , \mul_out7[0] ,
         \mul_out8[9] , \mul_out8[8] , \mul_out8[7] , \mul_out8[6] ,
         \mul_out8[5] , \mul_out8[4] , \mul_out8[3] , \mul_out8[2] ,
         \mul_out8[1] , \mul_out8[15] , \mul_out8[14] , \mul_out8[13] ,
         \mul_out8[12] , \mul_out8[11] , \mul_out8[10] , \mul_out8[0] ,
         \mul_out9[9] , \mul_out9[8] , \mul_out9[7] , \mul_out9[6] ,
         \mul_out9[5] , \mul_out9[4] , \mul_out9[3] , \mul_out9[2] ,
         \mul_out9[1] , \mul_out9[15] , \mul_out9[14] , \mul_out9[13] ,
         \mul_out9[12] , \mul_out9[11] , \mul_out9[10] , \mul_out9[0] ,
         \mul_out10[9] , \mul_out10[8] , \mul_out10[7] , \mul_out10[6] ,
         \mul_out10[5] , \mul_out10[4] , \mul_out10[3] , \mul_out10[2] ,
         \mul_out10[1] , \mul_out10[15] , \mul_out10[14] , \mul_out10[13] ,
         \mul_out10[12] , \mul_out10[11] , \mul_out10[10] , \mul_out10[0] ,
         \mul_out11[9] , \mul_out11[8] , \mul_out11[7] , \mul_out11[6] ,
         \mul_out11[5] , \mul_out11[4] , \mul_out11[3] , \mul_out11[2] ,
         \mul_out11[1] , \mul_out11[15] , \mul_out11[14] , \mul_out11[13] ,
         \mul_out11[12] , \mul_out11[11] , \mul_out11[10] , \mul_out11[0] ,
         \mul_out12[9] , \mul_out12[8] , \mul_out12[7] , \mul_out12[6] ,
         \mul_out12[5] , \mul_out12[4] , \mul_out12[3] , \mul_out12[2] ,
         \mul_out12[1] , \mul_out12[15] , \mul_out12[14] , \mul_out12[13] ,
         \mul_out12[12] , \mul_out12[11] , \mul_out12[10] , \mul_out12[0] ,
         \mul_out13[9] , \mul_out13[8] , \mul_out13[7] , \mul_out13[6] ,
         \mul_out13[5] , \mul_out13[4] , \mul_out13[3] , \mul_out13[2] ,
         \mul_out13[1] , \mul_out13[15] , \mul_out13[14] , \mul_out13[13] ,
         \mul_out13[12] , \mul_out13[11] , \mul_out13[10] , \mul_out13[0] ,
         \mul_out14[9] , \mul_out14[8] , \mul_out14[7] , \mul_out14[6] ,
         \mul_out14[5] , \mul_out14[4] , \mul_out14[3] , \mul_out14[2] ,
         \mul_out14[1] , \mul_out14[15] , \mul_out14[14] , \mul_out14[13] ,
         \mul_out14[12] , \mul_out14[11] , \mul_out14[10] , \mul_out14[0] ,
         \mul_out15[9] , \mul_out15[8] , \mul_out15[7] , \mul_out15[6] ,
         \mul_out15[5] , \mul_out15[4] , \mul_out15[3] , \mul_out15[2] ,
         \mul_out15[1] , \mul_out15[15] , \mul_out15[14] , \mul_out15[13] ,
         \mul_out15[12] , \mul_out15[11] , \mul_out15[10] , \mul_out15[0] ,
         \mul_out16[9] , \mul_out16[8] , \mul_out16[7] , \mul_out16[6] ,
         \mul_out16[5] , \mul_out16[4] , \mul_out16[3] , \mul_out16[2] ,
         \mul_out16[1] , \mul_out16[15] , \mul_out16[14] , \mul_out16[13] ,
         \mul_out16[12] , \mul_out16[11] , \mul_out16[10] , \mul_out16[0] ,
         \mul_out17[9] , \mul_out17[8] , \mul_out17[7] , \mul_out17[6] ,
         \mul_out17[5] , \mul_out17[4] , \mul_out17[3] , \mul_out17[2] ,
         \mul_out17[1] , \mul_out17[15] , \mul_out17[14] , \mul_out17[13] ,
         \mul_out17[12] , \mul_out17[11] , \mul_out17[10] , \mul_out17[0] ,
         \mul_out18[9] , \mul_out18[8] , \mul_out18[7] , \mul_out18[6] ,
         \mul_out18[5] , \mul_out18[4] , \mul_out18[3] , \mul_out18[2] ,
         \mul_out18[1] , \mul_out18[15] , \mul_out18[14] , \mul_out18[13] ,
         \mul_out18[12] , \mul_out18[11] , \mul_out18[10] , \mul_out18[0] ,
         \mul_out19[9] , \mul_out19[8] , \mul_out19[7] , \mul_out19[6] ,
         \mul_out19[5] , \mul_out19[4] , \mul_out19[3] , \mul_out19[2] ,
         \mul_out19[1] , \mul_out19[15] , \mul_out19[14] , \mul_out19[13] ,
         \mul_out19[12] , \mul_out19[11] , \mul_out19[10] , \mul_out19[0] ,
         \mul_out20[9] , \mul_out20[8] , \mul_out20[7] , \mul_out20[6] ,
         \mul_out20[5] , \mul_out20[4] , \mul_out20[3] , \mul_out20[2] ,
         \mul_out20[1] , \mul_out20[15] , \mul_out20[14] , \mul_out20[13] ,
         \mul_out20[12] , \mul_out20[11] , \mul_out20[10] , \mul_out20[0] ,
         \mul_out21[9] , \mul_out21[8] , \mul_out21[7] , \mul_out21[6] ,
         \mul_out21[5] , \mul_out21[4] , \mul_out21[3] , \mul_out21[2] ,
         \mul_out21[1] , \mul_out21[15] , \mul_out21[14] , \mul_out21[13] ,
         \mul_out21[12] , \mul_out21[11] , \mul_out21[10] , \mul_out21[0] ,
         \mul_out22[9] , \mul_out22[8] , \mul_out22[7] , \mul_out22[6] ,
         \mul_out22[5] , \mul_out22[4] , \mul_out22[3] , \mul_out22[2] ,
         \mul_out22[1] , \mul_out22[15] , \mul_out22[14] , \mul_out22[13] ,
         \mul_out22[12] , \mul_out22[11] , \mul_out22[10] , \mul_out22[0] ,
         \mul_out23[9] , \mul_out23[8] , \mul_out23[7] , \mul_out23[6] ,
         \mul_out23[5] , \mul_out23[4] , \mul_out23[3] , \mul_out23[2] ,
         \mul_out23[1] , \mul_out23[15] , \mul_out23[14] , \mul_out23[13] ,
         \mul_out23[12] , \mul_out23[11] , \mul_out23[10] , \mul_out23[0] ,
         \mul_out24[9] , \mul_out24[8] , \mul_out24[7] , \mul_out24[6] ,
         \mul_out24[5] , \mul_out24[4] , \mul_out24[3] , \mul_out24[2] ,
         \mul_out24[1] , \mul_out24[15] , \mul_out24[14] , \mul_out24[13] ,
         \mul_out24[12] , \mul_out24[11] , \mul_out24[10] , \mul_out24[0] ,
         \mul_out25[9] , \mul_out25[8] , \mul_out25[7] , \mul_out25[6] ,
         \mul_out25[5] , \mul_out25[4] , \mul_out25[3] , \mul_out25[2] ,
         \mul_out25[1] , \mul_out25[15] , \mul_out25[14] , \mul_out25[13] ,
         \mul_out25[12] , \mul_out25[11] , \mul_out25[10] , \mul_out25[0] ,
         \mul_out26[9] , \mul_out26[8] , \mul_out26[7] , \mul_out26[6] ,
         \mul_out26[5] , \mul_out26[4] , \mul_out26[3] , \mul_out26[2] ,
         \mul_out26[1] , \mul_out26[15] , \mul_out26[14] , \mul_out26[13] ,
         \mul_out26[12] , \mul_out26[11] , \mul_out26[10] , \mul_out26[0] ,
         \mul_out27[9] , \mul_out27[8] , \mul_out27[7] , \mul_out27[6] ,
         \mul_out27[5] , \mul_out27[4] , \mul_out27[3] , \mul_out27[2] ,
         \mul_out27[1] , \mul_out27[15] , \mul_out27[14] , \mul_out27[13] ,
         \mul_out27[12] , \mul_out27[11] , \mul_out27[10] , \mul_out27[0] ,
         \mul_out28[9] , \mul_out28[8] , \mul_out28[7] , \mul_out28[6] ,
         \mul_out28[5] , \mul_out28[4] , \mul_out28[3] , \mul_out28[2] ,
         \mul_out28[1] , \mul_out28[15] , \mul_out28[14] , \mul_out28[13] ,
         \mul_out28[12] , \mul_out28[11] , \mul_out28[10] , \mul_out28[0] ,
         \mul_out29[9] , \mul_out29[8] , \mul_out29[7] , \mul_out29[6] ,
         \mul_out29[5] , \mul_out29[4] , \mul_out29[3] , \mul_out29[2] ,
         \mul_out29[1] , \mul_out29[15] , \mul_out29[14] , \mul_out29[13] ,
         \mul_out29[12] , \mul_out29[11] , \mul_out29[10] , \mul_out29[0] ,
         \mul_out30[9] , \mul_out30[8] , \mul_out30[7] , \mul_out30[6] ,
         \mul_out30[5] , \mul_out30[4] , \mul_out30[3] , \mul_out30[2] ,
         \mul_out30[1] , \mul_out30[15] , \mul_out30[14] , \mul_out30[13] ,
         \mul_out30[12] , \mul_out30[11] , \mul_out30[10] , \mul_out30[0] ,
         \mul_out31[9] , \mul_out31[8] , \mul_out31[7] , \mul_out31[6] ,
         \mul_out31[5] , \mul_out31[4] , \mul_out31[3] , \mul_out31[2] ,
         \mul_out31[1] , \mul_out31[15] , \mul_out31[14] , \mul_out31[13] ,
         \mul_out31[12] , \mul_out31[11] , \mul_out31[10] , \mul_out31[0] ,
         \mul_out32[9] , \mul_out32[8] , \mul_out32[7] , \mul_out32[6] ,
         \mul_out32[5] , \mul_out32[4] , \mul_out32[3] , \mul_out32[2] ,
         \mul_out32[1] , \mul_out32[15] , \mul_out32[14] , \mul_out32[13] ,
         \mul_out32[12] , \mul_out32[11] , \mul_out32[10] , \mul_out32[0] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171;
  wire   [7:0] data_out_x;
  wire   [7:0] data_out_a1;
  wire   [7:0] data_out_a2;
  wire   [7:0] data_out_a3;
  wire   [7:0] data_out_a4;
  wire   [7:0] data_out_a5;
  wire   [7:0] data_out_a6;
  wire   [7:0] data_out_a7;
  wire   [7:0] data_out_a8;
  wire   [7:0] data_out_a9;
  wire   [7:0] data_out_a10;
  wire   [7:0] data_out_a11;
  wire   [7:0] data_out_a12;
  wire   [7:0] data_out_a13;
  wire   [7:0] data_out_a14;
  wire   [7:0] data_out_a15;
  wire   [7:0] data_out_a16;
  wire   [7:0] data_out_a17;
  wire   [7:0] data_out_a18;
  wire   [7:0] data_out_a19;
  wire   [7:0] data_out_a20;
  wire   [7:0] data_out_a21;
  wire   [7:0] data_out_a22;
  wire   [7:0] data_out_a23;
  wire   [7:0] data_out_a24;
  wire   [7:0] data_out_a25;
  wire   [7:0] data_out_a26;
  wire   [7:0] data_out_a27;
  wire   [7:0] data_out_a28;
  wire   [7:0] data_out_a29;
  wire   [7:0] data_out_a30;
  wire   [7:0] data_out_a31;
  wire   [7:0] data_out_a32;
  wire   [15:0] f;
  wire   [15:0] f1;
  wire   [15:0] f2;
  wire   [15:0] f3;
  wire   [15:0] f4;
  wire   [15:0] f5;
  wire   [15:0] f6;
  wire   [15:0] f7;
  wire   [15:0] f8;
  wire   [15:0] f9;
  wire   [15:0] f10;
  wire   [15:0] f11;
  wire   [15:0] f12;
  wire   [15:0] f13;
  wire   [15:0] f14;
  wire   [15:0] f15;
  wire   [15:0] f16;
  wire   [15:0] f17;
  wire   [15:0] f18;
  wire   [15:0] f19;
  wire   [15:0] f20;
  wire   [15:0] f21;
  wire   [15:0] f22;
  wire   [15:0] f23;
  wire   [15:0] f24;
  wire   [15:0] f25;
  wire   [15:0] f26;
  wire   [15:0] f27;
  wire   [15:0] f28;
  wire   [15:0] f29;
  wire   [15:0] f30;
  wire   [15:0] f31;
  wire   [15:0] f32;
  wire   [15:0] add_r1;
  wire   [15:0] add_r2;
  wire   [15:0] add_r3;
  wire   [15:0] add_r4;
  wire   [15:0] add_r5;
  wire   [15:0] add_r6;
  wire   [15:0] add_r7;
  wire   [15:0] add_r8;
  wire   [15:0] add_r9;
  wire   [15:0] add_r10;
  wire   [15:0] add_r11;
  wire   [15:0] add_r12;
  wire   [15:0] add_r13;
  wire   [15:0] add_r14;
  wire   [15:0] add_r15;
  wire   [15:0] add_r16;
  wire   [15:0] add_r17;
  wire   [15:0] add_r18;
  wire   [15:0] add_r19;
  wire   [15:0] add_r20;
  wire   [15:0] add_r21;
  wire   [15:0] add_r22;
  wire   [15:0] add_r23;
  wire   [15:0] add_r24;
  wire   [15:0] add_r25;
  wire   [15:0] add_r26;
  wire   [15:0] add_r27;
  wire   [15:0] add_r28;
  wire   [15:0] add_r29;
  wire   [15:0] add_r30;
  wire   [15:0] add_r31;
  wire   [15:0] add_r32;

  DFF_X1 \f1_reg[15]  ( .D(n2026), .CK(clk), .Q(f1[15]), .QN(n33) );
  DFF_X1 \f1_reg[14]  ( .D(n2025), .CK(clk), .Q(f1[14]), .QN(n34) );
  DFF_X1 \f1_reg[13]  ( .D(n2024), .CK(clk), .Q(f1[13]), .QN(n35) );
  DFF_X1 \f1_reg[12]  ( .D(n2023), .CK(clk), .Q(f1[12]), .QN(n36) );
  DFF_X1 \f1_reg[11]  ( .D(n2022), .CK(clk), .Q(f1[11]), .QN(n37) );
  DFF_X1 \f1_reg[10]  ( .D(n2021), .CK(clk), .Q(f1[10]), .QN(n38) );
  DFF_X1 \f1_reg[9]  ( .D(n2020), .CK(clk), .Q(f1[9]), .QN(n39) );
  DFF_X1 \f1_reg[8]  ( .D(n2019), .CK(clk), .Q(f1[8]), .QN(n40) );
  DFF_X1 \f1_reg[7]  ( .D(n2018), .CK(clk), .Q(f1[7]), .QN(n41) );
  DFF_X1 \f1_reg[6]  ( .D(n2017), .CK(clk), .Q(f1[6]), .QN(n42) );
  DFF_X1 \f1_reg[5]  ( .D(n2016), .CK(clk), .Q(f1[5]), .QN(n43) );
  DFF_X1 \f1_reg[4]  ( .D(n2015), .CK(clk), .Q(f1[4]), .QN(n44) );
  DFF_X1 \f1_reg[3]  ( .D(n2014), .CK(clk), .Q(f1[3]), .QN(n45) );
  DFF_X1 \f1_reg[2]  ( .D(n2013), .CK(clk), .Q(f1[2]), .QN(n46) );
  DFF_X1 \f1_reg[1]  ( .D(n2012), .CK(clk), .Q(f1[1]), .QN(n47) );
  DFF_X1 \f1_reg[0]  ( .D(n2011), .CK(clk), .Q(f1[0]), .QN(n48) );
  DFF_X1 \f2_reg[14]  ( .D(n2009), .CK(clk), .Q(f2[14]), .QN(n50) );
  DFF_X1 \f2_reg[13]  ( .D(n2008), .CK(clk), .Q(f2[13]), .QN(n51) );
  DFF_X1 \f2_reg[12]  ( .D(n2007), .CK(clk), .Q(f2[12]), .QN(n52) );
  DFF_X1 \f2_reg[11]  ( .D(n2006), .CK(clk), .Q(f2[11]), .QN(n53) );
  DFF_X1 \f2_reg[10]  ( .D(n2005), .CK(clk), .Q(f2[10]), .QN(n54) );
  DFF_X1 \f2_reg[9]  ( .D(n2004), .CK(clk), .Q(f2[9]), .QN(n55) );
  DFF_X1 \f2_reg[8]  ( .D(n2003), .CK(clk), .Q(f2[8]), .QN(n56) );
  DFF_X1 \f2_reg[7]  ( .D(n2002), .CK(clk), .Q(f2[7]), .QN(n57) );
  DFF_X1 \f2_reg[6]  ( .D(n2001), .CK(clk), .Q(f2[6]), .QN(n58) );
  DFF_X1 \f2_reg[5]  ( .D(n2000), .CK(clk), .Q(f2[5]), .QN(n59) );
  DFF_X1 \f2_reg[4]  ( .D(n1999), .CK(clk), .Q(f2[4]), .QN(n60) );
  DFF_X1 \f2_reg[3]  ( .D(n1998), .CK(clk), .Q(f2[3]), .QN(n61) );
  DFF_X1 \f2_reg[2]  ( .D(n1997), .CK(clk), .Q(f2[2]), .QN(n62) );
  DFF_X1 \f2_reg[1]  ( .D(n1996), .CK(clk), .Q(f2[1]), .QN(n63) );
  DFF_X1 \f2_reg[0]  ( .D(n1995), .CK(clk), .Q(f2[0]), .QN(n64) );
  DFF_X1 \f3_reg[14]  ( .D(n1993), .CK(clk), .Q(f3[14]), .QN(n66) );
  DFF_X1 \f3_reg[13]  ( .D(n1992), .CK(clk), .Q(f3[13]), .QN(n67) );
  DFF_X1 \f3_reg[12]  ( .D(n1991), .CK(clk), .Q(f3[12]), .QN(n68) );
  DFF_X1 \f3_reg[11]  ( .D(n1990), .CK(clk), .Q(f3[11]), .QN(n69) );
  DFF_X1 \f3_reg[10]  ( .D(n1989), .CK(clk), .Q(f3[10]), .QN(n70) );
  DFF_X1 \f3_reg[9]  ( .D(n1988), .CK(clk), .Q(f3[9]), .QN(n71) );
  DFF_X1 \f3_reg[8]  ( .D(n1987), .CK(clk), .Q(f3[8]), .QN(n72) );
  DFF_X1 \f3_reg[7]  ( .D(n1986), .CK(clk), .Q(f3[7]), .QN(n73) );
  DFF_X1 \f3_reg[6]  ( .D(n1985), .CK(clk), .Q(f3[6]), .QN(n74) );
  DFF_X1 \f3_reg[5]  ( .D(n1984), .CK(clk), .Q(f3[5]), .QN(n75) );
  DFF_X1 \f3_reg[4]  ( .D(n1983), .CK(clk), .Q(f3[4]), .QN(n76) );
  DFF_X1 \f3_reg[3]  ( .D(n1982), .CK(clk), .Q(f3[3]), .QN(n77) );
  DFF_X1 \f3_reg[2]  ( .D(n1981), .CK(clk), .Q(f3[2]), .QN(n78) );
  DFF_X1 \f3_reg[1]  ( .D(n1980), .CK(clk), .Q(f3[1]), .QN(n79) );
  DFF_X1 \f3_reg[0]  ( .D(n1979), .CK(clk), .Q(f3[0]), .QN(n80) );
  DFF_X1 \f4_reg[15]  ( .D(n1978), .CK(clk), .Q(f4[15]), .QN(n81) );
  DFF_X1 \f4_reg[14]  ( .D(n1977), .CK(clk), .Q(f4[14]), .QN(n82) );
  DFF_X1 \f4_reg[13]  ( .D(n1976), .CK(clk), .Q(f4[13]), .QN(n83) );
  DFF_X1 \f4_reg[12]  ( .D(n1975), .CK(clk), .Q(f4[12]), .QN(n84) );
  DFF_X1 \f4_reg[11]  ( .D(n1974), .CK(clk), .Q(f4[11]), .QN(n85) );
  DFF_X1 \f4_reg[10]  ( .D(n1973), .CK(clk), .Q(f4[10]), .QN(n86) );
  DFF_X1 \f4_reg[9]  ( .D(n1972), .CK(clk), .Q(f4[9]), .QN(n87) );
  DFF_X1 \f4_reg[8]  ( .D(n1971), .CK(clk), .Q(f4[8]), .QN(n88) );
  DFF_X1 \f4_reg[7]  ( .D(n1970), .CK(clk), .Q(f4[7]), .QN(n89) );
  DFF_X1 \f4_reg[6]  ( .D(n1969), .CK(clk), .Q(f4[6]), .QN(n90) );
  DFF_X1 \f4_reg[5]  ( .D(n1968), .CK(clk), .Q(f4[5]), .QN(n91) );
  DFF_X1 \f4_reg[4]  ( .D(n1967), .CK(clk), .Q(f4[4]), .QN(n92) );
  DFF_X1 \f4_reg[3]  ( .D(n1966), .CK(clk), .Q(f4[3]), .QN(n93) );
  DFF_X1 \f4_reg[2]  ( .D(n1965), .CK(clk), .Q(f4[2]), .QN(n94) );
  DFF_X1 \f4_reg[1]  ( .D(n1964), .CK(clk), .Q(f4[1]), .QN(n95) );
  DFF_X1 \f4_reg[0]  ( .D(n1963), .CK(clk), .Q(f4[0]), .QN(n96) );
  DFF_X1 \f5_reg[14]  ( .D(n1961), .CK(clk), .Q(f5[14]), .QN(n98) );
  DFF_X1 \f5_reg[13]  ( .D(n1960), .CK(clk), .Q(f5[13]), .QN(n99) );
  DFF_X1 \f5_reg[12]  ( .D(n1959), .CK(clk), .Q(f5[12]), .QN(n100) );
  DFF_X1 \f5_reg[11]  ( .D(n1958), .CK(clk), .Q(f5[11]), .QN(n101) );
  DFF_X1 \f5_reg[10]  ( .D(n1957), .CK(clk), .Q(f5[10]), .QN(n102) );
  DFF_X1 \f5_reg[9]  ( .D(n1956), .CK(clk), .Q(f5[9]), .QN(n103) );
  DFF_X1 \f5_reg[8]  ( .D(n1955), .CK(clk), .Q(f5[8]), .QN(n104) );
  DFF_X1 \f5_reg[7]  ( .D(n1954), .CK(clk), .Q(f5[7]), .QN(n105) );
  DFF_X1 \f5_reg[6]  ( .D(n1953), .CK(clk), .Q(f5[6]), .QN(n106) );
  DFF_X1 \f5_reg[5]  ( .D(n1952), .CK(clk), .Q(f5[5]), .QN(n107) );
  DFF_X1 \f5_reg[4]  ( .D(n1951), .CK(clk), .Q(f5[4]), .QN(n108) );
  DFF_X1 \f5_reg[3]  ( .D(n1950), .CK(clk), .Q(f5[3]), .QN(n109) );
  DFF_X1 \f5_reg[2]  ( .D(n1949), .CK(clk), .Q(f5[2]), .QN(n110) );
  DFF_X1 \f5_reg[1]  ( .D(n1948), .CK(clk), .Q(f5[1]), .QN(n111) );
  DFF_X1 \f5_reg[0]  ( .D(n1947), .CK(clk), .Q(f5[0]), .QN(n112) );
  DFF_X1 \f6_reg[14]  ( .D(n1945), .CK(clk), .Q(f6[14]), .QN(n114) );
  DFF_X1 \f6_reg[13]  ( .D(n1944), .CK(clk), .Q(f6[13]), .QN(n115) );
  DFF_X1 \f6_reg[12]  ( .D(n1943), .CK(clk), .Q(f6[12]), .QN(n116) );
  DFF_X1 \f6_reg[11]  ( .D(n1942), .CK(clk), .Q(f6[11]), .QN(n117) );
  DFF_X1 \f6_reg[10]  ( .D(n1941), .CK(clk), .Q(f6[10]), .QN(n118) );
  DFF_X1 \f6_reg[9]  ( .D(n1940), .CK(clk), .Q(f6[9]), .QN(n119) );
  DFF_X1 \f6_reg[8]  ( .D(n1939), .CK(clk), .Q(f6[8]), .QN(n120) );
  DFF_X1 \f6_reg[7]  ( .D(n1938), .CK(clk), .Q(f6[7]), .QN(n121) );
  DFF_X1 \f6_reg[6]  ( .D(n1937), .CK(clk), .Q(f6[6]), .QN(n122) );
  DFF_X1 \f6_reg[5]  ( .D(n1936), .CK(clk), .Q(f6[5]), .QN(n123) );
  DFF_X1 \f6_reg[4]  ( .D(n1935), .CK(clk), .Q(f6[4]), .QN(n124) );
  DFF_X1 \f6_reg[3]  ( .D(n1934), .CK(clk), .Q(f6[3]), .QN(n125) );
  DFF_X1 \f6_reg[2]  ( .D(n1933), .CK(clk), .Q(f6[2]), .QN(n126) );
  DFF_X1 \f6_reg[1]  ( .D(n1932), .CK(clk), .Q(f6[1]), .QN(n127) );
  DFF_X1 \f6_reg[0]  ( .D(n1931), .CK(clk), .Q(f6[0]), .QN(n128) );
  DFF_X1 \f7_reg[14]  ( .D(n1929), .CK(clk), .Q(f7[14]), .QN(n130) );
  DFF_X1 \f7_reg[13]  ( .D(n1928), .CK(clk), .Q(f7[13]), .QN(n131) );
  DFF_X1 \f7_reg[12]  ( .D(n1927), .CK(clk), .Q(f7[12]), .QN(n132) );
  DFF_X1 \f7_reg[11]  ( .D(n1926), .CK(clk), .Q(f7[11]), .QN(n133) );
  DFF_X1 \f7_reg[10]  ( .D(n1925), .CK(clk), .Q(f7[10]), .QN(n134) );
  DFF_X1 \f7_reg[9]  ( .D(n1924), .CK(clk), .Q(f7[9]), .QN(n135) );
  DFF_X1 \f7_reg[8]  ( .D(n1923), .CK(clk), .Q(f7[8]), .QN(n136) );
  DFF_X1 \f7_reg[7]  ( .D(n1922), .CK(clk), .Q(f7[7]), .QN(n137) );
  DFF_X1 \f7_reg[6]  ( .D(n1921), .CK(clk), .Q(f7[6]), .QN(n138) );
  DFF_X1 \f7_reg[5]  ( .D(n1920), .CK(clk), .Q(f7[5]), .QN(n139) );
  DFF_X1 \f7_reg[4]  ( .D(n1919), .CK(clk), .Q(f7[4]), .QN(n140) );
  DFF_X1 \f7_reg[3]  ( .D(n1918), .CK(clk), .Q(f7[3]), .QN(n141) );
  DFF_X1 \f7_reg[2]  ( .D(n1917), .CK(clk), .Q(f7[2]), .QN(n142) );
  DFF_X1 \f7_reg[1]  ( .D(n1916), .CK(clk), .Q(f7[1]), .QN(n143) );
  DFF_X1 \f7_reg[0]  ( .D(n1915), .CK(clk), .Q(f7[0]), .QN(n144) );
  DFF_X1 \f8_reg[15]  ( .D(n1914), .CK(clk), .Q(f8[15]), .QN(n145) );
  DFF_X1 \f8_reg[14]  ( .D(n1913), .CK(clk), .Q(f8[14]), .QN(n146) );
  DFF_X1 \f8_reg[13]  ( .D(n1912), .CK(clk), .Q(f8[13]), .QN(n147) );
  DFF_X1 \f8_reg[12]  ( .D(n1911), .CK(clk), .Q(f8[12]), .QN(n148) );
  DFF_X1 \f8_reg[11]  ( .D(n1910), .CK(clk), .Q(f8[11]), .QN(n149) );
  DFF_X1 \f8_reg[10]  ( .D(n1909), .CK(clk), .Q(f8[10]), .QN(n150) );
  DFF_X1 \f8_reg[9]  ( .D(n1908), .CK(clk), .Q(f8[9]), .QN(n151) );
  DFF_X1 \f8_reg[8]  ( .D(n1907), .CK(clk), .Q(f8[8]), .QN(n152) );
  DFF_X1 \f8_reg[7]  ( .D(n1906), .CK(clk), .Q(f8[7]), .QN(n153) );
  DFF_X1 \f8_reg[6]  ( .D(n1905), .CK(clk), .Q(f8[6]), .QN(n154) );
  DFF_X1 \f8_reg[5]  ( .D(n1904), .CK(clk), .Q(f8[5]), .QN(n155) );
  DFF_X1 \f8_reg[4]  ( .D(n1903), .CK(clk), .Q(f8[4]), .QN(n156) );
  DFF_X1 \f8_reg[3]  ( .D(n1902), .CK(clk), .Q(f8[3]), .QN(n157) );
  DFF_X1 \f8_reg[2]  ( .D(n1901), .CK(clk), .Q(f8[2]), .QN(n158) );
  DFF_X1 \f8_reg[1]  ( .D(n1900), .CK(clk), .Q(f8[1]), .QN(n159) );
  DFF_X1 \f8_reg[0]  ( .D(n1899), .CK(clk), .Q(f8[0]), .QN(n160) );
  DFF_X1 \f9_reg[14]  ( .D(n1897), .CK(clk), .Q(f9[14]), .QN(n162) );
  DFF_X1 \f9_reg[13]  ( .D(n1896), .CK(clk), .Q(f9[13]), .QN(n163) );
  DFF_X1 \f9_reg[12]  ( .D(n1895), .CK(clk), .Q(f9[12]), .QN(n164) );
  DFF_X1 \f9_reg[11]  ( .D(n1894), .CK(clk), .Q(f9[11]), .QN(n165) );
  DFF_X1 \f9_reg[10]  ( .D(n1893), .CK(clk), .Q(f9[10]), .QN(n166) );
  DFF_X1 \f9_reg[9]  ( .D(n1892), .CK(clk), .Q(f9[9]), .QN(n167) );
  DFF_X1 \f9_reg[8]  ( .D(n1891), .CK(clk), .Q(f9[8]), .QN(n168) );
  DFF_X1 \f9_reg[7]  ( .D(n1890), .CK(clk), .Q(f9[7]), .QN(n169) );
  DFF_X1 \f9_reg[6]  ( .D(n1889), .CK(clk), .Q(f9[6]), .QN(n170) );
  DFF_X1 \f9_reg[5]  ( .D(n1888), .CK(clk), .Q(f9[5]), .QN(n171) );
  DFF_X1 \f9_reg[4]  ( .D(n1887), .CK(clk), .Q(f9[4]), .QN(n172) );
  DFF_X1 \f9_reg[3]  ( .D(n1886), .CK(clk), .Q(f9[3]), .QN(n173) );
  DFF_X1 \f9_reg[2]  ( .D(n1885), .CK(clk), .Q(f9[2]), .QN(n174) );
  DFF_X1 \f9_reg[1]  ( .D(n1884), .CK(clk), .Q(f9[1]), .QN(n175) );
  DFF_X1 \f9_reg[0]  ( .D(n1883), .CK(clk), .Q(f9[0]), .QN(n176) );
  DFF_X1 \f10_reg[14]  ( .D(n1881), .CK(clk), .Q(f10[14]), .QN(n178) );
  DFF_X1 \f10_reg[13]  ( .D(n1880), .CK(clk), .Q(f10[13]), .QN(n179) );
  DFF_X1 \f10_reg[12]  ( .D(n1879), .CK(clk), .Q(f10[12]), .QN(n180) );
  DFF_X1 \f10_reg[11]  ( .D(n1878), .CK(clk), .Q(f10[11]), .QN(n181) );
  DFF_X1 \f10_reg[10]  ( .D(n1877), .CK(clk), .Q(f10[10]), .QN(n182) );
  DFF_X1 \f10_reg[9]  ( .D(n1876), .CK(clk), .Q(f10[9]), .QN(n183) );
  DFF_X1 \f10_reg[8]  ( .D(n1875), .CK(clk), .Q(f10[8]), .QN(n184) );
  DFF_X1 \f10_reg[7]  ( .D(n1874), .CK(clk), .Q(f10[7]), .QN(n185) );
  DFF_X1 \f10_reg[6]  ( .D(n1873), .CK(clk), .Q(f10[6]), .QN(n186) );
  DFF_X1 \f10_reg[5]  ( .D(n1872), .CK(clk), .Q(f10[5]), .QN(n187) );
  DFF_X1 \f10_reg[4]  ( .D(n1871), .CK(clk), .Q(f10[4]), .QN(n188) );
  DFF_X1 \f10_reg[3]  ( .D(n1870), .CK(clk), .Q(f10[3]), .QN(n189) );
  DFF_X1 \f10_reg[2]  ( .D(n1869), .CK(clk), .Q(f10[2]), .QN(n190) );
  DFF_X1 \f10_reg[1]  ( .D(n1868), .CK(clk), .Q(f10[1]), .QN(n191) );
  DFF_X1 \f10_reg[0]  ( .D(n1867), .CK(clk), .Q(f10[0]), .QN(n192) );
  DFF_X1 \f11_reg[15]  ( .D(n1866), .CK(clk), .Q(f11[15]), .QN(n193) );
  DFF_X1 \f11_reg[14]  ( .D(n1865), .CK(clk), .Q(f11[14]), .QN(n194) );
  DFF_X1 \f11_reg[13]  ( .D(n1864), .CK(clk), .Q(f11[13]), .QN(n195) );
  DFF_X1 \f11_reg[12]  ( .D(n1863), .CK(clk), .Q(f11[12]), .QN(n196) );
  DFF_X1 \f11_reg[11]  ( .D(n1862), .CK(clk), .Q(f11[11]), .QN(n197) );
  DFF_X1 \f11_reg[10]  ( .D(n1861), .CK(clk), .Q(f11[10]), .QN(n198) );
  DFF_X1 \f11_reg[9]  ( .D(n1860), .CK(clk), .Q(f11[9]), .QN(n199) );
  DFF_X1 \f11_reg[8]  ( .D(n1859), .CK(clk), .Q(f11[8]), .QN(n200) );
  DFF_X1 \f11_reg[7]  ( .D(n1858), .CK(clk), .Q(f11[7]), .QN(n201) );
  DFF_X1 \f11_reg[6]  ( .D(n1857), .CK(clk), .Q(f11[6]), .QN(n202) );
  DFF_X1 \f11_reg[5]  ( .D(n1856), .CK(clk), .Q(f11[5]), .QN(n203) );
  DFF_X1 \f11_reg[4]  ( .D(n1855), .CK(clk), .Q(f11[4]), .QN(n204) );
  DFF_X1 \f11_reg[3]  ( .D(n1854), .CK(clk), .Q(f11[3]), .QN(n205) );
  DFF_X1 \f11_reg[2]  ( .D(n1853), .CK(clk), .Q(f11[2]), .QN(n206) );
  DFF_X1 \f11_reg[1]  ( .D(n1852), .CK(clk), .Q(f11[1]), .QN(n207) );
  DFF_X1 \f11_reg[0]  ( .D(n1851), .CK(clk), .Q(f11[0]), .QN(n208) );
  DFF_X1 \f12_reg[14]  ( .D(n1849), .CK(clk), .Q(f12[14]), .QN(n210) );
  DFF_X1 \f12_reg[13]  ( .D(n1848), .CK(clk), .Q(f12[13]), .QN(n211) );
  DFF_X1 \f12_reg[12]  ( .D(n1847), .CK(clk), .Q(f12[12]), .QN(n212) );
  DFF_X1 \f12_reg[11]  ( .D(n1846), .CK(clk), .Q(f12[11]), .QN(n213) );
  DFF_X1 \f12_reg[10]  ( .D(n1845), .CK(clk), .Q(f12[10]), .QN(n214) );
  DFF_X1 \f12_reg[9]  ( .D(n1844), .CK(clk), .Q(f12[9]), .QN(n215) );
  DFF_X1 \f12_reg[8]  ( .D(n1843), .CK(clk), .Q(f12[8]), .QN(n216) );
  DFF_X1 \f12_reg[7]  ( .D(n1842), .CK(clk), .Q(f12[7]), .QN(n217) );
  DFF_X1 \f12_reg[6]  ( .D(n1841), .CK(clk), .Q(f12[6]), .QN(n218) );
  DFF_X1 \f12_reg[5]  ( .D(n1840), .CK(clk), .Q(f12[5]), .QN(n219) );
  DFF_X1 \f12_reg[4]  ( .D(n1839), .CK(clk), .Q(f12[4]), .QN(n220) );
  DFF_X1 \f12_reg[3]  ( .D(n1838), .CK(clk), .Q(f12[3]), .QN(n221) );
  DFF_X1 \f12_reg[2]  ( .D(n1837), .CK(clk), .Q(f12[2]), .QN(n222) );
  DFF_X1 \f12_reg[1]  ( .D(n1836), .CK(clk), .Q(f12[1]), .QN(n223) );
  DFF_X1 \f12_reg[0]  ( .D(n1835), .CK(clk), .Q(f12[0]), .QN(n224) );
  DFF_X1 \f13_reg[14]  ( .D(n1833), .CK(clk), .Q(f13[14]), .QN(n226) );
  DFF_X1 \f13_reg[13]  ( .D(n1832), .CK(clk), .Q(f13[13]), .QN(n227) );
  DFF_X1 \f13_reg[12]  ( .D(n1831), .CK(clk), .Q(f13[12]), .QN(n228) );
  DFF_X1 \f13_reg[11]  ( .D(n1830), .CK(clk), .Q(f13[11]), .QN(n229) );
  DFF_X1 \f13_reg[10]  ( .D(n1829), .CK(clk), .Q(f13[10]), .QN(n230) );
  DFF_X1 \f13_reg[9]  ( .D(n1828), .CK(clk), .Q(f13[9]), .QN(n231) );
  DFF_X1 \f13_reg[8]  ( .D(n1827), .CK(clk), .Q(f13[8]), .QN(n232) );
  DFF_X1 \f13_reg[7]  ( .D(n1826), .CK(clk), .Q(f13[7]), .QN(n233) );
  DFF_X1 \f13_reg[6]  ( .D(n1825), .CK(clk), .Q(f13[6]), .QN(n234) );
  DFF_X1 \f13_reg[5]  ( .D(n1824), .CK(clk), .Q(f13[5]), .QN(n235) );
  DFF_X1 \f13_reg[4]  ( .D(n1823), .CK(clk), .Q(f13[4]), .QN(n236) );
  DFF_X1 \f13_reg[3]  ( .D(n1822), .CK(clk), .Q(f13[3]), .QN(n237) );
  DFF_X1 \f13_reg[2]  ( .D(n1821), .CK(clk), .Q(f13[2]), .QN(n238) );
  DFF_X1 \f13_reg[1]  ( .D(n1820), .CK(clk), .Q(f13[1]), .QN(n239) );
  DFF_X1 \f13_reg[0]  ( .D(n1819), .CK(clk), .Q(f13[0]), .QN(n240) );
  DFF_X1 \f14_reg[14]  ( .D(n1817), .CK(clk), .Q(f14[14]), .QN(n242) );
  DFF_X1 \f14_reg[13]  ( .D(n1816), .CK(clk), .Q(f14[13]), .QN(n243) );
  DFF_X1 \f14_reg[12]  ( .D(n1815), .CK(clk), .Q(f14[12]), .QN(n244) );
  DFF_X1 \f14_reg[11]  ( .D(n1814), .CK(clk), .Q(f14[11]), .QN(n245) );
  DFF_X1 \f14_reg[10]  ( .D(n1813), .CK(clk), .Q(f14[10]), .QN(n246) );
  DFF_X1 \f14_reg[9]  ( .D(n1812), .CK(clk), .Q(f14[9]), .QN(n247) );
  DFF_X1 \f14_reg[8]  ( .D(n1811), .CK(clk), .Q(f14[8]), .QN(n248) );
  DFF_X1 \f14_reg[7]  ( .D(n1810), .CK(clk), .Q(f14[7]), .QN(n249) );
  DFF_X1 \f14_reg[6]  ( .D(n1809), .CK(clk), .Q(f14[6]), .QN(n250) );
  DFF_X1 \f14_reg[5]  ( .D(n1808), .CK(clk), .Q(f14[5]), .QN(n251) );
  DFF_X1 \f14_reg[4]  ( .D(n1807), .CK(clk), .Q(f14[4]), .QN(n252) );
  DFF_X1 \f14_reg[3]  ( .D(n1806), .CK(clk), .Q(f14[3]), .QN(n253) );
  DFF_X1 \f14_reg[2]  ( .D(n1805), .CK(clk), .Q(f14[2]), .QN(n254) );
  DFF_X1 \f14_reg[1]  ( .D(n1804), .CK(clk), .Q(f14[1]), .QN(n255) );
  DFF_X1 \f14_reg[0]  ( .D(n1803), .CK(clk), .Q(f14[0]), .QN(n256) );
  DFF_X1 \f15_reg[14]  ( .D(n1801), .CK(clk), .Q(f15[14]), .QN(n258) );
  DFF_X1 \f15_reg[13]  ( .D(n1800), .CK(clk), .Q(f15[13]), .QN(n259) );
  DFF_X1 \f15_reg[12]  ( .D(n1799), .CK(clk), .Q(f15[12]), .QN(n260) );
  DFF_X1 \f15_reg[11]  ( .D(n1798), .CK(clk), .Q(f15[11]), .QN(n261) );
  DFF_X1 \f15_reg[10]  ( .D(n1797), .CK(clk), .Q(f15[10]), .QN(n262) );
  DFF_X1 \f15_reg[9]  ( .D(n1796), .CK(clk), .Q(f15[9]), .QN(n263) );
  DFF_X1 \f15_reg[8]  ( .D(n1795), .CK(clk), .Q(f15[8]), .QN(n264) );
  DFF_X1 \f15_reg[7]  ( .D(n1794), .CK(clk), .Q(f15[7]), .QN(n265) );
  DFF_X1 \f15_reg[6]  ( .D(n1793), .CK(clk), .Q(f15[6]), .QN(n266) );
  DFF_X1 \f15_reg[5]  ( .D(n1792), .CK(clk), .Q(f15[5]), .QN(n267) );
  DFF_X1 \f15_reg[4]  ( .D(n1791), .CK(clk), .Q(f15[4]), .QN(n268) );
  DFF_X1 \f15_reg[3]  ( .D(n1790), .CK(clk), .Q(f15[3]), .QN(n269) );
  DFF_X1 \f15_reg[2]  ( .D(n1789), .CK(clk), .Q(f15[2]), .QN(n270) );
  DFF_X1 \f15_reg[1]  ( .D(n1788), .CK(clk), .Q(f15[1]), .QN(n271) );
  DFF_X1 \f15_reg[0]  ( .D(n1787), .CK(clk), .Q(f15[0]), .QN(n272) );
  DFF_X1 \f16_reg[15]  ( .D(n1786), .CK(clk), .Q(f16[15]), .QN(n273) );
  DFF_X1 \f16_reg[13]  ( .D(n1784), .CK(clk), .Q(f16[13]), .QN(n275) );
  DFF_X1 \f16_reg[12]  ( .D(n1783), .CK(clk), .Q(f16[12]), .QN(n276) );
  DFF_X1 \f16_reg[11]  ( .D(n1782), .CK(clk), .Q(f16[11]), .QN(n277) );
  DFF_X1 \f16_reg[10]  ( .D(n1781), .CK(clk), .Q(f16[10]), .QN(n278) );
  DFF_X1 \f16_reg[9]  ( .D(n1780), .CK(clk), .Q(f16[9]), .QN(n279) );
  DFF_X1 \f16_reg[8]  ( .D(n1779), .CK(clk), .Q(f16[8]), .QN(n280) );
  DFF_X1 \f16_reg[7]  ( .D(n1778), .CK(clk), .Q(f16[7]), .QN(n281) );
  DFF_X1 \f16_reg[6]  ( .D(n1777), .CK(clk), .Q(f16[6]), .QN(n282) );
  DFF_X1 \f16_reg[5]  ( .D(n1776), .CK(clk), .Q(f16[5]), .QN(n283) );
  DFF_X1 \f16_reg[4]  ( .D(n1775), .CK(clk), .Q(f16[4]), .QN(n284) );
  DFF_X1 \f16_reg[3]  ( .D(n1774), .CK(clk), .Q(f16[3]), .QN(n285) );
  DFF_X1 \f16_reg[2]  ( .D(n1773), .CK(clk), .Q(f16[2]), .QN(n286) );
  DFF_X1 \f16_reg[1]  ( .D(n1772), .CK(clk), .Q(f16[1]), .QN(n287) );
  DFF_X1 \f16_reg[0]  ( .D(n1771), .CK(clk), .Q(f16[0]), .QN(n288) );
  DFF_X1 \f17_reg[14]  ( .D(n1769), .CK(clk), .Q(f17[14]), .QN(n290) );
  DFF_X1 \f17_reg[13]  ( .D(n1768), .CK(clk), .Q(f17[13]), .QN(n291) );
  DFF_X1 \f17_reg[12]  ( .D(n1767), .CK(clk), .Q(f17[12]), .QN(n292) );
  DFF_X1 \f17_reg[11]  ( .D(n1766), .CK(clk), .Q(f17[11]), .QN(n293) );
  DFF_X1 \f17_reg[10]  ( .D(n1765), .CK(clk), .Q(f17[10]), .QN(n294) );
  DFF_X1 \f17_reg[9]  ( .D(n1764), .CK(clk), .Q(f17[9]), .QN(n295) );
  DFF_X1 \f17_reg[8]  ( .D(n1763), .CK(clk), .Q(f17[8]), .QN(n296) );
  DFF_X1 \f17_reg[7]  ( .D(n1762), .CK(clk), .Q(f17[7]), .QN(n297) );
  DFF_X1 \f17_reg[6]  ( .D(n1761), .CK(clk), .Q(f17[6]), .QN(n298) );
  DFF_X1 \f17_reg[5]  ( .D(n1760), .CK(clk), .Q(f17[5]), .QN(n299) );
  DFF_X1 \f17_reg[4]  ( .D(n1759), .CK(clk), .Q(f17[4]), .QN(n300) );
  DFF_X1 \f17_reg[3]  ( .D(n1758), .CK(clk), .Q(f17[3]), .QN(n301) );
  DFF_X1 \f17_reg[2]  ( .D(n1757), .CK(clk), .Q(f17[2]), .QN(n302) );
  DFF_X1 \f17_reg[1]  ( .D(n1756), .CK(clk), .Q(f17[1]), .QN(n303) );
  DFF_X1 \f17_reg[0]  ( .D(n1755), .CK(clk), .Q(f17[0]), .QN(n304) );
  DFF_X1 \f18_reg[14]  ( .D(n1753), .CK(clk), .Q(f18[14]), .QN(n306) );
  DFF_X1 \f18_reg[13]  ( .D(n1752), .CK(clk), .Q(f18[13]), .QN(n307) );
  DFF_X1 \f18_reg[12]  ( .D(n1751), .CK(clk), .Q(f18[12]), .QN(n308) );
  DFF_X1 \f18_reg[11]  ( .D(n1750), .CK(clk), .Q(f18[11]), .QN(n309) );
  DFF_X1 \f18_reg[10]  ( .D(n1749), .CK(clk), .Q(f18[10]), .QN(n310) );
  DFF_X1 \f18_reg[9]  ( .D(n1748), .CK(clk), .Q(f18[9]), .QN(n311) );
  DFF_X1 \f18_reg[8]  ( .D(n1747), .CK(clk), .Q(f18[8]), .QN(n312) );
  DFF_X1 \f18_reg[7]  ( .D(n1746), .CK(clk), .Q(f18[7]), .QN(n313) );
  DFF_X1 \f18_reg[6]  ( .D(n1745), .CK(clk), .Q(f18[6]), .QN(n314) );
  DFF_X1 \f18_reg[5]  ( .D(n1744), .CK(clk), .Q(f18[5]), .QN(n315) );
  DFF_X1 \f18_reg[4]  ( .D(n1743), .CK(clk), .Q(f18[4]), .QN(n316) );
  DFF_X1 \f18_reg[3]  ( .D(n1742), .CK(clk), .Q(f18[3]), .QN(n317) );
  DFF_X1 \f18_reg[2]  ( .D(n1741), .CK(clk), .Q(f18[2]), .QN(n318) );
  DFF_X1 \f18_reg[1]  ( .D(n1740), .CK(clk), .Q(f18[1]), .QN(n319) );
  DFF_X1 \f18_reg[0]  ( .D(n1739), .CK(clk), .Q(f18[0]), .QN(n320) );
  DFF_X1 \f19_reg[14]  ( .D(n1737), .CK(clk), .Q(f19[14]), .QN(n322) );
  DFF_X1 \f19_reg[13]  ( .D(n1736), .CK(clk), .Q(f19[13]), .QN(n323) );
  DFF_X1 \f19_reg[12]  ( .D(n1735), .CK(clk), .Q(f19[12]), .QN(n324) );
  DFF_X1 \f19_reg[11]  ( .D(n1734), .CK(clk), .Q(f19[11]), .QN(n325) );
  DFF_X1 \f19_reg[10]  ( .D(n1733), .CK(clk), .Q(f19[10]), .QN(n326) );
  DFF_X1 \f19_reg[9]  ( .D(n1732), .CK(clk), .Q(f19[9]), .QN(n327) );
  DFF_X1 \f19_reg[8]  ( .D(n1731), .CK(clk), .Q(f19[8]), .QN(n328) );
  DFF_X1 \f19_reg[7]  ( .D(n1730), .CK(clk), .Q(f19[7]), .QN(n329) );
  DFF_X1 \f19_reg[6]  ( .D(n1729), .CK(clk), .Q(f19[6]), .QN(n330) );
  DFF_X1 \f19_reg[5]  ( .D(n1728), .CK(clk), .Q(f19[5]), .QN(n331) );
  DFF_X1 \f19_reg[4]  ( .D(n1727), .CK(clk), .Q(f19[4]), .QN(n332) );
  DFF_X1 \f19_reg[3]  ( .D(n1726), .CK(clk), .Q(f19[3]), .QN(n333) );
  DFF_X1 \f19_reg[2]  ( .D(n1725), .CK(clk), .Q(f19[2]), .QN(n334) );
  DFF_X1 \f19_reg[1]  ( .D(n1724), .CK(clk), .Q(f19[1]), .QN(n335) );
  DFF_X1 \f19_reg[0]  ( .D(n1723), .CK(clk), .Q(f19[0]), .QN(n336) );
  DFF_X1 \f20_reg[14]  ( .D(n1721), .CK(clk), .Q(f20[14]), .QN(n338) );
  DFF_X1 \f20_reg[13]  ( .D(n1720), .CK(clk), .Q(f20[13]), .QN(n339) );
  DFF_X1 \f20_reg[12]  ( .D(n1719), .CK(clk), .Q(f20[12]), .QN(n340) );
  DFF_X1 \f20_reg[11]  ( .D(n1718), .CK(clk), .Q(f20[11]), .QN(n341) );
  DFF_X1 \f20_reg[10]  ( .D(n1717), .CK(clk), .Q(f20[10]), .QN(n342) );
  DFF_X1 \f20_reg[9]  ( .D(n1716), .CK(clk), .Q(f20[9]), .QN(n343) );
  DFF_X1 \f20_reg[8]  ( .D(n1715), .CK(clk), .Q(f20[8]), .QN(n344) );
  DFF_X1 \f20_reg[7]  ( .D(n1714), .CK(clk), .Q(f20[7]), .QN(n345) );
  DFF_X1 \f20_reg[6]  ( .D(n1713), .CK(clk), .Q(f20[6]), .QN(n346) );
  DFF_X1 \f20_reg[5]  ( .D(n1712), .CK(clk), .Q(f20[5]), .QN(n347) );
  DFF_X1 \f20_reg[4]  ( .D(n1711), .CK(clk), .Q(f20[4]), .QN(n348) );
  DFF_X1 \f20_reg[3]  ( .D(n1710), .CK(clk), .Q(f20[3]), .QN(n349) );
  DFF_X1 \f20_reg[2]  ( .D(n1709), .CK(clk), .Q(f20[2]), .QN(n350) );
  DFF_X1 \f20_reg[1]  ( .D(n1708), .CK(clk), .Q(f20[1]), .QN(n351) );
  DFF_X1 \f20_reg[0]  ( .D(n1707), .CK(clk), .Q(f20[0]), .QN(n352) );
  DFF_X1 \f21_reg[14]  ( .D(n1705), .CK(clk), .Q(f21[14]), .QN(n354) );
  DFF_X1 \f21_reg[13]  ( .D(n1704), .CK(clk), .Q(f21[13]), .QN(n355) );
  DFF_X1 \f21_reg[12]  ( .D(n1703), .CK(clk), .Q(f21[12]), .QN(n356) );
  DFF_X1 \f21_reg[11]  ( .D(n1702), .CK(clk), .Q(f21[11]), .QN(n357) );
  DFF_X1 \f21_reg[10]  ( .D(n1701), .CK(clk), .Q(f21[10]), .QN(n358) );
  DFF_X1 \f21_reg[9]  ( .D(n1700), .CK(clk), .Q(f21[9]), .QN(n359) );
  DFF_X1 \f21_reg[8]  ( .D(n1699), .CK(clk), .Q(f21[8]), .QN(n360) );
  DFF_X1 \f21_reg[7]  ( .D(n1698), .CK(clk), .Q(f21[7]), .QN(n361) );
  DFF_X1 \f21_reg[6]  ( .D(n1697), .CK(clk), .Q(f21[6]), .QN(n362) );
  DFF_X1 \f21_reg[5]  ( .D(n1696), .CK(clk), .Q(f21[5]), .QN(n363) );
  DFF_X1 \f21_reg[4]  ( .D(n1695), .CK(clk), .Q(f21[4]), .QN(n364) );
  DFF_X1 \f21_reg[3]  ( .D(n1694), .CK(clk), .Q(f21[3]), .QN(n365) );
  DFF_X1 \f21_reg[2]  ( .D(n1693), .CK(clk), .Q(f21[2]), .QN(n366) );
  DFF_X1 \f21_reg[1]  ( .D(n1692), .CK(clk), .Q(f21[1]), .QN(n367) );
  DFF_X1 \f21_reg[0]  ( .D(n1691), .CK(clk), .Q(f21[0]), .QN(n368) );
  DFF_X1 \f22_reg[14]  ( .D(n1689), .CK(clk), .Q(f22[14]), .QN(n370) );
  DFF_X1 \f22_reg[13]  ( .D(n1688), .CK(clk), .Q(f22[13]), .QN(n371) );
  DFF_X1 \f22_reg[12]  ( .D(n1687), .CK(clk), .Q(f22[12]), .QN(n372) );
  DFF_X1 \f22_reg[11]  ( .D(n1686), .CK(clk), .Q(f22[11]), .QN(n373) );
  DFF_X1 \f22_reg[10]  ( .D(n1685), .CK(clk), .Q(f22[10]), .QN(n374) );
  DFF_X1 \f22_reg[9]  ( .D(n1684), .CK(clk), .Q(f22[9]), .QN(n375) );
  DFF_X1 \f22_reg[8]  ( .D(n1683), .CK(clk), .Q(f22[8]), .QN(n376) );
  DFF_X1 \f22_reg[7]  ( .D(n1682), .CK(clk), .Q(f22[7]), .QN(n377) );
  DFF_X1 \f22_reg[6]  ( .D(n1681), .CK(clk), .Q(f22[6]), .QN(n378) );
  DFF_X1 \f22_reg[5]  ( .D(n1680), .CK(clk), .Q(f22[5]), .QN(n379) );
  DFF_X1 \f22_reg[4]  ( .D(n1679), .CK(clk), .Q(f22[4]), .QN(n380) );
  DFF_X1 \f22_reg[3]  ( .D(n1678), .CK(clk), .Q(f22[3]), .QN(n381) );
  DFF_X1 \f22_reg[2]  ( .D(n1677), .CK(clk), .Q(f22[2]), .QN(n382) );
  DFF_X1 \f22_reg[1]  ( .D(n1676), .CK(clk), .Q(f22[1]), .QN(n383) );
  DFF_X1 \f22_reg[0]  ( .D(n1675), .CK(clk), .Q(f22[0]), .QN(n384) );
  DFF_X1 \f23_reg[15]  ( .D(n1674), .CK(clk), .Q(f23[15]), .QN(n385) );
  DFF_X1 \f23_reg[14]  ( .D(n1673), .CK(clk), .Q(f23[14]), .QN(n386) );
  DFF_X1 \f23_reg[13]  ( .D(n1672), .CK(clk), .Q(f23[13]), .QN(n387) );
  DFF_X1 \f23_reg[12]  ( .D(n1671), .CK(clk), .Q(f23[12]), .QN(n388) );
  DFF_X1 \f23_reg[11]  ( .D(n1670), .CK(clk), .Q(f23[11]), .QN(n389) );
  DFF_X1 \f23_reg[10]  ( .D(n1669), .CK(clk), .Q(f23[10]), .QN(n390) );
  DFF_X1 \f23_reg[9]  ( .D(n1668), .CK(clk), .Q(f23[9]), .QN(n391) );
  DFF_X1 \f23_reg[8]  ( .D(n1667), .CK(clk), .Q(f23[8]), .QN(n392) );
  DFF_X1 \f23_reg[7]  ( .D(n1666), .CK(clk), .Q(f23[7]), .QN(n393) );
  DFF_X1 \f23_reg[6]  ( .D(n1665), .CK(clk), .Q(f23[6]), .QN(n394) );
  DFF_X1 \f23_reg[5]  ( .D(n1664), .CK(clk), .Q(f23[5]), .QN(n395) );
  DFF_X1 \f23_reg[4]  ( .D(n1663), .CK(clk), .Q(f23[4]), .QN(n396) );
  DFF_X1 \f23_reg[3]  ( .D(n1662), .CK(clk), .Q(f23[3]), .QN(n397) );
  DFF_X1 \f23_reg[2]  ( .D(n1661), .CK(clk), .Q(f23[2]), .QN(n398) );
  DFF_X1 \f23_reg[1]  ( .D(n1660), .CK(clk), .Q(f23[1]), .QN(n399) );
  DFF_X1 \f23_reg[0]  ( .D(n1659), .CK(clk), .Q(f23[0]), .QN(n400) );
  DFF_X1 \f24_reg[15]  ( .D(n1658), .CK(clk), .Q(f24[15]), .QN(n401) );
  DFF_X1 \f24_reg[14]  ( .D(n1657), .CK(clk), .Q(f24[14]), .QN(n402) );
  DFF_X1 \f24_reg[13]  ( .D(n1656), .CK(clk), .Q(f24[13]), .QN(n403) );
  DFF_X1 \f24_reg[12]  ( .D(n1655), .CK(clk), .Q(f24[12]), .QN(n404) );
  DFF_X1 \f24_reg[11]  ( .D(n1654), .CK(clk), .Q(f24[11]), .QN(n405) );
  DFF_X1 \f24_reg[10]  ( .D(n1653), .CK(clk), .Q(f24[10]), .QN(n406) );
  DFF_X1 \f24_reg[9]  ( .D(n1652), .CK(clk), .Q(f24[9]), .QN(n407) );
  DFF_X1 \f24_reg[8]  ( .D(n1651), .CK(clk), .Q(f24[8]), .QN(n408) );
  DFF_X1 \f24_reg[7]  ( .D(n1650), .CK(clk), .Q(f24[7]), .QN(n409) );
  DFF_X1 \f24_reg[6]  ( .D(n1649), .CK(clk), .Q(f24[6]), .QN(n410) );
  DFF_X1 \f24_reg[5]  ( .D(n1648), .CK(clk), .Q(f24[5]), .QN(n411) );
  DFF_X1 \f24_reg[4]  ( .D(n1647), .CK(clk), .Q(f24[4]), .QN(n412) );
  DFF_X1 \f24_reg[3]  ( .D(n1646), .CK(clk), .Q(f24[3]), .QN(n413) );
  DFF_X1 \f24_reg[2]  ( .D(n1645), .CK(clk), .Q(f24[2]), .QN(n414) );
  DFF_X1 \f24_reg[1]  ( .D(n1644), .CK(clk), .Q(f24[1]), .QN(n415) );
  DFF_X1 \f24_reg[0]  ( .D(n1643), .CK(clk), .Q(f24[0]), .QN(n416) );
  DFF_X1 \f25_reg[14]  ( .D(n1641), .CK(clk), .Q(f25[14]), .QN(n418) );
  DFF_X1 \f25_reg[13]  ( .D(n1640), .CK(clk), .Q(f25[13]), .QN(n419) );
  DFF_X1 \f25_reg[12]  ( .D(n1639), .CK(clk), .Q(f25[12]), .QN(n420) );
  DFF_X1 \f25_reg[11]  ( .D(n1638), .CK(clk), .Q(f25[11]), .QN(n421) );
  DFF_X1 \f25_reg[10]  ( .D(n1637), .CK(clk), .Q(f25[10]), .QN(n422) );
  DFF_X1 \f25_reg[9]  ( .D(n1636), .CK(clk), .Q(f25[9]), .QN(n423) );
  DFF_X1 \f25_reg[8]  ( .D(n1635), .CK(clk), .Q(f25[8]), .QN(n424) );
  DFF_X1 \f25_reg[7]  ( .D(n1634), .CK(clk), .Q(f25[7]), .QN(n425) );
  DFF_X1 \f25_reg[6]  ( .D(n1633), .CK(clk), .Q(f25[6]), .QN(n426) );
  DFF_X1 \f25_reg[5]  ( .D(n1632), .CK(clk), .Q(f25[5]), .QN(n427) );
  DFF_X1 \f25_reg[4]  ( .D(n1631), .CK(clk), .Q(f25[4]), .QN(n428) );
  DFF_X1 \f25_reg[3]  ( .D(n1630), .CK(clk), .Q(f25[3]), .QN(n429) );
  DFF_X1 \f25_reg[2]  ( .D(n1629), .CK(clk), .Q(f25[2]), .QN(n430) );
  DFF_X1 \f25_reg[1]  ( .D(n1628), .CK(clk), .Q(f25[1]), .QN(n431) );
  DFF_X1 \f25_reg[0]  ( .D(n1627), .CK(clk), .Q(f25[0]), .QN(n432) );
  DFF_X1 \f26_reg[14]  ( .D(n1625), .CK(clk), .Q(f26[14]), .QN(n434) );
  DFF_X1 \f26_reg[13]  ( .D(n1624), .CK(clk), .Q(f26[13]), .QN(n435) );
  DFF_X1 \f26_reg[12]  ( .D(n1623), .CK(clk), .Q(f26[12]), .QN(n436) );
  DFF_X1 \f26_reg[11]  ( .D(n1622), .CK(clk), .Q(f26[11]), .QN(n437) );
  DFF_X1 \f26_reg[10]  ( .D(n1621), .CK(clk), .Q(f26[10]), .QN(n438) );
  DFF_X1 \f26_reg[9]  ( .D(n1620), .CK(clk), .Q(f26[9]), .QN(n439) );
  DFF_X1 \f26_reg[8]  ( .D(n1619), .CK(clk), .Q(f26[8]), .QN(n440) );
  DFF_X1 \f26_reg[7]  ( .D(n1618), .CK(clk), .Q(f26[7]), .QN(n441) );
  DFF_X1 \f26_reg[6]  ( .D(n1617), .CK(clk), .Q(f26[6]), .QN(n442) );
  DFF_X1 \f26_reg[5]  ( .D(n1616), .CK(clk), .Q(f26[5]), .QN(n443) );
  DFF_X1 \f26_reg[4]  ( .D(n1615), .CK(clk), .Q(f26[4]), .QN(n444) );
  DFF_X1 \f26_reg[3]  ( .D(n1614), .CK(clk), .Q(f26[3]), .QN(n445) );
  DFF_X1 \f26_reg[2]  ( .D(n1613), .CK(clk), .Q(f26[2]), .QN(n446) );
  DFF_X1 \f26_reg[1]  ( .D(n1612), .CK(clk), .Q(f26[1]), .QN(n447) );
  DFF_X1 \f26_reg[0]  ( .D(n1611), .CK(clk), .Q(f26[0]), .QN(n448) );
  DFF_X1 \f27_reg[15]  ( .D(n1610), .CK(clk), .Q(f27[15]), .QN(n449) );
  DFF_X1 \f27_reg[14]  ( .D(n1609), .CK(clk), .Q(f27[14]), .QN(n450) );
  DFF_X1 \f27_reg[13]  ( .D(n1608), .CK(clk), .Q(f27[13]), .QN(n451) );
  DFF_X1 \f27_reg[12]  ( .D(n1607), .CK(clk), .Q(f27[12]), .QN(n452) );
  DFF_X1 \f27_reg[11]  ( .D(n1606), .CK(clk), .Q(f27[11]), .QN(n453) );
  DFF_X1 \f27_reg[10]  ( .D(n1605), .CK(clk), .Q(f27[10]), .QN(n454) );
  DFF_X1 \f27_reg[9]  ( .D(n1604), .CK(clk), .Q(f27[9]), .QN(n455) );
  DFF_X1 \f27_reg[8]  ( .D(n1603), .CK(clk), .Q(f27[8]), .QN(n456) );
  DFF_X1 \f27_reg[7]  ( .D(n1602), .CK(clk), .Q(f27[7]), .QN(n457) );
  DFF_X1 \f27_reg[6]  ( .D(n1601), .CK(clk), .Q(f27[6]), .QN(n458) );
  DFF_X1 \f27_reg[5]  ( .D(n1600), .CK(clk), .Q(f27[5]), .QN(n459) );
  DFF_X1 \f27_reg[4]  ( .D(n1599), .CK(clk), .Q(f27[4]), .QN(n460) );
  DFF_X1 \f27_reg[3]  ( .D(n1598), .CK(clk), .Q(f27[3]), .QN(n461) );
  DFF_X1 \f27_reg[2]  ( .D(n1597), .CK(clk), .Q(f27[2]), .QN(n462) );
  DFF_X1 \f27_reg[1]  ( .D(n1596), .CK(clk), .Q(f27[1]), .QN(n463) );
  DFF_X1 \f27_reg[0]  ( .D(n1595), .CK(clk), .Q(f27[0]), .QN(n464) );
  DFF_X1 \f28_reg[15]  ( .D(n1594), .CK(clk), .Q(f28[15]), .QN(n465) );
  DFF_X1 \f28_reg[14]  ( .D(n1593), .CK(clk), .Q(f28[14]), .QN(n466) );
  DFF_X1 \f28_reg[13]  ( .D(n1592), .CK(clk), .Q(f28[13]), .QN(n467) );
  DFF_X1 \f28_reg[12]  ( .D(n1591), .CK(clk), .Q(f28[12]), .QN(n468) );
  DFF_X1 \f28_reg[11]  ( .D(n1590), .CK(clk), .Q(f28[11]), .QN(n469) );
  DFF_X1 \f28_reg[10]  ( .D(n1589), .CK(clk), .Q(f28[10]), .QN(n470) );
  DFF_X1 \f28_reg[9]  ( .D(n1588), .CK(clk), .Q(f28[9]), .QN(n471) );
  DFF_X1 \f28_reg[8]  ( .D(n1587), .CK(clk), .Q(f28[8]), .QN(n472) );
  DFF_X1 \f28_reg[7]  ( .D(n1586), .CK(clk), .Q(f28[7]), .QN(n473) );
  DFF_X1 \f28_reg[6]  ( .D(n1585), .CK(clk), .Q(f28[6]), .QN(n474) );
  DFF_X1 \f28_reg[5]  ( .D(n1584), .CK(clk), .Q(f28[5]), .QN(n475) );
  DFF_X1 \f28_reg[4]  ( .D(n1583), .CK(clk), .Q(f28[4]), .QN(n476) );
  DFF_X1 \f28_reg[3]  ( .D(n1582), .CK(clk), .Q(f28[3]), .QN(n477) );
  DFF_X1 \f28_reg[2]  ( .D(n1581), .CK(clk), .Q(f28[2]), .QN(n478) );
  DFF_X1 \f28_reg[1]  ( .D(n1580), .CK(clk), .Q(f28[1]), .QN(n479) );
  DFF_X1 \f28_reg[0]  ( .D(n1579), .CK(clk), .Q(f28[0]), .QN(n480) );
  DFF_X1 \f29_reg[14]  ( .D(n1577), .CK(clk), .Q(f29[14]), .QN(n482) );
  DFF_X1 \f29_reg[13]  ( .D(n1576), .CK(clk), .Q(f29[13]), .QN(n483) );
  DFF_X1 \f29_reg[12]  ( .D(n1575), .CK(clk), .Q(f29[12]), .QN(n484) );
  DFF_X1 \f29_reg[11]  ( .D(n1574), .CK(clk), .Q(f29[11]), .QN(n485) );
  DFF_X1 \f29_reg[10]  ( .D(n1573), .CK(clk), .Q(f29[10]), .QN(n486) );
  DFF_X1 \f29_reg[9]  ( .D(n1572), .CK(clk), .Q(f29[9]), .QN(n487) );
  DFF_X1 \f29_reg[8]  ( .D(n1571), .CK(clk), .Q(f29[8]), .QN(n488) );
  DFF_X1 \f29_reg[7]  ( .D(n1570), .CK(clk), .Q(f29[7]), .QN(n489) );
  DFF_X1 \f29_reg[6]  ( .D(n1569), .CK(clk), .Q(f29[6]), .QN(n490) );
  DFF_X1 \f29_reg[5]  ( .D(n1568), .CK(clk), .Q(f29[5]), .QN(n491) );
  DFF_X1 \f29_reg[4]  ( .D(n1567), .CK(clk), .Q(f29[4]), .QN(n492) );
  DFF_X1 \f29_reg[3]  ( .D(n1566), .CK(clk), .Q(f29[3]), .QN(n493) );
  DFF_X1 \f29_reg[2]  ( .D(n1565), .CK(clk), .Q(f29[2]), .QN(n494) );
  DFF_X1 \f29_reg[1]  ( .D(n1564), .CK(clk), .Q(f29[1]), .QN(n495) );
  DFF_X1 \f29_reg[0]  ( .D(n1563), .CK(clk), .Q(f29[0]), .QN(n496) );
  DFF_X1 \f30_reg[14]  ( .D(n1561), .CK(clk), .Q(f30[14]), .QN(n498) );
  DFF_X1 \f30_reg[13]  ( .D(n1560), .CK(clk), .Q(f30[13]), .QN(n499) );
  DFF_X1 \f30_reg[12]  ( .D(n1559), .CK(clk), .Q(f30[12]), .QN(n500) );
  DFF_X1 \f30_reg[11]  ( .D(n1558), .CK(clk), .Q(f30[11]), .QN(n501) );
  DFF_X1 \f30_reg[10]  ( .D(n1557), .CK(clk), .Q(f30[10]), .QN(n502) );
  DFF_X1 \f30_reg[9]  ( .D(n1556), .CK(clk), .Q(f30[9]), .QN(n503) );
  DFF_X1 \f30_reg[8]  ( .D(n1555), .CK(clk), .Q(f30[8]), .QN(n504) );
  DFF_X1 \f30_reg[7]  ( .D(n1554), .CK(clk), .Q(f30[7]), .QN(n505) );
  DFF_X1 \f30_reg[6]  ( .D(n1553), .CK(clk), .Q(f30[6]), .QN(n506) );
  DFF_X1 \f30_reg[5]  ( .D(n1552), .CK(clk), .Q(f30[5]), .QN(n507) );
  DFF_X1 \f30_reg[4]  ( .D(n1551), .CK(clk), .Q(f30[4]), .QN(n508) );
  DFF_X1 \f30_reg[3]  ( .D(n1550), .CK(clk), .Q(f30[3]), .QN(n509) );
  DFF_X1 \f30_reg[2]  ( .D(n1549), .CK(clk), .Q(f30[2]), .QN(n510) );
  DFF_X1 \f30_reg[1]  ( .D(n1548), .CK(clk), .Q(f30[1]), .QN(n511) );
  DFF_X1 \f30_reg[0]  ( .D(n1547), .CK(clk), .Q(f30[0]), .QN(n512) );
  DFF_X1 \f31_reg[14]  ( .D(n1545), .CK(clk), .Q(f31[14]), .QN(n514) );
  DFF_X1 \f31_reg[13]  ( .D(n1544), .CK(clk), .Q(f31[13]), .QN(n515) );
  DFF_X1 \f31_reg[12]  ( .D(n1543), .CK(clk), .Q(f31[12]), .QN(n516) );
  DFF_X1 \f31_reg[11]  ( .D(n1542), .CK(clk), .Q(f31[11]), .QN(n517) );
  DFF_X1 \f31_reg[10]  ( .D(n1541), .CK(clk), .Q(f31[10]), .QN(n518) );
  DFF_X1 \f31_reg[9]  ( .D(n1540), .CK(clk), .Q(f31[9]), .QN(n519) );
  DFF_X1 \f31_reg[8]  ( .D(n1539), .CK(clk), .Q(f31[8]), .QN(n520) );
  DFF_X1 \f31_reg[7]  ( .D(n1538), .CK(clk), .Q(f31[7]), .QN(n521) );
  DFF_X1 \f31_reg[6]  ( .D(n1537), .CK(clk), .Q(f31[6]), .QN(n522) );
  DFF_X1 \f31_reg[5]  ( .D(n1536), .CK(clk), .Q(f31[5]), .QN(n523) );
  DFF_X1 \f31_reg[4]  ( .D(n1535), .CK(clk), .Q(f31[4]), .QN(n524) );
  DFF_X1 \f31_reg[3]  ( .D(n1534), .CK(clk), .Q(f31[3]), .QN(n525) );
  DFF_X1 \f31_reg[2]  ( .D(n1533), .CK(clk), .Q(f31[2]), .QN(n526) );
  DFF_X1 \f31_reg[1]  ( .D(n1532), .CK(clk), .Q(f31[1]), .QN(n527) );
  DFF_X1 \f31_reg[0]  ( .D(n1531), .CK(clk), .Q(f31[0]), .QN(n528) );
  DFF_X1 \f32_reg[15]  ( .D(n1530), .CK(clk), .Q(f32[15]), .QN(n529) );
  DFF_X1 \f_reg[15]  ( .D(n1499), .CK(clk), .Q(f[15]) );
  DFF_X1 \f32_reg[14]  ( .D(n1529), .CK(clk), .Q(f32[14]), .QN(n530) );
  DFF_X1 \f_reg[14]  ( .D(n1500), .CK(clk), .Q(f[14]) );
  DFF_X1 \f32_reg[13]  ( .D(n1528), .CK(clk), .Q(f32[13]), .QN(n531) );
  DFF_X1 \f_reg[13]  ( .D(n1501), .CK(clk), .Q(f[13]) );
  DFF_X1 \f32_reg[12]  ( .D(n1527), .CK(clk), .Q(f32[12]), .QN(n532) );
  DFF_X1 \f_reg[12]  ( .D(n1502), .CK(clk), .Q(f[12]) );
  DFF_X1 \f32_reg[11]  ( .D(n1526), .CK(clk), .Q(f32[11]), .QN(n533) );
  DFF_X1 \f_reg[11]  ( .D(n1503), .CK(clk), .Q(f[11]) );
  DFF_X1 \f32_reg[10]  ( .D(n1525), .CK(clk), .Q(f32[10]), .QN(n534) );
  DFF_X1 \f_reg[10]  ( .D(n1504), .CK(clk), .Q(f[10]) );
  DFF_X1 \f32_reg[9]  ( .D(n1524), .CK(clk), .Q(f32[9]), .QN(n535) );
  DFF_X1 \f_reg[9]  ( .D(n1505), .CK(clk), .Q(f[9]) );
  DFF_X1 \f32_reg[8]  ( .D(n1523), .CK(clk), .Q(f32[8]), .QN(n536) );
  DFF_X1 \f_reg[8]  ( .D(n1506), .CK(clk), .Q(f[8]) );
  DFF_X1 \f32_reg[7]  ( .D(n1522), .CK(clk), .Q(f32[7]), .QN(n537) );
  DFF_X1 \f_reg[7]  ( .D(n1507), .CK(clk), .Q(f[7]) );
  DFF_X1 \f32_reg[6]  ( .D(n1521), .CK(clk), .Q(f32[6]), .QN(n538) );
  DFF_X1 \f_reg[6]  ( .D(n1508), .CK(clk), .Q(f[6]) );
  DFF_X1 \f32_reg[5]  ( .D(n1520), .CK(clk), .Q(f32[5]), .QN(n539) );
  DFF_X1 \f_reg[5]  ( .D(n1509), .CK(clk), .Q(f[5]) );
  DFF_X1 \f32_reg[4]  ( .D(n1519), .CK(clk), .Q(f32[4]), .QN(n540) );
  DFF_X1 \f_reg[4]  ( .D(n1510), .CK(clk), .Q(f[4]) );
  DFF_X1 \f32_reg[3]  ( .D(n1518), .CK(clk), .Q(f32[3]), .QN(n541) );
  DFF_X1 \f_reg[3]  ( .D(n1511), .CK(clk), .Q(f[3]) );
  DFF_X1 \f32_reg[2]  ( .D(n1517), .CK(clk), .Q(f32[2]), .QN(n542) );
  DFF_X1 \f_reg[2]  ( .D(n1512), .CK(clk), .Q(f[2]) );
  DFF_X1 \f32_reg[1]  ( .D(n1516), .CK(clk), .Q(f32[1]), .QN(n543) );
  DFF_X1 \f_reg[1]  ( .D(n1513), .CK(clk), .Q(f[1]) );
  DFF_X1 \f32_reg[0]  ( .D(n1515), .CK(clk), .Q(f32[0]), .QN(n544) );
  DFF_X1 \f_reg[0]  ( .D(n1514), .CK(clk), .Q(f[0]) );
  NAND3_X1 U1483 ( .A1(n982), .A2(n1002), .A3(add_r31[0]), .ZN(n1001) );
  memory_WIDTH8_SIZE32_LOGSIZE5_0 mem_x ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_x), .addr(addr_x), .wr_en(wr_en_x) );
  memory_WIDTH8_SIZE32_LOGSIZE5_32 mem_a1 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a1), .addr(addr_a1), .wr_en(wr_en_a1) );
  memory_WIDTH8_SIZE32_LOGSIZE5_31 mem_a2 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a2), .addr(addr_a2), .wr_en(wr_en_a2) );
  memory_WIDTH8_SIZE32_LOGSIZE5_30 mem_a3 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a3), .addr(addr_a3), .wr_en(wr_en_a3) );
  memory_WIDTH8_SIZE32_LOGSIZE5_29 mem_a4 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a4), .addr(addr_a4), .wr_en(wr_en_a4) );
  memory_WIDTH8_SIZE32_LOGSIZE5_28 mem_a5 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a5), .addr(addr_a5), .wr_en(wr_en_a5) );
  memory_WIDTH8_SIZE32_LOGSIZE5_27 mem_a6 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a6), .addr(addr_a6), .wr_en(wr_en_a6) );
  memory_WIDTH8_SIZE32_LOGSIZE5_26 mem_a7 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a7), .addr(addr_a7), .wr_en(wr_en_a7) );
  memory_WIDTH8_SIZE32_LOGSIZE5_25 mem_a8 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a8), .addr(addr_a8), .wr_en(wr_en_a8) );
  memory_WIDTH8_SIZE32_LOGSIZE5_24 mem_a9 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a9), .addr(addr_a9), .wr_en(wr_en_a9) );
  memory_WIDTH8_SIZE32_LOGSIZE5_23 mem_a10 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a10), .addr(addr_a10), .wr_en(wr_en_a10) );
  memory_WIDTH8_SIZE32_LOGSIZE5_22 mem_a11 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a11), .addr(addr_a11), .wr_en(wr_en_a11) );
  memory_WIDTH8_SIZE32_LOGSIZE5_21 mem_a12 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a12), .addr(addr_a12), .wr_en(wr_en_a12) );
  memory_WIDTH8_SIZE32_LOGSIZE5_20 mem_a13 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a13), .addr(addr_a13), .wr_en(wr_en_a13) );
  memory_WIDTH8_SIZE32_LOGSIZE5_19 mem_a14 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a14), .addr(addr_a14), .wr_en(wr_en_a14) );
  memory_WIDTH8_SIZE32_LOGSIZE5_18 mem_a15 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a15), .addr(addr_a15), .wr_en(wr_en_a15) );
  memory_WIDTH8_SIZE32_LOGSIZE5_17 mem_a16 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a16), .addr(addr_a16), .wr_en(wr_en_a16) );
  memory_WIDTH8_SIZE32_LOGSIZE5_16 mem_a17 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a17), .addr(addr_a17), .wr_en(wr_en_a17) );
  memory_WIDTH8_SIZE32_LOGSIZE5_15 mem_a18 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a18), .addr(addr_a18), .wr_en(wr_en_a18) );
  memory_WIDTH8_SIZE32_LOGSIZE5_14 mem_a19 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a19), .addr(addr_a19), .wr_en(wr_en_a19) );
  memory_WIDTH8_SIZE32_LOGSIZE5_13 mem_a20 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a20), .addr(addr_a20), .wr_en(wr_en_a20) );
  memory_WIDTH8_SIZE32_LOGSIZE5_12 mem_a21 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a21), .addr(addr_a21), .wr_en(wr_en_a21) );
  memory_WIDTH8_SIZE32_LOGSIZE5_11 mem_a22 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a22), .addr(addr_a22), .wr_en(wr_en_a22) );
  memory_WIDTH8_SIZE32_LOGSIZE5_10 mem_a23 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a23), .addr(addr_a23), .wr_en(wr_en_a23) );
  memory_WIDTH8_SIZE32_LOGSIZE5_9 mem_a24 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a24), .addr(addr_a24), .wr_en(wr_en_a24) );
  memory_WIDTH8_SIZE32_LOGSIZE5_8 mem_a25 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a25), .addr(addr_a25), .wr_en(wr_en_a25) );
  memory_WIDTH8_SIZE32_LOGSIZE5_7 mem_a26 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a26), .addr(addr_a26), .wr_en(wr_en_a26) );
  memory_WIDTH8_SIZE32_LOGSIZE5_6 mem_a27 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a27), .addr(addr_a27), .wr_en(wr_en_a27) );
  memory_WIDTH8_SIZE32_LOGSIZE5_5 mem_a28 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a28), .addr(addr_a28), .wr_en(wr_en_a28) );
  memory_WIDTH8_SIZE32_LOGSIZE5_4 mem_a29 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a29), .addr(addr_a29), .wr_en(wr_en_a29) );
  memory_WIDTH8_SIZE32_LOGSIZE5_3 mem_a30 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a30), .addr(addr_a30), .wr_en(wr_en_a30) );
  memory_WIDTH8_SIZE32_LOGSIZE5_2 mem_a31 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a31), .addr(addr_a31), .wr_en(wr_en_a31) );
  memory_WIDTH8_SIZE32_LOGSIZE5_1 mem_a32 ( .clk(clk), .data_in(data_in), 
        .data_out(data_out_a32), .addr(addr_a32), .wr_en(wr_en_a32) );
  memory_WIDTH16_SIZE32_LOGSIZE5 mem_y ( .clk(clk), .data_in(f), .data_out(
        data_out), .addr(addr_y), .wr_en(wr_en_y) );
  datapath_DW_mult_tc_31 mult_108 ( .a(data_out_a1), .b({n2144, n2141, n2138, 
        n2135, n558, n571, n2124, n2121}), .product({\mul_out1[15] , 
        \mul_out1[14] , \mul_out1[13] , \mul_out1[12] , \mul_out1[11] , 
        \mul_out1[10] , \mul_out1[9] , \mul_out1[8] , \mul_out1[7] , 
        \mul_out1[6] , \mul_out1[5] , \mul_out1[4] , \mul_out1[3] , 
        \mul_out1[2] , \mul_out1[1] , \mul_out1[0] }) );
  datapath_DW01_add_31 add_109 ( .A(f1), .B({\mul_out1[15] , \mul_out1[14] , 
        \mul_out1[13] , \mul_out1[12] , \mul_out1[11] , \mul_out1[10] , 
        \mul_out1[9] , \mul_out1[8] , \mul_out1[7] , \mul_out1[6] , 
        \mul_out1[5] , \mul_out1[4] , \mul_out1[3] , \mul_out1[2] , 
        \mul_out1[1] , \mul_out1[0] }), .CI(1'b0), .SUM(add_r1) );
  datapath_DW_mult_tc_30 mult_110 ( .a(data_out_a2), .b({n2144, n2141, n2138, 
        n2133, n557, n570, n2124, n2123}), .product({\mul_out2[15] , 
        \mul_out2[14] , \mul_out2[13] , \mul_out2[12] , \mul_out2[11] , 
        \mul_out2[10] , \mul_out2[9] , \mul_out2[8] , \mul_out2[7] , 
        \mul_out2[6] , \mul_out2[5] , \mul_out2[4] , \mul_out2[3] , 
        \mul_out2[2] , \mul_out2[1] , \mul_out2[0] }) );
  datapath_DW01_add_30 add_111 ( .A(f2), .B({\mul_out2[15] , \mul_out2[14] , 
        \mul_out2[13] , \mul_out2[12] , \mul_out2[11] , \mul_out2[10] , 
        \mul_out2[9] , \mul_out2[8] , \mul_out2[7] , \mul_out2[6] , 
        \mul_out2[5] , \mul_out2[4] , \mul_out2[3] , \mul_out2[2] , 
        \mul_out2[1] , \mul_out2[0] }), .CI(1'b0), .SUM(add_r2) );
  datapath_DW_mult_tc_29 mult_112 ( .a(data_out_a3), .b({n2144, n2141, n2138, 
        n2135, n2132, n570, n2029, n2121}), .product({\mul_out3[15] , 
        \mul_out3[14] , \mul_out3[13] , \mul_out3[12] , \mul_out3[11] , 
        \mul_out3[10] , \mul_out3[9] , \mul_out3[8] , \mul_out3[7] , 
        \mul_out3[6] , \mul_out3[5] , \mul_out3[4] , \mul_out3[3] , 
        \mul_out3[2] , \mul_out3[1] , \mul_out3[0] }) );
  datapath_DW01_add_29 add_113 ( .A(f3), .B({\mul_out3[15] , \mul_out3[14] , 
        \mul_out3[13] , \mul_out3[12] , \mul_out3[11] , \mul_out3[10] , 
        \mul_out3[9] , \mul_out3[8] , \mul_out3[7] , \mul_out3[6] , 
        \mul_out3[5] , \mul_out3[4] , \mul_out3[3] , \mul_out3[2] , 
        \mul_out3[1] , \mul_out3[0] }), .CI(1'b0), .SUM(add_r3) );
  datapath_DW_mult_tc_28 mult_114 ( .a(data_out_a4), .b({n2144, n2141, n2138, 
        n2, n557, n570, n27, n2123}), .product({\mul_out4[15] , \mul_out4[14] , 
        \mul_out4[13] , \mul_out4[12] , \mul_out4[11] , \mul_out4[10] , 
        \mul_out4[9] , \mul_out4[8] , \mul_out4[7] , \mul_out4[6] , 
        \mul_out4[5] , \mul_out4[4] , \mul_out4[3] , \mul_out4[2] , 
        \mul_out4[1] , \mul_out4[0] }) );
  datapath_DW01_add_28 add_115 ( .A(f4), .B({\mul_out4[15] , \mul_out4[14] , 
        \mul_out4[13] , \mul_out4[12] , \mul_out4[11] , \mul_out4[10] , 
        \mul_out4[9] , \mul_out4[8] , \mul_out4[7] , \mul_out4[6] , 
        \mul_out4[5] , \mul_out4[4] , \mul_out4[3] , \mul_out4[2] , 
        \mul_out4[1] , \mul_out4[0] }), .CI(1'b0), .SUM(add_r4) );
  datapath_DW_mult_tc_27 mult_116 ( .a(data_out_a5), .b({n2144, n2141, n2138, 
        n2, n2132, n9, n2028, n2122}), .product({\mul_out5[15] , 
        \mul_out5[14] , \mul_out5[13] , \mul_out5[12] , \mul_out5[11] , 
        \mul_out5[10] , \mul_out5[9] , \mul_out5[8] , \mul_out5[7] , 
        \mul_out5[6] , \mul_out5[5] , \mul_out5[4] , \mul_out5[3] , 
        \mul_out5[2] , \mul_out5[1] , \mul_out5[0] }) );
  datapath_DW01_add_27 add_117 ( .A(f5), .B({\mul_out5[15] , \mul_out5[14] , 
        \mul_out5[13] , \mul_out5[12] , \mul_out5[11] , \mul_out5[10] , 
        \mul_out5[9] , \mul_out5[8] , \mul_out5[7] , \mul_out5[6] , 
        \mul_out5[5] , \mul_out5[4] , \mul_out5[3] , \mul_out5[2] , 
        \mul_out5[1] , \mul_out5[0] }), .CI(1'b0), .SUM(add_r5) );
  datapath_DW_mult_tc_26 mult_118 ( .a(data_out_a6), .b({n2144, n2141, n2138, 
        n2, n2131, n571, n2032, n2123}), .product({\mul_out6[15] , 
        \mul_out6[14] , \mul_out6[13] , \mul_out6[12] , \mul_out6[11] , 
        \mul_out6[10] , \mul_out6[9] , \mul_out6[8] , \mul_out6[7] , 
        \mul_out6[6] , \mul_out6[5] , \mul_out6[4] , \mul_out6[3] , 
        \mul_out6[2] , \mul_out6[1] , \mul_out6[0] }) );
  datapath_DW01_add_26 add_119 ( .A(f6), .B({\mul_out6[15] , \mul_out6[14] , 
        \mul_out6[13] , \mul_out6[12] , \mul_out6[11] , \mul_out6[10] , 
        \mul_out6[9] , \mul_out6[8] , \mul_out6[7] , \mul_out6[6] , 
        \mul_out6[5] , \mul_out6[4] , \mul_out6[3] , \mul_out6[2] , 
        \mul_out6[1] , \mul_out6[0] }), .CI(1'b0), .SUM(add_r6) );
  datapath_DW_mult_tc_25 mult_120 ( .a(data_out_a7), .b({n2144, n2141, n2138, 
        n2134, n558, n9, n2126, n2121}), .product({\mul_out7[15] , 
        \mul_out7[14] , \mul_out7[13] , \mul_out7[12] , \mul_out7[11] , 
        \mul_out7[10] , \mul_out7[9] , \mul_out7[8] , \mul_out7[7] , 
        \mul_out7[6] , \mul_out7[5] , \mul_out7[4] , \mul_out7[3] , 
        \mul_out7[2] , \mul_out7[1] , \mul_out7[0] }) );
  datapath_DW01_add_25 add_121 ( .A(f7), .B({\mul_out7[15] , \mul_out7[14] , 
        \mul_out7[13] , \mul_out7[12] , \mul_out7[11] , \mul_out7[10] , 
        \mul_out7[9] , \mul_out7[8] , \mul_out7[7] , \mul_out7[6] , 
        \mul_out7[5] , \mul_out7[4] , \mul_out7[3] , \mul_out7[2] , 
        \mul_out7[1] , \mul_out7[0] }), .CI(1'b0), .SUM(add_r7) );
  datapath_DW_mult_tc_24 mult_122 ( .a(data_out_a8), .b({n2144, n2141, n2138, 
        n2133, n558, n571, n2124, n2121}), .product({\mul_out8[15] , 
        \mul_out8[14] , \mul_out8[13] , \mul_out8[12] , \mul_out8[11] , 
        \mul_out8[10] , \mul_out8[9] , \mul_out8[8] , \mul_out8[7] , 
        \mul_out8[6] , \mul_out8[5] , \mul_out8[4] , \mul_out8[3] , 
        \mul_out8[2] , \mul_out8[1] , \mul_out8[0] }) );
  datapath_DW01_add_24 add_123 ( .A(f8), .B({\mul_out8[15] , \mul_out8[14] , 
        \mul_out8[13] , \mul_out8[12] , \mul_out8[11] , \mul_out8[10] , 
        \mul_out8[9] , \mul_out8[8] , \mul_out8[7] , \mul_out8[6] , 
        \mul_out8[5] , \mul_out8[4] , \mul_out8[3] , \mul_out8[2] , 
        \mul_out8[1] , \mul_out8[0] }), .CI(1'b0), .SUM(add_r8) );
  datapath_DW_mult_tc_23 mult_124 ( .a(data_out_a9), .b({n2143, n2140, n2137, 
        n2135, n2132, n19, n2034, n2123}), .product({\mul_out9[15] , 
        \mul_out9[14] , \mul_out9[13] , \mul_out9[12] , \mul_out9[11] , 
        \mul_out9[10] , \mul_out9[9] , \mul_out9[8] , \mul_out9[7] , 
        \mul_out9[6] , \mul_out9[5] , \mul_out9[4] , \mul_out9[3] , 
        \mul_out9[2] , \mul_out9[1] , \mul_out9[0] }) );
  datapath_DW01_add_23 add_125 ( .A(f9), .B({\mul_out9[15] , \mul_out9[14] , 
        \mul_out9[13] , \mul_out9[12] , \mul_out9[11] , \mul_out9[10] , 
        \mul_out9[9] , \mul_out9[8] , \mul_out9[7] , \mul_out9[6] , 
        \mul_out9[5] , \mul_out9[4] , \mul_out9[3] , \mul_out9[2] , 
        \mul_out9[1] , \mul_out9[0] }), .CI(1'b0), .SUM(add_r9) );
  datapath_DW_mult_tc_22 mult_126 ( .a(data_out_a10), .b({n2143, n2140, n2137, 
        n2134, n2131, n20, n2034, n2121}), .product({\mul_out10[15] , 
        \mul_out10[14] , \mul_out10[13] , \mul_out10[12] , \mul_out10[11] , 
        \mul_out10[10] , \mul_out10[9] , \mul_out10[8] , \mul_out10[7] , 
        \mul_out10[6] , \mul_out10[5] , \mul_out10[4] , \mul_out10[3] , 
        \mul_out10[2] , \mul_out10[1] , \mul_out10[0] }) );
  datapath_DW01_add_22 add_127 ( .A(f10), .B({\mul_out10[15] , \mul_out10[14] , 
        \mul_out10[13] , \mul_out10[12] , \mul_out10[11] , \mul_out10[10] , 
        \mul_out10[9] , \mul_out10[8] , \mul_out10[7] , \mul_out10[6] , 
        \mul_out10[5] , \mul_out10[4] , \mul_out10[3] , \mul_out10[2] , 
        \mul_out10[1] , \mul_out10[0] }), .CI(1'b0), .SUM(add_r10) );
  datapath_DW_mult_tc_21 mult_128 ( .a(data_out_a11), .b({n2143, n2140, n2137, 
        n2133, n557, n32, n2032, n2123}), .product({\mul_out11[15] , 
        \mul_out11[14] , \mul_out11[13] , \mul_out11[12] , \mul_out11[11] , 
        \mul_out11[10] , \mul_out11[9] , \mul_out11[8] , \mul_out11[7] , 
        \mul_out11[6] , \mul_out11[5] , \mul_out11[4] , \mul_out11[3] , 
        \mul_out11[2] , \mul_out11[1] , \mul_out11[0] }) );
  datapath_DW01_add_21 add_129 ( .A(f11), .B({\mul_out11[15] , \mul_out11[14] , 
        \mul_out11[13] , \mul_out11[12] , \mul_out11[11] , \mul_out11[10] , 
        \mul_out11[9] , \mul_out11[8] , \mul_out11[7] , \mul_out11[6] , 
        \mul_out11[5] , \mul_out11[4] , \mul_out11[3] , \mul_out11[2] , 
        \mul_out11[1] , \mul_out11[0] }), .CI(1'b0), .SUM(add_r11) );
  datapath_DW_mult_tc_20 mult_130 ( .a(data_out_a12), .b({n2143, n2140, n2137, 
        n2, n16, n32, n2027, n2122}), .product({\mul_out12[15] , 
        \mul_out12[14] , \mul_out12[13] , \mul_out12[12] , \mul_out12[11] , 
        \mul_out12[10] , \mul_out12[9] , \mul_out12[8] , \mul_out12[7] , 
        \mul_out12[6] , \mul_out12[5] , \mul_out12[4] , \mul_out12[3] , 
        \mul_out12[2] , \mul_out12[1] , \mul_out12[0] }) );
  datapath_DW01_add_20 add_131 ( .A(f12), .B({\mul_out12[15] , \mul_out12[14] , 
        \mul_out12[13] , \mul_out12[12] , \mul_out12[11] , \mul_out12[10] , 
        \mul_out12[9] , \mul_out12[8] , \mul_out12[7] , \mul_out12[6] , 
        \mul_out12[5] , \mul_out12[4] , \mul_out12[3] , \mul_out12[2] , 
        \mul_out12[1] , \mul_out12[0] }), .CI(1'b0), .SUM(add_r12) );
  datapath_DW_mult_tc_19 mult_132 ( .a(data_out_a13), .b({n2143, n2140, n2137, 
        n2133, n558, n19, n2126, n2123}), .product({\mul_out13[15] , 
        \mul_out13[14] , \mul_out13[13] , \mul_out13[12] , \mul_out13[11] , 
        \mul_out13[10] , \mul_out13[9] , \mul_out13[8] , \mul_out13[7] , 
        \mul_out13[6] , \mul_out13[5] , \mul_out13[4] , \mul_out13[3] , 
        \mul_out13[2] , \mul_out13[1] , \mul_out13[0] }) );
  datapath_DW01_add_19 add_133 ( .A(f13), .B({\mul_out13[15] , \mul_out13[14] , 
        \mul_out13[13] , \mul_out13[12] , \mul_out13[11] , \mul_out13[10] , 
        \mul_out13[9] , \mul_out13[8] , \mul_out13[7] , \mul_out13[6] , 
        \mul_out13[5] , \mul_out13[4] , \mul_out13[3] , \mul_out13[2] , 
        \mul_out13[1] , \mul_out13[0] }), .CI(1'b0), .SUM(add_r13) );
  datapath_DW_mult_tc_18 mult_134 ( .a(data_out_a14), .b({n2143, n2140, n2137, 
        n2135, n2131, n19, n2027, n2123}), .product({\mul_out14[15] , 
        \mul_out14[14] , \mul_out14[13] , \mul_out14[12] , \mul_out14[11] , 
        \mul_out14[10] , \mul_out14[9] , \mul_out14[8] , \mul_out14[7] , 
        \mul_out14[6] , \mul_out14[5] , \mul_out14[4] , \mul_out14[3] , 
        \mul_out14[2] , \mul_out14[1] , \mul_out14[0] }) );
  datapath_DW01_add_18 add_135 ( .A(f14), .B({\mul_out14[15] , \mul_out14[14] , 
        \mul_out14[13] , \mul_out14[12] , \mul_out14[11] , \mul_out14[10] , 
        \mul_out14[9] , \mul_out14[8] , \mul_out14[7] , \mul_out14[6] , 
        \mul_out14[5] , \mul_out14[4] , \mul_out14[3] , \mul_out14[2] , 
        \mul_out14[1] , \mul_out14[0] }), .CI(1'b0), .SUM(add_r14) );
  datapath_DW_mult_tc_17 mult_136 ( .a(data_out_a15), .b({n2143, n2140, n2137, 
        n2, n17, n32, n4, n2122}), .product({\mul_out15[15] , \mul_out15[14] , 
        \mul_out15[13] , \mul_out15[12] , \mul_out15[11] , \mul_out15[10] , 
        \mul_out15[9] , \mul_out15[8] , \mul_out15[7] , \mul_out15[6] , 
        \mul_out15[5] , \mul_out15[4] , \mul_out15[3] , \mul_out15[2] , 
        \mul_out15[1] , \mul_out15[0] }) );
  datapath_DW01_add_17 add_137 ( .A(f15), .B({\mul_out15[15] , \mul_out15[14] , 
        \mul_out15[13] , \mul_out15[12] , \mul_out15[11] , \mul_out15[10] , 
        \mul_out15[9] , \mul_out15[8] , \mul_out15[7] , \mul_out15[6] , 
        \mul_out15[5] , \mul_out15[4] , \mul_out15[3] , \mul_out15[2] , 
        \mul_out15[1] , \mul_out15[0] }), .CI(1'b0), .SUM(add_r15) );
  datapath_DW_mult_tc_16 mult_138 ( .a(data_out_a16), .b({n2143, n2140, n2137, 
        n2, n16, n545, n2028, n2121}), .product({\mul_out16[15] , 
        \mul_out16[14] , \mul_out16[13] , \mul_out16[12] , \mul_out16[11] , 
        \mul_out16[10] , \mul_out16[9] , \mul_out16[8] , \mul_out16[7] , 
        \mul_out16[6] , \mul_out16[5] , \mul_out16[4] , \mul_out16[3] , 
        \mul_out16[2] , \mul_out16[1] , \mul_out16[0] }) );
  datapath_DW01_add_16 add_139 ( .A(f16), .B({\mul_out16[15] , \mul_out16[14] , 
        \mul_out16[13] , \mul_out16[12] , \mul_out16[11] , \mul_out16[10] , 
        \mul_out16[9] , \mul_out16[8] , \mul_out16[7] , \mul_out16[6] , 
        \mul_out16[5] , \mul_out16[4] , \mul_out16[3] , \mul_out16[2] , 
        \mul_out16[1] , \mul_out16[0] }), .CI(1'b0), .SUM(add_r16) );
  datapath_DW_mult_tc_15 mult_140 ( .a(data_out_a17), .b({n2143, n2140, n2137, 
        n2134, n2132, n19, n2032, n2121}), .product({\mul_out17[15] , 
        \mul_out17[14] , \mul_out17[13] , \mul_out17[12] , \mul_out17[11] , 
        \mul_out17[10] , \mul_out17[9] , \mul_out17[8] , \mul_out17[7] , 
        \mul_out17[6] , \mul_out17[5] , \mul_out17[4] , \mul_out17[3] , 
        \mul_out17[2] , \mul_out17[1] , \mul_out17[0] }) );
  datapath_DW01_add_15 add_141 ( .A(f17), .B({\mul_out17[15] , \mul_out17[14] , 
        \mul_out17[13] , \mul_out17[12] , \mul_out17[11] , \mul_out17[10] , 
        \mul_out17[9] , \mul_out17[8] , \mul_out17[7] , \mul_out17[6] , 
        \mul_out17[5] , \mul_out17[4] , \mul_out17[3] , \mul_out17[2] , 
        \mul_out17[1] , \mul_out17[0] }), .CI(1'b0), .SUM(add_r17) );
  datapath_DW_mult_tc_14 mult_142 ( .a(data_out_a18), .b({n2143, n2140, n2137, 
        n2135, n16, n545, n2033, n2123}), .product({\mul_out18[15] , 
        \mul_out18[14] , \mul_out18[13] , \mul_out18[12] , \mul_out18[11] , 
        \mul_out18[10] , \mul_out18[9] , \mul_out18[8] , \mul_out18[7] , 
        \mul_out18[6] , \mul_out18[5] , \mul_out18[4] , \mul_out18[3] , 
        \mul_out18[2] , \mul_out18[1] , \mul_out18[0] }) );
  datapath_DW01_add_14 add_143 ( .A(f18), .B({\mul_out18[15] , \mul_out18[14] , 
        \mul_out18[13] , \mul_out18[12] , \mul_out18[11] , \mul_out18[10] , 
        \mul_out18[9] , \mul_out18[8] , \mul_out18[7] , \mul_out18[6] , 
        \mul_out18[5] , \mul_out18[4] , \mul_out18[3] , \mul_out18[2] , 
        \mul_out18[1] , \mul_out18[0] }), .CI(1'b0), .SUM(add_r18) );
  datapath_DW_mult_tc_13 mult_144 ( .a(data_out_a19), .b({n2143, n2140, n2137, 
        n2135, n2131, n20, n2033, n2122}), .product({\mul_out19[15] , 
        \mul_out19[14] , \mul_out19[13] , \mul_out19[12] , \mul_out19[11] , 
        \mul_out19[10] , \mul_out19[9] , \mul_out19[8] , \mul_out19[7] , 
        \mul_out19[6] , \mul_out19[5] , \mul_out19[4] , \mul_out19[3] , 
        \mul_out19[2] , \mul_out19[1] , \mul_out19[0] }) );
  datapath_DW01_add_13 add_145 ( .A(f19), .B({\mul_out19[15] , \mul_out19[14] , 
        \mul_out19[13] , \mul_out19[12] , \mul_out19[11] , \mul_out19[10] , 
        \mul_out19[9] , \mul_out19[8] , \mul_out19[7] , \mul_out19[6] , 
        \mul_out19[5] , \mul_out19[4] , \mul_out19[3] , \mul_out19[2] , 
        \mul_out19[1] , \mul_out19[0] }), .CI(1'b0), .SUM(add_r19) );
  datapath_DW_mult_tc_12 mult_146 ( .a(data_out_a20), .b({n2143, n2140, n2137, 
        n2135, n557, n545, n2027, n2122}), .product({\mul_out20[15] , 
        \mul_out20[14] , \mul_out20[13] , \mul_out20[12] , \mul_out20[11] , 
        \mul_out20[10] , \mul_out20[9] , \mul_out20[8] , \mul_out20[7] , 
        \mul_out20[6] , \mul_out20[5] , \mul_out20[4] , \mul_out20[3] , 
        \mul_out20[2] , \mul_out20[1] , \mul_out20[0] }) );
  datapath_DW01_add_12 add_147 ( .A(f20), .B({\mul_out20[15] , \mul_out20[14] , 
        \mul_out20[13] , \mul_out20[12] , \mul_out20[11] , \mul_out20[10] , 
        \mul_out20[9] , \mul_out20[8] , \mul_out20[7] , \mul_out20[6] , 
        \mul_out20[5] , \mul_out20[4] , \mul_out20[3] , \mul_out20[2] , 
        \mul_out20[1] , \mul_out20[0] }), .CI(1'b0), .SUM(add_r20) );
  datapath_DW_mult_tc_11 mult_148 ( .a(data_out_a21), .b({n2142, n2139, n2136, 
        n2134, n15, n23, n2029, n2123}), .product({\mul_out21[15] , 
        \mul_out21[14] , \mul_out21[13] , \mul_out21[12] , \mul_out21[11] , 
        \mul_out21[10] , \mul_out21[9] , \mul_out21[8] , \mul_out21[7] , 
        \mul_out21[6] , \mul_out21[5] , \mul_out21[4] , \mul_out21[3] , 
        \mul_out21[2] , \mul_out21[1] , \mul_out21[0] }) );
  datapath_DW01_add_11 add_149 ( .A(f21), .B({\mul_out21[15] , \mul_out21[14] , 
        \mul_out21[13] , \mul_out21[12] , \mul_out21[11] , \mul_out21[10] , 
        \mul_out21[9] , \mul_out21[8] , \mul_out21[7] , \mul_out21[6] , 
        \mul_out21[5] , \mul_out21[4] , \mul_out21[3] , \mul_out21[2] , 
        \mul_out21[1] , \mul_out21[0] }), .CI(1'b0), .SUM(add_r21) );
  datapath_DW_mult_tc_10 mult_150 ( .a(data_out_a22), .b({n2142, n2139, n2136, 
        n2134, n2132, n23, n2124, n2122}), .product({\mul_out22[15] , 
        \mul_out22[14] , \mul_out22[13] , \mul_out22[12] , \mul_out22[11] , 
        \mul_out22[10] , \mul_out22[9] , \mul_out22[8] , \mul_out22[7] , 
        \mul_out22[6] , \mul_out22[5] , \mul_out22[4] , \mul_out22[3] , 
        \mul_out22[2] , \mul_out22[1] , \mul_out22[0] }) );
  datapath_DW01_add_10 add_151 ( .A(f22), .B({\mul_out22[15] , \mul_out22[14] , 
        \mul_out22[13] , \mul_out22[12] , \mul_out22[11] , \mul_out22[10] , 
        \mul_out22[9] , \mul_out22[8] , \mul_out22[7] , \mul_out22[6] , 
        \mul_out22[5] , \mul_out22[4] , \mul_out22[3] , \mul_out22[2] , 
        \mul_out22[1] , \mul_out22[0] }), .CI(1'b0), .SUM(add_r22) );
  datapath_DW_mult_tc_9 mult_152 ( .a(data_out_a23), .b({n2142, n2139, n2136, 
        n2133, n557, n9, n2029, n2122}), .product({\mul_out23[15] , 
        \mul_out23[14] , \mul_out23[13] , \mul_out23[12] , \mul_out23[11] , 
        \mul_out23[10] , \mul_out23[9] , \mul_out23[8] , \mul_out23[7] , 
        \mul_out23[6] , \mul_out23[5] , \mul_out23[4] , \mul_out23[3] , 
        \mul_out23[2] , \mul_out23[1] , \mul_out23[0] }) );
  datapath_DW01_add_9 add_153 ( .A(f23), .B({\mul_out23[15] , \mul_out23[14] , 
        \mul_out23[13] , \mul_out23[12] , \mul_out23[11] , \mul_out23[10] , 
        \mul_out23[9] , \mul_out23[8] , \mul_out23[7] , \mul_out23[6] , 
        \mul_out23[5] , \mul_out23[4] , \mul_out23[3] , \mul_out23[2] , 
        \mul_out23[1] , \mul_out23[0] }), .CI(1'b0), .SUM(add_r23) );
  datapath_DW_mult_tc_8 mult_154 ( .a(data_out_a24), .b({n2142, n2139, n2136, 
        n2133, n557, n24, n2028, n2121}), .product({\mul_out24[15] , 
        \mul_out24[14] , \mul_out24[13] , \mul_out24[12] , \mul_out24[11] , 
        \mul_out24[10] , \mul_out24[9] , \mul_out24[8] , \mul_out24[7] , 
        \mul_out24[6] , \mul_out24[5] , \mul_out24[4] , \mul_out24[3] , 
        \mul_out24[2] , \mul_out24[1] , \mul_out24[0] }) );
  datapath_DW01_add_8 add_155 ( .A(f24), .B({\mul_out24[15] , \mul_out24[14] , 
        \mul_out24[13] , \mul_out24[12] , \mul_out24[11] , \mul_out24[10] , 
        \mul_out24[9] , \mul_out24[8] , \mul_out24[7] , \mul_out24[6] , 
        \mul_out24[5] , \mul_out24[4] , \mul_out24[3] , \mul_out24[2] , 
        \mul_out24[1] , \mul_out24[0] }), .CI(1'b0), .SUM(add_r24) );
  datapath_DW_mult_tc_7 mult_156 ( .a(data_out_a25), .b({n2142, n2139, n2136, 
        n2133, n2131, n24, n2028, n2121}), .product({\mul_out25[15] , 
        \mul_out25[14] , \mul_out25[13] , \mul_out25[12] , \mul_out25[11] , 
        \mul_out25[10] , \mul_out25[9] , \mul_out25[8] , \mul_out25[7] , 
        \mul_out25[6] , \mul_out25[5] , \mul_out25[4] , \mul_out25[3] , 
        \mul_out25[2] , \mul_out25[1] , \mul_out25[0] }) );
  datapath_DW01_add_7 add_157 ( .A(f25), .B({\mul_out25[15] , \mul_out25[14] , 
        \mul_out25[13] , \mul_out25[12] , \mul_out25[11] , \mul_out25[10] , 
        \mul_out25[9] , \mul_out25[8] , \mul_out25[7] , \mul_out25[6] , 
        \mul_out25[5] , \mul_out25[4] , \mul_out25[3] , \mul_out25[2] , 
        \mul_out25[1] , \mul_out25[0] }), .CI(1'b0), .SUM(add_r25) );
  datapath_DW_mult_tc_6 mult_158 ( .a(data_out_a26), .b({n2142, n2139, n2136, 
        n2133, n558, n20, n2126, n2123}), .product({\mul_out26[15] , 
        \mul_out26[14] , \mul_out26[13] , \mul_out26[12] , \mul_out26[11] , 
        \mul_out26[10] , \mul_out26[9] , \mul_out26[8] , \mul_out26[7] , 
        \mul_out26[6] , \mul_out26[5] , \mul_out26[4] , \mul_out26[3] , 
        \mul_out26[2] , \mul_out26[1] , \mul_out26[0] }) );
  datapath_DW01_add_6 add_159 ( .A(f26), .B({\mul_out26[15] , \mul_out26[14] , 
        \mul_out26[13] , \mul_out26[12] , \mul_out26[11] , \mul_out26[10] , 
        \mul_out26[9] , \mul_out26[8] , \mul_out26[7] , \mul_out26[6] , 
        \mul_out26[5] , \mul_out26[4] , \mul_out26[3] , \mul_out26[2] , 
        \mul_out26[1] , \mul_out26[0] }), .CI(1'b0), .SUM(add_r26) );
  datapath_DW_mult_tc_5 mult_160 ( .a(data_out_a27), .b({n2142, n2139, n2136, 
        n2134, n17, n25, n2034, n2122}), .product({\mul_out27[15] , 
        \mul_out27[14] , \mul_out27[13] , \mul_out27[12] , \mul_out27[11] , 
        \mul_out27[10] , \mul_out27[9] , \mul_out27[8] , \mul_out27[7] , 
        \mul_out27[6] , \mul_out27[5] , \mul_out27[4] , \mul_out27[3] , 
        \mul_out27[2] , \mul_out27[1] , \mul_out27[0] }) );
  datapath_DW01_add_5 add_161 ( .A(f27), .B({\mul_out27[15] , \mul_out27[14] , 
        \mul_out27[13] , \mul_out27[12] , \mul_out27[11] , \mul_out27[10] , 
        \mul_out27[9] , \mul_out27[8] , \mul_out27[7] , \mul_out27[6] , 
        \mul_out27[5] , \mul_out27[4] , \mul_out27[3] , \mul_out27[2] , 
        \mul_out27[1] , \mul_out27[0] }), .CI(1'b0), .SUM(add_r27) );
  datapath_DW_mult_tc_4 mult_162 ( .a(data_out_a28), .b({n2142, n2139, n2136, 
        n2133, n2132, n5, n2126, n2121}), .product({\mul_out28[15] , 
        \mul_out28[14] , \mul_out28[13] , \mul_out28[12] , \mul_out28[11] , 
        \mul_out28[10] , \mul_out28[9] , \mul_out28[8] , \mul_out28[7] , 
        \mul_out28[6] , \mul_out28[5] , \mul_out28[4] , \mul_out28[3] , 
        \mul_out28[2] , \mul_out28[1] , \mul_out28[0] }) );
  datapath_DW01_add_4 add_163 ( .A(f28), .B({\mul_out28[15] , \mul_out28[14] , 
        \mul_out28[13] , \mul_out28[12] , \mul_out28[11] , \mul_out28[10] , 
        \mul_out28[9] , \mul_out28[8] , \mul_out28[7] , \mul_out28[6] , 
        \mul_out28[5] , \mul_out28[4] , \mul_out28[3] , \mul_out28[2] , 
        \mul_out28[1] , \mul_out28[0] }), .CI(1'b0), .SUM(add_r28) );
  datapath_DW_mult_tc_3 mult_164 ( .a(data_out_a29), .b({n2142, n2139, n2136, 
        n2134, n17, n5, n2033, n2122}), .product({\mul_out29[15] , 
        \mul_out29[14] , \mul_out29[13] , \mul_out29[12] , \mul_out29[11] , 
        \mul_out29[10] , \mul_out29[9] , \mul_out29[8] , \mul_out29[7] , 
        \mul_out29[6] , \mul_out29[5] , \mul_out29[4] , \mul_out29[3] , 
        \mul_out29[2] , \mul_out29[1] , \mul_out29[0] }) );
  datapath_DW01_add_3 add_165 ( .A(f29), .B({\mul_out29[15] , \mul_out29[14] , 
        \mul_out29[13] , \mul_out29[12] , \mul_out29[11] , \mul_out29[10] , 
        \mul_out29[9] , \mul_out29[8] , \mul_out29[7] , \mul_out29[6] , 
        \mul_out29[5] , \mul_out29[4] , \mul_out29[3] , \mul_out29[2] , 
        \mul_out29[1] , \mul_out29[0] }), .CI(1'b0), .SUM(add_r29) );
  datapath_DW_mult_tc_2 mult_166 ( .a(data_out_a30), .b({n2142, n2139, n2136, 
        n2135, n558, n25, n2029, n2123}), .product({\mul_out30[15] , 
        \mul_out30[14] , \mul_out30[13] , \mul_out30[12] , \mul_out30[11] , 
        \mul_out30[10] , \mul_out30[9] , \mul_out30[8] , \mul_out30[7] , 
        \mul_out30[6] , \mul_out30[5] , \mul_out30[4] , \mul_out30[3] , 
        \mul_out30[2] , \mul_out30[1] , \mul_out30[0] }) );
  datapath_DW01_add_2 add_167 ( .A(f30), .B({\mul_out30[15] , \mul_out30[14] , 
        \mul_out30[13] , \mul_out30[12] , \mul_out30[11] , \mul_out30[10] , 
        \mul_out30[9] , \mul_out30[8] , \mul_out30[7] , \mul_out30[6] , 
        \mul_out30[5] , \mul_out30[4] , \mul_out30[3] , \mul_out30[2] , 
        \mul_out30[1] , \mul_out30[0] }), .CI(1'b0), .SUM(add_r30) );
  datapath_DW_mult_tc_1 mult_168 ( .a(data_out_a31), .b({n2142, n2139, n2136, 
        n2, n558, n5, n2126, n2122}), .product({\mul_out31[15] , 
        \mul_out31[14] , \mul_out31[13] , \mul_out31[12] , \mul_out31[11] , 
        \mul_out31[10] , \mul_out31[9] , \mul_out31[8] , \mul_out31[7] , 
        \mul_out31[6] , \mul_out31[5] , \mul_out31[4] , \mul_out31[3] , 
        \mul_out31[2] , \mul_out31[1] , \mul_out31[0] }) );
  datapath_DW01_add_1 add_169 ( .A(f31), .B({\mul_out31[15] , \mul_out31[14] , 
        \mul_out31[13] , \mul_out31[12] , \mul_out31[11] , \mul_out31[10] , 
        \mul_out31[9] , \mul_out31[8] , \mul_out31[7] , \mul_out31[6] , 
        \mul_out31[5] , \mul_out31[4] , \mul_out31[3] , \mul_out31[2] , 
        \mul_out31[1] , \mul_out31[0] }), .CI(1'b0), .SUM(add_r31) );
  datapath_DW_mult_tc_0 mult_170 ( .a(data_out_a32), .b({n2142, n2139, n2136, 
        n2, n2131, n23, n2032, n2123}), .product({\mul_out32[15] , 
        \mul_out32[14] , \mul_out32[13] , \mul_out32[12] , \mul_out32[11] , 
        \mul_out32[10] , \mul_out32[9] , \mul_out32[8] , \mul_out32[7] , 
        \mul_out32[6] , \mul_out32[5] , \mul_out32[4] , \mul_out32[3] , 
        \mul_out32[2] , \mul_out32[1] , \mul_out32[0] }) );
  datapath_DW01_add_0 add_171 ( .A(f32), .B({\mul_out32[15] , \mul_out32[14] , 
        \mul_out32[13] , \mul_out32[12] , \mul_out32[11] , \mul_out32[10] , 
        \mul_out32[9] , \mul_out32[8] , \mul_out32[7] , \mul_out32[6] , 
        \mul_out32[5] , \mul_out32[4] , \mul_out32[3] , \mul_out32[2] , 
        \mul_out32[1] , \mul_out32[0] }), .CI(1'b0), .SUM(add_r32) );
  DFF_X1 \f31_reg[15]  ( .D(n1546), .CK(clk), .Q(f31[15]), .QN(n513) );
  DFF_X1 \f6_reg[15]  ( .D(n1946), .CK(clk), .Q(f6[15]), .QN(n113) );
  DFF_X1 \f17_reg[15]  ( .D(n1770), .CK(clk), .Q(f17[15]), .QN(n289) );
  DFF_X1 \f3_reg[15]  ( .D(n1994), .CK(clk), .Q(f3[15]), .QN(n65) );
  DFF_X1 \f2_reg[15]  ( .D(n2010), .CK(clk), .Q(f2[15]), .QN(n49) );
  DFF_X1 \f30_reg[15]  ( .D(n1562), .CK(clk), .Q(f30[15]), .QN(n497) );
  DFF_X1 \f7_reg[15]  ( .D(n1930), .CK(clk), .Q(f7[15]), .QN(n129) );
  DFF_X1 \f15_reg[15]  ( .D(n1802), .CK(clk), .Q(f15[15]), .QN(n257) );
  DFF_X1 \f20_reg[15]  ( .D(n1722), .CK(clk), .Q(f20[15]), .QN(n337) );
  DFF_X1 \f10_reg[15]  ( .D(n1882), .CK(clk), .Q(f10[15]), .QN(n177) );
  DFF_X1 \f9_reg[15]  ( .D(n1898), .CK(clk), .Q(f9[15]), .QN(n161) );
  DFF_X1 \f19_reg[15]  ( .D(n1738), .CK(clk), .Q(f19[15]), .QN(n321) );
  DFF_X1 \f14_reg[15]  ( .D(n1818), .CK(clk), .Q(f14[15]), .QN(n241) );
  DFF_X1 \f18_reg[15]  ( .D(n1754), .CK(clk), .Q(f18[15]), .QN(n305) );
  DFF_X1 \f13_reg[15]  ( .D(n1834), .CK(clk), .Q(f13[15]), .QN(n225) );
  DFF_X1 \f29_reg[15]  ( .D(n1578), .CK(clk), .Q(f29[15]), .QN(n481) );
  DFF_X1 \f12_reg[15]  ( .D(n1850), .CK(clk), .Q(f12[15]), .QN(n209) );
  DFF_X1 \f22_reg[15]  ( .D(n1690), .CK(clk), .Q(f22[15]), .QN(n369) );
  DFF_X1 \f21_reg[15]  ( .D(n1706), .CK(clk), .Q(f21[15]), .QN(n353) );
  DFF_X1 \f26_reg[15]  ( .D(n1626), .CK(clk), .Q(f26[15]), .QN(n433) );
  DFF_X1 \f5_reg[15]  ( .D(n1962), .CK(clk), .Q(f5[15]), .QN(n97) );
  DFF_X1 \f16_reg[14]  ( .D(n1785), .CK(clk), .Q(f16[14]), .QN(n274) );
  DFF_X1 \f25_reg[15]  ( .D(n1642), .CK(clk), .Q(f25[15]), .QN(n417) );
  CLKBUF_X3 U3 ( .A(n2129), .Z(n570) );
  CLKBUF_X3 U4 ( .A(n2125), .Z(n2033) );
  BUF_X2 U5 ( .A(data_out_x[1]), .Z(n2125) );
  BUF_X1 U6 ( .A(data_out_x[2]), .Z(n2129) );
  BUF_X2 U7 ( .A(n2128), .Z(n545) );
  NOR2_X1 U8 ( .A1(n2149), .A2(addr_y[0]), .ZN(n947) );
  BUF_X2 U9 ( .A(n2127), .Z(n25) );
  CLKBUF_X3 U10 ( .A(n2128), .Z(n19) );
  CLKBUF_X3 U11 ( .A(n2129), .Z(n571) );
  OR2_X1 U12 ( .A1(n2091), .A2(n497), .ZN(n21) );
  OR2_X1 U13 ( .A1(n2112), .A2(n113), .ZN(n26) );
  OR2_X1 U14 ( .A1(n2094), .A2(n466), .ZN(n8) );
  OR2_X1 U15 ( .A1(n2095), .A2(n449), .ZN(n12) );
  OR2_X1 U16 ( .A1(n2097), .A2(n434), .ZN(n7) );
  OR2_X1 U17 ( .A1(n2099), .A2(n401), .ZN(n547) );
  OR2_X1 U18 ( .A1(n2101), .A2(n386), .ZN(n13) );
  OR2_X1 U19 ( .A1(n2108), .A2(n290), .ZN(n11) );
  OR2_X1 U20 ( .A1(n2112), .A2(n226), .ZN(n6) );
  OR2_X1 U21 ( .A1(n2117), .A2(n145), .ZN(n550) );
  AND2_X1 U22 ( .A1(n982), .A2(n1002), .ZN(n1) );
  BUF_X4 U23 ( .A(data_out_x[4]), .Z(n2133) );
  BUF_X4 U24 ( .A(data_out_x[4]), .Z(n2) );
  CLKBUF_X3 U25 ( .A(n2129), .Z(n9) );
  BUF_X2 U26 ( .A(n2029), .Z(n4) );
  BUF_X4 U27 ( .A(data_out_x[5]), .Z(n2138) );
  CLKBUF_X3 U28 ( .A(n2127), .Z(n24) );
  BUF_X1 U29 ( .A(n2029), .Z(n27) );
  BUF_X8 U30 ( .A(data_out_x[5]), .Z(n2136) );
  BUF_X4 U31 ( .A(data_out_x[4]), .Z(n2134) );
  OR2_X1 U32 ( .A1(n2098), .A2(n418), .ZN(n3) );
  NAND2_X1 U33 ( .A1(n3), .A2(n1113), .ZN(n1641) );
  BUF_X4 U34 ( .A(data_out_x[6]), .Z(n2141) );
  BUF_X8 U35 ( .A(data_out_x[6]), .Z(n2139) );
  BUF_X2 U36 ( .A(data_out_x[2]), .Z(n2128) );
  CLKBUF_X3 U37 ( .A(data_out_x[3]), .Z(n2131) );
  CLKBUF_X3 U38 ( .A(data_out_x[3]), .Z(n557) );
  CLKBUF_X3 U39 ( .A(data_out_x[3]), .Z(n2132) );
  CLKBUF_X1 U40 ( .A(data_out_x[3]), .Z(n2130) );
  BUF_X1 U41 ( .A(data_out_x[2]), .Z(n2127) );
  CLKBUF_X3 U42 ( .A(n2127), .Z(n5) );
  NAND2_X1 U43 ( .A1(n6), .A2(n1305), .ZN(n1833) );
  CLKBUF_X3 U44 ( .A(data_out_x[0]), .Z(n2123) );
  NAND2_X1 U45 ( .A1(n7), .A2(n1097), .ZN(n1625) );
  CLKBUF_X3 U46 ( .A(n2125), .Z(n2027) );
  NAND2_X1 U47 ( .A1(n8), .A2(n1065), .ZN(n1593) );
  OR2_X1 U48 ( .A1(n2090), .A2(n514), .ZN(n10) );
  NAND2_X1 U49 ( .A1(n1016), .A2(n10), .ZN(n1545) );
  NAND2_X1 U50 ( .A1(n11), .A2(n1241), .ZN(n1769) );
  BUF_X4 U51 ( .A(data_out_x[4]), .Z(n2135) );
  BUF_X4 U52 ( .A(data_out_x[3]), .Z(n558) );
  NAND2_X1 U53 ( .A1(n1082), .A2(n12), .ZN(n1610) );
  CLKBUF_X3 U54 ( .A(n2128), .Z(n20) );
  CLKBUF_X3 U55 ( .A(n2128), .Z(n32) );
  CLKBUF_X3 U56 ( .A(n2127), .Z(n23) );
  NAND2_X1 U57 ( .A1(n13), .A2(n1145), .ZN(n1673) );
  OR2_X1 U58 ( .A1(n2095), .A2(n450), .ZN(n14) );
  NAND2_X1 U59 ( .A1(n1081), .A2(n14), .ZN(n1609) );
  CLKBUF_X1 U60 ( .A(n2130), .Z(n15) );
  CLKBUF_X3 U61 ( .A(n2130), .Z(n16) );
  CLKBUF_X3 U62 ( .A(n2130), .Z(n17) );
  OR2_X1 U63 ( .A1(n2091), .A2(n498), .ZN(n18) );
  NAND2_X1 U64 ( .A1(n1033), .A2(n18), .ZN(n1561) );
  CLKBUF_X3 U65 ( .A(data_out_x[1]), .Z(n2126) );
  CLKBUF_X3 U66 ( .A(n2125), .Z(n2032) );
  NAND2_X1 U67 ( .A1(n1034), .A2(n21), .ZN(n1562) );
  CLKBUF_X3 U68 ( .A(n2125), .Z(n2034) );
  OR2_X1 U69 ( .A1(n2109), .A2(n274), .ZN(n22) );
  NAND2_X1 U70 ( .A1(n1257), .A2(n22), .ZN(n1785) );
  NAND2_X1 U71 ( .A1(n1418), .A2(n26), .ZN(n1946) );
  CLKBUF_X3 U72 ( .A(data_out_x[0]), .Z(n2122) );
  CLKBUF_X3 U73 ( .A(data_out_x[0]), .Z(n2121) );
  OR2_X1 U74 ( .A1(n2119), .A2(n81), .ZN(n28) );
  NAND2_X1 U75 ( .A1(n1450), .A2(n28), .ZN(n1978) );
  CLKBUF_X3 U76 ( .A(data_out_x[1]), .Z(n2029) );
  OR2_X1 U77 ( .A1(n2094), .A2(n465), .ZN(n29) );
  NAND2_X1 U78 ( .A1(n1066), .A2(n29), .ZN(n1594) );
  OR2_X1 U79 ( .A1(n2101), .A2(n385), .ZN(n30) );
  NAND2_X1 U80 ( .A1(n1146), .A2(n30), .ZN(n1674) );
  OR2_X1 U81 ( .A1(n2094), .A2(n97), .ZN(n31) );
  NAND2_X1 U82 ( .A1(n1434), .A2(n31), .ZN(n1962) );
  OR2_X1 U83 ( .A1(n2084), .A2(n33), .ZN(n546) );
  NAND2_X1 U84 ( .A1(n1498), .A2(n546), .ZN(n2026) );
  NAND2_X1 U85 ( .A1(n1130), .A2(n547), .ZN(n1658) );
  OR2_X1 U86 ( .A1(n2089), .A2(n529), .ZN(n548) );
  NAND2_X1 U87 ( .A1(n1000), .A2(n548), .ZN(n1530) );
  OR2_X1 U88 ( .A1(n2120), .A2(n65), .ZN(n549) );
  NAND2_X1 U89 ( .A1(n1466), .A2(n549), .ZN(n1994) );
  NAND2_X1 U90 ( .A1(n1386), .A2(n550), .ZN(n1914) );
  OR2_X1 U91 ( .A1(n2120), .A2(n49), .ZN(n551) );
  NAND2_X1 U92 ( .A1(n1482), .A2(n551), .ZN(n2010) );
  OR2_X1 U93 ( .A1(n2098), .A2(n417), .ZN(n552) );
  NAND2_X1 U94 ( .A1(n1114), .A2(n552), .ZN(n1642) );
  OR2_X1 U95 ( .A1(n2093), .A2(n481), .ZN(n553) );
  NAND2_X1 U96 ( .A1(n1050), .A2(n553), .ZN(n1578) );
  OR2_X1 U97 ( .A1(n2097), .A2(n433), .ZN(n554) );
  NAND2_X1 U98 ( .A1(n1098), .A2(n554), .ZN(n1626) );
  OR2_X1 U99 ( .A1(n2103), .A2(n353), .ZN(n555) );
  NAND2_X1 U100 ( .A1(n1178), .A2(n555), .ZN(n1706) );
  OR2_X1 U101 ( .A1(n2102), .A2(n369), .ZN(n556) );
  NAND2_X1 U102 ( .A1(n1162), .A2(n556), .ZN(n1690) );
  OR2_X1 U103 ( .A1(n2107), .A2(n305), .ZN(n559) );
  NAND2_X1 U104 ( .A1(n1226), .A2(n559), .ZN(n1754) );
  OR2_X1 U105 ( .A1(n2111), .A2(n241), .ZN(n560) );
  NAND2_X1 U106 ( .A1(n1290), .A2(n560), .ZN(n1818) );
  OR2_X1 U107 ( .A1(n2106), .A2(n321), .ZN(n561) );
  NAND2_X1 U108 ( .A1(n1210), .A2(n561), .ZN(n1738) );
  OR2_X1 U109 ( .A1(n2115), .A2(n161), .ZN(n562) );
  NAND2_X1 U110 ( .A1(n1370), .A2(n562), .ZN(n1898) );
  OR2_X1 U111 ( .A1(n2114), .A2(n177), .ZN(n563) );
  NAND2_X1 U112 ( .A1(n1354), .A2(n563), .ZN(n1882) );
  OR2_X1 U113 ( .A1(n2112), .A2(n225), .ZN(n564) );
  NAND2_X1 U114 ( .A1(n1306), .A2(n564), .ZN(n1834) );
  OR2_X1 U115 ( .A1(n2120), .A2(n209), .ZN(n565) );
  NAND2_X1 U116 ( .A1(n1322), .A2(n565), .ZN(n1850) );
  OR2_X1 U117 ( .A1(n2109), .A2(n273), .ZN(n566) );
  NAND2_X1 U118 ( .A1(n1258), .A2(n566), .ZN(n1786) );
  OR2_X1 U119 ( .A1(n2108), .A2(n289), .ZN(n567) );
  NAND2_X1 U120 ( .A1(n1242), .A2(n567), .ZN(n1770) );
  OR2_X1 U121 ( .A1(n2105), .A2(n337), .ZN(n568) );
  NAND2_X1 U122 ( .A1(n1194), .A2(n568), .ZN(n1722) );
  OR2_X1 U123 ( .A1(n2120), .A2(n257), .ZN(n569) );
  NAND2_X1 U124 ( .A1(n1274), .A2(n569), .ZN(n1802) );
  INV_X1 U125 ( .A(n966), .ZN(n2151) );
  BUF_X1 U126 ( .A(n2042), .Z(n2077) );
  BUF_X1 U127 ( .A(n2042), .Z(n2073) );
  BUF_X1 U128 ( .A(n2041), .Z(n2069) );
  BUF_X1 U129 ( .A(n2040), .Z(n2067) );
  BUF_X1 U130 ( .A(n2039), .Z(n2066) );
  BUF_X1 U131 ( .A(n2039), .Z(n2062) );
  BUF_X1 U132 ( .A(n2038), .Z(n2058) );
  BUF_X1 U133 ( .A(n2037), .Z(n2054) );
  BUF_X1 U134 ( .A(n2036), .Z(n2050) );
  BUF_X1 U135 ( .A(n2043), .Z(n2078) );
  BUF_X1 U136 ( .A(n2042), .Z(n2076) );
  BUF_X1 U137 ( .A(n2042), .Z(n2075) );
  BUF_X1 U138 ( .A(n2042), .Z(n2074) );
  BUF_X1 U139 ( .A(n2041), .Z(n2072) );
  BUF_X1 U140 ( .A(n2041), .Z(n2071) );
  BUF_X1 U141 ( .A(n2041), .Z(n2070) );
  BUF_X1 U142 ( .A(n2041), .Z(n2068) );
  BUF_X1 U143 ( .A(n2039), .Z(n2065) );
  BUF_X1 U144 ( .A(n2039), .Z(n2064) );
  BUF_X1 U145 ( .A(n2039), .Z(n2063) );
  BUF_X1 U146 ( .A(n2038), .Z(n2061) );
  BUF_X1 U147 ( .A(n2038), .Z(n2060) );
  BUF_X1 U148 ( .A(n2038), .Z(n2059) );
  BUF_X1 U149 ( .A(n2038), .Z(n2057) );
  BUF_X1 U150 ( .A(n2037), .Z(n2056) );
  BUF_X1 U151 ( .A(n2037), .Z(n2055) );
  BUF_X1 U152 ( .A(n2037), .Z(n2053) );
  BUF_X1 U153 ( .A(n2037), .Z(n2052) );
  BUF_X1 U154 ( .A(n2036), .Z(n2051) );
  BUF_X1 U155 ( .A(n2036), .Z(n2049) );
  BUF_X1 U156 ( .A(n2036), .Z(n2048) );
  BUF_X1 U157 ( .A(n2036), .Z(n2047) );
  BUF_X1 U158 ( .A(n2043), .Z(n2079) );
  BUF_X1 U159 ( .A(n2082), .Z(n2096) );
  BUF_X1 U160 ( .A(n2083), .Z(n2100) );
  BUF_X1 U161 ( .A(n2084), .Z(n2104) );
  BUF_X1 U162 ( .A(n2086), .Z(n2110) );
  BUF_X1 U163 ( .A(n2081), .Z(n2088) );
  BUF_X1 U164 ( .A(n2081), .Z(n2092) );
  BUF_X1 U165 ( .A(n2086), .Z(n2113) );
  BUF_X1 U166 ( .A(n2085), .Z(n2116) );
  BUF_X1 U167 ( .A(n2082), .Z(n2093) );
  BUF_X1 U168 ( .A(n2082), .Z(n2094) );
  BUF_X1 U169 ( .A(n2082), .Z(n2095) );
  BUF_X1 U170 ( .A(n2082), .Z(n2097) );
  BUF_X1 U171 ( .A(n2083), .Z(n2098) );
  BUF_X1 U172 ( .A(n2083), .Z(n2099) );
  BUF_X1 U173 ( .A(n2083), .Z(n2101) );
  BUF_X1 U174 ( .A(n2083), .Z(n2102) );
  BUF_X1 U175 ( .A(n2084), .Z(n2103) );
  BUF_X1 U176 ( .A(n2084), .Z(n2105) );
  BUF_X1 U177 ( .A(n2084), .Z(n2106) );
  BUF_X1 U178 ( .A(n2084), .Z(n2107) );
  BUF_X1 U179 ( .A(n2083), .Z(n2108) );
  BUF_X1 U180 ( .A(n2081), .Z(n2109) );
  BUF_X1 U181 ( .A(n2085), .Z(n2119) );
  BUF_X1 U182 ( .A(n2086), .Z(n2120) );
  BUF_X1 U183 ( .A(n2081), .Z(n2089) );
  BUF_X1 U184 ( .A(n2081), .Z(n2091) );
  BUF_X1 U185 ( .A(n2087), .Z(n2111) );
  BUF_X1 U186 ( .A(n2086), .Z(n2112) );
  BUF_X1 U187 ( .A(n2085), .Z(n2114) );
  BUF_X1 U188 ( .A(n2085), .Z(n2115) );
  BUF_X1 U189 ( .A(n2085), .Z(n2117) );
  AND2_X1 U190 ( .A1(n950), .A2(n2145), .ZN(n615) );
  NAND2_X1 U191 ( .A1(n949), .A2(n2145), .ZN(n602) );
  AND4_X1 U192 ( .A1(n940), .A2(n939), .A3(n941), .A4(n944), .ZN(n589) );
  NOR4_X1 U193 ( .A1(n2168), .A2(n2162), .A3(n583), .A4(n582), .ZN(n944) );
  INV_X1 U194 ( .A(n585), .ZN(n2168) );
  INV_X1 U195 ( .A(n586), .ZN(n2162) );
  INV_X1 U196 ( .A(n940), .ZN(n2166) );
  INV_X1 U197 ( .A(n955), .ZN(n2159) );
  INV_X1 U198 ( .A(n941), .ZN(n2167) );
  INV_X1 U199 ( .A(n954), .ZN(n2164) );
  INV_X1 U200 ( .A(n939), .ZN(n2161) );
  INV_X1 U201 ( .A(n975), .ZN(n2153) );
  BUF_X1 U202 ( .A(n2044), .Z(n2042) );
  BUF_X1 U203 ( .A(n2044), .Z(n2041) );
  BUF_X1 U204 ( .A(n2045), .Z(n2040) );
  BUF_X1 U205 ( .A(n2045), .Z(n2039) );
  BUF_X1 U206 ( .A(n2046), .Z(n2038) );
  BUF_X1 U207 ( .A(n2046), .Z(n2037) );
  BUF_X1 U208 ( .A(n2046), .Z(n2036) );
  NAND2_X1 U209 ( .A1(n945), .A2(n2145), .ZN(n966) );
  BUF_X1 U210 ( .A(n2044), .Z(n2043) );
  BUF_X1 U211 ( .A(n2087), .Z(n2082) );
  BUF_X1 U212 ( .A(n2087), .Z(n2083) );
  BUF_X1 U213 ( .A(n2086), .Z(n2084) );
  BUF_X1 U214 ( .A(n2087), .Z(n2085) );
  BUF_X1 U215 ( .A(n2087), .Z(n2081) );
  NAND4_X1 U216 ( .A1(n976), .A2(n975), .A3(n617), .A4(n977), .ZN(n618) );
  NOR4_X1 U217 ( .A1(n2155), .A2(n2152), .A3(n616), .A4(n615), .ZN(n977) );
  INV_X1 U218 ( .A(n612), .ZN(n2152) );
  INV_X1 U219 ( .A(n613), .ZN(n2155) );
  NAND2_X1 U220 ( .A1(n948), .A2(n2145), .ZN(n606) );
  NAND2_X1 U221 ( .A1(n957), .A2(n2145), .ZN(n612) );
  NAND2_X1 U222 ( .A1(n957), .A2(n947), .ZN(n590) );
  AND2_X1 U223 ( .A1(n945), .A2(n947), .ZN(n583) );
  AND2_X1 U224 ( .A1(n958), .A2(n947), .ZN(n593) );
  AND2_X1 U225 ( .A1(n969), .A2(n2145), .ZN(n605) );
  NAND2_X1 U226 ( .A1(n948), .A2(n946), .ZN(n586) );
  NAND2_X1 U227 ( .A1(n949), .A2(n947), .ZN(n585) );
  AND2_X1 U228 ( .A1(n945), .A2(n946), .ZN(n582) );
  NAND2_X1 U229 ( .A1(n958), .A2(n946), .ZN(n591) );
  NAND2_X1 U230 ( .A1(n979), .A2(n2158), .ZN(n572) );
  INV_X1 U231 ( .A(n980), .ZN(n2158) );
  NAND4_X1 U232 ( .A1(n966), .A2(n965), .A3(n606), .A4(n967), .ZN(n608) );
  NOR4_X1 U233 ( .A1(n605), .A2(n604), .A3(n2150), .A4(n2157), .ZN(n967) );
  INV_X1 U234 ( .A(n602), .ZN(n2150) );
  INV_X1 U235 ( .A(n601), .ZN(n2157) );
  AND2_X1 U236 ( .A1(n946), .A2(n957), .ZN(n594) );
  INV_X1 U237 ( .A(n976), .ZN(n2154) );
  INV_X1 U238 ( .A(n965), .ZN(n2156) );
  INV_X1 U239 ( .A(addr_y[0]), .ZN(n2145) );
  AND2_X1 U240 ( .A1(n979), .A2(n980), .ZN(n575) );
  NOR2_X1 U241 ( .A1(addr_y[1]), .A2(addr_y[2]), .ZN(n959) );
  AND2_X1 U242 ( .A1(n957), .A2(addr_y[3]), .ZN(n949) );
  NAND2_X1 U243 ( .A1(n969), .A2(n947), .ZN(n981) );
  AND2_X1 U244 ( .A1(n978), .A2(addr_y[2]), .ZN(n950) );
  NAND2_X1 U245 ( .A1(n950), .A2(n947), .ZN(n941) );
  NAND2_X1 U246 ( .A1(n959), .A2(n947), .ZN(n954) );
  NAND2_X1 U247 ( .A1(n948), .A2(n947), .ZN(n940) );
  NAND2_X1 U248 ( .A1(n950), .A2(n946), .ZN(n939) );
  NAND2_X1 U249 ( .A1(n958), .A2(n2145), .ZN(n975) );
  NAND2_X1 U250 ( .A1(n959), .A2(n946), .ZN(n955) );
  NAND2_X1 U251 ( .A1(n949), .A2(n946), .ZN(n980) );
  NAND4_X1 U252 ( .A1(n955), .A2(n954), .A3(n595), .A4(n956), .ZN(n597) );
  NOR4_X1 U253 ( .A1(n594), .A2(n593), .A3(n2160), .A4(n2165), .ZN(n956) );
  INV_X1 U254 ( .A(n590), .ZN(n2165) );
  INV_X1 U255 ( .A(n591), .ZN(n2160) );
  AND2_X1 U256 ( .A1(n970), .A2(addr_y[1]), .ZN(n945) );
  BUF_X1 U257 ( .A(n985), .Z(n2044) );
  BUF_X1 U258 ( .A(n985), .Z(n2045) );
  BUF_X1 U259 ( .A(n985), .Z(n2046) );
  INV_X1 U260 ( .A(n932), .ZN(n2169) );
  BUF_X1 U261 ( .A(n983), .Z(n2087) );
  BUF_X1 U262 ( .A(n983), .Z(n2086) );
  NAND2_X1 U263 ( .A1(n968), .A2(n969), .ZN(n595) );
  NAND2_X1 U264 ( .A1(n959), .A2(n968), .ZN(n617) );
  NAND2_X1 U265 ( .A1(n968), .A2(n949), .ZN(n601) );
  AND2_X1 U266 ( .A1(n968), .A2(n945), .ZN(n604) );
  NOR2_X2 U267 ( .A1(n933), .A2(n981), .ZN(n620) );
  AND2_X1 U268 ( .A1(n968), .A2(n957), .ZN(n616) );
  NAND2_X1 U269 ( .A1(n968), .A2(n950), .ZN(n613) );
  NOR2_X1 U270 ( .A1(n2145), .A2(n2149), .ZN(n946) );
  NOR3_X1 U271 ( .A1(n2147), .A2(n2146), .A3(n2148), .ZN(n969) );
  NOR2_X1 U272 ( .A1(n2147), .A2(addr_y[1]), .ZN(n957) );
  NAND2_X1 U273 ( .A1(n968), .A2(n948), .ZN(n965) );
  NOR2_X1 U274 ( .A1(n933), .A2(n2163), .ZN(n979) );
  INV_X1 U275 ( .A(n981), .ZN(n2163) );
  NOR2_X1 U276 ( .A1(n2148), .A2(addr_y[2]), .ZN(n970) );
  AND2_X1 U277 ( .A1(n970), .A2(n2146), .ZN(n948) );
  NAND2_X1 U278 ( .A1(n1018), .A2(n2170), .ZN(n932) );
  NAND2_X1 U279 ( .A1(n958), .A2(n968), .ZN(n976) );
  AND2_X1 U280 ( .A1(n978), .A2(n2147), .ZN(n958) );
  NOR2_X1 U281 ( .A1(n2146), .A2(addr_y[3]), .ZN(n978) );
  AND2_X1 U282 ( .A1(n983), .A2(n2170), .ZN(n985) );
  AND2_X1 U283 ( .A1(n1002), .A2(n932), .ZN(n983) );
  AND2_X1 U284 ( .A1(n932), .A2(n933), .ZN(n577) );
  NOR2_X1 U285 ( .A1(n2145), .A2(addr_y[4]), .ZN(n968) );
  BUF_X4 U286 ( .A(data_out_x[7]), .Z(n2143) );
  BUF_X4 U287 ( .A(data_out_x[7]), .Z(n2142) );
  AOI221_X1 U288 ( .B1(f29[0]), .B2(n582), .C1(f28[0]), .C2(n583), .A(n938), 
        .ZN(n937) );
  OAI22_X1 U289 ( .A1(n585), .A2(n512), .B1(n586), .B2(n464), .ZN(n938) );
  AOI221_X1 U290 ( .B1(f29[1]), .B2(n582), .C1(f28[1]), .C2(n583), .A(n914), 
        .ZN(n913) );
  OAI22_X1 U291 ( .A1(n585), .A2(n511), .B1(n586), .B2(n463), .ZN(n914) );
  AOI221_X1 U292 ( .B1(f29[2]), .B2(n582), .C1(f28[2]), .C2(n583), .A(n892), 
        .ZN(n891) );
  OAI22_X1 U293 ( .A1(n585), .A2(n510), .B1(n586), .B2(n462), .ZN(n892) );
  AOI221_X1 U294 ( .B1(f29[3]), .B2(n582), .C1(f28[3]), .C2(n583), .A(n870), 
        .ZN(n869) );
  OAI22_X1 U295 ( .A1(n585), .A2(n509), .B1(n586), .B2(n461), .ZN(n870) );
  AOI221_X1 U296 ( .B1(f29[4]), .B2(n582), .C1(f28[4]), .C2(n583), .A(n848), 
        .ZN(n847) );
  OAI22_X1 U297 ( .A1(n585), .A2(n508), .B1(n586), .B2(n460), .ZN(n848) );
  AOI221_X1 U298 ( .B1(f29[5]), .B2(n582), .C1(f28[5]), .C2(n583), .A(n826), 
        .ZN(n825) );
  OAI22_X1 U299 ( .A1(n585), .A2(n507), .B1(n586), .B2(n459), .ZN(n826) );
  AOI221_X1 U300 ( .B1(f29[6]), .B2(n582), .C1(f28[6]), .C2(n583), .A(n804), 
        .ZN(n803) );
  OAI22_X1 U301 ( .A1(n585), .A2(n506), .B1(n586), .B2(n458), .ZN(n804) );
  AOI221_X1 U302 ( .B1(f29[7]), .B2(n582), .C1(f28[7]), .C2(n583), .A(n782), 
        .ZN(n781) );
  OAI22_X1 U303 ( .A1(n585), .A2(n505), .B1(n586), .B2(n457), .ZN(n782) );
  AOI221_X1 U304 ( .B1(f29[8]), .B2(n582), .C1(f28[8]), .C2(n583), .A(n760), 
        .ZN(n759) );
  OAI22_X1 U305 ( .A1(n585), .A2(n504), .B1(n586), .B2(n456), .ZN(n760) );
  AOI221_X1 U306 ( .B1(f29[9]), .B2(n582), .C1(f28[9]), .C2(n583), .A(n738), 
        .ZN(n737) );
  OAI22_X1 U307 ( .A1(n585), .A2(n503), .B1(n586), .B2(n455), .ZN(n738) );
  AOI221_X1 U308 ( .B1(f29[10]), .B2(n582), .C1(f28[10]), .C2(n583), .A(n716), 
        .ZN(n715) );
  OAI22_X1 U309 ( .A1(n585), .A2(n502), .B1(n586), .B2(n454), .ZN(n716) );
  AOI221_X1 U310 ( .B1(f29[11]), .B2(n582), .C1(f28[11]), .C2(n583), .A(n694), 
        .ZN(n693) );
  OAI22_X1 U311 ( .A1(n585), .A2(n501), .B1(n586), .B2(n453), .ZN(n694) );
  AOI221_X1 U312 ( .B1(f29[12]), .B2(n582), .C1(f28[12]), .C2(n583), .A(n672), 
        .ZN(n671) );
  OAI22_X1 U313 ( .A1(n585), .A2(n500), .B1(n586), .B2(n452), .ZN(n672) );
  AOI221_X1 U314 ( .B1(f29[13]), .B2(n582), .C1(f28[13]), .C2(n583), .A(n650), 
        .ZN(n649) );
  OAI22_X1 U315 ( .A1(n585), .A2(n499), .B1(n586), .B2(n451), .ZN(n650) );
  AOI221_X1 U316 ( .B1(f29[14]), .B2(n582), .C1(f28[14]), .C2(n583), .A(n628), 
        .ZN(n627) );
  OAI22_X1 U317 ( .A1(n585), .A2(n498), .B1(n586), .B2(n450), .ZN(n628) );
  AOI221_X1 U318 ( .B1(f29[15]), .B2(n582), .C1(f28[15]), .C2(n583), .A(n584), 
        .ZN(n581) );
  OAI22_X1 U319 ( .A1(n585), .A2(n497), .B1(n586), .B2(n449), .ZN(n584) );
  AOI22_X1 U320 ( .A1(f5[0]), .A2(n2154), .B1(f4[0]), .B2(n2153), .ZN(n974) );
  AOI22_X1 U321 ( .A1(f5[1]), .A2(n2154), .B1(f4[1]), .B2(n2153), .ZN(n928) );
  AOI22_X1 U322 ( .A1(f5[2]), .A2(n2154), .B1(f4[2]), .B2(n2153), .ZN(n906) );
  AOI22_X1 U323 ( .A1(f5[3]), .A2(n2154), .B1(f4[3]), .B2(n2153), .ZN(n884) );
  AOI22_X1 U324 ( .A1(f5[4]), .A2(n2154), .B1(f4[4]), .B2(n2153), .ZN(n862) );
  AOI22_X1 U325 ( .A1(f5[5]), .A2(n2154), .B1(f4[5]), .B2(n2153), .ZN(n840) );
  AOI22_X1 U326 ( .A1(f5[6]), .A2(n2154), .B1(f4[6]), .B2(n2153), .ZN(n818) );
  AOI22_X1 U327 ( .A1(f5[7]), .A2(n2154), .B1(f4[7]), .B2(n2153), .ZN(n796) );
  AOI22_X1 U328 ( .A1(f5[8]), .A2(n2154), .B1(f4[8]), .B2(n2153), .ZN(n774) );
  AOI22_X1 U329 ( .A1(f5[9]), .A2(n2154), .B1(f4[9]), .B2(n2153), .ZN(n752) );
  AOI22_X1 U330 ( .A1(f5[10]), .A2(n2154), .B1(f4[10]), .B2(n2153), .ZN(n730)
         );
  AOI22_X1 U331 ( .A1(f5[11]), .A2(n2154), .B1(f4[11]), .B2(n2153), .ZN(n708)
         );
  AOI22_X1 U332 ( .A1(f5[12]), .A2(n2154), .B1(f4[12]), .B2(n2153), .ZN(n686)
         );
  AOI22_X1 U333 ( .A1(f5[13]), .A2(n2154), .B1(f4[13]), .B2(n2153), .ZN(n664)
         );
  AOI22_X1 U334 ( .A1(f5[14]), .A2(n2154), .B1(f4[14]), .B2(n2153), .ZN(n642)
         );
  AOI22_X1 U335 ( .A1(f5[15]), .A2(n2154), .B1(f4[15]), .B2(n2153), .ZN(n619)
         );
  AOI22_X1 U336 ( .A1(f19[0]), .A2(n2159), .B1(f18[0]), .B2(n2164), .ZN(n953)
         );
  AOI22_X1 U337 ( .A1(f19[1]), .A2(n2159), .B1(f18[1]), .B2(n2164), .ZN(n919)
         );
  AOI22_X1 U338 ( .A1(f19[2]), .A2(n2159), .B1(f18[2]), .B2(n2164), .ZN(n897)
         );
  AOI22_X1 U339 ( .A1(f19[3]), .A2(n2159), .B1(f18[3]), .B2(n2164), .ZN(n875)
         );
  AOI22_X1 U340 ( .A1(f19[4]), .A2(n2159), .B1(f18[4]), .B2(n2164), .ZN(n853)
         );
  AOI22_X1 U341 ( .A1(f19[5]), .A2(n2159), .B1(f18[5]), .B2(n2164), .ZN(n831)
         );
  AOI22_X1 U342 ( .A1(f19[6]), .A2(n2159), .B1(f18[6]), .B2(n2164), .ZN(n809)
         );
  AOI22_X1 U343 ( .A1(f19[7]), .A2(n2159), .B1(f18[7]), .B2(n2164), .ZN(n787)
         );
  AOI22_X1 U344 ( .A1(f19[8]), .A2(n2159), .B1(f18[8]), .B2(n2164), .ZN(n765)
         );
  AOI22_X1 U345 ( .A1(f19[9]), .A2(n2159), .B1(f18[9]), .B2(n2164), .ZN(n743)
         );
  AOI22_X1 U346 ( .A1(f19[10]), .A2(n2159), .B1(f18[10]), .B2(n2164), .ZN(n721) );
  AOI22_X1 U347 ( .A1(f19[11]), .A2(n2159), .B1(f18[11]), .B2(n2164), .ZN(n699) );
  AOI22_X1 U348 ( .A1(f19[12]), .A2(n2159), .B1(f18[12]), .B2(n2164), .ZN(n677) );
  AOI22_X1 U349 ( .A1(f19[13]), .A2(n2159), .B1(f18[13]), .B2(n2164), .ZN(n655) );
  AOI22_X1 U350 ( .A1(f19[14]), .A2(n2159), .B1(f18[14]), .B2(n2164), .ZN(n633) );
  AOI22_X1 U351 ( .A1(f19[15]), .A2(n2159), .B1(f18[15]), .B2(n2164), .ZN(n598) );
  AOI22_X1 U352 ( .A1(f12[0]), .A2(n2151), .B1(f11[0]), .B2(n2156), .ZN(n964)
         );
  AOI22_X1 U353 ( .A1(f12[1]), .A2(n2151), .B1(f11[1]), .B2(n2156), .ZN(n924)
         );
  AOI22_X1 U354 ( .A1(f12[2]), .A2(n2151), .B1(f11[2]), .B2(n2156), .ZN(n902)
         );
  AOI22_X1 U355 ( .A1(f12[3]), .A2(n2151), .B1(f11[3]), .B2(n2156), .ZN(n880)
         );
  AOI22_X1 U356 ( .A1(f12[4]), .A2(n2151), .B1(f11[4]), .B2(n2156), .ZN(n858)
         );
  AOI22_X1 U357 ( .A1(f12[5]), .A2(n2151), .B1(f11[5]), .B2(n2156), .ZN(n836)
         );
  AOI22_X1 U358 ( .A1(f12[6]), .A2(n2151), .B1(f11[6]), .B2(n2156), .ZN(n814)
         );
  AOI22_X1 U359 ( .A1(f12[7]), .A2(n2151), .B1(f11[7]), .B2(n2156), .ZN(n792)
         );
  AOI22_X1 U360 ( .A1(f12[8]), .A2(n2151), .B1(f11[8]), .B2(n2156), .ZN(n770)
         );
  AOI22_X1 U361 ( .A1(f12[9]), .A2(n2151), .B1(f11[9]), .B2(n2156), .ZN(n748)
         );
  AOI22_X1 U362 ( .A1(f12[10]), .A2(n2151), .B1(f11[10]), .B2(n2156), .ZN(n726) );
  AOI22_X1 U363 ( .A1(f12[11]), .A2(n2151), .B1(f11[11]), .B2(n2156), .ZN(n704) );
  AOI22_X1 U364 ( .A1(f12[12]), .A2(n2151), .B1(f11[12]), .B2(n2156), .ZN(n682) );
  AOI22_X1 U365 ( .A1(f12[13]), .A2(n2151), .B1(f11[13]), .B2(n2156), .ZN(n660) );
  AOI22_X1 U366 ( .A1(f12[14]), .A2(n2151), .B1(f11[14]), .B2(n2156), .ZN(n638) );
  AOI22_X1 U367 ( .A1(f12[15]), .A2(n2151), .B1(f11[15]), .B2(n2156), .ZN(n609) );
  AOI22_X1 U368 ( .A1(f26[0]), .A2(n2166), .B1(f25[0]), .B2(n2161), .ZN(n936)
         );
  AOI22_X1 U369 ( .A1(f26[1]), .A2(n2166), .B1(f25[1]), .B2(n2161), .ZN(n912)
         );
  AOI22_X1 U370 ( .A1(f26[2]), .A2(n2166), .B1(f25[2]), .B2(n2161), .ZN(n890)
         );
  AOI22_X1 U371 ( .A1(f26[3]), .A2(n2166), .B1(f25[3]), .B2(n2161), .ZN(n868)
         );
  AOI22_X1 U372 ( .A1(f26[4]), .A2(n2166), .B1(f25[4]), .B2(n2161), .ZN(n846)
         );
  AOI22_X1 U373 ( .A1(f26[5]), .A2(n2166), .B1(f25[5]), .B2(n2161), .ZN(n824)
         );
  AOI22_X1 U374 ( .A1(f26[6]), .A2(n2166), .B1(f25[6]), .B2(n2161), .ZN(n802)
         );
  AOI22_X1 U375 ( .A1(f26[7]), .A2(n2166), .B1(f25[7]), .B2(n2161), .ZN(n780)
         );
  AOI22_X1 U376 ( .A1(f26[8]), .A2(n2166), .B1(f25[8]), .B2(n2161), .ZN(n758)
         );
  AOI22_X1 U377 ( .A1(f26[9]), .A2(n2166), .B1(f25[9]), .B2(n2161), .ZN(n736)
         );
  AOI22_X1 U378 ( .A1(f26[10]), .A2(n2166), .B1(f25[10]), .B2(n2161), .ZN(n714) );
  AOI22_X1 U379 ( .A1(f26[11]), .A2(n2166), .B1(f25[11]), .B2(n2161), .ZN(n692) );
  AOI22_X1 U380 ( .A1(f26[12]), .A2(n2166), .B1(f25[12]), .B2(n2161), .ZN(n670) );
  AOI22_X1 U381 ( .A1(f26[13]), .A2(n2166), .B1(f25[13]), .B2(n2161), .ZN(n648) );
  AOI22_X1 U382 ( .A1(f26[14]), .A2(n2166), .B1(f25[14]), .B2(n2161), .ZN(n626) );
  AOI22_X1 U383 ( .A1(f26[15]), .A2(n2166), .B1(f25[15]), .B2(n2161), .ZN(n580) );
  OAI211_X1 U384 ( .C1(n572), .C2(n528), .A(n929), .B(n930), .ZN(n1514) );
  AOI22_X1 U385 ( .A1(f1[0]), .A2(n2169), .B1(f32[0]), .B2(n620), .ZN(n929) );
  AOI22_X1 U386 ( .A1(n575), .A2(n931), .B1(f[0]), .B2(n577), .ZN(n930) );
  NAND4_X1 U387 ( .A1(n934), .A2(n935), .A3(n936), .A4(n937), .ZN(n931) );
  OAI211_X1 U388 ( .C1(n572), .C2(n527), .A(n907), .B(n908), .ZN(n1513) );
  AOI22_X1 U389 ( .A1(f1[1]), .A2(n2169), .B1(f32[1]), .B2(n620), .ZN(n907) );
  AOI22_X1 U390 ( .A1(n575), .A2(n909), .B1(f[1]), .B2(n577), .ZN(n908) );
  NAND4_X1 U391 ( .A1(n910), .A2(n911), .A3(n912), .A4(n913), .ZN(n909) );
  OAI211_X1 U392 ( .C1(n572), .C2(n526), .A(n885), .B(n886), .ZN(n1512) );
  AOI22_X1 U393 ( .A1(f1[2]), .A2(n2169), .B1(f32[2]), .B2(n620), .ZN(n885) );
  AOI22_X1 U394 ( .A1(n575), .A2(n887), .B1(f[2]), .B2(n577), .ZN(n886) );
  NAND4_X1 U395 ( .A1(n888), .A2(n889), .A3(n890), .A4(n891), .ZN(n887) );
  OAI211_X1 U396 ( .C1(n572), .C2(n525), .A(n863), .B(n864), .ZN(n1511) );
  AOI22_X1 U397 ( .A1(f1[3]), .A2(n2169), .B1(f32[3]), .B2(n620), .ZN(n863) );
  AOI22_X1 U398 ( .A1(n575), .A2(n865), .B1(f[3]), .B2(n577), .ZN(n864) );
  NAND4_X1 U399 ( .A1(n866), .A2(n867), .A3(n868), .A4(n869), .ZN(n865) );
  OAI211_X1 U400 ( .C1(n572), .C2(n524), .A(n841), .B(n842), .ZN(n1510) );
  AOI22_X1 U401 ( .A1(f1[4]), .A2(n2169), .B1(f32[4]), .B2(n620), .ZN(n841) );
  AOI22_X1 U402 ( .A1(n575), .A2(n843), .B1(f[4]), .B2(n577), .ZN(n842) );
  NAND4_X1 U403 ( .A1(n844), .A2(n845), .A3(n846), .A4(n847), .ZN(n843) );
  OAI211_X1 U404 ( .C1(n572), .C2(n523), .A(n819), .B(n820), .ZN(n1509) );
  AOI22_X1 U405 ( .A1(f1[5]), .A2(n2169), .B1(f32[5]), .B2(n620), .ZN(n819) );
  AOI22_X1 U406 ( .A1(n575), .A2(n821), .B1(f[5]), .B2(n577), .ZN(n820) );
  NAND4_X1 U407 ( .A1(n822), .A2(n823), .A3(n824), .A4(n825), .ZN(n821) );
  OAI211_X1 U408 ( .C1(n572), .C2(n522), .A(n797), .B(n798), .ZN(n1508) );
  AOI22_X1 U409 ( .A1(f1[6]), .A2(n2169), .B1(f32[6]), .B2(n620), .ZN(n797) );
  AOI22_X1 U410 ( .A1(n575), .A2(n799), .B1(f[6]), .B2(n577), .ZN(n798) );
  NAND4_X1 U411 ( .A1(n800), .A2(n801), .A3(n802), .A4(n803), .ZN(n799) );
  OAI211_X1 U412 ( .C1(n572), .C2(n521), .A(n775), .B(n776), .ZN(n1507) );
  AOI22_X1 U413 ( .A1(f1[7]), .A2(n2169), .B1(f32[7]), .B2(n620), .ZN(n775) );
  AOI22_X1 U414 ( .A1(n575), .A2(n777), .B1(f[7]), .B2(n577), .ZN(n776) );
  NAND4_X1 U415 ( .A1(n778), .A2(n779), .A3(n780), .A4(n781), .ZN(n777) );
  OAI211_X1 U416 ( .C1(n572), .C2(n520), .A(n753), .B(n754), .ZN(n1506) );
  AOI22_X1 U417 ( .A1(f1[8]), .A2(n2169), .B1(f32[8]), .B2(n620), .ZN(n753) );
  AOI22_X1 U418 ( .A1(n575), .A2(n755), .B1(f[8]), .B2(n577), .ZN(n754) );
  NAND4_X1 U419 ( .A1(n756), .A2(n757), .A3(n758), .A4(n759), .ZN(n755) );
  OAI211_X1 U420 ( .C1(n572), .C2(n519), .A(n731), .B(n732), .ZN(n1505) );
  AOI22_X1 U421 ( .A1(f1[9]), .A2(n2169), .B1(f32[9]), .B2(n620), .ZN(n731) );
  AOI22_X1 U422 ( .A1(n575), .A2(n733), .B1(f[9]), .B2(n577), .ZN(n732) );
  NAND4_X1 U423 ( .A1(n734), .A2(n735), .A3(n736), .A4(n737), .ZN(n733) );
  OAI211_X1 U424 ( .C1(n572), .C2(n518), .A(n709), .B(n710), .ZN(n1504) );
  AOI22_X1 U425 ( .A1(f1[10]), .A2(n2169), .B1(f32[10]), .B2(n620), .ZN(n709)
         );
  AOI22_X1 U426 ( .A1(n575), .A2(n711), .B1(f[10]), .B2(n577), .ZN(n710) );
  NAND4_X1 U427 ( .A1(n712), .A2(n713), .A3(n714), .A4(n715), .ZN(n711) );
  OAI211_X1 U428 ( .C1(n572), .C2(n517), .A(n687), .B(n688), .ZN(n1503) );
  AOI22_X1 U429 ( .A1(f1[11]), .A2(n2169), .B1(f32[11]), .B2(n620), .ZN(n687)
         );
  AOI22_X1 U430 ( .A1(n575), .A2(n689), .B1(f[11]), .B2(n577), .ZN(n688) );
  NAND4_X1 U431 ( .A1(n690), .A2(n691), .A3(n692), .A4(n693), .ZN(n689) );
  OAI211_X1 U432 ( .C1(n572), .C2(n516), .A(n665), .B(n666), .ZN(n1502) );
  AOI22_X1 U433 ( .A1(f1[12]), .A2(n2169), .B1(f32[12]), .B2(n620), .ZN(n665)
         );
  AOI22_X1 U434 ( .A1(n575), .A2(n667), .B1(f[12]), .B2(n577), .ZN(n666) );
  NAND4_X1 U435 ( .A1(n668), .A2(n669), .A3(n670), .A4(n671), .ZN(n667) );
  OAI211_X1 U436 ( .C1(n572), .C2(n515), .A(n643), .B(n644), .ZN(n1501) );
  AOI22_X1 U437 ( .A1(f1[13]), .A2(n2169), .B1(f32[13]), .B2(n620), .ZN(n643)
         );
  AOI22_X1 U438 ( .A1(n575), .A2(n645), .B1(f[13]), .B2(n577), .ZN(n644) );
  NAND4_X1 U439 ( .A1(n646), .A2(n647), .A3(n648), .A4(n649), .ZN(n645) );
  OAI211_X1 U440 ( .C1(n572), .C2(n514), .A(n621), .B(n622), .ZN(n1500) );
  AOI22_X1 U441 ( .A1(f1[14]), .A2(n2169), .B1(f32[14]), .B2(n620), .ZN(n621)
         );
  AOI22_X1 U442 ( .A1(n575), .A2(n623), .B1(f[14]), .B2(n577), .ZN(n622) );
  NAND4_X1 U443 ( .A1(n624), .A2(n625), .A3(n626), .A4(n627), .ZN(n623) );
  OAI211_X1 U444 ( .C1(n572), .C2(n513), .A(n573), .B(n574), .ZN(n1499) );
  AOI22_X1 U445 ( .A1(f1[15]), .A2(n2169), .B1(f32[15]), .B2(n620), .ZN(n573)
         );
  AOI22_X1 U446 ( .A1(n575), .A2(n576), .B1(f[15]), .B2(n577), .ZN(n574) );
  NAND4_X1 U447 ( .A1(n578), .A2(n579), .A3(n580), .A4(n581), .ZN(n576) );
  OAI21_X1 U448 ( .B1(n2090), .B2(n518), .A(n1012), .ZN(n1541) );
  NAND2_X1 U449 ( .A1(add_r31[10]), .A2(n2078), .ZN(n1012) );
  OAI21_X1 U450 ( .B1(n2090), .B2(n517), .A(n1013), .ZN(n1542) );
  NAND2_X1 U451 ( .A1(add_r31[11]), .A2(n2078), .ZN(n1013) );
  OAI21_X1 U452 ( .B1(n2118), .B2(n134), .A(n1397), .ZN(n1925) );
  NAND2_X1 U453 ( .A1(add_r7[10]), .A2(n2055), .ZN(n1397) );
  OAI21_X1 U454 ( .B1(n2118), .B2(n133), .A(n1398), .ZN(n1926) );
  NAND2_X1 U455 ( .A1(add_r7[11]), .A2(n2055), .ZN(n1398) );
  OAI21_X1 U456 ( .B1(n2118), .B2(n130), .A(n1401), .ZN(n1929) );
  NAND2_X1 U457 ( .A1(add_r7[14]), .A2(n2055), .ZN(n1401) );
  NAND2_X1 U458 ( .A1(add_r31[14]), .A2(n2078), .ZN(n1016) );
  OAI21_X1 U459 ( .B1(n2120), .B2(n194), .A(n1337), .ZN(n1865) );
  NAND2_X1 U460 ( .A1(add_r11[14]), .A2(n2060), .ZN(n1337) );
  OAI21_X1 U461 ( .B1(n2118), .B2(n131), .A(n1400), .ZN(n1928) );
  NAND2_X1 U462 ( .A1(add_r7[13]), .A2(n2055), .ZN(n1400) );
  OAI21_X1 U463 ( .B1(n2090), .B2(n515), .A(n1015), .ZN(n1544) );
  NAND2_X1 U464 ( .A1(add_r31[13]), .A2(n2078), .ZN(n1015) );
  OAI21_X1 U465 ( .B1(n2120), .B2(n195), .A(n1336), .ZN(n1864) );
  NAND2_X1 U466 ( .A1(add_r11[13]), .A2(n2060), .ZN(n1336) );
  OAI21_X1 U467 ( .B1(n2118), .B2(n132), .A(n1399), .ZN(n1927) );
  NAND2_X1 U468 ( .A1(add_r7[12]), .A2(n2055), .ZN(n1399) );
  OAI21_X1 U469 ( .B1(n2090), .B2(n516), .A(n1014), .ZN(n1543) );
  NAND2_X1 U470 ( .A1(add_r31[12]), .A2(n2078), .ZN(n1014) );
  OAI21_X1 U471 ( .B1(n2110), .B2(n196), .A(n1335), .ZN(n1863) );
  NAND2_X1 U472 ( .A1(add_r11[12]), .A2(n2060), .ZN(n1335) );
  OAI21_X1 U473 ( .B1(n2090), .B2(n520), .A(n1010), .ZN(n1539) );
  NAND2_X1 U474 ( .A1(add_r31[8]), .A2(n2078), .ZN(n1010) );
  OAI21_X1 U475 ( .B1(n2090), .B2(n519), .A(n1011), .ZN(n1540) );
  NAND2_X1 U476 ( .A1(add_r31[9]), .A2(n2078), .ZN(n1011) );
  OAI21_X1 U477 ( .B1(n2090), .B2(n512), .A(n1019), .ZN(n1547) );
  NAND2_X1 U478 ( .A1(add_r30[0]), .A2(n2077), .ZN(n1019) );
  OAI21_X1 U479 ( .B1(n2090), .B2(n511), .A(n1020), .ZN(n1548) );
  NAND2_X1 U480 ( .A1(add_r30[1]), .A2(n2077), .ZN(n1020) );
  OAI21_X1 U481 ( .B1(n2090), .B2(n510), .A(n1021), .ZN(n1549) );
  NAND2_X1 U482 ( .A1(add_r30[2]), .A2(n2077), .ZN(n1021) );
  OAI21_X1 U483 ( .B1(n2090), .B2(n509), .A(n1022), .ZN(n1550) );
  NAND2_X1 U484 ( .A1(add_r30[3]), .A2(n2077), .ZN(n1022) );
  OAI21_X1 U485 ( .B1(n2120), .B2(n192), .A(n1339), .ZN(n1867) );
  NAND2_X1 U486 ( .A1(add_r10[0]), .A2(n2060), .ZN(n1339) );
  OAI21_X1 U487 ( .B1(n2120), .B2(n191), .A(n1340), .ZN(n1868) );
  NAND2_X1 U488 ( .A1(add_r10[1]), .A2(n2060), .ZN(n1340) );
  OAI21_X1 U489 ( .B1(n2110), .B2(n190), .A(n1341), .ZN(n1869) );
  NAND2_X1 U490 ( .A1(add_r10[2]), .A2(n2060), .ZN(n1341) );
  OAI21_X1 U491 ( .B1(n2120), .B2(n189), .A(n1342), .ZN(n1870) );
  NAND2_X1 U492 ( .A1(add_r10[3]), .A2(n2060), .ZN(n1342) );
  OAI21_X1 U493 ( .B1(n2110), .B2(n188), .A(n1343), .ZN(n1871) );
  NAND2_X1 U494 ( .A1(add_r10[4]), .A2(n2059), .ZN(n1343) );
  OAI21_X1 U495 ( .B1(n2120), .B2(n187), .A(n1344), .ZN(n1872) );
  NAND2_X1 U496 ( .A1(add_r10[5]), .A2(n2059), .ZN(n1344) );
  OAI21_X1 U497 ( .B1(n2110), .B2(n186), .A(n1345), .ZN(n1873) );
  NAND2_X1 U498 ( .A1(add_r10[6]), .A2(n2059), .ZN(n1345) );
  OAI21_X1 U499 ( .B1(n2120), .B2(n185), .A(n1346), .ZN(n1874) );
  NAND2_X1 U500 ( .A1(add_r10[7]), .A2(n2059), .ZN(n1346) );
  OAI21_X1 U501 ( .B1(n2118), .B2(n136), .A(n1395), .ZN(n1923) );
  NAND2_X1 U502 ( .A1(add_r7[8]), .A2(n2055), .ZN(n1395) );
  OAI21_X1 U503 ( .B1(n2118), .B2(n135), .A(n1396), .ZN(n1924) );
  NAND2_X1 U504 ( .A1(add_r7[9]), .A2(n2055), .ZN(n1396) );
  OAI21_X1 U505 ( .B1(n2118), .B2(n128), .A(n1403), .ZN(n1931) );
  NAND2_X1 U506 ( .A1(add_r6[0]), .A2(n2054), .ZN(n1403) );
  OAI21_X1 U507 ( .B1(n2118), .B2(n127), .A(n1404), .ZN(n1932) );
  NAND2_X1 U508 ( .A1(add_r6[1]), .A2(n2054), .ZN(n1404) );
  OAI21_X1 U509 ( .B1(n2118), .B2(n126), .A(n1405), .ZN(n1933) );
  NAND2_X1 U510 ( .A1(add_r6[2]), .A2(n2054), .ZN(n1405) );
  OAI21_X1 U511 ( .B1(n2118), .B2(n125), .A(n1406), .ZN(n1934) );
  NAND2_X1 U512 ( .A1(add_r6[3]), .A2(n2054), .ZN(n1406) );
  NOR2_X1 U513 ( .A1(n2171), .A2(clc1), .ZN(n1018) );
  INV_X1 U514 ( .A(clc), .ZN(n2171) );
  OAI21_X1 U515 ( .B1(n942), .B2(n943), .A(n589), .ZN(n934) );
  OAI221_X1 U516 ( .B1(n590), .B2(n384), .C1(n591), .C2(n368), .A(n951), .ZN(
        n943) );
  OAI221_X1 U517 ( .B1(n595), .B2(n304), .C1(n952), .C2(n597), .A(n953), .ZN(
        n942) );
  AOI22_X1 U518 ( .A1(f20[0]), .A2(n593), .B1(f23[0]), .B2(n594), .ZN(n951) );
  OAI21_X1 U519 ( .B1(n915), .B2(n916), .A(n589), .ZN(n910) );
  OAI221_X1 U520 ( .B1(n590), .B2(n383), .C1(n591), .C2(n367), .A(n917), .ZN(
        n916) );
  OAI221_X1 U521 ( .B1(n595), .B2(n303), .C1(n918), .C2(n597), .A(n919), .ZN(
        n915) );
  AOI22_X1 U522 ( .A1(f20[1]), .A2(n593), .B1(f23[1]), .B2(n594), .ZN(n917) );
  OAI21_X1 U523 ( .B1(n893), .B2(n894), .A(n589), .ZN(n888) );
  OAI221_X1 U524 ( .B1(n590), .B2(n382), .C1(n591), .C2(n366), .A(n895), .ZN(
        n894) );
  OAI221_X1 U525 ( .B1(n595), .B2(n302), .C1(n896), .C2(n597), .A(n897), .ZN(
        n893) );
  AOI22_X1 U526 ( .A1(f20[2]), .A2(n593), .B1(f23[2]), .B2(n594), .ZN(n895) );
  OAI21_X1 U527 ( .B1(n871), .B2(n872), .A(n589), .ZN(n866) );
  OAI221_X1 U528 ( .B1(n590), .B2(n381), .C1(n591), .C2(n365), .A(n873), .ZN(
        n872) );
  OAI221_X1 U529 ( .B1(n595), .B2(n301), .C1(n874), .C2(n597), .A(n875), .ZN(
        n871) );
  AOI22_X1 U530 ( .A1(f20[3]), .A2(n593), .B1(f23[3]), .B2(n594), .ZN(n873) );
  OAI21_X1 U531 ( .B1(n849), .B2(n850), .A(n589), .ZN(n844) );
  OAI221_X1 U532 ( .B1(n590), .B2(n380), .C1(n591), .C2(n364), .A(n851), .ZN(
        n850) );
  OAI221_X1 U533 ( .B1(n595), .B2(n300), .C1(n852), .C2(n597), .A(n853), .ZN(
        n849) );
  AOI22_X1 U534 ( .A1(f20[4]), .A2(n593), .B1(f23[4]), .B2(n594), .ZN(n851) );
  OAI21_X1 U535 ( .B1(n827), .B2(n828), .A(n589), .ZN(n822) );
  OAI221_X1 U536 ( .B1(n590), .B2(n379), .C1(n591), .C2(n363), .A(n829), .ZN(
        n828) );
  OAI221_X1 U537 ( .B1(n595), .B2(n299), .C1(n830), .C2(n597), .A(n831), .ZN(
        n827) );
  AOI22_X1 U538 ( .A1(f20[5]), .A2(n593), .B1(f23[5]), .B2(n594), .ZN(n829) );
  OAI21_X1 U539 ( .B1(n805), .B2(n806), .A(n589), .ZN(n800) );
  OAI221_X1 U540 ( .B1(n590), .B2(n378), .C1(n591), .C2(n362), .A(n807), .ZN(
        n806) );
  OAI221_X1 U541 ( .B1(n595), .B2(n298), .C1(n808), .C2(n597), .A(n809), .ZN(
        n805) );
  AOI22_X1 U542 ( .A1(f20[6]), .A2(n593), .B1(f23[6]), .B2(n594), .ZN(n807) );
  OAI21_X1 U543 ( .B1(n783), .B2(n784), .A(n589), .ZN(n778) );
  OAI221_X1 U544 ( .B1(n590), .B2(n377), .C1(n591), .C2(n361), .A(n785), .ZN(
        n784) );
  OAI221_X1 U545 ( .B1(n595), .B2(n297), .C1(n786), .C2(n597), .A(n787), .ZN(
        n783) );
  AOI22_X1 U546 ( .A1(f20[7]), .A2(n593), .B1(f23[7]), .B2(n594), .ZN(n785) );
  OAI21_X1 U547 ( .B1(n761), .B2(n762), .A(n589), .ZN(n756) );
  OAI221_X1 U548 ( .B1(n590), .B2(n376), .C1(n591), .C2(n360), .A(n763), .ZN(
        n762) );
  OAI221_X1 U549 ( .B1(n595), .B2(n296), .C1(n764), .C2(n597), .A(n765), .ZN(
        n761) );
  AOI22_X1 U550 ( .A1(f20[8]), .A2(n593), .B1(f23[8]), .B2(n594), .ZN(n763) );
  OAI21_X1 U551 ( .B1(n739), .B2(n740), .A(n589), .ZN(n734) );
  OAI221_X1 U552 ( .B1(n590), .B2(n375), .C1(n591), .C2(n359), .A(n741), .ZN(
        n740) );
  OAI221_X1 U553 ( .B1(n595), .B2(n295), .C1(n742), .C2(n597), .A(n743), .ZN(
        n739) );
  AOI22_X1 U554 ( .A1(f20[9]), .A2(n593), .B1(f23[9]), .B2(n594), .ZN(n741) );
  OAI21_X1 U555 ( .B1(n717), .B2(n718), .A(n589), .ZN(n712) );
  OAI221_X1 U556 ( .B1(n590), .B2(n374), .C1(n591), .C2(n358), .A(n719), .ZN(
        n718) );
  OAI221_X1 U557 ( .B1(n595), .B2(n294), .C1(n720), .C2(n597), .A(n721), .ZN(
        n717) );
  AOI22_X1 U558 ( .A1(f20[10]), .A2(n593), .B1(f23[10]), .B2(n594), .ZN(n719)
         );
  OAI21_X1 U559 ( .B1(n695), .B2(n696), .A(n589), .ZN(n690) );
  OAI221_X1 U560 ( .B1(n590), .B2(n373), .C1(n591), .C2(n357), .A(n697), .ZN(
        n696) );
  OAI221_X1 U561 ( .B1(n595), .B2(n293), .C1(n698), .C2(n597), .A(n699), .ZN(
        n695) );
  AOI22_X1 U562 ( .A1(f20[11]), .A2(n593), .B1(f23[11]), .B2(n594), .ZN(n697)
         );
  OAI21_X1 U563 ( .B1(n673), .B2(n674), .A(n589), .ZN(n668) );
  OAI221_X1 U564 ( .B1(n590), .B2(n372), .C1(n591), .C2(n356), .A(n675), .ZN(
        n674) );
  OAI221_X1 U565 ( .B1(n595), .B2(n292), .C1(n676), .C2(n597), .A(n677), .ZN(
        n673) );
  AOI22_X1 U566 ( .A1(f20[12]), .A2(n593), .B1(f23[12]), .B2(n594), .ZN(n675)
         );
  OAI21_X1 U567 ( .B1(n651), .B2(n652), .A(n589), .ZN(n646) );
  OAI221_X1 U568 ( .B1(n590), .B2(n371), .C1(n591), .C2(n355), .A(n653), .ZN(
        n652) );
  OAI221_X1 U569 ( .B1(n595), .B2(n291), .C1(n654), .C2(n597), .A(n655), .ZN(
        n651) );
  AOI22_X1 U570 ( .A1(f20[13]), .A2(n593), .B1(f23[13]), .B2(n594), .ZN(n653)
         );
  OAI21_X1 U571 ( .B1(n629), .B2(n630), .A(n589), .ZN(n624) );
  OAI221_X1 U572 ( .B1(n590), .B2(n370), .C1(n591), .C2(n354), .A(n631), .ZN(
        n630) );
  OAI221_X1 U573 ( .B1(n595), .B2(n290), .C1(n632), .C2(n597), .A(n633), .ZN(
        n629) );
  AOI22_X1 U574 ( .A1(f20[14]), .A2(n593), .B1(f23[14]), .B2(n594), .ZN(n631)
         );
  OAI21_X1 U575 ( .B1(n587), .B2(n588), .A(n589), .ZN(n578) );
  OAI221_X1 U576 ( .B1(n590), .B2(n369), .C1(n591), .C2(n353), .A(n592), .ZN(
        n588) );
  OAI221_X1 U577 ( .B1(n595), .B2(n289), .C1(n596), .C2(n597), .A(n598), .ZN(
        n587) );
  AOI22_X1 U578 ( .A1(f20[15]), .A2(n593), .B1(f23[15]), .B2(n594), .ZN(n592)
         );
  NOR2_X1 U579 ( .A1(n960), .A2(n961), .ZN(n952) );
  OAI221_X1 U580 ( .B1(n601), .B2(n272), .C1(n602), .C2(n256), .A(n962), .ZN(
        n961) );
  OAI221_X1 U581 ( .B1(n606), .B2(n192), .C1(n963), .C2(n608), .A(n964), .ZN(
        n960) );
  AOI22_X1 U582 ( .A1(f13[0]), .A2(n604), .B1(f16[0]), .B2(n605), .ZN(n962) );
  NOR2_X1 U583 ( .A1(n920), .A2(n921), .ZN(n918) );
  OAI221_X1 U584 ( .B1(n601), .B2(n271), .C1(n602), .C2(n255), .A(n922), .ZN(
        n921) );
  OAI221_X1 U585 ( .B1(n606), .B2(n191), .C1(n923), .C2(n608), .A(n924), .ZN(
        n920) );
  AOI22_X1 U586 ( .A1(f13[1]), .A2(n604), .B1(f16[1]), .B2(n605), .ZN(n922) );
  NOR2_X1 U587 ( .A1(n898), .A2(n899), .ZN(n896) );
  OAI221_X1 U588 ( .B1(n601), .B2(n270), .C1(n602), .C2(n254), .A(n900), .ZN(
        n899) );
  OAI221_X1 U589 ( .B1(n606), .B2(n190), .C1(n901), .C2(n608), .A(n902), .ZN(
        n898) );
  AOI22_X1 U590 ( .A1(f13[2]), .A2(n604), .B1(f16[2]), .B2(n605), .ZN(n900) );
  NOR2_X1 U591 ( .A1(n876), .A2(n877), .ZN(n874) );
  OAI221_X1 U592 ( .B1(n601), .B2(n269), .C1(n602), .C2(n253), .A(n878), .ZN(
        n877) );
  OAI221_X1 U593 ( .B1(n606), .B2(n189), .C1(n879), .C2(n608), .A(n880), .ZN(
        n876) );
  AOI22_X1 U594 ( .A1(f13[3]), .A2(n604), .B1(f16[3]), .B2(n605), .ZN(n878) );
  NOR2_X1 U595 ( .A1(n854), .A2(n855), .ZN(n852) );
  OAI221_X1 U596 ( .B1(n601), .B2(n268), .C1(n602), .C2(n252), .A(n856), .ZN(
        n855) );
  OAI221_X1 U597 ( .B1(n606), .B2(n188), .C1(n857), .C2(n608), .A(n858), .ZN(
        n854) );
  AOI22_X1 U598 ( .A1(f13[4]), .A2(n604), .B1(f16[4]), .B2(n605), .ZN(n856) );
  NOR2_X1 U599 ( .A1(n832), .A2(n833), .ZN(n830) );
  OAI221_X1 U600 ( .B1(n601), .B2(n267), .C1(n602), .C2(n251), .A(n834), .ZN(
        n833) );
  OAI221_X1 U601 ( .B1(n606), .B2(n187), .C1(n835), .C2(n608), .A(n836), .ZN(
        n832) );
  AOI22_X1 U602 ( .A1(f13[5]), .A2(n604), .B1(f16[5]), .B2(n605), .ZN(n834) );
  NOR2_X1 U603 ( .A1(n810), .A2(n811), .ZN(n808) );
  OAI221_X1 U604 ( .B1(n601), .B2(n266), .C1(n602), .C2(n250), .A(n812), .ZN(
        n811) );
  OAI221_X1 U605 ( .B1(n606), .B2(n186), .C1(n813), .C2(n608), .A(n814), .ZN(
        n810) );
  AOI22_X1 U606 ( .A1(f13[6]), .A2(n604), .B1(f16[6]), .B2(n605), .ZN(n812) );
  NOR2_X1 U607 ( .A1(n788), .A2(n789), .ZN(n786) );
  OAI221_X1 U608 ( .B1(n601), .B2(n265), .C1(n602), .C2(n249), .A(n790), .ZN(
        n789) );
  OAI221_X1 U609 ( .B1(n606), .B2(n185), .C1(n791), .C2(n608), .A(n792), .ZN(
        n788) );
  AOI22_X1 U610 ( .A1(f13[7]), .A2(n604), .B1(f16[7]), .B2(n605), .ZN(n790) );
  NOR2_X1 U611 ( .A1(n766), .A2(n767), .ZN(n764) );
  OAI221_X1 U612 ( .B1(n601), .B2(n264), .C1(n602), .C2(n248), .A(n768), .ZN(
        n767) );
  OAI221_X1 U613 ( .B1(n606), .B2(n184), .C1(n769), .C2(n608), .A(n770), .ZN(
        n766) );
  AOI22_X1 U614 ( .A1(f13[8]), .A2(n604), .B1(f16[8]), .B2(n605), .ZN(n768) );
  NOR2_X1 U615 ( .A1(n744), .A2(n745), .ZN(n742) );
  OAI221_X1 U616 ( .B1(n601), .B2(n263), .C1(n602), .C2(n247), .A(n746), .ZN(
        n745) );
  OAI221_X1 U617 ( .B1(n606), .B2(n183), .C1(n747), .C2(n608), .A(n748), .ZN(
        n744) );
  AOI22_X1 U618 ( .A1(f13[9]), .A2(n604), .B1(f16[9]), .B2(n605), .ZN(n746) );
  NOR2_X1 U619 ( .A1(n722), .A2(n723), .ZN(n720) );
  OAI221_X1 U620 ( .B1(n601), .B2(n262), .C1(n602), .C2(n246), .A(n724), .ZN(
        n723) );
  OAI221_X1 U621 ( .B1(n606), .B2(n182), .C1(n725), .C2(n608), .A(n726), .ZN(
        n722) );
  AOI22_X1 U622 ( .A1(f13[10]), .A2(n604), .B1(f16[10]), .B2(n605), .ZN(n724)
         );
  NOR2_X1 U623 ( .A1(n700), .A2(n701), .ZN(n698) );
  OAI221_X1 U624 ( .B1(n601), .B2(n261), .C1(n602), .C2(n245), .A(n702), .ZN(
        n701) );
  OAI221_X1 U625 ( .B1(n606), .B2(n181), .C1(n703), .C2(n608), .A(n704), .ZN(
        n700) );
  AOI22_X1 U626 ( .A1(f13[11]), .A2(n604), .B1(f16[11]), .B2(n605), .ZN(n702)
         );
  NOR2_X1 U627 ( .A1(n678), .A2(n679), .ZN(n676) );
  OAI221_X1 U628 ( .B1(n601), .B2(n260), .C1(n602), .C2(n244), .A(n680), .ZN(
        n679) );
  OAI221_X1 U629 ( .B1(n606), .B2(n180), .C1(n681), .C2(n608), .A(n682), .ZN(
        n678) );
  AOI22_X1 U630 ( .A1(f13[12]), .A2(n604), .B1(f16[12]), .B2(n605), .ZN(n680)
         );
  NOR2_X1 U631 ( .A1(n656), .A2(n657), .ZN(n654) );
  OAI221_X1 U632 ( .B1(n601), .B2(n259), .C1(n602), .C2(n243), .A(n658), .ZN(
        n657) );
  OAI221_X1 U633 ( .B1(n606), .B2(n179), .C1(n659), .C2(n608), .A(n660), .ZN(
        n656) );
  AOI22_X1 U634 ( .A1(f13[13]), .A2(n604), .B1(f16[13]), .B2(n605), .ZN(n658)
         );
  NOR2_X1 U635 ( .A1(n634), .A2(n635), .ZN(n632) );
  OAI221_X1 U636 ( .B1(n601), .B2(n258), .C1(n602), .C2(n242), .A(n636), .ZN(
        n635) );
  OAI221_X1 U637 ( .B1(n606), .B2(n178), .C1(n637), .C2(n608), .A(n638), .ZN(
        n634) );
  AOI22_X1 U638 ( .A1(f13[14]), .A2(n604), .B1(f16[14]), .B2(n605), .ZN(n636)
         );
  NOR2_X1 U639 ( .A1(n599), .A2(n600), .ZN(n596) );
  OAI221_X1 U640 ( .B1(n601), .B2(n257), .C1(n602), .C2(n241), .A(n603), .ZN(
        n600) );
  OAI221_X1 U641 ( .B1(n606), .B2(n177), .C1(n607), .C2(n608), .A(n609), .ZN(
        n599) );
  AOI22_X1 U642 ( .A1(f13[15]), .A2(n604), .B1(f16[15]), .B2(n605), .ZN(n603)
         );
  NOR2_X1 U643 ( .A1(n971), .A2(n972), .ZN(n963) );
  OAI221_X1 U644 ( .B1(n612), .B2(n128), .C1(n613), .C2(n176), .A(n973), .ZN(
        n972) );
  OAI221_X1 U645 ( .B1(n617), .B2(n80), .C1(n618), .C2(n64), .A(n974), .ZN(
        n971) );
  AOI22_X1 U646 ( .A1(f8[0]), .A2(n615), .B1(f7[0]), .B2(n616), .ZN(n973) );
  NOR2_X1 U647 ( .A1(n925), .A2(n926), .ZN(n923) );
  OAI221_X1 U648 ( .B1(n612), .B2(n127), .C1(n613), .C2(n175), .A(n927), .ZN(
        n926) );
  OAI221_X1 U649 ( .B1(n617), .B2(n79), .C1(n618), .C2(n63), .A(n928), .ZN(
        n925) );
  AOI22_X1 U650 ( .A1(f8[1]), .A2(n615), .B1(f7[1]), .B2(n616), .ZN(n927) );
  NOR2_X1 U651 ( .A1(n903), .A2(n904), .ZN(n901) );
  OAI221_X1 U652 ( .B1(n612), .B2(n126), .C1(n613), .C2(n174), .A(n905), .ZN(
        n904) );
  OAI221_X1 U653 ( .B1(n617), .B2(n78), .C1(n618), .C2(n62), .A(n906), .ZN(
        n903) );
  AOI22_X1 U654 ( .A1(f8[2]), .A2(n615), .B1(f7[2]), .B2(n616), .ZN(n905) );
  NOR2_X1 U655 ( .A1(n881), .A2(n882), .ZN(n879) );
  OAI221_X1 U656 ( .B1(n612), .B2(n125), .C1(n613), .C2(n173), .A(n883), .ZN(
        n882) );
  OAI221_X1 U657 ( .B1(n617), .B2(n77), .C1(n618), .C2(n61), .A(n884), .ZN(
        n881) );
  AOI22_X1 U658 ( .A1(f8[3]), .A2(n615), .B1(f7[3]), .B2(n616), .ZN(n883) );
  NOR2_X1 U659 ( .A1(n859), .A2(n860), .ZN(n857) );
  OAI221_X1 U660 ( .B1(n612), .B2(n124), .C1(n613), .C2(n172), .A(n861), .ZN(
        n860) );
  OAI221_X1 U661 ( .B1(n617), .B2(n76), .C1(n618), .C2(n60), .A(n862), .ZN(
        n859) );
  AOI22_X1 U662 ( .A1(f8[4]), .A2(n615), .B1(f7[4]), .B2(n616), .ZN(n861) );
  NOR2_X1 U663 ( .A1(n837), .A2(n838), .ZN(n835) );
  OAI221_X1 U664 ( .B1(n612), .B2(n123), .C1(n613), .C2(n171), .A(n839), .ZN(
        n838) );
  OAI221_X1 U665 ( .B1(n617), .B2(n75), .C1(n618), .C2(n59), .A(n840), .ZN(
        n837) );
  AOI22_X1 U666 ( .A1(f8[5]), .A2(n615), .B1(f7[5]), .B2(n616), .ZN(n839) );
  NOR2_X1 U667 ( .A1(n815), .A2(n816), .ZN(n813) );
  OAI221_X1 U668 ( .B1(n612), .B2(n122), .C1(n613), .C2(n170), .A(n817), .ZN(
        n816) );
  OAI221_X1 U669 ( .B1(n617), .B2(n74), .C1(n618), .C2(n58), .A(n818), .ZN(
        n815) );
  AOI22_X1 U670 ( .A1(f8[6]), .A2(n615), .B1(f7[6]), .B2(n616), .ZN(n817) );
  NOR2_X1 U671 ( .A1(n793), .A2(n794), .ZN(n791) );
  OAI221_X1 U672 ( .B1(n612), .B2(n121), .C1(n613), .C2(n169), .A(n795), .ZN(
        n794) );
  OAI221_X1 U673 ( .B1(n617), .B2(n73), .C1(n618), .C2(n57), .A(n796), .ZN(
        n793) );
  AOI22_X1 U674 ( .A1(f8[7]), .A2(n615), .B1(f7[7]), .B2(n616), .ZN(n795) );
  NOR2_X1 U675 ( .A1(n771), .A2(n772), .ZN(n769) );
  OAI221_X1 U676 ( .B1(n612), .B2(n120), .C1(n613), .C2(n168), .A(n773), .ZN(
        n772) );
  OAI221_X1 U677 ( .B1(n617), .B2(n72), .C1(n618), .C2(n56), .A(n774), .ZN(
        n771) );
  AOI22_X1 U678 ( .A1(f8[8]), .A2(n615), .B1(f7[8]), .B2(n616), .ZN(n773) );
  NOR2_X1 U679 ( .A1(n749), .A2(n750), .ZN(n747) );
  OAI221_X1 U680 ( .B1(n612), .B2(n119), .C1(n613), .C2(n167), .A(n751), .ZN(
        n750) );
  OAI221_X1 U681 ( .B1(n617), .B2(n71), .C1(n618), .C2(n55), .A(n752), .ZN(
        n749) );
  AOI22_X1 U682 ( .A1(f8[9]), .A2(n615), .B1(f7[9]), .B2(n616), .ZN(n751) );
  NOR2_X1 U683 ( .A1(n727), .A2(n728), .ZN(n725) );
  OAI221_X1 U684 ( .B1(n612), .B2(n118), .C1(n613), .C2(n166), .A(n729), .ZN(
        n728) );
  OAI221_X1 U685 ( .B1(n617), .B2(n70), .C1(n618), .C2(n54), .A(n730), .ZN(
        n727) );
  AOI22_X1 U686 ( .A1(f8[10]), .A2(n615), .B1(f7[10]), .B2(n616), .ZN(n729) );
  NOR2_X1 U687 ( .A1(n705), .A2(n706), .ZN(n703) );
  OAI221_X1 U688 ( .B1(n612), .B2(n117), .C1(n613), .C2(n165), .A(n707), .ZN(
        n706) );
  OAI221_X1 U689 ( .B1(n617), .B2(n69), .C1(n618), .C2(n53), .A(n708), .ZN(
        n705) );
  AOI22_X1 U690 ( .A1(f8[11]), .A2(n615), .B1(f7[11]), .B2(n616), .ZN(n707) );
  NOR2_X1 U691 ( .A1(n683), .A2(n684), .ZN(n681) );
  OAI221_X1 U692 ( .B1(n612), .B2(n116), .C1(n613), .C2(n164), .A(n685), .ZN(
        n684) );
  OAI221_X1 U693 ( .B1(n617), .B2(n68), .C1(n618), .C2(n52), .A(n686), .ZN(
        n683) );
  AOI22_X1 U694 ( .A1(f8[12]), .A2(n615), .B1(f7[12]), .B2(n616), .ZN(n685) );
  NOR2_X1 U695 ( .A1(n661), .A2(n662), .ZN(n659) );
  OAI221_X1 U696 ( .B1(n612), .B2(n115), .C1(n613), .C2(n163), .A(n663), .ZN(
        n662) );
  OAI221_X1 U697 ( .B1(n617), .B2(n67), .C1(n618), .C2(n51), .A(n664), .ZN(
        n661) );
  AOI22_X1 U698 ( .A1(f8[13]), .A2(n615), .B1(f7[13]), .B2(n616), .ZN(n663) );
  NOR2_X1 U699 ( .A1(n639), .A2(n640), .ZN(n637) );
  OAI221_X1 U700 ( .B1(n612), .B2(n114), .C1(n613), .C2(n162), .A(n641), .ZN(
        n640) );
  OAI221_X1 U701 ( .B1(n617), .B2(n66), .C1(n618), .C2(n50), .A(n642), .ZN(
        n639) );
  AOI22_X1 U702 ( .A1(f8[14]), .A2(n615), .B1(f7[14]), .B2(n616), .ZN(n641) );
  NOR2_X1 U703 ( .A1(n610), .A2(n611), .ZN(n607) );
  OAI221_X1 U704 ( .B1(n612), .B2(n113), .C1(n613), .C2(n161), .A(n614), .ZN(
        n611) );
  OAI221_X1 U705 ( .B1(n617), .B2(n65), .C1(n618), .C2(n49), .A(n619), .ZN(
        n610) );
  AOI22_X1 U706 ( .A1(f8[15]), .A2(n615), .B1(f7[15]), .B2(n616), .ZN(n614) );
  INV_X1 U707 ( .A(addr_y[1]), .ZN(n2146) );
  INV_X1 U708 ( .A(addr_y[2]), .ZN(n2147) );
  OAI21_X1 U709 ( .B1(n2096), .B2(n438), .A(n1093), .ZN(n1621) );
  NAND2_X1 U710 ( .A1(add_r26[10]), .A2(n2071), .ZN(n1093) );
  OAI21_X1 U711 ( .B1(n2096), .B2(n437), .A(n1094), .ZN(n1622) );
  NAND2_X1 U712 ( .A1(add_r26[11]), .A2(n2071), .ZN(n1094) );
  OAI21_X1 U713 ( .B1(n2100), .B2(n390), .A(n1141), .ZN(n1669) );
  NAND2_X1 U714 ( .A1(add_r23[10]), .A2(n2040), .ZN(n1141) );
  OAI21_X1 U715 ( .B1(n2100), .B2(n389), .A(n1142), .ZN(n1670) );
  NAND2_X1 U716 ( .A1(add_r23[11]), .A2(n2038), .ZN(n1142) );
  OAI21_X1 U717 ( .B1(n2104), .B2(n342), .A(n1189), .ZN(n1717) );
  NAND2_X1 U718 ( .A1(add_r20[10]), .A2(n2080), .ZN(n1189) );
  OAI21_X1 U719 ( .B1(n2104), .B2(n341), .A(n1190), .ZN(n1718) );
  NAND2_X1 U720 ( .A1(add_r20[11]), .A2(n2046), .ZN(n1190) );
  OAI21_X1 U721 ( .B1(n2111), .B2(n294), .A(n1237), .ZN(n1765) );
  NAND2_X1 U722 ( .A1(add_r17[10]), .A2(n2043), .ZN(n1237) );
  OAI21_X1 U723 ( .B1(n2112), .B2(n293), .A(n1238), .ZN(n1766) );
  NAND2_X1 U724 ( .A1(add_r17[11]), .A2(n2046), .ZN(n1238) );
  OAI21_X1 U725 ( .B1(n2110), .B2(n246), .A(n1285), .ZN(n1813) );
  NAND2_X1 U726 ( .A1(add_r14[10]), .A2(n2064), .ZN(n1285) );
  OAI21_X1 U727 ( .B1(n2110), .B2(n245), .A(n1286), .ZN(n1814) );
  NAND2_X1 U728 ( .A1(add_r14[11]), .A2(n2064), .ZN(n1286) );
  OAI21_X1 U729 ( .B1(n2096), .B2(n102), .A(n1429), .ZN(n1957) );
  NAND2_X1 U730 ( .A1(add_r5[10]), .A2(n2052), .ZN(n1429) );
  OAI21_X1 U731 ( .B1(n2100), .B2(n101), .A(n1430), .ZN(n1958) );
  NAND2_X1 U732 ( .A1(add_r5[11]), .A2(n2052), .ZN(n1430) );
  OAI21_X1 U733 ( .B1(n2096), .B2(n448), .A(n1083), .ZN(n1611) );
  NAND2_X1 U734 ( .A1(add_r26[0]), .A2(n2072), .ZN(n1083) );
  OAI21_X1 U735 ( .B1(n2096), .B2(n447), .A(n1084), .ZN(n1612) );
  NAND2_X1 U736 ( .A1(add_r26[1]), .A2(n2072), .ZN(n1084) );
  OAI21_X1 U737 ( .B1(n2096), .B2(n446), .A(n1085), .ZN(n1613) );
  NAND2_X1 U738 ( .A1(add_r26[2]), .A2(n2072), .ZN(n1085) );
  OAI21_X1 U739 ( .B1(n2096), .B2(n445), .A(n1086), .ZN(n1614) );
  NAND2_X1 U740 ( .A1(add_r26[3]), .A2(n2072), .ZN(n1086) );
  OAI21_X1 U741 ( .B1(n2096), .B2(n444), .A(n1087), .ZN(n1615) );
  NAND2_X1 U742 ( .A1(add_r26[4]), .A2(n2072), .ZN(n1087) );
  OAI21_X1 U743 ( .B1(n2096), .B2(n443), .A(n1088), .ZN(n1616) );
  NAND2_X1 U744 ( .A1(add_r26[5]), .A2(n2072), .ZN(n1088) );
  OAI21_X1 U745 ( .B1(n2096), .B2(n442), .A(n1089), .ZN(n1617) );
  NAND2_X1 U746 ( .A1(add_r26[6]), .A2(n2072), .ZN(n1089) );
  OAI21_X1 U747 ( .B1(n2096), .B2(n441), .A(n1090), .ZN(n1618) );
  NAND2_X1 U748 ( .A1(add_r26[7]), .A2(n2072), .ZN(n1090) );
  OAI21_X1 U749 ( .B1(n2096), .B2(n440), .A(n1091), .ZN(n1619) );
  NAND2_X1 U750 ( .A1(add_r26[8]), .A2(n2071), .ZN(n1091) );
  OAI21_X1 U751 ( .B1(n2096), .B2(n439), .A(n1092), .ZN(n1620) );
  NAND2_X1 U752 ( .A1(add_r26[9]), .A2(n2071), .ZN(n1092) );
  OAI21_X1 U753 ( .B1(n2100), .B2(n400), .A(n1131), .ZN(n1659) );
  NAND2_X1 U754 ( .A1(add_r23[0]), .A2(n2068), .ZN(n1131) );
  OAI21_X1 U755 ( .B1(n2100), .B2(n399), .A(n1132), .ZN(n1660) );
  NAND2_X1 U756 ( .A1(add_r23[1]), .A2(n2068), .ZN(n1132) );
  OAI21_X1 U757 ( .B1(n2100), .B2(n398), .A(n1133), .ZN(n1661) );
  NAND2_X1 U758 ( .A1(add_r23[2]), .A2(n2068), .ZN(n1133) );
  OAI21_X1 U759 ( .B1(n2100), .B2(n397), .A(n1134), .ZN(n1662) );
  NAND2_X1 U760 ( .A1(add_r23[3]), .A2(n2068), .ZN(n1134) );
  OAI21_X1 U761 ( .B1(n2100), .B2(n396), .A(n1135), .ZN(n1663) );
  NAND2_X1 U762 ( .A1(add_r23[4]), .A2(n2068), .ZN(n1135) );
  OAI21_X1 U763 ( .B1(n2100), .B2(n395), .A(n1136), .ZN(n1664) );
  NAND2_X1 U764 ( .A1(add_r23[5]), .A2(n2068), .ZN(n1136) );
  OAI21_X1 U765 ( .B1(n2100), .B2(n394), .A(n1137), .ZN(n1665) );
  NAND2_X1 U766 ( .A1(add_r23[6]), .A2(n2068), .ZN(n1137) );
  OAI21_X1 U767 ( .B1(n2100), .B2(n393), .A(n1138), .ZN(n1666) );
  NAND2_X1 U768 ( .A1(add_r23[7]), .A2(n2068), .ZN(n1138) );
  OAI21_X1 U769 ( .B1(n2100), .B2(n392), .A(n1139), .ZN(n1667) );
  NAND2_X1 U770 ( .A1(add_r23[8]), .A2(n2037), .ZN(n1139) );
  OAI21_X1 U771 ( .B1(n2100), .B2(n391), .A(n1140), .ZN(n1668) );
  NAND2_X1 U772 ( .A1(add_r23[9]), .A2(n2036), .ZN(n1140) );
  OAI21_X1 U773 ( .B1(n2104), .B2(n352), .A(n1179), .ZN(n1707) );
  NAND2_X1 U774 ( .A1(add_r20[0]), .A2(n2040), .ZN(n1179) );
  OAI21_X1 U775 ( .B1(n2104), .B2(n351), .A(n1180), .ZN(n1708) );
  NAND2_X1 U776 ( .A1(add_r20[1]), .A2(n2045), .ZN(n1180) );
  OAI21_X1 U777 ( .B1(n2104), .B2(n350), .A(n1181), .ZN(n1709) );
  NAND2_X1 U778 ( .A1(add_r20[2]), .A2(n2040), .ZN(n1181) );
  OAI21_X1 U779 ( .B1(n2104), .B2(n349), .A(n1182), .ZN(n1710) );
  NAND2_X1 U780 ( .A1(add_r20[3]), .A2(n2043), .ZN(n1182) );
  OAI21_X1 U781 ( .B1(n2104), .B2(n348), .A(n1183), .ZN(n1711) );
  NAND2_X1 U782 ( .A1(add_r20[4]), .A2(n2045), .ZN(n1183) );
  OAI21_X1 U783 ( .B1(n2104), .B2(n347), .A(n1184), .ZN(n1712) );
  NAND2_X1 U784 ( .A1(add_r20[5]), .A2(n2045), .ZN(n1184) );
  OAI21_X1 U785 ( .B1(n2104), .B2(n346), .A(n1185), .ZN(n1713) );
  NAND2_X1 U786 ( .A1(add_r20[6]), .A2(n2046), .ZN(n1185) );
  OAI21_X1 U787 ( .B1(n2104), .B2(n345), .A(n1186), .ZN(n1714) );
  NAND2_X1 U788 ( .A1(add_r20[7]), .A2(n2041), .ZN(n1186) );
  OAI21_X1 U789 ( .B1(n2104), .B2(n344), .A(n1187), .ZN(n1715) );
  NAND2_X1 U790 ( .A1(add_r20[8]), .A2(n2043), .ZN(n1187) );
  OAI21_X1 U791 ( .B1(n2104), .B2(n343), .A(n1188), .ZN(n1716) );
  NAND2_X1 U792 ( .A1(add_r20[9]), .A2(n2046), .ZN(n1188) );
  OAI21_X1 U793 ( .B1(n2111), .B2(n304), .A(n1227), .ZN(n1755) );
  NAND2_X1 U794 ( .A1(add_r17[0]), .A2(n2045), .ZN(n1227) );
  OAI21_X1 U795 ( .B1(n2112), .B2(n303), .A(n1228), .ZN(n1756) );
  NAND2_X1 U796 ( .A1(add_r17[1]), .A2(n2040), .ZN(n1228) );
  OAI21_X1 U797 ( .B1(n2113), .B2(n302), .A(n1229), .ZN(n1757) );
  NAND2_X1 U798 ( .A1(add_r17[2]), .A2(n2039), .ZN(n1229) );
  OAI21_X1 U799 ( .B1(n2111), .B2(n301), .A(n1230), .ZN(n1758) );
  NAND2_X1 U800 ( .A1(add_r17[3]), .A2(n2041), .ZN(n1230) );
  OAI21_X1 U801 ( .B1(n2112), .B2(n300), .A(n1231), .ZN(n1759) );
  NAND2_X1 U802 ( .A1(add_r17[4]), .A2(n2040), .ZN(n1231) );
  OAI21_X1 U803 ( .B1(n2113), .B2(n299), .A(n1232), .ZN(n1760) );
  NAND2_X1 U804 ( .A1(add_r17[5]), .A2(n2045), .ZN(n1232) );
  OAI21_X1 U805 ( .B1(n2111), .B2(n298), .A(n1233), .ZN(n1761) );
  NAND2_X1 U806 ( .A1(add_r17[6]), .A2(n2080), .ZN(n1233) );
  OAI21_X1 U807 ( .B1(n2112), .B2(n297), .A(n1234), .ZN(n1762) );
  NAND2_X1 U808 ( .A1(add_r17[7]), .A2(n2080), .ZN(n1234) );
  OAI21_X1 U809 ( .B1(n2113), .B2(n296), .A(n1235), .ZN(n1763) );
  NAND2_X1 U810 ( .A1(add_r17[8]), .A2(n2041), .ZN(n1235) );
  OAI21_X1 U811 ( .B1(n2111), .B2(n295), .A(n1236), .ZN(n1764) );
  NAND2_X1 U812 ( .A1(add_r17[9]), .A2(n2042), .ZN(n1236) );
  OAI21_X1 U813 ( .B1(n2110), .B2(n256), .A(n1275), .ZN(n1803) );
  NAND2_X1 U814 ( .A1(add_r14[0]), .A2(n2065), .ZN(n1275) );
  OAI21_X1 U815 ( .B1(n2110), .B2(n255), .A(n1276), .ZN(n1804) );
  NAND2_X1 U816 ( .A1(add_r14[1]), .A2(n2065), .ZN(n1276) );
  OAI21_X1 U817 ( .B1(n2110), .B2(n254), .A(n1277), .ZN(n1805) );
  NAND2_X1 U818 ( .A1(add_r14[2]), .A2(n2065), .ZN(n1277) );
  OAI21_X1 U819 ( .B1(n2110), .B2(n253), .A(n1278), .ZN(n1806) );
  NAND2_X1 U820 ( .A1(add_r14[3]), .A2(n2065), .ZN(n1278) );
  OAI21_X1 U821 ( .B1(n2110), .B2(n252), .A(n1279), .ZN(n1807) );
  NAND2_X1 U822 ( .A1(add_r14[4]), .A2(n2065), .ZN(n1279) );
  OAI21_X1 U823 ( .B1(n2110), .B2(n250), .A(n1281), .ZN(n1809) );
  NAND2_X1 U824 ( .A1(add_r14[6]), .A2(n2065), .ZN(n1281) );
  OAI21_X1 U825 ( .B1(n2110), .B2(n249), .A(n1282), .ZN(n1810) );
  NAND2_X1 U826 ( .A1(add_r14[7]), .A2(n2065), .ZN(n1282) );
  OAI21_X1 U827 ( .B1(n2110), .B2(n248), .A(n1283), .ZN(n1811) );
  NAND2_X1 U828 ( .A1(add_r14[8]), .A2(n2064), .ZN(n1283) );
  OAI21_X1 U829 ( .B1(n2110), .B2(n247), .A(n1284), .ZN(n1812) );
  NAND2_X1 U830 ( .A1(add_r14[9]), .A2(n2064), .ZN(n1284) );
  OAI21_X1 U831 ( .B1(n2088), .B2(n112), .A(n1419), .ZN(n1947) );
  NAND2_X1 U832 ( .A1(add_r5[0]), .A2(n2053), .ZN(n1419) );
  OAI21_X1 U833 ( .B1(n2092), .B2(n111), .A(n1420), .ZN(n1948) );
  NAND2_X1 U834 ( .A1(add_r5[1]), .A2(n2053), .ZN(n1420) );
  OAI21_X1 U835 ( .B1(n2104), .B2(n110), .A(n1421), .ZN(n1949) );
  NAND2_X1 U836 ( .A1(add_r5[2]), .A2(n2053), .ZN(n1421) );
  OAI21_X1 U837 ( .B1(n2112), .B2(n109), .A(n1422), .ZN(n1950) );
  NAND2_X1 U838 ( .A1(add_r5[3]), .A2(n2053), .ZN(n1422) );
  OAI21_X1 U839 ( .B1(n2110), .B2(n108), .A(n1423), .ZN(n1951) );
  NAND2_X1 U840 ( .A1(add_r5[4]), .A2(n2053), .ZN(n1423) );
  OAI21_X1 U841 ( .B1(n2116), .B2(n107), .A(n1424), .ZN(n1952) );
  NAND2_X1 U842 ( .A1(add_r5[5]), .A2(n2053), .ZN(n1424) );
  OAI21_X1 U843 ( .B1(n2113), .B2(n106), .A(n1425), .ZN(n1953) );
  NAND2_X1 U844 ( .A1(add_r5[6]), .A2(n2053), .ZN(n1425) );
  OAI21_X1 U845 ( .B1(n2116), .B2(n105), .A(n1426), .ZN(n1954) );
  NAND2_X1 U846 ( .A1(add_r5[7]), .A2(n2053), .ZN(n1426) );
  OAI21_X1 U847 ( .B1(n2096), .B2(n104), .A(n1427), .ZN(n1955) );
  NAND2_X1 U848 ( .A1(add_r5[8]), .A2(n2052), .ZN(n1427) );
  OAI21_X1 U849 ( .B1(n2100), .B2(n103), .A(n1428), .ZN(n1956) );
  NAND2_X1 U850 ( .A1(add_r5[9]), .A2(n2052), .ZN(n1428) );
  OAI21_X1 U851 ( .B1(n2088), .B2(n534), .A(n995), .ZN(n1525) );
  NAND2_X1 U852 ( .A1(add_r32[10]), .A2(n2079), .ZN(n995) );
  OAI21_X1 U853 ( .B1(n2088), .B2(n533), .A(n996), .ZN(n1526) );
  NAND2_X1 U854 ( .A1(add_r32[11]), .A2(n2079), .ZN(n996) );
  OAI21_X1 U855 ( .B1(n2092), .B2(n486), .A(n1045), .ZN(n1573) );
  NAND2_X1 U856 ( .A1(add_r29[10]), .A2(n2075), .ZN(n1045) );
  OAI21_X1 U857 ( .B1(n2092), .B2(n485), .A(n1046), .ZN(n1574) );
  NAND2_X1 U858 ( .A1(add_r29[11]), .A2(n2075), .ZN(n1046) );
  OAI21_X1 U859 ( .B1(n2113), .B2(n198), .A(n1333), .ZN(n1861) );
  NAND2_X1 U860 ( .A1(add_r11[10]), .A2(n2060), .ZN(n1333) );
  OAI21_X1 U861 ( .B1(n2113), .B2(n197), .A(n1334), .ZN(n1862) );
  NAND2_X1 U862 ( .A1(add_r11[11]), .A2(n2060), .ZN(n1334) );
  OAI21_X1 U863 ( .B1(n2116), .B2(n150), .A(n1381), .ZN(n1909) );
  NAND2_X1 U864 ( .A1(add_r8[10]), .A2(n2056), .ZN(n1381) );
  OAI21_X1 U865 ( .B1(n2116), .B2(n149), .A(n1382), .ZN(n1910) );
  NAND2_X1 U866 ( .A1(add_r8[11]), .A2(n2056), .ZN(n1382) );
  OAI21_X1 U867 ( .B1(n2088), .B2(n544), .A(n984), .ZN(n1515) );
  NAND2_X1 U868 ( .A1(add_r32[0]), .A2(n2080), .ZN(n984) );
  OAI21_X1 U869 ( .B1(n2088), .B2(n543), .A(n986), .ZN(n1516) );
  NAND2_X1 U870 ( .A1(add_r32[1]), .A2(n2080), .ZN(n986) );
  OAI21_X1 U871 ( .B1(n2088), .B2(n542), .A(n987), .ZN(n1517) );
  NAND2_X1 U872 ( .A1(add_r32[2]), .A2(n2080), .ZN(n987) );
  OAI21_X1 U873 ( .B1(n2088), .B2(n541), .A(n988), .ZN(n1518) );
  NAND2_X1 U874 ( .A1(add_r32[3]), .A2(n2080), .ZN(n988) );
  OAI21_X1 U875 ( .B1(n2088), .B2(n540), .A(n989), .ZN(n1519) );
  NAND2_X1 U876 ( .A1(add_r32[4]), .A2(n2080), .ZN(n989) );
  OAI21_X1 U877 ( .B1(n2088), .B2(n539), .A(n990), .ZN(n1520) );
  NAND2_X1 U878 ( .A1(add_r32[5]), .A2(n2080), .ZN(n990) );
  OAI21_X1 U879 ( .B1(n2088), .B2(n538), .A(n991), .ZN(n1521) );
  NAND2_X1 U880 ( .A1(add_r32[6]), .A2(n2079), .ZN(n991) );
  OAI21_X1 U881 ( .B1(n2088), .B2(n537), .A(n992), .ZN(n1522) );
  NAND2_X1 U882 ( .A1(add_r32[7]), .A2(n2079), .ZN(n992) );
  OAI21_X1 U883 ( .B1(n2088), .B2(n536), .A(n993), .ZN(n1523) );
  NAND2_X1 U884 ( .A1(add_r32[8]), .A2(n2079), .ZN(n993) );
  OAI21_X1 U885 ( .B1(n2088), .B2(n535), .A(n994), .ZN(n1524) );
  NAND2_X1 U886 ( .A1(add_r32[9]), .A2(n2079), .ZN(n994) );
  OAI21_X1 U887 ( .B1(n2092), .B2(n496), .A(n1035), .ZN(n1563) );
  NAND2_X1 U888 ( .A1(add_r29[0]), .A2(n2076), .ZN(n1035) );
  OAI21_X1 U889 ( .B1(n2092), .B2(n495), .A(n1036), .ZN(n1564) );
  NAND2_X1 U890 ( .A1(add_r29[1]), .A2(n2076), .ZN(n1036) );
  OAI21_X1 U891 ( .B1(n2092), .B2(n494), .A(n1037), .ZN(n1565) );
  NAND2_X1 U892 ( .A1(add_r29[2]), .A2(n2076), .ZN(n1037) );
  OAI21_X1 U893 ( .B1(n2092), .B2(n493), .A(n1038), .ZN(n1566) );
  NAND2_X1 U894 ( .A1(add_r29[3]), .A2(n2076), .ZN(n1038) );
  OAI21_X1 U895 ( .B1(n2092), .B2(n492), .A(n1039), .ZN(n1567) );
  NAND2_X1 U896 ( .A1(add_r29[4]), .A2(n2076), .ZN(n1039) );
  OAI21_X1 U897 ( .B1(n2092), .B2(n491), .A(n1040), .ZN(n1568) );
  NAND2_X1 U898 ( .A1(add_r29[5]), .A2(n2076), .ZN(n1040) );
  OAI21_X1 U899 ( .B1(n2092), .B2(n490), .A(n1041), .ZN(n1569) );
  NAND2_X1 U900 ( .A1(add_r29[6]), .A2(n2076), .ZN(n1041) );
  OAI21_X1 U901 ( .B1(n2092), .B2(n489), .A(n1042), .ZN(n1570) );
  NAND2_X1 U902 ( .A1(add_r29[7]), .A2(n2076), .ZN(n1042) );
  OAI21_X1 U903 ( .B1(n2092), .B2(n488), .A(n1043), .ZN(n1571) );
  NAND2_X1 U904 ( .A1(add_r29[8]), .A2(n2075), .ZN(n1043) );
  OAI21_X1 U905 ( .B1(n2092), .B2(n487), .A(n1044), .ZN(n1572) );
  NAND2_X1 U906 ( .A1(add_r29[9]), .A2(n2075), .ZN(n1044) );
  OAI21_X1 U907 ( .B1(n2113), .B2(n208), .A(n1323), .ZN(n1851) );
  NAND2_X1 U908 ( .A1(add_r11[0]), .A2(n2061), .ZN(n1323) );
  OAI21_X1 U909 ( .B1(n2113), .B2(n207), .A(n1324), .ZN(n1852) );
  NAND2_X1 U910 ( .A1(add_r11[1]), .A2(n2061), .ZN(n1324) );
  OAI21_X1 U911 ( .B1(n2113), .B2(n206), .A(n1325), .ZN(n1853) );
  NAND2_X1 U912 ( .A1(add_r11[2]), .A2(n2061), .ZN(n1325) );
  OAI21_X1 U913 ( .B1(n2113), .B2(n205), .A(n1326), .ZN(n1854) );
  NAND2_X1 U914 ( .A1(add_r11[3]), .A2(n2061), .ZN(n1326) );
  OAI21_X1 U915 ( .B1(n2113), .B2(n204), .A(n1327), .ZN(n1855) );
  NAND2_X1 U916 ( .A1(add_r11[4]), .A2(n2061), .ZN(n1327) );
  OAI21_X1 U917 ( .B1(n2113), .B2(n202), .A(n1329), .ZN(n1857) );
  NAND2_X1 U918 ( .A1(add_r11[6]), .A2(n2061), .ZN(n1329) );
  OAI21_X1 U919 ( .B1(n2113), .B2(n201), .A(n1330), .ZN(n1858) );
  NAND2_X1 U920 ( .A1(add_r11[7]), .A2(n2061), .ZN(n1330) );
  OAI21_X1 U921 ( .B1(n2113), .B2(n200), .A(n1331), .ZN(n1859) );
  NAND2_X1 U922 ( .A1(add_r11[8]), .A2(n2060), .ZN(n1331) );
  OAI21_X1 U923 ( .B1(n2113), .B2(n199), .A(n1332), .ZN(n1860) );
  NAND2_X1 U924 ( .A1(add_r11[9]), .A2(n2060), .ZN(n1332) );
  OAI21_X1 U925 ( .B1(n2116), .B2(n160), .A(n1371), .ZN(n1899) );
  NAND2_X1 U926 ( .A1(add_r8[0]), .A2(n2057), .ZN(n1371) );
  OAI21_X1 U927 ( .B1(n2116), .B2(n159), .A(n1372), .ZN(n1900) );
  NAND2_X1 U928 ( .A1(add_r8[1]), .A2(n2057), .ZN(n1372) );
  OAI21_X1 U929 ( .B1(n2116), .B2(n158), .A(n1373), .ZN(n1901) );
  NAND2_X1 U930 ( .A1(add_r8[2]), .A2(n2057), .ZN(n1373) );
  OAI21_X1 U931 ( .B1(n2116), .B2(n157), .A(n1374), .ZN(n1902) );
  NAND2_X1 U932 ( .A1(add_r8[3]), .A2(n2057), .ZN(n1374) );
  OAI21_X1 U933 ( .B1(n2116), .B2(n156), .A(n1375), .ZN(n1903) );
  NAND2_X1 U934 ( .A1(add_r8[4]), .A2(n2057), .ZN(n1375) );
  OAI21_X1 U935 ( .B1(n2116), .B2(n155), .A(n1376), .ZN(n1904) );
  NAND2_X1 U936 ( .A1(add_r8[5]), .A2(n2057), .ZN(n1376) );
  OAI21_X1 U937 ( .B1(n2116), .B2(n154), .A(n1377), .ZN(n1905) );
  NAND2_X1 U938 ( .A1(add_r8[6]), .A2(n2057), .ZN(n1377) );
  OAI21_X1 U939 ( .B1(n2116), .B2(n153), .A(n1378), .ZN(n1906) );
  NAND2_X1 U940 ( .A1(add_r8[7]), .A2(n2057), .ZN(n1378) );
  OAI21_X1 U941 ( .B1(n2116), .B2(n152), .A(n1379), .ZN(n1907) );
  NAND2_X1 U942 ( .A1(add_r8[8]), .A2(n2056), .ZN(n1379) );
  OAI21_X1 U943 ( .B1(n2116), .B2(n151), .A(n1380), .ZN(n1908) );
  NAND2_X1 U944 ( .A1(add_r8[9]), .A2(n2056), .ZN(n1380) );
  OAI21_X1 U945 ( .B1(n2094), .B2(n54), .A(n1477), .ZN(n2005) );
  NAND2_X1 U946 ( .A1(add_r2[10]), .A2(n2048), .ZN(n1477) );
  OAI21_X1 U947 ( .B1(n2095), .B2(n53), .A(n1478), .ZN(n2006) );
  NAND2_X1 U948 ( .A1(add_r2[11]), .A2(n2048), .ZN(n1478) );
  OAI21_X1 U949 ( .B1(n2097), .B2(n64), .A(n1467), .ZN(n1995) );
  NAND2_X1 U950 ( .A1(add_r2[0]), .A2(n2049), .ZN(n1467) );
  OAI21_X1 U951 ( .B1(n2098), .B2(n63), .A(n1468), .ZN(n1996) );
  NAND2_X1 U952 ( .A1(add_r2[1]), .A2(n2049), .ZN(n1468) );
  OAI21_X1 U953 ( .B1(n2101), .B2(n62), .A(n1469), .ZN(n1997) );
  NAND2_X1 U954 ( .A1(add_r2[2]), .A2(n2049), .ZN(n1469) );
  OAI21_X1 U955 ( .B1(n2091), .B2(n61), .A(n1470), .ZN(n1998) );
  NAND2_X1 U956 ( .A1(add_r2[3]), .A2(n2049), .ZN(n1470) );
  OAI21_X1 U957 ( .B1(n2108), .B2(n60), .A(n1471), .ZN(n1999) );
  NAND2_X1 U958 ( .A1(add_r2[4]), .A2(n2049), .ZN(n1471) );
  OAI21_X1 U959 ( .B1(n2109), .B2(n59), .A(n1472), .ZN(n2000) );
  NAND2_X1 U960 ( .A1(add_r2[5]), .A2(n2049), .ZN(n1472) );
  OAI21_X1 U961 ( .B1(n2112), .B2(n58), .A(n1473), .ZN(n2001) );
  NAND2_X1 U962 ( .A1(add_r2[6]), .A2(n2049), .ZN(n1473) );
  OAI21_X1 U963 ( .B1(n2090), .B2(n57), .A(n1474), .ZN(n2002) );
  NAND2_X1 U964 ( .A1(add_r2[7]), .A2(n2049), .ZN(n1474) );
  OAI21_X1 U965 ( .B1(n2096), .B2(n56), .A(n1475), .ZN(n2003) );
  NAND2_X1 U966 ( .A1(add_r2[8]), .A2(n2048), .ZN(n1475) );
  OAI21_X1 U967 ( .B1(n2085), .B2(n55), .A(n1476), .ZN(n2004) );
  NAND2_X1 U968 ( .A1(add_r2[9]), .A2(n2048), .ZN(n1476) );
  OAI21_X1 U969 ( .B1(n2094), .B2(n470), .A(n1061), .ZN(n1589) );
  NAND2_X1 U970 ( .A1(add_r28[10]), .A2(n2074), .ZN(n1061) );
  OAI21_X1 U971 ( .B1(n2094), .B2(n469), .A(n1062), .ZN(n1590) );
  NAND2_X1 U972 ( .A1(add_r28[11]), .A2(n2074), .ZN(n1062) );
  OAI21_X1 U973 ( .B1(n2095), .B2(n454), .A(n1077), .ZN(n1605) );
  NAND2_X1 U974 ( .A1(add_r27[10]), .A2(n2073), .ZN(n1077) );
  OAI21_X1 U975 ( .B1(n2095), .B2(n453), .A(n1078), .ZN(n1606) );
  NAND2_X1 U976 ( .A1(add_r27[11]), .A2(n2073), .ZN(n1078) );
  OAI21_X1 U977 ( .B1(n2098), .B2(n422), .A(n1109), .ZN(n1637) );
  NAND2_X1 U978 ( .A1(add_r25[10]), .A2(n2070), .ZN(n1109) );
  OAI21_X1 U979 ( .B1(n2098), .B2(n421), .A(n1110), .ZN(n1638) );
  NAND2_X1 U980 ( .A1(add_r25[11]), .A2(n2070), .ZN(n1110) );
  OAI21_X1 U981 ( .B1(n2099), .B2(n406), .A(n1125), .ZN(n1653) );
  NAND2_X1 U982 ( .A1(add_r24[10]), .A2(n2069), .ZN(n1125) );
  OAI21_X1 U983 ( .B1(n2099), .B2(n405), .A(n1126), .ZN(n1654) );
  NAND2_X1 U984 ( .A1(add_r24[11]), .A2(n2069), .ZN(n1126) );
  OAI21_X1 U985 ( .B1(n2102), .B2(n374), .A(n1157), .ZN(n1685) );
  NAND2_X1 U986 ( .A1(add_r22[10]), .A2(n2043), .ZN(n1157) );
  OAI21_X1 U987 ( .B1(n2102), .B2(n373), .A(n1158), .ZN(n1686) );
  NAND2_X1 U988 ( .A1(add_r22[11]), .A2(n2043), .ZN(n1158) );
  OAI21_X1 U989 ( .B1(n2103), .B2(n358), .A(n1173), .ZN(n1701) );
  NAND2_X1 U990 ( .A1(add_r21[10]), .A2(n2067), .ZN(n1173) );
  OAI21_X1 U991 ( .B1(n2103), .B2(n357), .A(n1174), .ZN(n1702) );
  NAND2_X1 U992 ( .A1(add_r21[11]), .A2(n2067), .ZN(n1174) );
  OAI21_X1 U993 ( .B1(n2106), .B2(n326), .A(n1205), .ZN(n1733) );
  NAND2_X1 U994 ( .A1(add_r19[10]), .A2(n2041), .ZN(n1205) );
  OAI21_X1 U995 ( .B1(n2106), .B2(n325), .A(n1206), .ZN(n1734) );
  NAND2_X1 U996 ( .A1(add_r19[11]), .A2(n2042), .ZN(n1206) );
  OAI21_X1 U997 ( .B1(n2107), .B2(n310), .A(n1221), .ZN(n1749) );
  NAND2_X1 U998 ( .A1(add_r18[10]), .A2(n2042), .ZN(n1221) );
  OAI21_X1 U999 ( .B1(n2107), .B2(n309), .A(n1222), .ZN(n1750) );
  NAND2_X1 U1000 ( .A1(add_r18[11]), .A2(n2044), .ZN(n1222) );
  OAI21_X1 U1001 ( .B1(n2109), .B2(n278), .A(n1253), .ZN(n1781) );
  NAND2_X1 U1002 ( .A1(add_r16[10]), .A2(n985), .ZN(n1253) );
  OAI21_X1 U1003 ( .B1(n2109), .B2(n277), .A(n1254), .ZN(n1782) );
  NAND2_X1 U1004 ( .A1(add_r16[11]), .A2(n985), .ZN(n1254) );
  OAI21_X1 U1005 ( .B1(n2113), .B2(n262), .A(n1269), .ZN(n1797) );
  NAND2_X1 U1006 ( .A1(add_r15[10]), .A2(n2066), .ZN(n1269) );
  OAI21_X1 U1007 ( .B1(n2112), .B2(n261), .A(n1270), .ZN(n1798) );
  NAND2_X1 U1008 ( .A1(add_r15[11]), .A2(n2066), .ZN(n1270) );
  OAI21_X1 U1009 ( .B1(n2116), .B2(n118), .A(n1413), .ZN(n1941) );
  NAND2_X1 U1010 ( .A1(add_r6[10]), .A2(n2054), .ZN(n1413) );
  OAI21_X1 U1011 ( .B1(n2113), .B2(n117), .A(n1414), .ZN(n1942) );
  NAND2_X1 U1012 ( .A1(add_r6[11]), .A2(n2054), .ZN(n1414) );
  OAI21_X1 U1013 ( .B1(n2119), .B2(n86), .A(n1445), .ZN(n1973) );
  NAND2_X1 U1014 ( .A1(add_r4[10]), .A2(n2051), .ZN(n1445) );
  OAI21_X1 U1015 ( .B1(n2119), .B2(n85), .A(n1446), .ZN(n1974) );
  NAND2_X1 U1016 ( .A1(add_r4[11]), .A2(n2051), .ZN(n1446) );
  OAI21_X1 U1017 ( .B1(n2120), .B2(n70), .A(n1461), .ZN(n1989) );
  NAND2_X1 U1018 ( .A1(add_r3[10]), .A2(n2050), .ZN(n1461) );
  OAI21_X1 U1019 ( .B1(n2120), .B2(n69), .A(n1462), .ZN(n1990) );
  NAND2_X1 U1020 ( .A1(add_r3[11]), .A2(n2050), .ZN(n1462) );
  NAND2_X1 U1021 ( .A1(add_r28[14]), .A2(n2074), .ZN(n1065) );
  NAND2_X1 U1022 ( .A1(add_r17[14]), .A2(n2044), .ZN(n1241) );
  OAI21_X1 U1023 ( .B1(n2103), .B2(n354), .A(n1177), .ZN(n1705) );
  NAND2_X1 U1024 ( .A1(add_r21[14]), .A2(n2042), .ZN(n1177) );
  OAI21_X1 U1025 ( .B1(n2102), .B2(n370), .A(n1161), .ZN(n1689) );
  NAND2_X1 U1026 ( .A1(add_r22[14]), .A2(n2040), .ZN(n1161) );
  NAND2_X1 U1027 ( .A1(add_r26[14]), .A2(n2071), .ZN(n1097) );
  OAI21_X1 U1028 ( .B1(n2107), .B2(n306), .A(n1225), .ZN(n1753) );
  NAND2_X1 U1029 ( .A1(add_r18[14]), .A2(n2045), .ZN(n1225) );
  OAI21_X1 U1030 ( .B1(n2106), .B2(n322), .A(n1209), .ZN(n1737) );
  NAND2_X1 U1031 ( .A1(add_r19[14]), .A2(n2044), .ZN(n1209) );
  OAI21_X1 U1032 ( .B1(n2110), .B2(n258), .A(n1273), .ZN(n1801) );
  NAND2_X1 U1033 ( .A1(add_r15[14]), .A2(n2065), .ZN(n1273) );
  OAI21_X1 U1034 ( .B1(n2099), .B2(n402), .A(n1129), .ZN(n1657) );
  NAND2_X1 U1035 ( .A1(add_r24[14]), .A2(n2068), .ZN(n1129) );
  OAI21_X1 U1036 ( .B1(n2105), .B2(n338), .A(n1193), .ZN(n1721) );
  NAND2_X1 U1037 ( .A1(add_r20[14]), .A2(n2040), .ZN(n1193) );
  NAND2_X1 U1038 ( .A1(add_r16[14]), .A2(n2046), .ZN(n1257) );
  NAND2_X1 U1039 ( .A1(add_r27[14]), .A2(n2072), .ZN(n1081) );
  OAI21_X1 U1040 ( .B1(n2093), .B2(n482), .A(n1049), .ZN(n1577) );
  NAND2_X1 U1041 ( .A1(add_r29[14]), .A2(n2075), .ZN(n1049) );
  NAND2_X1 U1042 ( .A1(add_r25[14]), .A2(n2070), .ZN(n1113) );
  NAND2_X1 U1043 ( .A1(add_r23[14]), .A2(n2039), .ZN(n1145) );
  OAI21_X1 U1044 ( .B1(n2120), .B2(n66), .A(n1465), .ZN(n1993) );
  NAND2_X1 U1045 ( .A1(add_r3[14]), .A2(n2049), .ZN(n1465) );
  OAI21_X1 U1046 ( .B1(n2119), .B2(n82), .A(n1449), .ZN(n1977) );
  NAND2_X1 U1047 ( .A1(add_r4[14]), .A2(n2051), .ZN(n1449) );
  OAI21_X1 U1048 ( .B1(n2116), .B2(n114), .A(n1417), .ZN(n1945) );
  NAND2_X1 U1049 ( .A1(add_r6[14]), .A2(n2053), .ZN(n1417) );
  OAI21_X1 U1050 ( .B1(n2112), .B2(n98), .A(n1433), .ZN(n1961) );
  NAND2_X1 U1051 ( .A1(add_r5[14]), .A2(n2052), .ZN(n1433) );
  OAI21_X1 U1052 ( .B1(n2094), .B2(n467), .A(n1064), .ZN(n1592) );
  NAND2_X1 U1053 ( .A1(add_r28[13]), .A2(n2074), .ZN(n1064) );
  OAI21_X1 U1054 ( .B1(n2108), .B2(n291), .A(n1240), .ZN(n1768) );
  NAND2_X1 U1055 ( .A1(add_r17[13]), .A2(n2044), .ZN(n1240) );
  OAI21_X1 U1056 ( .B1(n2103), .B2(n355), .A(n1176), .ZN(n1704) );
  NAND2_X1 U1057 ( .A1(add_r21[13]), .A2(n2044), .ZN(n1176) );
  OAI21_X1 U1058 ( .B1(n2106), .B2(n323), .A(n1208), .ZN(n1736) );
  NAND2_X1 U1059 ( .A1(add_r19[13]), .A2(n2038), .ZN(n1208) );
  OAI21_X1 U1060 ( .B1(n2107), .B2(n307), .A(n1224), .ZN(n1752) );
  NAND2_X1 U1061 ( .A1(add_r18[13]), .A2(n2043), .ZN(n1224) );
  OAI21_X1 U1062 ( .B1(n2104), .B2(n259), .A(n1272), .ZN(n1800) );
  NAND2_X1 U1063 ( .A1(add_r15[13]), .A2(n2065), .ZN(n1272) );
  OAI21_X1 U1064 ( .B1(n2102), .B2(n371), .A(n1160), .ZN(n1688) );
  NAND2_X1 U1065 ( .A1(add_r22[13]), .A2(n2041), .ZN(n1160) );
  OAI21_X1 U1066 ( .B1(n2097), .B2(n435), .A(n1096), .ZN(n1624) );
  NAND2_X1 U1067 ( .A1(add_r26[13]), .A2(n2071), .ZN(n1096) );
  OAI21_X1 U1068 ( .B1(n2099), .B2(n403), .A(n1128), .ZN(n1656) );
  NAND2_X1 U1069 ( .A1(add_r24[13]), .A2(n2068), .ZN(n1128) );
  OAI21_X1 U1070 ( .B1(n2105), .B2(n339), .A(n1192), .ZN(n1720) );
  NAND2_X1 U1071 ( .A1(add_r20[13]), .A2(n2039), .ZN(n1192) );
  OAI21_X1 U1072 ( .B1(n2109), .B2(n275), .A(n1256), .ZN(n1784) );
  NAND2_X1 U1073 ( .A1(add_r16[13]), .A2(n2039), .ZN(n1256) );
  OAI21_X1 U1074 ( .B1(n2095), .B2(n451), .A(n1080), .ZN(n1608) );
  NAND2_X1 U1075 ( .A1(add_r27[13]), .A2(n2072), .ZN(n1080) );
  OAI21_X1 U1076 ( .B1(n2093), .B2(n483), .A(n1048), .ZN(n1576) );
  NAND2_X1 U1077 ( .A1(add_r29[13]), .A2(n2075), .ZN(n1048) );
  OAI21_X1 U1078 ( .B1(n2098), .B2(n419), .A(n1112), .ZN(n1640) );
  NAND2_X1 U1079 ( .A1(add_r25[13]), .A2(n2070), .ZN(n1112) );
  OAI21_X1 U1080 ( .B1(n2101), .B2(n387), .A(n1144), .ZN(n1672) );
  NAND2_X1 U1081 ( .A1(add_r23[13]), .A2(n2038), .ZN(n1144) );
  OAI21_X1 U1082 ( .B1(n2120), .B2(n67), .A(n1464), .ZN(n1992) );
  NAND2_X1 U1083 ( .A1(add_r3[13]), .A2(n2049), .ZN(n1464) );
  OAI21_X1 U1084 ( .B1(n2119), .B2(n83), .A(n1448), .ZN(n1976) );
  NAND2_X1 U1085 ( .A1(add_r4[13]), .A2(n2051), .ZN(n1448) );
  OAI21_X1 U1086 ( .B1(n2104), .B2(n115), .A(n1416), .ZN(n1944) );
  NAND2_X1 U1087 ( .A1(add_r6[13]), .A2(n2053), .ZN(n1416) );
  OAI21_X1 U1088 ( .B1(n2110), .B2(n99), .A(n1432), .ZN(n1960) );
  NAND2_X1 U1089 ( .A1(add_r5[13]), .A2(n2052), .ZN(n1432) );
  OAI21_X1 U1090 ( .B1(n2094), .B2(n468), .A(n1063), .ZN(n1591) );
  NAND2_X1 U1091 ( .A1(add_r28[12]), .A2(n2074), .ZN(n1063) );
  OAI21_X1 U1092 ( .B1(n2108), .B2(n292), .A(n1239), .ZN(n1767) );
  NAND2_X1 U1093 ( .A1(add_r17[12]), .A2(n2039), .ZN(n1239) );
  OAI21_X1 U1094 ( .B1(n2103), .B2(n356), .A(n1175), .ZN(n1703) );
  NAND2_X1 U1095 ( .A1(add_r21[12]), .A2(n2045), .ZN(n1175) );
  OAI21_X1 U1096 ( .B1(n2106), .B2(n324), .A(n1207), .ZN(n1735) );
  NAND2_X1 U1097 ( .A1(add_r19[12]), .A2(n2037), .ZN(n1207) );
  OAI21_X1 U1098 ( .B1(n2107), .B2(n308), .A(n1223), .ZN(n1751) );
  NAND2_X1 U1099 ( .A1(add_r18[12]), .A2(n2041), .ZN(n1223) );
  OAI21_X1 U1100 ( .B1(n2092), .B2(n260), .A(n1271), .ZN(n1799) );
  NAND2_X1 U1101 ( .A1(add_r15[12]), .A2(n2065), .ZN(n1271) );
  OAI21_X1 U1102 ( .B1(n2102), .B2(n372), .A(n1159), .ZN(n1687) );
  NAND2_X1 U1103 ( .A1(add_r22[12]), .A2(n2042), .ZN(n1159) );
  OAI21_X1 U1104 ( .B1(n2097), .B2(n436), .A(n1095), .ZN(n1623) );
  NAND2_X1 U1105 ( .A1(add_r26[12]), .A2(n2071), .ZN(n1095) );
  OAI21_X1 U1106 ( .B1(n2099), .B2(n404), .A(n1127), .ZN(n1655) );
  NAND2_X1 U1107 ( .A1(add_r24[12]), .A2(n2068), .ZN(n1127) );
  OAI21_X1 U1108 ( .B1(n2105), .B2(n340), .A(n1191), .ZN(n1719) );
  NAND2_X1 U1109 ( .A1(add_r20[12]), .A2(n2044), .ZN(n1191) );
  OAI21_X1 U1110 ( .B1(n2109), .B2(n276), .A(n1255), .ZN(n1783) );
  NAND2_X1 U1111 ( .A1(add_r16[12]), .A2(n2046), .ZN(n1255) );
  OAI21_X1 U1112 ( .B1(n2095), .B2(n452), .A(n1079), .ZN(n1607) );
  NAND2_X1 U1113 ( .A1(add_r27[12]), .A2(n2072), .ZN(n1079) );
  OAI21_X1 U1114 ( .B1(n2093), .B2(n484), .A(n1047), .ZN(n1575) );
  NAND2_X1 U1115 ( .A1(add_r29[12]), .A2(n2075), .ZN(n1047) );
  OAI21_X1 U1116 ( .B1(n2098), .B2(n420), .A(n1111), .ZN(n1639) );
  NAND2_X1 U1117 ( .A1(add_r25[12]), .A2(n2070), .ZN(n1111) );
  OAI21_X1 U1118 ( .B1(n2101), .B2(n388), .A(n1143), .ZN(n1671) );
  NAND2_X1 U1119 ( .A1(add_r23[12]), .A2(n2037), .ZN(n1143) );
  OAI21_X1 U1120 ( .B1(n2120), .B2(n68), .A(n1463), .ZN(n1991) );
  NAND2_X1 U1121 ( .A1(add_r3[12]), .A2(n2049), .ZN(n1463) );
  OAI21_X1 U1122 ( .B1(n2119), .B2(n84), .A(n1447), .ZN(n1975) );
  NAND2_X1 U1123 ( .A1(add_r4[12]), .A2(n2051), .ZN(n1447) );
  OAI21_X1 U1124 ( .B1(n2096), .B2(n116), .A(n1415), .ZN(n1943) );
  NAND2_X1 U1125 ( .A1(add_r6[12]), .A2(n2053), .ZN(n1415) );
  OAI21_X1 U1126 ( .B1(n2113), .B2(n100), .A(n1431), .ZN(n1959) );
  NAND2_X1 U1127 ( .A1(add_r5[12]), .A2(n2052), .ZN(n1431) );
  OAI21_X1 U1128 ( .B1(n2093), .B2(n480), .A(n1051), .ZN(n1579) );
  NAND2_X1 U1129 ( .A1(add_r28[0]), .A2(n2075), .ZN(n1051) );
  OAI21_X1 U1130 ( .B1(n2093), .B2(n479), .A(n1052), .ZN(n1580) );
  NAND2_X1 U1131 ( .A1(add_r28[1]), .A2(n2075), .ZN(n1052) );
  OAI21_X1 U1132 ( .B1(n2093), .B2(n478), .A(n1053), .ZN(n1581) );
  NAND2_X1 U1133 ( .A1(add_r28[2]), .A2(n2075), .ZN(n1053) );
  OAI21_X1 U1134 ( .B1(n2093), .B2(n477), .A(n1054), .ZN(n1582) );
  NAND2_X1 U1135 ( .A1(add_r28[3]), .A2(n2075), .ZN(n1054) );
  OAI21_X1 U1136 ( .B1(n2093), .B2(n476), .A(n1055), .ZN(n1583) );
  NAND2_X1 U1137 ( .A1(add_r28[4]), .A2(n2074), .ZN(n1055) );
  OAI21_X1 U1138 ( .B1(n2093), .B2(n475), .A(n1056), .ZN(n1584) );
  NAND2_X1 U1139 ( .A1(add_r28[5]), .A2(n2074), .ZN(n1056) );
  OAI21_X1 U1140 ( .B1(n2093), .B2(n474), .A(n1057), .ZN(n1585) );
  NAND2_X1 U1141 ( .A1(add_r28[6]), .A2(n2074), .ZN(n1057) );
  OAI21_X1 U1142 ( .B1(n2093), .B2(n473), .A(n1058), .ZN(n1586) );
  NAND2_X1 U1143 ( .A1(add_r28[7]), .A2(n2074), .ZN(n1058) );
  OAI21_X1 U1144 ( .B1(n2094), .B2(n472), .A(n1059), .ZN(n1587) );
  NAND2_X1 U1145 ( .A1(add_r28[8]), .A2(n2074), .ZN(n1059) );
  OAI21_X1 U1146 ( .B1(n2094), .B2(n471), .A(n1060), .ZN(n1588) );
  NAND2_X1 U1147 ( .A1(add_r28[9]), .A2(n2074), .ZN(n1060) );
  OAI21_X1 U1148 ( .B1(n2094), .B2(n464), .A(n1067), .ZN(n1595) );
  NAND2_X1 U1149 ( .A1(add_r27[0]), .A2(n2073), .ZN(n1067) );
  OAI21_X1 U1150 ( .B1(n2094), .B2(n463), .A(n1068), .ZN(n1596) );
  NAND2_X1 U1151 ( .A1(add_r27[1]), .A2(n2073), .ZN(n1068) );
  OAI21_X1 U1152 ( .B1(n2094), .B2(n462), .A(n1069), .ZN(n1597) );
  NAND2_X1 U1153 ( .A1(add_r27[2]), .A2(n2073), .ZN(n1069) );
  OAI21_X1 U1154 ( .B1(n2094), .B2(n461), .A(n1070), .ZN(n1598) );
  NAND2_X1 U1155 ( .A1(add_r27[3]), .A2(n2073), .ZN(n1070) );
  OAI21_X1 U1156 ( .B1(n2095), .B2(n460), .A(n1071), .ZN(n1599) );
  NAND2_X1 U1157 ( .A1(add_r27[4]), .A2(n2073), .ZN(n1071) );
  OAI21_X1 U1158 ( .B1(n2095), .B2(n459), .A(n1072), .ZN(n1600) );
  NAND2_X1 U1159 ( .A1(add_r27[5]), .A2(n2073), .ZN(n1072) );
  OAI21_X1 U1160 ( .B1(n2095), .B2(n458), .A(n1073), .ZN(n1601) );
  NAND2_X1 U1161 ( .A1(add_r27[6]), .A2(n2073), .ZN(n1073) );
  OAI21_X1 U1162 ( .B1(n2095), .B2(n457), .A(n1074), .ZN(n1602) );
  NAND2_X1 U1163 ( .A1(add_r27[7]), .A2(n2073), .ZN(n1074) );
  OAI21_X1 U1164 ( .B1(n2095), .B2(n456), .A(n1075), .ZN(n1603) );
  NAND2_X1 U1165 ( .A1(add_r27[8]), .A2(n2073), .ZN(n1075) );
  OAI21_X1 U1166 ( .B1(n2095), .B2(n455), .A(n1076), .ZN(n1604) );
  NAND2_X1 U1167 ( .A1(add_r27[9]), .A2(n2073), .ZN(n1076) );
  OAI21_X1 U1168 ( .B1(n2097), .B2(n432), .A(n1099), .ZN(n1627) );
  NAND2_X1 U1169 ( .A1(add_r25[0]), .A2(n2071), .ZN(n1099) );
  OAI21_X1 U1170 ( .B1(n2097), .B2(n431), .A(n1100), .ZN(n1628) );
  NAND2_X1 U1171 ( .A1(add_r25[1]), .A2(n2071), .ZN(n1100) );
  OAI21_X1 U1172 ( .B1(n2097), .B2(n430), .A(n1101), .ZN(n1629) );
  NAND2_X1 U1173 ( .A1(add_r25[2]), .A2(n2071), .ZN(n1101) );
  OAI21_X1 U1174 ( .B1(n2097), .B2(n429), .A(n1102), .ZN(n1630) );
  NAND2_X1 U1175 ( .A1(add_r25[3]), .A2(n2071), .ZN(n1102) );
  OAI21_X1 U1176 ( .B1(n2097), .B2(n428), .A(n1103), .ZN(n1631) );
  NAND2_X1 U1177 ( .A1(add_r25[4]), .A2(n2070), .ZN(n1103) );
  OAI21_X1 U1178 ( .B1(n2097), .B2(n427), .A(n1104), .ZN(n1632) );
  NAND2_X1 U1179 ( .A1(add_r25[5]), .A2(n2070), .ZN(n1104) );
  OAI21_X1 U1180 ( .B1(n2097), .B2(n426), .A(n1105), .ZN(n1633) );
  NAND2_X1 U1181 ( .A1(add_r25[6]), .A2(n2070), .ZN(n1105) );
  OAI21_X1 U1182 ( .B1(n2097), .B2(n425), .A(n1106), .ZN(n1634) );
  NAND2_X1 U1183 ( .A1(add_r25[7]), .A2(n2070), .ZN(n1106) );
  OAI21_X1 U1184 ( .B1(n2098), .B2(n424), .A(n1107), .ZN(n1635) );
  NAND2_X1 U1185 ( .A1(add_r25[8]), .A2(n2070), .ZN(n1107) );
  OAI21_X1 U1186 ( .B1(n2098), .B2(n423), .A(n1108), .ZN(n1636) );
  NAND2_X1 U1187 ( .A1(add_r25[9]), .A2(n2070), .ZN(n1108) );
  OAI21_X1 U1188 ( .B1(n2098), .B2(n416), .A(n1115), .ZN(n1643) );
  NAND2_X1 U1189 ( .A1(add_r24[0]), .A2(n2069), .ZN(n1115) );
  OAI21_X1 U1190 ( .B1(n2098), .B2(n415), .A(n1116), .ZN(n1644) );
  NAND2_X1 U1191 ( .A1(add_r24[1]), .A2(n2069), .ZN(n1116) );
  OAI21_X1 U1192 ( .B1(n2098), .B2(n414), .A(n1117), .ZN(n1645) );
  NAND2_X1 U1193 ( .A1(add_r24[2]), .A2(n2069), .ZN(n1117) );
  OAI21_X1 U1194 ( .B1(n2098), .B2(n413), .A(n1118), .ZN(n1646) );
  NAND2_X1 U1195 ( .A1(add_r24[3]), .A2(n2069), .ZN(n1118) );
  OAI21_X1 U1196 ( .B1(n2099), .B2(n412), .A(n1119), .ZN(n1647) );
  NAND2_X1 U1197 ( .A1(add_r24[4]), .A2(n2069), .ZN(n1119) );
  OAI21_X1 U1198 ( .B1(n2099), .B2(n411), .A(n1120), .ZN(n1648) );
  NAND2_X1 U1199 ( .A1(add_r24[5]), .A2(n2069), .ZN(n1120) );
  OAI21_X1 U1200 ( .B1(n2099), .B2(n410), .A(n1121), .ZN(n1649) );
  NAND2_X1 U1201 ( .A1(add_r24[6]), .A2(n2069), .ZN(n1121) );
  OAI21_X1 U1202 ( .B1(n2099), .B2(n409), .A(n1122), .ZN(n1650) );
  NAND2_X1 U1203 ( .A1(add_r24[7]), .A2(n2069), .ZN(n1122) );
  OAI21_X1 U1204 ( .B1(n2099), .B2(n408), .A(n1123), .ZN(n1651) );
  NAND2_X1 U1205 ( .A1(add_r24[8]), .A2(n2069), .ZN(n1123) );
  OAI21_X1 U1206 ( .B1(n2099), .B2(n407), .A(n1124), .ZN(n1652) );
  NAND2_X1 U1207 ( .A1(add_r24[9]), .A2(n2069), .ZN(n1124) );
  OAI21_X1 U1208 ( .B1(n2101), .B2(n384), .A(n1147), .ZN(n1675) );
  NAND2_X1 U1209 ( .A1(add_r22[0]), .A2(n2036), .ZN(n1147) );
  OAI21_X1 U1210 ( .B1(n2101), .B2(n383), .A(n1148), .ZN(n1676) );
  NAND2_X1 U1211 ( .A1(add_r22[1]), .A2(n2046), .ZN(n1148) );
  OAI21_X1 U1212 ( .B1(n2101), .B2(n382), .A(n1149), .ZN(n1677) );
  NAND2_X1 U1213 ( .A1(add_r22[2]), .A2(n2080), .ZN(n1149) );
  OAI21_X1 U1214 ( .B1(n2101), .B2(n381), .A(n1150), .ZN(n1678) );
  NAND2_X1 U1215 ( .A1(add_r22[3]), .A2(n2040), .ZN(n1150) );
  OAI21_X1 U1216 ( .B1(n2101), .B2(n380), .A(n1151), .ZN(n1679) );
  NAND2_X1 U1217 ( .A1(add_r22[4]), .A2(n2039), .ZN(n1151) );
  OAI21_X1 U1218 ( .B1(n2101), .B2(n379), .A(n1152), .ZN(n1680) );
  NAND2_X1 U1219 ( .A1(add_r22[5]), .A2(n2036), .ZN(n1152) );
  OAI21_X1 U1220 ( .B1(n2101), .B2(n378), .A(n1153), .ZN(n1681) );
  NAND2_X1 U1221 ( .A1(add_r22[6]), .A2(n2043), .ZN(n1153) );
  OAI21_X1 U1222 ( .B1(n2101), .B2(n377), .A(n1154), .ZN(n1682) );
  NAND2_X1 U1223 ( .A1(add_r22[7]), .A2(n2044), .ZN(n1154) );
  OAI21_X1 U1224 ( .B1(n2102), .B2(n376), .A(n1155), .ZN(n1683) );
  NAND2_X1 U1225 ( .A1(add_r22[8]), .A2(n2038), .ZN(n1155) );
  OAI21_X1 U1226 ( .B1(n2102), .B2(n375), .A(n1156), .ZN(n1684) );
  NAND2_X1 U1227 ( .A1(add_r22[9]), .A2(n2037), .ZN(n1156) );
  OAI21_X1 U1228 ( .B1(n2102), .B2(n368), .A(n1163), .ZN(n1691) );
  NAND2_X1 U1229 ( .A1(add_r21[0]), .A2(n2067), .ZN(n1163) );
  OAI21_X1 U1230 ( .B1(n2102), .B2(n367), .A(n1164), .ZN(n1692) );
  NAND2_X1 U1231 ( .A1(add_r21[1]), .A2(n2067), .ZN(n1164) );
  OAI21_X1 U1232 ( .B1(n2102), .B2(n366), .A(n1165), .ZN(n1693) );
  NAND2_X1 U1233 ( .A1(add_r21[2]), .A2(n2067), .ZN(n1165) );
  OAI21_X1 U1234 ( .B1(n2102), .B2(n365), .A(n1166), .ZN(n1694) );
  NAND2_X1 U1235 ( .A1(add_r21[3]), .A2(n2067), .ZN(n1166) );
  OAI21_X1 U1236 ( .B1(n2103), .B2(n364), .A(n1167), .ZN(n1695) );
  NAND2_X1 U1237 ( .A1(add_r21[4]), .A2(n2067), .ZN(n1167) );
  OAI21_X1 U1238 ( .B1(n2103), .B2(n363), .A(n1168), .ZN(n1696) );
  NAND2_X1 U1239 ( .A1(add_r21[5]), .A2(n2067), .ZN(n1168) );
  OAI21_X1 U1240 ( .B1(n2103), .B2(n362), .A(n1169), .ZN(n1697) );
  NAND2_X1 U1241 ( .A1(add_r21[6]), .A2(n2067), .ZN(n1169) );
  OAI21_X1 U1242 ( .B1(n2103), .B2(n361), .A(n1170), .ZN(n1698) );
  NAND2_X1 U1243 ( .A1(add_r21[7]), .A2(n2067), .ZN(n1170) );
  OAI21_X1 U1244 ( .B1(n2103), .B2(n360), .A(n1171), .ZN(n1699) );
  NAND2_X1 U1245 ( .A1(add_r21[8]), .A2(n2067), .ZN(n1171) );
  OAI21_X1 U1246 ( .B1(n2103), .B2(n359), .A(n1172), .ZN(n1700) );
  NAND2_X1 U1247 ( .A1(add_r21[9]), .A2(n2067), .ZN(n1172) );
  OAI21_X1 U1248 ( .B1(n2105), .B2(n336), .A(n1195), .ZN(n1723) );
  NAND2_X1 U1249 ( .A1(add_r19[0]), .A2(n2046), .ZN(n1195) );
  OAI21_X1 U1250 ( .B1(n2105), .B2(n335), .A(n1196), .ZN(n1724) );
  NAND2_X1 U1251 ( .A1(add_r19[1]), .A2(n2040), .ZN(n1196) );
  OAI21_X1 U1252 ( .B1(n2105), .B2(n334), .A(n1197), .ZN(n1725) );
  NAND2_X1 U1253 ( .A1(add_r19[2]), .A2(n2044), .ZN(n1197) );
  OAI21_X1 U1254 ( .B1(n2105), .B2(n333), .A(n1198), .ZN(n1726) );
  NAND2_X1 U1255 ( .A1(add_r19[3]), .A2(n2039), .ZN(n1198) );
  OAI21_X1 U1256 ( .B1(n2105), .B2(n332), .A(n1199), .ZN(n1727) );
  NAND2_X1 U1257 ( .A1(add_r19[4]), .A2(n2036), .ZN(n1199) );
  OAI21_X1 U1258 ( .B1(n2105), .B2(n330), .A(n1201), .ZN(n1729) );
  NAND2_X1 U1259 ( .A1(add_r19[6]), .A2(n2046), .ZN(n1201) );
  OAI21_X1 U1260 ( .B1(n2105), .B2(n329), .A(n1202), .ZN(n1730) );
  NAND2_X1 U1261 ( .A1(add_r19[7]), .A2(n2044), .ZN(n1202) );
  OAI21_X1 U1262 ( .B1(n2106), .B2(n328), .A(n1203), .ZN(n1731) );
  NAND2_X1 U1263 ( .A1(add_r19[8]), .A2(n985), .ZN(n1203) );
  OAI21_X1 U1264 ( .B1(n2106), .B2(n327), .A(n1204), .ZN(n1732) );
  NAND2_X1 U1265 ( .A1(add_r19[9]), .A2(n2045), .ZN(n1204) );
  OAI21_X1 U1266 ( .B1(n2106), .B2(n320), .A(n1211), .ZN(n1739) );
  NAND2_X1 U1267 ( .A1(add_r18[0]), .A2(n2040), .ZN(n1211) );
  OAI21_X1 U1268 ( .B1(n2106), .B2(n319), .A(n1212), .ZN(n1740) );
  NAND2_X1 U1269 ( .A1(add_r18[1]), .A2(n2039), .ZN(n1212) );
  OAI21_X1 U1270 ( .B1(n2106), .B2(n318), .A(n1213), .ZN(n1741) );
  NAND2_X1 U1271 ( .A1(add_r18[2]), .A2(n2045), .ZN(n1213) );
  OAI21_X1 U1272 ( .B1(n2106), .B2(n317), .A(n1214), .ZN(n1742) );
  NAND2_X1 U1273 ( .A1(add_r18[3]), .A2(n2044), .ZN(n1214) );
  OAI21_X1 U1274 ( .B1(n2107), .B2(n316), .A(n1215), .ZN(n1743) );
  NAND2_X1 U1275 ( .A1(add_r18[4]), .A2(n2038), .ZN(n1215) );
  OAI21_X1 U1276 ( .B1(n2107), .B2(n314), .A(n1217), .ZN(n1745) );
  NAND2_X1 U1277 ( .A1(add_r18[6]), .A2(n2037), .ZN(n1217) );
  OAI21_X1 U1278 ( .B1(n2107), .B2(n313), .A(n1218), .ZN(n1746) );
  NAND2_X1 U1279 ( .A1(add_r18[7]), .A2(n2036), .ZN(n1218) );
  OAI21_X1 U1280 ( .B1(n2107), .B2(n312), .A(n1219), .ZN(n1747) );
  NAND2_X1 U1281 ( .A1(add_r18[8]), .A2(n985), .ZN(n1219) );
  OAI21_X1 U1282 ( .B1(n2107), .B2(n311), .A(n1220), .ZN(n1748) );
  NAND2_X1 U1283 ( .A1(add_r18[9]), .A2(n985), .ZN(n1220) );
  OAI21_X1 U1284 ( .B1(n2108), .B2(n288), .A(n1243), .ZN(n1771) );
  NAND2_X1 U1285 ( .A1(add_r16[0]), .A2(n985), .ZN(n1243) );
  OAI21_X1 U1286 ( .B1(n2108), .B2(n287), .A(n1244), .ZN(n1772) );
  NAND2_X1 U1287 ( .A1(add_r16[1]), .A2(n2038), .ZN(n1244) );
  OAI21_X1 U1288 ( .B1(n2108), .B2(n286), .A(n1245), .ZN(n1773) );
  NAND2_X1 U1289 ( .A1(add_r16[2]), .A2(n2037), .ZN(n1245) );
  OAI21_X1 U1290 ( .B1(n2108), .B2(n285), .A(n1246), .ZN(n1774) );
  NAND2_X1 U1291 ( .A1(add_r16[3]), .A2(n2036), .ZN(n1246) );
  OAI21_X1 U1292 ( .B1(n2108), .B2(n284), .A(n1247), .ZN(n1775) );
  NAND2_X1 U1293 ( .A1(add_r16[4]), .A2(n2080), .ZN(n1247) );
  OAI21_X1 U1294 ( .B1(n2108), .B2(n283), .A(n1248), .ZN(n1776) );
  NAND2_X1 U1295 ( .A1(add_r16[5]), .A2(n2040), .ZN(n1248) );
  OAI21_X1 U1296 ( .B1(n2108), .B2(n282), .A(n1249), .ZN(n1777) );
  NAND2_X1 U1297 ( .A1(add_r16[6]), .A2(n985), .ZN(n1249) );
  OAI21_X1 U1298 ( .B1(n2108), .B2(n281), .A(n1250), .ZN(n1778) );
  NAND2_X1 U1299 ( .A1(add_r16[7]), .A2(n2045), .ZN(n1250) );
  OAI21_X1 U1300 ( .B1(n2109), .B2(n280), .A(n1251), .ZN(n1779) );
  NAND2_X1 U1301 ( .A1(add_r16[8]), .A2(n2041), .ZN(n1251) );
  OAI21_X1 U1302 ( .B1(n2109), .B2(n279), .A(n1252), .ZN(n1780) );
  NAND2_X1 U1303 ( .A1(add_r16[9]), .A2(n2042), .ZN(n1252) );
  OAI21_X1 U1304 ( .B1(n2109), .B2(n272), .A(n1259), .ZN(n1787) );
  NAND2_X1 U1305 ( .A1(add_r15[0]), .A2(n2066), .ZN(n1259) );
  OAI21_X1 U1306 ( .B1(n2109), .B2(n271), .A(n1260), .ZN(n1788) );
  NAND2_X1 U1307 ( .A1(add_r15[1]), .A2(n2066), .ZN(n1260) );
  OAI21_X1 U1308 ( .B1(n2109), .B2(n270), .A(n1261), .ZN(n1789) );
  NAND2_X1 U1309 ( .A1(add_r15[2]), .A2(n2066), .ZN(n1261) );
  OAI21_X1 U1310 ( .B1(n2109), .B2(n269), .A(n1262), .ZN(n1790) );
  NAND2_X1 U1311 ( .A1(add_r15[3]), .A2(n2066), .ZN(n1262) );
  OAI21_X1 U1312 ( .B1(n2088), .B2(n268), .A(n1263), .ZN(n1791) );
  NAND2_X1 U1313 ( .A1(add_r15[4]), .A2(n2066), .ZN(n1263) );
  OAI21_X1 U1314 ( .B1(n2100), .B2(n266), .A(n1265), .ZN(n1793) );
  NAND2_X1 U1315 ( .A1(add_r15[6]), .A2(n2066), .ZN(n1265) );
  OAI21_X1 U1316 ( .B1(n2113), .B2(n265), .A(n1266), .ZN(n1794) );
  NAND2_X1 U1317 ( .A1(add_r15[7]), .A2(n2066), .ZN(n1266) );
  OAI21_X1 U1318 ( .B1(n2111), .B2(n264), .A(n1267), .ZN(n1795) );
  NAND2_X1 U1319 ( .A1(add_r15[8]), .A2(n2066), .ZN(n1267) );
  OAI21_X1 U1320 ( .B1(n2110), .B2(n263), .A(n1268), .ZN(n1796) );
  NAND2_X1 U1321 ( .A1(add_r15[9]), .A2(n2066), .ZN(n1268) );
  OAI21_X1 U1322 ( .B1(n2100), .B2(n124), .A(n1407), .ZN(n1935) );
  NAND2_X1 U1323 ( .A1(add_r6[4]), .A2(n2054), .ZN(n1407) );
  OAI21_X1 U1324 ( .B1(n2088), .B2(n123), .A(n1408), .ZN(n1936) );
  NAND2_X1 U1325 ( .A1(add_r6[5]), .A2(n2054), .ZN(n1408) );
  OAI21_X1 U1326 ( .B1(n2092), .B2(n122), .A(n1409), .ZN(n1937) );
  NAND2_X1 U1327 ( .A1(add_r6[6]), .A2(n2054), .ZN(n1409) );
  OAI21_X1 U1328 ( .B1(n2104), .B2(n121), .A(n1410), .ZN(n1938) );
  NAND2_X1 U1329 ( .A1(add_r6[7]), .A2(n2054), .ZN(n1410) );
  OAI21_X1 U1330 ( .B1(n2111), .B2(n120), .A(n1411), .ZN(n1939) );
  NAND2_X1 U1331 ( .A1(add_r6[8]), .A2(n2054), .ZN(n1411) );
  OAI21_X1 U1332 ( .B1(n2110), .B2(n119), .A(n1412), .ZN(n1940) );
  NAND2_X1 U1333 ( .A1(add_r6[9]), .A2(n2054), .ZN(n1412) );
  OAI21_X1 U1334 ( .B1(n2096), .B2(n96), .A(n1435), .ZN(n1963) );
  NAND2_X1 U1335 ( .A1(add_r4[0]), .A2(n2052), .ZN(n1435) );
  OAI21_X1 U1336 ( .B1(n2100), .B2(n95), .A(n1436), .ZN(n1964) );
  NAND2_X1 U1337 ( .A1(add_r4[1]), .A2(n2052), .ZN(n1436) );
  OAI21_X1 U1338 ( .B1(n2088), .B2(n94), .A(n1437), .ZN(n1965) );
  NAND2_X1 U1339 ( .A1(add_r4[2]), .A2(n2052), .ZN(n1437) );
  OAI21_X1 U1340 ( .B1(n2092), .B2(n93), .A(n1438), .ZN(n1966) );
  NAND2_X1 U1341 ( .A1(add_r4[3]), .A2(n2052), .ZN(n1438) );
  OAI21_X1 U1342 ( .B1(n2104), .B2(n92), .A(n1439), .ZN(n1967) );
  NAND2_X1 U1343 ( .A1(add_r4[4]), .A2(n2051), .ZN(n1439) );
  OAI21_X1 U1344 ( .B1(n2113), .B2(n91), .A(n1440), .ZN(n1968) );
  NAND2_X1 U1345 ( .A1(add_r4[5]), .A2(n2051), .ZN(n1440) );
  OAI21_X1 U1346 ( .B1(n2110), .B2(n90), .A(n1441), .ZN(n1969) );
  NAND2_X1 U1347 ( .A1(add_r4[6]), .A2(n2051), .ZN(n1441) );
  OAI21_X1 U1348 ( .B1(n2113), .B2(n89), .A(n1442), .ZN(n1970) );
  NAND2_X1 U1349 ( .A1(add_r4[7]), .A2(n2051), .ZN(n1442) );
  OAI21_X1 U1350 ( .B1(n2119), .B2(n88), .A(n1443), .ZN(n1971) );
  NAND2_X1 U1351 ( .A1(add_r4[8]), .A2(n2051), .ZN(n1443) );
  OAI21_X1 U1352 ( .B1(n2119), .B2(n87), .A(n1444), .ZN(n1972) );
  NAND2_X1 U1353 ( .A1(add_r4[9]), .A2(n2051), .ZN(n1444) );
  OAI21_X1 U1354 ( .B1(n2119), .B2(n80), .A(n1451), .ZN(n1979) );
  NAND2_X1 U1355 ( .A1(add_r3[0]), .A2(n2050), .ZN(n1451) );
  OAI21_X1 U1356 ( .B1(n2119), .B2(n79), .A(n1452), .ZN(n1980) );
  NAND2_X1 U1357 ( .A1(add_r3[1]), .A2(n2050), .ZN(n1452) );
  OAI21_X1 U1358 ( .B1(n2119), .B2(n78), .A(n1453), .ZN(n1981) );
  NAND2_X1 U1359 ( .A1(add_r3[2]), .A2(n2050), .ZN(n1453) );
  OAI21_X1 U1360 ( .B1(n2119), .B2(n77), .A(n1454), .ZN(n1982) );
  NAND2_X1 U1361 ( .A1(add_r3[3]), .A2(n2050), .ZN(n1454) );
  OAI21_X1 U1362 ( .B1(n2120), .B2(n76), .A(n1455), .ZN(n1983) );
  NAND2_X1 U1363 ( .A1(add_r3[4]), .A2(n2050), .ZN(n1455) );
  OAI21_X1 U1364 ( .B1(n2120), .B2(n75), .A(n1456), .ZN(n1984) );
  NAND2_X1 U1365 ( .A1(add_r3[5]), .A2(n2050), .ZN(n1456) );
  OAI21_X1 U1366 ( .B1(n2120), .B2(n74), .A(n1457), .ZN(n1985) );
  NAND2_X1 U1367 ( .A1(add_r3[6]), .A2(n2050), .ZN(n1457) );
  OAI21_X1 U1368 ( .B1(n2120), .B2(n73), .A(n1458), .ZN(n1986) );
  NAND2_X1 U1369 ( .A1(add_r3[7]), .A2(n2050), .ZN(n1458) );
  OAI21_X1 U1370 ( .B1(n2120), .B2(n72), .A(n1459), .ZN(n1987) );
  NAND2_X1 U1371 ( .A1(add_r3[8]), .A2(n2050), .ZN(n1459) );
  OAI21_X1 U1372 ( .B1(n2120), .B2(n71), .A(n1460), .ZN(n1988) );
  NAND2_X1 U1373 ( .A1(add_r3[9]), .A2(n2050), .ZN(n1460) );
  OAI21_X1 U1374 ( .B1(n2091), .B2(n502), .A(n1029), .ZN(n1557) );
  NAND2_X1 U1375 ( .A1(add_r30[10]), .A2(n2077), .ZN(n1029) );
  OAI21_X1 U1376 ( .B1(n2091), .B2(n501), .A(n1030), .ZN(n1558) );
  NAND2_X1 U1377 ( .A1(add_r30[11]), .A2(n2077), .ZN(n1030) );
  OAI21_X1 U1378 ( .B1(n2112), .B2(n230), .A(n1301), .ZN(n1829) );
  NAND2_X1 U1379 ( .A1(add_r13[10]), .A2(n2063), .ZN(n1301) );
  OAI21_X1 U1380 ( .B1(n2112), .B2(n229), .A(n1302), .ZN(n1830) );
  NAND2_X1 U1381 ( .A1(add_r13[11]), .A2(n2063), .ZN(n1302) );
  OAI21_X1 U1382 ( .B1(n2106), .B2(n214), .A(n1317), .ZN(n1845) );
  NAND2_X1 U1383 ( .A1(add_r12[10]), .A2(n2062), .ZN(n1317) );
  OAI21_X1 U1384 ( .B1(n2103), .B2(n213), .A(n1318), .ZN(n1846) );
  NAND2_X1 U1385 ( .A1(add_r12[11]), .A2(n2062), .ZN(n1318) );
  OAI21_X1 U1386 ( .B1(n2114), .B2(n182), .A(n1349), .ZN(n1877) );
  NAND2_X1 U1387 ( .A1(add_r10[10]), .A2(n2059), .ZN(n1349) );
  OAI21_X1 U1388 ( .B1(n2114), .B2(n181), .A(n1350), .ZN(n1878) );
  NAND2_X1 U1389 ( .A1(add_r10[11]), .A2(n2059), .ZN(n1350) );
  OAI21_X1 U1390 ( .B1(n2115), .B2(n166), .A(n1365), .ZN(n1893) );
  NAND2_X1 U1391 ( .A1(add_r9[10]), .A2(n2058), .ZN(n1365) );
  OAI21_X1 U1392 ( .B1(n2115), .B2(n165), .A(n1366), .ZN(n1894) );
  NAND2_X1 U1393 ( .A1(add_r9[11]), .A2(n2058), .ZN(n1366) );
  OAI21_X1 U1394 ( .B1(n2115), .B2(n162), .A(n1369), .ZN(n1897) );
  NAND2_X1 U1395 ( .A1(add_r9[14]), .A2(n2057), .ZN(n1369) );
  OAI21_X1 U1396 ( .B1(n2114), .B2(n178), .A(n1353), .ZN(n1881) );
  NAND2_X1 U1397 ( .A1(add_r10[14]), .A2(n2059), .ZN(n1353) );
  OAI21_X1 U1398 ( .B1(n2111), .B2(n242), .A(n1289), .ZN(n1817) );
  NAND2_X1 U1399 ( .A1(add_r14[14]), .A2(n2064), .ZN(n1289) );
  NAND2_X1 U1400 ( .A1(add_r13[14]), .A2(n2063), .ZN(n1305) );
  OAI21_X1 U1401 ( .B1(n2105), .B2(n210), .A(n1321), .ZN(n1849) );
  NAND2_X1 U1402 ( .A1(add_r12[14]), .A2(n2061), .ZN(n1321) );
  NAND2_X1 U1403 ( .A1(add_r30[14]), .A2(n2076), .ZN(n1033) );
  OAI21_X1 U1404 ( .B1(n2089), .B2(n530), .A(n999), .ZN(n1529) );
  NAND2_X1 U1405 ( .A1(add_r32[14]), .A2(n2079), .ZN(n999) );
  OAI21_X1 U1406 ( .B1(n2117), .B2(n146), .A(n1385), .ZN(n1913) );
  NAND2_X1 U1407 ( .A1(add_r8[14]), .A2(n2056), .ZN(n1385) );
  OAI21_X1 U1408 ( .B1(n2115), .B2(n163), .A(n1368), .ZN(n1896) );
  NAND2_X1 U1409 ( .A1(add_r9[13]), .A2(n2057), .ZN(n1368) );
  OAI21_X1 U1410 ( .B1(n2114), .B2(n179), .A(n1352), .ZN(n1880) );
  NAND2_X1 U1411 ( .A1(add_r10[13]), .A2(n2059), .ZN(n1352) );
  OAI21_X1 U1412 ( .B1(n2111), .B2(n243), .A(n1288), .ZN(n1816) );
  NAND2_X1 U1413 ( .A1(add_r14[13]), .A2(n2064), .ZN(n1288) );
  OAI21_X1 U1414 ( .B1(n2112), .B2(n227), .A(n1304), .ZN(n1832) );
  NAND2_X1 U1415 ( .A1(add_r13[13]), .A2(n2063), .ZN(n1304) );
  OAI21_X1 U1416 ( .B1(n2107), .B2(n211), .A(n1320), .ZN(n1848) );
  NAND2_X1 U1417 ( .A1(add_r12[13]), .A2(n2061), .ZN(n1320) );
  OAI21_X1 U1418 ( .B1(n2091), .B2(n499), .A(n1032), .ZN(n1560) );
  NAND2_X1 U1419 ( .A1(add_r30[13]), .A2(n2076), .ZN(n1032) );
  OAI21_X1 U1420 ( .B1(n2089), .B2(n531), .A(n998), .ZN(n1528) );
  NAND2_X1 U1421 ( .A1(add_r32[13]), .A2(n2079), .ZN(n998) );
  OAI21_X1 U1422 ( .B1(n2117), .B2(n147), .A(n1384), .ZN(n1912) );
  NAND2_X1 U1423 ( .A1(add_r8[13]), .A2(n2056), .ZN(n1384) );
  OAI21_X1 U1424 ( .B1(n2115), .B2(n164), .A(n1367), .ZN(n1895) );
  NAND2_X1 U1425 ( .A1(add_r9[12]), .A2(n2057), .ZN(n1367) );
  OAI21_X1 U1426 ( .B1(n2114), .B2(n180), .A(n1351), .ZN(n1879) );
  NAND2_X1 U1427 ( .A1(add_r10[12]), .A2(n2059), .ZN(n1351) );
  OAI21_X1 U1428 ( .B1(n2111), .B2(n244), .A(n1287), .ZN(n1815) );
  NAND2_X1 U1429 ( .A1(add_r14[12]), .A2(n2064), .ZN(n1287) );
  OAI21_X1 U1430 ( .B1(n2112), .B2(n228), .A(n1303), .ZN(n1831) );
  NAND2_X1 U1431 ( .A1(add_r13[12]), .A2(n2063), .ZN(n1303) );
  OAI21_X1 U1432 ( .B1(n2097), .B2(n212), .A(n1319), .ZN(n1847) );
  NAND2_X1 U1433 ( .A1(add_r12[12]), .A2(n2061), .ZN(n1319) );
  OAI21_X1 U1434 ( .B1(n2091), .B2(n500), .A(n1031), .ZN(n1559) );
  NAND2_X1 U1435 ( .A1(add_r30[12]), .A2(n2076), .ZN(n1031) );
  OAI21_X1 U1436 ( .B1(n2089), .B2(n532), .A(n997), .ZN(n1527) );
  NAND2_X1 U1437 ( .A1(add_r32[12]), .A2(n2079), .ZN(n997) );
  OAI21_X1 U1438 ( .B1(n2117), .B2(n148), .A(n1383), .ZN(n1911) );
  NAND2_X1 U1439 ( .A1(add_r8[12]), .A2(n2056), .ZN(n1383) );
  OAI21_X1 U1440 ( .B1(n2089), .B2(n527), .A(n1003), .ZN(n1532) );
  NAND2_X1 U1441 ( .A1(add_r31[1]), .A2(n2079), .ZN(n1003) );
  OAI21_X1 U1442 ( .B1(n2089), .B2(n526), .A(n1004), .ZN(n1533) );
  NAND2_X1 U1443 ( .A1(add_r31[2]), .A2(n2079), .ZN(n1004) );
  OAI21_X1 U1444 ( .B1(n2089), .B2(n525), .A(n1005), .ZN(n1534) );
  NAND2_X1 U1445 ( .A1(add_r31[3]), .A2(n2078), .ZN(n1005) );
  OAI21_X1 U1446 ( .B1(n2089), .B2(n524), .A(n1006), .ZN(n1535) );
  NAND2_X1 U1447 ( .A1(add_r31[4]), .A2(n2078), .ZN(n1006) );
  OAI21_X1 U1448 ( .B1(n2089), .B2(n523), .A(n1007), .ZN(n1536) );
  NAND2_X1 U1449 ( .A1(add_r31[5]), .A2(n2078), .ZN(n1007) );
  OAI21_X1 U1450 ( .B1(n2089), .B2(n522), .A(n1008), .ZN(n1537) );
  NAND2_X1 U1451 ( .A1(add_r31[6]), .A2(n2078), .ZN(n1008) );
  OAI21_X1 U1452 ( .B1(n2089), .B2(n521), .A(n1009), .ZN(n1538) );
  NAND2_X1 U1453 ( .A1(add_r31[7]), .A2(n2078), .ZN(n1009) );
  OAI21_X1 U1454 ( .B1(n2091), .B2(n508), .A(n1023), .ZN(n1551) );
  NAND2_X1 U1455 ( .A1(add_r30[4]), .A2(n2077), .ZN(n1023) );
  OAI21_X1 U1456 ( .B1(n2091), .B2(n507), .A(n1024), .ZN(n1552) );
  NAND2_X1 U1457 ( .A1(add_r30[5]), .A2(n2077), .ZN(n1024) );
  OAI21_X1 U1458 ( .B1(n2091), .B2(n506), .A(n1025), .ZN(n1553) );
  NAND2_X1 U1459 ( .A1(add_r30[6]), .A2(n2077), .ZN(n1025) );
  OAI21_X1 U1460 ( .B1(n2091), .B2(n505), .A(n1026), .ZN(n1554) );
  NAND2_X1 U1461 ( .A1(add_r30[7]), .A2(n2077), .ZN(n1026) );
  OAI21_X1 U1462 ( .B1(n2091), .B2(n504), .A(n1027), .ZN(n1555) );
  NAND2_X1 U1463 ( .A1(add_r30[8]), .A2(n2077), .ZN(n1027) );
  OAI21_X1 U1464 ( .B1(n2091), .B2(n503), .A(n1028), .ZN(n1556) );
  NAND2_X1 U1465 ( .A1(add_r30[9]), .A2(n2077), .ZN(n1028) );
  OAI21_X1 U1466 ( .B1(n2111), .B2(n240), .A(n1291), .ZN(n1819) );
  NAND2_X1 U1467 ( .A1(add_r13[0]), .A2(n2064), .ZN(n1291) );
  OAI21_X1 U1468 ( .B1(n2111), .B2(n239), .A(n1292), .ZN(n1820) );
  NAND2_X1 U1469 ( .A1(add_r13[1]), .A2(n2064), .ZN(n1292) );
  OAI21_X1 U1470 ( .B1(n2111), .B2(n238), .A(n1293), .ZN(n1821) );
  NAND2_X1 U1471 ( .A1(add_r13[2]), .A2(n2064), .ZN(n1293) );
  OAI21_X1 U1472 ( .B1(n2111), .B2(n237), .A(n1294), .ZN(n1822) );
  NAND2_X1 U1473 ( .A1(add_r13[3]), .A2(n2064), .ZN(n1294) );
  OAI21_X1 U1474 ( .B1(n2111), .B2(n236), .A(n1295), .ZN(n1823) );
  NAND2_X1 U1475 ( .A1(add_r13[4]), .A2(n2063), .ZN(n1295) );
  OAI21_X1 U1476 ( .B1(n2111), .B2(n234), .A(n1297), .ZN(n1825) );
  NAND2_X1 U1477 ( .A1(add_r13[6]), .A2(n2063), .ZN(n1297) );
  OAI21_X1 U1478 ( .B1(n2111), .B2(n233), .A(n1298), .ZN(n1826) );
  NAND2_X1 U1479 ( .A1(add_r13[7]), .A2(n2063), .ZN(n1298) );
  OAI21_X1 U1480 ( .B1(n2112), .B2(n232), .A(n1299), .ZN(n1827) );
  NAND2_X1 U1481 ( .A1(add_r13[8]), .A2(n2063), .ZN(n1299) );
  OAI21_X1 U1482 ( .B1(n2112), .B2(n231), .A(n1300), .ZN(n1828) );
  NAND2_X1 U1484 ( .A1(add_r13[9]), .A2(n2063), .ZN(n1300) );
  OAI21_X1 U1485 ( .B1(n2112), .B2(n224), .A(n1307), .ZN(n1835) );
  NAND2_X1 U1486 ( .A1(add_r12[0]), .A2(n2062), .ZN(n1307) );
  OAI21_X1 U1487 ( .B1(n2112), .B2(n223), .A(n1308), .ZN(n1836) );
  NAND2_X1 U1488 ( .A1(add_r12[1]), .A2(n2062), .ZN(n1308) );
  OAI21_X1 U1489 ( .B1(n2112), .B2(n222), .A(n1309), .ZN(n1837) );
  NAND2_X1 U1490 ( .A1(add_r12[2]), .A2(n2062), .ZN(n1309) );
  OAI21_X1 U1491 ( .B1(n2112), .B2(n221), .A(n1310), .ZN(n1838) );
  NAND2_X1 U1492 ( .A1(add_r12[3]), .A2(n2062), .ZN(n1310) );
  OAI21_X1 U1493 ( .B1(n2095), .B2(n220), .A(n1311), .ZN(n1839) );
  NAND2_X1 U1494 ( .A1(add_r12[4]), .A2(n2062), .ZN(n1311) );
  OAI21_X1 U1495 ( .B1(n2093), .B2(n219), .A(n1312), .ZN(n1840) );
  NAND2_X1 U1496 ( .A1(add_r12[5]), .A2(n2062), .ZN(n1312) );
  OAI21_X1 U1497 ( .B1(n2120), .B2(n218), .A(n1313), .ZN(n1841) );
  NAND2_X1 U1498 ( .A1(add_r12[6]), .A2(n2062), .ZN(n1313) );
  OAI21_X1 U1499 ( .B1(n2096), .B2(n217), .A(n1314), .ZN(n1842) );
  NAND2_X1 U1500 ( .A1(add_r12[7]), .A2(n2062), .ZN(n1314) );
  OAI21_X1 U1501 ( .B1(n2106), .B2(n216), .A(n1315), .ZN(n1843) );
  NAND2_X1 U1502 ( .A1(add_r12[8]), .A2(n2062), .ZN(n1315) );
  OAI21_X1 U1503 ( .B1(n2103), .B2(n215), .A(n1316), .ZN(n1844) );
  NAND2_X1 U1504 ( .A1(add_r12[9]), .A2(n2062), .ZN(n1316) );
  OAI21_X1 U1505 ( .B1(n2114), .B2(n184), .A(n1347), .ZN(n1875) );
  NAND2_X1 U1506 ( .A1(add_r10[8]), .A2(n2059), .ZN(n1347) );
  OAI21_X1 U1507 ( .B1(n2114), .B2(n183), .A(n1348), .ZN(n1876) );
  NAND2_X1 U1508 ( .A1(add_r10[9]), .A2(n2059), .ZN(n1348) );
  OAI21_X1 U1509 ( .B1(n2114), .B2(n176), .A(n1355), .ZN(n1883) );
  NAND2_X1 U1510 ( .A1(add_r9[0]), .A2(n2058), .ZN(n1355) );
  OAI21_X1 U1511 ( .B1(n2114), .B2(n175), .A(n1356), .ZN(n1884) );
  NAND2_X1 U1512 ( .A1(add_r9[1]), .A2(n2058), .ZN(n1356) );
  OAI21_X1 U1513 ( .B1(n2114), .B2(n174), .A(n1357), .ZN(n1885) );
  NAND2_X1 U1514 ( .A1(add_r9[2]), .A2(n2058), .ZN(n1357) );
  OAI21_X1 U1515 ( .B1(n2114), .B2(n173), .A(n1358), .ZN(n1886) );
  NAND2_X1 U1516 ( .A1(add_r9[3]), .A2(n2058), .ZN(n1358) );
  OAI21_X1 U1517 ( .B1(n2115), .B2(n172), .A(n1359), .ZN(n1887) );
  NAND2_X1 U1518 ( .A1(add_r9[4]), .A2(n2058), .ZN(n1359) );
  OAI21_X1 U1519 ( .B1(n2115), .B2(n171), .A(n1360), .ZN(n1888) );
  NAND2_X1 U1520 ( .A1(add_r9[5]), .A2(n2058), .ZN(n1360) );
  OAI21_X1 U1521 ( .B1(n2115), .B2(n170), .A(n1361), .ZN(n1889) );
  NAND2_X1 U1522 ( .A1(add_r9[6]), .A2(n2058), .ZN(n1361) );
  OAI21_X1 U1523 ( .B1(n2115), .B2(n169), .A(n1362), .ZN(n1890) );
  NAND2_X1 U1524 ( .A1(add_r9[7]), .A2(n2058), .ZN(n1362) );
  OAI21_X1 U1525 ( .B1(n2115), .B2(n168), .A(n1363), .ZN(n1891) );
  NAND2_X1 U1526 ( .A1(add_r9[8]), .A2(n2058), .ZN(n1363) );
  OAI21_X1 U1527 ( .B1(n2115), .B2(n167), .A(n1364), .ZN(n1892) );
  NAND2_X1 U1528 ( .A1(add_r9[9]), .A2(n2058), .ZN(n1364) );
  OAI21_X1 U1529 ( .B1(n2117), .B2(n144), .A(n1387), .ZN(n1915) );
  NAND2_X1 U1530 ( .A1(add_r7[0]), .A2(n2056), .ZN(n1387) );
  OAI21_X1 U1531 ( .B1(n2117), .B2(n143), .A(n1388), .ZN(n1916) );
  NAND2_X1 U1532 ( .A1(add_r7[1]), .A2(n2056), .ZN(n1388) );
  OAI21_X1 U1533 ( .B1(n2117), .B2(n142), .A(n1389), .ZN(n1917) );
  NAND2_X1 U1534 ( .A1(add_r7[2]), .A2(n2056), .ZN(n1389) );
  OAI21_X1 U1535 ( .B1(n2117), .B2(n141), .A(n1390), .ZN(n1918) );
  NAND2_X1 U1536 ( .A1(add_r7[3]), .A2(n2056), .ZN(n1390) );
  OAI21_X1 U1537 ( .B1(n2117), .B2(n140), .A(n1391), .ZN(n1919) );
  NAND2_X1 U1538 ( .A1(add_r7[4]), .A2(n2055), .ZN(n1391) );
  OAI21_X1 U1539 ( .B1(n2117), .B2(n139), .A(n1392), .ZN(n1920) );
  NAND2_X1 U1540 ( .A1(add_r7[5]), .A2(n2055), .ZN(n1392) );
  OAI21_X1 U1541 ( .B1(n2117), .B2(n138), .A(n1393), .ZN(n1921) );
  NAND2_X1 U1542 ( .A1(add_r7[6]), .A2(n2055), .ZN(n1393) );
  OAI21_X1 U1543 ( .B1(n2117), .B2(n137), .A(n1394), .ZN(n1922) );
  NAND2_X1 U1544 ( .A1(add_r7[7]), .A2(n2055), .ZN(n1394) );
  OAI21_X1 U1545 ( .B1(n2096), .B2(n50), .A(n1481), .ZN(n2009) );
  NAND2_X1 U1546 ( .A1(add_r2[14]), .A2(n2048), .ZN(n1481) );
  OAI21_X1 U1547 ( .B1(n2088), .B2(n51), .A(n1480), .ZN(n2008) );
  NAND2_X1 U1548 ( .A1(add_r2[13]), .A2(n2048), .ZN(n1480) );
  OAI21_X1 U1549 ( .B1(n2092), .B2(n52), .A(n1479), .ZN(n2007) );
  NAND2_X1 U1550 ( .A1(add_r2[12]), .A2(n2048), .ZN(n1479) );
  OAI21_X1 U1551 ( .B1(n2104), .B2(n48), .A(n1483), .ZN(n2011) );
  NAND2_X1 U1552 ( .A1(add_r1[0]), .A2(n2048), .ZN(n1483) );
  OAI21_X1 U1553 ( .B1(n2113), .B2(n47), .A(n1484), .ZN(n2012) );
  NAND2_X1 U1554 ( .A1(add_r1[1]), .A2(n2048), .ZN(n1484) );
  OAI21_X1 U1555 ( .B1(n2110), .B2(n46), .A(n1485), .ZN(n2013) );
  NAND2_X1 U1556 ( .A1(add_r1[2]), .A2(n2048), .ZN(n1485) );
  OAI21_X1 U1557 ( .B1(n2113), .B2(n45), .A(n1486), .ZN(n2014) );
  NAND2_X1 U1558 ( .A1(add_r1[3]), .A2(n2048), .ZN(n1486) );
  OAI21_X1 U1559 ( .B1(n2116), .B2(n44), .A(n1487), .ZN(n2015) );
  NAND2_X1 U1560 ( .A1(add_r1[4]), .A2(n2047), .ZN(n1487) );
  OAI21_X1 U1561 ( .B1(n2100), .B2(n43), .A(n1488), .ZN(n2016) );
  NAND2_X1 U1562 ( .A1(add_r1[5]), .A2(n2047), .ZN(n1488) );
  OAI21_X1 U1563 ( .B1(n2088), .B2(n42), .A(n1489), .ZN(n2017) );
  NAND2_X1 U1564 ( .A1(add_r1[6]), .A2(n2047), .ZN(n1489) );
  OAI21_X1 U1565 ( .B1(n2092), .B2(n41), .A(n1490), .ZN(n2018) );
  NAND2_X1 U1566 ( .A1(add_r1[7]), .A2(n2047), .ZN(n1490) );
  INV_X1 U1567 ( .A(addr_y[3]), .ZN(n2148) );
  OAI21_X1 U1568 ( .B1(n2093), .B2(n38), .A(n1493), .ZN(n2021) );
  NAND2_X1 U1569 ( .A1(add_r1[10]), .A2(n2047), .ZN(n1493) );
  OAI21_X1 U1570 ( .B1(n2099), .B2(n37), .A(n1494), .ZN(n2022) );
  NAND2_X1 U1571 ( .A1(add_r1[11]), .A2(n2047), .ZN(n1494) );
  OAI21_X1 U1572 ( .B1(n2102), .B2(n34), .A(n1497), .ZN(n2025) );
  NAND2_X1 U1573 ( .A1(add_r1[14]), .A2(n2047), .ZN(n1497) );
  OAI21_X1 U1574 ( .B1(n2089), .B2(n35), .A(n1496), .ZN(n2024) );
  NAND2_X1 U1575 ( .A1(add_r1[13]), .A2(n2047), .ZN(n1496) );
  OAI21_X1 U1576 ( .B1(n2111), .B2(n36), .A(n1495), .ZN(n2023) );
  NAND2_X1 U1577 ( .A1(add_r1[12]), .A2(n2047), .ZN(n1495) );
  OAI21_X1 U1578 ( .B1(n2111), .B2(n40), .A(n1491), .ZN(n2019) );
  NAND2_X1 U1579 ( .A1(add_r1[8]), .A2(n2047), .ZN(n1491) );
  OAI21_X1 U1580 ( .B1(n2110), .B2(n39), .A(n1492), .ZN(n2020) );
  NAND2_X1 U1581 ( .A1(add_r1[9]), .A2(n2047), .ZN(n1492) );
  INV_X1 U1582 ( .A(clear_acc), .ZN(n2170) );
  NAND2_X1 U1583 ( .A1(f24[0]), .A2(n2167), .ZN(n935) );
  NAND2_X1 U1584 ( .A1(f24[1]), .A2(n2167), .ZN(n911) );
  NAND2_X1 U1585 ( .A1(f24[2]), .A2(n2167), .ZN(n889) );
  NAND2_X1 U1586 ( .A1(f24[3]), .A2(n2167), .ZN(n867) );
  NAND2_X1 U1587 ( .A1(f24[4]), .A2(n2167), .ZN(n845) );
  NAND2_X1 U1588 ( .A1(f24[5]), .A2(n2167), .ZN(n823) );
  NAND2_X1 U1589 ( .A1(f24[6]), .A2(n2167), .ZN(n801) );
  NAND2_X1 U1590 ( .A1(f24[7]), .A2(n2167), .ZN(n779) );
  NAND2_X1 U1591 ( .A1(f24[8]), .A2(n2167), .ZN(n757) );
  NAND2_X1 U1592 ( .A1(f24[9]), .A2(n2167), .ZN(n735) );
  NAND2_X1 U1593 ( .A1(f24[10]), .A2(n2167), .ZN(n713) );
  NAND2_X1 U1594 ( .A1(f24[11]), .A2(n2167), .ZN(n691) );
  NAND2_X1 U1595 ( .A1(f24[12]), .A2(n2167), .ZN(n669) );
  NAND2_X1 U1596 ( .A1(f24[13]), .A2(n2167), .ZN(n647) );
  NAND2_X1 U1597 ( .A1(f24[14]), .A2(n2167), .ZN(n625) );
  NAND2_X1 U1598 ( .A1(f24[15]), .A2(n2167), .ZN(n579) );
  OAI21_X1 U1599 ( .B1(n2107), .B2(n315), .A(n1216), .ZN(n1744) );
  NAND2_X1 U1600 ( .A1(add_r18[5]), .A2(n985), .ZN(n1216) );
  OAI21_X1 U1601 ( .B1(n2110), .B2(n267), .A(n1264), .ZN(n1792) );
  NAND2_X1 U1602 ( .A1(add_r15[5]), .A2(n2066), .ZN(n1264) );
  OAI21_X1 U1603 ( .B1(n2105), .B2(n331), .A(n1200), .ZN(n1728) );
  NAND2_X1 U1604 ( .A1(add_r19[5]), .A2(n2043), .ZN(n1200) );
  OAI21_X1 U1605 ( .B1(n2110), .B2(n251), .A(n1280), .ZN(n1808) );
  NAND2_X1 U1606 ( .A1(add_r14[5]), .A2(n2065), .ZN(n1280) );
  OAI21_X1 U1607 ( .B1(n2111), .B2(n235), .A(n1296), .ZN(n1824) );
  NAND2_X1 U1608 ( .A1(add_r13[5]), .A2(n2063), .ZN(n1296) );
  OAI21_X1 U1609 ( .B1(n2113), .B2(n203), .A(n1328), .ZN(n1856) );
  NAND2_X1 U1610 ( .A1(add_r11[5]), .A2(n2061), .ZN(n1328) );
  NAND2_X1 U1611 ( .A1(clc1), .A2(n982), .ZN(n933) );
  OAI21_X1 U1612 ( .B1(n2089), .B2(n528), .A(n1001), .ZN(n1531) );
  CLKBUF_X3 U1613 ( .A(data_out_x[1]), .Z(n2028) );
  CLKBUF_X3 U1614 ( .A(data_out_x[1]), .Z(n2124) );
  OR2_X1 U1615 ( .A1(n2120), .A2(n193), .ZN(n2030) );
  NAND2_X1 U1616 ( .A1(n1338), .A2(n2030), .ZN(n1866) );
  OR2_X1 U1617 ( .A1(n2118), .A2(n129), .ZN(n2031) );
  NAND2_X1 U1618 ( .A1(n1402), .A2(n2031), .ZN(n1930) );
  BUF_X1 U1619 ( .A(n2085), .Z(n2118) );
  NAND2_X1 U1620 ( .A1(add_r31[15]), .A2(n1), .ZN(n1017) );
  NOR2_X1 U1621 ( .A1(n1018), .A2(clear_acc), .ZN(n982) );
  NAND2_X1 U1622 ( .A1(clc1), .A2(n2170), .ZN(n1002) );
  OR2_X1 U1623 ( .A1(n2090), .A2(n513), .ZN(n2035) );
  NAND2_X1 U1624 ( .A1(n1017), .A2(n2035), .ZN(n1546) );
  BUF_X1 U1625 ( .A(n2081), .Z(n2090) );
  NAND2_X1 U1626 ( .A1(add_r1[15]), .A2(n2047), .ZN(n1498) );
  NAND2_X1 U1627 ( .A1(add_r32[15]), .A2(n2079), .ZN(n1000) );
  NAND2_X1 U1628 ( .A1(add_r2[15]), .A2(n2048), .ZN(n1482) );
  NAND2_X1 U1629 ( .A1(add_r3[15]), .A2(n2049), .ZN(n1466) );
  NAND2_X1 U1630 ( .A1(add_r4[15]), .A2(n2051), .ZN(n1450) );
  NAND2_X1 U1631 ( .A1(add_r5[15]), .A2(n2052), .ZN(n1434) );
  NAND2_X1 U1632 ( .A1(add_r6[15]), .A2(n2053), .ZN(n1418) );
  NAND2_X1 U1633 ( .A1(add_r7[15]), .A2(n2055), .ZN(n1402) );
  NAND2_X1 U1634 ( .A1(add_r8[15]), .A2(n2056), .ZN(n1386) );
  NAND2_X1 U1635 ( .A1(add_r9[15]), .A2(n2057), .ZN(n1370) );
  NAND2_X1 U1636 ( .A1(add_r10[15]), .A2(n2059), .ZN(n1354) );
  NAND2_X1 U1637 ( .A1(add_r11[15]), .A2(n2060), .ZN(n1338) );
  NAND2_X1 U1638 ( .A1(add_r12[15]), .A2(n2061), .ZN(n1322) );
  NAND2_X1 U1639 ( .A1(add_r13[15]), .A2(n2063), .ZN(n1306) );
  NAND2_X1 U1640 ( .A1(add_r14[15]), .A2(n2064), .ZN(n1290) );
  NAND2_X1 U1641 ( .A1(add_r15[15]), .A2(n2065), .ZN(n1274) );
  NAND2_X1 U1642 ( .A1(add_r16[15]), .A2(n985), .ZN(n1258) );
  NAND2_X1 U1643 ( .A1(add_r17[15]), .A2(n2046), .ZN(n1242) );
  NAND2_X1 U1644 ( .A1(add_r18[15]), .A2(n2042), .ZN(n1226) );
  NAND2_X1 U1645 ( .A1(add_r19[15]), .A2(n2046), .ZN(n1210) );
  NAND2_X1 U1646 ( .A1(add_r20[15]), .A2(n985), .ZN(n1194) );
  NAND2_X1 U1647 ( .A1(add_r21[15]), .A2(n985), .ZN(n1178) );
  NAND2_X1 U1648 ( .A1(add_r22[15]), .A2(n2046), .ZN(n1162) );
  NAND2_X1 U1649 ( .A1(add_r23[15]), .A2(n2045), .ZN(n1146) );
  NAND2_X1 U1650 ( .A1(add_r24[15]), .A2(n2068), .ZN(n1130) );
  NAND2_X1 U1651 ( .A1(add_r25[15]), .A2(n2070), .ZN(n1114) );
  NAND2_X1 U1652 ( .A1(add_r26[15]), .A2(n2071), .ZN(n1098) );
  NAND2_X1 U1653 ( .A1(add_r27[15]), .A2(n2072), .ZN(n1082) );
  NAND2_X1 U1654 ( .A1(add_r28[15]), .A2(n2074), .ZN(n1066) );
  NAND2_X1 U1655 ( .A1(add_r29[15]), .A2(n2075), .ZN(n1050) );
  NAND2_X1 U1656 ( .A1(add_r30[15]), .A2(n2076), .ZN(n1034) );
  BUF_X8 U1657 ( .A(data_out_x[5]), .Z(n2137) );
  BUF_X8 U1658 ( .A(data_out_x[6]), .Z(n2140) );
  CLKBUF_X1 U1659 ( .A(n2043), .Z(n2080) );
  CLKBUF_X3 U1660 ( .A(data_out_x[7]), .Z(n2144) );
  INV_X1 U1661 ( .A(addr_y[4]), .ZN(n2149) );
endmodule


module ctrlpath ( clk, reset, start, addr_x, wr_en_x, addr_a1, addr_a2, 
        addr_a3, addr_a4, addr_a5, addr_a6, addr_a7, addr_a8, addr_a9, 
        addr_a10, addr_a11, addr_a12, addr_a13, addr_a14, addr_a15, addr_a16, 
        addr_a17, addr_a18, addr_a19, addr_a20, addr_a21, addr_a22, addr_a23, 
        addr_a24, addr_a25, addr_a26, addr_a27, addr_a28, addr_a29, addr_a30, 
        addr_a31, addr_a32, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, 
        wr_en_a6, wr_en_a7, wr_en_a8, wr_en_a9, wr_en_a10, wr_en_a11, 
        wr_en_a12, wr_en_a13, wr_en_a14, wr_en_a15, wr_en_a16, wr_en_a17, 
        wr_en_a18, wr_en_a19, wr_en_a20, wr_en_a21, wr_en_a22, wr_en_a23, 
        wr_en_a24, wr_en_a25, wr_en_a26, wr_en_a27, wr_en_a28, wr_en_a29, 
        wr_en_a30, wr_en_a31, wr_en_a32, clear_acc, clc, clc1, addr_y, wr_en_y, 
        done, loadMatrix, loadVector );
  output [4:0] addr_x;
  output [4:0] addr_a1;
  output [4:0] addr_a2;
  output [4:0] addr_a3;
  output [4:0] addr_a4;
  output [4:0] addr_a5;
  output [4:0] addr_a6;
  output [4:0] addr_a7;
  output [4:0] addr_a8;
  output [4:0] addr_a9;
  output [4:0] addr_a10;
  output [4:0] addr_a11;
  output [4:0] addr_a12;
  output [4:0] addr_a13;
  output [4:0] addr_a14;
  output [4:0] addr_a15;
  output [4:0] addr_a16;
  output [4:0] addr_a17;
  output [4:0] addr_a18;
  output [4:0] addr_a19;
  output [4:0] addr_a20;
  output [4:0] addr_a21;
  output [4:0] addr_a22;
  output [4:0] addr_a23;
  output [4:0] addr_a24;
  output [4:0] addr_a25;
  output [4:0] addr_a26;
  output [4:0] addr_a27;
  output [4:0] addr_a28;
  output [4:0] addr_a29;
  output [4:0] addr_a30;
  output [4:0] addr_a31;
  output [4:0] addr_a32;
  output [4:0] addr_y;
  input clk, reset, start, loadMatrix, loadVector;
  output wr_en_x, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6,
         wr_en_a7, wr_en_a8, wr_en_a9, wr_en_a10, wr_en_a11, wr_en_a12,
         wr_en_a13, wr_en_a14, wr_en_a15, wr_en_a16, wr_en_a17, wr_en_a18,
         wr_en_a19, wr_en_a20, wr_en_a21, wr_en_a22, wr_en_a23, wr_en_a24,
         wr_en_a25, wr_en_a26, wr_en_a27, wr_en_a28, wr_en_a29, wr_en_a30,
         wr_en_a31, wr_en_a32, clear_acc, clc, clc1, wr_en_y, done;
  wire   N80, N81, N82, N83, N84, N85, N86, N91, N92, N93, N94, N106, N107,
         N108, N109, N121, N122, N123, N124, N136, N137, N138, N139, N151,
         N152, N153, N154, N166, N167, N168, N169, N181, N182, N183, N184,
         N196, N197, N198, N199, N211, N212, N213, N214, N226, N227, N228,
         N229, N241, N242, N243, N244, N256, N257, N258, N259, N271, N272,
         N273, N274, N286, N287, N288, N289, N301, N302, N303, N304, N316,
         N317, N318, N319, N331, N332, N333, N334, N346, N347, N348, N349,
         N361, N362, N363, N364, N376, N377, N378, N379, N391, N392, N393,
         N394, N406, N407, N408, N409, N421, N422, N423, N424, N436, N437,
         N438, N439, N451, N452, N453, N454, N466, N467, N468, N469, N481,
         N482, N483, N484, N496, N497, N498, N499, N511, N512, N513, N514,
         N526, N527, N528, N529, N541, N542, N543, N544, N556, N557, N558,
         N559, N570, N571, N572, N573, N574, N575, N576, N577, N578, N584,
         N585, N586, N587, N595, N596, N597, N604, N606, N608, N610, N612,
         N614, N616, N618, N620, N622, N624, N626, N628, N630, N632, N634,
         N636, N638, N640, N642, N644, N646, N648, N650, N652, N654, N656,
         N658, N660, N662, N664, N666, N668, N674, n321, n354, n355, n358,
         n359, n360, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, \add_501/carry[4] , \add_501/carry[3] ,
         \add_501/carry[2] , \add_494/carry[4] , \add_494/carry[3] ,
         \add_494/carry[2] , \add_485/carry[4] , \add_485/carry[3] ,
         \add_485/carry[2] , \add_476/carry[4] , \add_476/carry[3] ,
         \add_476/carry[2] , \add_467/carry[4] , \add_467/carry[3] ,
         \add_467/carry[2] , \add_458/carry[4] , \add_458/carry[3] ,
         \add_458/carry[2] , \add_449/carry[4] , \add_449/carry[3] ,
         \add_449/carry[2] , \add_440/carry[4] , \add_440/carry[3] ,
         \add_440/carry[2] , \add_431/carry[4] , \add_431/carry[3] ,
         \add_431/carry[2] , \add_422/carry[4] , \add_422/carry[3] ,
         \add_422/carry[2] , \add_413/carry[4] , \add_413/carry[3] ,
         \add_413/carry[2] , \add_404/carry[4] , \add_404/carry[3] ,
         \add_404/carry[2] , \add_395/carry[4] , \add_395/carry[3] ,
         \add_395/carry[2] , \add_386/carry[4] , \add_386/carry[3] ,
         \add_386/carry[2] , \add_377/carry[4] , \add_377/carry[3] ,
         \add_377/carry[2] , \add_368/carry[4] , \add_368/carry[3] ,
         \add_368/carry[2] , \add_359/carry[4] , \add_359/carry[3] ,
         \add_359/carry[2] , \add_350/carry[4] , \add_350/carry[3] ,
         \add_350/carry[2] , \add_341/carry[4] , \add_341/carry[3] ,
         \add_341/carry[2] , \add_332/carry[4] , \add_332/carry[3] ,
         \add_332/carry[2] , \add_323/carry[4] , \add_323/carry[3] ,
         \add_323/carry[2] , \add_314/carry[4] , \add_314/carry[3] ,
         \add_314/carry[2] , \add_305/carry[4] , \add_305/carry[3] ,
         \add_305/carry[2] , \add_296/carry[4] , \add_296/carry[3] ,
         \add_296/carry[2] , \add_287/carry[4] , \add_287/carry[3] ,
         \add_287/carry[2] , \add_278/carry[4] , \add_278/carry[3] ,
         \add_278/carry[2] , \add_269/carry[4] , \add_269/carry[3] ,
         \add_269/carry[2] , \add_260/carry[4] , \add_260/carry[3] ,
         \add_260/carry[2] , \add_251/carry[4] , \add_251/carry[3] ,
         \add_251/carry[2] , \add_242/carry[4] , \add_242/carry[3] ,
         \add_242/carry[2] , \add_233/carry[4] , \add_233/carry[3] ,
         \add_233/carry[2] , \add_224/carry[4] , \add_224/carry[3] ,
         \add_224/carry[2] , \add_215/carry[4] , \add_215/carry[3] ,
         \add_215/carry[2] , \add_206/carry[4] , \add_206/carry[3] ,
         \add_206/carry[2] , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340;
  wire   [5:0] state;

  DFF_X1 \addr_y_reg[0]  ( .D(n113), .CK(clk), .Q(addr_y[0]), .QN(n49) );
  DFF_X1 \addr_y_reg[4]  ( .D(n117), .CK(clk), .Q(addr_y[4]) );
  DFF_X1 done_reg ( .D(N86), .CK(clk), .Q(done) );
  DFF_X1 \state_reg[1]  ( .D(N81), .CK(clk), .Q(state[1]), .QN(n359) );
  DFF_X1 \addr_a25_reg[0]  ( .D(n217), .CK(clk), .Q(addr_a25[0]), .QN(n44) );
  DFF_X1 \addr_a25_reg[4]  ( .D(n221), .CK(clk), .Q(addr_a25[4]) );
  DFF_X1 \state_reg[2]  ( .D(N82), .CK(clk), .Q(state[2]), .QN(n358) );
  DFF_X1 \addr_a25_reg[3]  ( .D(n220), .CK(clk), .Q(addr_a25[3]) );
  DFF_X1 \addr_a25_reg[2]  ( .D(n219), .CK(clk), .Q(addr_a25[2]) );
  DFF_X1 \addr_a25_reg[1]  ( .D(n218), .CK(clk), .Q(addr_a25[1]) );
  DFF_X1 \addr_a2_reg[0]  ( .D(n137), .CK(clk), .Q(addr_a2[0]), .QN(n35) );
  DFF_X1 \addr_a2_reg[1]  ( .D(n138), .CK(clk), .Q(addr_a2[1]) );
  DFF_X1 \addr_a2_reg[2]  ( .D(n139), .CK(clk), .Q(addr_a2[2]) );
  DFF_X1 \addr_a2_reg[3]  ( .D(n140), .CK(clk), .Q(addr_a2[3]) );
  DFF_X1 \addr_a2_reg[4]  ( .D(n141), .CK(clk), .Q(addr_a2[4]) );
  DFF_X1 \state_reg[0]  ( .D(N80), .CK(clk), .Q(state[0]), .QN(n360) );
  DFF_X1 \addr_a5_reg[0]  ( .D(n238), .CK(clk), .Q(addr_a5[0]), .QN(n67) );
  DFF_X1 \addr_a5_reg[1]  ( .D(n239), .CK(clk), .Q(addr_a5[1]) );
  DFF_X1 \addr_a5_reg[2]  ( .D(n240), .CK(clk), .Q(addr_a5[2]) );
  DFF_X1 \addr_a5_reg[3]  ( .D(n241), .CK(clk), .Q(addr_a5[3]) );
  DFF_X1 \addr_a5_reg[4]  ( .D(n242), .CK(clk), .Q(addr_a5[4]) );
  DFF_X1 \state_reg[3]  ( .D(N83), .CK(clk), .Q(state[3]), .QN(n355) );
  DFF_X1 \addr_x_reg[0]  ( .D(N574), .CK(clk), .Q(addr_x[0]), .QN(n68) );
  DFF_X1 \addr_x_reg[1]  ( .D(N575), .CK(clk), .Q(addr_x[1]) );
  DFF_X1 \addr_x_reg[2]  ( .D(N576), .CK(clk), .Q(addr_x[2]) );
  DFF_X1 \addr_x_reg[3]  ( .D(N577), .CK(clk), .Q(addr_x[3]) );
  DFF_X1 \addr_x_reg[4]  ( .D(N578), .CK(clk), .Q(addr_x[4]) );
  DFF_X1 \addr_a32_reg[0]  ( .D(n132), .CK(clk), .Q(addr_a32[0]), .QN(n43) );
  DFF_X1 \addr_a32_reg[1]  ( .D(n133), .CK(clk), .Q(addr_a32[1]) );
  DFF_X1 \addr_a32_reg[2]  ( .D(n134), .CK(clk), .Q(addr_a32[2]) );
  DFF_X1 \addr_a32_reg[3]  ( .D(n135), .CK(clk), .Q(addr_a32[3]) );
  DFF_X1 \addr_a32_reg[4]  ( .D(n136), .CK(clk), .Q(addr_a32[4]) );
  DFF_X1 \state_reg[5]  ( .D(N85), .CK(clk), .Q(state[5]), .QN(n321) );
  DFF_X1 \state_reg[4]  ( .D(N84), .CK(clk), .Q(state[4]), .QN(n354) );
  DFF_X1 \addr_a20_reg[0]  ( .D(n147), .CK(clk), .Q(addr_a20[0]), .QN(n66) );
  DFF_X1 \addr_a20_reg[1]  ( .D(n148), .CK(clk), .Q(addr_a20[1]) );
  DFF_X1 \addr_a20_reg[2]  ( .D(n149), .CK(clk), .Q(addr_a20[2]) );
  DFF_X1 \addr_a20_reg[3]  ( .D(n150), .CK(clk), .Q(addr_a20[3]) );
  DFF_X1 \addr_a20_reg[4]  ( .D(n151), .CK(clk), .Q(addr_a20[4]) );
  DFF_X1 \addr_a19_reg[0]  ( .D(n152), .CK(clk), .Q(addr_a19[0]), .QN(n65) );
  DFF_X1 \addr_a19_reg[1]  ( .D(n153), .CK(clk), .Q(addr_a19[1]) );
  DFF_X1 \addr_a19_reg[2]  ( .D(n154), .CK(clk), .Q(addr_a19[2]) );
  DFF_X1 \addr_a19_reg[3]  ( .D(n155), .CK(clk), .Q(addr_a19[3]) );
  DFF_X1 \addr_a19_reg[4]  ( .D(n156), .CK(clk), .Q(addr_a19[4]) );
  DFF_X1 \addr_a18_reg[0]  ( .D(n142), .CK(clk), .Q(addr_a18[0]), .QN(n64) );
  DFF_X1 \addr_a18_reg[1]  ( .D(n143), .CK(clk), .Q(addr_a18[1]) );
  DFF_X1 \addr_a18_reg[2]  ( .D(n144), .CK(clk), .Q(addr_a18[2]) );
  DFF_X1 \addr_a18_reg[3]  ( .D(n145), .CK(clk), .Q(addr_a18[3]) );
  DFF_X1 \addr_a18_reg[4]  ( .D(n146), .CK(clk), .Q(addr_a18[4]) );
  DFF_X1 \addr_a14_reg[0]  ( .D(n157), .CK(clk), .Q(addr_a14[0]), .QN(n63) );
  DFF_X1 \addr_a14_reg[1]  ( .D(n158), .CK(clk), .Q(addr_a14[1]) );
  DFF_X1 \addr_a14_reg[2]  ( .D(n159), .CK(clk), .Q(addr_a14[2]) );
  DFF_X1 \addr_a14_reg[3]  ( .D(n160), .CK(clk), .Q(addr_a14[3]) );
  DFF_X1 \addr_a14_reg[4]  ( .D(n161), .CK(clk), .Q(addr_a14[4]) );
  DFF_X1 \addr_a17_reg[0]  ( .D(n172), .CK(clk), .Q(addr_a17[0]), .QN(n62) );
  DFF_X1 \addr_a17_reg[1]  ( .D(n173), .CK(clk), .Q(addr_a17[1]) );
  DFF_X1 \addr_a17_reg[2]  ( .D(n174), .CK(clk), .Q(addr_a17[2]) );
  DFF_X1 \addr_a17_reg[3]  ( .D(n175), .CK(clk), .Q(addr_a17[3]) );
  DFF_X1 \addr_a17_reg[4]  ( .D(n176), .CK(clk), .Q(addr_a17[4]) );
  DFF_X1 \addr_a16_reg[0]  ( .D(n167), .CK(clk), .Q(addr_a16[0]), .QN(n61) );
  DFF_X1 \addr_a16_reg[1]  ( .D(n168), .CK(clk), .Q(addr_a16[1]) );
  DFF_X1 \addr_a16_reg[2]  ( .D(n169), .CK(clk), .Q(addr_a16[2]) );
  DFF_X1 \addr_a16_reg[3]  ( .D(n170), .CK(clk), .Q(addr_a16[3]) );
  DFF_X1 \addr_a16_reg[4]  ( .D(n171), .CK(clk), .Q(addr_a16[4]) );
  DFF_X1 \addr_a15_reg[0]  ( .D(n162), .CK(clk), .Q(addr_a15[0]), .QN(n60) );
  DFF_X1 \addr_a15_reg[1]  ( .D(n163), .CK(clk), .Q(addr_a15[1]) );
  DFF_X1 \addr_a15_reg[2]  ( .D(n164), .CK(clk), .Q(addr_a15[2]) );
  DFF_X1 \addr_a15_reg[3]  ( .D(n165), .CK(clk), .Q(addr_a15[3]) );
  DFF_X1 \addr_a15_reg[4]  ( .D(n166), .CK(clk), .Q(addr_a15[4]) );
  DFF_X1 \addr_a13_reg[0]  ( .D(n187), .CK(clk), .Q(addr_a13[0]), .QN(n48) );
  DFF_X1 \addr_a13_reg[1]  ( .D(n188), .CK(clk), .Q(addr_a13[1]) );
  DFF_X1 \addr_a13_reg[2]  ( .D(n189), .CK(clk), .Q(addr_a13[2]) );
  DFF_X1 \addr_a13_reg[3]  ( .D(n190), .CK(clk), .Q(addr_a13[3]) );
  DFF_X1 \addr_a13_reg[4]  ( .D(n191), .CK(clk), .Q(addr_a13[4]) );
  DFF_X1 \addr_a23_reg[0]  ( .D(n182), .CK(clk), .Q(addr_a23[0]), .QN(n42) );
  DFF_X1 \addr_a23_reg[1]  ( .D(n183), .CK(clk), .Q(addr_a23[1]) );
  DFF_X1 \addr_a23_reg[2]  ( .D(n184), .CK(clk), .Q(addr_a23[2]) );
  DFF_X1 \addr_a23_reg[3]  ( .D(n185), .CK(clk), .Q(addr_a23[3]) );
  DFF_X1 \addr_a23_reg[4]  ( .D(n186), .CK(clk), .Q(addr_a23[4]) );
  DFF_X1 \addr_a22_reg[0]  ( .D(n177), .CK(clk), .Q(addr_a22[0]), .QN(n47) );
  DFF_X1 \addr_a22_reg[1]  ( .D(n178), .CK(clk), .Q(addr_a22[1]) );
  DFF_X1 \addr_a22_reg[2]  ( .D(n179), .CK(clk), .Q(addr_a22[2]) );
  DFF_X1 \addr_a22_reg[3]  ( .D(n180), .CK(clk), .Q(addr_a22[3]) );
  DFF_X1 \addr_a22_reg[4]  ( .D(n181), .CK(clk), .Q(addr_a22[4]) );
  DFF_X1 \addr_a21_reg[0]  ( .D(n192), .CK(clk), .Q(addr_a21[0]), .QN(n46) );
  DFF_X1 \addr_a21_reg[1]  ( .D(n193), .CK(clk), .Q(addr_a21[1]) );
  DFF_X1 \addr_a21_reg[2]  ( .D(n194), .CK(clk), .Q(addr_a21[2]) );
  DFF_X1 \addr_a21_reg[3]  ( .D(n195), .CK(clk), .Q(addr_a21[3]) );
  DFF_X1 \addr_a21_reg[4]  ( .D(n196), .CK(clk), .Q(addr_a21[4]) );
  DFF_X1 \addr_a29_reg[0]  ( .D(n222), .CK(clk), .Q(addr_a29[0]), .QN(n41) );
  DFF_X1 \addr_a29_reg[1]  ( .D(n223), .CK(clk), .Q(addr_a29[1]) );
  DFF_X1 \addr_a29_reg[2]  ( .D(n224), .CK(clk), .Q(addr_a29[2]) );
  DFF_X1 \addr_a29_reg[3]  ( .D(n225), .CK(clk), .Q(addr_a29[3]) );
  DFF_X1 \addr_a29_reg[4]  ( .D(n226), .CK(clk), .Q(addr_a29[4]) );
  DFF_X1 \addr_a27_reg[0]  ( .D(n212), .CK(clk), .Q(addr_a27[0]), .QN(n40) );
  DFF_X1 \addr_a27_reg[1]  ( .D(n213), .CK(clk), .Q(addr_a27[1]) );
  DFF_X1 \addr_a27_reg[2]  ( .D(n214), .CK(clk), .Q(addr_a27[2]) );
  DFF_X1 \addr_a27_reg[3]  ( .D(n215), .CK(clk), .Q(addr_a27[3]) );
  DFF_X1 \addr_a27_reg[4]  ( .D(n216), .CK(clk), .Q(addr_a27[4]) );
  DFF_X1 \addr_a24_reg[0]  ( .D(n207), .CK(clk), .Q(addr_a24[0]), .QN(n39) );
  DFF_X1 \addr_a24_reg[1]  ( .D(n208), .CK(clk), .Q(addr_a24[1]) );
  DFF_X1 \addr_a24_reg[2]  ( .D(n209), .CK(clk), .Q(addr_a24[2]) );
  DFF_X1 \addr_a24_reg[3]  ( .D(n210), .CK(clk), .Q(addr_a24[3]) );
  DFF_X1 \addr_a24_reg[4]  ( .D(n211), .CK(clk), .Q(addr_a24[4]) );
  DFF_X1 \addr_a28_reg[0]  ( .D(n202), .CK(clk), .Q(addr_a28[0]), .QN(n59) );
  DFF_X1 \addr_a28_reg[1]  ( .D(n203), .CK(clk), .Q(addr_a28[1]) );
  DFF_X1 \addr_a28_reg[2]  ( .D(n204), .CK(clk), .Q(addr_a28[2]) );
  DFF_X1 \addr_a28_reg[3]  ( .D(n205), .CK(clk), .Q(addr_a28[3]) );
  DFF_X1 \addr_a28_reg[4]  ( .D(n206), .CK(clk), .Q(addr_a28[4]) );
  DFF_X1 \addr_a26_reg[0]  ( .D(n197), .CK(clk), .Q(addr_a26[0]), .QN(n58) );
  DFF_X1 \addr_a26_reg[1]  ( .D(n198), .CK(clk), .Q(addr_a26[1]) );
  DFF_X1 \addr_a26_reg[2]  ( .D(n199), .CK(clk), .Q(addr_a26[2]) );
  DFF_X1 \addr_a26_reg[3]  ( .D(n200), .CK(clk), .Q(addr_a26[3]) );
  DFF_X1 \addr_a26_reg[4]  ( .D(n201), .CK(clk), .Q(addr_a26[4]) );
  DFF_X1 \addr_a1_reg[0]  ( .D(n279), .CK(clk), .Q(addr_a1[0]), .QN(n45) );
  DFF_X1 \addr_a1_reg[1]  ( .D(n280), .CK(clk), .Q(addr_a1[1]) );
  DFF_X1 \addr_a1_reg[2]  ( .D(n281), .CK(clk), .Q(addr_a1[2]) );
  DFF_X1 \addr_a1_reg[3]  ( .D(n282), .CK(clk), .Q(addr_a1[3]) );
  DFF_X1 \addr_a1_reg[4]  ( .D(n283), .CK(clk), .Q(addr_a1[4]) );
  DFF_X1 \addr_a4_reg[0]  ( .D(n233), .CK(clk), .Q(addr_a4[0]), .QN(n57) );
  DFF_X1 \addr_a4_reg[1]  ( .D(n234), .CK(clk), .Q(addr_a4[1]) );
  DFF_X1 \addr_a4_reg[2]  ( .D(n235), .CK(clk), .Q(addr_a4[2]) );
  DFF_X1 \addr_a4_reg[3]  ( .D(n236), .CK(clk), .Q(addr_a4[3]) );
  DFF_X1 \addr_a4_reg[4]  ( .D(n237), .CK(clk), .Q(addr_a4[4]) );
  DFF_X1 \addr_a31_reg[0]  ( .D(n127), .CK(clk), .Q(addr_a31[0]), .QN(n38) );
  DFF_X1 \addr_a31_reg[1]  ( .D(n128), .CK(clk), .Q(addr_a31[1]) );
  DFF_X1 \addr_a31_reg[2]  ( .D(n129), .CK(clk), .Q(addr_a31[2]) );
  DFF_X1 \addr_a31_reg[3]  ( .D(n130), .CK(clk), .Q(addr_a31[3]) );
  DFF_X1 \addr_a31_reg[4]  ( .D(n131), .CK(clk), .Q(addr_a31[4]) );
  DFF_X1 \addr_a30_reg[0]  ( .D(n122), .CK(clk), .Q(addr_a30[0]), .QN(n37) );
  DFF_X1 \addr_a30_reg[1]  ( .D(n123), .CK(clk), .Q(addr_a30[1]) );
  DFF_X1 \addr_a30_reg[2]  ( .D(n124), .CK(clk), .Q(addr_a30[2]) );
  DFF_X1 \addr_a30_reg[3]  ( .D(n125), .CK(clk), .Q(addr_a30[3]) );
  DFF_X1 \addr_a30_reg[4]  ( .D(n126), .CK(clk), .Q(addr_a30[4]) );
  DFF_X1 \addr_a7_reg[0]  ( .D(n274), .CK(clk), .Q(addr_a7[0]), .QN(n56) );
  DFF_X1 \addr_a7_reg[1]  ( .D(n275), .CK(clk), .Q(addr_a7[1]) );
  DFF_X1 \addr_a7_reg[2]  ( .D(n276), .CK(clk), .Q(addr_a7[2]) );
  DFF_X1 \addr_a7_reg[3]  ( .D(n277), .CK(clk), .Q(addr_a7[3]) );
  DFF_X1 \addr_a7_reg[4]  ( .D(n278), .CK(clk), .Q(addr_a7[4]) );
  DFF_X1 \addr_a8_reg[0]  ( .D(n269), .CK(clk), .Q(addr_a8[0]), .QN(n55) );
  DFF_X1 \addr_a8_reg[1]  ( .D(n270), .CK(clk), .Q(addr_a8[1]) );
  DFF_X1 \addr_a8_reg[2]  ( .D(n271), .CK(clk), .Q(addr_a8[2]) );
  DFF_X1 \addr_a8_reg[3]  ( .D(n272), .CK(clk), .Q(addr_a8[3]) );
  DFF_X1 \addr_a8_reg[4]  ( .D(n273), .CK(clk), .Q(addr_a8[4]) );
  DFF_X1 \addr_a11_reg[0]  ( .D(n264), .CK(clk), .Q(addr_a11[0]), .QN(n54) );
  DFF_X1 \addr_a11_reg[1]  ( .D(n265), .CK(clk), .Q(addr_a11[1]) );
  DFF_X1 \addr_a11_reg[2]  ( .D(n266), .CK(clk), .Q(addr_a11[2]) );
  DFF_X1 \addr_a11_reg[3]  ( .D(n267), .CK(clk), .Q(addr_a11[3]) );
  DFF_X1 \addr_a11_reg[4]  ( .D(n268), .CK(clk), .Q(addr_a11[4]) );
  DFF_X1 \addr_a12_reg[0]  ( .D(n259), .CK(clk), .Q(addr_a12[0]), .QN(n53) );
  DFF_X1 \addr_a12_reg[1]  ( .D(n260), .CK(clk), .Q(addr_a12[1]) );
  DFF_X1 \addr_a12_reg[2]  ( .D(n261), .CK(clk), .Q(addr_a12[2]) );
  DFF_X1 \addr_a12_reg[3]  ( .D(n262), .CK(clk), .Q(addr_a12[3]) );
  DFF_X1 \addr_a12_reg[4]  ( .D(n263), .CK(clk), .Q(addr_a12[4]) );
  DFF_X1 \addr_a10_reg[0]  ( .D(n254), .CK(clk), .Q(addr_a10[0]), .QN(n52) );
  DFF_X1 \addr_a10_reg[1]  ( .D(n255), .CK(clk), .Q(addr_a10[1]) );
  DFF_X1 \addr_a10_reg[2]  ( .D(n256), .CK(clk), .Q(addr_a10[2]) );
  DFF_X1 \addr_a10_reg[3]  ( .D(n257), .CK(clk), .Q(addr_a10[3]) );
  DFF_X1 \addr_a10_reg[4]  ( .D(n258), .CK(clk), .Q(addr_a10[4]) );
  DFF_X1 \addr_a9_reg[0]  ( .D(n249), .CK(clk), .Q(addr_a9[0]), .QN(n51) );
  DFF_X1 \addr_a9_reg[1]  ( .D(n250), .CK(clk), .Q(addr_a9[1]) );
  DFF_X1 \addr_a9_reg[2]  ( .D(n251), .CK(clk), .Q(addr_a9[2]) );
  DFF_X1 \addr_a9_reg[3]  ( .D(n252), .CK(clk), .Q(addr_a9[3]) );
  DFF_X1 \addr_a9_reg[4]  ( .D(n253), .CK(clk), .Q(addr_a9[4]) );
  DFF_X1 \addr_a6_reg[0]  ( .D(n244), .CK(clk), .Q(addr_a6[0]), .QN(n50) );
  DFF_X1 \addr_a6_reg[1]  ( .D(n245), .CK(clk), .Q(addr_a6[1]) );
  DFF_X1 \addr_a6_reg[2]  ( .D(n246), .CK(clk), .Q(addr_a6[2]) );
  DFF_X1 \addr_a6_reg[3]  ( .D(n247), .CK(clk), .Q(addr_a6[3]) );
  DFF_X1 \addr_a6_reg[4]  ( .D(n248), .CK(clk), .Q(addr_a6[4]) );
  DFF_X1 \addr_a3_reg[0]  ( .D(n228), .CK(clk), .Q(addr_a3[0]), .QN(n36) );
  DFF_X1 \addr_a3_reg[1]  ( .D(n229), .CK(clk), .Q(addr_a3[1]) );
  DFF_X1 \addr_a3_reg[2]  ( .D(n230), .CK(clk), .Q(addr_a3[2]) );
  DFF_X1 \addr_a3_reg[3]  ( .D(n231), .CK(clk), .Q(addr_a3[3]) );
  DFF_X1 \addr_a3_reg[4]  ( .D(n232), .CK(clk), .Q(addr_a3[4]) );
  DFF_X1 \addr_y_reg[3]  ( .D(n116), .CK(clk), .Q(addr_y[3]) );
  DFF_X1 \addr_y_reg[2]  ( .D(n115), .CK(clk), .Q(addr_y[2]) );
  DFF_X1 \addr_y_reg[1]  ( .D(n114), .CK(clk), .Q(addr_y[1]) );
  DFF_X1 clear_acc_reg ( .D(N595), .CK(clk), .Q(clear_acc) );
  DFF_X1 clc_reg ( .D(N596), .CK(clk), .Q(clc) );
  DFF_X1 clc1_reg ( .D(N597), .CK(clk), .Q(clc1) );
  NAND3_X1 U720 ( .A1(n419), .A2(n298), .A3(n420), .ZN(n418) );
  NAND3_X1 U721 ( .A1(n444), .A2(n295), .A3(n298), .ZN(n441) );
  NAND3_X1 U722 ( .A1(n454), .A2(n340), .A3(loadVector), .ZN(n452) );
  NAND3_X1 U723 ( .A1(n354), .A2(n321), .A3(n492), .ZN(n491) );
  NAND3_X1 U724 ( .A1(state[2]), .A2(n493), .A3(n328), .ZN(n490) );
  NAND3_X1 U725 ( .A1(N666), .A2(n313), .A3(n502), .ZN(n501) );
  NAND3_X1 U726 ( .A1(n534), .A2(n391), .A3(N658), .ZN(n533) );
  NAND3_X1 U727 ( .A1(n303), .A2(n391), .A3(n542), .ZN(n541) );
  NAND3_X1 U728 ( .A1(n534), .A2(n389), .A3(N654), .ZN(n550) );
  NAND3_X1 U729 ( .A1(n542), .A2(n444), .A3(N650), .ZN(n564) );
  NAND3_X1 U730 ( .A1(n292), .A2(n400), .A3(n598), .ZN(n605) );
  NAND3_X1 U731 ( .A1(n614), .A2(n624), .A3(N630), .ZN(n647) );
  NAND3_X1 U732 ( .A1(n287), .A2(n590), .A3(n574), .ZN(n654) );
  NAND3_X1 U733 ( .A1(n294), .A2(n408), .A3(n664), .ZN(n671) );
  NAND3_X1 U734 ( .A1(N620), .A2(n381), .A3(n689), .ZN(n688) );
  NAND3_X1 U735 ( .A1(N618), .A2(n680), .A3(n697), .ZN(n696) );
  NAND3_X1 U736 ( .A1(n689), .A2(n378), .A3(N614), .ZN(n715) );
  NAND3_X1 U737 ( .A1(n427), .A2(n383), .A3(n243), .ZN(n722) );
  NAND3_X1 U738 ( .A1(n243), .A2(n420), .A3(N610), .ZN(n730) );
  NAND3_X1 U739 ( .A1(n409), .A2(n387), .A3(n419), .ZN(n708) );
  NAND3_X1 U740 ( .A1(n517), .A2(n750), .A3(N606), .ZN(n747) );
  NAND3_X1 U741 ( .A1(n420), .A2(n739), .A3(n755), .ZN(n749) );
  NAND3_X1 U742 ( .A1(n761), .A2(n354), .A3(state[3]), .ZN(n760) );
  NAND3_X1 U743 ( .A1(n681), .A2(n380), .A3(n295), .ZN(n723) );
  NAND3_X1 U744 ( .A1(n407), .A2(n406), .A3(n408), .ZN(n698) );
  NAND3_X1 U745 ( .A1(n392), .A2(n388), .A3(n526), .ZN(n424) );
  NAND3_X1 U746 ( .A1(n360), .A2(n358), .A3(state[1]), .ZN(n772) );
  HA_X1 \add_501/U1_1_1  ( .A(addr_y[1]), .B(addr_y[0]), .CO(
        \add_501/carry[2] ), .S(N584) );
  HA_X1 \add_501/U1_1_2  ( .A(addr_y[2]), .B(\add_501/carry[2] ), .CO(
        \add_501/carry[3] ), .S(N585) );
  HA_X1 \add_501/U1_1_3  ( .A(addr_y[3]), .B(\add_501/carry[3] ), .CO(
        \add_501/carry[4] ), .S(N586) );
  HA_X1 \add_494/U1_1_1  ( .A(addr_x[1]), .B(addr_x[0]), .CO(
        \add_494/carry[2] ), .S(N570) );
  HA_X1 \add_494/U1_1_2  ( .A(addr_x[2]), .B(\add_494/carry[2] ), .CO(
        \add_494/carry[3] ), .S(N571) );
  HA_X1 \add_494/U1_1_3  ( .A(addr_x[3]), .B(\add_494/carry[3] ), .CO(
        \add_494/carry[4] ), .S(N572) );
  HA_X1 \add_485/U1_1_1  ( .A(addr_a32[1]), .B(addr_a32[0]), .CO(
        \add_485/carry[2] ), .S(N556) );
  HA_X1 \add_485/U1_1_2  ( .A(addr_a32[2]), .B(\add_485/carry[2] ), .CO(
        \add_485/carry[3] ), .S(N557) );
  HA_X1 \add_485/U1_1_3  ( .A(addr_a32[3]), .B(\add_485/carry[3] ), .CO(
        \add_485/carry[4] ), .S(N558) );
  HA_X1 \add_476/U1_1_1  ( .A(addr_a31[1]), .B(addr_a31[0]), .CO(
        \add_476/carry[2] ), .S(N541) );
  HA_X1 \add_476/U1_1_2  ( .A(addr_a31[2]), .B(\add_476/carry[2] ), .CO(
        \add_476/carry[3] ), .S(N542) );
  HA_X1 \add_476/U1_1_3  ( .A(addr_a31[3]), .B(\add_476/carry[3] ), .CO(
        \add_476/carry[4] ), .S(N543) );
  HA_X1 \add_467/U1_1_1  ( .A(addr_a30[1]), .B(addr_a30[0]), .CO(
        \add_467/carry[2] ), .S(N526) );
  HA_X1 \add_467/U1_1_2  ( .A(addr_a30[2]), .B(\add_467/carry[2] ), .CO(
        \add_467/carry[3] ), .S(N527) );
  HA_X1 \add_467/U1_1_3  ( .A(addr_a30[3]), .B(\add_467/carry[3] ), .CO(
        \add_467/carry[4] ), .S(N528) );
  HA_X1 \add_458/U1_1_1  ( .A(addr_a29[1]), .B(addr_a29[0]), .CO(
        \add_458/carry[2] ), .S(N511) );
  HA_X1 \add_458/U1_1_2  ( .A(addr_a29[2]), .B(\add_458/carry[2] ), .CO(
        \add_458/carry[3] ), .S(N512) );
  HA_X1 \add_458/U1_1_3  ( .A(addr_a29[3]), .B(\add_458/carry[3] ), .CO(
        \add_458/carry[4] ), .S(N513) );
  HA_X1 \add_449/U1_1_1  ( .A(addr_a28[1]), .B(addr_a28[0]), .CO(
        \add_449/carry[2] ), .S(N496) );
  HA_X1 \add_449/U1_1_2  ( .A(addr_a28[2]), .B(\add_449/carry[2] ), .CO(
        \add_449/carry[3] ), .S(N497) );
  HA_X1 \add_449/U1_1_3  ( .A(addr_a28[3]), .B(\add_449/carry[3] ), .CO(
        \add_449/carry[4] ), .S(N498) );
  HA_X1 \add_440/U1_1_1  ( .A(addr_a27[1]), .B(addr_a27[0]), .CO(
        \add_440/carry[2] ), .S(N481) );
  HA_X1 \add_440/U1_1_2  ( .A(addr_a27[2]), .B(\add_440/carry[2] ), .CO(
        \add_440/carry[3] ), .S(N482) );
  HA_X1 \add_440/U1_1_3  ( .A(addr_a27[3]), .B(\add_440/carry[3] ), .CO(
        \add_440/carry[4] ), .S(N483) );
  HA_X1 \add_431/U1_1_1  ( .A(addr_a26[1]), .B(addr_a26[0]), .CO(
        \add_431/carry[2] ), .S(N466) );
  HA_X1 \add_431/U1_1_2  ( .A(addr_a26[2]), .B(\add_431/carry[2] ), .CO(
        \add_431/carry[3] ), .S(N467) );
  HA_X1 \add_431/U1_1_3  ( .A(addr_a26[3]), .B(\add_431/carry[3] ), .CO(
        \add_431/carry[4] ), .S(N468) );
  HA_X1 \add_422/U1_1_1  ( .A(addr_a25[1]), .B(addr_a25[0]), .CO(
        \add_422/carry[2] ), .S(N451) );
  HA_X1 \add_422/U1_1_2  ( .A(addr_a25[2]), .B(\add_422/carry[2] ), .CO(
        \add_422/carry[3] ), .S(N452) );
  HA_X1 \add_422/U1_1_3  ( .A(addr_a25[3]), .B(\add_422/carry[3] ), .CO(
        \add_422/carry[4] ), .S(N453) );
  HA_X1 \add_413/U1_1_1  ( .A(addr_a24[1]), .B(addr_a24[0]), .CO(
        \add_413/carry[2] ), .S(N436) );
  HA_X1 \add_413/U1_1_2  ( .A(addr_a24[2]), .B(\add_413/carry[2] ), .CO(
        \add_413/carry[3] ), .S(N437) );
  HA_X1 \add_413/U1_1_3  ( .A(addr_a24[3]), .B(\add_413/carry[3] ), .CO(
        \add_413/carry[4] ), .S(N438) );
  HA_X1 \add_404/U1_1_1  ( .A(addr_a23[1]), .B(addr_a23[0]), .CO(
        \add_404/carry[2] ), .S(N421) );
  HA_X1 \add_404/U1_1_2  ( .A(addr_a23[2]), .B(\add_404/carry[2] ), .CO(
        \add_404/carry[3] ), .S(N422) );
  HA_X1 \add_404/U1_1_3  ( .A(addr_a23[3]), .B(\add_404/carry[3] ), .CO(
        \add_404/carry[4] ), .S(N423) );
  HA_X1 \add_395/U1_1_1  ( .A(addr_a22[1]), .B(addr_a22[0]), .CO(
        \add_395/carry[2] ), .S(N406) );
  HA_X1 \add_395/U1_1_2  ( .A(addr_a22[2]), .B(\add_395/carry[2] ), .CO(
        \add_395/carry[3] ), .S(N407) );
  HA_X1 \add_395/U1_1_3  ( .A(addr_a22[3]), .B(\add_395/carry[3] ), .CO(
        \add_395/carry[4] ), .S(N408) );
  HA_X1 \add_386/U1_1_1  ( .A(addr_a21[1]), .B(addr_a21[0]), .CO(
        \add_386/carry[2] ), .S(N391) );
  HA_X1 \add_386/U1_1_2  ( .A(addr_a21[2]), .B(\add_386/carry[2] ), .CO(
        \add_386/carry[3] ), .S(N392) );
  HA_X1 \add_386/U1_1_3  ( .A(addr_a21[3]), .B(\add_386/carry[3] ), .CO(
        \add_386/carry[4] ), .S(N393) );
  HA_X1 \add_377/U1_1_1  ( .A(addr_a20[1]), .B(addr_a20[0]), .CO(
        \add_377/carry[2] ), .S(N376) );
  HA_X1 \add_377/U1_1_2  ( .A(addr_a20[2]), .B(\add_377/carry[2] ), .CO(
        \add_377/carry[3] ), .S(N377) );
  HA_X1 \add_377/U1_1_3  ( .A(addr_a20[3]), .B(\add_377/carry[3] ), .CO(
        \add_377/carry[4] ), .S(N378) );
  HA_X1 \add_368/U1_1_1  ( .A(addr_a19[1]), .B(addr_a19[0]), .CO(
        \add_368/carry[2] ), .S(N361) );
  HA_X1 \add_368/U1_1_2  ( .A(addr_a19[2]), .B(\add_368/carry[2] ), .CO(
        \add_368/carry[3] ), .S(N362) );
  HA_X1 \add_368/U1_1_3  ( .A(addr_a19[3]), .B(\add_368/carry[3] ), .CO(
        \add_368/carry[4] ), .S(N363) );
  HA_X1 \add_359/U1_1_1  ( .A(addr_a18[1]), .B(addr_a18[0]), .CO(
        \add_359/carry[2] ), .S(N346) );
  HA_X1 \add_359/U1_1_2  ( .A(addr_a18[2]), .B(\add_359/carry[2] ), .CO(
        \add_359/carry[3] ), .S(N347) );
  HA_X1 \add_359/U1_1_3  ( .A(addr_a18[3]), .B(\add_359/carry[3] ), .CO(
        \add_359/carry[4] ), .S(N348) );
  HA_X1 \add_350/U1_1_1  ( .A(addr_a17[1]), .B(addr_a17[0]), .CO(
        \add_350/carry[2] ), .S(N331) );
  HA_X1 \add_350/U1_1_2  ( .A(addr_a17[2]), .B(\add_350/carry[2] ), .CO(
        \add_350/carry[3] ), .S(N332) );
  HA_X1 \add_350/U1_1_3  ( .A(addr_a17[3]), .B(\add_350/carry[3] ), .CO(
        \add_350/carry[4] ), .S(N333) );
  HA_X1 \add_341/U1_1_1  ( .A(addr_a16[1]), .B(addr_a16[0]), .CO(
        \add_341/carry[2] ), .S(N316) );
  HA_X1 \add_341/U1_1_2  ( .A(addr_a16[2]), .B(\add_341/carry[2] ), .CO(
        \add_341/carry[3] ), .S(N317) );
  HA_X1 \add_341/U1_1_3  ( .A(addr_a16[3]), .B(\add_341/carry[3] ), .CO(
        \add_341/carry[4] ), .S(N318) );
  HA_X1 \add_332/U1_1_1  ( .A(addr_a15[1]), .B(addr_a15[0]), .CO(
        \add_332/carry[2] ), .S(N301) );
  HA_X1 \add_332/U1_1_2  ( .A(addr_a15[2]), .B(\add_332/carry[2] ), .CO(
        \add_332/carry[3] ), .S(N302) );
  HA_X1 \add_332/U1_1_3  ( .A(addr_a15[3]), .B(\add_332/carry[3] ), .CO(
        \add_332/carry[4] ), .S(N303) );
  HA_X1 \add_323/U1_1_1  ( .A(addr_a14[1]), .B(addr_a14[0]), .CO(
        \add_323/carry[2] ), .S(N286) );
  HA_X1 \add_323/U1_1_2  ( .A(addr_a14[2]), .B(\add_323/carry[2] ), .CO(
        \add_323/carry[3] ), .S(N287) );
  HA_X1 \add_323/U1_1_3  ( .A(addr_a14[3]), .B(\add_323/carry[3] ), .CO(
        \add_323/carry[4] ), .S(N288) );
  HA_X1 \add_314/U1_1_1  ( .A(addr_a13[1]), .B(addr_a13[0]), .CO(
        \add_314/carry[2] ), .S(N271) );
  HA_X1 \add_314/U1_1_2  ( .A(addr_a13[2]), .B(\add_314/carry[2] ), .CO(
        \add_314/carry[3] ), .S(N272) );
  HA_X1 \add_314/U1_1_3  ( .A(addr_a13[3]), .B(\add_314/carry[3] ), .CO(
        \add_314/carry[4] ), .S(N273) );
  HA_X1 \add_305/U1_1_1  ( .A(addr_a12[1]), .B(addr_a12[0]), .CO(
        \add_305/carry[2] ), .S(N256) );
  HA_X1 \add_305/U1_1_2  ( .A(addr_a12[2]), .B(\add_305/carry[2] ), .CO(
        \add_305/carry[3] ), .S(N257) );
  HA_X1 \add_305/U1_1_3  ( .A(addr_a12[3]), .B(\add_305/carry[3] ), .CO(
        \add_305/carry[4] ), .S(N258) );
  HA_X1 \add_296/U1_1_1  ( .A(addr_a11[1]), .B(addr_a11[0]), .CO(
        \add_296/carry[2] ), .S(N241) );
  HA_X1 \add_296/U1_1_2  ( .A(addr_a11[2]), .B(\add_296/carry[2] ), .CO(
        \add_296/carry[3] ), .S(N242) );
  HA_X1 \add_296/U1_1_3  ( .A(addr_a11[3]), .B(\add_296/carry[3] ), .CO(
        \add_296/carry[4] ), .S(N243) );
  HA_X1 \add_287/U1_1_1  ( .A(addr_a10[1]), .B(addr_a10[0]), .CO(
        \add_287/carry[2] ), .S(N226) );
  HA_X1 \add_287/U1_1_2  ( .A(addr_a10[2]), .B(\add_287/carry[2] ), .CO(
        \add_287/carry[3] ), .S(N227) );
  HA_X1 \add_287/U1_1_3  ( .A(addr_a10[3]), .B(\add_287/carry[3] ), .CO(
        \add_287/carry[4] ), .S(N228) );
  HA_X1 \add_278/U1_1_1  ( .A(addr_a9[1]), .B(addr_a9[0]), .CO(
        \add_278/carry[2] ), .S(N211) );
  HA_X1 \add_278/U1_1_2  ( .A(addr_a9[2]), .B(\add_278/carry[2] ), .CO(
        \add_278/carry[3] ), .S(N212) );
  HA_X1 \add_278/U1_1_3  ( .A(addr_a9[3]), .B(\add_278/carry[3] ), .CO(
        \add_278/carry[4] ), .S(N213) );
  HA_X1 \add_269/U1_1_1  ( .A(addr_a8[1]), .B(addr_a8[0]), .CO(
        \add_269/carry[2] ), .S(N196) );
  HA_X1 \add_269/U1_1_2  ( .A(addr_a8[2]), .B(\add_269/carry[2] ), .CO(
        \add_269/carry[3] ), .S(N197) );
  HA_X1 \add_269/U1_1_3  ( .A(addr_a8[3]), .B(\add_269/carry[3] ), .CO(
        \add_269/carry[4] ), .S(N198) );
  HA_X1 \add_260/U1_1_1  ( .A(addr_a7[1]), .B(addr_a7[0]), .CO(
        \add_260/carry[2] ), .S(N181) );
  HA_X1 \add_260/U1_1_2  ( .A(addr_a7[2]), .B(\add_260/carry[2] ), .CO(
        \add_260/carry[3] ), .S(N182) );
  HA_X1 \add_260/U1_1_3  ( .A(addr_a7[3]), .B(\add_260/carry[3] ), .CO(
        \add_260/carry[4] ), .S(N183) );
  HA_X1 \add_251/U1_1_1  ( .A(addr_a6[1]), .B(addr_a6[0]), .CO(
        \add_251/carry[2] ), .S(N166) );
  HA_X1 \add_251/U1_1_2  ( .A(addr_a6[2]), .B(\add_251/carry[2] ), .CO(
        \add_251/carry[3] ), .S(N167) );
  HA_X1 \add_251/U1_1_3  ( .A(addr_a6[3]), .B(\add_251/carry[3] ), .CO(
        \add_251/carry[4] ), .S(N168) );
  HA_X1 \add_242/U1_1_1  ( .A(addr_a5[1]), .B(addr_a5[0]), .CO(
        \add_242/carry[2] ), .S(N151) );
  HA_X1 \add_242/U1_1_2  ( .A(addr_a5[2]), .B(\add_242/carry[2] ), .CO(
        \add_242/carry[3] ), .S(N152) );
  HA_X1 \add_242/U1_1_3  ( .A(addr_a5[3]), .B(\add_242/carry[3] ), .CO(
        \add_242/carry[4] ), .S(N153) );
  HA_X1 \add_233/U1_1_1  ( .A(addr_a4[1]), .B(addr_a4[0]), .CO(
        \add_233/carry[2] ), .S(N136) );
  HA_X1 \add_233/U1_1_2  ( .A(addr_a4[2]), .B(\add_233/carry[2] ), .CO(
        \add_233/carry[3] ), .S(N137) );
  HA_X1 \add_233/U1_1_3  ( .A(addr_a4[3]), .B(\add_233/carry[3] ), .CO(
        \add_233/carry[4] ), .S(N138) );
  HA_X1 \add_224/U1_1_1  ( .A(addr_a3[1]), .B(addr_a3[0]), .CO(
        \add_224/carry[2] ), .S(N121) );
  HA_X1 \add_224/U1_1_2  ( .A(addr_a3[2]), .B(\add_224/carry[2] ), .CO(
        \add_224/carry[3] ), .S(N122) );
  HA_X1 \add_224/U1_1_3  ( .A(addr_a3[3]), .B(\add_224/carry[3] ), .CO(
        \add_224/carry[4] ), .S(N123) );
  HA_X1 \add_215/U1_1_1  ( .A(addr_a2[1]), .B(addr_a2[0]), .CO(
        \add_215/carry[2] ), .S(N106) );
  HA_X1 \add_215/U1_1_2  ( .A(addr_a2[2]), .B(\add_215/carry[2] ), .CO(
        \add_215/carry[3] ), .S(N107) );
  HA_X1 \add_215/U1_1_3  ( .A(addr_a2[3]), .B(\add_215/carry[3] ), .CO(
        \add_215/carry[4] ), .S(N108) );
  HA_X1 \add_206/U1_1_1  ( .A(addr_a1[1]), .B(addr_a1[0]), .CO(
        \add_206/carry[2] ), .S(N91) );
  HA_X1 \add_206/U1_1_2  ( .A(addr_a1[2]), .B(\add_206/carry[2] ), .CO(
        \add_206/carry[3] ), .S(N92) );
  HA_X1 \add_206/U1_1_3  ( .A(addr_a1[3]), .B(\add_206/carry[3] ), .CO(
        \add_206/carry[4] ), .S(N93) );
  NOR3_X1 U3 ( .A1(n360), .A2(state[2]), .A3(n359), .ZN(n761) );
  NOR2_X1 U4 ( .A1(n424), .A2(n433), .ZN(n589) );
  NOR3_X1 U5 ( .A1(n707), .A2(n316), .A3(n708), .ZN(n680) );
  NOR2_X1 U6 ( .A1(n749), .A2(n227), .ZN(n566) );
  INV_X1 U7 ( .A(n740), .ZN(n227) );
  NOR2_X1 U8 ( .A1(n310), .A2(n314), .ZN(n623) );
  BUF_X1 U9 ( .A(n411), .Z(n73) );
  BUF_X1 U10 ( .A(n70), .Z(n74) );
  BUF_X1 U11 ( .A(n411), .Z(n71) );
  BUF_X1 U12 ( .A(n70), .Z(n72) );
  BUF_X1 U13 ( .A(n70), .Z(n75) );
  BUF_X1 U14 ( .A(n417), .Z(n69) );
  NOR2_X1 U15 ( .A1(n723), .A2(n301), .ZN(n420) );
  NOR2_X1 U16 ( .A1(n423), .A2(n322), .ZN(n750) );
  INV_X1 U17 ( .A(n428), .ZN(n286) );
  AND3_X1 U18 ( .A1(n565), .A2(n307), .A3(n566), .ZN(n525) );
  INV_X1 U19 ( .A(n433), .ZN(n307) );
  INV_X1 U20 ( .A(n698), .ZN(n295) );
  AND2_X1 U21 ( .A1(n680), .A2(n681), .ZN(n664) );
  INV_X1 U22 ( .A(n708), .ZN(n243) );
  AND3_X1 U23 ( .A1(n565), .A2(n289), .A3(n566), .ZN(n517) );
  INV_X1 U24 ( .A(n424), .ZN(n289) );
  NOR3_X1 U25 ( .A1(n284), .A2(N597), .A3(n432), .ZN(n740) );
  OAI21_X1 U26 ( .B1(n377), .B2(n329), .A(n69), .ZN(n494) );
  NAND2_X1 U27 ( .A1(n324), .A2(n328), .ZN(n377) );
  NOR2_X1 U28 ( .A1(reset), .A2(n392), .ZN(wr_en_a25) );
  NOR2_X1 U29 ( .A1(reset), .A2(n384), .ZN(wr_en_a32) );
  NOR2_X1 U30 ( .A1(reset), .A2(n385), .ZN(wr_en_a31) );
  NAND2_X1 U31 ( .A1(n417), .A2(n588), .ZN(n583) );
  NAND4_X1 U32 ( .A1(n566), .A2(n300), .A3(n589), .A4(n286), .ZN(n588) );
  INV_X1 U33 ( .A(n425), .ZN(n300) );
  NOR2_X1 U34 ( .A1(reset), .A2(n401), .ZN(wr_en_a17) );
  NOR2_X1 U35 ( .A1(reset), .A2(n399), .ZN(wr_en_a19) );
  NOR2_X1 U36 ( .A1(reset), .A2(n407), .ZN(wr_en_a11) );
  NOR2_X1 U37 ( .A1(reset), .A2(n402), .ZN(wr_en_a16) );
  NOR2_X1 U38 ( .A1(reset), .A2(n393), .ZN(wr_en_a24) );
  NOR2_X1 U39 ( .A1(reset), .A2(n386), .ZN(wr_en_a30) );
  NOR2_X1 U40 ( .A1(reset), .A2(n383), .ZN(wr_en_a4) );
  NOR2_X1 U41 ( .A1(reset), .A2(n378), .ZN(wr_en_a9) );
  NAND2_X1 U42 ( .A1(n417), .A2(n621), .ZN(n616) );
  NAND4_X1 U43 ( .A1(n622), .A2(n288), .A3(n623), .A4(n402), .ZN(n621) );
  INV_X1 U44 ( .A(n442), .ZN(n288) );
  NOR2_X1 U45 ( .A1(reset), .A2(n377), .ZN(wr_en_x) );
  NOR2_X1 U46 ( .A1(reset), .A2(n398), .ZN(wr_en_a2) );
  NAND2_X1 U47 ( .A1(n417), .A2(n671), .ZN(n666) );
  NAND2_X1 U48 ( .A1(n69), .A2(n418), .ZN(n412) );
  NAND2_X1 U49 ( .A1(n69), .A2(n541), .ZN(n536) );
  NAND2_X1 U50 ( .A1(n417), .A2(n654), .ZN(n649) );
  NAND2_X1 U51 ( .A1(n417), .A2(n605), .ZN(n600) );
  NAND2_X1 U52 ( .A1(n417), .A2(n722), .ZN(n717) );
  NOR2_X1 U53 ( .A1(reset), .A2(n387), .ZN(wr_en_a3) );
  NOR2_X1 U54 ( .A1(reset), .A2(n397), .ZN(wr_en_a20) );
  NOR2_X1 U55 ( .A1(reset), .A2(n388), .ZN(wr_en_a29) );
  NOR2_X1 U56 ( .A1(reset), .A2(n400), .ZN(wr_en_a18) );
  NOR2_X1 U57 ( .A1(reset), .A2(n408), .ZN(wr_en_a10) );
  NOR2_X1 U58 ( .A1(reset), .A2(n409), .ZN(wr_en_a1) );
  NOR2_X1 U59 ( .A1(reset), .A2(n379), .ZN(wr_en_a8) );
  NOR2_X1 U60 ( .A1(reset), .A2(n396), .ZN(wr_en_a21) );
  NOR2_X1 U61 ( .A1(reset), .A2(n403), .ZN(wr_en_a15) );
  NOR2_X1 U62 ( .A1(reset), .A2(n406), .ZN(wr_en_a12) );
  NOR2_X1 U63 ( .A1(reset), .A2(n405), .ZN(wr_en_a13) );
  NOR2_X1 U64 ( .A1(reset), .A2(n404), .ZN(wr_en_a14) );
  NOR2_X1 U65 ( .A1(reset), .A2(n394), .ZN(wr_en_a23) );
  NOR2_X1 U66 ( .A1(reset), .A2(n389), .ZN(wr_en_a28) );
  NOR2_X1 U67 ( .A1(reset), .A2(n390), .ZN(wr_en_a27) );
  NOR2_X1 U68 ( .A1(reset), .A2(n382), .ZN(wr_en_a5) );
  NOR2_X1 U69 ( .A1(reset), .A2(n381), .ZN(wr_en_a6) );
  NOR2_X1 U70 ( .A1(reset), .A2(n380), .ZN(wr_en_a7) );
  NOR2_X1 U71 ( .A1(reset), .A2(n395), .ZN(wr_en_a22) );
  NOR2_X1 U72 ( .A1(reset), .A2(n391), .ZN(wr_en_a26) );
  NAND4_X1 U73 ( .A1(n589), .A2(n466), .A3(n565), .A4(n748), .ZN(n417) );
  NOR2_X1 U74 ( .A1(n749), .A2(n76), .ZN(n748) );
  NOR2_X1 U75 ( .A1(reset), .A2(n376), .ZN(wr_en_y) );
  AND3_X1 U76 ( .A1(n409), .A2(n383), .A3(n387), .ZN(n755) );
  AND3_X1 U77 ( .A1(n590), .A2(n405), .A3(n574), .ZN(n622) );
  NAND2_X1 U78 ( .A1(n386), .A2(n385), .ZN(n423) );
  NAND2_X1 U79 ( .A1(n750), .A2(n398), .ZN(n433) );
  AND3_X1 U80 ( .A1(n589), .A2(n396), .A3(n566), .ZN(n574) );
  AND3_X1 U81 ( .A1(n286), .A2(n396), .A3(n590), .ZN(n565) );
  NAND2_X1 U82 ( .A1(n383), .A2(n382), .ZN(n707) );
  INV_X1 U83 ( .A(n384), .ZN(n322) );
  NAND2_X1 U84 ( .A1(n466), .A2(n376), .ZN(N597) );
  NAND2_X1 U85 ( .A1(n417), .A2(n639), .ZN(n634) );
  NAND4_X1 U86 ( .A1(n622), .A2(n315), .A3(n632), .A4(n404), .ZN(n639) );
  INV_X1 U87 ( .A(n754), .ZN(n284) );
  NAND2_X1 U88 ( .A1(n477), .A2(n435), .ZN(n454) );
  INV_X1 U89 ( .A(n382), .ZN(n301) );
  AND2_X1 U90 ( .A1(n624), .A2(n401), .ZN(n632) );
  AND2_X1 U91 ( .A1(n395), .A2(n394), .ZN(n590) );
  AND2_X1 U92 ( .A1(n444), .A2(n393), .ZN(n526) );
  AND3_X1 U93 ( .A1(n379), .A2(n378), .A3(n381), .ZN(n681) );
  AND3_X1 U94 ( .A1(n399), .A2(n397), .A3(n400), .ZN(n624) );
  AND2_X1 U95 ( .A1(n614), .A2(n404), .ZN(n598) );
  AND2_X1 U96 ( .A1(n517), .A2(n398), .ZN(n502) );
  NAND2_X1 U97 ( .A1(n656), .A2(n405), .ZN(n428) );
  AND3_X1 U98 ( .A1(n632), .A2(n402), .A3(n623), .ZN(n656) );
  INV_X1 U99 ( .A(n378), .ZN(n290) );
  AND3_X1 U100 ( .A1(n392), .A2(n388), .A3(n525), .ZN(n542) );
  AND3_X1 U101 ( .A1(n390), .A2(n389), .A3(n391), .ZN(n444) );
  INV_X1 U102 ( .A(n403), .ZN(n314) );
  INV_X1 U103 ( .A(n396), .ZN(n299) );
  AND4_X1 U104 ( .A1(n565), .A2(n589), .A3(n739), .A4(n740), .ZN(n419) );
  NAND2_X1 U105 ( .A1(n377), .A2(n435), .ZN(N595) );
  INV_X1 U106 ( .A(n404), .ZN(n310) );
  INV_X1 U107 ( .A(n380), .ZN(n316) );
  AND3_X1 U108 ( .A1(n295), .A2(n379), .A3(n680), .ZN(n689) );
  AND3_X1 U109 ( .A1(n393), .A2(n390), .A3(n542), .ZN(n534) );
  INV_X1 U110 ( .A(N86), .ZN(n118) );
  AND4_X1 U111 ( .A1(n622), .A2(n403), .A3(n402), .A4(n401), .ZN(n614) );
  INV_X1 U112 ( .A(n409), .ZN(n319) );
  BUF_X1 U113 ( .A(n411), .Z(n70) );
  INV_X1 U114 ( .A(n476), .ZN(n296) );
  AOI211_X1 U115 ( .C1(n329), .C2(n284), .A(n306), .B(N597), .ZN(n440) );
  INV_X1 U116 ( .A(n398), .ZN(n306) );
  INV_X1 U117 ( .A(n381), .ZN(n311) );
  INV_X1 U118 ( .A(n385), .ZN(n320) );
  AOI221_X1 U119 ( .B1(N636), .B2(n285), .C1(N620), .C2(n290), .A(n443), .ZN(
        n473) );
  INV_X1 U120 ( .A(n401), .ZN(n285) );
  OAI211_X1 U121 ( .C1(n405), .C2(n332), .A(n436), .B(n474), .ZN(n443) );
  INV_X1 U122 ( .A(N628), .ZN(n332) );
  AOI221_X1 U123 ( .B1(N660), .B2(n302), .C1(N674), .C2(n475), .A(n296), .ZN(
        n474) );
  INV_X1 U124 ( .A(n388), .ZN(n302) );
  INV_X1 U125 ( .A(n481), .ZN(n328) );
  OAI221_X1 U126 ( .B1(N606), .B2(n398), .C1(n409), .C2(n335), .A(n120), .ZN(
        n470) );
  INV_X1 U127 ( .A(N604), .ZN(n335) );
  OAI221_X1 U128 ( .B1(n394), .B2(n333), .C1(N646), .C2(n395), .A(n293), .ZN(
        n460) );
  INV_X1 U129 ( .A(N648), .ZN(n333) );
  INV_X1 U130 ( .A(n461), .ZN(n293) );
  OAI22_X1 U131 ( .A1(n397), .A2(N642), .B1(n330), .B2(n399), .ZN(n461) );
  OAI21_X1 U132 ( .B1(n772), .B2(n482), .A(n455), .ZN(n432) );
  AOI22_X1 U133 ( .A1(n301), .A2(N612), .B1(n299), .B2(N644), .ZN(n436) );
  OAI21_X1 U134 ( .B1(N644), .B2(n396), .A(n590), .ZN(n425) );
  NAND2_X1 U135 ( .A1(n757), .A2(n327), .ZN(n383) );
  OAI21_X1 U136 ( .B1(N636), .B2(n401), .A(n624), .ZN(n442) );
  NAND2_X1 U137 ( .A1(n770), .A2(n756), .ZN(n399) );
  NAND2_X1 U138 ( .A1(n763), .A2(n756), .ZN(n407) );
  NAND2_X1 U139 ( .A1(n770), .A2(n324), .ZN(n402) );
  NOR2_X1 U140 ( .A1(n376), .A2(N674), .ZN(N86) );
  OAI221_X1 U141 ( .B1(N610), .B2(n383), .C1(n387), .C2(n339), .A(n478), .ZN(
        n469) );
  INV_X1 U142 ( .A(N608), .ZN(n339) );
  AOI22_X1 U143 ( .A1(N616), .A2(n316), .B1(n311), .B2(n338), .ZN(n478) );
  INV_X1 U144 ( .A(N614), .ZN(n338) );
  NAND2_X1 U145 ( .A1(n764), .A2(n761), .ZN(n392) );
  AOI21_X1 U146 ( .B1(n438), .B2(n121), .A(reset), .ZN(N82) );
  INV_X1 U147 ( .A(n439), .ZN(n121) );
  NOR3_X1 U148 ( .A1(n441), .A2(n442), .A3(n443), .ZN(n438) );
  OAI221_X1 U149 ( .B1(n392), .B2(N652), .C1(n378), .C2(N620), .A(n440), .ZN(
        n439) );
  NAND2_X1 U150 ( .A1(n69), .A2(n501), .ZN(n496) );
  INV_X1 U151 ( .A(n423), .ZN(n313) );
  NAND2_X1 U152 ( .A1(n752), .A2(n324), .ZN(n384) );
  NAND2_X1 U153 ( .A1(n768), .A2(n767), .ZN(n388) );
  NAND2_X1 U154 ( .A1(n417), .A2(n663), .ZN(n658) );
  NAND4_X1 U155 ( .A1(N626), .A2(n664), .A3(n408), .A4(n407), .ZN(n663) );
  NAND2_X1 U156 ( .A1(n417), .A2(n613), .ZN(n608) );
  NAND4_X1 U157 ( .A1(N638), .A2(n598), .A3(n399), .A4(n397), .ZN(n613) );
  NAND2_X1 U158 ( .A1(n417), .A2(n679), .ZN(n674) );
  NAND4_X1 U159 ( .A1(N622), .A2(n664), .A3(n407), .A4(n406), .ZN(n679) );
  NAND2_X1 U160 ( .A1(n417), .A2(n597), .ZN(n592) );
  NAND4_X1 U161 ( .A1(N642), .A2(n598), .A3(n400), .A4(n399), .ZN(n597) );
  NAND2_X1 U162 ( .A1(n69), .A2(n516), .ZN(n511) );
  NAND4_X1 U163 ( .A1(N662), .A2(n502), .A3(n385), .A4(n384), .ZN(n516) );
  NAND2_X1 U164 ( .A1(n417), .A2(n581), .ZN(n576) );
  NAND4_X1 U165 ( .A1(N646), .A2(n574), .A3(n286), .A4(n394), .ZN(n581) );
  NAND2_X1 U166 ( .A1(n417), .A2(n631), .ZN(n626) );
  NAND4_X1 U167 ( .A1(N634), .A2(n622), .A3(n623), .A4(n632), .ZN(n631) );
  NAND2_X1 U168 ( .A1(n69), .A2(n573), .ZN(n568) );
  NAND4_X1 U169 ( .A1(n574), .A2(N648), .A3(n286), .A4(n395), .ZN(n573) );
  NAND2_X1 U170 ( .A1(n69), .A2(n557), .ZN(n552) );
  NAND4_X1 U171 ( .A1(n525), .A2(N652), .A3(n526), .A4(n388), .ZN(n557) );
  NAND2_X1 U172 ( .A1(n69), .A2(n737), .ZN(n732) );
  NAND4_X1 U173 ( .A1(n297), .A2(N608), .A3(n738), .A4(n419), .ZN(n737) );
  INV_X1 U174 ( .A(n707), .ZN(n297) );
  NOR2_X1 U175 ( .A1(n319), .A2(n723), .ZN(n738) );
  NAND2_X1 U176 ( .A1(n69), .A2(n524), .ZN(n519) );
  NAND4_X1 U177 ( .A1(n525), .A2(N660), .A3(n526), .A4(n392), .ZN(n524) );
  NAND2_X1 U178 ( .A1(n417), .A2(n688), .ZN(n683) );
  NAND2_X1 U179 ( .A1(n69), .A2(n509), .ZN(n504) );
  NAND4_X1 U180 ( .A1(n502), .A2(N664), .A3(n386), .A4(n384), .ZN(n509) );
  NAND2_X1 U181 ( .A1(n417), .A2(n705), .ZN(n700) );
  NAND4_X1 U182 ( .A1(n295), .A2(n681), .A3(N616), .A4(n706), .ZN(n705) );
  NOR2_X1 U183 ( .A1(n707), .A2(n708), .ZN(n706) );
  NAND2_X1 U184 ( .A1(n417), .A2(n696), .ZN(n691) );
  NOR3_X1 U185 ( .A1(n698), .A2(n290), .A3(n311), .ZN(n697) );
  INV_X1 U186 ( .A(N668), .ZN(n329) );
  NAND2_X1 U187 ( .A1(n417), .A2(n715), .ZN(n710) );
  NAND2_X1 U188 ( .A1(n417), .A2(n730), .ZN(n725) );
  NAND2_X1 U189 ( .A1(n69), .A2(n550), .ZN(n545) );
  NAND2_X1 U190 ( .A1(n69), .A2(n533), .ZN(n528) );
  NAND2_X1 U191 ( .A1(n417), .A2(n647), .ZN(n642) );
  NAND2_X1 U192 ( .A1(n747), .A2(n69), .ZN(n742) );
  AOI21_X1 U193 ( .B1(n326), .B2(n301), .A(n723), .ZN(n427) );
  INV_X1 U194 ( .A(N612), .ZN(n326) );
  INV_X1 U195 ( .A(n482), .ZN(n327) );
  NAND2_X1 U196 ( .A1(n328), .A2(n756), .ZN(n376) );
  NAND2_X1 U197 ( .A1(n752), .A2(n753), .ZN(n385) );
  NAND2_X1 U198 ( .A1(n327), .A2(n756), .ZN(n387) );
  NAND2_X1 U199 ( .A1(n753), .A2(n328), .ZN(n409) );
  INV_X1 U200 ( .A(n746), .ZN(n137) );
  AOI22_X1 U201 ( .A1(addr_a2[0]), .A2(n76), .B1(n35), .B2(n742), .ZN(n746) );
  INV_X1 U202 ( .A(n772), .ZN(n324) );
  NAND2_X1 U203 ( .A1(n770), .A2(n761), .ZN(n401) );
  NAND2_X1 U204 ( .A1(n768), .A2(n769), .ZN(n394) );
  INV_X1 U205 ( .A(n490), .ZN(n119) );
  INV_X1 U206 ( .A(n736), .ZN(n228) );
  AOI22_X1 U207 ( .A1(addr_a3[0]), .A2(n75), .B1(n36), .B2(n732), .ZN(n736) );
  INV_X1 U208 ( .A(n515), .ZN(n122) );
  AOI22_X1 U209 ( .A1(addr_a30[0]), .A2(n70), .B1(n37), .B2(n511), .ZN(n515)
         );
  INV_X1 U210 ( .A(n508), .ZN(n127) );
  AOI22_X1 U211 ( .A1(addr_a31[0]), .A2(n75), .B1(n38), .B2(n504), .ZN(n508)
         );
  INV_X1 U212 ( .A(n563), .ZN(n207) );
  AOI22_X1 U213 ( .A1(addr_a24[0]), .A2(n73), .B1(n39), .B2(n559), .ZN(n563)
         );
  INV_X1 U214 ( .A(n540), .ZN(n212) );
  AOI22_X1 U215 ( .A1(addr_a27[0]), .A2(n70), .B1(n40), .B2(n536), .ZN(n540)
         );
  INV_X1 U216 ( .A(n523), .ZN(n222) );
  AOI22_X1 U217 ( .A1(addr_a29[0]), .A2(n75), .B1(n41), .B2(n519), .ZN(n523)
         );
  INV_X1 U218 ( .A(n572), .ZN(n182) );
  AOI22_X1 U219 ( .A1(addr_a23[0]), .A2(n73), .B1(n42), .B2(n568), .ZN(n572)
         );
  INV_X1 U220 ( .A(n500), .ZN(n132) );
  AOI22_X1 U221 ( .A1(addr_a32[0]), .A2(n71), .B1(n43), .B2(n496), .ZN(n500)
         );
  INV_X1 U222 ( .A(n556), .ZN(n217) );
  AOI22_X1 U223 ( .A1(addr_a25[0]), .A2(n72), .B1(n44), .B2(n552), .ZN(n556)
         );
  INV_X1 U224 ( .A(n416), .ZN(n279) );
  AOI22_X1 U225 ( .A1(addr_a1[0]), .A2(n71), .B1(n45), .B2(n412), .ZN(n416) );
  INV_X1 U226 ( .A(n587), .ZN(n192) );
  AOI22_X1 U227 ( .A1(addr_a21[0]), .A2(n74), .B1(n46), .B2(n583), .ZN(n587)
         );
  INV_X1 U228 ( .A(n580), .ZN(n177) );
  AOI22_X1 U229 ( .A1(addr_a22[0]), .A2(n73), .B1(n47), .B2(n576), .ZN(n580)
         );
  INV_X1 U230 ( .A(n653), .ZN(n187) );
  AOI22_X1 U231 ( .A1(addr_a13[0]), .A2(n73), .B1(n48), .B2(n649), .ZN(n653)
         );
  NAND2_X1 U232 ( .A1(n757), .A2(n763), .ZN(n406) );
  INV_X1 U233 ( .A(n489), .ZN(n113) );
  AOI22_X1 U234 ( .A1(addr_y[0]), .A2(n485), .B1(n49), .B2(n119), .ZN(n489) );
  NAND2_X1 U235 ( .A1(n770), .A2(n757), .ZN(n397) );
  NAND2_X1 U236 ( .A1(n751), .A2(n327), .ZN(n398) );
  NAND2_X1 U237 ( .A1(n762), .A2(n763), .ZN(n405) );
  NAND2_X1 U238 ( .A1(n764), .A2(n324), .ZN(n393) );
  INV_X1 U239 ( .A(n640), .ZN(n315) );
  OAI21_X1 U240 ( .B1(N632), .B2(n403), .A(n402), .ZN(n640) );
  NAND2_X1 U241 ( .A1(n752), .A2(n492), .ZN(n386) );
  NAND2_X1 U242 ( .A1(n763), .A2(n761), .ZN(n378) );
  NAND2_X1 U243 ( .A1(n751), .A2(n763), .ZN(n408) );
  NAND2_X1 U244 ( .A1(n751), .A2(n770), .ZN(n400) );
  NAND2_X1 U245 ( .A1(n761), .A2(n328), .ZN(n754) );
  NAND2_X1 U246 ( .A1(n763), .A2(n324), .ZN(n379) );
  NAND2_X1 U247 ( .A1(n770), .A2(n762), .ZN(n396) );
  NAND2_X1 U248 ( .A1(n765), .A2(n767), .ZN(n389) );
  NAND2_X1 U249 ( .A1(n768), .A2(n766), .ZN(n390) );
  NAND2_X1 U250 ( .A1(n770), .A2(n753), .ZN(n403) );
  NAND2_X1 U251 ( .A1(n69), .A2(n564), .ZN(n559) );
  NAND2_X1 U252 ( .A1(n770), .A2(n492), .ZN(n404) );
  NAND2_X1 U253 ( .A1(n765), .A2(n769), .ZN(n395) );
  NAND2_X1 U254 ( .A1(n765), .A2(n766), .ZN(n391) );
  NAND2_X1 U255 ( .A1(n327), .A2(n753), .ZN(n435) );
  NAND2_X1 U256 ( .A1(n753), .A2(n763), .ZN(n380) );
  NAND2_X1 U257 ( .A1(n492), .A2(n763), .ZN(n381) );
  NAND2_X1 U258 ( .A1(n327), .A2(n762), .ZN(n382) );
  NAND2_X1 U259 ( .A1(n327), .A2(n492), .ZN(n466) );
  NAND4_X1 U260 ( .A1(n120), .A2(n303), .A3(n294), .A4(n315), .ZN(n450) );
  AOI21_X1 U261 ( .B1(n426), .B2(n427), .A(reset), .ZN(N84) );
  AOI21_X1 U262 ( .B1(N644), .B2(n299), .A(n428), .ZN(n426) );
  AOI21_X1 U263 ( .B1(n456), .B2(n457), .A(reset), .ZN(N80) );
  NOR4_X1 U264 ( .A1(n111), .A2(n458), .A3(n459), .A4(n460), .ZN(n457) );
  NOR4_X1 U265 ( .A1(n467), .A2(n468), .A3(n469), .A4(n470), .ZN(n456) );
  OAI221_X1 U266 ( .B1(N658), .B2(n389), .C1(n390), .C2(n334), .A(n309), .ZN(
        n459) );
  NAND2_X1 U267 ( .A1(n751), .A2(n328), .ZN(n455) );
  INV_X1 U268 ( .A(n766), .ZN(n308) );
  INV_X1 U269 ( .A(N640), .ZN(n330) );
  NAND2_X1 U270 ( .A1(n757), .A2(n328), .ZN(n476) );
  INV_X1 U271 ( .A(N674), .ZN(n112) );
  NAND2_X1 U272 ( .A1(n492), .A2(n328), .ZN(n477) );
  AND2_X1 U273 ( .A1(n762), .A2(n328), .ZN(n475) );
  INV_X1 U274 ( .A(n445), .ZN(n298) );
  OAI211_X1 U275 ( .C1(N604), .C2(n409), .A(n387), .B(n383), .ZN(n445) );
  NOR2_X1 U276 ( .A1(reset), .A2(n429), .ZN(N83) );
  NOR4_X1 U277 ( .A1(n430), .A2(n431), .A3(n432), .A4(n433), .ZN(n429) );
  OAI221_X1 U278 ( .B1(N668), .B2(n377), .C1(N660), .C2(n388), .A(n434), .ZN(
        n431) );
  NAND4_X1 U279 ( .A1(n287), .A2(n436), .A3(n298), .A4(n291), .ZN(n430) );
  NOR2_X1 U280 ( .A1(reset), .A2(n446), .ZN(N81) );
  NOR4_X1 U281 ( .A1(n447), .A2(n448), .A3(n449), .A4(n450), .ZN(n446) );
  OAI211_X1 U282 ( .C1(N608), .C2(n387), .A(n292), .B(n317), .ZN(n449) );
  NAND4_X1 U283 ( .A1(n455), .A2(n383), .A3(n379), .A4(n118), .ZN(n447) );
  AND4_X1 U284 ( .A1(n477), .A2(n318), .A3(n476), .A4(n758), .ZN(n739) );
  NOR2_X1 U285 ( .A1(n475), .A2(n437), .ZN(n758) );
  INV_X1 U286 ( .A(N595), .ZN(n318) );
  INV_X1 U287 ( .A(n543), .ZN(n303) );
  OAI211_X1 U288 ( .C1(N656), .C2(n390), .A(n393), .B(n389), .ZN(n543) );
  INV_X1 U289 ( .A(n672), .ZN(n294) );
  OAI21_X1 U290 ( .B1(N624), .B2(n407), .A(n406), .ZN(n672) );
  INV_X1 U291 ( .A(n606), .ZN(n292) );
  OAI21_X1 U292 ( .B1(N640), .B2(n399), .A(n397), .ZN(n606) );
  INV_X1 U293 ( .A(n655), .ZN(n287) );
  OAI21_X1 U294 ( .B1(N628), .B2(n405), .A(n656), .ZN(n655) );
  OAI211_X1 U295 ( .C1(N668), .C2(n754), .A(n376), .B(n304), .ZN(n411) );
  INV_X1 U296 ( .A(n432), .ZN(n304) );
  AND2_X1 U297 ( .A1(N572), .A2(n494), .ZN(N577) );
  AND2_X1 U298 ( .A1(N571), .A2(n494), .ZN(N576) );
  AND2_X1 U299 ( .A1(N570), .A2(n494), .ZN(N575) );
  AND2_X1 U300 ( .A1(n68), .A2(n494), .ZN(N574) );
  INV_X1 U301 ( .A(n714), .ZN(n244) );
  AOI22_X1 U302 ( .A1(addr_a6[0]), .A2(n70), .B1(n50), .B2(n710), .ZN(n714) );
  INV_X1 U303 ( .A(n687), .ZN(n249) );
  AOI22_X1 U304 ( .A1(addr_a9[0]), .A2(n73), .B1(n51), .B2(n683), .ZN(n687) );
  INV_X1 U305 ( .A(n678), .ZN(n254) );
  AOI22_X1 U306 ( .A1(addr_a10[0]), .A2(n74), .B1(n52), .B2(n674), .ZN(n678)
         );
  INV_X1 U307 ( .A(n662), .ZN(n259) );
  AOI22_X1 U308 ( .A1(addr_a12[0]), .A2(n74), .B1(n53), .B2(n658), .ZN(n662)
         );
  INV_X1 U309 ( .A(n670), .ZN(n264) );
  AOI22_X1 U310 ( .A1(addr_a11[0]), .A2(n71), .B1(n54), .B2(n666), .ZN(n670)
         );
  INV_X1 U311 ( .A(n695), .ZN(n269) );
  AOI22_X1 U312 ( .A1(addr_a8[0]), .A2(n74), .B1(n55), .B2(n691), .ZN(n695) );
  INV_X1 U313 ( .A(n704), .ZN(n274) );
  AOI22_X1 U314 ( .A1(addr_a7[0]), .A2(n70), .B1(n56), .B2(n700), .ZN(n704) );
  INV_X1 U315 ( .A(n729), .ZN(n233) );
  AOI22_X1 U316 ( .A1(addr_a4[0]), .A2(n75), .B1(n57), .B2(n725), .ZN(n729) );
  INV_X1 U317 ( .A(n549), .ZN(n197) );
  AOI22_X1 U318 ( .A1(addr_a26[0]), .A2(n72), .B1(n58), .B2(n545), .ZN(n549)
         );
  INV_X1 U319 ( .A(n532), .ZN(n202) );
  AOI22_X1 U320 ( .A1(addr_a28[0]), .A2(n70), .B1(n59), .B2(n528), .ZN(n532)
         );
  INV_X1 U321 ( .A(n638), .ZN(n162) );
  AOI22_X1 U322 ( .A1(addr_a15[0]), .A2(n73), .B1(n60), .B2(n634), .ZN(n638)
         );
  INV_X1 U323 ( .A(n630), .ZN(n167) );
  AOI22_X1 U324 ( .A1(addr_a16[0]), .A2(n74), .B1(n61), .B2(n626), .ZN(n630)
         );
  INV_X1 U325 ( .A(n620), .ZN(n172) );
  AOI22_X1 U326 ( .A1(addr_a17[0]), .A2(n73), .B1(n62), .B2(n616), .ZN(n620)
         );
  INV_X1 U327 ( .A(n646), .ZN(n157) );
  AOI22_X1 U328 ( .A1(addr_a14[0]), .A2(n74), .B1(n63), .B2(n642), .ZN(n646)
         );
  INV_X1 U329 ( .A(n612), .ZN(n142) );
  AOI22_X1 U330 ( .A1(addr_a18[0]), .A2(n73), .B1(n64), .B2(n608), .ZN(n612)
         );
  INV_X1 U331 ( .A(n604), .ZN(n152) );
  AOI22_X1 U332 ( .A1(addr_a19[0]), .A2(n71), .B1(n65), .B2(n600), .ZN(n604)
         );
  INV_X1 U333 ( .A(n596), .ZN(n147) );
  AOI22_X1 U334 ( .A1(addr_a20[0]), .A2(n74), .B1(n66), .B2(n592), .ZN(n596)
         );
  INV_X1 U335 ( .A(n721), .ZN(n238) );
  AOI22_X1 U336 ( .A1(addr_a5[0]), .A2(n75), .B1(n67), .B2(n717), .ZN(n721) );
  OAI221_X1 U337 ( .B1(N626), .B2(n406), .C1(n407), .C2(n337), .A(n305), .ZN(
        n468) );
  INV_X1 U338 ( .A(N624), .ZN(n337) );
  INV_X1 U339 ( .A(n479), .ZN(n305) );
  OAI22_X1 U340 ( .A1(n408), .A2(N622), .B1(n379), .B2(N618), .ZN(n479) );
  OAI221_X1 U341 ( .B1(n385), .B2(n336), .C1(N662), .C2(n386), .A(n323), .ZN(
        n458) );
  INV_X1 U342 ( .A(n463), .ZN(n323) );
  OAI22_X1 U343 ( .A1(n377), .A2(N668), .B1(n384), .B2(N666), .ZN(n463) );
  OAI221_X1 U344 ( .B1(N638), .B2(n400), .C1(N634), .C2(n402), .A(n480), .ZN(
        n467) );
  AOI22_X1 U345 ( .A1(N632), .A2(n314), .B1(n310), .B2(n331), .ZN(n480) );
  INV_X1 U346 ( .A(N630), .ZN(n331) );
  INV_X1 U347 ( .A(N664), .ZN(n336) );
  AOI21_X1 U348 ( .B1(n421), .B2(n422), .A(reset), .ZN(N85) );
  AOI21_X1 U349 ( .B1(N666), .B2(n322), .A(n423), .ZN(n422) );
  NOR2_X1 U350 ( .A1(n424), .A2(n425), .ZN(n421) );
  INV_X1 U351 ( .A(N656), .ZN(n334) );
  INV_X1 U352 ( .A(n437), .ZN(n291) );
  INV_X1 U353 ( .A(n451), .ZN(n317) );
  OAI22_X1 U354 ( .A1(n394), .A2(N648), .B1(n380), .B2(N616), .ZN(n451) );
  INV_X1 U355 ( .A(n462), .ZN(n309) );
  OAI22_X1 U356 ( .A1(n391), .A2(N654), .B1(n393), .B2(N650), .ZN(n462) );
  NOR3_X1 U357 ( .A1(state[3]), .A2(state[4]), .A3(n321), .ZN(n764) );
  NOR3_X1 U358 ( .A1(n355), .A2(state[4]), .A3(n321), .ZN(n752) );
  NOR2_X1 U359 ( .A1(n360), .A2(n308), .ZN(n756) );
  NOR2_X1 U360 ( .A1(n308), .A2(state[0]), .ZN(n751) );
  AND2_X1 U361 ( .A1(state[4]), .A2(n771), .ZN(n763) );
  INV_X1 U362 ( .A(n464), .ZN(n111) );
  AOI211_X1 U363 ( .C1(n454), .C2(loadMatrix), .A(n312), .B(n465), .ZN(n464)
         );
  INV_X1 U364 ( .A(n466), .ZN(n312) );
  OAI22_X1 U365 ( .A1(n112), .A2(n376), .B1(n435), .B2(loadVector), .ZN(n465)
         );
  AND2_X1 U366 ( .A1(n773), .A2(state[4]), .ZN(n770) );
  NOR2_X1 U367 ( .A1(n359), .A2(n358), .ZN(n767) );
  NOR2_X1 U368 ( .A1(state[2]), .A2(state[1]), .ZN(n769) );
  NOR2_X1 U369 ( .A1(n358), .A2(state[1]), .ZN(n766) );
  OAI21_X1 U370 ( .B1(n759), .B2(n321), .A(n760), .ZN(n437) );
  AOI21_X1 U371 ( .B1(state[3]), .B2(state[2]), .A(state[4]), .ZN(n759) );
  AND2_X1 U372 ( .A1(n769), .A2(n360), .ZN(n492) );
  AND3_X1 U373 ( .A1(n490), .A2(n118), .A3(n491), .ZN(n485) );
  INV_X1 U374 ( .A(n744), .ZN(n139) );
  AOI22_X1 U375 ( .A1(addr_a2[2]), .A2(n76), .B1(N107), .B2(n742), .ZN(n744)
         );
  INV_X1 U376 ( .A(n745), .ZN(n138) );
  AOI22_X1 U377 ( .A1(addr_a2[1]), .A2(n76), .B1(N106), .B2(n742), .ZN(n745)
         );
  INV_X1 U378 ( .A(n731), .ZN(n232) );
  AOI22_X1 U379 ( .A1(addr_a3[4]), .A2(n75), .B1(N124), .B2(n732), .ZN(n731)
         );
  INV_X1 U380 ( .A(n510), .ZN(n126) );
  AOI22_X1 U381 ( .A1(addr_a30[4]), .A2(n70), .B1(N529), .B2(n511), .ZN(n510)
         );
  INV_X1 U382 ( .A(n503), .ZN(n131) );
  AOI22_X1 U383 ( .A1(addr_a31[4]), .A2(n71), .B1(N544), .B2(n504), .ZN(n503)
         );
  INV_X1 U384 ( .A(n410), .ZN(n283) );
  AOI22_X1 U385 ( .A1(addr_a1[4]), .A2(n71), .B1(N94), .B2(n412), .ZN(n410) );
  INV_X1 U386 ( .A(n535), .ZN(n216) );
  AOI22_X1 U387 ( .A1(addr_a27[4]), .A2(n70), .B1(N484), .B2(n536), .ZN(n535)
         );
  INV_X1 U388 ( .A(n518), .ZN(n226) );
  AOI22_X1 U389 ( .A1(addr_a29[4]), .A2(n75), .B1(N514), .B2(n519), .ZN(n518)
         );
  INV_X1 U390 ( .A(n582), .ZN(n196) );
  AOI22_X1 U391 ( .A1(addr_a21[4]), .A2(n74), .B1(N394), .B2(n583), .ZN(n582)
         );
  INV_X1 U392 ( .A(n575), .ZN(n181) );
  AOI22_X1 U393 ( .A1(addr_a22[4]), .A2(n73), .B1(N409), .B2(n576), .ZN(n575)
         );
  INV_X1 U394 ( .A(n567), .ZN(n186) );
  AOI22_X1 U395 ( .A1(addr_a23[4]), .A2(n73), .B1(N424), .B2(n568), .ZN(n567)
         );
  INV_X1 U396 ( .A(n648), .ZN(n191) );
  AOI22_X1 U397 ( .A1(addr_a13[4]), .A2(n411), .B1(N274), .B2(n649), .ZN(n648)
         );
  INV_X1 U398 ( .A(n495), .ZN(n136) );
  AOI22_X1 U399 ( .A1(addr_a32[4]), .A2(n71), .B1(N559), .B2(n496), .ZN(n495)
         );
  INV_X1 U400 ( .A(n551), .ZN(n221) );
  AOI22_X1 U401 ( .A1(addr_a25[4]), .A2(n72), .B1(N454), .B2(n552), .ZN(n551)
         );
  INV_X1 U402 ( .A(n734), .ZN(n230) );
  AOI22_X1 U403 ( .A1(addr_a3[2]), .A2(n75), .B1(N122), .B2(n732), .ZN(n734)
         );
  INV_X1 U404 ( .A(n735), .ZN(n229) );
  AOI22_X1 U405 ( .A1(addr_a3[1]), .A2(n75), .B1(N121), .B2(n732), .ZN(n735)
         );
  INV_X1 U406 ( .A(n506), .ZN(n129) );
  AOI22_X1 U407 ( .A1(addr_a31[2]), .A2(n75), .B1(N542), .B2(n504), .ZN(n506)
         );
  INV_X1 U408 ( .A(n507), .ZN(n128) );
  AOI22_X1 U409 ( .A1(addr_a31[1]), .A2(n70), .B1(N541), .B2(n504), .ZN(n507)
         );
  INV_X1 U410 ( .A(n521), .ZN(n224) );
  AOI22_X1 U411 ( .A1(addr_a29[2]), .A2(n75), .B1(N512), .B2(n519), .ZN(n521)
         );
  INV_X1 U412 ( .A(n522), .ZN(n223) );
  AOI22_X1 U413 ( .A1(addr_a29[1]), .A2(n75), .B1(N511), .B2(n519), .ZN(n522)
         );
  INV_X1 U414 ( .A(n570), .ZN(n184) );
  AOI22_X1 U415 ( .A1(addr_a23[2]), .A2(n73), .B1(N422), .B2(n568), .ZN(n570)
         );
  INV_X1 U416 ( .A(n571), .ZN(n183) );
  AOI22_X1 U417 ( .A1(addr_a23[1]), .A2(n73), .B1(N421), .B2(n568), .ZN(n571)
         );
  INV_X1 U418 ( .A(n498), .ZN(n134) );
  AOI22_X1 U419 ( .A1(addr_a32[2]), .A2(n71), .B1(N557), .B2(n496), .ZN(n498)
         );
  INV_X1 U420 ( .A(n499), .ZN(n133) );
  AOI22_X1 U421 ( .A1(addr_a32[1]), .A2(n71), .B1(N556), .B2(n496), .ZN(n499)
         );
  INV_X1 U422 ( .A(n555), .ZN(n218) );
  AOI22_X1 U423 ( .A1(addr_a25[1]), .A2(n72), .B1(N451), .B2(n552), .ZN(n555)
         );
  INV_X1 U424 ( .A(n554), .ZN(n219) );
  AOI22_X1 U425 ( .A1(addr_a25[2]), .A2(n72), .B1(N452), .B2(n552), .ZN(n554)
         );
  INV_X1 U426 ( .A(n414), .ZN(n281) );
  AOI22_X1 U427 ( .A1(addr_a1[2]), .A2(n71), .B1(N92), .B2(n412), .ZN(n414) );
  INV_X1 U428 ( .A(n415), .ZN(n280) );
  AOI22_X1 U429 ( .A1(addr_a1[1]), .A2(n71), .B1(N91), .B2(n412), .ZN(n415) );
  INV_X1 U430 ( .A(n585), .ZN(n194) );
  AOI22_X1 U431 ( .A1(addr_a21[2]), .A2(n74), .B1(N392), .B2(n583), .ZN(n585)
         );
  INV_X1 U432 ( .A(n586), .ZN(n193) );
  AOI22_X1 U433 ( .A1(addr_a21[1]), .A2(n74), .B1(N391), .B2(n583), .ZN(n586)
         );
  INV_X1 U434 ( .A(n578), .ZN(n179) );
  AOI22_X1 U435 ( .A1(addr_a22[2]), .A2(n73), .B1(N407), .B2(n576), .ZN(n578)
         );
  INV_X1 U436 ( .A(n579), .ZN(n178) );
  AOI22_X1 U437 ( .A1(addr_a22[1]), .A2(n73), .B1(N406), .B2(n576), .ZN(n579)
         );
  INV_X1 U438 ( .A(n651), .ZN(n189) );
  AOI22_X1 U439 ( .A1(addr_a13[2]), .A2(n71), .B1(N272), .B2(n649), .ZN(n651)
         );
  INV_X1 U440 ( .A(n652), .ZN(n188) );
  AOI22_X1 U441 ( .A1(addr_a13[1]), .A2(n72), .B1(N271), .B2(n649), .ZN(n652)
         );
  AND2_X1 U442 ( .A1(n769), .A2(state[0]), .ZN(n753) );
  OAI211_X1 U443 ( .C1(n377), .C2(n329), .A(n452), .B(n453), .ZN(n448) );
  AOI22_X1 U444 ( .A1(N666), .A2(n322), .B1(n320), .B2(n336), .ZN(n453) );
  INV_X1 U445 ( .A(loadMatrix), .ZN(n340) );
  OAI21_X1 U446 ( .B1(N86), .B2(n360), .A(n359), .ZN(n493) );
  AND2_X1 U447 ( .A1(n767), .A2(n360), .ZN(n757) );
  NOR2_X1 U448 ( .A1(state[5]), .A2(state[3]), .ZN(n771) );
  NOR2_X1 U449 ( .A1(n355), .A2(state[5]), .ZN(n773) );
  AND2_X1 U450 ( .A1(n767), .A2(state[0]), .ZN(n762) );
  NAND2_X1 U451 ( .A1(n773), .A2(n354), .ZN(n482) );
  AND2_X1 U452 ( .A1(n764), .A2(state[0]), .ZN(n768) );
  AND2_X1 U453 ( .A1(n764), .A2(n360), .ZN(n765) );
  NAND2_X1 U454 ( .A1(n771), .A2(n354), .ZN(n481) );
  INV_X1 U455 ( .A(n471), .ZN(n120) );
  OAI211_X1 U456 ( .C1(n392), .C2(n325), .A(n472), .B(n473), .ZN(n471) );
  INV_X1 U457 ( .A(N652), .ZN(n325) );
  AOI22_X1 U458 ( .A1(start), .A2(n454), .B1(N668), .B2(n284), .ZN(n472) );
  INV_X1 U459 ( .A(n733), .ZN(n231) );
  AOI22_X1 U460 ( .A1(addr_a3[3]), .A2(n75), .B1(N123), .B2(n732), .ZN(n733)
         );
  INV_X1 U461 ( .A(n711), .ZN(n247) );
  AOI22_X1 U462 ( .A1(addr_a6[3]), .A2(n70), .B1(N168), .B2(n710), .ZN(n711)
         );
  INV_X1 U463 ( .A(n684), .ZN(n252) );
  AOI22_X1 U464 ( .A1(addr_a9[3]), .A2(n71), .B1(N213), .B2(n683), .ZN(n684)
         );
  INV_X1 U465 ( .A(n675), .ZN(n257) );
  AOI22_X1 U466 ( .A1(addr_a10[3]), .A2(n411), .B1(N228), .B2(n674), .ZN(n675)
         );
  INV_X1 U467 ( .A(n659), .ZN(n262) );
  AOI22_X1 U468 ( .A1(addr_a12[3]), .A2(n70), .B1(N258), .B2(n658), .ZN(n659)
         );
  INV_X1 U469 ( .A(n667), .ZN(n267) );
  AOI22_X1 U470 ( .A1(addr_a11[3]), .A2(n71), .B1(N243), .B2(n666), .ZN(n667)
         );
  INV_X1 U471 ( .A(n692), .ZN(n272) );
  AOI22_X1 U472 ( .A1(addr_a8[3]), .A2(n72), .B1(N198), .B2(n691), .ZN(n692)
         );
  INV_X1 U473 ( .A(n701), .ZN(n277) );
  AOI22_X1 U474 ( .A1(addr_a7[3]), .A2(n72), .B1(N183), .B2(n700), .ZN(n701)
         );
  INV_X1 U475 ( .A(n512), .ZN(n125) );
  AOI22_X1 U476 ( .A1(addr_a30[3]), .A2(n75), .B1(N528), .B2(n511), .ZN(n512)
         );
  INV_X1 U477 ( .A(n505), .ZN(n130) );
  AOI22_X1 U478 ( .A1(addr_a31[3]), .A2(n71), .B1(N543), .B2(n504), .ZN(n505)
         );
  INV_X1 U479 ( .A(n726), .ZN(n236) );
  AOI22_X1 U480 ( .A1(addr_a4[3]), .A2(n75), .B1(N138), .B2(n725), .ZN(n726)
         );
  INV_X1 U481 ( .A(n413), .ZN(n282) );
  AOI22_X1 U482 ( .A1(addr_a1[3]), .A2(n71), .B1(N93), .B2(n412), .ZN(n413) );
  INV_X1 U483 ( .A(n546), .ZN(n200) );
  AOI22_X1 U484 ( .A1(addr_a26[3]), .A2(n72), .B1(N468), .B2(n545), .ZN(n546)
         );
  INV_X1 U485 ( .A(n529), .ZN(n205) );
  AOI22_X1 U486 ( .A1(addr_a28[3]), .A2(n75), .B1(N498), .B2(n528), .ZN(n529)
         );
  INV_X1 U487 ( .A(n560), .ZN(n210) );
  AOI22_X1 U488 ( .A1(addr_a24[3]), .A2(n72), .B1(N438), .B2(n559), .ZN(n560)
         );
  INV_X1 U489 ( .A(n537), .ZN(n215) );
  AOI22_X1 U490 ( .A1(addr_a27[3]), .A2(n75), .B1(N483), .B2(n536), .ZN(n537)
         );
  INV_X1 U491 ( .A(n520), .ZN(n225) );
  AOI22_X1 U492 ( .A1(addr_a29[3]), .A2(n75), .B1(N513), .B2(n519), .ZN(n520)
         );
  INV_X1 U493 ( .A(n584), .ZN(n195) );
  AOI22_X1 U494 ( .A1(addr_a21[3]), .A2(n74), .B1(N393), .B2(n583), .ZN(n584)
         );
  INV_X1 U495 ( .A(n577), .ZN(n180) );
  AOI22_X1 U496 ( .A1(addr_a22[3]), .A2(n73), .B1(N408), .B2(n576), .ZN(n577)
         );
  INV_X1 U497 ( .A(n569), .ZN(n185) );
  AOI22_X1 U498 ( .A1(addr_a23[3]), .A2(n73), .B1(N423), .B2(n568), .ZN(n569)
         );
  INV_X1 U499 ( .A(n650), .ZN(n190) );
  AOI22_X1 U500 ( .A1(addr_a13[3]), .A2(n71), .B1(N273), .B2(n649), .ZN(n650)
         );
  INV_X1 U501 ( .A(n635), .ZN(n165) );
  AOI22_X1 U502 ( .A1(addr_a15[3]), .A2(n72), .B1(N303), .B2(n634), .ZN(n635)
         );
  INV_X1 U503 ( .A(n627), .ZN(n170) );
  AOI22_X1 U504 ( .A1(addr_a16[3]), .A2(n70), .B1(N318), .B2(n626), .ZN(n627)
         );
  INV_X1 U505 ( .A(n617), .ZN(n175) );
  AOI22_X1 U506 ( .A1(addr_a17[3]), .A2(n73), .B1(N333), .B2(n616), .ZN(n617)
         );
  INV_X1 U507 ( .A(n643), .ZN(n160) );
  AOI22_X1 U508 ( .A1(addr_a14[3]), .A2(n72), .B1(N288), .B2(n642), .ZN(n643)
         );
  INV_X1 U509 ( .A(n609), .ZN(n145) );
  AOI22_X1 U510 ( .A1(addr_a18[3]), .A2(n71), .B1(N348), .B2(n608), .ZN(n609)
         );
  INV_X1 U511 ( .A(n601), .ZN(n155) );
  AOI22_X1 U512 ( .A1(addr_a19[3]), .A2(n74), .B1(N363), .B2(n600), .ZN(n601)
         );
  INV_X1 U513 ( .A(n593), .ZN(n150) );
  AOI22_X1 U514 ( .A1(addr_a20[3]), .A2(n74), .B1(N378), .B2(n592), .ZN(n593)
         );
  INV_X1 U515 ( .A(n497), .ZN(n135) );
  AOI22_X1 U516 ( .A1(addr_a32[3]), .A2(n71), .B1(N558), .B2(n496), .ZN(n497)
         );
  INV_X1 U517 ( .A(n718), .ZN(n241) );
  AOI22_X1 U518 ( .A1(addr_a5[3]), .A2(n70), .B1(N153), .B2(n717), .ZN(n718)
         );
  INV_X1 U519 ( .A(n743), .ZN(n140) );
  AOI22_X1 U520 ( .A1(addr_a2[3]), .A2(n76), .B1(N108), .B2(n742), .ZN(n743)
         );
  INV_X1 U521 ( .A(n553), .ZN(n220) );
  AOI22_X1 U522 ( .A1(addr_a25[3]), .A2(n72), .B1(N453), .B2(n552), .ZN(n553)
         );
  INV_X1 U523 ( .A(n709), .ZN(n248) );
  AOI22_X1 U524 ( .A1(addr_a6[4]), .A2(n70), .B1(N169), .B2(n710), .ZN(n709)
         );
  INV_X1 U525 ( .A(n682), .ZN(n253) );
  AOI22_X1 U526 ( .A1(addr_a9[4]), .A2(n71), .B1(N214), .B2(n683), .ZN(n682)
         );
  INV_X1 U527 ( .A(n673), .ZN(n258) );
  AOI22_X1 U528 ( .A1(addr_a10[4]), .A2(n72), .B1(N229), .B2(n674), .ZN(n673)
         );
  INV_X1 U529 ( .A(n657), .ZN(n263) );
  AOI22_X1 U530 ( .A1(addr_a12[4]), .A2(n73), .B1(N259), .B2(n658), .ZN(n657)
         );
  INV_X1 U531 ( .A(n665), .ZN(n268) );
  AOI22_X1 U532 ( .A1(addr_a11[4]), .A2(n73), .B1(N244), .B2(n666), .ZN(n665)
         );
  INV_X1 U533 ( .A(n690), .ZN(n273) );
  AOI22_X1 U534 ( .A1(addr_a8[4]), .A2(n72), .B1(N199), .B2(n691), .ZN(n690)
         );
  INV_X1 U535 ( .A(n699), .ZN(n278) );
  AOI22_X1 U536 ( .A1(addr_a7[4]), .A2(n73), .B1(N184), .B2(n700), .ZN(n699)
         );
  INV_X1 U537 ( .A(n724), .ZN(n237) );
  AOI22_X1 U538 ( .A1(addr_a4[4]), .A2(n75), .B1(N139), .B2(n725), .ZN(n724)
         );
  INV_X1 U539 ( .A(n544), .ZN(n201) );
  AOI22_X1 U540 ( .A1(addr_a26[4]), .A2(n75), .B1(N469), .B2(n545), .ZN(n544)
         );
  INV_X1 U541 ( .A(n527), .ZN(n206) );
  AOI22_X1 U542 ( .A1(addr_a28[4]), .A2(n70), .B1(N499), .B2(n528), .ZN(n527)
         );
  INV_X1 U543 ( .A(n558), .ZN(n211) );
  AOI22_X1 U544 ( .A1(addr_a24[4]), .A2(n72), .B1(N439), .B2(n559), .ZN(n558)
         );
  INV_X1 U545 ( .A(n633), .ZN(n166) );
  AOI22_X1 U546 ( .A1(addr_a15[4]), .A2(n411), .B1(N304), .B2(n634), .ZN(n633)
         );
  INV_X1 U547 ( .A(n625), .ZN(n171) );
  AOI22_X1 U548 ( .A1(addr_a16[4]), .A2(n72), .B1(N319), .B2(n626), .ZN(n625)
         );
  INV_X1 U549 ( .A(n615), .ZN(n176) );
  AOI22_X1 U550 ( .A1(addr_a17[4]), .A2(n72), .B1(N334), .B2(n616), .ZN(n615)
         );
  INV_X1 U551 ( .A(n641), .ZN(n161) );
  AOI22_X1 U552 ( .A1(addr_a14[4]), .A2(n73), .B1(N289), .B2(n642), .ZN(n641)
         );
  INV_X1 U553 ( .A(n607), .ZN(n146) );
  AOI22_X1 U554 ( .A1(addr_a18[4]), .A2(n73), .B1(N349), .B2(n608), .ZN(n607)
         );
  INV_X1 U555 ( .A(n599), .ZN(n156) );
  AOI22_X1 U556 ( .A1(addr_a19[4]), .A2(n74), .B1(N364), .B2(n600), .ZN(n599)
         );
  INV_X1 U557 ( .A(n591), .ZN(n151) );
  AOI22_X1 U558 ( .A1(addr_a20[4]), .A2(n74), .B1(N379), .B2(n592), .ZN(n591)
         );
  INV_X1 U559 ( .A(n716), .ZN(n242) );
  AOI22_X1 U560 ( .A1(addr_a5[4]), .A2(n70), .B1(N154), .B2(n717), .ZN(n716)
         );
  INV_X1 U561 ( .A(n741), .ZN(n141) );
  AOI22_X1 U562 ( .A1(addr_a2[4]), .A2(n75), .B1(N109), .B2(n742), .ZN(n741)
         );
  INV_X1 U563 ( .A(n484), .ZN(n117) );
  AOI22_X1 U564 ( .A1(addr_y[4]), .A2(n485), .B1(N587), .B2(n119), .ZN(n484)
         );
  INV_X1 U565 ( .A(n712), .ZN(n246) );
  AOI22_X1 U566 ( .A1(addr_a6[2]), .A2(n70), .B1(N167), .B2(n710), .ZN(n712)
         );
  INV_X1 U567 ( .A(n685), .ZN(n251) );
  AOI22_X1 U568 ( .A1(addr_a9[2]), .A2(n74), .B1(N212), .B2(n683), .ZN(n685)
         );
  INV_X1 U569 ( .A(n676), .ZN(n256) );
  AOI22_X1 U570 ( .A1(addr_a10[2]), .A2(n74), .B1(N227), .B2(n674), .ZN(n676)
         );
  INV_X1 U571 ( .A(n660), .ZN(n261) );
  AOI22_X1 U572 ( .A1(addr_a12[2]), .A2(n74), .B1(N257), .B2(n658), .ZN(n660)
         );
  INV_X1 U573 ( .A(n668), .ZN(n266) );
  AOI22_X1 U574 ( .A1(addr_a11[2]), .A2(n71), .B1(N242), .B2(n666), .ZN(n668)
         );
  INV_X1 U575 ( .A(n693), .ZN(n271) );
  AOI22_X1 U576 ( .A1(addr_a8[2]), .A2(n71), .B1(N197), .B2(n691), .ZN(n693)
         );
  INV_X1 U577 ( .A(n702), .ZN(n276) );
  AOI22_X1 U578 ( .A1(addr_a7[2]), .A2(n73), .B1(N182), .B2(n700), .ZN(n702)
         );
  INV_X1 U579 ( .A(n513), .ZN(n124) );
  AOI22_X1 U580 ( .A1(addr_a30[2]), .A2(n70), .B1(N527), .B2(n511), .ZN(n513)
         );
  INV_X1 U581 ( .A(n727), .ZN(n235) );
  AOI22_X1 U582 ( .A1(addr_a4[2]), .A2(n75), .B1(N137), .B2(n725), .ZN(n727)
         );
  INV_X1 U583 ( .A(n547), .ZN(n199) );
  AOI22_X1 U584 ( .A1(addr_a26[2]), .A2(n72), .B1(N467), .B2(n545), .ZN(n547)
         );
  INV_X1 U585 ( .A(n530), .ZN(n204) );
  AOI22_X1 U586 ( .A1(addr_a28[2]), .A2(n70), .B1(N497), .B2(n528), .ZN(n530)
         );
  INV_X1 U587 ( .A(n561), .ZN(n209) );
  AOI22_X1 U588 ( .A1(addr_a24[2]), .A2(n72), .B1(N437), .B2(n559), .ZN(n561)
         );
  INV_X1 U589 ( .A(n538), .ZN(n214) );
  AOI22_X1 U590 ( .A1(addr_a27[2]), .A2(n75), .B1(N482), .B2(n536), .ZN(n538)
         );
  INV_X1 U591 ( .A(n636), .ZN(n164) );
  AOI22_X1 U592 ( .A1(addr_a15[2]), .A2(n74), .B1(N302), .B2(n634), .ZN(n636)
         );
  INV_X1 U593 ( .A(n628), .ZN(n169) );
  AOI22_X1 U594 ( .A1(addr_a16[2]), .A2(n71), .B1(N317), .B2(n626), .ZN(n628)
         );
  INV_X1 U595 ( .A(n618), .ZN(n174) );
  AOI22_X1 U596 ( .A1(addr_a17[2]), .A2(n74), .B1(N332), .B2(n616), .ZN(n618)
         );
  INV_X1 U597 ( .A(n644), .ZN(n159) );
  AOI22_X1 U598 ( .A1(addr_a14[2]), .A2(n411), .B1(N287), .B2(n642), .ZN(n644)
         );
  INV_X1 U599 ( .A(n610), .ZN(n144) );
  AOI22_X1 U600 ( .A1(addr_a18[2]), .A2(n70), .B1(N347), .B2(n608), .ZN(n610)
         );
  INV_X1 U601 ( .A(n602), .ZN(n154) );
  AOI22_X1 U602 ( .A1(addr_a19[2]), .A2(n411), .B1(N362), .B2(n600), .ZN(n602)
         );
  INV_X1 U603 ( .A(n594), .ZN(n149) );
  AOI22_X1 U604 ( .A1(addr_a20[2]), .A2(n74), .B1(N377), .B2(n592), .ZN(n594)
         );
  INV_X1 U605 ( .A(n719), .ZN(n240) );
  AOI22_X1 U606 ( .A1(addr_a5[2]), .A2(n74), .B1(N152), .B2(n717), .ZN(n719)
         );
  AND2_X1 U607 ( .A1(N573), .A2(n494), .ZN(N578) );
  INV_X1 U608 ( .A(n488), .ZN(n114) );
  AOI22_X1 U609 ( .A1(addr_y[1]), .A2(n485), .B1(N584), .B2(n119), .ZN(n488)
         );
  INV_X1 U610 ( .A(n713), .ZN(n245) );
  AOI22_X1 U611 ( .A1(addr_a6[1]), .A2(n71), .B1(N166), .B2(n710), .ZN(n713)
         );
  INV_X1 U612 ( .A(n686), .ZN(n250) );
  AOI22_X1 U613 ( .A1(addr_a9[1]), .A2(n72), .B1(N211), .B2(n683), .ZN(n686)
         );
  INV_X1 U614 ( .A(n677), .ZN(n255) );
  AOI22_X1 U615 ( .A1(addr_a10[1]), .A2(n72), .B1(N226), .B2(n674), .ZN(n677)
         );
  INV_X1 U616 ( .A(n661), .ZN(n260) );
  AOI22_X1 U617 ( .A1(addr_a12[1]), .A2(n73), .B1(N256), .B2(n658), .ZN(n661)
         );
  INV_X1 U618 ( .A(n669), .ZN(n265) );
  AOI22_X1 U619 ( .A1(addr_a11[1]), .A2(n70), .B1(N241), .B2(n666), .ZN(n669)
         );
  INV_X1 U620 ( .A(n694), .ZN(n270) );
  AOI22_X1 U621 ( .A1(addr_a8[1]), .A2(n411), .B1(N196), .B2(n691), .ZN(n694)
         );
  INV_X1 U622 ( .A(n703), .ZN(n275) );
  AOI22_X1 U623 ( .A1(addr_a7[1]), .A2(n72), .B1(N181), .B2(n700), .ZN(n703)
         );
  INV_X1 U624 ( .A(n514), .ZN(n123) );
  AOI22_X1 U625 ( .A1(addr_a30[1]), .A2(n75), .B1(N526), .B2(n511), .ZN(n514)
         );
  INV_X1 U626 ( .A(n728), .ZN(n234) );
  AOI22_X1 U627 ( .A1(addr_a4[1]), .A2(n75), .B1(N136), .B2(n725), .ZN(n728)
         );
  INV_X1 U628 ( .A(n548), .ZN(n198) );
  AOI22_X1 U629 ( .A1(addr_a26[1]), .A2(n72), .B1(N466), .B2(n545), .ZN(n548)
         );
  INV_X1 U630 ( .A(n531), .ZN(n203) );
  AOI22_X1 U631 ( .A1(addr_a28[1]), .A2(n70), .B1(N496), .B2(n528), .ZN(n531)
         );
  INV_X1 U632 ( .A(n562), .ZN(n208) );
  AOI22_X1 U633 ( .A1(addr_a24[1]), .A2(n73), .B1(N436), .B2(n559), .ZN(n562)
         );
  INV_X1 U634 ( .A(n539), .ZN(n213) );
  AOI22_X1 U635 ( .A1(addr_a27[1]), .A2(n70), .B1(N481), .B2(n536), .ZN(n539)
         );
  INV_X1 U636 ( .A(n637), .ZN(n163) );
  AOI22_X1 U637 ( .A1(addr_a15[1]), .A2(n411), .B1(N301), .B2(n634), .ZN(n637)
         );
  INV_X1 U638 ( .A(n629), .ZN(n168) );
  AOI22_X1 U639 ( .A1(addr_a16[1]), .A2(n74), .B1(N316), .B2(n626), .ZN(n629)
         );
  INV_X1 U640 ( .A(n619), .ZN(n173) );
  AOI22_X1 U641 ( .A1(addr_a17[1]), .A2(n74), .B1(N331), .B2(n616), .ZN(n619)
         );
  INV_X1 U642 ( .A(n645), .ZN(n158) );
  AOI22_X1 U643 ( .A1(addr_a14[1]), .A2(n72), .B1(N286), .B2(n642), .ZN(n645)
         );
  INV_X1 U644 ( .A(n611), .ZN(n143) );
  AOI22_X1 U645 ( .A1(addr_a18[1]), .A2(n71), .B1(N346), .B2(n608), .ZN(n611)
         );
  INV_X1 U646 ( .A(n603), .ZN(n153) );
  AOI22_X1 U647 ( .A1(addr_a19[1]), .A2(n411), .B1(N361), .B2(n600), .ZN(n603)
         );
  INV_X1 U648 ( .A(n595), .ZN(n148) );
  AOI22_X1 U649 ( .A1(addr_a20[1]), .A2(n74), .B1(N376), .B2(n592), .ZN(n595)
         );
  INV_X1 U650 ( .A(n720), .ZN(n239) );
  AOI22_X1 U651 ( .A1(addr_a5[1]), .A2(n411), .B1(N151), .B2(n717), .ZN(n720)
         );
  INV_X1 U652 ( .A(n487), .ZN(n115) );
  AOI22_X1 U653 ( .A1(addr_y[2]), .A2(n485), .B1(N585), .B2(n119), .ZN(n487)
         );
  INV_X1 U654 ( .A(n486), .ZN(n116) );
  AOI22_X1 U655 ( .A1(addr_y[3]), .A2(n485), .B1(N586), .B2(n119), .ZN(n486)
         );
  OAI22_X1 U656 ( .A1(n308), .A2(n481), .B1(n482), .B2(n483), .ZN(N596) );
  NAND2_X1 U657 ( .A1(n360), .A2(n358), .ZN(n483) );
  OR4_X1 U658 ( .A1(n435), .A2(loadMatrix), .A3(loadVector), .A4(start), .ZN(
        n434) );
  CLKBUF_X1 U659 ( .A(n70), .Z(n76) );
  XOR2_X1 U660 ( .A(\add_206/carry[4] ), .B(addr_a1[4]), .Z(N94) );
  XOR2_X1 U661 ( .A(\add_215/carry[4] ), .B(addr_a2[4]), .Z(N109) );
  XOR2_X1 U662 ( .A(\add_224/carry[4] ), .B(addr_a3[4]), .Z(N124) );
  XOR2_X1 U663 ( .A(\add_233/carry[4] ), .B(addr_a4[4]), .Z(N139) );
  XOR2_X1 U664 ( .A(\add_242/carry[4] ), .B(addr_a5[4]), .Z(N154) );
  XOR2_X1 U665 ( .A(\add_251/carry[4] ), .B(addr_a6[4]), .Z(N169) );
  XOR2_X1 U666 ( .A(\add_260/carry[4] ), .B(addr_a7[4]), .Z(N184) );
  XOR2_X1 U667 ( .A(\add_269/carry[4] ), .B(addr_a8[4]), .Z(N199) );
  XOR2_X1 U668 ( .A(\add_278/carry[4] ), .B(addr_a9[4]), .Z(N214) );
  XOR2_X1 U669 ( .A(\add_287/carry[4] ), .B(addr_a10[4]), .Z(N229) );
  XOR2_X1 U670 ( .A(\add_296/carry[4] ), .B(addr_a11[4]), .Z(N244) );
  XOR2_X1 U671 ( .A(\add_305/carry[4] ), .B(addr_a12[4]), .Z(N259) );
  XOR2_X1 U672 ( .A(\add_314/carry[4] ), .B(addr_a13[4]), .Z(N274) );
  XOR2_X1 U673 ( .A(\add_323/carry[4] ), .B(addr_a14[4]), .Z(N289) );
  XOR2_X1 U674 ( .A(\add_332/carry[4] ), .B(addr_a15[4]), .Z(N304) );
  XOR2_X1 U675 ( .A(\add_341/carry[4] ), .B(addr_a16[4]), .Z(N319) );
  XOR2_X1 U676 ( .A(\add_350/carry[4] ), .B(addr_a17[4]), .Z(N334) );
  XOR2_X1 U677 ( .A(\add_359/carry[4] ), .B(addr_a18[4]), .Z(N349) );
  XOR2_X1 U678 ( .A(\add_368/carry[4] ), .B(addr_a19[4]), .Z(N364) );
  XOR2_X1 U679 ( .A(\add_377/carry[4] ), .B(addr_a20[4]), .Z(N379) );
  XOR2_X1 U680 ( .A(\add_386/carry[4] ), .B(addr_a21[4]), .Z(N394) );
  XOR2_X1 U681 ( .A(\add_395/carry[4] ), .B(addr_a22[4]), .Z(N409) );
  XOR2_X1 U682 ( .A(\add_404/carry[4] ), .B(addr_a23[4]), .Z(N424) );
  XOR2_X1 U683 ( .A(\add_413/carry[4] ), .B(addr_a24[4]), .Z(N439) );
  XOR2_X1 U684 ( .A(\add_422/carry[4] ), .B(addr_a25[4]), .Z(N454) );
  XOR2_X1 U685 ( .A(\add_431/carry[4] ), .B(addr_a26[4]), .Z(N469) );
  XOR2_X1 U686 ( .A(\add_440/carry[4] ), .B(addr_a27[4]), .Z(N484) );
  XOR2_X1 U687 ( .A(\add_449/carry[4] ), .B(addr_a28[4]), .Z(N499) );
  XOR2_X1 U688 ( .A(\add_458/carry[4] ), .B(addr_a29[4]), .Z(N514) );
  XOR2_X1 U689 ( .A(\add_467/carry[4] ), .B(addr_a30[4]), .Z(N529) );
  XOR2_X1 U690 ( .A(\add_476/carry[4] ), .B(addr_a31[4]), .Z(N544) );
  XOR2_X1 U691 ( .A(\add_485/carry[4] ), .B(addr_a32[4]), .Z(N559) );
  XOR2_X1 U692 ( .A(\add_494/carry[4] ), .B(addr_x[4]), .Z(N573) );
  XOR2_X1 U693 ( .A(\add_501/carry[4] ), .B(addr_y[4]), .Z(N587) );
  AND2_X1 U694 ( .A1(addr_x[1]), .A2(addr_x[0]), .ZN(n77) );
  NAND4_X1 U695 ( .A1(addr_x[4]), .A2(addr_x[3]), .A3(n77), .A4(addr_x[2]), 
        .ZN(N668) );
  AND2_X1 U696 ( .A1(addr_y[1]), .A2(addr_y[0]), .ZN(n78) );
  NAND4_X1 U697 ( .A1(addr_y[4]), .A2(addr_y[3]), .A3(n78), .A4(addr_y[2]), 
        .ZN(N674) );
  AND2_X1 U698 ( .A1(addr_a1[1]), .A2(addr_a1[0]), .ZN(n79) );
  NAND4_X1 U699 ( .A1(addr_a1[4]), .A2(addr_a1[3]), .A3(n79), .A4(addr_a1[2]), 
        .ZN(N604) );
  AND2_X1 U700 ( .A1(addr_a2[1]), .A2(addr_a2[0]), .ZN(n80) );
  NAND4_X1 U701 ( .A1(addr_a2[4]), .A2(addr_a2[3]), .A3(n80), .A4(addr_a2[2]), 
        .ZN(N606) );
  AND2_X1 U702 ( .A1(addr_a3[1]), .A2(addr_a3[0]), .ZN(n81) );
  NAND4_X1 U703 ( .A1(addr_a3[4]), .A2(addr_a3[3]), .A3(n81), .A4(addr_a3[2]), 
        .ZN(N608) );
  AND2_X1 U704 ( .A1(addr_a4[1]), .A2(addr_a4[0]), .ZN(n82) );
  NAND4_X1 U705 ( .A1(addr_a4[4]), .A2(addr_a4[3]), .A3(n82), .A4(addr_a4[2]), 
        .ZN(N610) );
  AND2_X1 U706 ( .A1(addr_a5[1]), .A2(addr_a5[0]), .ZN(n83) );
  NAND4_X1 U707 ( .A1(addr_a5[4]), .A2(addr_a5[3]), .A3(n83), .A4(addr_a5[2]), 
        .ZN(N612) );
  AND2_X1 U708 ( .A1(addr_a6[1]), .A2(addr_a6[0]), .ZN(n84) );
  NAND4_X1 U709 ( .A1(addr_a6[4]), .A2(addr_a6[3]), .A3(n84), .A4(addr_a6[2]), 
        .ZN(N614) );
  AND2_X1 U710 ( .A1(addr_a7[1]), .A2(addr_a7[0]), .ZN(n85) );
  NAND4_X1 U711 ( .A1(addr_a7[4]), .A2(addr_a7[3]), .A3(n85), .A4(addr_a7[2]), 
        .ZN(N616) );
  AND2_X1 U712 ( .A1(addr_a8[1]), .A2(addr_a8[0]), .ZN(n86) );
  NAND4_X1 U713 ( .A1(addr_a8[4]), .A2(addr_a8[3]), .A3(n86), .A4(addr_a8[2]), 
        .ZN(N618) );
  AND2_X1 U714 ( .A1(addr_a9[1]), .A2(addr_a9[0]), .ZN(n87) );
  NAND4_X1 U715 ( .A1(addr_a9[4]), .A2(addr_a9[3]), .A3(n87), .A4(addr_a9[2]), 
        .ZN(N620) );
  AND2_X1 U716 ( .A1(addr_a10[1]), .A2(addr_a10[0]), .ZN(n88) );
  NAND4_X1 U717 ( .A1(addr_a10[4]), .A2(addr_a10[3]), .A3(n88), .A4(
        addr_a10[2]), .ZN(N622) );
  AND2_X1 U718 ( .A1(addr_a11[1]), .A2(addr_a11[0]), .ZN(n89) );
  NAND4_X1 U719 ( .A1(addr_a11[4]), .A2(addr_a11[3]), .A3(n89), .A4(
        addr_a11[2]), .ZN(N624) );
  AND2_X1 U747 ( .A1(addr_a12[1]), .A2(addr_a12[0]), .ZN(n90) );
  NAND4_X1 U748 ( .A1(addr_a12[4]), .A2(addr_a12[3]), .A3(n90), .A4(
        addr_a12[2]), .ZN(N626) );
  AND2_X1 U749 ( .A1(addr_a13[1]), .A2(addr_a13[0]), .ZN(n91) );
  NAND4_X1 U750 ( .A1(addr_a13[4]), .A2(addr_a13[3]), .A3(n91), .A4(
        addr_a13[2]), .ZN(N628) );
  AND2_X1 U751 ( .A1(addr_a14[1]), .A2(addr_a14[0]), .ZN(n92) );
  NAND4_X1 U752 ( .A1(addr_a14[4]), .A2(addr_a14[3]), .A3(n92), .A4(
        addr_a14[2]), .ZN(N630) );
  AND2_X1 U753 ( .A1(addr_a15[1]), .A2(addr_a15[0]), .ZN(n93) );
  NAND4_X1 U754 ( .A1(addr_a15[4]), .A2(addr_a15[3]), .A3(n93), .A4(
        addr_a15[2]), .ZN(N632) );
  AND2_X1 U755 ( .A1(addr_a16[1]), .A2(addr_a16[0]), .ZN(n94) );
  NAND4_X1 U756 ( .A1(addr_a16[4]), .A2(addr_a16[3]), .A3(n94), .A4(
        addr_a16[2]), .ZN(N634) );
  AND2_X1 U757 ( .A1(addr_a17[1]), .A2(addr_a17[0]), .ZN(n95) );
  NAND4_X1 U758 ( .A1(addr_a17[4]), .A2(addr_a17[3]), .A3(n95), .A4(
        addr_a17[2]), .ZN(N636) );
  AND2_X1 U759 ( .A1(addr_a18[1]), .A2(addr_a18[0]), .ZN(n96) );
  NAND4_X1 U760 ( .A1(addr_a18[4]), .A2(addr_a18[3]), .A3(n96), .A4(
        addr_a18[2]), .ZN(N638) );
  AND2_X1 U761 ( .A1(addr_a19[1]), .A2(addr_a19[0]), .ZN(n97) );
  NAND4_X1 U762 ( .A1(addr_a19[4]), .A2(addr_a19[3]), .A3(n97), .A4(
        addr_a19[2]), .ZN(N640) );
  AND2_X1 U763 ( .A1(addr_a20[1]), .A2(addr_a20[0]), .ZN(n98) );
  NAND4_X1 U764 ( .A1(addr_a20[4]), .A2(addr_a20[3]), .A3(n98), .A4(
        addr_a20[2]), .ZN(N642) );
  AND2_X1 U765 ( .A1(addr_a21[1]), .A2(addr_a21[0]), .ZN(n99) );
  NAND4_X1 U766 ( .A1(addr_a21[4]), .A2(addr_a21[3]), .A3(n99), .A4(
        addr_a21[2]), .ZN(N644) );
  AND2_X1 U767 ( .A1(addr_a22[1]), .A2(addr_a22[0]), .ZN(n100) );
  NAND4_X1 U768 ( .A1(addr_a22[4]), .A2(addr_a22[3]), .A3(n100), .A4(
        addr_a22[2]), .ZN(N646) );
  AND2_X1 U769 ( .A1(addr_a23[1]), .A2(addr_a23[0]), .ZN(n101) );
  NAND4_X1 U770 ( .A1(addr_a23[4]), .A2(addr_a23[3]), .A3(n101), .A4(
        addr_a23[2]), .ZN(N648) );
  AND2_X1 U771 ( .A1(addr_a24[1]), .A2(addr_a24[0]), .ZN(n102) );
  NAND4_X1 U772 ( .A1(addr_a24[4]), .A2(addr_a24[3]), .A3(n102), .A4(
        addr_a24[2]), .ZN(N650) );
  AND2_X1 U773 ( .A1(addr_a25[1]), .A2(addr_a25[0]), .ZN(n103) );
  NAND4_X1 U774 ( .A1(addr_a25[4]), .A2(addr_a25[3]), .A3(n103), .A4(
        addr_a25[2]), .ZN(N652) );
  AND2_X1 U775 ( .A1(addr_a26[1]), .A2(addr_a26[0]), .ZN(n104) );
  NAND4_X1 U776 ( .A1(addr_a26[4]), .A2(addr_a26[3]), .A3(n104), .A4(
        addr_a26[2]), .ZN(N654) );
  AND2_X1 U777 ( .A1(addr_a27[1]), .A2(addr_a27[0]), .ZN(n105) );
  NAND4_X1 U778 ( .A1(addr_a27[4]), .A2(addr_a27[3]), .A3(n105), .A4(
        addr_a27[2]), .ZN(N656) );
  AND2_X1 U779 ( .A1(addr_a28[1]), .A2(addr_a28[0]), .ZN(n106) );
  NAND4_X1 U780 ( .A1(addr_a28[4]), .A2(addr_a28[3]), .A3(n106), .A4(
        addr_a28[2]), .ZN(N658) );
  AND2_X1 U781 ( .A1(addr_a29[1]), .A2(addr_a29[0]), .ZN(n107) );
  NAND4_X1 U782 ( .A1(addr_a29[4]), .A2(addr_a29[3]), .A3(n107), .A4(
        addr_a29[2]), .ZN(N660) );
  AND2_X1 U783 ( .A1(addr_a30[1]), .A2(addr_a30[0]), .ZN(n108) );
  NAND4_X1 U784 ( .A1(addr_a30[4]), .A2(addr_a30[3]), .A3(n108), .A4(
        addr_a30[2]), .ZN(N662) );
  AND2_X1 U785 ( .A1(addr_a31[1]), .A2(addr_a31[0]), .ZN(n109) );
  NAND4_X1 U786 ( .A1(addr_a31[4]), .A2(addr_a31[3]), .A3(n109), .A4(
        addr_a31[2]), .ZN(N664) );
  AND2_X1 U787 ( .A1(addr_a32[1]), .A2(addr_a32[0]), .ZN(n110) );
  NAND4_X1 U788 ( .A1(addr_a32[4]), .A2(addr_a32[3]), .A3(n110), .A4(
        addr_a32[2]), .ZN(N666) );
endmodule


module mvm_32_32_8_1 ( clk, reset, loadMatrix, loadVector, start, done, 
        data_in, data_out );
  input [7:0] data_in;
  output [15:0] data_out;
  input clk, reset, loadMatrix, loadVector, start;
  output done;
  wire   wr_en_x, wr_en_a1, wr_en_a2, wr_en_a3, wr_en_a4, wr_en_a5, wr_en_a6,
         wr_en_a7, wr_en_a8, wr_en_a9, wr_en_a10, wr_en_a11, wr_en_a12,
         wr_en_a13, wr_en_a14, wr_en_a15, wr_en_a16, wr_en_a17, wr_en_a18,
         wr_en_a19, wr_en_a20, wr_en_a21, wr_en_a22, wr_en_a23, wr_en_a24,
         wr_en_a25, wr_en_a26, wr_en_a27, wr_en_a28, wr_en_a29, wr_en_a30,
         wr_en_a31, wr_en_a32, wr_en_y, clear_acc, clc, clc1;
  wire   [4:0] addr_x;
  wire   [4:0] addr_a1;
  wire   [4:0] addr_a2;
  wire   [4:0] addr_a3;
  wire   [4:0] addr_a4;
  wire   [4:0] addr_a5;
  wire   [4:0] addr_a6;
  wire   [4:0] addr_a7;
  wire   [4:0] addr_a8;
  wire   [4:0] addr_a9;
  wire   [4:0] addr_a10;
  wire   [4:0] addr_a11;
  wire   [4:0] addr_a12;
  wire   [4:0] addr_a13;
  wire   [4:0] addr_a14;
  wire   [4:0] addr_a15;
  wire   [4:0] addr_a16;
  wire   [4:0] addr_a17;
  wire   [4:0] addr_a18;
  wire   [4:0] addr_a19;
  wire   [4:0] addr_a20;
  wire   [4:0] addr_a21;
  wire   [4:0] addr_a22;
  wire   [4:0] addr_a23;
  wire   [4:0] addr_a24;
  wire   [4:0] addr_a25;
  wire   [4:0] addr_a26;
  wire   [4:0] addr_a27;
  wire   [4:0] addr_a28;
  wire   [4:0] addr_a29;
  wire   [4:0] addr_a30;
  wire   [4:0] addr_a31;
  wire   [4:0] addr_a32;
  wire   [4:0] addr_y;

  datapath d ( .clk(clk), .data_in(data_in), .addr_x(addr_x), .wr_en_x(wr_en_x), .addr_a1(addr_a1), .addr_a2(addr_a2), .addr_a3(addr_a3), .addr_a4(addr_a4), 
        .addr_a5(addr_a5), .addr_a6(addr_a6), .addr_a7(addr_a7), .addr_a8(
        addr_a8), .addr_a9(addr_a9), .addr_a10(addr_a10), .addr_a11(addr_a11), 
        .addr_a12(addr_a12), .addr_a13(addr_a13), .addr_a14(addr_a14), 
        .addr_a15(addr_a15), .addr_a16(addr_a16), .addr_a17(addr_a17), 
        .addr_a18(addr_a18), .addr_a19(addr_a19), .addr_a20(addr_a20), 
        .addr_a21(addr_a21), .addr_a22(addr_a22), .addr_a23(addr_a23), 
        .addr_a24(addr_a24), .addr_a25(addr_a25), .addr_a26(addr_a26), 
        .addr_a27(addr_a27), .addr_a28(addr_a28), .addr_a29(addr_a29), 
        .addr_a30(addr_a30), .addr_a31(addr_a31), .addr_a32(addr_a32), 
        .wr_en_a1(wr_en_a1), .wr_en_a2(wr_en_a2), .wr_en_a3(wr_en_a3), 
        .wr_en_a4(wr_en_a4), .wr_en_a5(wr_en_a5), .wr_en_a6(wr_en_a6), 
        .wr_en_a7(wr_en_a7), .wr_en_a8(wr_en_a8), .wr_en_a9(wr_en_a9), 
        .wr_en_a10(wr_en_a10), .wr_en_a11(wr_en_a11), .wr_en_a12(wr_en_a12), 
        .wr_en_a13(wr_en_a13), .wr_en_a14(wr_en_a14), .wr_en_a15(wr_en_a15), 
        .wr_en_a16(wr_en_a16), .wr_en_a17(wr_en_a17), .wr_en_a18(wr_en_a18), 
        .wr_en_a19(wr_en_a19), .wr_en_a20(wr_en_a20), .wr_en_a21(wr_en_a21), 
        .wr_en_a22(wr_en_a22), .wr_en_a23(wr_en_a23), .wr_en_a24(wr_en_a24), 
        .wr_en_a25(wr_en_a25), .wr_en_a26(wr_en_a26), .wr_en_a27(wr_en_a27), 
        .wr_en_a28(wr_en_a28), .wr_en_a29(wr_en_a29), .wr_en_a30(wr_en_a30), 
        .wr_en_a31(wr_en_a31), .wr_en_a32(wr_en_a32), .addr_y(addr_y), 
        .wr_en_y(wr_en_y), .clear_acc(clear_acc), .clc(clc), .clc1(clc1), 
        .data_out(data_out) );
  ctrlpath c ( .clk(clk), .reset(reset), .start(start), .addr_x(addr_x), 
        .wr_en_x(wr_en_x), .addr_a1(addr_a1), .addr_a2(addr_a2), .addr_a3(
        addr_a3), .addr_a4(addr_a4), .addr_a5(addr_a5), .addr_a6(addr_a6), 
        .addr_a7(addr_a7), .addr_a8(addr_a8), .addr_a9(addr_a9), .addr_a10(
        addr_a10), .addr_a11(addr_a11), .addr_a12(addr_a12), .addr_a13(
        addr_a13), .addr_a14(addr_a14), .addr_a15(addr_a15), .addr_a16(
        addr_a16), .addr_a17(addr_a17), .addr_a18(addr_a18), .addr_a19(
        addr_a19), .addr_a20(addr_a20), .addr_a21(addr_a21), .addr_a22(
        addr_a22), .addr_a23(addr_a23), .addr_a24(addr_a24), .addr_a25(
        addr_a25), .addr_a26(addr_a26), .addr_a27(addr_a27), .addr_a28(
        addr_a28), .addr_a29(addr_a29), .addr_a30(addr_a30), .addr_a31(
        addr_a31), .addr_a32(addr_a32), .wr_en_a1(wr_en_a1), .wr_en_a2(
        wr_en_a2), .wr_en_a3(wr_en_a3), .wr_en_a4(wr_en_a4), .wr_en_a5(
        wr_en_a5), .wr_en_a6(wr_en_a6), .wr_en_a7(wr_en_a7), .wr_en_a8(
        wr_en_a8), .wr_en_a9(wr_en_a9), .wr_en_a10(wr_en_a10), .wr_en_a11(
        wr_en_a11), .wr_en_a12(wr_en_a12), .wr_en_a13(wr_en_a13), .wr_en_a14(
        wr_en_a14), .wr_en_a15(wr_en_a15), .wr_en_a16(wr_en_a16), .wr_en_a17(
        wr_en_a17), .wr_en_a18(wr_en_a18), .wr_en_a19(wr_en_a19), .wr_en_a20(
        wr_en_a20), .wr_en_a21(wr_en_a21), .wr_en_a22(wr_en_a22), .wr_en_a23(
        wr_en_a23), .wr_en_a24(wr_en_a24), .wr_en_a25(wr_en_a25), .wr_en_a26(
        wr_en_a26), .wr_en_a27(wr_en_a27), .wr_en_a28(wr_en_a28), .wr_en_a29(
        wr_en_a29), .wr_en_a30(wr_en_a30), .wr_en_a31(wr_en_a31), .wr_en_a32(
        wr_en_a32), .clear_acc(clear_acc), .clc(clc), .clc1(clc1), .addr_y(
        addr_y), .wr_en_y(wr_en_y), .done(done), .loadMatrix(loadMatrix), 
        .loadVector(loadVector) );
endmodule

